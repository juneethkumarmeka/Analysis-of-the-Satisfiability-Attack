module basic_2000_20000_2500_4_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_106,In_1636);
xor U1 (N_1,In_1199,In_651);
nor U2 (N_2,In_420,In_358);
and U3 (N_3,In_1723,In_425);
nand U4 (N_4,In_245,In_179);
or U5 (N_5,In_599,In_1255);
xor U6 (N_6,In_923,In_399);
and U7 (N_7,In_491,In_1050);
or U8 (N_8,In_950,In_926);
and U9 (N_9,In_1475,In_240);
or U10 (N_10,In_828,In_474);
and U11 (N_11,In_521,In_1813);
or U12 (N_12,In_1566,In_1720);
or U13 (N_13,In_137,In_1510);
nor U14 (N_14,In_843,In_1184);
nand U15 (N_15,In_1450,In_708);
nand U16 (N_16,In_91,In_1150);
nor U17 (N_17,In_1030,In_647);
or U18 (N_18,In_1552,In_1954);
or U19 (N_19,In_263,In_1346);
and U20 (N_20,In_753,In_359);
and U21 (N_21,In_1920,In_1085);
and U22 (N_22,In_682,In_1539);
nand U23 (N_23,In_104,In_1138);
nand U24 (N_24,In_951,In_1489);
nand U25 (N_25,In_1296,In_173);
xor U26 (N_26,In_204,In_591);
or U27 (N_27,In_1998,In_47);
nand U28 (N_28,In_1188,In_631);
nor U29 (N_29,In_1322,In_1559);
or U30 (N_30,In_1575,In_1758);
nand U31 (N_31,In_95,In_1205);
or U32 (N_32,In_1187,In_1598);
or U33 (N_33,In_1061,In_52);
and U34 (N_34,In_1816,In_1573);
or U35 (N_35,In_632,In_852);
nand U36 (N_36,In_1166,In_900);
or U37 (N_37,In_219,In_449);
nor U38 (N_38,In_601,In_1502);
or U39 (N_39,In_692,In_1135);
and U40 (N_40,In_54,In_954);
nor U41 (N_41,In_1049,In_987);
and U42 (N_42,In_927,In_341);
nand U43 (N_43,In_518,In_360);
and U44 (N_44,In_1057,In_1206);
or U45 (N_45,In_1756,In_1499);
nor U46 (N_46,In_70,In_571);
or U47 (N_47,In_198,In_1417);
and U48 (N_48,In_1679,In_1970);
or U49 (N_49,In_1807,In_1103);
and U50 (N_50,In_1655,In_1618);
or U51 (N_51,In_1545,In_853);
nand U52 (N_52,In_93,In_1880);
nor U53 (N_53,In_654,In_1314);
nand U54 (N_54,In_1226,In_1044);
or U55 (N_55,In_722,In_635);
nor U56 (N_56,In_1121,In_959);
nor U57 (N_57,In_11,In_803);
and U58 (N_58,In_97,In_344);
and U59 (N_59,In_423,In_439);
nor U60 (N_60,In_1113,In_533);
nand U61 (N_61,In_1752,In_1143);
or U62 (N_62,In_740,In_1481);
or U63 (N_63,In_1436,In_1717);
nand U64 (N_64,In_1520,In_880);
nor U65 (N_65,In_250,In_1691);
nor U66 (N_66,In_1458,In_300);
and U67 (N_67,In_442,In_98);
or U68 (N_68,In_1556,In_1656);
nand U69 (N_69,In_662,In_1392);
and U70 (N_70,In_258,In_897);
nand U71 (N_71,In_226,In_553);
nor U72 (N_72,In_1038,In_924);
nor U73 (N_73,In_484,In_977);
nor U74 (N_74,In_731,In_408);
nand U75 (N_75,In_166,In_1531);
nor U76 (N_76,In_225,In_62);
nor U77 (N_77,In_319,In_1710);
or U78 (N_78,In_638,In_1628);
and U79 (N_79,In_574,In_1214);
nor U80 (N_80,In_1411,In_373);
or U81 (N_81,In_383,In_1385);
and U82 (N_82,In_1240,In_279);
and U83 (N_83,In_535,In_497);
and U84 (N_84,In_1682,In_1429);
nor U85 (N_85,In_809,In_906);
nand U86 (N_86,In_693,In_1785);
or U87 (N_87,In_1796,In_770);
and U88 (N_88,In_794,In_1620);
nor U89 (N_89,In_308,In_89);
or U90 (N_90,In_560,In_808);
nor U91 (N_91,In_1939,In_1021);
nand U92 (N_92,In_610,In_515);
nor U93 (N_93,In_1399,In_1662);
and U94 (N_94,In_548,In_832);
nand U95 (N_95,In_134,In_694);
nand U96 (N_96,In_1716,In_1955);
or U97 (N_97,In_278,In_63);
and U98 (N_98,In_1344,In_288);
and U99 (N_99,In_1151,In_1430);
xnor U100 (N_100,In_757,In_685);
and U101 (N_101,In_1276,In_1607);
nand U102 (N_102,In_277,In_1200);
and U103 (N_103,In_846,In_939);
nor U104 (N_104,In_86,In_1791);
nor U105 (N_105,In_435,In_1553);
or U106 (N_106,In_1833,In_1039);
nand U107 (N_107,In_1705,In_626);
nor U108 (N_108,In_642,In_686);
nor U109 (N_109,In_144,In_71);
or U110 (N_110,In_320,In_1660);
nand U111 (N_111,In_778,In_1515);
nor U112 (N_112,In_816,In_1830);
nor U113 (N_113,In_1068,In_1852);
or U114 (N_114,In_1605,In_716);
and U115 (N_115,In_1145,In_139);
and U116 (N_116,In_588,In_1459);
nand U117 (N_117,In_130,In_1357);
and U118 (N_118,In_1086,In_863);
nor U119 (N_119,In_337,In_266);
or U120 (N_120,In_1131,In_1674);
or U121 (N_121,In_94,In_490);
nand U122 (N_122,In_1882,In_1183);
nand U123 (N_123,In_1104,In_909);
nor U124 (N_124,In_1002,In_671);
or U125 (N_125,In_721,In_646);
or U126 (N_126,In_371,In_100);
and U127 (N_127,In_1786,In_176);
nor U128 (N_128,In_958,In_103);
nor U129 (N_129,In_121,In_1944);
nor U130 (N_130,In_1555,In_568);
nand U131 (N_131,In_46,In_232);
nor U132 (N_132,In_1733,In_965);
nand U133 (N_133,In_325,In_1498);
or U134 (N_134,In_1164,In_1902);
nor U135 (N_135,In_1310,In_1161);
nor U136 (N_136,In_340,In_223);
nand U137 (N_137,In_1088,In_291);
or U138 (N_138,In_1697,In_723);
nand U139 (N_139,In_1087,In_554);
nor U140 (N_140,In_1870,In_613);
and U141 (N_141,In_1007,In_0);
and U142 (N_142,In_1117,In_164);
and U143 (N_143,In_1380,In_437);
nor U144 (N_144,In_1953,In_1141);
nand U145 (N_145,In_1378,In_339);
nand U146 (N_146,In_1529,In_516);
nor U147 (N_147,In_1316,In_1389);
nor U148 (N_148,In_573,In_1174);
or U149 (N_149,In_985,In_1129);
and U150 (N_150,In_1783,In_583);
nand U151 (N_151,In_1726,In_899);
nor U152 (N_152,In_962,In_1695);
or U153 (N_153,In_156,In_1744);
nand U154 (N_154,In_108,In_294);
or U155 (N_155,In_1988,In_877);
nor U156 (N_156,In_1198,In_1779);
nor U157 (N_157,In_921,In_1402);
and U158 (N_158,In_1915,In_1884);
or U159 (N_159,In_931,In_1926);
xnor U160 (N_160,In_1640,In_1275);
or U161 (N_161,In_189,In_650);
and U162 (N_162,In_23,In_1839);
nor U163 (N_163,In_1631,In_1362);
nand U164 (N_164,In_1290,In_868);
or U165 (N_165,In_760,In_1163);
or U166 (N_166,In_124,In_717);
or U167 (N_167,In_188,In_1425);
nor U168 (N_168,In_1672,In_318);
nand U169 (N_169,In_367,In_1751);
and U170 (N_170,In_656,In_1230);
or U171 (N_171,In_744,In_1175);
nand U172 (N_172,In_1757,In_1619);
nor U173 (N_173,In_1629,In_1702);
nor U174 (N_174,In_145,In_1949);
nor U175 (N_175,In_1587,In_1651);
or U176 (N_176,In_1196,In_1648);
or U177 (N_177,In_1516,In_504);
nor U178 (N_178,In_624,In_1806);
nand U179 (N_179,In_80,In_1537);
or U180 (N_180,In_305,In_1464);
nor U181 (N_181,In_180,In_1118);
or U182 (N_182,In_218,In_697);
nand U183 (N_183,In_1558,In_1601);
nor U184 (N_184,In_1673,In_32);
and U185 (N_185,In_1313,In_904);
xnor U186 (N_186,In_1860,In_57);
or U187 (N_187,In_202,In_274);
nor U188 (N_188,In_1147,In_1289);
or U189 (N_189,In_1112,In_1423);
and U190 (N_190,In_643,In_1202);
or U191 (N_191,In_1019,In_995);
xnor U192 (N_192,In_947,In_1484);
nor U193 (N_193,In_310,In_1937);
nand U194 (N_194,In_409,In_990);
or U195 (N_195,In_614,In_641);
nand U196 (N_196,In_881,In_1784);
nand U197 (N_197,In_454,In_737);
nand U198 (N_198,In_1259,In_1023);
nand U199 (N_199,In_823,In_764);
nand U200 (N_200,In_1773,In_1521);
nor U201 (N_201,In_860,In_256);
nand U202 (N_202,In_1356,In_384);
nand U203 (N_203,In_306,In_1480);
nor U204 (N_204,In_1031,In_1506);
or U205 (N_205,In_84,In_1795);
nor U206 (N_206,In_353,In_578);
nor U207 (N_207,In_1540,In_1476);
nor U208 (N_208,In_749,In_1060);
or U209 (N_209,In_658,In_1856);
nor U210 (N_210,In_1277,In_728);
and U211 (N_211,In_151,In_527);
and U212 (N_212,In_824,In_1445);
or U213 (N_213,In_1582,In_311);
and U214 (N_214,In_605,In_1438);
nor U215 (N_215,In_1868,In_679);
or U216 (N_216,In_856,In_362);
or U217 (N_217,In_798,In_1097);
nand U218 (N_218,In_249,In_1886);
and U219 (N_219,In_72,In_494);
nor U220 (N_220,In_627,In_1419);
and U221 (N_221,In_1251,In_1467);
nand U222 (N_222,In_1216,In_514);
or U223 (N_223,In_858,In_862);
and U224 (N_224,In_251,In_1070);
or U225 (N_225,In_1913,In_791);
or U226 (N_226,In_1133,In_968);
and U227 (N_227,In_35,In_1343);
or U228 (N_228,In_470,In_1584);
nand U229 (N_229,In_1832,In_855);
nor U230 (N_230,In_676,In_1272);
and U231 (N_231,In_467,In_175);
or U232 (N_232,In_1869,In_406);
nand U233 (N_233,In_1879,In_1471);
or U234 (N_234,In_1741,In_428);
nand U235 (N_235,In_471,In_257);
nand U236 (N_236,In_73,In_670);
or U237 (N_237,In_304,In_1659);
or U238 (N_238,In_1446,In_589);
nand U239 (N_239,In_1243,In_1986);
nor U240 (N_240,In_1534,In_620);
nand U241 (N_241,In_891,In_1286);
or U242 (N_242,In_1130,In_411);
and U243 (N_243,In_405,In_390);
nand U244 (N_244,In_133,In_1325);
nor U245 (N_245,In_1291,In_259);
or U246 (N_246,In_276,In_674);
or U247 (N_247,In_978,In_1114);
nand U248 (N_248,In_1212,In_640);
or U249 (N_249,In_532,In_530);
or U250 (N_250,In_7,In_1013);
nor U251 (N_251,In_562,In_1981);
nor U252 (N_252,In_413,In_1488);
nor U253 (N_253,In_612,In_1172);
or U254 (N_254,In_719,In_815);
nand U255 (N_255,In_243,In_1627);
xor U256 (N_256,In_40,In_1403);
or U257 (N_257,In_876,In_1678);
or U258 (N_258,In_349,In_1854);
or U259 (N_259,In_1606,In_1055);
and U260 (N_260,In_167,In_1509);
and U261 (N_261,In_368,In_505);
nand U262 (N_262,In_827,In_431);
nor U263 (N_263,In_1336,In_5);
nand U264 (N_264,In_1588,In_1689);
nor U265 (N_265,In_1638,In_1805);
nor U266 (N_266,In_1543,In_1765);
and U267 (N_267,In_922,In_1707);
nand U268 (N_268,In_338,In_769);
and U269 (N_269,In_508,In_865);
and U270 (N_270,In_168,In_919);
nor U271 (N_271,In_804,In_157);
and U272 (N_272,In_1302,In_512);
and U273 (N_273,In_236,In_460);
and U274 (N_274,In_285,In_31);
nand U275 (N_275,In_1401,In_1919);
nor U276 (N_276,In_1352,In_1787);
nand U277 (N_277,In_1195,In_1452);
or U278 (N_278,In_440,In_811);
nand U279 (N_279,In_109,In_988);
or U280 (N_280,In_1326,In_1661);
nor U281 (N_281,In_374,In_49);
nor U282 (N_282,In_1406,In_1728);
or U283 (N_283,In_476,In_1181);
or U284 (N_284,In_1080,In_1747);
and U285 (N_285,In_298,In_683);
and U286 (N_286,In_1797,In_25);
or U287 (N_287,In_1612,In_1461);
or U288 (N_288,In_607,In_1979);
nor U289 (N_289,In_659,In_487);
nor U290 (N_290,In_1846,In_1862);
or U291 (N_291,In_1084,In_1924);
nand U292 (N_292,In_1367,In_981);
or U293 (N_293,In_520,In_871);
or U294 (N_294,In_938,In_1692);
nor U295 (N_295,In_1664,In_1729);
nand U296 (N_296,In_1338,In_220);
nand U297 (N_297,In_443,In_1256);
and U298 (N_298,In_1665,In_1615);
or U299 (N_299,In_441,In_382);
nand U300 (N_300,In_1081,In_1447);
nor U301 (N_301,In_1825,In_1912);
nor U302 (N_302,In_1224,In_1448);
nand U303 (N_303,In_1867,In_943);
nor U304 (N_304,In_1646,In_265);
nand U305 (N_305,In_732,In_314);
nor U306 (N_306,In_1412,In_1761);
and U307 (N_307,In_81,In_892);
nand U308 (N_308,In_710,In_229);
or U309 (N_309,In_1091,In_970);
nor U310 (N_310,In_436,In_814);
and U311 (N_311,In_766,In_83);
nand U312 (N_312,In_639,In_1398);
nand U313 (N_313,In_112,In_864);
and U314 (N_314,In_765,In_172);
or U315 (N_315,In_1696,In_1887);
nor U316 (N_316,In_422,In_1693);
nand U317 (N_317,In_459,In_1388);
and U318 (N_318,In_1148,In_129);
nand U319 (N_319,In_247,In_1279);
nor U320 (N_320,In_1064,In_1273);
or U321 (N_321,In_1236,In_1991);
or U322 (N_322,In_1743,In_1951);
nor U323 (N_323,In_1822,In_1257);
nand U324 (N_324,In_1560,In_1153);
or U325 (N_325,In_1883,In_1144);
or U326 (N_326,In_569,In_1441);
nand U327 (N_327,In_1234,In_1456);
and U328 (N_328,In_1847,In_1564);
nor U329 (N_329,In_1641,In_1134);
nand U330 (N_330,In_1897,In_1532);
nor U331 (N_331,In_1999,In_1719);
or U332 (N_332,In_385,In_1254);
and U333 (N_333,In_1600,In_1826);
and U334 (N_334,In_1810,In_500);
nor U335 (N_335,In_598,In_1185);
nand U336 (N_336,In_838,In_844);
nand U337 (N_337,In_1051,In_1278);
nor U338 (N_338,In_297,In_1442);
and U339 (N_339,In_594,In_149);
nand U340 (N_340,In_473,In_478);
and U341 (N_341,In_564,In_1293);
nand U342 (N_342,In_107,In_1871);
nor U343 (N_343,In_1386,In_1162);
nand U344 (N_344,In_1350,In_397);
nand U345 (N_345,In_17,In_570);
nand U346 (N_346,In_1611,In_252);
or U347 (N_347,In_689,In_1177);
nand U348 (N_348,In_131,In_664);
nor U349 (N_349,In_1,In_275);
or U350 (N_350,In_1770,In_1576);
or U351 (N_351,In_1680,In_966);
nand U352 (N_352,In_1197,In_577);
nand U353 (N_353,In_1217,In_1769);
and U354 (N_354,In_1345,In_1123);
xnor U355 (N_355,In_185,In_1063);
nor U356 (N_356,In_547,In_941);
or U357 (N_357,In_170,In_1045);
and U358 (N_358,In_894,In_580);
nor U359 (N_359,In_1963,In_1505);
and U360 (N_360,In_465,In_1514);
nor U361 (N_361,In_667,In_78);
and U362 (N_362,In_1579,In_1683);
and U363 (N_363,In_830,In_556);
nand U364 (N_364,In_833,In_1004);
or U365 (N_365,In_681,In_1300);
nand U366 (N_366,In_1229,In_355);
and U367 (N_367,In_1213,In_1985);
nor U368 (N_368,In_1046,In_1223);
nor U369 (N_369,In_1811,In_418);
and U370 (N_370,In_261,In_1984);
or U371 (N_371,In_1969,In_392);
or U372 (N_372,In_956,In_636);
and U373 (N_373,In_720,In_1809);
nor U374 (N_374,In_1128,In_1863);
or U375 (N_375,In_1396,In_56);
or U376 (N_376,In_1483,In_648);
nand U377 (N_377,In_1207,In_1268);
nand U378 (N_378,In_848,In_724);
and U379 (N_379,In_1889,In_1959);
and U380 (N_380,In_1011,In_324);
or U381 (N_381,In_1075,In_543);
nor U382 (N_382,In_1708,In_187);
and U383 (N_383,In_545,In_59);
or U384 (N_384,In_1898,In_429);
nor U385 (N_385,In_128,In_738);
and U386 (N_386,In_1602,In_1895);
nand U387 (N_387,In_1432,In_1592);
or U388 (N_388,In_1252,In_464);
and U389 (N_389,In_1815,In_1341);
and U390 (N_390,In_1171,In_1101);
and U391 (N_391,In_53,In_1434);
nand U392 (N_392,In_1440,In_905);
and U393 (N_393,In_463,In_1443);
or U394 (N_394,In_1368,In_1652);
nor U395 (N_395,In_586,In_1740);
or U396 (N_396,In_1125,In_41);
and U397 (N_397,In_1265,In_933);
and U398 (N_398,In_1261,In_1533);
nand U399 (N_399,In_1950,In_596);
and U400 (N_400,In_1544,In_445);
and U401 (N_401,In_1961,In_321);
nor U402 (N_402,In_1323,In_949);
nand U403 (N_403,In_1712,In_537);
nor U404 (N_404,In_1590,In_143);
or U405 (N_405,In_557,In_789);
nand U406 (N_406,In_834,In_1760);
and U407 (N_407,In_1715,In_1333);
nand U408 (N_408,In_1557,In_39);
nor U409 (N_409,In_105,In_948);
or U410 (N_410,In_1394,In_540);
or U411 (N_411,In_136,In_1749);
or U412 (N_412,In_1000,In_1542);
or U413 (N_413,In_434,In_1792);
nand U414 (N_414,In_1062,In_1339);
nor U415 (N_415,In_1078,In_608);
or U416 (N_416,In_1977,In_998);
nand U417 (N_417,In_742,In_851);
nor U418 (N_418,In_678,In_1995);
nand U419 (N_419,In_785,In_343);
or U420 (N_420,In_1909,In_1709);
or U421 (N_421,In_119,In_1320);
and U422 (N_422,In_1119,In_825);
nor U423 (N_423,In_1059,In_391);
nor U424 (N_424,In_602,In_645);
nor U425 (N_425,In_178,In_1058);
and U426 (N_426,In_1982,In_96);
nand U427 (N_427,In_1663,In_902);
or U428 (N_428,In_1347,In_793);
nor U429 (N_429,In_403,In_1098);
or U430 (N_430,In_1965,In_1933);
or U431 (N_431,In_388,In_684);
and U432 (N_432,In_1156,In_1288);
and U433 (N_433,In_1793,In_419);
nor U434 (N_434,In_616,In_779);
and U435 (N_435,In_404,In_486);
or U436 (N_436,In_1634,In_1759);
or U437 (N_437,In_499,In_957);
nand U438 (N_438,In_123,In_1983);
and U439 (N_439,In_1517,In_1437);
nor U440 (N_440,In_579,In_1580);
and U441 (N_441,In_1838,In_706);
nand U442 (N_442,In_1083,In_707);
or U443 (N_443,In_600,In_529);
or U444 (N_444,In_1428,In_394);
or U445 (N_445,In_313,In_203);
nand U446 (N_446,In_1650,In_363);
nand U447 (N_447,In_996,In_417);
and U448 (N_448,In_1633,In_364);
nor U449 (N_449,In_604,In_839);
nand U450 (N_450,In_186,In_1987);
or U451 (N_451,In_369,In_929);
and U452 (N_452,In_351,In_82);
nand U453 (N_453,In_531,In_378);
and U454 (N_454,In_912,In_160);
nand U455 (N_455,In_210,In_751);
nor U456 (N_456,In_493,In_1821);
and U457 (N_457,In_675,In_193);
nand U458 (N_458,In_1158,In_925);
nand U459 (N_459,In_528,In_85);
nor U460 (N_460,In_356,In_1029);
and U461 (N_461,In_750,In_1092);
or U462 (N_462,In_907,In_1492);
nand U463 (N_463,In_283,In_739);
or U464 (N_464,In_316,In_637);
nand U465 (N_465,In_51,In_1859);
or U466 (N_466,In_784,In_88);
nor U467 (N_467,In_1996,In_696);
or U468 (N_468,In_212,In_1096);
nor U469 (N_469,In_1836,In_857);
nand U470 (N_470,In_1801,In_216);
or U471 (N_471,In_1610,In_1124);
nor U472 (N_472,In_332,In_1943);
nand U473 (N_473,In_971,In_1928);
and U474 (N_474,In_1666,In_908);
nand U475 (N_475,In_623,In_336);
and U476 (N_476,In_611,In_609);
nand U477 (N_477,In_983,In_1227);
or U478 (N_478,In_930,In_1735);
nor U479 (N_479,In_1043,In_1015);
nand U480 (N_480,In_792,In_1146);
nand U481 (N_481,In_150,In_1414);
and U482 (N_482,In_1922,In_1473);
and U483 (N_483,In_254,In_1873);
nand U484 (N_484,In_433,In_1768);
and U485 (N_485,In_847,In_19);
nand U486 (N_486,In_669,In_524);
nor U487 (N_487,In_867,In_754);
nor U488 (N_488,In_335,In_264);
xnor U489 (N_489,In_606,In_485);
nor U490 (N_490,In_268,In_1245);
or U491 (N_491,In_1511,In_1585);
nand U492 (N_492,In_1767,In_767);
nand U493 (N_493,In_773,In_1875);
and U494 (N_494,In_327,In_118);
nor U495 (N_495,In_1753,In_376);
nand U496 (N_496,In_745,In_1215);
nand U497 (N_497,In_690,In_1952);
xnor U498 (N_498,In_1024,In_1415);
nor U499 (N_499,In_841,In_1377);
nor U500 (N_500,In_1005,In_1155);
and U501 (N_501,In_1292,In_1755);
and U502 (N_502,In_1318,In_169);
nand U503 (N_503,In_1957,In_13);
and U504 (N_504,In_1617,In_699);
and U505 (N_505,In_114,In_829);
nor U506 (N_506,In_303,In_282);
nand U507 (N_507,In_1945,In_1704);
and U508 (N_508,In_482,In_1775);
nand U509 (N_509,In_1072,In_1191);
and U510 (N_510,In_331,In_893);
or U511 (N_511,In_1508,In_1485);
nand U512 (N_512,In_248,In_48);
nand U513 (N_513,In_116,In_181);
nor U514 (N_514,In_1899,In_1827);
or U515 (N_515,In_999,In_1025);
and U516 (N_516,In_1154,In_1287);
and U517 (N_517,In_698,In_182);
nor U518 (N_518,In_1725,In_1681);
nor U519 (N_519,In_1281,In_1921);
nand U520 (N_520,In_1035,In_190);
and U521 (N_521,In_330,In_913);
nand U522 (N_522,In_1418,In_125);
nor U523 (N_523,In_1349,In_1237);
or U524 (N_524,In_1376,In_550);
nor U525 (N_525,In_1244,In_1894);
and U526 (N_526,In_869,In_77);
xor U527 (N_527,In_1746,In_1032);
and U528 (N_528,In_797,In_657);
nand U529 (N_529,In_628,In_1327);
or U530 (N_530,In_152,In_937);
nor U531 (N_531,In_634,In_174);
or U532 (N_532,In_1306,In_979);
nand U533 (N_533,In_700,In_1722);
nor U534 (N_534,In_952,In_974);
xnor U535 (N_535,In_8,In_111);
nor U536 (N_536,In_884,In_99);
nand U537 (N_537,In_705,In_1365);
and U538 (N_538,In_184,In_1501);
nor U539 (N_539,In_1359,In_295);
nand U540 (N_540,In_1160,In_1095);
or U541 (N_541,In_1844,In_1053);
nor U542 (N_542,In_1554,In_1820);
nand U543 (N_543,In_630,In_1668);
and U544 (N_544,In_842,In_1570);
or U545 (N_545,In_1303,In_1009);
nand U546 (N_546,In_1017,In_389);
and U547 (N_547,In_747,In_1126);
or U548 (N_548,In_982,In_90);
or U549 (N_549,In_115,In_895);
nand U550 (N_550,In_1637,In_1968);
nand U551 (N_551,In_618,In_1190);
nor U552 (N_552,In_835,In_713);
nor U553 (N_553,In_140,In_1210);
and U554 (N_554,In_237,In_1108);
nand U555 (N_555,In_1684,In_1892);
or U556 (N_556,In_165,In_1690);
nor U557 (N_557,In_1503,In_633);
nor U558 (N_558,In_1623,In_522);
nor U559 (N_559,In_1858,In_102);
or U560 (N_560,In_661,In_963);
nor U561 (N_561,In_806,In_1850);
or U562 (N_562,In_1591,In_126);
nor U563 (N_563,In_1319,In_1270);
nor U564 (N_564,In_972,In_1421);
xor U565 (N_565,In_448,In_715);
nor U566 (N_566,In_1940,In_1997);
or U567 (N_567,In_1593,In_994);
nand U568 (N_568,In_1453,In_1548);
nand U569 (N_569,In_4,In_328);
and U570 (N_570,In_1835,In_366);
nor U571 (N_571,In_1614,In_346);
nor U572 (N_572,In_354,In_1204);
nand U573 (N_573,In_567,In_489);
nor U574 (N_574,In_461,In_525);
or U575 (N_575,In_22,In_718);
nor U576 (N_576,In_1393,In_269);
and U577 (N_577,In_233,In_1644);
nor U578 (N_578,In_762,In_1120);
nor U579 (N_579,In_122,In_727);
and U580 (N_580,In_1321,In_1837);
and U581 (N_581,In_768,In_1903);
or U582 (N_582,In_866,In_565);
nor U583 (N_583,In_36,In_65);
or U584 (N_584,In_1687,In_1971);
and U585 (N_585,In_1688,In_1624);
or U586 (N_586,In_1706,In_673);
nor U587 (N_587,In_1972,In_398);
nand U588 (N_588,In_44,In_1422);
nand U589 (N_589,In_1139,In_162);
nor U590 (N_590,In_1893,In_1383);
nor U591 (N_591,In_299,In_854);
or U592 (N_592,In_1841,In_1541);
nor U593 (N_593,In_726,In_207);
xnor U594 (N_594,In_1028,In_790);
nor U595 (N_595,In_1235,In_58);
nor U596 (N_596,In_1149,In_1572);
nor U597 (N_597,In_1375,In_444);
and U598 (N_598,In_523,In_309);
nand U599 (N_599,In_886,In_1596);
nor U600 (N_600,In_911,In_1828);
or U601 (N_601,In_381,In_1936);
nand U602 (N_602,In_1469,In_976);
nand U603 (N_603,In_1036,In_1208);
nand U604 (N_604,In_1069,In_1109);
or U605 (N_605,In_469,In_859);
and U606 (N_606,In_414,In_1366);
or U607 (N_607,In_1890,In_315);
and U608 (N_608,In_1258,In_1914);
nor U609 (N_609,In_622,In_101);
or U610 (N_610,In_1799,In_781);
nor U611 (N_611,In_69,In_1878);
or U612 (N_612,In_542,In_468);
or U613 (N_613,In_1220,In_1397);
xor U614 (N_614,In_1478,In_347);
and U615 (N_615,In_1027,In_1829);
or U616 (N_616,In_1335,In_1304);
and U617 (N_617,In_1294,In_457);
xor U618 (N_618,In_1881,In_1494);
nor U619 (N_619,In_882,In_221);
and U620 (N_620,In_1609,In_33);
and U621 (N_621,In_301,In_1264);
or U622 (N_622,In_1616,In_1718);
xnor U623 (N_623,In_1006,In_807);
nor U624 (N_624,In_1910,In_511);
and U625 (N_625,In_1395,In_1635);
nor U626 (N_626,In_1703,In_787);
or U627 (N_627,In_1781,In_701);
and U628 (N_628,In_1363,In_329);
and U629 (N_629,In_393,In_1625);
nor U630 (N_630,In_280,In_127);
nand U631 (N_631,In_1877,In_1493);
or U632 (N_632,In_584,In_711);
and U633 (N_633,In_1789,In_1507);
or U634 (N_634,In_214,In_171);
nor U635 (N_635,In_244,In_1731);
nand U636 (N_636,In_222,In_1865);
and U637 (N_637,In_1384,In_704);
nand U638 (N_638,In_60,In_191);
or U639 (N_639,In_585,In_66);
nor U640 (N_640,In_1354,In_1930);
nor U641 (N_641,In_898,In_975);
nor U642 (N_642,In_1932,In_1449);
and U643 (N_643,In_1358,In_450);
nand U644 (N_644,In_1253,In_582);
nor U645 (N_645,In_1479,In_1565);
nand U646 (N_646,In_649,In_1218);
and U647 (N_647,In_1737,In_1033);
or U648 (N_648,In_672,In_680);
or U649 (N_649,In_1331,In_1823);
nor U650 (N_650,In_1427,In_771);
nor U651 (N_651,In_415,In_307);
or U652 (N_652,In_1929,In_810);
nand U653 (N_653,In_1916,In_55);
or U654 (N_654,In_617,In_1100);
and U655 (N_655,In_1460,In_1840);
and U656 (N_656,In_1111,In_289);
nor U657 (N_657,In_1340,In_1280);
and U658 (N_658,In_1698,In_1431);
nor U659 (N_659,In_1482,In_496);
and U660 (N_660,In_488,In_840);
or U661 (N_661,In_1701,In_555);
or U662 (N_662,In_1405,In_287);
or U663 (N_663,In_590,In_1232);
xnor U664 (N_664,In_644,In_271);
or U665 (N_665,In_479,In_1048);
nand U666 (N_666,In_1872,In_477);
nand U667 (N_667,In_1569,In_1496);
nor U668 (N_668,In_695,In_1667);
nand U669 (N_669,In_915,In_61);
and U670 (N_670,In_1671,In_1420);
nor U671 (N_671,In_3,In_293);
and U672 (N_672,In_163,In_1577);
and U673 (N_673,In_1905,In_817);
or U674 (N_674,In_412,In_758);
nand U675 (N_675,In_322,In_1042);
or U676 (N_676,In_1976,In_1778);
and U677 (N_677,In_1106,In_703);
or U678 (N_678,In_292,In_1948);
and U679 (N_679,In_1231,In_16);
nor U680 (N_680,In_1713,In_1201);
and U681 (N_681,In_92,In_1241);
xnor U682 (N_682,In_350,In_763);
and U683 (N_683,In_1621,In_1474);
nand U684 (N_684,In_993,In_158);
nand U685 (N_685,In_290,In_1180);
and U686 (N_686,In_1538,In_517);
nor U687 (N_687,In_194,In_1677);
and U688 (N_688,In_1186,In_914);
nand U689 (N_689,In_1700,In_836);
or U690 (N_690,In_141,In_1561);
nand U691 (N_691,In_775,In_1608);
or U692 (N_692,In_1906,In_1387);
nand U693 (N_693,In_372,In_1907);
nand U694 (N_694,In_967,In_1848);
nor U695 (N_695,In_68,In_426);
xor U696 (N_696,In_597,In_940);
nor U697 (N_697,In_1853,In_1176);
and U698 (N_698,In_1992,In_24);
nand U699 (N_699,In_1536,In_1630);
or U700 (N_700,In_1917,In_1165);
xnor U701 (N_701,In_296,In_581);
or U702 (N_702,In_1896,In_1518);
or U703 (N_703,In_10,In_1209);
nand U704 (N_704,In_1274,In_748);
and U705 (N_705,In_1639,In_1754);
and U706 (N_706,In_64,In_1400);
nand U707 (N_707,In_1528,In_1562);
nand U708 (N_708,In_725,In_67);
nand U709 (N_709,In_215,In_1433);
nor U710 (N_710,In_668,In_1686);
nor U711 (N_711,In_883,In_1861);
or U712 (N_712,In_1269,In_1127);
nand U713 (N_713,In_117,In_1105);
nor U714 (N_714,In_424,In_228);
or U715 (N_715,In_483,In_752);
nand U716 (N_716,In_799,In_1504);
nor U717 (N_717,In_1927,In_1764);
xor U718 (N_718,In_625,In_735);
nand U719 (N_719,In_402,In_788);
nand U720 (N_720,In_677,In_1724);
nand U721 (N_721,In_666,In_1159);
or U722 (N_722,In_42,In_1457);
nand U723 (N_723,In_845,In_262);
and U724 (N_724,In_1056,In_916);
nand U725 (N_725,In_238,In_1649);
and U726 (N_726,In_1364,In_37);
or U727 (N_727,In_246,In_1330);
and U728 (N_728,In_709,In_217);
nand U729 (N_729,In_1632,In_688);
or U730 (N_730,In_1077,In_1947);
nor U731 (N_731,In_209,In_1563);
nand U732 (N_732,In_192,In_1312);
nand U733 (N_733,In_730,In_850);
and U734 (N_734,In_1066,In_1851);
nor U735 (N_735,In_805,In_1800);
or U736 (N_736,In_702,In_935);
nor U737 (N_737,In_552,In_1074);
and U738 (N_738,In_446,In_110);
or U739 (N_739,In_885,In_874);
or U740 (N_740,In_1849,In_1925);
and U741 (N_741,In_1470,In_462);
nand U742 (N_742,In_1990,In_438);
or U743 (N_743,In_629,In_777);
or U744 (N_744,In_989,In_928);
nor U745 (N_745,In_1547,In_1093);
nor U746 (N_746,In_453,In_395);
and U747 (N_747,In_687,In_1931);
nand U748 (N_748,In_1390,In_1022);
nor U749 (N_749,In_1486,In_1010);
or U750 (N_750,In_1221,In_1819);
and U751 (N_751,In_352,In_802);
nand U752 (N_752,In_1714,In_1361);
and U753 (N_753,In_861,In_1727);
nor U754 (N_754,In_714,In_1382);
nor U755 (N_755,In_501,In_1079);
and U756 (N_756,In_1817,In_334);
nand U757 (N_757,In_230,In_1242);
nor U758 (N_758,In_1067,In_1571);
and U759 (N_759,In_242,In_1332);
or U760 (N_760,In_1738,In_1594);
and U761 (N_761,In_1018,In_1842);
and U762 (N_762,In_161,In_1178);
nor U763 (N_763,In_132,In_45);
or U764 (N_764,In_1802,In_944);
and U765 (N_765,In_960,In_1526);
nand U766 (N_766,In_961,In_401);
or U767 (N_767,In_146,In_878);
and U768 (N_768,In_563,In_1465);
or U769 (N_769,In_456,In_1675);
nand U770 (N_770,In_1003,In_224);
nor U771 (N_771,In_873,In_270);
or U772 (N_772,In_1054,In_1578);
or U773 (N_773,In_147,In_213);
or U774 (N_774,In_1189,In_1843);
or U775 (N_775,In_1581,In_1934);
or U776 (N_776,In_1524,In_1297);
nand U777 (N_777,In_377,In_1962);
nor U778 (N_778,In_1568,In_1989);
and U779 (N_779,In_1519,In_386);
and U780 (N_780,In_1299,In_1413);
and U781 (N_781,In_901,In_800);
or U782 (N_782,In_1595,In_1745);
nor U783 (N_783,In_1857,In_655);
or U784 (N_784,In_1094,In_1642);
or U785 (N_785,In_379,In_1379);
nor U786 (N_786,In_38,In_416);
nor U787 (N_787,In_1864,In_1994);
or U788 (N_788,In_1891,In_619);
or U789 (N_789,In_743,In_986);
nand U790 (N_790,In_1946,In_918);
and U791 (N_791,In_1211,In_317);
and U792 (N_792,In_312,In_427);
or U793 (N_793,In_1203,In_396);
xor U794 (N_794,In_756,In_889);
nand U795 (N_795,In_796,In_991);
and U796 (N_796,In_27,In_1535);
xor U797 (N_797,In_1102,In_1250);
or U798 (N_798,In_1305,In_1956);
nand U799 (N_799,In_795,In_1271);
or U800 (N_800,In_1298,In_1685);
nand U801 (N_801,In_1451,In_1381);
nor U802 (N_802,In_1604,In_1522);
nand U803 (N_803,In_1041,In_430);
xnor U804 (N_804,In_466,In_955);
nand U805 (N_805,In_1173,In_1834);
or U806 (N_806,In_1512,In_15);
nand U807 (N_807,In_1249,In_1408);
and U808 (N_808,In_1142,In_113);
nor U809 (N_809,In_903,In_21);
nand U810 (N_810,In_432,In_492);
nand U811 (N_811,In_621,In_1170);
nand U812 (N_812,In_1904,In_1657);
or U813 (N_813,In_1122,In_1317);
xnor U814 (N_814,In_196,In_1699);
nand U815 (N_815,In_1324,In_1348);
or U816 (N_816,In_1374,In_822);
or U817 (N_817,In_964,In_818);
and U818 (N_818,In_831,In_572);
nor U819 (N_819,In_1613,In_1676);
or U820 (N_820,In_1157,In_1966);
nor U821 (N_821,In_1034,In_1052);
nor U822 (N_822,In_1222,In_345);
nor U823 (N_823,In_79,In_549);
nor U824 (N_824,In_495,In_801);
nor U825 (N_825,In_286,In_1750);
and U826 (N_826,In_1309,In_1658);
or U827 (N_827,In_1495,In_890);
nor U828 (N_828,In_120,In_1455);
nor U829 (N_829,In_451,In_660);
nor U830 (N_830,In_1167,In_761);
or U831 (N_831,In_1169,In_1466);
and U832 (N_832,In_593,In_9);
or U833 (N_833,In_138,In_1040);
and U834 (N_834,In_774,In_879);
and U835 (N_835,In_74,In_849);
nand U836 (N_836,In_1525,In_387);
nor U837 (N_837,In_1360,In_1490);
nor U838 (N_838,In_1247,In_1391);
nand U839 (N_839,In_1477,In_183);
nor U840 (N_840,In_200,In_1876);
or U841 (N_841,In_576,In_455);
nand U842 (N_842,In_201,In_1283);
or U843 (N_843,In_195,In_1669);
xnor U844 (N_844,In_1342,In_1012);
or U845 (N_845,In_1487,In_813);
xor U846 (N_846,In_503,In_1530);
nor U847 (N_847,In_34,In_973);
or U848 (N_848,In_1424,In_323);
nand U849 (N_849,In_513,In_780);
and U850 (N_850,In_1980,In_400);
nand U851 (N_851,In_421,In_253);
nor U852 (N_852,In_20,In_365);
or U853 (N_853,In_1527,In_472);
or U854 (N_854,In_510,In_712);
nand U855 (N_855,In_1228,In_821);
nor U856 (N_856,In_260,In_326);
and U857 (N_857,In_592,In_1001);
nor U858 (N_858,In_932,In_1409);
or U859 (N_859,In_1763,In_1831);
nor U860 (N_860,In_746,In_348);
nor U861 (N_861,In_652,In_1462);
nor U862 (N_862,In_1788,In_410);
and U863 (N_863,In_1116,In_1964);
nand U864 (N_864,In_1370,In_1885);
and U865 (N_865,In_357,In_1804);
and U866 (N_866,In_1654,In_1372);
nand U867 (N_867,In_159,In_458);
or U868 (N_868,In_1426,In_1026);
nand U869 (N_869,In_1497,In_870);
and U870 (N_870,In_1308,In_1225);
nor U871 (N_871,In_1282,In_1284);
nor U872 (N_872,In_1777,In_281);
and U873 (N_873,In_142,In_1721);
nand U874 (N_874,In_1780,In_772);
or U875 (N_875,In_43,In_1307);
and U876 (N_876,In_1295,In_980);
and U877 (N_877,In_1301,In_239);
nand U878 (N_878,In_782,In_1855);
nand U879 (N_879,In_1047,In_603);
or U880 (N_880,In_733,In_407);
or U881 (N_881,In_1901,In_615);
and U882 (N_882,In_1808,In_1246);
or U883 (N_883,In_526,In_1239);
or U884 (N_884,In_1329,In_812);
nor U885 (N_885,In_969,In_1016);
and U886 (N_886,In_953,In_1285);
nand U887 (N_887,In_1766,In_211);
nand U888 (N_888,In_6,In_587);
or U889 (N_889,In_1812,In_1734);
nand U890 (N_890,In_1194,In_1110);
nor U891 (N_891,In_1866,In_1439);
or U892 (N_892,In_235,In_1546);
nand U893 (N_893,In_1908,In_1938);
nor U894 (N_894,In_544,In_837);
or U895 (N_895,In_872,In_231);
nor U896 (N_896,In_197,In_663);
or U897 (N_897,In_1551,In_1774);
nor U898 (N_898,In_1958,In_1404);
nor U899 (N_899,In_1942,In_1444);
xor U900 (N_900,In_786,In_1014);
and U901 (N_901,In_1597,In_361);
or U902 (N_902,In_1334,In_1550);
nand U903 (N_903,In_936,In_1974);
or U904 (N_904,In_984,In_1410);
and U905 (N_905,In_1739,In_1960);
nor U906 (N_906,In_1794,In_1115);
or U907 (N_907,In_14,In_826);
and U908 (N_908,In_272,In_875);
and U909 (N_909,In_917,In_1694);
or U910 (N_910,In_888,In_559);
or U911 (N_911,In_481,In_1454);
or U912 (N_912,In_1923,In_1037);
or U913 (N_913,In_1248,In_1567);
or U914 (N_914,In_541,In_1748);
nor U915 (N_915,In_29,In_30);
nand U916 (N_916,In_1790,In_370);
and U917 (N_917,In_1730,In_1152);
or U918 (N_918,In_50,In_1975);
and U919 (N_919,In_820,In_1435);
or U920 (N_920,In_1647,In_1993);
and U921 (N_921,In_1267,In_1643);
or U922 (N_922,In_1586,In_1351);
or U923 (N_923,In_1941,In_1099);
nor U924 (N_924,In_1711,In_1782);
nor U925 (N_925,In_1967,In_1603);
nand U926 (N_926,In_199,In_1020);
nand U927 (N_927,In_284,In_155);
nor U928 (N_928,In_2,In_1168);
or U929 (N_929,In_946,In_1192);
nor U930 (N_930,In_87,In_819);
nor U931 (N_931,In_551,In_148);
nand U932 (N_932,In_1845,In_665);
and U933 (N_933,In_1670,In_1065);
nand U934 (N_934,In_1771,In_1589);
nand U935 (N_935,In_509,In_1416);
nand U936 (N_936,In_741,In_1140);
and U937 (N_937,In_1179,In_12);
nor U938 (N_938,In_759,In_534);
nand U939 (N_939,In_1082,In_1491);
nand U940 (N_940,In_1742,In_206);
and U941 (N_941,In_342,In_1583);
and U942 (N_942,In_507,In_480);
nor U943 (N_943,In_1090,In_153);
and U944 (N_944,In_1798,In_1653);
nand U945 (N_945,In_1973,In_519);
nor U946 (N_946,In_896,In_1089);
nand U947 (N_947,In_595,In_920);
nor U948 (N_948,In_942,In_1918);
or U949 (N_949,In_241,In_76);
and U950 (N_950,In_561,In_910);
and U951 (N_951,In_1818,In_267);
and U952 (N_952,In_1513,In_1233);
and U953 (N_953,In_205,In_255);
nand U954 (N_954,In_1266,In_1824);
and U955 (N_955,In_475,In_135);
nor U956 (N_956,In_997,In_1468);
nor U957 (N_957,In_28,In_1935);
nand U958 (N_958,In_1353,In_1219);
nor U959 (N_959,In_1814,In_1071);
and U960 (N_960,In_1622,In_502);
nor U961 (N_961,In_1337,In_18);
or U962 (N_962,In_1328,In_1888);
and U963 (N_963,In_1369,In_1073);
nand U964 (N_964,In_1136,In_1107);
and U965 (N_965,In_1732,In_945);
or U966 (N_966,In_1736,In_755);
nand U967 (N_967,In_566,In_1373);
nand U968 (N_968,In_227,In_558);
and U969 (N_969,In_783,In_452);
nand U970 (N_970,In_1803,In_1900);
nor U971 (N_971,In_302,In_691);
nand U972 (N_972,In_1263,In_934);
and U973 (N_973,In_1874,In_498);
and U974 (N_974,In_1776,In_1260);
nand U975 (N_975,In_177,In_447);
or U976 (N_976,In_208,In_1472);
or U977 (N_977,In_1315,In_734);
nor U978 (N_978,In_26,In_1371);
nand U979 (N_979,In_653,In_333);
or U980 (N_980,In_1262,In_1599);
or U981 (N_981,In_1193,In_1772);
nand U982 (N_982,In_575,In_1645);
or U983 (N_983,In_75,In_154);
and U984 (N_984,In_1500,In_1463);
or U985 (N_985,In_729,In_538);
nand U986 (N_986,In_1407,In_539);
or U987 (N_987,In_1311,In_506);
nor U988 (N_988,In_234,In_1182);
nor U989 (N_989,In_1762,In_1978);
nor U990 (N_990,In_887,In_1132);
and U991 (N_991,In_736,In_375);
nand U992 (N_992,In_546,In_1626);
nand U993 (N_993,In_776,In_1076);
and U994 (N_994,In_1137,In_1355);
nor U995 (N_995,In_992,In_1911);
nor U996 (N_996,In_1238,In_536);
or U997 (N_997,In_1008,In_1523);
or U998 (N_998,In_1549,In_1574);
or U999 (N_999,In_273,In_380);
nor U1000 (N_1000,In_1678,In_702);
and U1001 (N_1001,In_1955,In_276);
nor U1002 (N_1002,In_869,In_1820);
and U1003 (N_1003,In_203,In_672);
and U1004 (N_1004,In_1259,In_1201);
and U1005 (N_1005,In_804,In_1685);
or U1006 (N_1006,In_568,In_1359);
nand U1007 (N_1007,In_1713,In_1203);
nand U1008 (N_1008,In_1726,In_1281);
or U1009 (N_1009,In_1537,In_1314);
or U1010 (N_1010,In_1269,In_535);
and U1011 (N_1011,In_1626,In_13);
nor U1012 (N_1012,In_429,In_941);
nor U1013 (N_1013,In_1530,In_1783);
nand U1014 (N_1014,In_927,In_130);
and U1015 (N_1015,In_556,In_1819);
nor U1016 (N_1016,In_1952,In_358);
or U1017 (N_1017,In_952,In_1440);
nor U1018 (N_1018,In_369,In_1392);
nor U1019 (N_1019,In_1382,In_1408);
xor U1020 (N_1020,In_389,In_1286);
nor U1021 (N_1021,In_1698,In_373);
and U1022 (N_1022,In_8,In_942);
nor U1023 (N_1023,In_1346,In_1009);
and U1024 (N_1024,In_1338,In_96);
nor U1025 (N_1025,In_1330,In_1512);
or U1026 (N_1026,In_1742,In_1537);
nand U1027 (N_1027,In_988,In_738);
nor U1028 (N_1028,In_818,In_358);
or U1029 (N_1029,In_1000,In_369);
and U1030 (N_1030,In_1500,In_1758);
nor U1031 (N_1031,In_1814,In_558);
and U1032 (N_1032,In_1458,In_1360);
nor U1033 (N_1033,In_409,In_627);
nand U1034 (N_1034,In_40,In_536);
nand U1035 (N_1035,In_1878,In_778);
and U1036 (N_1036,In_377,In_943);
or U1037 (N_1037,In_683,In_488);
nand U1038 (N_1038,In_737,In_404);
nor U1039 (N_1039,In_1522,In_1381);
or U1040 (N_1040,In_611,In_1934);
xor U1041 (N_1041,In_915,In_1906);
and U1042 (N_1042,In_336,In_218);
nor U1043 (N_1043,In_15,In_1303);
or U1044 (N_1044,In_581,In_1643);
nand U1045 (N_1045,In_1206,In_1388);
and U1046 (N_1046,In_1954,In_419);
or U1047 (N_1047,In_1392,In_345);
or U1048 (N_1048,In_653,In_16);
nand U1049 (N_1049,In_980,In_1144);
nand U1050 (N_1050,In_1134,In_568);
nor U1051 (N_1051,In_780,In_1136);
nor U1052 (N_1052,In_858,In_872);
nand U1053 (N_1053,In_1095,In_870);
or U1054 (N_1054,In_149,In_277);
and U1055 (N_1055,In_1568,In_915);
or U1056 (N_1056,In_759,In_124);
and U1057 (N_1057,In_1883,In_1899);
or U1058 (N_1058,In_1870,In_547);
or U1059 (N_1059,In_841,In_380);
nor U1060 (N_1060,In_70,In_325);
nand U1061 (N_1061,In_1224,In_892);
and U1062 (N_1062,In_1151,In_141);
nor U1063 (N_1063,In_591,In_1218);
or U1064 (N_1064,In_1767,In_109);
or U1065 (N_1065,In_1181,In_90);
and U1066 (N_1066,In_1270,In_313);
and U1067 (N_1067,In_191,In_1513);
and U1068 (N_1068,In_988,In_635);
or U1069 (N_1069,In_760,In_675);
nor U1070 (N_1070,In_1522,In_1119);
nand U1071 (N_1071,In_31,In_842);
or U1072 (N_1072,In_620,In_1459);
nand U1073 (N_1073,In_1251,In_1503);
and U1074 (N_1074,In_1767,In_311);
nor U1075 (N_1075,In_1133,In_1298);
or U1076 (N_1076,In_958,In_1274);
nor U1077 (N_1077,In_719,In_1860);
or U1078 (N_1078,In_1537,In_1852);
xor U1079 (N_1079,In_301,In_1165);
and U1080 (N_1080,In_750,In_690);
or U1081 (N_1081,In_1602,In_1907);
nor U1082 (N_1082,In_113,In_42);
nand U1083 (N_1083,In_293,In_1055);
nor U1084 (N_1084,In_1468,In_1401);
xor U1085 (N_1085,In_1962,In_986);
and U1086 (N_1086,In_1901,In_1615);
nand U1087 (N_1087,In_1968,In_642);
nor U1088 (N_1088,In_1704,In_217);
xnor U1089 (N_1089,In_1516,In_1949);
or U1090 (N_1090,In_365,In_724);
nor U1091 (N_1091,In_900,In_1227);
and U1092 (N_1092,In_1577,In_1208);
nor U1093 (N_1093,In_1107,In_1750);
nor U1094 (N_1094,In_1349,In_850);
xnor U1095 (N_1095,In_404,In_1541);
and U1096 (N_1096,In_860,In_98);
or U1097 (N_1097,In_1524,In_1135);
and U1098 (N_1098,In_893,In_162);
and U1099 (N_1099,In_427,In_26);
or U1100 (N_1100,In_1099,In_1850);
nor U1101 (N_1101,In_1919,In_1917);
or U1102 (N_1102,In_953,In_1050);
nor U1103 (N_1103,In_811,In_954);
nand U1104 (N_1104,In_1430,In_1881);
nand U1105 (N_1105,In_1287,In_683);
nand U1106 (N_1106,In_870,In_174);
and U1107 (N_1107,In_1312,In_593);
nor U1108 (N_1108,In_1788,In_1173);
nor U1109 (N_1109,In_454,In_1652);
or U1110 (N_1110,In_871,In_1872);
or U1111 (N_1111,In_341,In_1619);
nor U1112 (N_1112,In_273,In_1491);
or U1113 (N_1113,In_1922,In_1360);
nand U1114 (N_1114,In_1273,In_443);
nor U1115 (N_1115,In_255,In_291);
nand U1116 (N_1116,In_527,In_914);
nor U1117 (N_1117,In_1579,In_189);
nor U1118 (N_1118,In_1130,In_971);
nor U1119 (N_1119,In_1274,In_441);
nand U1120 (N_1120,In_1902,In_500);
or U1121 (N_1121,In_1551,In_1042);
and U1122 (N_1122,In_632,In_177);
nand U1123 (N_1123,In_995,In_1670);
nor U1124 (N_1124,In_210,In_1037);
nand U1125 (N_1125,In_184,In_1067);
or U1126 (N_1126,In_1447,In_825);
nor U1127 (N_1127,In_743,In_598);
or U1128 (N_1128,In_1737,In_1648);
nor U1129 (N_1129,In_1993,In_1453);
nand U1130 (N_1130,In_1619,In_1851);
xor U1131 (N_1131,In_1715,In_1347);
and U1132 (N_1132,In_1884,In_605);
or U1133 (N_1133,In_1868,In_1423);
nand U1134 (N_1134,In_885,In_276);
and U1135 (N_1135,In_1917,In_1673);
or U1136 (N_1136,In_89,In_334);
or U1137 (N_1137,In_1576,In_1271);
and U1138 (N_1138,In_643,In_1854);
and U1139 (N_1139,In_898,In_1469);
xnor U1140 (N_1140,In_1406,In_292);
or U1141 (N_1141,In_1367,In_1819);
or U1142 (N_1142,In_427,In_187);
nor U1143 (N_1143,In_107,In_480);
nor U1144 (N_1144,In_244,In_181);
and U1145 (N_1145,In_1284,In_624);
nand U1146 (N_1146,In_1730,In_54);
nand U1147 (N_1147,In_938,In_1228);
nand U1148 (N_1148,In_442,In_429);
and U1149 (N_1149,In_125,In_1182);
and U1150 (N_1150,In_381,In_1624);
nor U1151 (N_1151,In_1627,In_1350);
or U1152 (N_1152,In_1388,In_751);
nand U1153 (N_1153,In_1450,In_949);
and U1154 (N_1154,In_1212,In_1062);
and U1155 (N_1155,In_743,In_1328);
nand U1156 (N_1156,In_1195,In_721);
or U1157 (N_1157,In_684,In_275);
nor U1158 (N_1158,In_1130,In_1835);
and U1159 (N_1159,In_666,In_1663);
nor U1160 (N_1160,In_1515,In_1757);
nand U1161 (N_1161,In_1400,In_1525);
or U1162 (N_1162,In_24,In_1483);
and U1163 (N_1163,In_1858,In_819);
or U1164 (N_1164,In_750,In_314);
or U1165 (N_1165,In_1092,In_1645);
nor U1166 (N_1166,In_904,In_1966);
nand U1167 (N_1167,In_966,In_1325);
nor U1168 (N_1168,In_1751,In_34);
or U1169 (N_1169,In_1029,In_128);
or U1170 (N_1170,In_163,In_581);
nor U1171 (N_1171,In_1801,In_1989);
nand U1172 (N_1172,In_1561,In_1495);
and U1173 (N_1173,In_1460,In_1999);
nand U1174 (N_1174,In_1911,In_1802);
and U1175 (N_1175,In_1412,In_936);
nor U1176 (N_1176,In_1740,In_324);
nor U1177 (N_1177,In_1243,In_1192);
or U1178 (N_1178,In_1079,In_407);
and U1179 (N_1179,In_860,In_892);
nand U1180 (N_1180,In_353,In_871);
and U1181 (N_1181,In_1141,In_483);
nand U1182 (N_1182,In_1830,In_1827);
and U1183 (N_1183,In_774,In_1031);
nand U1184 (N_1184,In_675,In_436);
and U1185 (N_1185,In_1819,In_1294);
or U1186 (N_1186,In_177,In_1816);
nor U1187 (N_1187,In_547,In_1108);
or U1188 (N_1188,In_1682,In_1021);
nand U1189 (N_1189,In_1977,In_64);
nand U1190 (N_1190,In_980,In_1665);
nor U1191 (N_1191,In_1275,In_400);
and U1192 (N_1192,In_1035,In_134);
and U1193 (N_1193,In_237,In_571);
and U1194 (N_1194,In_198,In_1268);
nand U1195 (N_1195,In_1370,In_1577);
and U1196 (N_1196,In_717,In_1428);
or U1197 (N_1197,In_1452,In_744);
nand U1198 (N_1198,In_1507,In_468);
nor U1199 (N_1199,In_1502,In_52);
xor U1200 (N_1200,In_1100,In_826);
or U1201 (N_1201,In_1186,In_705);
and U1202 (N_1202,In_1731,In_611);
or U1203 (N_1203,In_1577,In_1406);
nor U1204 (N_1204,In_1615,In_1711);
and U1205 (N_1205,In_1690,In_340);
nand U1206 (N_1206,In_1304,In_914);
or U1207 (N_1207,In_1174,In_642);
nor U1208 (N_1208,In_555,In_1623);
or U1209 (N_1209,In_1329,In_1221);
nor U1210 (N_1210,In_1558,In_579);
and U1211 (N_1211,In_1851,In_625);
and U1212 (N_1212,In_624,In_1724);
or U1213 (N_1213,In_416,In_994);
and U1214 (N_1214,In_442,In_385);
and U1215 (N_1215,In_23,In_1533);
or U1216 (N_1216,In_754,In_13);
and U1217 (N_1217,In_160,In_782);
nor U1218 (N_1218,In_764,In_870);
or U1219 (N_1219,In_114,In_768);
and U1220 (N_1220,In_289,In_1627);
nor U1221 (N_1221,In_621,In_802);
and U1222 (N_1222,In_215,In_332);
nor U1223 (N_1223,In_624,In_1403);
nand U1224 (N_1224,In_335,In_1891);
nand U1225 (N_1225,In_173,In_957);
nand U1226 (N_1226,In_1255,In_1581);
nor U1227 (N_1227,In_69,In_1903);
nor U1228 (N_1228,In_536,In_96);
nand U1229 (N_1229,In_762,In_612);
nor U1230 (N_1230,In_1429,In_1859);
or U1231 (N_1231,In_1122,In_26);
nand U1232 (N_1232,In_533,In_1618);
or U1233 (N_1233,In_1747,In_1464);
nand U1234 (N_1234,In_185,In_569);
nand U1235 (N_1235,In_1268,In_44);
or U1236 (N_1236,In_410,In_1924);
xnor U1237 (N_1237,In_366,In_1082);
and U1238 (N_1238,In_1879,In_1);
nor U1239 (N_1239,In_1645,In_780);
nor U1240 (N_1240,In_373,In_1443);
or U1241 (N_1241,In_91,In_1709);
or U1242 (N_1242,In_836,In_151);
or U1243 (N_1243,In_909,In_898);
and U1244 (N_1244,In_228,In_1324);
xnor U1245 (N_1245,In_37,In_965);
or U1246 (N_1246,In_321,In_1389);
and U1247 (N_1247,In_1,In_1716);
and U1248 (N_1248,In_254,In_156);
xor U1249 (N_1249,In_1254,In_863);
nand U1250 (N_1250,In_1602,In_1531);
or U1251 (N_1251,In_1623,In_576);
and U1252 (N_1252,In_380,In_1832);
and U1253 (N_1253,In_1500,In_426);
nand U1254 (N_1254,In_616,In_1073);
nand U1255 (N_1255,In_675,In_440);
or U1256 (N_1256,In_1312,In_179);
nand U1257 (N_1257,In_350,In_3);
and U1258 (N_1258,In_1167,In_1969);
or U1259 (N_1259,In_1250,In_612);
and U1260 (N_1260,In_1309,In_1933);
and U1261 (N_1261,In_1177,In_1413);
nand U1262 (N_1262,In_1863,In_662);
or U1263 (N_1263,In_1998,In_878);
or U1264 (N_1264,In_109,In_1698);
nand U1265 (N_1265,In_354,In_970);
and U1266 (N_1266,In_1605,In_656);
and U1267 (N_1267,In_554,In_937);
or U1268 (N_1268,In_1632,In_1582);
nor U1269 (N_1269,In_511,In_1373);
nand U1270 (N_1270,In_1998,In_1972);
or U1271 (N_1271,In_1646,In_1422);
nor U1272 (N_1272,In_535,In_940);
and U1273 (N_1273,In_715,In_852);
or U1274 (N_1274,In_417,In_898);
and U1275 (N_1275,In_755,In_540);
or U1276 (N_1276,In_1260,In_1758);
nor U1277 (N_1277,In_422,In_1376);
nor U1278 (N_1278,In_121,In_1647);
and U1279 (N_1279,In_1796,In_411);
or U1280 (N_1280,In_547,In_761);
nand U1281 (N_1281,In_1289,In_587);
nand U1282 (N_1282,In_11,In_17);
and U1283 (N_1283,In_574,In_1187);
or U1284 (N_1284,In_195,In_887);
nand U1285 (N_1285,In_1178,In_1342);
nor U1286 (N_1286,In_33,In_1114);
nand U1287 (N_1287,In_1357,In_383);
nand U1288 (N_1288,In_1542,In_210);
xnor U1289 (N_1289,In_655,In_16);
nand U1290 (N_1290,In_992,In_1445);
or U1291 (N_1291,In_1940,In_1179);
or U1292 (N_1292,In_1906,In_1077);
or U1293 (N_1293,In_1136,In_1715);
xor U1294 (N_1294,In_1279,In_661);
and U1295 (N_1295,In_53,In_84);
nand U1296 (N_1296,In_669,In_1011);
or U1297 (N_1297,In_1003,In_918);
or U1298 (N_1298,In_199,In_4);
nor U1299 (N_1299,In_1294,In_1552);
nor U1300 (N_1300,In_333,In_867);
or U1301 (N_1301,In_1508,In_1731);
nand U1302 (N_1302,In_1680,In_1196);
and U1303 (N_1303,In_1108,In_1547);
or U1304 (N_1304,In_419,In_1184);
xor U1305 (N_1305,In_1692,In_457);
nand U1306 (N_1306,In_1774,In_998);
and U1307 (N_1307,In_1030,In_527);
nor U1308 (N_1308,In_439,In_134);
nand U1309 (N_1309,In_841,In_1051);
or U1310 (N_1310,In_1088,In_167);
or U1311 (N_1311,In_1680,In_373);
xor U1312 (N_1312,In_1804,In_1851);
nor U1313 (N_1313,In_979,In_1840);
xor U1314 (N_1314,In_314,In_1238);
nor U1315 (N_1315,In_1226,In_1367);
nor U1316 (N_1316,In_870,In_507);
and U1317 (N_1317,In_1536,In_182);
or U1318 (N_1318,In_1816,In_437);
nand U1319 (N_1319,In_1535,In_802);
and U1320 (N_1320,In_45,In_270);
and U1321 (N_1321,In_71,In_1227);
nand U1322 (N_1322,In_853,In_1264);
or U1323 (N_1323,In_1682,In_1524);
nand U1324 (N_1324,In_157,In_1222);
and U1325 (N_1325,In_7,In_1796);
nor U1326 (N_1326,In_552,In_1073);
nor U1327 (N_1327,In_1125,In_1320);
nand U1328 (N_1328,In_1153,In_791);
or U1329 (N_1329,In_1336,In_727);
or U1330 (N_1330,In_1829,In_1859);
nand U1331 (N_1331,In_778,In_1532);
nand U1332 (N_1332,In_1580,In_139);
nor U1333 (N_1333,In_1219,In_1860);
nor U1334 (N_1334,In_891,In_1894);
or U1335 (N_1335,In_1707,In_424);
nand U1336 (N_1336,In_1291,In_1822);
or U1337 (N_1337,In_1438,In_420);
or U1338 (N_1338,In_983,In_1470);
or U1339 (N_1339,In_1279,In_1524);
nor U1340 (N_1340,In_1605,In_1547);
nor U1341 (N_1341,In_1152,In_1407);
and U1342 (N_1342,In_360,In_779);
nand U1343 (N_1343,In_380,In_332);
nor U1344 (N_1344,In_1713,In_733);
and U1345 (N_1345,In_1761,In_821);
nor U1346 (N_1346,In_611,In_1518);
or U1347 (N_1347,In_296,In_1911);
and U1348 (N_1348,In_1562,In_1219);
and U1349 (N_1349,In_1947,In_681);
and U1350 (N_1350,In_1222,In_457);
nor U1351 (N_1351,In_29,In_70);
xnor U1352 (N_1352,In_834,In_620);
nor U1353 (N_1353,In_250,In_211);
nand U1354 (N_1354,In_1058,In_1239);
nor U1355 (N_1355,In_616,In_1336);
nor U1356 (N_1356,In_39,In_956);
nand U1357 (N_1357,In_1621,In_285);
nor U1358 (N_1358,In_1850,In_531);
nor U1359 (N_1359,In_1541,In_657);
nor U1360 (N_1360,In_794,In_1118);
and U1361 (N_1361,In_1913,In_1600);
and U1362 (N_1362,In_258,In_748);
and U1363 (N_1363,In_1692,In_1697);
nor U1364 (N_1364,In_545,In_1594);
nor U1365 (N_1365,In_1353,In_1986);
and U1366 (N_1366,In_1174,In_1069);
or U1367 (N_1367,In_1541,In_1706);
nand U1368 (N_1368,In_575,In_1564);
nor U1369 (N_1369,In_1583,In_175);
and U1370 (N_1370,In_1258,In_992);
and U1371 (N_1371,In_1204,In_537);
nor U1372 (N_1372,In_90,In_1949);
xnor U1373 (N_1373,In_1768,In_1757);
nand U1374 (N_1374,In_872,In_857);
nor U1375 (N_1375,In_1787,In_93);
nor U1376 (N_1376,In_38,In_226);
or U1377 (N_1377,In_845,In_1430);
or U1378 (N_1378,In_146,In_65);
and U1379 (N_1379,In_1889,In_947);
and U1380 (N_1380,In_1236,In_219);
and U1381 (N_1381,In_83,In_1883);
or U1382 (N_1382,In_1486,In_1537);
nand U1383 (N_1383,In_1260,In_1247);
nor U1384 (N_1384,In_1866,In_920);
nor U1385 (N_1385,In_1990,In_56);
nand U1386 (N_1386,In_1008,In_1556);
and U1387 (N_1387,In_21,In_1849);
nor U1388 (N_1388,In_460,In_620);
and U1389 (N_1389,In_48,In_1741);
and U1390 (N_1390,In_505,In_347);
nand U1391 (N_1391,In_1387,In_837);
nand U1392 (N_1392,In_1861,In_1204);
and U1393 (N_1393,In_783,In_1043);
nand U1394 (N_1394,In_997,In_979);
or U1395 (N_1395,In_1183,In_1826);
nor U1396 (N_1396,In_1412,In_430);
or U1397 (N_1397,In_799,In_914);
nand U1398 (N_1398,In_1940,In_1096);
xnor U1399 (N_1399,In_422,In_455);
or U1400 (N_1400,In_21,In_172);
or U1401 (N_1401,In_350,In_404);
nand U1402 (N_1402,In_251,In_1388);
or U1403 (N_1403,In_1400,In_676);
and U1404 (N_1404,In_1059,In_1890);
nor U1405 (N_1405,In_1752,In_1935);
nand U1406 (N_1406,In_139,In_1522);
nand U1407 (N_1407,In_123,In_492);
or U1408 (N_1408,In_697,In_1901);
or U1409 (N_1409,In_328,In_1542);
nand U1410 (N_1410,In_1541,In_1704);
nand U1411 (N_1411,In_512,In_518);
and U1412 (N_1412,In_1553,In_851);
nand U1413 (N_1413,In_891,In_712);
and U1414 (N_1414,In_1029,In_465);
and U1415 (N_1415,In_1618,In_1510);
or U1416 (N_1416,In_1736,In_1719);
or U1417 (N_1417,In_163,In_454);
nor U1418 (N_1418,In_133,In_277);
and U1419 (N_1419,In_551,In_89);
nor U1420 (N_1420,In_177,In_544);
nand U1421 (N_1421,In_737,In_1587);
and U1422 (N_1422,In_857,In_751);
and U1423 (N_1423,In_1063,In_1472);
nand U1424 (N_1424,In_470,In_137);
nor U1425 (N_1425,In_421,In_603);
nor U1426 (N_1426,In_185,In_1446);
or U1427 (N_1427,In_1543,In_121);
and U1428 (N_1428,In_748,In_591);
nor U1429 (N_1429,In_1891,In_1978);
and U1430 (N_1430,In_701,In_1777);
nand U1431 (N_1431,In_443,In_1199);
and U1432 (N_1432,In_554,In_625);
or U1433 (N_1433,In_637,In_538);
nand U1434 (N_1434,In_962,In_123);
nor U1435 (N_1435,In_1067,In_421);
or U1436 (N_1436,In_725,In_1406);
and U1437 (N_1437,In_871,In_846);
nor U1438 (N_1438,In_479,In_41);
or U1439 (N_1439,In_1554,In_1784);
nor U1440 (N_1440,In_763,In_904);
or U1441 (N_1441,In_738,In_355);
nor U1442 (N_1442,In_766,In_302);
xnor U1443 (N_1443,In_210,In_601);
nand U1444 (N_1444,In_34,In_1372);
or U1445 (N_1445,In_1581,In_143);
nand U1446 (N_1446,In_1482,In_1014);
nor U1447 (N_1447,In_1696,In_1702);
or U1448 (N_1448,In_1852,In_328);
or U1449 (N_1449,In_1888,In_1660);
and U1450 (N_1450,In_106,In_579);
nand U1451 (N_1451,In_824,In_402);
nand U1452 (N_1452,In_1517,In_891);
nor U1453 (N_1453,In_1000,In_689);
nand U1454 (N_1454,In_1785,In_543);
nand U1455 (N_1455,In_1292,In_1151);
nand U1456 (N_1456,In_1000,In_1298);
and U1457 (N_1457,In_1952,In_1877);
and U1458 (N_1458,In_1662,In_1425);
and U1459 (N_1459,In_1155,In_120);
or U1460 (N_1460,In_1597,In_1327);
or U1461 (N_1461,In_476,In_112);
nor U1462 (N_1462,In_693,In_823);
nor U1463 (N_1463,In_1728,In_1621);
nor U1464 (N_1464,In_982,In_9);
and U1465 (N_1465,In_1653,In_737);
and U1466 (N_1466,In_338,In_1670);
nor U1467 (N_1467,In_206,In_858);
nand U1468 (N_1468,In_1045,In_1781);
nand U1469 (N_1469,In_728,In_1232);
and U1470 (N_1470,In_197,In_470);
or U1471 (N_1471,In_1991,In_1049);
or U1472 (N_1472,In_1255,In_743);
or U1473 (N_1473,In_395,In_1362);
nor U1474 (N_1474,In_1542,In_1103);
and U1475 (N_1475,In_1343,In_272);
and U1476 (N_1476,In_325,In_1073);
nand U1477 (N_1477,In_1714,In_1390);
or U1478 (N_1478,In_410,In_1115);
or U1479 (N_1479,In_1261,In_1475);
and U1480 (N_1480,In_1506,In_546);
nor U1481 (N_1481,In_1949,In_1196);
or U1482 (N_1482,In_435,In_1024);
or U1483 (N_1483,In_400,In_1301);
or U1484 (N_1484,In_1650,In_723);
or U1485 (N_1485,In_1893,In_63);
and U1486 (N_1486,In_1951,In_229);
nor U1487 (N_1487,In_164,In_1389);
nand U1488 (N_1488,In_455,In_1616);
nand U1489 (N_1489,In_1244,In_227);
or U1490 (N_1490,In_335,In_1963);
xor U1491 (N_1491,In_1794,In_303);
xor U1492 (N_1492,In_596,In_1468);
xnor U1493 (N_1493,In_31,In_546);
and U1494 (N_1494,In_1223,In_992);
or U1495 (N_1495,In_1128,In_1396);
and U1496 (N_1496,In_1153,In_1797);
nor U1497 (N_1497,In_1648,In_1288);
nor U1498 (N_1498,In_1287,In_672);
nand U1499 (N_1499,In_934,In_1826);
and U1500 (N_1500,In_625,In_109);
and U1501 (N_1501,In_30,In_610);
and U1502 (N_1502,In_443,In_868);
xor U1503 (N_1503,In_938,In_1686);
and U1504 (N_1504,In_198,In_1631);
or U1505 (N_1505,In_879,In_330);
nor U1506 (N_1506,In_1101,In_1108);
or U1507 (N_1507,In_556,In_1040);
and U1508 (N_1508,In_489,In_1302);
nand U1509 (N_1509,In_1242,In_1148);
and U1510 (N_1510,In_547,In_1785);
nor U1511 (N_1511,In_1774,In_666);
and U1512 (N_1512,In_775,In_1844);
or U1513 (N_1513,In_864,In_348);
and U1514 (N_1514,In_1186,In_1340);
and U1515 (N_1515,In_1964,In_1104);
nor U1516 (N_1516,In_1647,In_73);
nor U1517 (N_1517,In_813,In_1027);
nand U1518 (N_1518,In_1517,In_227);
nor U1519 (N_1519,In_940,In_1967);
and U1520 (N_1520,In_388,In_867);
nor U1521 (N_1521,In_1087,In_1904);
and U1522 (N_1522,In_1435,In_570);
or U1523 (N_1523,In_747,In_263);
nand U1524 (N_1524,In_1387,In_1667);
nand U1525 (N_1525,In_1656,In_1166);
or U1526 (N_1526,In_972,In_1532);
or U1527 (N_1527,In_522,In_18);
and U1528 (N_1528,In_119,In_1781);
nor U1529 (N_1529,In_1841,In_168);
xnor U1530 (N_1530,In_153,In_105);
and U1531 (N_1531,In_2,In_1181);
nor U1532 (N_1532,In_171,In_1000);
nor U1533 (N_1533,In_1412,In_681);
or U1534 (N_1534,In_309,In_1212);
nor U1535 (N_1535,In_1723,In_1154);
nor U1536 (N_1536,In_1180,In_320);
or U1537 (N_1537,In_1360,In_1573);
nor U1538 (N_1538,In_1677,In_335);
or U1539 (N_1539,In_885,In_854);
or U1540 (N_1540,In_1706,In_1583);
nor U1541 (N_1541,In_781,In_1626);
xnor U1542 (N_1542,In_80,In_1219);
and U1543 (N_1543,In_520,In_1118);
nand U1544 (N_1544,In_624,In_394);
and U1545 (N_1545,In_1331,In_1469);
and U1546 (N_1546,In_1746,In_239);
or U1547 (N_1547,In_1210,In_37);
nand U1548 (N_1548,In_718,In_786);
nor U1549 (N_1549,In_252,In_68);
nor U1550 (N_1550,In_1407,In_279);
or U1551 (N_1551,In_733,In_1705);
and U1552 (N_1552,In_1239,In_153);
or U1553 (N_1553,In_51,In_898);
nand U1554 (N_1554,In_959,In_1398);
nor U1555 (N_1555,In_1511,In_1205);
or U1556 (N_1556,In_102,In_1673);
nor U1557 (N_1557,In_514,In_1501);
or U1558 (N_1558,In_1311,In_1931);
nor U1559 (N_1559,In_917,In_876);
or U1560 (N_1560,In_1430,In_1406);
nand U1561 (N_1561,In_64,In_87);
xnor U1562 (N_1562,In_891,In_1006);
nand U1563 (N_1563,In_785,In_220);
xor U1564 (N_1564,In_1752,In_670);
and U1565 (N_1565,In_767,In_1309);
or U1566 (N_1566,In_1091,In_78);
nand U1567 (N_1567,In_1449,In_1227);
and U1568 (N_1568,In_785,In_459);
and U1569 (N_1569,In_1649,In_1570);
and U1570 (N_1570,In_534,In_944);
and U1571 (N_1571,In_494,In_535);
nor U1572 (N_1572,In_446,In_269);
and U1573 (N_1573,In_637,In_1827);
nor U1574 (N_1574,In_1968,In_157);
nor U1575 (N_1575,In_1009,In_1049);
and U1576 (N_1576,In_50,In_1977);
nand U1577 (N_1577,In_357,In_622);
and U1578 (N_1578,In_1708,In_1119);
or U1579 (N_1579,In_1784,In_1701);
nand U1580 (N_1580,In_590,In_1463);
or U1581 (N_1581,In_460,In_386);
and U1582 (N_1582,In_595,In_1814);
nor U1583 (N_1583,In_135,In_807);
nor U1584 (N_1584,In_244,In_790);
or U1585 (N_1585,In_339,In_1128);
nand U1586 (N_1586,In_412,In_1411);
or U1587 (N_1587,In_401,In_450);
nor U1588 (N_1588,In_1393,In_860);
nand U1589 (N_1589,In_1528,In_53);
nor U1590 (N_1590,In_379,In_1888);
nor U1591 (N_1591,In_514,In_970);
or U1592 (N_1592,In_1172,In_894);
nand U1593 (N_1593,In_848,In_1407);
nor U1594 (N_1594,In_1834,In_1044);
nand U1595 (N_1595,In_645,In_1999);
and U1596 (N_1596,In_221,In_1090);
nand U1597 (N_1597,In_112,In_403);
and U1598 (N_1598,In_1117,In_1860);
nor U1599 (N_1599,In_537,In_1843);
and U1600 (N_1600,In_1808,In_342);
nor U1601 (N_1601,In_1142,In_912);
nand U1602 (N_1602,In_573,In_1867);
nor U1603 (N_1603,In_1726,In_247);
xor U1604 (N_1604,In_520,In_1881);
nor U1605 (N_1605,In_421,In_737);
nand U1606 (N_1606,In_581,In_1900);
nand U1607 (N_1607,In_452,In_1556);
and U1608 (N_1608,In_1908,In_1289);
nor U1609 (N_1609,In_1372,In_638);
and U1610 (N_1610,In_1236,In_24);
and U1611 (N_1611,In_259,In_231);
nor U1612 (N_1612,In_1657,In_151);
nand U1613 (N_1613,In_1798,In_808);
or U1614 (N_1614,In_724,In_1921);
nor U1615 (N_1615,In_407,In_1516);
nor U1616 (N_1616,In_371,In_766);
nor U1617 (N_1617,In_307,In_553);
or U1618 (N_1618,In_1954,In_590);
or U1619 (N_1619,In_797,In_1551);
nor U1620 (N_1620,In_458,In_916);
and U1621 (N_1621,In_678,In_1933);
or U1622 (N_1622,In_996,In_1472);
or U1623 (N_1623,In_1423,In_1830);
nor U1624 (N_1624,In_1804,In_1787);
or U1625 (N_1625,In_172,In_1093);
and U1626 (N_1626,In_1020,In_1182);
nand U1627 (N_1627,In_557,In_1786);
or U1628 (N_1628,In_1423,In_1837);
or U1629 (N_1629,In_1827,In_1985);
and U1630 (N_1630,In_1626,In_825);
nor U1631 (N_1631,In_1052,In_409);
nand U1632 (N_1632,In_1157,In_627);
nand U1633 (N_1633,In_640,In_1218);
and U1634 (N_1634,In_415,In_483);
nand U1635 (N_1635,In_1074,In_1069);
nor U1636 (N_1636,In_603,In_1724);
nor U1637 (N_1637,In_1600,In_401);
nand U1638 (N_1638,In_750,In_1727);
or U1639 (N_1639,In_862,In_549);
nand U1640 (N_1640,In_368,In_1684);
nor U1641 (N_1641,In_1435,In_1331);
and U1642 (N_1642,In_337,In_907);
and U1643 (N_1643,In_528,In_1100);
or U1644 (N_1644,In_1387,In_645);
or U1645 (N_1645,In_562,In_763);
and U1646 (N_1646,In_123,In_1762);
or U1647 (N_1647,In_1771,In_374);
and U1648 (N_1648,In_1271,In_579);
nor U1649 (N_1649,In_1774,In_1284);
and U1650 (N_1650,In_1027,In_1746);
nand U1651 (N_1651,In_1431,In_268);
or U1652 (N_1652,In_1564,In_1572);
nor U1653 (N_1653,In_704,In_347);
nand U1654 (N_1654,In_16,In_995);
nand U1655 (N_1655,In_1965,In_545);
nand U1656 (N_1656,In_909,In_1492);
nand U1657 (N_1657,In_732,In_757);
and U1658 (N_1658,In_1095,In_1637);
nor U1659 (N_1659,In_1995,In_1448);
or U1660 (N_1660,In_991,In_1924);
nand U1661 (N_1661,In_1057,In_1768);
or U1662 (N_1662,In_1624,In_1707);
and U1663 (N_1663,In_1750,In_907);
nor U1664 (N_1664,In_606,In_1930);
or U1665 (N_1665,In_1435,In_84);
nand U1666 (N_1666,In_570,In_440);
or U1667 (N_1667,In_435,In_587);
nor U1668 (N_1668,In_1636,In_1119);
or U1669 (N_1669,In_1272,In_1484);
or U1670 (N_1670,In_408,In_697);
nor U1671 (N_1671,In_517,In_154);
or U1672 (N_1672,In_1416,In_1497);
nand U1673 (N_1673,In_918,In_1547);
nand U1674 (N_1674,In_1546,In_1323);
and U1675 (N_1675,In_251,In_1790);
xnor U1676 (N_1676,In_1124,In_944);
or U1677 (N_1677,In_1165,In_1384);
or U1678 (N_1678,In_1618,In_806);
and U1679 (N_1679,In_303,In_1970);
nor U1680 (N_1680,In_19,In_972);
or U1681 (N_1681,In_320,In_328);
and U1682 (N_1682,In_334,In_1760);
or U1683 (N_1683,In_1125,In_848);
or U1684 (N_1684,In_1745,In_1701);
nor U1685 (N_1685,In_1419,In_357);
nor U1686 (N_1686,In_1422,In_334);
nor U1687 (N_1687,In_840,In_1894);
nand U1688 (N_1688,In_1421,In_1407);
nor U1689 (N_1689,In_1430,In_429);
nor U1690 (N_1690,In_437,In_1589);
nor U1691 (N_1691,In_260,In_121);
nor U1692 (N_1692,In_1477,In_1383);
nand U1693 (N_1693,In_1709,In_1361);
and U1694 (N_1694,In_495,In_436);
or U1695 (N_1695,In_1012,In_78);
or U1696 (N_1696,In_1568,In_1077);
or U1697 (N_1697,In_1009,In_1716);
nand U1698 (N_1698,In_1045,In_417);
and U1699 (N_1699,In_776,In_1331);
nor U1700 (N_1700,In_190,In_398);
and U1701 (N_1701,In_490,In_1965);
and U1702 (N_1702,In_451,In_557);
nand U1703 (N_1703,In_426,In_1293);
nor U1704 (N_1704,In_1375,In_1556);
or U1705 (N_1705,In_1240,In_867);
nand U1706 (N_1706,In_1629,In_1595);
or U1707 (N_1707,In_912,In_1525);
and U1708 (N_1708,In_796,In_145);
or U1709 (N_1709,In_204,In_1982);
nor U1710 (N_1710,In_1872,In_381);
nor U1711 (N_1711,In_966,In_1252);
nor U1712 (N_1712,In_819,In_1634);
xnor U1713 (N_1713,In_736,In_1543);
and U1714 (N_1714,In_1984,In_1539);
nand U1715 (N_1715,In_1322,In_1415);
and U1716 (N_1716,In_259,In_1768);
and U1717 (N_1717,In_684,In_640);
nand U1718 (N_1718,In_706,In_576);
nor U1719 (N_1719,In_528,In_1781);
nand U1720 (N_1720,In_1410,In_1611);
and U1721 (N_1721,In_57,In_1420);
and U1722 (N_1722,In_1013,In_272);
and U1723 (N_1723,In_1853,In_1184);
and U1724 (N_1724,In_1340,In_1267);
nor U1725 (N_1725,In_270,In_1308);
or U1726 (N_1726,In_1899,In_1916);
or U1727 (N_1727,In_1727,In_1127);
and U1728 (N_1728,In_352,In_495);
or U1729 (N_1729,In_1635,In_627);
nand U1730 (N_1730,In_167,In_512);
nand U1731 (N_1731,In_49,In_1154);
nand U1732 (N_1732,In_1197,In_1809);
nand U1733 (N_1733,In_928,In_1795);
nand U1734 (N_1734,In_428,In_484);
or U1735 (N_1735,In_388,In_1237);
nor U1736 (N_1736,In_359,In_1775);
nor U1737 (N_1737,In_785,In_1768);
or U1738 (N_1738,In_716,In_862);
and U1739 (N_1739,In_41,In_1800);
nor U1740 (N_1740,In_1254,In_1824);
nor U1741 (N_1741,In_1058,In_617);
nand U1742 (N_1742,In_1964,In_403);
nand U1743 (N_1743,In_1624,In_861);
or U1744 (N_1744,In_1639,In_401);
and U1745 (N_1745,In_1479,In_342);
or U1746 (N_1746,In_36,In_1062);
nor U1747 (N_1747,In_1351,In_49);
nand U1748 (N_1748,In_1398,In_1312);
and U1749 (N_1749,In_1515,In_123);
and U1750 (N_1750,In_970,In_716);
or U1751 (N_1751,In_708,In_949);
and U1752 (N_1752,In_778,In_1701);
or U1753 (N_1753,In_1042,In_563);
nand U1754 (N_1754,In_202,In_1203);
nor U1755 (N_1755,In_8,In_1930);
and U1756 (N_1756,In_1642,In_539);
nand U1757 (N_1757,In_1557,In_1269);
or U1758 (N_1758,In_1574,In_1583);
or U1759 (N_1759,In_414,In_1417);
nor U1760 (N_1760,In_320,In_88);
and U1761 (N_1761,In_889,In_179);
nor U1762 (N_1762,In_1201,In_1290);
nand U1763 (N_1763,In_1913,In_1271);
nand U1764 (N_1764,In_125,In_127);
or U1765 (N_1765,In_311,In_723);
nand U1766 (N_1766,In_1,In_1613);
nand U1767 (N_1767,In_858,In_777);
or U1768 (N_1768,In_784,In_1993);
and U1769 (N_1769,In_35,In_444);
or U1770 (N_1770,In_1992,In_548);
nor U1771 (N_1771,In_1020,In_965);
nor U1772 (N_1772,In_1254,In_625);
xnor U1773 (N_1773,In_529,In_1421);
or U1774 (N_1774,In_991,In_112);
and U1775 (N_1775,In_1108,In_525);
and U1776 (N_1776,In_479,In_1797);
nor U1777 (N_1777,In_21,In_1606);
nor U1778 (N_1778,In_1945,In_268);
or U1779 (N_1779,In_1031,In_1532);
and U1780 (N_1780,In_337,In_1919);
nand U1781 (N_1781,In_4,In_13);
nor U1782 (N_1782,In_519,In_1820);
and U1783 (N_1783,In_413,In_361);
and U1784 (N_1784,In_570,In_1735);
nor U1785 (N_1785,In_919,In_1790);
and U1786 (N_1786,In_1038,In_18);
nor U1787 (N_1787,In_372,In_766);
and U1788 (N_1788,In_692,In_1341);
nor U1789 (N_1789,In_1355,In_1394);
nand U1790 (N_1790,In_1855,In_1845);
and U1791 (N_1791,In_265,In_1897);
nand U1792 (N_1792,In_299,In_344);
nor U1793 (N_1793,In_380,In_335);
nand U1794 (N_1794,In_354,In_1517);
and U1795 (N_1795,In_1111,In_1447);
nand U1796 (N_1796,In_1567,In_1629);
nor U1797 (N_1797,In_520,In_952);
and U1798 (N_1798,In_7,In_1489);
nor U1799 (N_1799,In_1059,In_580);
or U1800 (N_1800,In_1486,In_790);
and U1801 (N_1801,In_647,In_1613);
and U1802 (N_1802,In_50,In_881);
nor U1803 (N_1803,In_1818,In_134);
nand U1804 (N_1804,In_804,In_816);
nor U1805 (N_1805,In_1362,In_1160);
nand U1806 (N_1806,In_1869,In_236);
and U1807 (N_1807,In_576,In_815);
nor U1808 (N_1808,In_739,In_1064);
nor U1809 (N_1809,In_175,In_158);
nor U1810 (N_1810,In_447,In_428);
or U1811 (N_1811,In_630,In_1792);
nand U1812 (N_1812,In_1565,In_1526);
nor U1813 (N_1813,In_407,In_1173);
nor U1814 (N_1814,In_1556,In_733);
or U1815 (N_1815,In_1638,In_1233);
nand U1816 (N_1816,In_1305,In_395);
or U1817 (N_1817,In_723,In_1970);
or U1818 (N_1818,In_1720,In_1464);
nand U1819 (N_1819,In_908,In_610);
and U1820 (N_1820,In_584,In_582);
xnor U1821 (N_1821,In_1212,In_1807);
nand U1822 (N_1822,In_1235,In_697);
nand U1823 (N_1823,In_345,In_1558);
or U1824 (N_1824,In_116,In_38);
nand U1825 (N_1825,In_1672,In_241);
and U1826 (N_1826,In_382,In_1103);
or U1827 (N_1827,In_779,In_1363);
and U1828 (N_1828,In_834,In_698);
and U1829 (N_1829,In_522,In_1390);
nand U1830 (N_1830,In_1245,In_559);
nand U1831 (N_1831,In_480,In_1353);
and U1832 (N_1832,In_568,In_1437);
nand U1833 (N_1833,In_12,In_91);
nand U1834 (N_1834,In_1754,In_1375);
nand U1835 (N_1835,In_230,In_1467);
nand U1836 (N_1836,In_174,In_201);
nor U1837 (N_1837,In_1446,In_1913);
or U1838 (N_1838,In_1638,In_1063);
nand U1839 (N_1839,In_1611,In_1752);
nand U1840 (N_1840,In_1018,In_804);
and U1841 (N_1841,In_1015,In_264);
nor U1842 (N_1842,In_97,In_866);
nor U1843 (N_1843,In_200,In_1534);
or U1844 (N_1844,In_503,In_1296);
nand U1845 (N_1845,In_725,In_1096);
or U1846 (N_1846,In_1233,In_1652);
and U1847 (N_1847,In_1172,In_867);
and U1848 (N_1848,In_1395,In_1971);
or U1849 (N_1849,In_1904,In_47);
and U1850 (N_1850,In_1413,In_1559);
nor U1851 (N_1851,In_1916,In_1557);
and U1852 (N_1852,In_674,In_197);
or U1853 (N_1853,In_1968,In_867);
nor U1854 (N_1854,In_229,In_542);
or U1855 (N_1855,In_1310,In_846);
nor U1856 (N_1856,In_363,In_1343);
or U1857 (N_1857,In_1723,In_0);
and U1858 (N_1858,In_1430,In_164);
nor U1859 (N_1859,In_759,In_1467);
or U1860 (N_1860,In_258,In_761);
and U1861 (N_1861,In_1056,In_702);
or U1862 (N_1862,In_1037,In_744);
nand U1863 (N_1863,In_1150,In_89);
nor U1864 (N_1864,In_939,In_1122);
nand U1865 (N_1865,In_1210,In_1602);
and U1866 (N_1866,In_1957,In_773);
and U1867 (N_1867,In_61,In_473);
nor U1868 (N_1868,In_1438,In_867);
nor U1869 (N_1869,In_985,In_1971);
and U1870 (N_1870,In_781,In_1945);
and U1871 (N_1871,In_1666,In_779);
and U1872 (N_1872,In_1463,In_1181);
and U1873 (N_1873,In_1523,In_166);
and U1874 (N_1874,In_1494,In_1665);
or U1875 (N_1875,In_1313,In_402);
nand U1876 (N_1876,In_964,In_309);
nor U1877 (N_1877,In_254,In_938);
nor U1878 (N_1878,In_1449,In_79);
and U1879 (N_1879,In_1017,In_1369);
and U1880 (N_1880,In_1430,In_1266);
and U1881 (N_1881,In_523,In_798);
nor U1882 (N_1882,In_1012,In_518);
or U1883 (N_1883,In_1276,In_1574);
nand U1884 (N_1884,In_416,In_926);
and U1885 (N_1885,In_870,In_786);
xor U1886 (N_1886,In_823,In_1977);
nand U1887 (N_1887,In_917,In_1213);
nand U1888 (N_1888,In_1448,In_756);
nand U1889 (N_1889,In_404,In_1451);
nand U1890 (N_1890,In_1510,In_1038);
nor U1891 (N_1891,In_1726,In_1624);
nor U1892 (N_1892,In_1883,In_1199);
and U1893 (N_1893,In_1584,In_1464);
nand U1894 (N_1894,In_1624,In_1883);
and U1895 (N_1895,In_101,In_127);
nor U1896 (N_1896,In_164,In_819);
nor U1897 (N_1897,In_1752,In_252);
or U1898 (N_1898,In_1745,In_867);
nor U1899 (N_1899,In_1096,In_1661);
nand U1900 (N_1900,In_1629,In_1018);
nor U1901 (N_1901,In_1353,In_1328);
nor U1902 (N_1902,In_632,In_1894);
nor U1903 (N_1903,In_1838,In_1779);
and U1904 (N_1904,In_104,In_1980);
nor U1905 (N_1905,In_1561,In_1289);
and U1906 (N_1906,In_1200,In_1869);
or U1907 (N_1907,In_1191,In_1355);
nor U1908 (N_1908,In_471,In_1221);
and U1909 (N_1909,In_390,In_1178);
nand U1910 (N_1910,In_1688,In_320);
and U1911 (N_1911,In_733,In_268);
and U1912 (N_1912,In_575,In_1124);
or U1913 (N_1913,In_1592,In_813);
or U1914 (N_1914,In_919,In_1233);
nand U1915 (N_1915,In_1567,In_906);
nand U1916 (N_1916,In_1116,In_1432);
nor U1917 (N_1917,In_1434,In_1653);
and U1918 (N_1918,In_1234,In_1866);
and U1919 (N_1919,In_311,In_453);
nor U1920 (N_1920,In_114,In_601);
and U1921 (N_1921,In_1095,In_747);
nor U1922 (N_1922,In_805,In_1926);
nand U1923 (N_1923,In_464,In_1244);
nor U1924 (N_1924,In_1559,In_163);
nor U1925 (N_1925,In_89,In_1217);
and U1926 (N_1926,In_1715,In_76);
nand U1927 (N_1927,In_1204,In_363);
or U1928 (N_1928,In_1528,In_742);
and U1929 (N_1929,In_171,In_1988);
or U1930 (N_1930,In_218,In_613);
and U1931 (N_1931,In_1935,In_1948);
nand U1932 (N_1932,In_1927,In_799);
or U1933 (N_1933,In_387,In_1892);
nor U1934 (N_1934,In_717,In_1010);
and U1935 (N_1935,In_678,In_1615);
or U1936 (N_1936,In_1733,In_1255);
and U1937 (N_1937,In_1841,In_610);
or U1938 (N_1938,In_544,In_1591);
or U1939 (N_1939,In_77,In_601);
and U1940 (N_1940,In_436,In_613);
and U1941 (N_1941,In_1185,In_288);
and U1942 (N_1942,In_985,In_1864);
nor U1943 (N_1943,In_1532,In_1332);
or U1944 (N_1944,In_1014,In_256);
or U1945 (N_1945,In_1761,In_1531);
xor U1946 (N_1946,In_1108,In_1441);
and U1947 (N_1947,In_1,In_1780);
nand U1948 (N_1948,In_597,In_1215);
and U1949 (N_1949,In_328,In_711);
nor U1950 (N_1950,In_394,In_623);
or U1951 (N_1951,In_364,In_231);
nor U1952 (N_1952,In_1100,In_799);
or U1953 (N_1953,In_729,In_1367);
nand U1954 (N_1954,In_1381,In_335);
or U1955 (N_1955,In_1168,In_1703);
or U1956 (N_1956,In_75,In_1017);
or U1957 (N_1957,In_277,In_1112);
or U1958 (N_1958,In_1620,In_1951);
nor U1959 (N_1959,In_993,In_72);
nand U1960 (N_1960,In_1101,In_1420);
nand U1961 (N_1961,In_441,In_852);
or U1962 (N_1962,In_1660,In_312);
or U1963 (N_1963,In_243,In_594);
or U1964 (N_1964,In_1617,In_226);
or U1965 (N_1965,In_1595,In_1027);
xor U1966 (N_1966,In_1989,In_35);
nand U1967 (N_1967,In_1429,In_1474);
nand U1968 (N_1968,In_1318,In_295);
and U1969 (N_1969,In_1751,In_1468);
nand U1970 (N_1970,In_1235,In_1315);
and U1971 (N_1971,In_457,In_738);
nand U1972 (N_1972,In_1275,In_572);
or U1973 (N_1973,In_809,In_491);
or U1974 (N_1974,In_1888,In_1179);
and U1975 (N_1975,In_964,In_19);
and U1976 (N_1976,In_1211,In_1857);
nor U1977 (N_1977,In_555,In_1565);
nor U1978 (N_1978,In_1954,In_953);
nand U1979 (N_1979,In_868,In_1627);
nor U1980 (N_1980,In_373,In_715);
nor U1981 (N_1981,In_1930,In_1117);
xor U1982 (N_1982,In_1031,In_244);
or U1983 (N_1983,In_1115,In_639);
or U1984 (N_1984,In_1666,In_1266);
or U1985 (N_1985,In_295,In_8);
nand U1986 (N_1986,In_1733,In_1161);
or U1987 (N_1987,In_958,In_1362);
nor U1988 (N_1988,In_1365,In_893);
xor U1989 (N_1989,In_1368,In_1665);
and U1990 (N_1990,In_1257,In_1600);
or U1991 (N_1991,In_1267,In_1136);
and U1992 (N_1992,In_1427,In_1661);
nor U1993 (N_1993,In_614,In_1615);
or U1994 (N_1994,In_1159,In_1421);
and U1995 (N_1995,In_1427,In_111);
nor U1996 (N_1996,In_1410,In_1269);
and U1997 (N_1997,In_1982,In_456);
and U1998 (N_1998,In_352,In_1566);
xor U1999 (N_1999,In_1587,In_235);
nand U2000 (N_2000,In_1801,In_72);
nand U2001 (N_2001,In_1258,In_19);
nor U2002 (N_2002,In_1360,In_1415);
and U2003 (N_2003,In_517,In_926);
and U2004 (N_2004,In_938,In_727);
nor U2005 (N_2005,In_643,In_1377);
xnor U2006 (N_2006,In_262,In_1507);
or U2007 (N_2007,In_1242,In_691);
or U2008 (N_2008,In_1910,In_1906);
nor U2009 (N_2009,In_327,In_1383);
nand U2010 (N_2010,In_90,In_201);
nand U2011 (N_2011,In_552,In_852);
and U2012 (N_2012,In_1270,In_1436);
nor U2013 (N_2013,In_1751,In_192);
and U2014 (N_2014,In_926,In_1011);
and U2015 (N_2015,In_1106,In_1599);
nand U2016 (N_2016,In_1700,In_1645);
nand U2017 (N_2017,In_564,In_128);
and U2018 (N_2018,In_1920,In_837);
or U2019 (N_2019,In_21,In_1681);
nor U2020 (N_2020,In_398,In_306);
or U2021 (N_2021,In_1955,In_96);
or U2022 (N_2022,In_1149,In_652);
or U2023 (N_2023,In_1817,In_761);
nand U2024 (N_2024,In_478,In_1542);
nor U2025 (N_2025,In_772,In_1981);
nor U2026 (N_2026,In_1910,In_1159);
nor U2027 (N_2027,In_1101,In_1986);
nand U2028 (N_2028,In_521,In_1932);
and U2029 (N_2029,In_854,In_916);
or U2030 (N_2030,In_1880,In_1092);
and U2031 (N_2031,In_1841,In_175);
or U2032 (N_2032,In_1886,In_640);
nand U2033 (N_2033,In_948,In_546);
and U2034 (N_2034,In_1748,In_70);
nand U2035 (N_2035,In_438,In_755);
nand U2036 (N_2036,In_1603,In_20);
nand U2037 (N_2037,In_244,In_1856);
or U2038 (N_2038,In_827,In_724);
or U2039 (N_2039,In_1095,In_1953);
and U2040 (N_2040,In_361,In_730);
and U2041 (N_2041,In_1934,In_990);
nand U2042 (N_2042,In_691,In_1304);
and U2043 (N_2043,In_147,In_24);
or U2044 (N_2044,In_481,In_726);
or U2045 (N_2045,In_881,In_1411);
or U2046 (N_2046,In_787,In_1891);
and U2047 (N_2047,In_323,In_531);
nor U2048 (N_2048,In_211,In_1970);
nor U2049 (N_2049,In_699,In_40);
nand U2050 (N_2050,In_751,In_1209);
or U2051 (N_2051,In_685,In_1261);
or U2052 (N_2052,In_699,In_1858);
nor U2053 (N_2053,In_970,In_207);
or U2054 (N_2054,In_461,In_899);
and U2055 (N_2055,In_1062,In_1958);
and U2056 (N_2056,In_404,In_521);
nand U2057 (N_2057,In_1083,In_1267);
and U2058 (N_2058,In_1297,In_1151);
nand U2059 (N_2059,In_1964,In_1155);
xor U2060 (N_2060,In_969,In_359);
or U2061 (N_2061,In_1015,In_947);
xor U2062 (N_2062,In_457,In_1253);
or U2063 (N_2063,In_797,In_1881);
nor U2064 (N_2064,In_1581,In_1552);
and U2065 (N_2065,In_1758,In_399);
or U2066 (N_2066,In_114,In_1846);
xor U2067 (N_2067,In_1811,In_769);
or U2068 (N_2068,In_268,In_496);
nand U2069 (N_2069,In_1652,In_1010);
or U2070 (N_2070,In_1660,In_1110);
nor U2071 (N_2071,In_937,In_1030);
or U2072 (N_2072,In_338,In_577);
and U2073 (N_2073,In_850,In_1017);
nand U2074 (N_2074,In_483,In_1618);
and U2075 (N_2075,In_1556,In_1884);
nor U2076 (N_2076,In_329,In_578);
and U2077 (N_2077,In_773,In_1317);
nor U2078 (N_2078,In_1804,In_1091);
or U2079 (N_2079,In_998,In_1347);
or U2080 (N_2080,In_274,In_1089);
nor U2081 (N_2081,In_931,In_66);
and U2082 (N_2082,In_250,In_417);
or U2083 (N_2083,In_1355,In_926);
nand U2084 (N_2084,In_952,In_958);
nand U2085 (N_2085,In_1296,In_409);
nor U2086 (N_2086,In_1905,In_1066);
or U2087 (N_2087,In_1233,In_1062);
and U2088 (N_2088,In_1192,In_550);
nand U2089 (N_2089,In_1421,In_1251);
and U2090 (N_2090,In_616,In_887);
nor U2091 (N_2091,In_1530,In_1927);
and U2092 (N_2092,In_1157,In_1977);
or U2093 (N_2093,In_1905,In_130);
or U2094 (N_2094,In_466,In_1161);
nand U2095 (N_2095,In_219,In_1402);
or U2096 (N_2096,In_1454,In_504);
and U2097 (N_2097,In_1657,In_809);
or U2098 (N_2098,In_1714,In_1299);
and U2099 (N_2099,In_1455,In_579);
or U2100 (N_2100,In_1107,In_1867);
or U2101 (N_2101,In_934,In_1623);
nor U2102 (N_2102,In_1817,In_108);
nor U2103 (N_2103,In_1288,In_551);
or U2104 (N_2104,In_208,In_1037);
nor U2105 (N_2105,In_1820,In_3);
and U2106 (N_2106,In_1094,In_346);
xor U2107 (N_2107,In_1668,In_1754);
or U2108 (N_2108,In_1466,In_1070);
and U2109 (N_2109,In_71,In_1429);
and U2110 (N_2110,In_1358,In_1566);
nor U2111 (N_2111,In_891,In_1397);
or U2112 (N_2112,In_73,In_783);
xor U2113 (N_2113,In_79,In_1075);
nor U2114 (N_2114,In_1277,In_1041);
nand U2115 (N_2115,In_991,In_149);
nor U2116 (N_2116,In_807,In_1199);
and U2117 (N_2117,In_1576,In_145);
nor U2118 (N_2118,In_356,In_454);
or U2119 (N_2119,In_4,In_530);
and U2120 (N_2120,In_870,In_1207);
nor U2121 (N_2121,In_777,In_1986);
or U2122 (N_2122,In_1475,In_1083);
nor U2123 (N_2123,In_1987,In_1355);
nand U2124 (N_2124,In_1695,In_1283);
and U2125 (N_2125,In_283,In_156);
nor U2126 (N_2126,In_1455,In_153);
nor U2127 (N_2127,In_1741,In_71);
xor U2128 (N_2128,In_1763,In_1790);
or U2129 (N_2129,In_908,In_1972);
and U2130 (N_2130,In_370,In_1262);
nor U2131 (N_2131,In_1244,In_593);
nand U2132 (N_2132,In_894,In_670);
or U2133 (N_2133,In_1926,In_1641);
or U2134 (N_2134,In_1269,In_642);
nand U2135 (N_2135,In_862,In_325);
and U2136 (N_2136,In_229,In_270);
or U2137 (N_2137,In_1537,In_1300);
nand U2138 (N_2138,In_22,In_1830);
or U2139 (N_2139,In_1115,In_703);
nand U2140 (N_2140,In_88,In_1462);
nand U2141 (N_2141,In_418,In_1227);
or U2142 (N_2142,In_1806,In_306);
nor U2143 (N_2143,In_1590,In_1753);
nand U2144 (N_2144,In_89,In_519);
nor U2145 (N_2145,In_369,In_1428);
nand U2146 (N_2146,In_952,In_614);
or U2147 (N_2147,In_1695,In_1737);
nand U2148 (N_2148,In_1028,In_341);
nand U2149 (N_2149,In_453,In_607);
or U2150 (N_2150,In_179,In_1079);
and U2151 (N_2151,In_515,In_641);
and U2152 (N_2152,In_1036,In_286);
nor U2153 (N_2153,In_810,In_1184);
and U2154 (N_2154,In_1828,In_490);
nor U2155 (N_2155,In_449,In_597);
and U2156 (N_2156,In_80,In_375);
nor U2157 (N_2157,In_174,In_1856);
and U2158 (N_2158,In_552,In_1845);
or U2159 (N_2159,In_978,In_832);
or U2160 (N_2160,In_12,In_261);
and U2161 (N_2161,In_269,In_810);
or U2162 (N_2162,In_353,In_183);
or U2163 (N_2163,In_993,In_400);
nor U2164 (N_2164,In_1539,In_51);
and U2165 (N_2165,In_529,In_1022);
nand U2166 (N_2166,In_1489,In_1025);
or U2167 (N_2167,In_1283,In_1285);
or U2168 (N_2168,In_1412,In_546);
or U2169 (N_2169,In_1113,In_943);
nand U2170 (N_2170,In_1203,In_1152);
or U2171 (N_2171,In_148,In_1236);
or U2172 (N_2172,In_957,In_1781);
nor U2173 (N_2173,In_280,In_416);
or U2174 (N_2174,In_177,In_1890);
nand U2175 (N_2175,In_499,In_1215);
or U2176 (N_2176,In_1808,In_1030);
or U2177 (N_2177,In_1152,In_27);
nor U2178 (N_2178,In_1364,In_1234);
nand U2179 (N_2179,In_232,In_521);
or U2180 (N_2180,In_1984,In_1628);
nor U2181 (N_2181,In_1878,In_1897);
nand U2182 (N_2182,In_555,In_1761);
and U2183 (N_2183,In_404,In_418);
and U2184 (N_2184,In_1151,In_351);
nor U2185 (N_2185,In_204,In_1672);
nand U2186 (N_2186,In_1066,In_88);
nand U2187 (N_2187,In_600,In_1579);
nand U2188 (N_2188,In_389,In_1067);
or U2189 (N_2189,In_1954,In_1544);
nor U2190 (N_2190,In_1551,In_1374);
or U2191 (N_2191,In_203,In_1724);
nor U2192 (N_2192,In_1893,In_330);
xor U2193 (N_2193,In_574,In_1751);
nand U2194 (N_2194,In_717,In_1799);
nand U2195 (N_2195,In_1632,In_1231);
nor U2196 (N_2196,In_1422,In_1388);
or U2197 (N_2197,In_1245,In_748);
or U2198 (N_2198,In_1864,In_1523);
xor U2199 (N_2199,In_906,In_3);
nand U2200 (N_2200,In_208,In_581);
nor U2201 (N_2201,In_1949,In_1815);
or U2202 (N_2202,In_587,In_1940);
nor U2203 (N_2203,In_681,In_1440);
and U2204 (N_2204,In_1281,In_1587);
or U2205 (N_2205,In_891,In_731);
or U2206 (N_2206,In_1255,In_812);
or U2207 (N_2207,In_1626,In_820);
nand U2208 (N_2208,In_737,In_1103);
and U2209 (N_2209,In_532,In_958);
nand U2210 (N_2210,In_565,In_1835);
nor U2211 (N_2211,In_1561,In_1795);
or U2212 (N_2212,In_1025,In_1276);
or U2213 (N_2213,In_930,In_574);
or U2214 (N_2214,In_1608,In_176);
or U2215 (N_2215,In_541,In_778);
nand U2216 (N_2216,In_1928,In_1662);
nor U2217 (N_2217,In_1640,In_1649);
nand U2218 (N_2218,In_1384,In_431);
nor U2219 (N_2219,In_769,In_1851);
nand U2220 (N_2220,In_361,In_1891);
and U2221 (N_2221,In_1368,In_1827);
nand U2222 (N_2222,In_1257,In_665);
or U2223 (N_2223,In_1396,In_1652);
nand U2224 (N_2224,In_1681,In_1733);
and U2225 (N_2225,In_540,In_1583);
or U2226 (N_2226,In_913,In_1009);
and U2227 (N_2227,In_1807,In_1514);
or U2228 (N_2228,In_575,In_1267);
or U2229 (N_2229,In_1390,In_172);
or U2230 (N_2230,In_789,In_792);
and U2231 (N_2231,In_1600,In_450);
nand U2232 (N_2232,In_470,In_77);
or U2233 (N_2233,In_1952,In_1277);
nand U2234 (N_2234,In_806,In_1947);
nor U2235 (N_2235,In_1242,In_1558);
and U2236 (N_2236,In_960,In_1263);
or U2237 (N_2237,In_1810,In_1431);
and U2238 (N_2238,In_1498,In_546);
or U2239 (N_2239,In_1269,In_710);
and U2240 (N_2240,In_1959,In_1849);
and U2241 (N_2241,In_1000,In_233);
and U2242 (N_2242,In_866,In_833);
xnor U2243 (N_2243,In_747,In_228);
nor U2244 (N_2244,In_1676,In_1674);
nor U2245 (N_2245,In_1626,In_983);
nor U2246 (N_2246,In_1622,In_643);
or U2247 (N_2247,In_698,In_1815);
nand U2248 (N_2248,In_1882,In_1542);
nand U2249 (N_2249,In_865,In_275);
nor U2250 (N_2250,In_798,In_1537);
nor U2251 (N_2251,In_644,In_1892);
and U2252 (N_2252,In_1187,In_777);
or U2253 (N_2253,In_1041,In_1675);
and U2254 (N_2254,In_1313,In_116);
nor U2255 (N_2255,In_259,In_1425);
nor U2256 (N_2256,In_517,In_903);
or U2257 (N_2257,In_913,In_1701);
nand U2258 (N_2258,In_417,In_1180);
and U2259 (N_2259,In_225,In_1422);
or U2260 (N_2260,In_1942,In_1848);
or U2261 (N_2261,In_1426,In_1238);
xnor U2262 (N_2262,In_890,In_1816);
or U2263 (N_2263,In_1717,In_751);
and U2264 (N_2264,In_618,In_319);
nand U2265 (N_2265,In_298,In_746);
nor U2266 (N_2266,In_471,In_821);
or U2267 (N_2267,In_298,In_987);
and U2268 (N_2268,In_954,In_1200);
or U2269 (N_2269,In_439,In_1146);
and U2270 (N_2270,In_1130,In_440);
nand U2271 (N_2271,In_717,In_1961);
nand U2272 (N_2272,In_1644,In_1510);
nand U2273 (N_2273,In_477,In_1601);
or U2274 (N_2274,In_947,In_1020);
and U2275 (N_2275,In_723,In_1895);
or U2276 (N_2276,In_1898,In_87);
nor U2277 (N_2277,In_1749,In_1924);
and U2278 (N_2278,In_1901,In_1926);
nor U2279 (N_2279,In_1054,In_106);
and U2280 (N_2280,In_1567,In_277);
and U2281 (N_2281,In_1328,In_222);
and U2282 (N_2282,In_301,In_989);
nor U2283 (N_2283,In_655,In_1149);
and U2284 (N_2284,In_832,In_1305);
or U2285 (N_2285,In_1066,In_610);
or U2286 (N_2286,In_74,In_1537);
xnor U2287 (N_2287,In_502,In_671);
nor U2288 (N_2288,In_1898,In_229);
nand U2289 (N_2289,In_1345,In_189);
or U2290 (N_2290,In_1396,In_1907);
nand U2291 (N_2291,In_1277,In_1155);
and U2292 (N_2292,In_1669,In_1371);
xor U2293 (N_2293,In_1452,In_1507);
nor U2294 (N_2294,In_1268,In_195);
and U2295 (N_2295,In_177,In_519);
nand U2296 (N_2296,In_353,In_1074);
and U2297 (N_2297,In_1077,In_808);
nor U2298 (N_2298,In_1297,In_1733);
nor U2299 (N_2299,In_730,In_488);
nand U2300 (N_2300,In_121,In_123);
or U2301 (N_2301,In_143,In_1763);
and U2302 (N_2302,In_573,In_964);
and U2303 (N_2303,In_1863,In_1970);
xor U2304 (N_2304,In_154,In_471);
or U2305 (N_2305,In_776,In_187);
and U2306 (N_2306,In_1229,In_1003);
nor U2307 (N_2307,In_170,In_670);
nor U2308 (N_2308,In_277,In_355);
nand U2309 (N_2309,In_1625,In_1500);
nand U2310 (N_2310,In_1340,In_1648);
xnor U2311 (N_2311,In_779,In_1991);
and U2312 (N_2312,In_1288,In_1012);
nand U2313 (N_2313,In_1615,In_965);
nand U2314 (N_2314,In_1062,In_1359);
nand U2315 (N_2315,In_1016,In_364);
or U2316 (N_2316,In_1877,In_1288);
nor U2317 (N_2317,In_152,In_1377);
nand U2318 (N_2318,In_893,In_508);
or U2319 (N_2319,In_22,In_369);
nand U2320 (N_2320,In_1413,In_1664);
and U2321 (N_2321,In_172,In_1559);
nand U2322 (N_2322,In_174,In_1520);
or U2323 (N_2323,In_1074,In_428);
and U2324 (N_2324,In_1239,In_429);
nor U2325 (N_2325,In_1761,In_139);
nand U2326 (N_2326,In_521,In_1197);
nand U2327 (N_2327,In_465,In_1218);
xnor U2328 (N_2328,In_1889,In_1828);
and U2329 (N_2329,In_1034,In_1298);
xor U2330 (N_2330,In_1147,In_1414);
or U2331 (N_2331,In_733,In_1216);
nand U2332 (N_2332,In_1486,In_1901);
and U2333 (N_2333,In_900,In_1661);
or U2334 (N_2334,In_279,In_1694);
or U2335 (N_2335,In_1768,In_1601);
nand U2336 (N_2336,In_1381,In_359);
nor U2337 (N_2337,In_491,In_504);
and U2338 (N_2338,In_1251,In_1126);
xor U2339 (N_2339,In_1735,In_938);
nor U2340 (N_2340,In_1424,In_800);
nor U2341 (N_2341,In_1430,In_1100);
or U2342 (N_2342,In_410,In_57);
and U2343 (N_2343,In_1050,In_848);
xnor U2344 (N_2344,In_1683,In_881);
or U2345 (N_2345,In_385,In_1616);
nand U2346 (N_2346,In_1294,In_850);
nand U2347 (N_2347,In_1252,In_1932);
or U2348 (N_2348,In_938,In_1996);
or U2349 (N_2349,In_1564,In_634);
nor U2350 (N_2350,In_1411,In_1120);
and U2351 (N_2351,In_1186,In_876);
and U2352 (N_2352,In_1227,In_793);
or U2353 (N_2353,In_1197,In_853);
nand U2354 (N_2354,In_1854,In_332);
and U2355 (N_2355,In_1208,In_1854);
and U2356 (N_2356,In_999,In_796);
or U2357 (N_2357,In_420,In_693);
xnor U2358 (N_2358,In_142,In_879);
nand U2359 (N_2359,In_1563,In_664);
or U2360 (N_2360,In_878,In_114);
nor U2361 (N_2361,In_1041,In_1487);
or U2362 (N_2362,In_207,In_1804);
nor U2363 (N_2363,In_398,In_95);
nor U2364 (N_2364,In_1791,In_1776);
nand U2365 (N_2365,In_416,In_1003);
and U2366 (N_2366,In_413,In_1211);
nor U2367 (N_2367,In_959,In_289);
and U2368 (N_2368,In_1217,In_744);
nor U2369 (N_2369,In_574,In_262);
nor U2370 (N_2370,In_1165,In_1778);
and U2371 (N_2371,In_1945,In_1118);
and U2372 (N_2372,In_321,In_13);
nand U2373 (N_2373,In_1695,In_539);
and U2374 (N_2374,In_1227,In_432);
and U2375 (N_2375,In_1370,In_1156);
nor U2376 (N_2376,In_1530,In_1793);
nand U2377 (N_2377,In_1116,In_1562);
or U2378 (N_2378,In_828,In_283);
or U2379 (N_2379,In_930,In_1046);
and U2380 (N_2380,In_825,In_671);
nor U2381 (N_2381,In_1767,In_1985);
nand U2382 (N_2382,In_1113,In_1608);
or U2383 (N_2383,In_1304,In_231);
or U2384 (N_2384,In_179,In_1168);
or U2385 (N_2385,In_647,In_1320);
or U2386 (N_2386,In_1659,In_1187);
or U2387 (N_2387,In_1798,In_1536);
nand U2388 (N_2388,In_1593,In_1440);
or U2389 (N_2389,In_1466,In_1627);
nand U2390 (N_2390,In_139,In_1561);
nor U2391 (N_2391,In_1634,In_150);
nand U2392 (N_2392,In_1508,In_1837);
nor U2393 (N_2393,In_1739,In_1564);
or U2394 (N_2394,In_1566,In_985);
nand U2395 (N_2395,In_1105,In_17);
nand U2396 (N_2396,In_1906,In_542);
and U2397 (N_2397,In_1290,In_944);
and U2398 (N_2398,In_502,In_1704);
xor U2399 (N_2399,In_381,In_1021);
or U2400 (N_2400,In_1935,In_725);
and U2401 (N_2401,In_1526,In_591);
nand U2402 (N_2402,In_1841,In_632);
or U2403 (N_2403,In_545,In_928);
and U2404 (N_2404,In_1017,In_1860);
and U2405 (N_2405,In_1014,In_884);
nor U2406 (N_2406,In_1133,In_648);
or U2407 (N_2407,In_185,In_676);
or U2408 (N_2408,In_1402,In_1817);
or U2409 (N_2409,In_1099,In_1491);
nor U2410 (N_2410,In_1760,In_523);
nand U2411 (N_2411,In_912,In_1208);
or U2412 (N_2412,In_1694,In_1968);
and U2413 (N_2413,In_885,In_1740);
or U2414 (N_2414,In_1432,In_574);
nor U2415 (N_2415,In_1940,In_870);
or U2416 (N_2416,In_838,In_1832);
or U2417 (N_2417,In_558,In_1289);
nor U2418 (N_2418,In_510,In_822);
nor U2419 (N_2419,In_1004,In_1794);
nand U2420 (N_2420,In_1163,In_151);
and U2421 (N_2421,In_784,In_225);
xor U2422 (N_2422,In_160,In_1912);
nand U2423 (N_2423,In_100,In_464);
and U2424 (N_2424,In_706,In_297);
or U2425 (N_2425,In_1826,In_270);
nand U2426 (N_2426,In_356,In_1090);
nor U2427 (N_2427,In_512,In_1234);
nor U2428 (N_2428,In_90,In_1205);
and U2429 (N_2429,In_404,In_867);
nor U2430 (N_2430,In_1463,In_999);
and U2431 (N_2431,In_1480,In_438);
nand U2432 (N_2432,In_76,In_292);
nand U2433 (N_2433,In_1555,In_588);
and U2434 (N_2434,In_1110,In_1855);
nand U2435 (N_2435,In_129,In_1436);
nand U2436 (N_2436,In_138,In_106);
and U2437 (N_2437,In_132,In_1180);
nand U2438 (N_2438,In_336,In_1215);
or U2439 (N_2439,In_502,In_829);
nand U2440 (N_2440,In_1425,In_921);
and U2441 (N_2441,In_437,In_345);
xor U2442 (N_2442,In_1294,In_1432);
and U2443 (N_2443,In_1142,In_1064);
and U2444 (N_2444,In_249,In_1897);
or U2445 (N_2445,In_1238,In_72);
nor U2446 (N_2446,In_21,In_587);
nand U2447 (N_2447,In_934,In_1200);
and U2448 (N_2448,In_495,In_1101);
and U2449 (N_2449,In_594,In_925);
or U2450 (N_2450,In_130,In_1771);
or U2451 (N_2451,In_582,In_1230);
nand U2452 (N_2452,In_675,In_1540);
nand U2453 (N_2453,In_128,In_775);
or U2454 (N_2454,In_873,In_1131);
and U2455 (N_2455,In_1702,In_1782);
and U2456 (N_2456,In_893,In_1002);
and U2457 (N_2457,In_1545,In_957);
or U2458 (N_2458,In_1116,In_333);
nand U2459 (N_2459,In_1613,In_1871);
nor U2460 (N_2460,In_1951,In_884);
nor U2461 (N_2461,In_296,In_1065);
and U2462 (N_2462,In_1362,In_799);
and U2463 (N_2463,In_416,In_1864);
or U2464 (N_2464,In_706,In_1312);
and U2465 (N_2465,In_1304,In_565);
or U2466 (N_2466,In_1334,In_544);
xnor U2467 (N_2467,In_1846,In_377);
nand U2468 (N_2468,In_164,In_1622);
nand U2469 (N_2469,In_320,In_31);
and U2470 (N_2470,In_537,In_1272);
xnor U2471 (N_2471,In_1947,In_327);
or U2472 (N_2472,In_1544,In_1117);
nand U2473 (N_2473,In_924,In_1091);
and U2474 (N_2474,In_1729,In_1062);
or U2475 (N_2475,In_715,In_47);
or U2476 (N_2476,In_1258,In_364);
and U2477 (N_2477,In_1975,In_10);
and U2478 (N_2478,In_1144,In_791);
or U2479 (N_2479,In_1438,In_1928);
nand U2480 (N_2480,In_880,In_1687);
nor U2481 (N_2481,In_1297,In_1283);
nor U2482 (N_2482,In_477,In_856);
nor U2483 (N_2483,In_269,In_1074);
or U2484 (N_2484,In_52,In_145);
nor U2485 (N_2485,In_82,In_69);
nand U2486 (N_2486,In_1105,In_1070);
or U2487 (N_2487,In_1642,In_304);
or U2488 (N_2488,In_496,In_1096);
nor U2489 (N_2489,In_982,In_513);
or U2490 (N_2490,In_294,In_26);
nand U2491 (N_2491,In_453,In_497);
nand U2492 (N_2492,In_1393,In_272);
and U2493 (N_2493,In_56,In_1007);
or U2494 (N_2494,In_224,In_1237);
and U2495 (N_2495,In_865,In_1441);
nand U2496 (N_2496,In_315,In_1491);
or U2497 (N_2497,In_592,In_1800);
and U2498 (N_2498,In_11,In_1870);
and U2499 (N_2499,In_1511,In_790);
nor U2500 (N_2500,In_1598,In_989);
nor U2501 (N_2501,In_1316,In_1745);
or U2502 (N_2502,In_109,In_585);
and U2503 (N_2503,In_1593,In_1083);
xor U2504 (N_2504,In_20,In_1790);
and U2505 (N_2505,In_110,In_1259);
and U2506 (N_2506,In_1558,In_1270);
nand U2507 (N_2507,In_1679,In_1065);
nand U2508 (N_2508,In_307,In_538);
xor U2509 (N_2509,In_1970,In_909);
nor U2510 (N_2510,In_127,In_1849);
and U2511 (N_2511,In_557,In_1226);
and U2512 (N_2512,In_192,In_392);
nand U2513 (N_2513,In_1301,In_1575);
and U2514 (N_2514,In_1957,In_1907);
nor U2515 (N_2515,In_1484,In_1834);
nand U2516 (N_2516,In_924,In_1690);
or U2517 (N_2517,In_253,In_612);
and U2518 (N_2518,In_1279,In_1453);
and U2519 (N_2519,In_517,In_1427);
or U2520 (N_2520,In_502,In_1164);
nor U2521 (N_2521,In_1622,In_754);
nor U2522 (N_2522,In_732,In_739);
or U2523 (N_2523,In_95,In_1144);
nor U2524 (N_2524,In_851,In_1031);
nor U2525 (N_2525,In_1224,In_1452);
or U2526 (N_2526,In_634,In_552);
xor U2527 (N_2527,In_921,In_1182);
nor U2528 (N_2528,In_1830,In_1719);
or U2529 (N_2529,In_35,In_1970);
or U2530 (N_2530,In_144,In_40);
nor U2531 (N_2531,In_1056,In_1148);
and U2532 (N_2532,In_1814,In_777);
nor U2533 (N_2533,In_1530,In_1540);
nand U2534 (N_2534,In_140,In_1281);
or U2535 (N_2535,In_367,In_415);
nand U2536 (N_2536,In_150,In_196);
nand U2537 (N_2537,In_1154,In_1974);
xnor U2538 (N_2538,In_80,In_1862);
nor U2539 (N_2539,In_1129,In_372);
and U2540 (N_2540,In_824,In_1661);
nor U2541 (N_2541,In_1461,In_375);
nor U2542 (N_2542,In_1321,In_1335);
and U2543 (N_2543,In_1198,In_1825);
or U2544 (N_2544,In_1862,In_1143);
nor U2545 (N_2545,In_1455,In_857);
nand U2546 (N_2546,In_781,In_913);
nor U2547 (N_2547,In_223,In_815);
or U2548 (N_2548,In_703,In_995);
nand U2549 (N_2549,In_775,In_998);
or U2550 (N_2550,In_202,In_237);
and U2551 (N_2551,In_178,In_361);
and U2552 (N_2552,In_1950,In_975);
nand U2553 (N_2553,In_1474,In_1450);
nand U2554 (N_2554,In_38,In_1700);
nand U2555 (N_2555,In_584,In_1773);
and U2556 (N_2556,In_433,In_491);
xnor U2557 (N_2557,In_1649,In_1835);
or U2558 (N_2558,In_163,In_199);
and U2559 (N_2559,In_1793,In_1392);
or U2560 (N_2560,In_857,In_637);
and U2561 (N_2561,In_1208,In_1971);
or U2562 (N_2562,In_1708,In_1860);
or U2563 (N_2563,In_687,In_271);
or U2564 (N_2564,In_146,In_294);
nor U2565 (N_2565,In_1869,In_62);
and U2566 (N_2566,In_167,In_1318);
nand U2567 (N_2567,In_1587,In_538);
nor U2568 (N_2568,In_1425,In_1004);
or U2569 (N_2569,In_567,In_41);
or U2570 (N_2570,In_1832,In_443);
xor U2571 (N_2571,In_1398,In_1255);
nand U2572 (N_2572,In_820,In_397);
nand U2573 (N_2573,In_475,In_1077);
nand U2574 (N_2574,In_598,In_1684);
or U2575 (N_2575,In_480,In_1711);
or U2576 (N_2576,In_1296,In_732);
or U2577 (N_2577,In_507,In_1201);
or U2578 (N_2578,In_1810,In_1019);
nor U2579 (N_2579,In_1030,In_788);
xnor U2580 (N_2580,In_1962,In_1773);
and U2581 (N_2581,In_1023,In_1725);
nor U2582 (N_2582,In_1168,In_1660);
and U2583 (N_2583,In_15,In_558);
nand U2584 (N_2584,In_594,In_746);
nor U2585 (N_2585,In_722,In_1684);
and U2586 (N_2586,In_427,In_1946);
and U2587 (N_2587,In_1314,In_1489);
or U2588 (N_2588,In_337,In_303);
or U2589 (N_2589,In_618,In_463);
xnor U2590 (N_2590,In_265,In_1853);
or U2591 (N_2591,In_1975,In_1910);
or U2592 (N_2592,In_838,In_1249);
or U2593 (N_2593,In_1394,In_1124);
nor U2594 (N_2594,In_1955,In_1100);
nand U2595 (N_2595,In_57,In_67);
and U2596 (N_2596,In_457,In_556);
and U2597 (N_2597,In_973,In_1608);
nor U2598 (N_2598,In_1253,In_1876);
and U2599 (N_2599,In_114,In_1117);
nand U2600 (N_2600,In_349,In_1675);
nor U2601 (N_2601,In_137,In_458);
and U2602 (N_2602,In_56,In_1336);
nand U2603 (N_2603,In_1063,In_517);
and U2604 (N_2604,In_1020,In_784);
xor U2605 (N_2605,In_1077,In_1648);
nor U2606 (N_2606,In_125,In_987);
nor U2607 (N_2607,In_1622,In_510);
nor U2608 (N_2608,In_370,In_1952);
nor U2609 (N_2609,In_1082,In_1459);
or U2610 (N_2610,In_1610,In_1050);
and U2611 (N_2611,In_1725,In_1331);
nor U2612 (N_2612,In_985,In_850);
nor U2613 (N_2613,In_398,In_1578);
nand U2614 (N_2614,In_1044,In_284);
nand U2615 (N_2615,In_230,In_1849);
nand U2616 (N_2616,In_1238,In_1881);
nor U2617 (N_2617,In_287,In_1033);
nor U2618 (N_2618,In_512,In_428);
nor U2619 (N_2619,In_1063,In_1942);
and U2620 (N_2620,In_580,In_789);
or U2621 (N_2621,In_1359,In_1139);
nand U2622 (N_2622,In_963,In_1055);
and U2623 (N_2623,In_1986,In_1716);
or U2624 (N_2624,In_1749,In_896);
or U2625 (N_2625,In_1582,In_1194);
xor U2626 (N_2626,In_337,In_1580);
and U2627 (N_2627,In_1435,In_1133);
nor U2628 (N_2628,In_1103,In_1890);
nand U2629 (N_2629,In_1310,In_1661);
nand U2630 (N_2630,In_1434,In_1230);
or U2631 (N_2631,In_1990,In_1146);
nand U2632 (N_2632,In_22,In_791);
or U2633 (N_2633,In_1613,In_37);
or U2634 (N_2634,In_1402,In_1539);
nor U2635 (N_2635,In_539,In_1478);
nand U2636 (N_2636,In_1385,In_98);
or U2637 (N_2637,In_1429,In_1233);
or U2638 (N_2638,In_593,In_1254);
and U2639 (N_2639,In_572,In_246);
or U2640 (N_2640,In_776,In_1184);
nand U2641 (N_2641,In_83,In_1754);
or U2642 (N_2642,In_559,In_1314);
or U2643 (N_2643,In_335,In_1476);
and U2644 (N_2644,In_1039,In_642);
and U2645 (N_2645,In_1119,In_1939);
or U2646 (N_2646,In_654,In_395);
and U2647 (N_2647,In_337,In_557);
or U2648 (N_2648,In_691,In_429);
or U2649 (N_2649,In_1572,In_981);
nand U2650 (N_2650,In_806,In_1920);
and U2651 (N_2651,In_911,In_1447);
or U2652 (N_2652,In_26,In_517);
nand U2653 (N_2653,In_736,In_796);
nand U2654 (N_2654,In_1663,In_826);
nand U2655 (N_2655,In_1792,In_506);
nand U2656 (N_2656,In_1359,In_1560);
xnor U2657 (N_2657,In_1173,In_535);
and U2658 (N_2658,In_1174,In_715);
or U2659 (N_2659,In_641,In_900);
nand U2660 (N_2660,In_1359,In_389);
nor U2661 (N_2661,In_124,In_1241);
or U2662 (N_2662,In_1341,In_50);
and U2663 (N_2663,In_1712,In_103);
or U2664 (N_2664,In_1309,In_1612);
nand U2665 (N_2665,In_183,In_344);
nand U2666 (N_2666,In_1434,In_1125);
nor U2667 (N_2667,In_1731,In_1104);
nand U2668 (N_2668,In_377,In_1134);
nor U2669 (N_2669,In_312,In_64);
xnor U2670 (N_2670,In_1223,In_606);
or U2671 (N_2671,In_698,In_1366);
and U2672 (N_2672,In_1116,In_846);
or U2673 (N_2673,In_295,In_1263);
and U2674 (N_2674,In_127,In_301);
and U2675 (N_2675,In_753,In_183);
and U2676 (N_2676,In_792,In_134);
or U2677 (N_2677,In_534,In_643);
and U2678 (N_2678,In_517,In_936);
or U2679 (N_2679,In_281,In_646);
nor U2680 (N_2680,In_1109,In_798);
or U2681 (N_2681,In_1803,In_1246);
xor U2682 (N_2682,In_1791,In_1990);
and U2683 (N_2683,In_198,In_1692);
and U2684 (N_2684,In_1754,In_698);
nor U2685 (N_2685,In_108,In_1069);
nand U2686 (N_2686,In_670,In_1739);
and U2687 (N_2687,In_1523,In_533);
and U2688 (N_2688,In_1844,In_1690);
nor U2689 (N_2689,In_417,In_431);
xnor U2690 (N_2690,In_120,In_1174);
xor U2691 (N_2691,In_898,In_1915);
nor U2692 (N_2692,In_1263,In_1348);
and U2693 (N_2693,In_1931,In_320);
nand U2694 (N_2694,In_132,In_1845);
xor U2695 (N_2695,In_1977,In_1635);
or U2696 (N_2696,In_63,In_1575);
or U2697 (N_2697,In_1727,In_1900);
and U2698 (N_2698,In_834,In_701);
and U2699 (N_2699,In_776,In_1108);
and U2700 (N_2700,In_539,In_554);
and U2701 (N_2701,In_1233,In_1350);
nand U2702 (N_2702,In_1490,In_1926);
or U2703 (N_2703,In_33,In_1490);
or U2704 (N_2704,In_1798,In_882);
or U2705 (N_2705,In_111,In_147);
nand U2706 (N_2706,In_410,In_485);
or U2707 (N_2707,In_1197,In_906);
or U2708 (N_2708,In_59,In_1223);
or U2709 (N_2709,In_221,In_452);
nand U2710 (N_2710,In_960,In_1453);
and U2711 (N_2711,In_1012,In_1407);
or U2712 (N_2712,In_1398,In_331);
nor U2713 (N_2713,In_1458,In_128);
nor U2714 (N_2714,In_284,In_337);
nor U2715 (N_2715,In_1068,In_844);
and U2716 (N_2716,In_1250,In_769);
and U2717 (N_2717,In_1002,In_1387);
nand U2718 (N_2718,In_703,In_712);
nor U2719 (N_2719,In_1446,In_1715);
and U2720 (N_2720,In_925,In_1244);
nor U2721 (N_2721,In_684,In_118);
nand U2722 (N_2722,In_1787,In_1536);
or U2723 (N_2723,In_913,In_1231);
and U2724 (N_2724,In_1883,In_1655);
or U2725 (N_2725,In_1602,In_383);
or U2726 (N_2726,In_1702,In_1916);
nand U2727 (N_2727,In_702,In_160);
or U2728 (N_2728,In_654,In_849);
or U2729 (N_2729,In_1378,In_1798);
and U2730 (N_2730,In_732,In_568);
or U2731 (N_2731,In_1986,In_167);
nor U2732 (N_2732,In_1502,In_1390);
nor U2733 (N_2733,In_1309,In_1730);
nor U2734 (N_2734,In_1647,In_524);
or U2735 (N_2735,In_673,In_283);
or U2736 (N_2736,In_1367,In_487);
and U2737 (N_2737,In_1500,In_1461);
and U2738 (N_2738,In_1453,In_79);
nor U2739 (N_2739,In_1942,In_904);
or U2740 (N_2740,In_916,In_8);
or U2741 (N_2741,In_659,In_354);
nor U2742 (N_2742,In_299,In_1779);
nand U2743 (N_2743,In_1990,In_1821);
and U2744 (N_2744,In_1914,In_445);
or U2745 (N_2745,In_829,In_190);
nor U2746 (N_2746,In_1935,In_1967);
nand U2747 (N_2747,In_567,In_232);
nor U2748 (N_2748,In_338,In_1230);
and U2749 (N_2749,In_1862,In_562);
and U2750 (N_2750,In_1255,In_831);
or U2751 (N_2751,In_68,In_1622);
nor U2752 (N_2752,In_1752,In_1881);
nand U2753 (N_2753,In_1159,In_1683);
nand U2754 (N_2754,In_549,In_604);
nand U2755 (N_2755,In_537,In_1495);
and U2756 (N_2756,In_1497,In_1289);
nor U2757 (N_2757,In_917,In_1943);
and U2758 (N_2758,In_307,In_1279);
and U2759 (N_2759,In_474,In_1340);
and U2760 (N_2760,In_327,In_51);
nor U2761 (N_2761,In_1444,In_287);
and U2762 (N_2762,In_1712,In_733);
nor U2763 (N_2763,In_142,In_538);
or U2764 (N_2764,In_1674,In_569);
nor U2765 (N_2765,In_506,In_323);
xor U2766 (N_2766,In_455,In_1477);
or U2767 (N_2767,In_1432,In_143);
xnor U2768 (N_2768,In_368,In_1215);
nor U2769 (N_2769,In_1831,In_1371);
nand U2770 (N_2770,In_1989,In_1969);
and U2771 (N_2771,In_341,In_892);
nor U2772 (N_2772,In_218,In_1489);
nor U2773 (N_2773,In_342,In_684);
nand U2774 (N_2774,In_1529,In_968);
nand U2775 (N_2775,In_16,In_757);
nor U2776 (N_2776,In_1072,In_842);
nor U2777 (N_2777,In_1136,In_369);
and U2778 (N_2778,In_1386,In_1000);
and U2779 (N_2779,In_855,In_1614);
and U2780 (N_2780,In_930,In_559);
nand U2781 (N_2781,In_584,In_896);
or U2782 (N_2782,In_820,In_1771);
or U2783 (N_2783,In_709,In_971);
and U2784 (N_2784,In_1630,In_106);
or U2785 (N_2785,In_1503,In_3);
nor U2786 (N_2786,In_1282,In_1849);
and U2787 (N_2787,In_495,In_1301);
nand U2788 (N_2788,In_1047,In_283);
nand U2789 (N_2789,In_1272,In_1913);
or U2790 (N_2790,In_610,In_463);
nor U2791 (N_2791,In_1106,In_239);
nor U2792 (N_2792,In_1820,In_1302);
nor U2793 (N_2793,In_792,In_349);
or U2794 (N_2794,In_1564,In_1743);
nor U2795 (N_2795,In_1328,In_530);
nor U2796 (N_2796,In_577,In_1246);
nor U2797 (N_2797,In_580,In_929);
or U2798 (N_2798,In_1399,In_418);
nand U2799 (N_2799,In_35,In_1848);
nand U2800 (N_2800,In_416,In_1358);
and U2801 (N_2801,In_307,In_1909);
or U2802 (N_2802,In_1942,In_258);
nor U2803 (N_2803,In_1102,In_1013);
nand U2804 (N_2804,In_1288,In_1024);
or U2805 (N_2805,In_296,In_1778);
nand U2806 (N_2806,In_1843,In_145);
xnor U2807 (N_2807,In_1641,In_1073);
or U2808 (N_2808,In_1524,In_713);
and U2809 (N_2809,In_995,In_1828);
nor U2810 (N_2810,In_527,In_1810);
or U2811 (N_2811,In_503,In_1103);
or U2812 (N_2812,In_1431,In_1148);
or U2813 (N_2813,In_972,In_1284);
nor U2814 (N_2814,In_1863,In_1743);
or U2815 (N_2815,In_481,In_236);
or U2816 (N_2816,In_884,In_624);
and U2817 (N_2817,In_1046,In_1652);
or U2818 (N_2818,In_1589,In_1003);
or U2819 (N_2819,In_1037,In_804);
nand U2820 (N_2820,In_1379,In_1806);
nand U2821 (N_2821,In_865,In_363);
nor U2822 (N_2822,In_1470,In_1579);
nor U2823 (N_2823,In_1045,In_1133);
nand U2824 (N_2824,In_1694,In_1686);
nand U2825 (N_2825,In_128,In_1009);
and U2826 (N_2826,In_1530,In_1861);
nor U2827 (N_2827,In_630,In_1717);
or U2828 (N_2828,In_1558,In_967);
nand U2829 (N_2829,In_1637,In_1577);
and U2830 (N_2830,In_737,In_1435);
and U2831 (N_2831,In_1557,In_1482);
nand U2832 (N_2832,In_547,In_1107);
and U2833 (N_2833,In_1958,In_685);
nand U2834 (N_2834,In_500,In_1264);
nand U2835 (N_2835,In_947,In_1290);
nand U2836 (N_2836,In_913,In_1069);
nor U2837 (N_2837,In_1299,In_1972);
nor U2838 (N_2838,In_617,In_1510);
nor U2839 (N_2839,In_1938,In_736);
or U2840 (N_2840,In_1485,In_1169);
nand U2841 (N_2841,In_211,In_167);
xnor U2842 (N_2842,In_1694,In_1705);
or U2843 (N_2843,In_120,In_585);
or U2844 (N_2844,In_271,In_387);
nand U2845 (N_2845,In_735,In_1718);
or U2846 (N_2846,In_137,In_435);
nand U2847 (N_2847,In_1978,In_1929);
xnor U2848 (N_2848,In_727,In_1899);
nor U2849 (N_2849,In_847,In_744);
nand U2850 (N_2850,In_226,In_430);
nor U2851 (N_2851,In_362,In_1272);
nand U2852 (N_2852,In_834,In_217);
xor U2853 (N_2853,In_248,In_1335);
nand U2854 (N_2854,In_524,In_1433);
nor U2855 (N_2855,In_574,In_1622);
or U2856 (N_2856,In_699,In_47);
or U2857 (N_2857,In_1782,In_484);
or U2858 (N_2858,In_270,In_118);
and U2859 (N_2859,In_659,In_92);
nor U2860 (N_2860,In_34,In_1068);
and U2861 (N_2861,In_362,In_328);
and U2862 (N_2862,In_781,In_1802);
nand U2863 (N_2863,In_1138,In_926);
nor U2864 (N_2864,In_370,In_329);
and U2865 (N_2865,In_250,In_937);
or U2866 (N_2866,In_1824,In_1507);
nor U2867 (N_2867,In_108,In_1649);
nand U2868 (N_2868,In_96,In_1379);
nand U2869 (N_2869,In_895,In_999);
nand U2870 (N_2870,In_1914,In_1900);
or U2871 (N_2871,In_565,In_1298);
or U2872 (N_2872,In_1497,In_146);
nor U2873 (N_2873,In_332,In_1580);
nand U2874 (N_2874,In_1655,In_445);
nand U2875 (N_2875,In_1431,In_168);
and U2876 (N_2876,In_82,In_1047);
nor U2877 (N_2877,In_1430,In_1640);
or U2878 (N_2878,In_1106,In_1462);
or U2879 (N_2879,In_1737,In_1144);
nand U2880 (N_2880,In_1239,In_1264);
or U2881 (N_2881,In_1881,In_248);
and U2882 (N_2882,In_253,In_133);
nand U2883 (N_2883,In_1942,In_1855);
or U2884 (N_2884,In_536,In_507);
or U2885 (N_2885,In_404,In_86);
nand U2886 (N_2886,In_675,In_1258);
and U2887 (N_2887,In_1598,In_1522);
nor U2888 (N_2888,In_1287,In_961);
nand U2889 (N_2889,In_1674,In_225);
and U2890 (N_2890,In_1862,In_1434);
and U2891 (N_2891,In_1030,In_805);
or U2892 (N_2892,In_369,In_1137);
or U2893 (N_2893,In_368,In_1251);
or U2894 (N_2894,In_1054,In_171);
or U2895 (N_2895,In_1320,In_542);
or U2896 (N_2896,In_324,In_106);
and U2897 (N_2897,In_1596,In_1064);
and U2898 (N_2898,In_788,In_379);
nor U2899 (N_2899,In_1551,In_1441);
and U2900 (N_2900,In_458,In_221);
and U2901 (N_2901,In_835,In_1427);
or U2902 (N_2902,In_1548,In_647);
or U2903 (N_2903,In_1672,In_739);
nand U2904 (N_2904,In_528,In_1295);
nor U2905 (N_2905,In_1160,In_1946);
nor U2906 (N_2906,In_1263,In_999);
and U2907 (N_2907,In_984,In_340);
nor U2908 (N_2908,In_1439,In_542);
or U2909 (N_2909,In_1152,In_1605);
and U2910 (N_2910,In_1213,In_1233);
nand U2911 (N_2911,In_222,In_1872);
xor U2912 (N_2912,In_1002,In_710);
nor U2913 (N_2913,In_1461,In_980);
and U2914 (N_2914,In_695,In_1149);
or U2915 (N_2915,In_1111,In_25);
and U2916 (N_2916,In_712,In_737);
nand U2917 (N_2917,In_1999,In_1411);
nor U2918 (N_2918,In_296,In_828);
or U2919 (N_2919,In_1183,In_449);
nand U2920 (N_2920,In_768,In_1904);
nand U2921 (N_2921,In_1638,In_1311);
or U2922 (N_2922,In_1291,In_826);
or U2923 (N_2923,In_1359,In_1671);
or U2924 (N_2924,In_2,In_1309);
and U2925 (N_2925,In_788,In_147);
nand U2926 (N_2926,In_1932,In_1578);
or U2927 (N_2927,In_1444,In_28);
and U2928 (N_2928,In_502,In_1966);
and U2929 (N_2929,In_677,In_136);
nand U2930 (N_2930,In_1947,In_756);
and U2931 (N_2931,In_1772,In_937);
nor U2932 (N_2932,In_98,In_1796);
or U2933 (N_2933,In_633,In_1639);
nor U2934 (N_2934,In_175,In_293);
nor U2935 (N_2935,In_1826,In_1832);
and U2936 (N_2936,In_699,In_859);
nand U2937 (N_2937,In_345,In_1507);
nor U2938 (N_2938,In_294,In_526);
nand U2939 (N_2939,In_436,In_630);
nor U2940 (N_2940,In_414,In_961);
or U2941 (N_2941,In_1486,In_629);
and U2942 (N_2942,In_694,In_1200);
nor U2943 (N_2943,In_1022,In_546);
and U2944 (N_2944,In_814,In_950);
nor U2945 (N_2945,In_1915,In_1707);
nor U2946 (N_2946,In_1551,In_1151);
nor U2947 (N_2947,In_1589,In_1793);
and U2948 (N_2948,In_1158,In_1501);
or U2949 (N_2949,In_1610,In_1077);
nor U2950 (N_2950,In_21,In_1513);
and U2951 (N_2951,In_862,In_1053);
xor U2952 (N_2952,In_1178,In_482);
nand U2953 (N_2953,In_271,In_1027);
nand U2954 (N_2954,In_441,In_824);
nor U2955 (N_2955,In_1917,In_1664);
nor U2956 (N_2956,In_389,In_1956);
or U2957 (N_2957,In_1831,In_1458);
nand U2958 (N_2958,In_1466,In_533);
nand U2959 (N_2959,In_507,In_256);
and U2960 (N_2960,In_1900,In_499);
or U2961 (N_2961,In_1612,In_1506);
and U2962 (N_2962,In_1059,In_1995);
nor U2963 (N_2963,In_1931,In_1498);
nor U2964 (N_2964,In_1672,In_1986);
and U2965 (N_2965,In_963,In_1682);
nand U2966 (N_2966,In_1123,In_914);
or U2967 (N_2967,In_1341,In_1653);
nor U2968 (N_2968,In_6,In_1919);
nand U2969 (N_2969,In_1457,In_766);
or U2970 (N_2970,In_981,In_1184);
nor U2971 (N_2971,In_1663,In_1394);
or U2972 (N_2972,In_1204,In_1652);
nand U2973 (N_2973,In_700,In_1409);
and U2974 (N_2974,In_734,In_1848);
nand U2975 (N_2975,In_846,In_600);
nand U2976 (N_2976,In_494,In_841);
or U2977 (N_2977,In_1850,In_1181);
or U2978 (N_2978,In_842,In_155);
and U2979 (N_2979,In_1386,In_155);
and U2980 (N_2980,In_317,In_678);
nand U2981 (N_2981,In_1923,In_1647);
and U2982 (N_2982,In_280,In_828);
and U2983 (N_2983,In_1365,In_1245);
or U2984 (N_2984,In_1499,In_1880);
or U2985 (N_2985,In_416,In_1631);
or U2986 (N_2986,In_1650,In_1195);
nand U2987 (N_2987,In_1827,In_1551);
and U2988 (N_2988,In_467,In_1855);
or U2989 (N_2989,In_188,In_366);
nand U2990 (N_2990,In_1413,In_1009);
and U2991 (N_2991,In_1320,In_359);
or U2992 (N_2992,In_588,In_815);
nor U2993 (N_2993,In_796,In_576);
or U2994 (N_2994,In_1465,In_107);
nand U2995 (N_2995,In_688,In_1881);
and U2996 (N_2996,In_746,In_453);
nand U2997 (N_2997,In_235,In_1779);
or U2998 (N_2998,In_1375,In_902);
nor U2999 (N_2999,In_1175,In_167);
nand U3000 (N_3000,In_827,In_1862);
nand U3001 (N_3001,In_843,In_161);
nor U3002 (N_3002,In_732,In_381);
nor U3003 (N_3003,In_1718,In_396);
and U3004 (N_3004,In_1686,In_1571);
nor U3005 (N_3005,In_275,In_1876);
nor U3006 (N_3006,In_887,In_564);
nand U3007 (N_3007,In_321,In_754);
or U3008 (N_3008,In_1913,In_501);
and U3009 (N_3009,In_1224,In_476);
nand U3010 (N_3010,In_1465,In_495);
or U3011 (N_3011,In_630,In_995);
or U3012 (N_3012,In_1879,In_250);
and U3013 (N_3013,In_992,In_640);
nor U3014 (N_3014,In_711,In_1561);
or U3015 (N_3015,In_1287,In_411);
nand U3016 (N_3016,In_785,In_97);
nand U3017 (N_3017,In_492,In_666);
and U3018 (N_3018,In_1848,In_856);
and U3019 (N_3019,In_1497,In_1900);
and U3020 (N_3020,In_479,In_1554);
xor U3021 (N_3021,In_1061,In_1026);
nand U3022 (N_3022,In_754,In_433);
nor U3023 (N_3023,In_1101,In_375);
nor U3024 (N_3024,In_1105,In_13);
nand U3025 (N_3025,In_299,In_666);
or U3026 (N_3026,In_826,In_1579);
nand U3027 (N_3027,In_1629,In_1403);
xnor U3028 (N_3028,In_1112,In_4);
nor U3029 (N_3029,In_1992,In_1487);
and U3030 (N_3030,In_957,In_677);
nand U3031 (N_3031,In_1124,In_447);
or U3032 (N_3032,In_1051,In_561);
and U3033 (N_3033,In_495,In_1499);
and U3034 (N_3034,In_697,In_1565);
and U3035 (N_3035,In_221,In_1821);
nand U3036 (N_3036,In_164,In_1241);
and U3037 (N_3037,In_1033,In_1915);
nor U3038 (N_3038,In_1437,In_1048);
nand U3039 (N_3039,In_258,In_1374);
and U3040 (N_3040,In_96,In_1358);
nand U3041 (N_3041,In_899,In_846);
nor U3042 (N_3042,In_11,In_199);
nor U3043 (N_3043,In_552,In_1194);
and U3044 (N_3044,In_1840,In_1392);
nand U3045 (N_3045,In_5,In_1784);
nor U3046 (N_3046,In_1875,In_838);
nand U3047 (N_3047,In_375,In_1632);
or U3048 (N_3048,In_358,In_535);
nor U3049 (N_3049,In_235,In_1884);
nand U3050 (N_3050,In_1331,In_1573);
nand U3051 (N_3051,In_373,In_486);
nand U3052 (N_3052,In_951,In_260);
and U3053 (N_3053,In_1704,In_1507);
nor U3054 (N_3054,In_421,In_23);
and U3055 (N_3055,In_860,In_1305);
nor U3056 (N_3056,In_1961,In_1527);
and U3057 (N_3057,In_1802,In_430);
or U3058 (N_3058,In_116,In_1368);
nand U3059 (N_3059,In_875,In_1058);
nand U3060 (N_3060,In_949,In_1591);
xnor U3061 (N_3061,In_761,In_597);
or U3062 (N_3062,In_609,In_708);
nand U3063 (N_3063,In_1903,In_26);
and U3064 (N_3064,In_1968,In_164);
or U3065 (N_3065,In_1797,In_513);
and U3066 (N_3066,In_708,In_193);
or U3067 (N_3067,In_284,In_512);
or U3068 (N_3068,In_765,In_1106);
nor U3069 (N_3069,In_297,In_149);
nand U3070 (N_3070,In_266,In_296);
and U3071 (N_3071,In_61,In_100);
xnor U3072 (N_3072,In_1409,In_1197);
and U3073 (N_3073,In_1781,In_555);
nor U3074 (N_3074,In_1586,In_125);
and U3075 (N_3075,In_371,In_511);
or U3076 (N_3076,In_1284,In_731);
or U3077 (N_3077,In_1887,In_1697);
nand U3078 (N_3078,In_250,In_1319);
or U3079 (N_3079,In_493,In_1826);
and U3080 (N_3080,In_1588,In_1040);
nor U3081 (N_3081,In_170,In_567);
or U3082 (N_3082,In_463,In_1673);
or U3083 (N_3083,In_542,In_853);
or U3084 (N_3084,In_37,In_1019);
and U3085 (N_3085,In_38,In_920);
nor U3086 (N_3086,In_206,In_1686);
or U3087 (N_3087,In_1217,In_1152);
nor U3088 (N_3088,In_147,In_520);
nand U3089 (N_3089,In_1440,In_1876);
nand U3090 (N_3090,In_314,In_272);
nor U3091 (N_3091,In_76,In_679);
or U3092 (N_3092,In_1393,In_513);
nor U3093 (N_3093,In_1758,In_845);
nand U3094 (N_3094,In_1568,In_1144);
and U3095 (N_3095,In_386,In_1012);
xor U3096 (N_3096,In_1997,In_568);
and U3097 (N_3097,In_1710,In_465);
and U3098 (N_3098,In_619,In_127);
or U3099 (N_3099,In_1427,In_92);
and U3100 (N_3100,In_155,In_1750);
xnor U3101 (N_3101,In_1710,In_1350);
nor U3102 (N_3102,In_873,In_987);
or U3103 (N_3103,In_1719,In_134);
or U3104 (N_3104,In_716,In_1963);
nor U3105 (N_3105,In_1188,In_149);
or U3106 (N_3106,In_566,In_458);
or U3107 (N_3107,In_1883,In_1310);
nand U3108 (N_3108,In_1747,In_177);
nand U3109 (N_3109,In_1999,In_1014);
nand U3110 (N_3110,In_1751,In_1407);
xnor U3111 (N_3111,In_1659,In_1322);
nand U3112 (N_3112,In_468,In_1643);
and U3113 (N_3113,In_1766,In_1600);
or U3114 (N_3114,In_390,In_1724);
or U3115 (N_3115,In_10,In_29);
or U3116 (N_3116,In_1367,In_1380);
nand U3117 (N_3117,In_885,In_1412);
nor U3118 (N_3118,In_518,In_1160);
nand U3119 (N_3119,In_1293,In_573);
nor U3120 (N_3120,In_124,In_1986);
nor U3121 (N_3121,In_4,In_1339);
or U3122 (N_3122,In_541,In_823);
nand U3123 (N_3123,In_441,In_1621);
or U3124 (N_3124,In_21,In_1835);
or U3125 (N_3125,In_1751,In_678);
xor U3126 (N_3126,In_400,In_1221);
or U3127 (N_3127,In_874,In_1876);
nor U3128 (N_3128,In_322,In_1807);
and U3129 (N_3129,In_1229,In_1258);
nor U3130 (N_3130,In_569,In_927);
and U3131 (N_3131,In_1754,In_1448);
nand U3132 (N_3132,In_1877,In_1768);
and U3133 (N_3133,In_1796,In_508);
nor U3134 (N_3134,In_1999,In_572);
nand U3135 (N_3135,In_960,In_1648);
or U3136 (N_3136,In_1148,In_1514);
or U3137 (N_3137,In_476,In_1110);
or U3138 (N_3138,In_270,In_1850);
or U3139 (N_3139,In_87,In_891);
or U3140 (N_3140,In_730,In_1312);
and U3141 (N_3141,In_373,In_445);
xor U3142 (N_3142,In_103,In_248);
nor U3143 (N_3143,In_1616,In_1082);
nand U3144 (N_3144,In_1372,In_423);
nand U3145 (N_3145,In_1116,In_1760);
nor U3146 (N_3146,In_1840,In_1490);
or U3147 (N_3147,In_796,In_1707);
and U3148 (N_3148,In_1897,In_418);
nand U3149 (N_3149,In_1251,In_1735);
or U3150 (N_3150,In_1347,In_1950);
nor U3151 (N_3151,In_967,In_387);
and U3152 (N_3152,In_224,In_1513);
or U3153 (N_3153,In_1984,In_1447);
or U3154 (N_3154,In_743,In_1441);
nor U3155 (N_3155,In_140,In_949);
nor U3156 (N_3156,In_1390,In_1379);
and U3157 (N_3157,In_128,In_1489);
nand U3158 (N_3158,In_150,In_749);
or U3159 (N_3159,In_346,In_42);
nor U3160 (N_3160,In_1713,In_1695);
or U3161 (N_3161,In_234,In_1474);
nor U3162 (N_3162,In_716,In_127);
and U3163 (N_3163,In_1895,In_1872);
and U3164 (N_3164,In_640,In_1858);
nor U3165 (N_3165,In_281,In_914);
and U3166 (N_3166,In_1764,In_1899);
or U3167 (N_3167,In_1871,In_720);
nor U3168 (N_3168,In_1434,In_1082);
nor U3169 (N_3169,In_1459,In_441);
nand U3170 (N_3170,In_1137,In_1877);
or U3171 (N_3171,In_996,In_425);
or U3172 (N_3172,In_758,In_940);
and U3173 (N_3173,In_391,In_797);
nor U3174 (N_3174,In_15,In_484);
and U3175 (N_3175,In_391,In_124);
nor U3176 (N_3176,In_1780,In_1117);
and U3177 (N_3177,In_1559,In_845);
nand U3178 (N_3178,In_585,In_311);
or U3179 (N_3179,In_340,In_755);
nand U3180 (N_3180,In_1781,In_1773);
nand U3181 (N_3181,In_284,In_299);
or U3182 (N_3182,In_1924,In_185);
and U3183 (N_3183,In_1898,In_1097);
nand U3184 (N_3184,In_909,In_1117);
or U3185 (N_3185,In_1489,In_1416);
or U3186 (N_3186,In_849,In_157);
nor U3187 (N_3187,In_953,In_1451);
nand U3188 (N_3188,In_1656,In_1837);
nand U3189 (N_3189,In_792,In_1597);
nor U3190 (N_3190,In_1604,In_801);
or U3191 (N_3191,In_351,In_1388);
nand U3192 (N_3192,In_1264,In_1899);
nand U3193 (N_3193,In_99,In_1791);
nor U3194 (N_3194,In_1757,In_411);
and U3195 (N_3195,In_284,In_1925);
nor U3196 (N_3196,In_1103,In_129);
nor U3197 (N_3197,In_1428,In_1347);
and U3198 (N_3198,In_832,In_292);
and U3199 (N_3199,In_1177,In_1258);
nand U3200 (N_3200,In_814,In_120);
or U3201 (N_3201,In_1042,In_1312);
and U3202 (N_3202,In_1492,In_325);
and U3203 (N_3203,In_242,In_823);
or U3204 (N_3204,In_1838,In_1086);
and U3205 (N_3205,In_1332,In_1427);
and U3206 (N_3206,In_767,In_879);
nor U3207 (N_3207,In_1058,In_1988);
xor U3208 (N_3208,In_1707,In_535);
nand U3209 (N_3209,In_152,In_505);
nand U3210 (N_3210,In_103,In_742);
nor U3211 (N_3211,In_371,In_894);
and U3212 (N_3212,In_1877,In_620);
nor U3213 (N_3213,In_1620,In_1003);
and U3214 (N_3214,In_1006,In_1427);
and U3215 (N_3215,In_1037,In_438);
or U3216 (N_3216,In_1330,In_591);
nor U3217 (N_3217,In_1265,In_1082);
and U3218 (N_3218,In_1199,In_1633);
nand U3219 (N_3219,In_1803,In_1683);
nand U3220 (N_3220,In_1879,In_1821);
nor U3221 (N_3221,In_350,In_1890);
nor U3222 (N_3222,In_500,In_1286);
and U3223 (N_3223,In_215,In_272);
nor U3224 (N_3224,In_747,In_653);
xnor U3225 (N_3225,In_809,In_897);
or U3226 (N_3226,In_1889,In_511);
and U3227 (N_3227,In_1881,In_1845);
and U3228 (N_3228,In_213,In_707);
and U3229 (N_3229,In_1696,In_1819);
nand U3230 (N_3230,In_1496,In_1201);
or U3231 (N_3231,In_908,In_332);
or U3232 (N_3232,In_400,In_1862);
nand U3233 (N_3233,In_1961,In_1894);
and U3234 (N_3234,In_1629,In_1535);
or U3235 (N_3235,In_751,In_1546);
and U3236 (N_3236,In_100,In_1324);
or U3237 (N_3237,In_1194,In_83);
nand U3238 (N_3238,In_1497,In_744);
nor U3239 (N_3239,In_1000,In_637);
nand U3240 (N_3240,In_1747,In_794);
or U3241 (N_3241,In_855,In_185);
nand U3242 (N_3242,In_320,In_1921);
nand U3243 (N_3243,In_366,In_295);
nor U3244 (N_3244,In_852,In_1367);
nand U3245 (N_3245,In_1161,In_1936);
and U3246 (N_3246,In_1937,In_639);
nand U3247 (N_3247,In_1692,In_180);
or U3248 (N_3248,In_1029,In_1362);
nor U3249 (N_3249,In_1303,In_998);
and U3250 (N_3250,In_26,In_253);
or U3251 (N_3251,In_470,In_465);
or U3252 (N_3252,In_471,In_510);
nand U3253 (N_3253,In_428,In_1120);
nand U3254 (N_3254,In_1318,In_1142);
nand U3255 (N_3255,In_796,In_984);
nor U3256 (N_3256,In_1146,In_1963);
and U3257 (N_3257,In_746,In_737);
nand U3258 (N_3258,In_1721,In_1212);
nand U3259 (N_3259,In_97,In_983);
nor U3260 (N_3260,In_812,In_1552);
nor U3261 (N_3261,In_1497,In_1318);
and U3262 (N_3262,In_384,In_1089);
or U3263 (N_3263,In_265,In_1411);
and U3264 (N_3264,In_1884,In_565);
and U3265 (N_3265,In_536,In_600);
nand U3266 (N_3266,In_128,In_1614);
nor U3267 (N_3267,In_1789,In_1401);
nand U3268 (N_3268,In_823,In_1499);
nor U3269 (N_3269,In_1569,In_469);
nor U3270 (N_3270,In_1122,In_1434);
nand U3271 (N_3271,In_787,In_628);
and U3272 (N_3272,In_283,In_806);
and U3273 (N_3273,In_326,In_144);
and U3274 (N_3274,In_681,In_1284);
or U3275 (N_3275,In_774,In_106);
nand U3276 (N_3276,In_680,In_973);
or U3277 (N_3277,In_1882,In_477);
and U3278 (N_3278,In_189,In_1125);
or U3279 (N_3279,In_494,In_699);
and U3280 (N_3280,In_846,In_1429);
nor U3281 (N_3281,In_255,In_1680);
nand U3282 (N_3282,In_372,In_566);
or U3283 (N_3283,In_20,In_510);
and U3284 (N_3284,In_1104,In_1084);
nor U3285 (N_3285,In_249,In_272);
or U3286 (N_3286,In_85,In_117);
nor U3287 (N_3287,In_1740,In_868);
nand U3288 (N_3288,In_630,In_429);
or U3289 (N_3289,In_706,In_1042);
and U3290 (N_3290,In_964,In_1973);
nand U3291 (N_3291,In_444,In_1632);
nand U3292 (N_3292,In_511,In_1881);
nand U3293 (N_3293,In_1461,In_975);
and U3294 (N_3294,In_755,In_1744);
nor U3295 (N_3295,In_638,In_871);
nand U3296 (N_3296,In_1033,In_675);
or U3297 (N_3297,In_11,In_1373);
nand U3298 (N_3298,In_1227,In_1745);
or U3299 (N_3299,In_884,In_1675);
or U3300 (N_3300,In_299,In_840);
or U3301 (N_3301,In_512,In_163);
or U3302 (N_3302,In_176,In_1119);
nand U3303 (N_3303,In_35,In_1251);
or U3304 (N_3304,In_953,In_50);
nand U3305 (N_3305,In_1885,In_1045);
nand U3306 (N_3306,In_1545,In_1103);
or U3307 (N_3307,In_844,In_509);
and U3308 (N_3308,In_1623,In_625);
nand U3309 (N_3309,In_1019,In_1300);
or U3310 (N_3310,In_1654,In_987);
nand U3311 (N_3311,In_1397,In_1281);
and U3312 (N_3312,In_839,In_1017);
and U3313 (N_3313,In_82,In_1186);
or U3314 (N_3314,In_229,In_502);
nor U3315 (N_3315,In_1970,In_871);
xnor U3316 (N_3316,In_1497,In_11);
or U3317 (N_3317,In_10,In_882);
nor U3318 (N_3318,In_1213,In_26);
nand U3319 (N_3319,In_395,In_354);
nand U3320 (N_3320,In_1962,In_1985);
xor U3321 (N_3321,In_1871,In_531);
and U3322 (N_3322,In_1504,In_195);
nor U3323 (N_3323,In_1682,In_458);
or U3324 (N_3324,In_765,In_1589);
nand U3325 (N_3325,In_1294,In_521);
nor U3326 (N_3326,In_659,In_676);
or U3327 (N_3327,In_1539,In_482);
nand U3328 (N_3328,In_185,In_1060);
or U3329 (N_3329,In_1435,In_1780);
xor U3330 (N_3330,In_133,In_464);
nand U3331 (N_3331,In_181,In_446);
and U3332 (N_3332,In_1049,In_424);
or U3333 (N_3333,In_1991,In_760);
nor U3334 (N_3334,In_787,In_498);
xnor U3335 (N_3335,In_973,In_970);
and U3336 (N_3336,In_1466,In_821);
nand U3337 (N_3337,In_213,In_1679);
and U3338 (N_3338,In_79,In_571);
nor U3339 (N_3339,In_108,In_1715);
and U3340 (N_3340,In_1851,In_808);
and U3341 (N_3341,In_264,In_636);
and U3342 (N_3342,In_1828,In_341);
nand U3343 (N_3343,In_355,In_142);
nand U3344 (N_3344,In_1084,In_285);
or U3345 (N_3345,In_1751,In_1551);
nand U3346 (N_3346,In_1719,In_90);
and U3347 (N_3347,In_662,In_976);
nor U3348 (N_3348,In_1402,In_1076);
and U3349 (N_3349,In_1539,In_1427);
and U3350 (N_3350,In_368,In_1059);
and U3351 (N_3351,In_1867,In_1204);
or U3352 (N_3352,In_186,In_463);
nor U3353 (N_3353,In_594,In_599);
nor U3354 (N_3354,In_474,In_413);
and U3355 (N_3355,In_298,In_1855);
and U3356 (N_3356,In_1162,In_1725);
nand U3357 (N_3357,In_238,In_376);
or U3358 (N_3358,In_1569,In_1118);
nor U3359 (N_3359,In_284,In_1124);
nand U3360 (N_3360,In_742,In_1431);
or U3361 (N_3361,In_1263,In_596);
or U3362 (N_3362,In_574,In_1388);
xor U3363 (N_3363,In_1477,In_953);
or U3364 (N_3364,In_978,In_739);
xor U3365 (N_3365,In_599,In_1053);
nand U3366 (N_3366,In_560,In_475);
or U3367 (N_3367,In_1390,In_1284);
and U3368 (N_3368,In_1658,In_635);
nand U3369 (N_3369,In_1844,In_24);
nor U3370 (N_3370,In_1730,In_339);
or U3371 (N_3371,In_1852,In_441);
or U3372 (N_3372,In_1594,In_350);
and U3373 (N_3373,In_480,In_1009);
nand U3374 (N_3374,In_1540,In_821);
or U3375 (N_3375,In_1401,In_942);
nand U3376 (N_3376,In_1741,In_83);
nor U3377 (N_3377,In_260,In_482);
nor U3378 (N_3378,In_171,In_1356);
and U3379 (N_3379,In_27,In_560);
nand U3380 (N_3380,In_1252,In_1821);
nand U3381 (N_3381,In_963,In_754);
and U3382 (N_3382,In_464,In_899);
or U3383 (N_3383,In_939,In_755);
and U3384 (N_3384,In_392,In_1191);
nor U3385 (N_3385,In_169,In_145);
and U3386 (N_3386,In_75,In_1235);
nand U3387 (N_3387,In_887,In_907);
or U3388 (N_3388,In_1446,In_947);
nand U3389 (N_3389,In_205,In_162);
or U3390 (N_3390,In_1409,In_1846);
nand U3391 (N_3391,In_1350,In_105);
or U3392 (N_3392,In_1968,In_1916);
nand U3393 (N_3393,In_1580,In_60);
or U3394 (N_3394,In_155,In_306);
nand U3395 (N_3395,In_1238,In_713);
nor U3396 (N_3396,In_504,In_1819);
xnor U3397 (N_3397,In_1450,In_1947);
nand U3398 (N_3398,In_918,In_1101);
and U3399 (N_3399,In_1430,In_1626);
nor U3400 (N_3400,In_1712,In_926);
nand U3401 (N_3401,In_1327,In_1623);
or U3402 (N_3402,In_478,In_81);
or U3403 (N_3403,In_443,In_251);
nor U3404 (N_3404,In_49,In_1379);
nand U3405 (N_3405,In_795,In_1635);
nor U3406 (N_3406,In_1048,In_637);
nand U3407 (N_3407,In_724,In_149);
nand U3408 (N_3408,In_175,In_1345);
or U3409 (N_3409,In_1326,In_932);
or U3410 (N_3410,In_446,In_1410);
nor U3411 (N_3411,In_1625,In_355);
and U3412 (N_3412,In_1456,In_1616);
or U3413 (N_3413,In_1326,In_1844);
or U3414 (N_3414,In_999,In_1686);
nor U3415 (N_3415,In_1646,In_516);
or U3416 (N_3416,In_143,In_782);
nand U3417 (N_3417,In_760,In_674);
or U3418 (N_3418,In_1597,In_1707);
nor U3419 (N_3419,In_1606,In_1296);
and U3420 (N_3420,In_176,In_23);
nand U3421 (N_3421,In_1896,In_761);
and U3422 (N_3422,In_1236,In_1140);
nor U3423 (N_3423,In_1008,In_1003);
or U3424 (N_3424,In_1403,In_1910);
nor U3425 (N_3425,In_734,In_1840);
nor U3426 (N_3426,In_889,In_248);
nor U3427 (N_3427,In_1214,In_705);
nand U3428 (N_3428,In_813,In_1102);
or U3429 (N_3429,In_852,In_713);
nand U3430 (N_3430,In_524,In_1170);
or U3431 (N_3431,In_1192,In_567);
nand U3432 (N_3432,In_1099,In_1098);
and U3433 (N_3433,In_788,In_180);
nor U3434 (N_3434,In_1854,In_1780);
and U3435 (N_3435,In_1069,In_638);
or U3436 (N_3436,In_1517,In_512);
or U3437 (N_3437,In_138,In_234);
and U3438 (N_3438,In_103,In_1546);
and U3439 (N_3439,In_1588,In_1078);
nand U3440 (N_3440,In_1661,In_660);
nor U3441 (N_3441,In_644,In_400);
nor U3442 (N_3442,In_1655,In_94);
nand U3443 (N_3443,In_1243,In_1753);
and U3444 (N_3444,In_1326,In_1174);
nand U3445 (N_3445,In_1628,In_1461);
nand U3446 (N_3446,In_134,In_32);
or U3447 (N_3447,In_588,In_912);
and U3448 (N_3448,In_179,In_1683);
xor U3449 (N_3449,In_1308,In_1686);
nor U3450 (N_3450,In_1490,In_1353);
nor U3451 (N_3451,In_1691,In_921);
nor U3452 (N_3452,In_1751,In_611);
or U3453 (N_3453,In_910,In_1089);
nand U3454 (N_3454,In_88,In_71);
and U3455 (N_3455,In_1158,In_478);
nand U3456 (N_3456,In_426,In_772);
nand U3457 (N_3457,In_923,In_1958);
and U3458 (N_3458,In_591,In_857);
nor U3459 (N_3459,In_1773,In_536);
and U3460 (N_3460,In_662,In_230);
and U3461 (N_3461,In_130,In_1415);
and U3462 (N_3462,In_176,In_1862);
nand U3463 (N_3463,In_1907,In_599);
or U3464 (N_3464,In_1612,In_1168);
and U3465 (N_3465,In_1585,In_37);
nor U3466 (N_3466,In_160,In_1079);
nor U3467 (N_3467,In_1873,In_92);
nand U3468 (N_3468,In_91,In_832);
nor U3469 (N_3469,In_609,In_1300);
or U3470 (N_3470,In_1610,In_573);
xnor U3471 (N_3471,In_1668,In_1825);
nor U3472 (N_3472,In_549,In_42);
and U3473 (N_3473,In_1073,In_536);
nor U3474 (N_3474,In_85,In_259);
and U3475 (N_3475,In_963,In_1231);
and U3476 (N_3476,In_737,In_99);
nor U3477 (N_3477,In_221,In_1957);
nand U3478 (N_3478,In_811,In_1874);
and U3479 (N_3479,In_512,In_1635);
and U3480 (N_3480,In_932,In_1460);
and U3481 (N_3481,In_316,In_169);
xor U3482 (N_3482,In_1318,In_53);
nor U3483 (N_3483,In_1952,In_1649);
and U3484 (N_3484,In_1908,In_881);
and U3485 (N_3485,In_798,In_1891);
and U3486 (N_3486,In_1383,In_536);
or U3487 (N_3487,In_1596,In_78);
nor U3488 (N_3488,In_1090,In_912);
nor U3489 (N_3489,In_137,In_921);
and U3490 (N_3490,In_696,In_768);
and U3491 (N_3491,In_1925,In_1079);
or U3492 (N_3492,In_1682,In_859);
and U3493 (N_3493,In_354,In_1716);
and U3494 (N_3494,In_1627,In_1166);
or U3495 (N_3495,In_971,In_222);
nand U3496 (N_3496,In_284,In_1487);
or U3497 (N_3497,In_1567,In_515);
nor U3498 (N_3498,In_1351,In_464);
or U3499 (N_3499,In_1861,In_924);
nor U3500 (N_3500,In_861,In_916);
and U3501 (N_3501,In_404,In_1718);
nand U3502 (N_3502,In_943,In_524);
nor U3503 (N_3503,In_5,In_437);
nand U3504 (N_3504,In_1595,In_1139);
nor U3505 (N_3505,In_180,In_1757);
or U3506 (N_3506,In_1497,In_407);
xnor U3507 (N_3507,In_1079,In_794);
or U3508 (N_3508,In_1544,In_1339);
nand U3509 (N_3509,In_870,In_204);
and U3510 (N_3510,In_616,In_902);
or U3511 (N_3511,In_213,In_1102);
nor U3512 (N_3512,In_1854,In_1890);
nor U3513 (N_3513,In_856,In_673);
or U3514 (N_3514,In_74,In_272);
nand U3515 (N_3515,In_1631,In_908);
nor U3516 (N_3516,In_1654,In_1964);
and U3517 (N_3517,In_515,In_1358);
or U3518 (N_3518,In_444,In_765);
and U3519 (N_3519,In_528,In_280);
nand U3520 (N_3520,In_1597,In_618);
and U3521 (N_3521,In_605,In_1618);
nand U3522 (N_3522,In_755,In_1748);
nor U3523 (N_3523,In_13,In_525);
and U3524 (N_3524,In_534,In_1951);
and U3525 (N_3525,In_1389,In_1252);
nor U3526 (N_3526,In_375,In_1129);
xnor U3527 (N_3527,In_729,In_1932);
nor U3528 (N_3528,In_1312,In_866);
or U3529 (N_3529,In_17,In_187);
nor U3530 (N_3530,In_1496,In_46);
or U3531 (N_3531,In_1275,In_1693);
and U3532 (N_3532,In_1046,In_605);
or U3533 (N_3533,In_1645,In_1288);
and U3534 (N_3534,In_1962,In_98);
nor U3535 (N_3535,In_891,In_897);
nor U3536 (N_3536,In_1596,In_1960);
nand U3537 (N_3537,In_1979,In_725);
and U3538 (N_3538,In_1500,In_1843);
nor U3539 (N_3539,In_788,In_1644);
and U3540 (N_3540,In_761,In_1716);
nand U3541 (N_3541,In_1023,In_1761);
or U3542 (N_3542,In_434,In_1097);
or U3543 (N_3543,In_1903,In_380);
nor U3544 (N_3544,In_446,In_885);
nor U3545 (N_3545,In_1535,In_1784);
and U3546 (N_3546,In_248,In_1908);
and U3547 (N_3547,In_1445,In_88);
and U3548 (N_3548,In_423,In_18);
nand U3549 (N_3549,In_266,In_1004);
nand U3550 (N_3550,In_192,In_15);
nand U3551 (N_3551,In_1394,In_665);
xnor U3552 (N_3552,In_1157,In_434);
and U3553 (N_3553,In_1795,In_1119);
and U3554 (N_3554,In_739,In_1437);
nand U3555 (N_3555,In_1047,In_871);
nor U3556 (N_3556,In_1193,In_1586);
nand U3557 (N_3557,In_29,In_458);
nor U3558 (N_3558,In_15,In_885);
nand U3559 (N_3559,In_80,In_1677);
nor U3560 (N_3560,In_1401,In_1024);
and U3561 (N_3561,In_1651,In_94);
nand U3562 (N_3562,In_1480,In_30);
nor U3563 (N_3563,In_1605,In_1470);
or U3564 (N_3564,In_873,In_1179);
and U3565 (N_3565,In_1332,In_825);
or U3566 (N_3566,In_1510,In_1974);
nand U3567 (N_3567,In_1484,In_1572);
nor U3568 (N_3568,In_1141,In_1973);
nand U3569 (N_3569,In_253,In_1911);
nor U3570 (N_3570,In_1709,In_1324);
nor U3571 (N_3571,In_1734,In_1700);
nor U3572 (N_3572,In_218,In_1838);
nand U3573 (N_3573,In_26,In_153);
nand U3574 (N_3574,In_1639,In_1388);
nand U3575 (N_3575,In_1838,In_467);
nor U3576 (N_3576,In_1276,In_1710);
and U3577 (N_3577,In_151,In_74);
or U3578 (N_3578,In_1441,In_368);
nor U3579 (N_3579,In_740,In_1584);
and U3580 (N_3580,In_1283,In_1946);
xnor U3581 (N_3581,In_1900,In_43);
nor U3582 (N_3582,In_1271,In_281);
xnor U3583 (N_3583,In_1904,In_618);
nand U3584 (N_3584,In_1171,In_1123);
nand U3585 (N_3585,In_734,In_1178);
xnor U3586 (N_3586,In_702,In_1808);
and U3587 (N_3587,In_1055,In_1392);
or U3588 (N_3588,In_204,In_1590);
and U3589 (N_3589,In_197,In_160);
nand U3590 (N_3590,In_1965,In_538);
or U3591 (N_3591,In_764,In_1905);
nand U3592 (N_3592,In_1794,In_523);
nor U3593 (N_3593,In_291,In_1783);
nand U3594 (N_3594,In_926,In_368);
nand U3595 (N_3595,In_1617,In_785);
and U3596 (N_3596,In_263,In_1990);
nand U3597 (N_3597,In_1421,In_1222);
or U3598 (N_3598,In_621,In_699);
nor U3599 (N_3599,In_62,In_1370);
and U3600 (N_3600,In_1891,In_109);
and U3601 (N_3601,In_1703,In_678);
xor U3602 (N_3602,In_1617,In_815);
nor U3603 (N_3603,In_1992,In_1094);
nor U3604 (N_3604,In_1659,In_75);
and U3605 (N_3605,In_1485,In_1049);
nand U3606 (N_3606,In_1633,In_24);
nand U3607 (N_3607,In_1444,In_235);
nor U3608 (N_3608,In_1551,In_734);
or U3609 (N_3609,In_1241,In_1003);
and U3610 (N_3610,In_1426,In_1902);
or U3611 (N_3611,In_1706,In_1347);
nor U3612 (N_3612,In_777,In_1865);
nand U3613 (N_3613,In_201,In_1324);
nor U3614 (N_3614,In_992,In_1224);
nor U3615 (N_3615,In_1309,In_270);
nor U3616 (N_3616,In_1411,In_487);
nand U3617 (N_3617,In_852,In_1472);
and U3618 (N_3618,In_982,In_985);
nor U3619 (N_3619,In_1695,In_1177);
nand U3620 (N_3620,In_399,In_1430);
nor U3621 (N_3621,In_801,In_749);
or U3622 (N_3622,In_862,In_241);
and U3623 (N_3623,In_376,In_1645);
nor U3624 (N_3624,In_1732,In_1052);
and U3625 (N_3625,In_1607,In_1603);
nand U3626 (N_3626,In_879,In_658);
nand U3627 (N_3627,In_740,In_1057);
or U3628 (N_3628,In_725,In_1197);
or U3629 (N_3629,In_1660,In_340);
nor U3630 (N_3630,In_864,In_1792);
nor U3631 (N_3631,In_1305,In_1727);
nand U3632 (N_3632,In_414,In_1721);
xor U3633 (N_3633,In_1881,In_957);
nand U3634 (N_3634,In_221,In_1655);
or U3635 (N_3635,In_1660,In_1446);
and U3636 (N_3636,In_1657,In_1230);
nand U3637 (N_3637,In_1600,In_1979);
nand U3638 (N_3638,In_1755,In_768);
or U3639 (N_3639,In_356,In_1831);
and U3640 (N_3640,In_878,In_303);
and U3641 (N_3641,In_1191,In_790);
nand U3642 (N_3642,In_1754,In_1912);
nand U3643 (N_3643,In_1672,In_298);
and U3644 (N_3644,In_62,In_1148);
and U3645 (N_3645,In_55,In_1615);
or U3646 (N_3646,In_282,In_1912);
nand U3647 (N_3647,In_572,In_193);
nor U3648 (N_3648,In_923,In_1333);
or U3649 (N_3649,In_1812,In_1814);
xor U3650 (N_3650,In_765,In_917);
nor U3651 (N_3651,In_1137,In_531);
and U3652 (N_3652,In_1422,In_1336);
nand U3653 (N_3653,In_1688,In_1093);
and U3654 (N_3654,In_421,In_809);
nand U3655 (N_3655,In_1055,In_1618);
and U3656 (N_3656,In_1561,In_1919);
nand U3657 (N_3657,In_922,In_474);
and U3658 (N_3658,In_668,In_1595);
and U3659 (N_3659,In_1641,In_708);
nor U3660 (N_3660,In_908,In_1050);
or U3661 (N_3661,In_617,In_223);
nand U3662 (N_3662,In_753,In_581);
or U3663 (N_3663,In_73,In_380);
or U3664 (N_3664,In_368,In_443);
nor U3665 (N_3665,In_1760,In_1279);
nand U3666 (N_3666,In_1054,In_1268);
nand U3667 (N_3667,In_898,In_1980);
nand U3668 (N_3668,In_1345,In_836);
or U3669 (N_3669,In_906,In_244);
nand U3670 (N_3670,In_881,In_1558);
nand U3671 (N_3671,In_652,In_73);
nand U3672 (N_3672,In_1427,In_1640);
nand U3673 (N_3673,In_749,In_776);
nor U3674 (N_3674,In_1944,In_114);
nor U3675 (N_3675,In_1437,In_1043);
and U3676 (N_3676,In_438,In_505);
nand U3677 (N_3677,In_1547,In_796);
or U3678 (N_3678,In_982,In_1737);
xor U3679 (N_3679,In_1188,In_834);
nor U3680 (N_3680,In_1477,In_726);
or U3681 (N_3681,In_1176,In_1210);
nor U3682 (N_3682,In_376,In_1548);
nand U3683 (N_3683,In_645,In_1447);
nand U3684 (N_3684,In_1833,In_1197);
nand U3685 (N_3685,In_1655,In_35);
nor U3686 (N_3686,In_90,In_84);
and U3687 (N_3687,In_1810,In_1045);
or U3688 (N_3688,In_969,In_721);
nand U3689 (N_3689,In_970,In_81);
or U3690 (N_3690,In_1303,In_201);
nand U3691 (N_3691,In_1853,In_861);
nor U3692 (N_3692,In_1705,In_453);
xnor U3693 (N_3693,In_425,In_432);
or U3694 (N_3694,In_340,In_1663);
nor U3695 (N_3695,In_651,In_1985);
or U3696 (N_3696,In_1197,In_1690);
nor U3697 (N_3697,In_22,In_403);
or U3698 (N_3698,In_1688,In_781);
nand U3699 (N_3699,In_708,In_1277);
and U3700 (N_3700,In_490,In_1962);
nor U3701 (N_3701,In_576,In_183);
nor U3702 (N_3702,In_1288,In_461);
nand U3703 (N_3703,In_1003,In_849);
nand U3704 (N_3704,In_822,In_1077);
and U3705 (N_3705,In_323,In_227);
nor U3706 (N_3706,In_1469,In_998);
and U3707 (N_3707,In_795,In_1381);
or U3708 (N_3708,In_356,In_1443);
nand U3709 (N_3709,In_882,In_693);
nor U3710 (N_3710,In_1147,In_1320);
nor U3711 (N_3711,In_301,In_1704);
and U3712 (N_3712,In_969,In_1699);
nand U3713 (N_3713,In_563,In_1690);
and U3714 (N_3714,In_1867,In_1336);
or U3715 (N_3715,In_1942,In_198);
nor U3716 (N_3716,In_684,In_54);
or U3717 (N_3717,In_1476,In_1079);
nand U3718 (N_3718,In_1637,In_1243);
or U3719 (N_3719,In_952,In_797);
or U3720 (N_3720,In_235,In_1196);
and U3721 (N_3721,In_350,In_1652);
or U3722 (N_3722,In_871,In_1617);
and U3723 (N_3723,In_231,In_614);
nand U3724 (N_3724,In_1890,In_1332);
nand U3725 (N_3725,In_893,In_1161);
nand U3726 (N_3726,In_1402,In_1078);
or U3727 (N_3727,In_1678,In_1028);
or U3728 (N_3728,In_1136,In_1850);
or U3729 (N_3729,In_1388,In_1473);
and U3730 (N_3730,In_1345,In_208);
xor U3731 (N_3731,In_1211,In_739);
and U3732 (N_3732,In_1531,In_413);
and U3733 (N_3733,In_262,In_1088);
xnor U3734 (N_3734,In_1371,In_1389);
xnor U3735 (N_3735,In_1769,In_1524);
nor U3736 (N_3736,In_1022,In_316);
or U3737 (N_3737,In_83,In_1104);
or U3738 (N_3738,In_1320,In_750);
or U3739 (N_3739,In_96,In_238);
nor U3740 (N_3740,In_76,In_1404);
and U3741 (N_3741,In_1631,In_1753);
nor U3742 (N_3742,In_537,In_659);
nand U3743 (N_3743,In_659,In_1254);
or U3744 (N_3744,In_1698,In_690);
or U3745 (N_3745,In_1015,In_1198);
and U3746 (N_3746,In_927,In_1470);
or U3747 (N_3747,In_1207,In_1285);
nand U3748 (N_3748,In_1630,In_1537);
nand U3749 (N_3749,In_1746,In_1125);
or U3750 (N_3750,In_1045,In_1957);
nand U3751 (N_3751,In_1357,In_1424);
nor U3752 (N_3752,In_594,In_1104);
and U3753 (N_3753,In_747,In_1527);
or U3754 (N_3754,In_847,In_832);
or U3755 (N_3755,In_1370,In_65);
nand U3756 (N_3756,In_1665,In_614);
xor U3757 (N_3757,In_1752,In_383);
nand U3758 (N_3758,In_1038,In_1345);
or U3759 (N_3759,In_149,In_630);
and U3760 (N_3760,In_1690,In_1791);
or U3761 (N_3761,In_1351,In_827);
or U3762 (N_3762,In_1432,In_488);
or U3763 (N_3763,In_800,In_688);
or U3764 (N_3764,In_142,In_1015);
and U3765 (N_3765,In_1779,In_499);
or U3766 (N_3766,In_184,In_683);
nor U3767 (N_3767,In_107,In_420);
or U3768 (N_3768,In_81,In_848);
or U3769 (N_3769,In_1193,In_1933);
or U3770 (N_3770,In_1291,In_123);
or U3771 (N_3771,In_1539,In_406);
xor U3772 (N_3772,In_1361,In_1117);
and U3773 (N_3773,In_1088,In_451);
or U3774 (N_3774,In_168,In_1368);
and U3775 (N_3775,In_1875,In_1112);
nand U3776 (N_3776,In_1752,In_221);
or U3777 (N_3777,In_148,In_181);
or U3778 (N_3778,In_1088,In_207);
nor U3779 (N_3779,In_1365,In_1391);
nor U3780 (N_3780,In_483,In_834);
or U3781 (N_3781,In_1004,In_343);
and U3782 (N_3782,In_954,In_493);
or U3783 (N_3783,In_334,In_43);
or U3784 (N_3784,In_868,In_1068);
and U3785 (N_3785,In_1548,In_1060);
and U3786 (N_3786,In_1161,In_787);
nor U3787 (N_3787,In_1275,In_1321);
nor U3788 (N_3788,In_149,In_1373);
and U3789 (N_3789,In_1436,In_1359);
nor U3790 (N_3790,In_615,In_325);
or U3791 (N_3791,In_534,In_554);
nor U3792 (N_3792,In_1034,In_873);
and U3793 (N_3793,In_1332,In_990);
or U3794 (N_3794,In_1693,In_1943);
and U3795 (N_3795,In_195,In_345);
nand U3796 (N_3796,In_133,In_1960);
nor U3797 (N_3797,In_1675,In_39);
nor U3798 (N_3798,In_543,In_727);
nand U3799 (N_3799,In_1272,In_880);
nand U3800 (N_3800,In_1015,In_1963);
or U3801 (N_3801,In_1246,In_907);
nand U3802 (N_3802,In_1718,In_1536);
nand U3803 (N_3803,In_776,In_332);
and U3804 (N_3804,In_1129,In_1880);
or U3805 (N_3805,In_159,In_1621);
nor U3806 (N_3806,In_733,In_1808);
nor U3807 (N_3807,In_915,In_86);
and U3808 (N_3808,In_1728,In_412);
or U3809 (N_3809,In_1053,In_1947);
or U3810 (N_3810,In_1759,In_1805);
or U3811 (N_3811,In_445,In_1383);
nor U3812 (N_3812,In_869,In_1243);
nand U3813 (N_3813,In_185,In_1300);
and U3814 (N_3814,In_904,In_133);
or U3815 (N_3815,In_1483,In_646);
and U3816 (N_3816,In_409,In_301);
and U3817 (N_3817,In_691,In_567);
nor U3818 (N_3818,In_862,In_1077);
and U3819 (N_3819,In_1949,In_1618);
nor U3820 (N_3820,In_1255,In_721);
or U3821 (N_3821,In_822,In_173);
and U3822 (N_3822,In_1831,In_413);
nand U3823 (N_3823,In_1209,In_1805);
nor U3824 (N_3824,In_28,In_1117);
nand U3825 (N_3825,In_1440,In_1249);
or U3826 (N_3826,In_1504,In_1466);
and U3827 (N_3827,In_170,In_85);
and U3828 (N_3828,In_584,In_1014);
nand U3829 (N_3829,In_175,In_1682);
nand U3830 (N_3830,In_1998,In_1498);
nor U3831 (N_3831,In_1402,In_1541);
or U3832 (N_3832,In_1249,In_1549);
and U3833 (N_3833,In_1824,In_1525);
and U3834 (N_3834,In_132,In_499);
nand U3835 (N_3835,In_1573,In_706);
or U3836 (N_3836,In_1824,In_12);
nor U3837 (N_3837,In_1838,In_1459);
and U3838 (N_3838,In_1449,In_1725);
nor U3839 (N_3839,In_968,In_639);
or U3840 (N_3840,In_1031,In_1650);
xnor U3841 (N_3841,In_67,In_144);
and U3842 (N_3842,In_355,In_1214);
and U3843 (N_3843,In_857,In_459);
xor U3844 (N_3844,In_1324,In_1020);
nand U3845 (N_3845,In_1832,In_230);
or U3846 (N_3846,In_1961,In_1181);
nor U3847 (N_3847,In_203,In_1461);
or U3848 (N_3848,In_1602,In_180);
and U3849 (N_3849,In_742,In_1102);
nand U3850 (N_3850,In_1898,In_769);
and U3851 (N_3851,In_879,In_1519);
nor U3852 (N_3852,In_1186,In_783);
nor U3853 (N_3853,In_264,In_359);
or U3854 (N_3854,In_1062,In_311);
or U3855 (N_3855,In_76,In_1721);
nand U3856 (N_3856,In_131,In_890);
or U3857 (N_3857,In_1196,In_433);
and U3858 (N_3858,In_182,In_1753);
or U3859 (N_3859,In_95,In_1463);
nor U3860 (N_3860,In_326,In_1421);
xor U3861 (N_3861,In_778,In_1700);
or U3862 (N_3862,In_1883,In_779);
nand U3863 (N_3863,In_1962,In_166);
nand U3864 (N_3864,In_139,In_1086);
and U3865 (N_3865,In_1772,In_770);
nand U3866 (N_3866,In_207,In_220);
nand U3867 (N_3867,In_98,In_588);
nand U3868 (N_3868,In_1503,In_450);
or U3869 (N_3869,In_1657,In_1685);
nand U3870 (N_3870,In_1976,In_397);
and U3871 (N_3871,In_523,In_1676);
and U3872 (N_3872,In_279,In_1225);
nand U3873 (N_3873,In_811,In_1037);
nor U3874 (N_3874,In_32,In_1264);
nand U3875 (N_3875,In_803,In_1447);
and U3876 (N_3876,In_634,In_1035);
nor U3877 (N_3877,In_1441,In_1031);
and U3878 (N_3878,In_24,In_530);
nor U3879 (N_3879,In_1116,In_1596);
or U3880 (N_3880,In_1552,In_800);
or U3881 (N_3881,In_159,In_1429);
nand U3882 (N_3882,In_657,In_854);
and U3883 (N_3883,In_152,In_1423);
nor U3884 (N_3884,In_506,In_1182);
and U3885 (N_3885,In_1307,In_9);
nand U3886 (N_3886,In_1008,In_1076);
and U3887 (N_3887,In_1247,In_857);
nor U3888 (N_3888,In_730,In_1556);
and U3889 (N_3889,In_928,In_709);
or U3890 (N_3890,In_234,In_1692);
nand U3891 (N_3891,In_1780,In_139);
and U3892 (N_3892,In_473,In_1363);
or U3893 (N_3893,In_286,In_549);
or U3894 (N_3894,In_1905,In_1045);
nor U3895 (N_3895,In_68,In_352);
nor U3896 (N_3896,In_819,In_1983);
nor U3897 (N_3897,In_924,In_947);
and U3898 (N_3898,In_197,In_1883);
and U3899 (N_3899,In_1171,In_1858);
and U3900 (N_3900,In_921,In_1421);
xnor U3901 (N_3901,In_1375,In_899);
nand U3902 (N_3902,In_1072,In_647);
or U3903 (N_3903,In_1365,In_3);
and U3904 (N_3904,In_1274,In_920);
nor U3905 (N_3905,In_1944,In_1080);
nand U3906 (N_3906,In_448,In_1039);
nand U3907 (N_3907,In_1296,In_1759);
nor U3908 (N_3908,In_507,In_960);
or U3909 (N_3909,In_1001,In_677);
nor U3910 (N_3910,In_186,In_1107);
nand U3911 (N_3911,In_1593,In_1672);
or U3912 (N_3912,In_1918,In_1432);
and U3913 (N_3913,In_1673,In_835);
nand U3914 (N_3914,In_826,In_1751);
and U3915 (N_3915,In_1871,In_990);
nand U3916 (N_3916,In_1913,In_629);
and U3917 (N_3917,In_1160,In_1379);
nand U3918 (N_3918,In_980,In_1465);
nor U3919 (N_3919,In_1986,In_1935);
nand U3920 (N_3920,In_371,In_1505);
nor U3921 (N_3921,In_1682,In_1262);
or U3922 (N_3922,In_1124,In_1890);
or U3923 (N_3923,In_360,In_1125);
nand U3924 (N_3924,In_222,In_1645);
nor U3925 (N_3925,In_680,In_421);
nand U3926 (N_3926,In_1698,In_839);
nand U3927 (N_3927,In_1193,In_1594);
nand U3928 (N_3928,In_1709,In_7);
nand U3929 (N_3929,In_1879,In_1684);
nor U3930 (N_3930,In_1323,In_26);
nand U3931 (N_3931,In_420,In_517);
nand U3932 (N_3932,In_305,In_889);
nor U3933 (N_3933,In_1113,In_643);
or U3934 (N_3934,In_684,In_1312);
or U3935 (N_3935,In_268,In_293);
and U3936 (N_3936,In_122,In_1254);
nor U3937 (N_3937,In_891,In_1339);
and U3938 (N_3938,In_462,In_1312);
and U3939 (N_3939,In_391,In_1156);
nor U3940 (N_3940,In_1246,In_1136);
nand U3941 (N_3941,In_696,In_1251);
nor U3942 (N_3942,In_1501,In_314);
nand U3943 (N_3943,In_1568,In_1937);
nor U3944 (N_3944,In_558,In_810);
nor U3945 (N_3945,In_1734,In_85);
and U3946 (N_3946,In_201,In_551);
and U3947 (N_3947,In_393,In_1854);
or U3948 (N_3948,In_731,In_1806);
and U3949 (N_3949,In_1793,In_1730);
and U3950 (N_3950,In_881,In_1995);
nand U3951 (N_3951,In_512,In_1378);
or U3952 (N_3952,In_250,In_1456);
or U3953 (N_3953,In_836,In_1023);
nand U3954 (N_3954,In_1270,In_385);
xnor U3955 (N_3955,In_1852,In_417);
nand U3956 (N_3956,In_48,In_1062);
or U3957 (N_3957,In_1402,In_1712);
and U3958 (N_3958,In_452,In_1209);
or U3959 (N_3959,In_171,In_165);
nor U3960 (N_3960,In_955,In_362);
xnor U3961 (N_3961,In_1470,In_1320);
nand U3962 (N_3962,In_1535,In_298);
or U3963 (N_3963,In_1384,In_1674);
or U3964 (N_3964,In_1899,In_1518);
nand U3965 (N_3965,In_1289,In_1265);
nor U3966 (N_3966,In_1631,In_1929);
and U3967 (N_3967,In_1916,In_460);
nand U3968 (N_3968,In_1770,In_1545);
xor U3969 (N_3969,In_1108,In_1740);
or U3970 (N_3970,In_1459,In_1358);
nand U3971 (N_3971,In_215,In_147);
nor U3972 (N_3972,In_1458,In_1934);
nor U3973 (N_3973,In_1096,In_979);
nand U3974 (N_3974,In_1096,In_1618);
and U3975 (N_3975,In_1598,In_1567);
or U3976 (N_3976,In_1950,In_1491);
nor U3977 (N_3977,In_244,In_811);
or U3978 (N_3978,In_511,In_997);
and U3979 (N_3979,In_923,In_139);
nand U3980 (N_3980,In_381,In_1136);
nand U3981 (N_3981,In_904,In_1608);
and U3982 (N_3982,In_1805,In_1106);
nand U3983 (N_3983,In_1372,In_1290);
or U3984 (N_3984,In_1724,In_276);
nor U3985 (N_3985,In_1248,In_1139);
nand U3986 (N_3986,In_1042,In_1251);
or U3987 (N_3987,In_1886,In_1265);
and U3988 (N_3988,In_614,In_1883);
nor U3989 (N_3989,In_1936,In_1792);
nor U3990 (N_3990,In_1631,In_99);
nand U3991 (N_3991,In_529,In_1795);
nand U3992 (N_3992,In_1778,In_648);
nor U3993 (N_3993,In_1576,In_59);
or U3994 (N_3994,In_1170,In_898);
or U3995 (N_3995,In_1227,In_1676);
nand U3996 (N_3996,In_211,In_1982);
nand U3997 (N_3997,In_892,In_1907);
nor U3998 (N_3998,In_680,In_265);
or U3999 (N_3999,In_1016,In_439);
or U4000 (N_4000,In_1848,In_830);
and U4001 (N_4001,In_208,In_1377);
nand U4002 (N_4002,In_990,In_852);
nor U4003 (N_4003,In_222,In_476);
or U4004 (N_4004,In_553,In_897);
nor U4005 (N_4005,In_166,In_1662);
or U4006 (N_4006,In_1661,In_1961);
nor U4007 (N_4007,In_928,In_390);
nor U4008 (N_4008,In_898,In_1446);
or U4009 (N_4009,In_1480,In_616);
nand U4010 (N_4010,In_1598,In_940);
nand U4011 (N_4011,In_1140,In_731);
or U4012 (N_4012,In_1153,In_1870);
nor U4013 (N_4013,In_694,In_394);
nand U4014 (N_4014,In_550,In_1434);
and U4015 (N_4015,In_1489,In_1370);
nor U4016 (N_4016,In_216,In_824);
or U4017 (N_4017,In_1601,In_1725);
or U4018 (N_4018,In_1375,In_891);
and U4019 (N_4019,In_879,In_579);
nor U4020 (N_4020,In_542,In_253);
nand U4021 (N_4021,In_473,In_280);
and U4022 (N_4022,In_1885,In_1636);
nor U4023 (N_4023,In_105,In_1431);
nor U4024 (N_4024,In_1825,In_407);
nand U4025 (N_4025,In_1013,In_656);
nor U4026 (N_4026,In_1788,In_1548);
nor U4027 (N_4027,In_460,In_1595);
or U4028 (N_4028,In_370,In_434);
and U4029 (N_4029,In_732,In_411);
or U4030 (N_4030,In_1774,In_1594);
and U4031 (N_4031,In_818,In_966);
nand U4032 (N_4032,In_1051,In_475);
and U4033 (N_4033,In_818,In_27);
and U4034 (N_4034,In_179,In_1138);
and U4035 (N_4035,In_1631,In_1976);
nor U4036 (N_4036,In_1970,In_1214);
nand U4037 (N_4037,In_1442,In_586);
and U4038 (N_4038,In_1708,In_685);
or U4039 (N_4039,In_121,In_1686);
or U4040 (N_4040,In_1544,In_223);
or U4041 (N_4041,In_666,In_1526);
or U4042 (N_4042,In_1596,In_1279);
or U4043 (N_4043,In_1890,In_265);
nor U4044 (N_4044,In_1292,In_1560);
nor U4045 (N_4045,In_906,In_1644);
and U4046 (N_4046,In_286,In_80);
nor U4047 (N_4047,In_1705,In_1807);
or U4048 (N_4048,In_1255,In_1222);
nand U4049 (N_4049,In_743,In_1124);
nand U4050 (N_4050,In_1761,In_1065);
or U4051 (N_4051,In_1121,In_325);
nor U4052 (N_4052,In_607,In_671);
nor U4053 (N_4053,In_900,In_1700);
or U4054 (N_4054,In_499,In_502);
nor U4055 (N_4055,In_647,In_808);
nor U4056 (N_4056,In_1140,In_1795);
and U4057 (N_4057,In_1964,In_180);
or U4058 (N_4058,In_350,In_559);
or U4059 (N_4059,In_992,In_1290);
nor U4060 (N_4060,In_398,In_1542);
or U4061 (N_4061,In_615,In_1759);
and U4062 (N_4062,In_441,In_336);
nand U4063 (N_4063,In_976,In_467);
nor U4064 (N_4064,In_1396,In_1348);
xnor U4065 (N_4065,In_903,In_1195);
or U4066 (N_4066,In_348,In_1809);
and U4067 (N_4067,In_1959,In_975);
xor U4068 (N_4068,In_96,In_1349);
nor U4069 (N_4069,In_362,In_1678);
or U4070 (N_4070,In_251,In_1707);
nand U4071 (N_4071,In_1529,In_729);
nand U4072 (N_4072,In_1357,In_639);
nand U4073 (N_4073,In_1978,In_1749);
nand U4074 (N_4074,In_1974,In_244);
or U4075 (N_4075,In_1224,In_622);
or U4076 (N_4076,In_1579,In_1828);
or U4077 (N_4077,In_778,In_780);
or U4078 (N_4078,In_737,In_1770);
nor U4079 (N_4079,In_1872,In_345);
nand U4080 (N_4080,In_328,In_584);
or U4081 (N_4081,In_1431,In_1220);
and U4082 (N_4082,In_1413,In_1682);
and U4083 (N_4083,In_1215,In_974);
nor U4084 (N_4084,In_648,In_1828);
and U4085 (N_4085,In_760,In_873);
or U4086 (N_4086,In_1484,In_271);
nor U4087 (N_4087,In_498,In_1937);
and U4088 (N_4088,In_677,In_666);
and U4089 (N_4089,In_1103,In_913);
or U4090 (N_4090,In_138,In_1809);
or U4091 (N_4091,In_955,In_1565);
or U4092 (N_4092,In_484,In_1604);
nor U4093 (N_4093,In_1573,In_539);
and U4094 (N_4094,In_1162,In_1924);
nor U4095 (N_4095,In_702,In_494);
or U4096 (N_4096,In_1184,In_1941);
xor U4097 (N_4097,In_1389,In_1179);
nand U4098 (N_4098,In_528,In_1662);
nor U4099 (N_4099,In_1320,In_1256);
nand U4100 (N_4100,In_404,In_56);
and U4101 (N_4101,In_407,In_1252);
and U4102 (N_4102,In_1609,In_409);
nor U4103 (N_4103,In_1207,In_1640);
or U4104 (N_4104,In_1059,In_1654);
and U4105 (N_4105,In_840,In_1580);
or U4106 (N_4106,In_1196,In_1392);
and U4107 (N_4107,In_217,In_227);
and U4108 (N_4108,In_1473,In_1568);
nor U4109 (N_4109,In_440,In_1279);
or U4110 (N_4110,In_1898,In_777);
or U4111 (N_4111,In_300,In_1454);
and U4112 (N_4112,In_1449,In_1489);
xor U4113 (N_4113,In_75,In_176);
or U4114 (N_4114,In_537,In_845);
and U4115 (N_4115,In_349,In_436);
and U4116 (N_4116,In_1152,In_815);
or U4117 (N_4117,In_413,In_1680);
nand U4118 (N_4118,In_612,In_1478);
and U4119 (N_4119,In_1400,In_651);
nor U4120 (N_4120,In_1060,In_1496);
nor U4121 (N_4121,In_282,In_229);
nor U4122 (N_4122,In_1355,In_5);
nor U4123 (N_4123,In_124,In_362);
nor U4124 (N_4124,In_1379,In_772);
xnor U4125 (N_4125,In_770,In_1056);
nand U4126 (N_4126,In_724,In_901);
or U4127 (N_4127,In_1253,In_304);
and U4128 (N_4128,In_1958,In_1696);
nor U4129 (N_4129,In_174,In_237);
nor U4130 (N_4130,In_475,In_141);
and U4131 (N_4131,In_763,In_98);
and U4132 (N_4132,In_113,In_1930);
nor U4133 (N_4133,In_371,In_327);
and U4134 (N_4134,In_44,In_199);
nor U4135 (N_4135,In_1899,In_733);
nor U4136 (N_4136,In_7,In_532);
and U4137 (N_4137,In_352,In_766);
xor U4138 (N_4138,In_158,In_1129);
and U4139 (N_4139,In_718,In_672);
or U4140 (N_4140,In_806,In_1598);
or U4141 (N_4141,In_730,In_177);
or U4142 (N_4142,In_1578,In_524);
nand U4143 (N_4143,In_924,In_1636);
or U4144 (N_4144,In_220,In_265);
and U4145 (N_4145,In_1736,In_539);
nor U4146 (N_4146,In_1208,In_1637);
nor U4147 (N_4147,In_936,In_1246);
and U4148 (N_4148,In_1321,In_186);
nand U4149 (N_4149,In_1323,In_1969);
or U4150 (N_4150,In_394,In_1906);
or U4151 (N_4151,In_146,In_1180);
nor U4152 (N_4152,In_114,In_1737);
or U4153 (N_4153,In_634,In_1083);
nor U4154 (N_4154,In_1758,In_528);
nand U4155 (N_4155,In_541,In_497);
and U4156 (N_4156,In_1334,In_1967);
nand U4157 (N_4157,In_273,In_1249);
nand U4158 (N_4158,In_619,In_1584);
nand U4159 (N_4159,In_888,In_1587);
nor U4160 (N_4160,In_1936,In_544);
nor U4161 (N_4161,In_1706,In_369);
and U4162 (N_4162,In_1498,In_1794);
nor U4163 (N_4163,In_42,In_1328);
nor U4164 (N_4164,In_629,In_1350);
xor U4165 (N_4165,In_66,In_142);
nor U4166 (N_4166,In_1089,In_1657);
nand U4167 (N_4167,In_457,In_225);
or U4168 (N_4168,In_918,In_1182);
nand U4169 (N_4169,In_16,In_263);
nand U4170 (N_4170,In_1867,In_925);
nand U4171 (N_4171,In_218,In_813);
nand U4172 (N_4172,In_1597,In_1632);
and U4173 (N_4173,In_371,In_14);
or U4174 (N_4174,In_1899,In_187);
nor U4175 (N_4175,In_1716,In_155);
or U4176 (N_4176,In_135,In_1654);
nand U4177 (N_4177,In_148,In_565);
nor U4178 (N_4178,In_814,In_958);
nor U4179 (N_4179,In_1778,In_358);
and U4180 (N_4180,In_713,In_161);
nor U4181 (N_4181,In_196,In_1433);
nand U4182 (N_4182,In_1762,In_548);
or U4183 (N_4183,In_1273,In_1441);
nand U4184 (N_4184,In_74,In_1908);
or U4185 (N_4185,In_507,In_381);
or U4186 (N_4186,In_660,In_1980);
or U4187 (N_4187,In_1429,In_799);
nand U4188 (N_4188,In_1148,In_1600);
or U4189 (N_4189,In_1537,In_950);
nor U4190 (N_4190,In_1779,In_1918);
or U4191 (N_4191,In_1871,In_143);
or U4192 (N_4192,In_501,In_1955);
nor U4193 (N_4193,In_1102,In_918);
and U4194 (N_4194,In_646,In_591);
and U4195 (N_4195,In_1749,In_1650);
and U4196 (N_4196,In_1119,In_210);
nand U4197 (N_4197,In_1150,In_1114);
nand U4198 (N_4198,In_1185,In_1045);
nor U4199 (N_4199,In_716,In_1622);
nor U4200 (N_4200,In_988,In_681);
or U4201 (N_4201,In_1035,In_682);
nand U4202 (N_4202,In_410,In_403);
nand U4203 (N_4203,In_1223,In_424);
nor U4204 (N_4204,In_1630,In_81);
or U4205 (N_4205,In_1338,In_1992);
nand U4206 (N_4206,In_852,In_1678);
or U4207 (N_4207,In_1275,In_1007);
nand U4208 (N_4208,In_1938,In_1633);
or U4209 (N_4209,In_457,In_657);
and U4210 (N_4210,In_1118,In_1091);
or U4211 (N_4211,In_1290,In_1833);
or U4212 (N_4212,In_1332,In_513);
nor U4213 (N_4213,In_477,In_1734);
nand U4214 (N_4214,In_1645,In_335);
and U4215 (N_4215,In_79,In_1456);
nand U4216 (N_4216,In_508,In_946);
nor U4217 (N_4217,In_581,In_1953);
or U4218 (N_4218,In_199,In_1875);
or U4219 (N_4219,In_595,In_545);
or U4220 (N_4220,In_486,In_5);
nand U4221 (N_4221,In_96,In_1932);
or U4222 (N_4222,In_80,In_724);
nor U4223 (N_4223,In_1477,In_266);
or U4224 (N_4224,In_345,In_482);
or U4225 (N_4225,In_258,In_439);
and U4226 (N_4226,In_1834,In_1895);
nand U4227 (N_4227,In_1194,In_1695);
or U4228 (N_4228,In_1907,In_1818);
nor U4229 (N_4229,In_490,In_923);
nand U4230 (N_4230,In_1863,In_335);
or U4231 (N_4231,In_466,In_280);
or U4232 (N_4232,In_139,In_1352);
and U4233 (N_4233,In_198,In_115);
xor U4234 (N_4234,In_18,In_1433);
nor U4235 (N_4235,In_1070,In_1415);
and U4236 (N_4236,In_55,In_702);
nand U4237 (N_4237,In_1671,In_126);
nor U4238 (N_4238,In_1319,In_1447);
nor U4239 (N_4239,In_895,In_371);
and U4240 (N_4240,In_1536,In_1893);
or U4241 (N_4241,In_1311,In_703);
and U4242 (N_4242,In_1567,In_1735);
or U4243 (N_4243,In_903,In_1879);
and U4244 (N_4244,In_255,In_171);
xor U4245 (N_4245,In_1644,In_1617);
or U4246 (N_4246,In_803,In_82);
nand U4247 (N_4247,In_220,In_570);
nand U4248 (N_4248,In_1890,In_1694);
nor U4249 (N_4249,In_1142,In_1740);
and U4250 (N_4250,In_544,In_38);
nand U4251 (N_4251,In_1156,In_1333);
or U4252 (N_4252,In_1111,In_1379);
nor U4253 (N_4253,In_1915,In_1805);
nand U4254 (N_4254,In_976,In_802);
and U4255 (N_4255,In_1235,In_289);
nand U4256 (N_4256,In_504,In_656);
nor U4257 (N_4257,In_1713,In_1710);
or U4258 (N_4258,In_598,In_1358);
nand U4259 (N_4259,In_1515,In_966);
or U4260 (N_4260,In_1309,In_469);
nand U4261 (N_4261,In_774,In_994);
and U4262 (N_4262,In_1847,In_1446);
and U4263 (N_4263,In_261,In_1400);
nor U4264 (N_4264,In_1467,In_1137);
nor U4265 (N_4265,In_1046,In_142);
or U4266 (N_4266,In_454,In_55);
nand U4267 (N_4267,In_1475,In_1630);
or U4268 (N_4268,In_325,In_381);
nor U4269 (N_4269,In_989,In_1806);
nand U4270 (N_4270,In_1857,In_169);
nor U4271 (N_4271,In_68,In_736);
and U4272 (N_4272,In_101,In_1140);
and U4273 (N_4273,In_1475,In_1519);
or U4274 (N_4274,In_924,In_276);
or U4275 (N_4275,In_192,In_476);
nor U4276 (N_4276,In_1939,In_1786);
and U4277 (N_4277,In_1485,In_532);
or U4278 (N_4278,In_1083,In_191);
and U4279 (N_4279,In_1996,In_454);
nand U4280 (N_4280,In_902,In_768);
and U4281 (N_4281,In_187,In_794);
or U4282 (N_4282,In_442,In_772);
or U4283 (N_4283,In_1891,In_1010);
and U4284 (N_4284,In_1823,In_737);
or U4285 (N_4285,In_1987,In_343);
nor U4286 (N_4286,In_1072,In_307);
nand U4287 (N_4287,In_423,In_722);
or U4288 (N_4288,In_282,In_323);
and U4289 (N_4289,In_81,In_845);
nor U4290 (N_4290,In_1062,In_1227);
nand U4291 (N_4291,In_266,In_1201);
or U4292 (N_4292,In_785,In_1940);
nand U4293 (N_4293,In_413,In_298);
nand U4294 (N_4294,In_55,In_1069);
nor U4295 (N_4295,In_1706,In_1789);
and U4296 (N_4296,In_203,In_757);
or U4297 (N_4297,In_1232,In_288);
nor U4298 (N_4298,In_158,In_1449);
nor U4299 (N_4299,In_1003,In_339);
and U4300 (N_4300,In_720,In_831);
nor U4301 (N_4301,In_378,In_272);
nand U4302 (N_4302,In_1212,In_1975);
or U4303 (N_4303,In_1590,In_1116);
nand U4304 (N_4304,In_1462,In_1779);
and U4305 (N_4305,In_841,In_1062);
and U4306 (N_4306,In_810,In_1194);
nand U4307 (N_4307,In_14,In_654);
nand U4308 (N_4308,In_802,In_76);
nor U4309 (N_4309,In_1211,In_1865);
nand U4310 (N_4310,In_435,In_1662);
and U4311 (N_4311,In_442,In_846);
nor U4312 (N_4312,In_1193,In_624);
nand U4313 (N_4313,In_873,In_1945);
nand U4314 (N_4314,In_198,In_422);
and U4315 (N_4315,In_14,In_1645);
or U4316 (N_4316,In_1214,In_998);
xor U4317 (N_4317,In_1434,In_1395);
or U4318 (N_4318,In_379,In_1242);
and U4319 (N_4319,In_42,In_1650);
nand U4320 (N_4320,In_1014,In_252);
nor U4321 (N_4321,In_1311,In_1377);
nand U4322 (N_4322,In_112,In_412);
and U4323 (N_4323,In_1334,In_956);
xnor U4324 (N_4324,In_1929,In_1560);
nand U4325 (N_4325,In_322,In_482);
or U4326 (N_4326,In_1652,In_1780);
nor U4327 (N_4327,In_1984,In_817);
nor U4328 (N_4328,In_707,In_146);
and U4329 (N_4329,In_1982,In_1843);
or U4330 (N_4330,In_1779,In_455);
and U4331 (N_4331,In_766,In_643);
nor U4332 (N_4332,In_965,In_1409);
nor U4333 (N_4333,In_1250,In_1902);
or U4334 (N_4334,In_1630,In_675);
or U4335 (N_4335,In_1695,In_1171);
or U4336 (N_4336,In_539,In_225);
nand U4337 (N_4337,In_1284,In_1325);
and U4338 (N_4338,In_885,In_336);
or U4339 (N_4339,In_1129,In_795);
nand U4340 (N_4340,In_1417,In_262);
nor U4341 (N_4341,In_245,In_1562);
nand U4342 (N_4342,In_437,In_1631);
nand U4343 (N_4343,In_1594,In_1197);
nor U4344 (N_4344,In_1435,In_457);
or U4345 (N_4345,In_960,In_218);
and U4346 (N_4346,In_420,In_475);
or U4347 (N_4347,In_400,In_1139);
nor U4348 (N_4348,In_1759,In_1281);
nand U4349 (N_4349,In_446,In_381);
nor U4350 (N_4350,In_1243,In_279);
xnor U4351 (N_4351,In_677,In_547);
and U4352 (N_4352,In_232,In_1896);
nand U4353 (N_4353,In_877,In_343);
nand U4354 (N_4354,In_742,In_607);
nor U4355 (N_4355,In_639,In_512);
nor U4356 (N_4356,In_1470,In_1417);
nand U4357 (N_4357,In_1674,In_1956);
and U4358 (N_4358,In_1815,In_1698);
nand U4359 (N_4359,In_746,In_429);
or U4360 (N_4360,In_641,In_617);
xor U4361 (N_4361,In_1690,In_1012);
or U4362 (N_4362,In_1979,In_1507);
and U4363 (N_4363,In_192,In_777);
or U4364 (N_4364,In_913,In_605);
or U4365 (N_4365,In_1678,In_127);
and U4366 (N_4366,In_1074,In_1538);
and U4367 (N_4367,In_1074,In_828);
nand U4368 (N_4368,In_1063,In_1613);
and U4369 (N_4369,In_1221,In_1557);
or U4370 (N_4370,In_1193,In_295);
or U4371 (N_4371,In_695,In_140);
nand U4372 (N_4372,In_842,In_1434);
or U4373 (N_4373,In_1052,In_1338);
and U4374 (N_4374,In_959,In_1039);
xor U4375 (N_4375,In_1790,In_1915);
or U4376 (N_4376,In_1385,In_934);
or U4377 (N_4377,In_872,In_403);
or U4378 (N_4378,In_990,In_525);
and U4379 (N_4379,In_1921,In_506);
xnor U4380 (N_4380,In_540,In_1848);
or U4381 (N_4381,In_1917,In_1139);
nor U4382 (N_4382,In_1339,In_1506);
and U4383 (N_4383,In_1259,In_1632);
nor U4384 (N_4384,In_221,In_853);
or U4385 (N_4385,In_937,In_1124);
xor U4386 (N_4386,In_1877,In_164);
nand U4387 (N_4387,In_1173,In_1604);
nor U4388 (N_4388,In_875,In_1237);
nand U4389 (N_4389,In_188,In_1149);
and U4390 (N_4390,In_687,In_1671);
nor U4391 (N_4391,In_226,In_1961);
and U4392 (N_4392,In_1973,In_1093);
or U4393 (N_4393,In_181,In_1239);
and U4394 (N_4394,In_496,In_752);
nor U4395 (N_4395,In_928,In_1243);
and U4396 (N_4396,In_1208,In_108);
or U4397 (N_4397,In_417,In_1195);
nor U4398 (N_4398,In_1868,In_1570);
or U4399 (N_4399,In_1789,In_1499);
xnor U4400 (N_4400,In_1066,In_618);
nor U4401 (N_4401,In_794,In_765);
or U4402 (N_4402,In_223,In_284);
nand U4403 (N_4403,In_618,In_1591);
or U4404 (N_4404,In_1580,In_826);
nor U4405 (N_4405,In_1997,In_1562);
nand U4406 (N_4406,In_244,In_1174);
nor U4407 (N_4407,In_1266,In_197);
or U4408 (N_4408,In_1698,In_620);
nor U4409 (N_4409,In_601,In_1572);
or U4410 (N_4410,In_1306,In_1141);
or U4411 (N_4411,In_424,In_1230);
and U4412 (N_4412,In_1954,In_1098);
nand U4413 (N_4413,In_1804,In_832);
and U4414 (N_4414,In_623,In_1267);
nand U4415 (N_4415,In_218,In_450);
nand U4416 (N_4416,In_1851,In_1157);
and U4417 (N_4417,In_765,In_453);
and U4418 (N_4418,In_805,In_884);
or U4419 (N_4419,In_796,In_365);
nand U4420 (N_4420,In_1743,In_125);
or U4421 (N_4421,In_1825,In_769);
nor U4422 (N_4422,In_655,In_698);
and U4423 (N_4423,In_1648,In_1785);
nor U4424 (N_4424,In_1539,In_1207);
or U4425 (N_4425,In_501,In_211);
and U4426 (N_4426,In_1582,In_1137);
nand U4427 (N_4427,In_1534,In_1938);
nand U4428 (N_4428,In_1821,In_408);
nor U4429 (N_4429,In_527,In_630);
and U4430 (N_4430,In_440,In_1079);
and U4431 (N_4431,In_1353,In_769);
nor U4432 (N_4432,In_1984,In_993);
nor U4433 (N_4433,In_308,In_202);
nor U4434 (N_4434,In_1505,In_713);
or U4435 (N_4435,In_890,In_808);
or U4436 (N_4436,In_326,In_140);
and U4437 (N_4437,In_967,In_455);
nand U4438 (N_4438,In_772,In_58);
xor U4439 (N_4439,In_1344,In_767);
or U4440 (N_4440,In_83,In_1359);
nor U4441 (N_4441,In_224,In_1055);
nand U4442 (N_4442,In_809,In_1343);
or U4443 (N_4443,In_34,In_1096);
nor U4444 (N_4444,In_675,In_1921);
nor U4445 (N_4445,In_913,In_561);
nand U4446 (N_4446,In_744,In_297);
nand U4447 (N_4447,In_589,In_1797);
nor U4448 (N_4448,In_280,In_1738);
nor U4449 (N_4449,In_537,In_639);
nor U4450 (N_4450,In_1125,In_227);
or U4451 (N_4451,In_41,In_348);
nand U4452 (N_4452,In_1098,In_342);
and U4453 (N_4453,In_1618,In_1430);
or U4454 (N_4454,In_235,In_674);
nand U4455 (N_4455,In_1914,In_816);
nand U4456 (N_4456,In_183,In_909);
and U4457 (N_4457,In_1398,In_1532);
nand U4458 (N_4458,In_306,In_517);
xor U4459 (N_4459,In_1823,In_422);
and U4460 (N_4460,In_627,In_1288);
or U4461 (N_4461,In_92,In_657);
or U4462 (N_4462,In_132,In_644);
nor U4463 (N_4463,In_1823,In_1105);
nand U4464 (N_4464,In_1012,In_1538);
nand U4465 (N_4465,In_417,In_1996);
nand U4466 (N_4466,In_1553,In_1942);
nand U4467 (N_4467,In_1388,In_673);
or U4468 (N_4468,In_512,In_906);
and U4469 (N_4469,In_1476,In_1562);
or U4470 (N_4470,In_1861,In_977);
and U4471 (N_4471,In_129,In_1313);
and U4472 (N_4472,In_1701,In_498);
nand U4473 (N_4473,In_483,In_709);
nand U4474 (N_4474,In_1030,In_1409);
and U4475 (N_4475,In_1832,In_1886);
nor U4476 (N_4476,In_1951,In_1497);
and U4477 (N_4477,In_1221,In_899);
or U4478 (N_4478,In_1868,In_808);
nand U4479 (N_4479,In_257,In_622);
nand U4480 (N_4480,In_1299,In_1883);
nor U4481 (N_4481,In_126,In_698);
and U4482 (N_4482,In_115,In_1274);
or U4483 (N_4483,In_614,In_179);
or U4484 (N_4484,In_587,In_574);
nand U4485 (N_4485,In_1358,In_1468);
nand U4486 (N_4486,In_344,In_800);
nor U4487 (N_4487,In_1412,In_1823);
and U4488 (N_4488,In_1635,In_796);
nand U4489 (N_4489,In_726,In_1041);
and U4490 (N_4490,In_301,In_939);
xor U4491 (N_4491,In_68,In_925);
nand U4492 (N_4492,In_997,In_1226);
or U4493 (N_4493,In_601,In_507);
and U4494 (N_4494,In_1232,In_794);
nor U4495 (N_4495,In_1124,In_705);
and U4496 (N_4496,In_1209,In_719);
or U4497 (N_4497,In_1136,In_790);
or U4498 (N_4498,In_1997,In_1668);
or U4499 (N_4499,In_561,In_1929);
or U4500 (N_4500,In_142,In_1980);
nor U4501 (N_4501,In_754,In_855);
and U4502 (N_4502,In_273,In_1436);
nor U4503 (N_4503,In_478,In_432);
nand U4504 (N_4504,In_1712,In_188);
and U4505 (N_4505,In_261,In_889);
nor U4506 (N_4506,In_1021,In_687);
nor U4507 (N_4507,In_697,In_887);
and U4508 (N_4508,In_1312,In_185);
and U4509 (N_4509,In_1596,In_576);
or U4510 (N_4510,In_1494,In_564);
and U4511 (N_4511,In_1501,In_1529);
and U4512 (N_4512,In_968,In_273);
and U4513 (N_4513,In_107,In_1992);
or U4514 (N_4514,In_1512,In_1496);
or U4515 (N_4515,In_630,In_1484);
nand U4516 (N_4516,In_693,In_1512);
or U4517 (N_4517,In_1023,In_367);
or U4518 (N_4518,In_1794,In_970);
nor U4519 (N_4519,In_1372,In_1479);
nor U4520 (N_4520,In_732,In_58);
nand U4521 (N_4521,In_407,In_237);
nand U4522 (N_4522,In_325,In_1622);
xnor U4523 (N_4523,In_1417,In_1782);
or U4524 (N_4524,In_851,In_1624);
or U4525 (N_4525,In_1055,In_522);
or U4526 (N_4526,In_929,In_1044);
nand U4527 (N_4527,In_1570,In_1840);
nand U4528 (N_4528,In_427,In_1281);
or U4529 (N_4529,In_1881,In_31);
nand U4530 (N_4530,In_943,In_1022);
and U4531 (N_4531,In_241,In_1606);
nand U4532 (N_4532,In_499,In_593);
and U4533 (N_4533,In_553,In_405);
and U4534 (N_4534,In_1386,In_890);
nor U4535 (N_4535,In_1336,In_308);
nand U4536 (N_4536,In_1489,In_442);
or U4537 (N_4537,In_1954,In_506);
nand U4538 (N_4538,In_772,In_1183);
or U4539 (N_4539,In_674,In_757);
nand U4540 (N_4540,In_1625,In_1888);
and U4541 (N_4541,In_204,In_736);
and U4542 (N_4542,In_334,In_248);
nor U4543 (N_4543,In_1797,In_1330);
nor U4544 (N_4544,In_1240,In_1980);
nor U4545 (N_4545,In_1485,In_1649);
and U4546 (N_4546,In_1006,In_1716);
or U4547 (N_4547,In_1788,In_713);
and U4548 (N_4548,In_986,In_593);
nor U4549 (N_4549,In_984,In_1618);
and U4550 (N_4550,In_971,In_15);
xor U4551 (N_4551,In_1617,In_203);
nor U4552 (N_4552,In_743,In_268);
or U4553 (N_4553,In_1353,In_608);
nand U4554 (N_4554,In_274,In_1595);
or U4555 (N_4555,In_1846,In_198);
nand U4556 (N_4556,In_303,In_1187);
and U4557 (N_4557,In_1664,In_26);
nor U4558 (N_4558,In_748,In_1961);
nand U4559 (N_4559,In_641,In_152);
nor U4560 (N_4560,In_1865,In_1497);
and U4561 (N_4561,In_1314,In_769);
nor U4562 (N_4562,In_1838,In_1879);
nor U4563 (N_4563,In_431,In_863);
nor U4564 (N_4564,In_1141,In_276);
or U4565 (N_4565,In_1642,In_41);
nand U4566 (N_4566,In_295,In_782);
or U4567 (N_4567,In_1045,In_450);
or U4568 (N_4568,In_752,In_1587);
nor U4569 (N_4569,In_421,In_1909);
or U4570 (N_4570,In_732,In_1651);
and U4571 (N_4571,In_1351,In_1401);
and U4572 (N_4572,In_614,In_27);
nand U4573 (N_4573,In_508,In_162);
nand U4574 (N_4574,In_1656,In_77);
and U4575 (N_4575,In_1078,In_696);
nor U4576 (N_4576,In_794,In_1074);
nand U4577 (N_4577,In_1278,In_938);
and U4578 (N_4578,In_74,In_1002);
nand U4579 (N_4579,In_340,In_1927);
nor U4580 (N_4580,In_648,In_679);
xor U4581 (N_4581,In_786,In_1820);
or U4582 (N_4582,In_1825,In_291);
nand U4583 (N_4583,In_597,In_1984);
nand U4584 (N_4584,In_828,In_168);
and U4585 (N_4585,In_857,In_761);
nand U4586 (N_4586,In_1704,In_691);
nand U4587 (N_4587,In_541,In_1583);
nand U4588 (N_4588,In_1618,In_400);
nand U4589 (N_4589,In_987,In_871);
xor U4590 (N_4590,In_1284,In_589);
or U4591 (N_4591,In_1559,In_1145);
and U4592 (N_4592,In_1575,In_567);
nor U4593 (N_4593,In_1275,In_748);
and U4594 (N_4594,In_1492,In_921);
nand U4595 (N_4595,In_364,In_357);
nor U4596 (N_4596,In_1120,In_1054);
and U4597 (N_4597,In_1258,In_139);
and U4598 (N_4598,In_396,In_1866);
or U4599 (N_4599,In_867,In_974);
nand U4600 (N_4600,In_674,In_1030);
xor U4601 (N_4601,In_774,In_1722);
nor U4602 (N_4602,In_394,In_1575);
nor U4603 (N_4603,In_507,In_801);
or U4604 (N_4604,In_751,In_383);
nor U4605 (N_4605,In_327,In_1971);
or U4606 (N_4606,In_1542,In_803);
and U4607 (N_4607,In_1292,In_1172);
nor U4608 (N_4608,In_1613,In_944);
and U4609 (N_4609,In_906,In_990);
xor U4610 (N_4610,In_989,In_1374);
nand U4611 (N_4611,In_1431,In_1992);
or U4612 (N_4612,In_1962,In_885);
nor U4613 (N_4613,In_512,In_949);
nand U4614 (N_4614,In_1126,In_904);
nand U4615 (N_4615,In_298,In_1050);
nand U4616 (N_4616,In_245,In_1240);
or U4617 (N_4617,In_195,In_1905);
nand U4618 (N_4618,In_698,In_1654);
and U4619 (N_4619,In_1972,In_703);
or U4620 (N_4620,In_262,In_1637);
and U4621 (N_4621,In_323,In_77);
or U4622 (N_4622,In_789,In_972);
nand U4623 (N_4623,In_37,In_1406);
and U4624 (N_4624,In_1904,In_193);
or U4625 (N_4625,In_194,In_203);
or U4626 (N_4626,In_1836,In_454);
and U4627 (N_4627,In_845,In_1196);
nor U4628 (N_4628,In_654,In_1071);
and U4629 (N_4629,In_1595,In_155);
or U4630 (N_4630,In_324,In_680);
nor U4631 (N_4631,In_1259,In_1182);
nand U4632 (N_4632,In_540,In_8);
and U4633 (N_4633,In_615,In_1708);
or U4634 (N_4634,In_1312,In_659);
nand U4635 (N_4635,In_1991,In_26);
nand U4636 (N_4636,In_872,In_173);
nand U4637 (N_4637,In_1699,In_433);
xor U4638 (N_4638,In_155,In_1208);
nand U4639 (N_4639,In_2,In_16);
nor U4640 (N_4640,In_1035,In_373);
xnor U4641 (N_4641,In_285,In_1125);
nand U4642 (N_4642,In_1904,In_76);
nor U4643 (N_4643,In_739,In_1986);
nor U4644 (N_4644,In_1957,In_1163);
or U4645 (N_4645,In_331,In_160);
and U4646 (N_4646,In_1493,In_113);
nor U4647 (N_4647,In_992,In_1465);
or U4648 (N_4648,In_146,In_1434);
or U4649 (N_4649,In_1415,In_1487);
nand U4650 (N_4650,In_56,In_1198);
nand U4651 (N_4651,In_10,In_1339);
nor U4652 (N_4652,In_1349,In_369);
nor U4653 (N_4653,In_654,In_434);
and U4654 (N_4654,In_1328,In_1339);
nand U4655 (N_4655,In_883,In_1498);
and U4656 (N_4656,In_1869,In_457);
or U4657 (N_4657,In_1645,In_1808);
nand U4658 (N_4658,In_1656,In_319);
nand U4659 (N_4659,In_347,In_1383);
xnor U4660 (N_4660,In_759,In_1796);
or U4661 (N_4661,In_1225,In_649);
or U4662 (N_4662,In_278,In_883);
or U4663 (N_4663,In_933,In_1791);
and U4664 (N_4664,In_1011,In_765);
nand U4665 (N_4665,In_1298,In_876);
and U4666 (N_4666,In_404,In_1625);
nor U4667 (N_4667,In_1113,In_349);
and U4668 (N_4668,In_581,In_1437);
or U4669 (N_4669,In_1453,In_182);
or U4670 (N_4670,In_1099,In_388);
nand U4671 (N_4671,In_167,In_1959);
nor U4672 (N_4672,In_205,In_679);
or U4673 (N_4673,In_105,In_220);
or U4674 (N_4674,In_778,In_1232);
or U4675 (N_4675,In_1037,In_88);
nand U4676 (N_4676,In_871,In_1154);
nor U4677 (N_4677,In_718,In_927);
nor U4678 (N_4678,In_349,In_512);
or U4679 (N_4679,In_1786,In_644);
nand U4680 (N_4680,In_1225,In_432);
or U4681 (N_4681,In_880,In_516);
nand U4682 (N_4682,In_536,In_1335);
and U4683 (N_4683,In_554,In_1438);
and U4684 (N_4684,In_277,In_1432);
and U4685 (N_4685,In_1878,In_91);
nor U4686 (N_4686,In_1728,In_803);
nor U4687 (N_4687,In_155,In_1008);
nand U4688 (N_4688,In_555,In_1046);
nand U4689 (N_4689,In_509,In_1420);
nor U4690 (N_4690,In_1591,In_505);
nand U4691 (N_4691,In_72,In_1936);
and U4692 (N_4692,In_312,In_1533);
and U4693 (N_4693,In_736,In_1036);
nand U4694 (N_4694,In_1650,In_193);
nand U4695 (N_4695,In_1134,In_148);
nor U4696 (N_4696,In_1667,In_1994);
and U4697 (N_4697,In_883,In_1881);
nor U4698 (N_4698,In_701,In_1981);
and U4699 (N_4699,In_1469,In_709);
nor U4700 (N_4700,In_704,In_1887);
nand U4701 (N_4701,In_1165,In_1979);
nor U4702 (N_4702,In_865,In_1016);
nand U4703 (N_4703,In_1107,In_1688);
or U4704 (N_4704,In_1980,In_392);
nand U4705 (N_4705,In_1236,In_237);
nor U4706 (N_4706,In_473,In_1025);
nand U4707 (N_4707,In_1748,In_224);
nor U4708 (N_4708,In_980,In_478);
nor U4709 (N_4709,In_264,In_1497);
nand U4710 (N_4710,In_1459,In_1230);
nor U4711 (N_4711,In_288,In_1621);
nand U4712 (N_4712,In_1962,In_946);
nand U4713 (N_4713,In_1350,In_1204);
or U4714 (N_4714,In_749,In_1869);
nand U4715 (N_4715,In_1785,In_1981);
or U4716 (N_4716,In_1952,In_1884);
nor U4717 (N_4717,In_806,In_1500);
and U4718 (N_4718,In_111,In_1967);
nor U4719 (N_4719,In_746,In_872);
and U4720 (N_4720,In_1797,In_1518);
nand U4721 (N_4721,In_367,In_1105);
or U4722 (N_4722,In_1323,In_1813);
nor U4723 (N_4723,In_1869,In_916);
and U4724 (N_4724,In_1357,In_1367);
and U4725 (N_4725,In_415,In_231);
and U4726 (N_4726,In_1481,In_271);
and U4727 (N_4727,In_322,In_1175);
and U4728 (N_4728,In_423,In_1635);
nand U4729 (N_4729,In_1944,In_172);
or U4730 (N_4730,In_510,In_1211);
nand U4731 (N_4731,In_576,In_1976);
nor U4732 (N_4732,In_261,In_536);
nor U4733 (N_4733,In_1629,In_958);
nand U4734 (N_4734,In_1985,In_642);
and U4735 (N_4735,In_1905,In_1845);
nand U4736 (N_4736,In_1545,In_1144);
nand U4737 (N_4737,In_614,In_1005);
nand U4738 (N_4738,In_166,In_697);
and U4739 (N_4739,In_1566,In_525);
and U4740 (N_4740,In_1688,In_1682);
or U4741 (N_4741,In_721,In_1920);
or U4742 (N_4742,In_445,In_169);
or U4743 (N_4743,In_528,In_480);
nand U4744 (N_4744,In_192,In_746);
and U4745 (N_4745,In_485,In_1449);
nor U4746 (N_4746,In_617,In_135);
nor U4747 (N_4747,In_786,In_1348);
or U4748 (N_4748,In_824,In_1156);
or U4749 (N_4749,In_1797,In_1264);
nor U4750 (N_4750,In_1278,In_348);
nor U4751 (N_4751,In_848,In_338);
nand U4752 (N_4752,In_455,In_678);
nand U4753 (N_4753,In_916,In_1487);
nand U4754 (N_4754,In_1908,In_354);
and U4755 (N_4755,In_589,In_660);
xor U4756 (N_4756,In_1209,In_1617);
or U4757 (N_4757,In_1396,In_273);
nor U4758 (N_4758,In_1309,In_1539);
nor U4759 (N_4759,In_102,In_959);
and U4760 (N_4760,In_772,In_817);
xor U4761 (N_4761,In_1610,In_373);
and U4762 (N_4762,In_1981,In_638);
nand U4763 (N_4763,In_1477,In_825);
and U4764 (N_4764,In_1394,In_1462);
nand U4765 (N_4765,In_819,In_1739);
nor U4766 (N_4766,In_164,In_1040);
and U4767 (N_4767,In_1003,In_335);
or U4768 (N_4768,In_1361,In_1266);
nand U4769 (N_4769,In_338,In_893);
nor U4770 (N_4770,In_1709,In_1235);
nor U4771 (N_4771,In_1176,In_1683);
and U4772 (N_4772,In_220,In_276);
or U4773 (N_4773,In_1340,In_220);
nand U4774 (N_4774,In_754,In_978);
nand U4775 (N_4775,In_791,In_1388);
nor U4776 (N_4776,In_1908,In_1555);
nor U4777 (N_4777,In_1638,In_1391);
and U4778 (N_4778,In_838,In_898);
and U4779 (N_4779,In_1379,In_1782);
xor U4780 (N_4780,In_1304,In_605);
nor U4781 (N_4781,In_1282,In_629);
nand U4782 (N_4782,In_539,In_1964);
and U4783 (N_4783,In_1638,In_1200);
or U4784 (N_4784,In_515,In_264);
or U4785 (N_4785,In_339,In_1506);
and U4786 (N_4786,In_100,In_1155);
nand U4787 (N_4787,In_1056,In_1914);
or U4788 (N_4788,In_611,In_1919);
nand U4789 (N_4789,In_641,In_1386);
xnor U4790 (N_4790,In_527,In_718);
and U4791 (N_4791,In_1207,In_1637);
nand U4792 (N_4792,In_1025,In_1359);
nand U4793 (N_4793,In_1367,In_330);
nor U4794 (N_4794,In_1760,In_621);
and U4795 (N_4795,In_1923,In_488);
nor U4796 (N_4796,In_1561,In_1113);
nand U4797 (N_4797,In_1666,In_650);
nand U4798 (N_4798,In_1305,In_1179);
or U4799 (N_4799,In_978,In_1277);
or U4800 (N_4800,In_1063,In_1387);
or U4801 (N_4801,In_1651,In_306);
and U4802 (N_4802,In_624,In_1280);
or U4803 (N_4803,In_175,In_557);
nor U4804 (N_4804,In_1799,In_256);
and U4805 (N_4805,In_454,In_1206);
nand U4806 (N_4806,In_1117,In_347);
nor U4807 (N_4807,In_1878,In_1204);
or U4808 (N_4808,In_202,In_500);
or U4809 (N_4809,In_1232,In_1469);
or U4810 (N_4810,In_479,In_747);
and U4811 (N_4811,In_1685,In_327);
nor U4812 (N_4812,In_1447,In_1644);
nor U4813 (N_4813,In_757,In_113);
and U4814 (N_4814,In_1906,In_522);
nor U4815 (N_4815,In_1900,In_1886);
nor U4816 (N_4816,In_346,In_1534);
or U4817 (N_4817,In_875,In_556);
nand U4818 (N_4818,In_1294,In_122);
or U4819 (N_4819,In_1499,In_1884);
or U4820 (N_4820,In_1802,In_1893);
nor U4821 (N_4821,In_77,In_1126);
or U4822 (N_4822,In_548,In_852);
and U4823 (N_4823,In_227,In_1901);
or U4824 (N_4824,In_1649,In_1248);
xnor U4825 (N_4825,In_651,In_1449);
nand U4826 (N_4826,In_1195,In_302);
and U4827 (N_4827,In_789,In_1186);
nand U4828 (N_4828,In_772,In_929);
and U4829 (N_4829,In_728,In_877);
nand U4830 (N_4830,In_328,In_1675);
or U4831 (N_4831,In_1115,In_1467);
or U4832 (N_4832,In_1536,In_514);
nor U4833 (N_4833,In_175,In_1023);
nand U4834 (N_4834,In_1373,In_66);
nor U4835 (N_4835,In_1991,In_252);
nor U4836 (N_4836,In_112,In_466);
or U4837 (N_4837,In_544,In_484);
nor U4838 (N_4838,In_1104,In_908);
nand U4839 (N_4839,In_1058,In_1800);
or U4840 (N_4840,In_1830,In_791);
nand U4841 (N_4841,In_1410,In_505);
and U4842 (N_4842,In_1377,In_1252);
and U4843 (N_4843,In_1442,In_823);
and U4844 (N_4844,In_1532,In_834);
and U4845 (N_4845,In_1166,In_203);
and U4846 (N_4846,In_118,In_696);
and U4847 (N_4847,In_518,In_1115);
nand U4848 (N_4848,In_1220,In_295);
and U4849 (N_4849,In_1451,In_885);
nand U4850 (N_4850,In_914,In_706);
nor U4851 (N_4851,In_1333,In_1061);
nor U4852 (N_4852,In_367,In_586);
nor U4853 (N_4853,In_575,In_1048);
or U4854 (N_4854,In_904,In_1480);
nor U4855 (N_4855,In_1806,In_834);
nor U4856 (N_4856,In_21,In_1942);
nand U4857 (N_4857,In_1473,In_212);
nand U4858 (N_4858,In_1586,In_64);
or U4859 (N_4859,In_1276,In_399);
or U4860 (N_4860,In_546,In_492);
or U4861 (N_4861,In_1733,In_1057);
nor U4862 (N_4862,In_581,In_1281);
and U4863 (N_4863,In_1636,In_926);
and U4864 (N_4864,In_491,In_1106);
nand U4865 (N_4865,In_1929,In_203);
or U4866 (N_4866,In_1317,In_1846);
or U4867 (N_4867,In_1275,In_172);
nand U4868 (N_4868,In_1071,In_1250);
and U4869 (N_4869,In_1715,In_491);
or U4870 (N_4870,In_905,In_1030);
nand U4871 (N_4871,In_1283,In_1136);
and U4872 (N_4872,In_194,In_1973);
or U4873 (N_4873,In_913,In_712);
and U4874 (N_4874,In_942,In_486);
and U4875 (N_4875,In_1144,In_999);
and U4876 (N_4876,In_540,In_448);
or U4877 (N_4877,In_1804,In_47);
or U4878 (N_4878,In_1576,In_1180);
nand U4879 (N_4879,In_885,In_1781);
nor U4880 (N_4880,In_742,In_444);
and U4881 (N_4881,In_636,In_979);
nand U4882 (N_4882,In_1950,In_496);
and U4883 (N_4883,In_1100,In_1652);
nand U4884 (N_4884,In_704,In_653);
or U4885 (N_4885,In_616,In_179);
nand U4886 (N_4886,In_78,In_456);
nor U4887 (N_4887,In_1323,In_1203);
nor U4888 (N_4888,In_868,In_1921);
and U4889 (N_4889,In_1117,In_1769);
or U4890 (N_4890,In_1643,In_1205);
nor U4891 (N_4891,In_1261,In_1349);
nand U4892 (N_4892,In_4,In_841);
nand U4893 (N_4893,In_430,In_1505);
and U4894 (N_4894,In_1274,In_989);
nor U4895 (N_4895,In_1269,In_1902);
nor U4896 (N_4896,In_1349,In_1552);
nand U4897 (N_4897,In_1426,In_290);
and U4898 (N_4898,In_1932,In_1358);
or U4899 (N_4899,In_1249,In_1726);
and U4900 (N_4900,In_176,In_1598);
nor U4901 (N_4901,In_772,In_22);
nand U4902 (N_4902,In_1134,In_547);
xnor U4903 (N_4903,In_431,In_1005);
and U4904 (N_4904,In_1514,In_592);
nor U4905 (N_4905,In_77,In_1224);
and U4906 (N_4906,In_1489,In_1858);
nand U4907 (N_4907,In_567,In_1381);
nor U4908 (N_4908,In_1259,In_205);
and U4909 (N_4909,In_1004,In_794);
or U4910 (N_4910,In_1406,In_430);
nand U4911 (N_4911,In_1860,In_737);
or U4912 (N_4912,In_1652,In_143);
or U4913 (N_4913,In_842,In_816);
nand U4914 (N_4914,In_1967,In_607);
nor U4915 (N_4915,In_1535,In_1063);
nor U4916 (N_4916,In_826,In_1979);
nor U4917 (N_4917,In_1222,In_908);
or U4918 (N_4918,In_1877,In_927);
and U4919 (N_4919,In_725,In_1279);
and U4920 (N_4920,In_255,In_1774);
nor U4921 (N_4921,In_1623,In_394);
or U4922 (N_4922,In_826,In_1041);
and U4923 (N_4923,In_445,In_1984);
nand U4924 (N_4924,In_1924,In_774);
and U4925 (N_4925,In_1767,In_1287);
nand U4926 (N_4926,In_113,In_1352);
nand U4927 (N_4927,In_95,In_857);
nor U4928 (N_4928,In_1919,In_474);
nor U4929 (N_4929,In_1294,In_1768);
nand U4930 (N_4930,In_1510,In_1395);
and U4931 (N_4931,In_1190,In_97);
nand U4932 (N_4932,In_1710,In_623);
nand U4933 (N_4933,In_1287,In_1897);
or U4934 (N_4934,In_918,In_312);
nand U4935 (N_4935,In_915,In_610);
or U4936 (N_4936,In_650,In_516);
xor U4937 (N_4937,In_967,In_1563);
and U4938 (N_4938,In_629,In_538);
nor U4939 (N_4939,In_1231,In_396);
nor U4940 (N_4940,In_469,In_1173);
nor U4941 (N_4941,In_1338,In_583);
and U4942 (N_4942,In_988,In_1311);
and U4943 (N_4943,In_568,In_1595);
nand U4944 (N_4944,In_1906,In_1025);
nor U4945 (N_4945,In_756,In_555);
nand U4946 (N_4946,In_949,In_865);
and U4947 (N_4947,In_1068,In_69);
nand U4948 (N_4948,In_1877,In_808);
or U4949 (N_4949,In_201,In_214);
and U4950 (N_4950,In_463,In_1049);
or U4951 (N_4951,In_1527,In_219);
nand U4952 (N_4952,In_228,In_1310);
nand U4953 (N_4953,In_1375,In_1205);
or U4954 (N_4954,In_1672,In_1244);
or U4955 (N_4955,In_274,In_1329);
and U4956 (N_4956,In_668,In_1583);
nor U4957 (N_4957,In_397,In_1243);
nor U4958 (N_4958,In_110,In_1363);
nor U4959 (N_4959,In_894,In_173);
and U4960 (N_4960,In_956,In_1760);
or U4961 (N_4961,In_1531,In_827);
nor U4962 (N_4962,In_328,In_848);
and U4963 (N_4963,In_420,In_752);
nand U4964 (N_4964,In_624,In_1591);
and U4965 (N_4965,In_1594,In_1411);
nor U4966 (N_4966,In_186,In_1442);
nand U4967 (N_4967,In_834,In_1607);
and U4968 (N_4968,In_387,In_1326);
and U4969 (N_4969,In_1804,In_1632);
and U4970 (N_4970,In_987,In_1289);
nor U4971 (N_4971,In_634,In_71);
or U4972 (N_4972,In_1098,In_1307);
nand U4973 (N_4973,In_172,In_259);
nand U4974 (N_4974,In_1817,In_1791);
xnor U4975 (N_4975,In_730,In_529);
and U4976 (N_4976,In_1716,In_1848);
or U4977 (N_4977,In_761,In_1257);
nand U4978 (N_4978,In_165,In_744);
nand U4979 (N_4979,In_1910,In_200);
or U4980 (N_4980,In_1920,In_383);
and U4981 (N_4981,In_113,In_1002);
or U4982 (N_4982,In_1948,In_1410);
or U4983 (N_4983,In_1054,In_1617);
or U4984 (N_4984,In_319,In_1665);
nor U4985 (N_4985,In_638,In_1155);
nand U4986 (N_4986,In_1541,In_260);
and U4987 (N_4987,In_626,In_1034);
or U4988 (N_4988,In_1748,In_1072);
nand U4989 (N_4989,In_973,In_1461);
or U4990 (N_4990,In_1757,In_248);
nor U4991 (N_4991,In_934,In_1137);
xor U4992 (N_4992,In_1078,In_1830);
and U4993 (N_4993,In_125,In_1662);
or U4994 (N_4994,In_1394,In_1717);
or U4995 (N_4995,In_1888,In_1153);
and U4996 (N_4996,In_241,In_1553);
nand U4997 (N_4997,In_1433,In_440);
or U4998 (N_4998,In_259,In_251);
nor U4999 (N_4999,In_1967,In_1217);
or U5000 (N_5000,N_3435,N_4039);
and U5001 (N_5001,N_4562,N_3605);
nor U5002 (N_5002,N_1321,N_2052);
or U5003 (N_5003,N_2661,N_706);
or U5004 (N_5004,N_1331,N_349);
and U5005 (N_5005,N_1696,N_303);
or U5006 (N_5006,N_1698,N_1328);
nor U5007 (N_5007,N_2077,N_3464);
or U5008 (N_5008,N_4935,N_3453);
nand U5009 (N_5009,N_1621,N_2852);
nand U5010 (N_5010,N_4590,N_1928);
nand U5011 (N_5011,N_2873,N_2486);
nand U5012 (N_5012,N_4297,N_1388);
nand U5013 (N_5013,N_4051,N_3906);
nor U5014 (N_5014,N_528,N_1820);
and U5015 (N_5015,N_3897,N_604);
and U5016 (N_5016,N_533,N_748);
or U5017 (N_5017,N_2903,N_4691);
nand U5018 (N_5018,N_3245,N_3493);
nand U5019 (N_5019,N_1299,N_880);
and U5020 (N_5020,N_4711,N_4632);
or U5021 (N_5021,N_1064,N_925);
nor U5022 (N_5022,N_4263,N_3063);
nor U5023 (N_5023,N_685,N_3615);
nand U5024 (N_5024,N_832,N_4098);
nor U5025 (N_5025,N_1508,N_1493);
or U5026 (N_5026,N_3239,N_6);
nand U5027 (N_5027,N_301,N_2654);
nor U5028 (N_5028,N_2612,N_707);
and U5029 (N_5029,N_776,N_508);
nor U5030 (N_5030,N_3325,N_3940);
nor U5031 (N_5031,N_1226,N_2437);
or U5032 (N_5032,N_479,N_994);
or U5033 (N_5033,N_1941,N_1778);
nor U5034 (N_5034,N_1609,N_4316);
nor U5035 (N_5035,N_778,N_3002);
nand U5036 (N_5036,N_2453,N_3027);
nor U5037 (N_5037,N_518,N_3543);
nand U5038 (N_5038,N_3960,N_4778);
or U5039 (N_5039,N_2834,N_141);
or U5040 (N_5040,N_3748,N_1398);
or U5041 (N_5041,N_1133,N_4653);
and U5042 (N_5042,N_329,N_2559);
nand U5043 (N_5043,N_4492,N_4);
and U5044 (N_5044,N_1425,N_1247);
or U5045 (N_5045,N_784,N_2408);
and U5046 (N_5046,N_705,N_1402);
or U5047 (N_5047,N_2219,N_771);
nor U5048 (N_5048,N_1374,N_2091);
nand U5049 (N_5049,N_3875,N_1480);
nand U5050 (N_5050,N_1992,N_1617);
nand U5051 (N_5051,N_3070,N_3877);
nor U5052 (N_5052,N_3934,N_289);
and U5053 (N_5053,N_3354,N_4859);
or U5054 (N_5054,N_2829,N_215);
nand U5055 (N_5055,N_4088,N_4640);
or U5056 (N_5056,N_3386,N_4615);
and U5057 (N_5057,N_2763,N_869);
and U5058 (N_5058,N_4800,N_599);
nand U5059 (N_5059,N_1701,N_4998);
or U5060 (N_5060,N_2444,N_1918);
nand U5061 (N_5061,N_2622,N_905);
or U5062 (N_5062,N_4693,N_1187);
or U5063 (N_5063,N_2516,N_4795);
and U5064 (N_5064,N_4147,N_2773);
and U5065 (N_5065,N_4558,N_2276);
and U5066 (N_5066,N_1025,N_4247);
nor U5067 (N_5067,N_3333,N_722);
xnor U5068 (N_5068,N_4471,N_69);
nand U5069 (N_5069,N_4864,N_1189);
nor U5070 (N_5070,N_3633,N_4125);
nand U5071 (N_5071,N_4746,N_3872);
nor U5072 (N_5072,N_3620,N_4612);
or U5073 (N_5073,N_4172,N_3350);
and U5074 (N_5074,N_3943,N_4504);
nand U5075 (N_5075,N_2623,N_2391);
nand U5076 (N_5076,N_4973,N_3219);
or U5077 (N_5077,N_1379,N_4611);
and U5078 (N_5078,N_4194,N_1304);
or U5079 (N_5079,N_1969,N_98);
nor U5080 (N_5080,N_2495,N_1573);
and U5081 (N_5081,N_3295,N_1177);
or U5082 (N_5082,N_4095,N_2421);
nand U5083 (N_5083,N_1434,N_2772);
or U5084 (N_5084,N_1682,N_4610);
nor U5085 (N_5085,N_2123,N_3418);
or U5086 (N_5086,N_3792,N_2449);
nor U5087 (N_5087,N_1768,N_2619);
nand U5088 (N_5088,N_4774,N_4828);
and U5089 (N_5089,N_4390,N_836);
nor U5090 (N_5090,N_4292,N_3876);
or U5091 (N_5091,N_696,N_164);
and U5092 (N_5092,N_2196,N_2618);
nor U5093 (N_5093,N_2350,N_1399);
or U5094 (N_5094,N_2036,N_1950);
and U5095 (N_5095,N_3126,N_4555);
nand U5096 (N_5096,N_3360,N_3226);
and U5097 (N_5097,N_2053,N_2303);
and U5098 (N_5098,N_2041,N_1806);
and U5099 (N_5099,N_1454,N_4667);
and U5100 (N_5100,N_4265,N_1043);
nand U5101 (N_5101,N_3162,N_2329);
nor U5102 (N_5102,N_4344,N_4449);
nand U5103 (N_5103,N_4279,N_1515);
nor U5104 (N_5104,N_4979,N_3924);
and U5105 (N_5105,N_2293,N_473);
nor U5106 (N_5106,N_1579,N_4835);
nor U5107 (N_5107,N_2716,N_4284);
and U5108 (N_5108,N_4818,N_2318);
xnor U5109 (N_5109,N_2592,N_2469);
nand U5110 (N_5110,N_4443,N_3703);
nor U5111 (N_5111,N_3883,N_1156);
and U5112 (N_5112,N_1066,N_2093);
nand U5113 (N_5113,N_1204,N_4644);
nand U5114 (N_5114,N_4768,N_208);
nand U5115 (N_5115,N_758,N_3965);
nor U5116 (N_5116,N_1670,N_2784);
or U5117 (N_5117,N_4510,N_2693);
nand U5118 (N_5118,N_2989,N_583);
nor U5119 (N_5119,N_2346,N_4030);
nor U5120 (N_5120,N_75,N_3971);
and U5121 (N_5121,N_4628,N_4553);
nor U5122 (N_5122,N_4616,N_2107);
nand U5123 (N_5123,N_4081,N_2344);
nand U5124 (N_5124,N_3317,N_1717);
nand U5125 (N_5125,N_4484,N_2470);
and U5126 (N_5126,N_1245,N_1977);
nand U5127 (N_5127,N_3719,N_2328);
or U5128 (N_5128,N_921,N_1512);
nor U5129 (N_5129,N_413,N_1949);
and U5130 (N_5130,N_4210,N_1769);
and U5131 (N_5131,N_1875,N_325);
nand U5132 (N_5132,N_803,N_2889);
nor U5133 (N_5133,N_4270,N_614);
nor U5134 (N_5134,N_2151,N_782);
or U5135 (N_5135,N_4019,N_3429);
and U5136 (N_5136,N_4107,N_4097);
and U5137 (N_5137,N_894,N_1052);
or U5138 (N_5138,N_876,N_2322);
nor U5139 (N_5139,N_1632,N_1637);
or U5140 (N_5140,N_1711,N_3488);
nor U5141 (N_5141,N_4969,N_4026);
nand U5142 (N_5142,N_958,N_4021);
and U5143 (N_5143,N_1961,N_1087);
xnor U5144 (N_5144,N_3385,N_2259);
or U5145 (N_5145,N_2141,N_2451);
nor U5146 (N_5146,N_1881,N_4748);
or U5147 (N_5147,N_2922,N_3952);
nor U5148 (N_5148,N_3112,N_1577);
or U5149 (N_5149,N_3738,N_1239);
and U5150 (N_5150,N_527,N_1921);
nor U5151 (N_5151,N_4087,N_1240);
and U5152 (N_5152,N_452,N_1162);
nand U5153 (N_5153,N_1227,N_2617);
or U5154 (N_5154,N_1275,N_1415);
nor U5155 (N_5155,N_1751,N_3110);
nor U5156 (N_5156,N_1925,N_1793);
or U5157 (N_5157,N_1427,N_730);
nor U5158 (N_5158,N_1221,N_97);
nand U5159 (N_5159,N_4387,N_582);
and U5160 (N_5160,N_3309,N_1694);
nand U5161 (N_5161,N_3664,N_1663);
xor U5162 (N_5162,N_2728,N_1967);
and U5163 (N_5163,N_1652,N_2628);
and U5164 (N_5164,N_1269,N_3031);
or U5165 (N_5165,N_2058,N_4074);
or U5166 (N_5166,N_2285,N_2298);
and U5167 (N_5167,N_3292,N_3975);
nor U5168 (N_5168,N_1125,N_2472);
nand U5169 (N_5169,N_3989,N_1898);
and U5170 (N_5170,N_1785,N_3414);
or U5171 (N_5171,N_2103,N_2797);
and U5172 (N_5172,N_1497,N_3996);
nor U5173 (N_5173,N_4206,N_4617);
nand U5174 (N_5174,N_4092,N_857);
nor U5175 (N_5175,N_2717,N_3737);
or U5176 (N_5176,N_2020,N_1303);
or U5177 (N_5177,N_2651,N_2897);
or U5178 (N_5178,N_2425,N_4111);
nand U5179 (N_5179,N_2879,N_296);
nand U5180 (N_5180,N_1309,N_2589);
nand U5181 (N_5181,N_3697,N_1049);
or U5182 (N_5182,N_3713,N_761);
nor U5183 (N_5183,N_432,N_1702);
nor U5184 (N_5184,N_3571,N_1326);
or U5185 (N_5185,N_367,N_1510);
nor U5186 (N_5186,N_146,N_986);
and U5187 (N_5187,N_944,N_1722);
nor U5188 (N_5188,N_3206,N_711);
or U5189 (N_5189,N_265,N_603);
or U5190 (N_5190,N_879,N_1762);
nand U5191 (N_5191,N_4235,N_2815);
nand U5192 (N_5192,N_1438,N_3419);
nand U5193 (N_5193,N_4002,N_143);
nand U5194 (N_5194,N_4636,N_295);
nor U5195 (N_5195,N_350,N_1693);
nand U5196 (N_5196,N_2070,N_4150);
nor U5197 (N_5197,N_3136,N_2663);
nand U5198 (N_5198,N_4905,N_3577);
and U5199 (N_5199,N_4239,N_459);
and U5200 (N_5200,N_131,N_922);
or U5201 (N_5201,N_4065,N_4465);
nor U5202 (N_5202,N_554,N_2975);
nor U5203 (N_5203,N_42,N_1562);
nor U5204 (N_5204,N_2527,N_2251);
nor U5205 (N_5205,N_3567,N_1863);
or U5206 (N_5206,N_3831,N_4756);
or U5207 (N_5207,N_4280,N_4333);
and U5208 (N_5208,N_4418,N_3562);
and U5209 (N_5209,N_3362,N_4241);
nand U5210 (N_5210,N_3217,N_1552);
and U5211 (N_5211,N_3452,N_4363);
nand U5212 (N_5212,N_86,N_4583);
nand U5213 (N_5213,N_2664,N_4603);
or U5214 (N_5214,N_109,N_2398);
and U5215 (N_5215,N_1138,N_1832);
or U5216 (N_5216,N_1404,N_1885);
nor U5217 (N_5217,N_1850,N_1350);
and U5218 (N_5218,N_2809,N_485);
or U5219 (N_5219,N_2767,N_3424);
nor U5220 (N_5220,N_1031,N_2241);
nor U5221 (N_5221,N_2094,N_223);
nand U5222 (N_5222,N_1345,N_4971);
or U5223 (N_5223,N_2340,N_4378);
nor U5224 (N_5224,N_87,N_1292);
nor U5225 (N_5225,N_2330,N_3997);
and U5226 (N_5226,N_1000,N_1947);
or U5227 (N_5227,N_1014,N_46);
nand U5228 (N_5228,N_1942,N_4910);
nor U5229 (N_5229,N_2867,N_2524);
nand U5230 (N_5230,N_3866,N_196);
or U5231 (N_5231,N_472,N_3769);
nand U5232 (N_5232,N_4729,N_4461);
nor U5233 (N_5233,N_3428,N_268);
or U5234 (N_5234,N_3828,N_1758);
or U5235 (N_5235,N_2890,N_3098);
and U5236 (N_5236,N_4004,N_1712);
and U5237 (N_5237,N_4837,N_826);
nor U5238 (N_5238,N_3051,N_2000);
nor U5239 (N_5239,N_4139,N_2500);
or U5240 (N_5240,N_3169,N_2082);
or U5241 (N_5241,N_1598,N_2836);
nand U5242 (N_5242,N_2505,N_4500);
and U5243 (N_5243,N_2703,N_1645);
or U5244 (N_5244,N_1470,N_962);
nand U5245 (N_5245,N_949,N_1092);
and U5246 (N_5246,N_3534,N_3016);
or U5247 (N_5247,N_968,N_1101);
nor U5248 (N_5248,N_3705,N_201);
or U5249 (N_5249,N_3968,N_4089);
or U5250 (N_5250,N_105,N_1644);
or U5251 (N_5251,N_3237,N_2439);
nor U5252 (N_5252,N_1161,N_3793);
and U5253 (N_5253,N_3691,N_4319);
and U5254 (N_5254,N_1914,N_4442);
nand U5255 (N_5255,N_2277,N_2125);
nand U5256 (N_5256,N_4996,N_3330);
nor U5257 (N_5257,N_65,N_4517);
nor U5258 (N_5258,N_2962,N_2980);
or U5259 (N_5259,N_1365,N_58);
or U5260 (N_5260,N_3393,N_1267);
nand U5261 (N_5261,N_1211,N_1951);
or U5262 (N_5262,N_0,N_1894);
or U5263 (N_5263,N_1877,N_992);
and U5264 (N_5264,N_2129,N_4062);
or U5265 (N_5265,N_3326,N_3732);
or U5266 (N_5266,N_794,N_875);
and U5267 (N_5267,N_1990,N_563);
and U5268 (N_5268,N_2598,N_2976);
and U5269 (N_5269,N_1217,N_738);
xor U5270 (N_5270,N_1098,N_187);
and U5271 (N_5271,N_2173,N_3505);
and U5272 (N_5272,N_1647,N_1513);
nand U5273 (N_5273,N_3653,N_61);
or U5274 (N_5274,N_1551,N_3670);
or U5275 (N_5275,N_305,N_1416);
nand U5276 (N_5276,N_1686,N_2168);
nor U5277 (N_5277,N_2228,N_48);
nor U5278 (N_5278,N_1650,N_974);
nand U5279 (N_5279,N_4976,N_602);
xor U5280 (N_5280,N_3467,N_100);
or U5281 (N_5281,N_418,N_1729);
nor U5282 (N_5282,N_167,N_155);
and U5283 (N_5283,N_1447,N_4601);
and U5284 (N_5284,N_3927,N_2163);
and U5285 (N_5285,N_420,N_1165);
and U5286 (N_5286,N_2939,N_3291);
nand U5287 (N_5287,N_3764,N_2011);
nor U5288 (N_5288,N_3778,N_2206);
xnor U5289 (N_5289,N_2378,N_1371);
or U5290 (N_5290,N_1126,N_2088);
and U5291 (N_5291,N_3434,N_2209);
or U5292 (N_5292,N_3377,N_2419);
nor U5293 (N_5293,N_4080,N_4991);
nand U5294 (N_5294,N_3728,N_1063);
or U5295 (N_5295,N_3057,N_4790);
nor U5296 (N_5296,N_2427,N_4650);
nor U5297 (N_5297,N_4665,N_848);
xnor U5298 (N_5298,N_3391,N_1400);
or U5299 (N_5299,N_1593,N_1131);
xnor U5300 (N_5300,N_1665,N_3984);
nand U5301 (N_5301,N_1003,N_3029);
nand U5302 (N_5302,N_2267,N_4811);
and U5303 (N_5303,N_898,N_2543);
or U5304 (N_5304,N_4382,N_866);
or U5305 (N_5305,N_3521,N_4103);
and U5306 (N_5306,N_4001,N_1506);
and U5307 (N_5307,N_3053,N_487);
nor U5308 (N_5308,N_2512,N_4096);
nor U5309 (N_5309,N_3545,N_3671);
and U5310 (N_5310,N_2878,N_3932);
nand U5311 (N_5311,N_342,N_2357);
and U5312 (N_5312,N_3928,N_4470);
nor U5313 (N_5313,N_4779,N_3539);
or U5314 (N_5314,N_3089,N_2002);
nor U5315 (N_5315,N_4178,N_3014);
nand U5316 (N_5316,N_2802,N_207);
xnor U5317 (N_5317,N_3179,N_4475);
nor U5318 (N_5318,N_157,N_525);
nand U5319 (N_5319,N_3912,N_883);
nand U5320 (N_5320,N_2819,N_4788);
or U5321 (N_5321,N_4827,N_2429);
nor U5322 (N_5322,N_3529,N_645);
or U5323 (N_5323,N_3035,N_2682);
and U5324 (N_5324,N_2739,N_1219);
xor U5325 (N_5325,N_2926,N_1305);
nor U5326 (N_5326,N_2952,N_3969);
and U5327 (N_5327,N_3269,N_1730);
or U5328 (N_5328,N_4924,N_1413);
and U5329 (N_5329,N_4507,N_503);
or U5330 (N_5330,N_2216,N_328);
or U5331 (N_5331,N_2407,N_482);
and U5332 (N_5332,N_2128,N_122);
nor U5333 (N_5333,N_3420,N_1796);
xnor U5334 (N_5334,N_1608,N_2462);
nand U5335 (N_5335,N_1869,N_363);
and U5336 (N_5336,N_4389,N_3022);
nor U5337 (N_5337,N_2030,N_3716);
and U5338 (N_5338,N_2687,N_3403);
nor U5339 (N_5339,N_3225,N_4686);
or U5340 (N_5340,N_2409,N_4057);
nor U5341 (N_5341,N_4900,N_1005);
and U5342 (N_5342,N_2669,N_723);
and U5343 (N_5343,N_3967,N_3398);
and U5344 (N_5344,N_4295,N_1818);
or U5345 (N_5345,N_2971,N_1756);
and U5346 (N_5346,N_1073,N_2230);
and U5347 (N_5347,N_4894,N_3357);
and U5348 (N_5348,N_2447,N_2465);
nand U5349 (N_5349,N_222,N_4656);
and U5350 (N_5350,N_4540,N_2231);
and U5351 (N_5351,N_1143,N_756);
or U5352 (N_5352,N_3525,N_2627);
nand U5353 (N_5353,N_4011,N_3131);
or U5354 (N_5354,N_3258,N_3494);
and U5355 (N_5355,N_202,N_3595);
and U5356 (N_5356,N_797,N_3880);
nand U5357 (N_5357,N_4276,N_2014);
or U5358 (N_5358,N_1018,N_3966);
or U5359 (N_5359,N_4256,N_806);
nor U5360 (N_5360,N_3367,N_127);
nand U5361 (N_5361,N_559,N_1278);
nor U5362 (N_5362,N_1798,N_545);
nand U5363 (N_5363,N_3954,N_1822);
and U5364 (N_5364,N_2837,N_951);
nand U5365 (N_5365,N_2672,N_137);
and U5366 (N_5366,N_933,N_1106);
nor U5367 (N_5367,N_1514,N_4414);
xnor U5368 (N_5368,N_1774,N_3617);
nand U5369 (N_5369,N_3686,N_4183);
and U5370 (N_5370,N_1103,N_4320);
and U5371 (N_5371,N_911,N_1554);
and U5372 (N_5372,N_1386,N_1021);
nand U5373 (N_5373,N_4977,N_3129);
or U5374 (N_5374,N_125,N_3644);
nand U5375 (N_5375,N_2306,N_3817);
or U5376 (N_5376,N_1629,N_3819);
nor U5377 (N_5377,N_3701,N_1528);
or U5378 (N_5378,N_38,N_2951);
xor U5379 (N_5379,N_3284,N_192);
or U5380 (N_5380,N_644,N_313);
nand U5381 (N_5381,N_3754,N_547);
nor U5382 (N_5382,N_4660,N_2822);
nor U5383 (N_5383,N_4668,N_4338);
and U5384 (N_5384,N_4834,N_3865);
or U5385 (N_5385,N_4544,N_4791);
or U5386 (N_5386,N_1668,N_2028);
nand U5387 (N_5387,N_501,N_913);
nand U5388 (N_5388,N_32,N_1910);
nand U5389 (N_5389,N_1418,N_4619);
nand U5390 (N_5390,N_340,N_4933);
and U5391 (N_5391,N_926,N_1998);
or U5392 (N_5392,N_3992,N_2558);
or U5393 (N_5393,N_4411,N_3918);
nor U5394 (N_5394,N_3550,N_2586);
and U5395 (N_5395,N_1489,N_4993);
nand U5396 (N_5396,N_4873,N_1993);
and U5397 (N_5397,N_4780,N_1195);
or U5398 (N_5398,N_3840,N_18);
nor U5399 (N_5399,N_128,N_4877);
nand U5400 (N_5400,N_1482,N_1924);
nand U5401 (N_5401,N_4375,N_4516);
and U5402 (N_5402,N_2475,N_834);
nor U5403 (N_5403,N_1812,N_22);
nand U5404 (N_5404,N_3765,N_3800);
nor U5405 (N_5405,N_4867,N_461);
or U5406 (N_5406,N_2245,N_2790);
and U5407 (N_5407,N_2203,N_421);
and U5408 (N_5408,N_3849,N_1842);
xnor U5409 (N_5409,N_2489,N_136);
nand U5410 (N_5410,N_3387,N_4523);
and U5411 (N_5411,N_4505,N_2426);
nand U5412 (N_5412,N_388,N_236);
nor U5413 (N_5413,N_3,N_788);
and U5414 (N_5414,N_759,N_1128);
nand U5415 (N_5415,N_3805,N_914);
nor U5416 (N_5416,N_2670,N_2326);
and U5417 (N_5417,N_333,N_2616);
nand U5418 (N_5418,N_4661,N_2263);
nor U5419 (N_5419,N_1307,N_3776);
or U5420 (N_5420,N_1630,N_2354);
nor U5421 (N_5421,N_2096,N_1873);
nor U5422 (N_5422,N_1892,N_1680);
nor U5423 (N_5423,N_70,N_2813);
or U5424 (N_5424,N_181,N_3739);
and U5425 (N_5425,N_1886,N_3830);
or U5426 (N_5426,N_2458,N_2424);
or U5427 (N_5427,N_3478,N_1273);
or U5428 (N_5428,N_1755,N_4416);
or U5429 (N_5429,N_2801,N_209);
nor U5430 (N_5430,N_1611,N_1596);
nand U5431 (N_5431,N_2395,N_2700);
nor U5432 (N_5432,N_4671,N_271);
nand U5433 (N_5433,N_1794,N_2713);
nor U5434 (N_5434,N_3353,N_3599);
nand U5435 (N_5435,N_2864,N_4369);
and U5436 (N_5436,N_2550,N_1580);
or U5437 (N_5437,N_3685,N_4824);
or U5438 (N_5438,N_386,N_4497);
nor U5439 (N_5439,N_2831,N_248);
nor U5440 (N_5440,N_855,N_3196);
nand U5441 (N_5441,N_2707,N_4807);
xnor U5442 (N_5442,N_1265,N_657);
and U5443 (N_5443,N_117,N_4953);
nand U5444 (N_5444,N_2861,N_4219);
nor U5445 (N_5445,N_4849,N_2781);
or U5446 (N_5446,N_1594,N_4865);
xor U5447 (N_5447,N_3889,N_4306);
nor U5448 (N_5448,N_4897,N_2587);
or U5449 (N_5449,N_1393,N_4005);
nor U5450 (N_5450,N_2862,N_4052);
nor U5451 (N_5451,N_627,N_2174);
nor U5452 (N_5452,N_4196,N_3695);
xor U5453 (N_5453,N_410,N_1656);
or U5454 (N_5454,N_624,N_495);
nor U5455 (N_5455,N_2810,N_1889);
nand U5456 (N_5456,N_3829,N_252);
nor U5457 (N_5457,N_3389,N_4980);
nor U5458 (N_5458,N_2051,N_2721);
nand U5459 (N_5459,N_1041,N_3036);
or U5460 (N_5460,N_2396,N_2715);
and U5461 (N_5461,N_453,N_1801);
and U5462 (N_5462,N_4250,N_1811);
or U5463 (N_5463,N_2363,N_1212);
nor U5464 (N_5464,N_2909,N_4793);
or U5465 (N_5465,N_3510,N_2032);
nor U5466 (N_5466,N_2624,N_3808);
nor U5467 (N_5467,N_3263,N_3751);
nand U5468 (N_5468,N_668,N_601);
nand U5469 (N_5469,N_3709,N_4329);
nand U5470 (N_5470,N_767,N_2215);
nand U5471 (N_5471,N_1097,N_2657);
or U5472 (N_5472,N_2441,N_3540);
or U5473 (N_5473,N_3816,N_2648);
nor U5474 (N_5474,N_3652,N_76);
or U5475 (N_5475,N_2742,N_2261);
nand U5476 (N_5476,N_2588,N_4137);
or U5477 (N_5477,N_3706,N_1370);
nor U5478 (N_5478,N_2918,N_2748);
xor U5479 (N_5479,N_4741,N_889);
nor U5480 (N_5480,N_2957,N_3852);
or U5481 (N_5481,N_725,N_4243);
nand U5482 (N_5482,N_3844,N_1727);
nor U5483 (N_5483,N_860,N_1406);
nand U5484 (N_5484,N_3444,N_4215);
or U5485 (N_5485,N_1684,N_3548);
or U5486 (N_5486,N_2001,N_1456);
nand U5487 (N_5487,N_139,N_4548);
nand U5488 (N_5488,N_1464,N_3841);
and U5489 (N_5489,N_912,N_4022);
or U5490 (N_5490,N_4623,N_4832);
and U5491 (N_5491,N_4045,N_1649);
or U5492 (N_5492,N_3366,N_2908);
or U5493 (N_5493,N_3188,N_4967);
nand U5494 (N_5494,N_3980,N_2750);
or U5495 (N_5495,N_3970,N_4621);
nor U5496 (N_5496,N_1657,N_4133);
nand U5497 (N_5497,N_4703,N_4447);
nor U5498 (N_5498,N_1688,N_688);
and U5499 (N_5499,N_2579,N_4645);
nand U5500 (N_5500,N_3724,N_2863);
nor U5501 (N_5501,N_116,N_3915);
nand U5502 (N_5502,N_2949,N_3504);
or U5503 (N_5503,N_1991,N_572);
and U5504 (N_5504,N_564,N_1347);
nand U5505 (N_5505,N_3375,N_2888);
and U5506 (N_5506,N_2756,N_1207);
or U5507 (N_5507,N_339,N_3007);
nor U5508 (N_5508,N_4132,N_4909);
nor U5509 (N_5509,N_15,N_4020);
nand U5510 (N_5510,N_1311,N_1495);
and U5511 (N_5511,N_203,N_4639);
or U5512 (N_5512,N_3455,N_2319);
nand U5513 (N_5513,N_4261,N_1184);
nand U5514 (N_5514,N_3437,N_4543);
or U5515 (N_5515,N_2385,N_997);
nand U5516 (N_5516,N_854,N_2540);
or U5517 (N_5517,N_244,N_2611);
nand U5518 (N_5518,N_1412,N_808);
nand U5519 (N_5519,N_2502,N_290);
and U5520 (N_5520,N_2643,N_1074);
and U5521 (N_5521,N_2887,N_475);
or U5522 (N_5522,N_352,N_2175);
or U5523 (N_5523,N_138,N_2358);
or U5524 (N_5524,N_4951,N_3516);
and U5525 (N_5525,N_2234,N_1527);
nor U5526 (N_5526,N_3544,N_3138);
or U5527 (N_5527,N_2600,N_4036);
nor U5528 (N_5528,N_4386,N_1270);
nand U5529 (N_5529,N_4407,N_3116);
nand U5530 (N_5530,N_2379,N_1159);
nor U5531 (N_5531,N_4293,N_2959);
nor U5532 (N_5532,N_190,N_3948);
nand U5533 (N_5533,N_3018,N_2921);
nand U5534 (N_5534,N_344,N_3365);
nor U5535 (N_5535,N_4579,N_2401);
nand U5536 (N_5536,N_489,N_3784);
nand U5537 (N_5537,N_4232,N_998);
and U5538 (N_5538,N_612,N_3827);
xnor U5539 (N_5539,N_2432,N_2392);
and U5540 (N_5540,N_3983,N_2953);
or U5541 (N_5541,N_924,N_710);
and U5542 (N_5542,N_1648,N_4207);
nand U5543 (N_5543,N_3072,N_755);
or U5544 (N_5544,N_4949,N_4229);
or U5545 (N_5545,N_2254,N_2383);
nor U5546 (N_5546,N_2060,N_4275);
or U5547 (N_5547,N_434,N_3068);
nor U5548 (N_5548,N_3340,N_4184);
and U5549 (N_5549,N_4554,N_689);
and U5550 (N_5550,N_3472,N_3950);
or U5551 (N_5551,N_3320,N_3355);
or U5552 (N_5552,N_2433,N_3720);
or U5553 (N_5553,N_1011,N_3541);
nand U5554 (N_5554,N_391,N_1653);
nor U5555 (N_5555,N_4752,N_1449);
and U5556 (N_5556,N_548,N_1054);
and U5557 (N_5557,N_1932,N_4773);
and U5558 (N_5558,N_825,N_2450);
nor U5559 (N_5559,N_835,N_780);
and U5560 (N_5560,N_1973,N_4010);
nand U5561 (N_5561,N_286,N_4545);
or U5562 (N_5562,N_3107,N_1276);
or U5563 (N_5563,N_4160,N_1254);
nor U5564 (N_5564,N_148,N_3448);
xnor U5565 (N_5565,N_121,N_3371);
nor U5566 (N_5566,N_3886,N_4538);
nor U5567 (N_5567,N_2481,N_4866);
and U5568 (N_5568,N_4921,N_4079);
nand U5569 (N_5569,N_2325,N_2800);
and U5570 (N_5570,N_1086,N_920);
nand U5571 (N_5571,N_2662,N_94);
nor U5572 (N_5572,N_3923,N_1809);
nand U5573 (N_5573,N_4913,N_3369);
and U5574 (N_5574,N_3458,N_2402);
and U5575 (N_5575,N_524,N_245);
or U5576 (N_5576,N_1341,N_1566);
nor U5577 (N_5577,N_3958,N_4076);
and U5578 (N_5578,N_4959,N_474);
or U5579 (N_5579,N_71,N_273);
nor U5580 (N_5580,N_4428,N_3105);
nor U5581 (N_5581,N_1968,N_3603);
and U5582 (N_5582,N_721,N_40);
nand U5583 (N_5583,N_1164,N_1529);
or U5584 (N_5584,N_732,N_3526);
and U5585 (N_5585,N_1752,N_3461);
and U5586 (N_5586,N_3580,N_3693);
and U5587 (N_5587,N_2296,N_335);
nor U5588 (N_5588,N_1900,N_3694);
or U5589 (N_5589,N_2114,N_1639);
and U5590 (N_5590,N_2595,N_2795);
and U5591 (N_5591,N_3204,N_1078);
nand U5592 (N_5592,N_3314,N_625);
nand U5593 (N_5593,N_2603,N_172);
nor U5594 (N_5594,N_2178,N_1601);
or U5595 (N_5595,N_1825,N_182);
and U5596 (N_5596,N_3628,N_4049);
or U5597 (N_5597,N_5,N_4754);
nor U5598 (N_5598,N_447,N_4736);
xnor U5599 (N_5599,N_2725,N_4986);
nand U5600 (N_5600,N_355,N_1251);
and U5601 (N_5601,N_1996,N_4972);
and U5602 (N_5602,N_3207,N_3408);
nand U5603 (N_5603,N_3262,N_1671);
or U5604 (N_5604,N_1606,N_1038);
and U5605 (N_5605,N_3988,N_1249);
or U5606 (N_5606,N_4217,N_4377);
nand U5607 (N_5607,N_4869,N_322);
nand U5608 (N_5608,N_1330,N_973);
nor U5609 (N_5609,N_589,N_963);
and U5610 (N_5610,N_4189,N_2180);
nor U5611 (N_5611,N_1380,N_358);
nor U5612 (N_5612,N_1897,N_1481);
xnor U5613 (N_5613,N_830,N_1109);
nor U5614 (N_5614,N_1548,N_2381);
and U5615 (N_5615,N_51,N_1290);
or U5616 (N_5616,N_839,N_372);
nand U5617 (N_5617,N_1337,N_3184);
and U5618 (N_5618,N_4804,N_145);
and U5619 (N_5619,N_4842,N_2714);
nor U5620 (N_5620,N_4156,N_2964);
and U5621 (N_5621,N_356,N_1966);
nand U5622 (N_5622,N_1995,N_4388);
nand U5623 (N_5623,N_4481,N_846);
nand U5624 (N_5624,N_3904,N_2720);
and U5625 (N_5625,N_4187,N_2824);
and U5626 (N_5626,N_2753,N_2347);
and U5627 (N_5627,N_648,N_1051);
and U5628 (N_5628,N_762,N_3982);
nand U5629 (N_5629,N_3596,N_2494);
and U5630 (N_5630,N_3822,N_3399);
and U5631 (N_5631,N_731,N_3358);
or U5632 (N_5632,N_2641,N_2256);
nand U5633 (N_5633,N_1659,N_2655);
or U5634 (N_5634,N_1655,N_1252);
nand U5635 (N_5635,N_2906,N_2596);
or U5636 (N_5636,N_4974,N_1716);
nor U5637 (N_5637,N_406,N_2899);
nor U5638 (N_5638,N_1059,N_2724);
or U5639 (N_5639,N_1300,N_807);
nor U5640 (N_5640,N_2264,N_694);
nand U5641 (N_5641,N_3673,N_2877);
and U5642 (N_5642,N_1302,N_28);
xnor U5643 (N_5643,N_2299,N_2061);
nor U5644 (N_5644,N_2710,N_1797);
or U5645 (N_5645,N_197,N_3884);
nand U5646 (N_5646,N_2062,N_1732);
and U5647 (N_5647,N_3078,N_4696);
or U5648 (N_5648,N_39,N_3205);
nand U5649 (N_5649,N_4536,N_642);
nand U5650 (N_5650,N_2403,N_3807);
nor U5651 (N_5651,N_3468,N_4770);
and U5652 (N_5652,N_3240,N_4798);
or U5653 (N_5653,N_3231,N_174);
and U5654 (N_5654,N_4374,N_2712);
nor U5655 (N_5655,N_4954,N_1286);
and U5656 (N_5656,N_2198,N_4075);
or U5657 (N_5657,N_4456,N_2804);
nor U5658 (N_5658,N_1363,N_4647);
nor U5659 (N_5659,N_2799,N_3283);
nor U5660 (N_5660,N_2138,N_2923);
nand U5661 (N_5661,N_397,N_60);
nor U5662 (N_5662,N_1916,N_2079);
or U5663 (N_5663,N_4888,N_4573);
or U5664 (N_5664,N_4450,N_1430);
xnor U5665 (N_5665,N_1646,N_740);
nand U5666 (N_5666,N_3171,N_1641);
nor U5667 (N_5667,N_4956,N_1333);
nand U5668 (N_5668,N_3278,N_1190);
nor U5669 (N_5669,N_2690,N_1520);
nand U5670 (N_5670,N_3048,N_4483);
nor U5671 (N_5671,N_2118,N_4528);
nor U5672 (N_5672,N_2993,N_2202);
nor U5673 (N_5673,N_2526,N_1354);
and U5674 (N_5674,N_3842,N_4216);
or U5675 (N_5675,N_2482,N_3288);
nor U5676 (N_5676,N_4466,N_3492);
nor U5677 (N_5677,N_4044,N_1642);
nor U5678 (N_5678,N_3380,N_1127);
or U5679 (N_5679,N_838,N_733);
nor U5680 (N_5680,N_633,N_1872);
or U5681 (N_5681,N_3017,N_1385);
nor U5682 (N_5682,N_2930,N_2916);
xnor U5683 (N_5683,N_2099,N_1009);
or U5684 (N_5684,N_2842,N_458);
or U5685 (N_5685,N_1234,N_813);
nor U5686 (N_5686,N_2005,N_1075);
and U5687 (N_5687,N_1202,N_184);
nand U5688 (N_5688,N_2006,N_2268);
nand U5689 (N_5689,N_2384,N_3094);
xnor U5690 (N_5690,N_4240,N_1258);
and U5691 (N_5691,N_3061,N_2634);
nor U5692 (N_5692,N_1056,N_4708);
nor U5693 (N_5693,N_3749,N_1395);
nand U5694 (N_5694,N_1335,N_4162);
xnor U5695 (N_5695,N_2187,N_956);
and U5696 (N_5696,N_4874,N_4907);
nor U5697 (N_5697,N_683,N_3307);
and U5698 (N_5698,N_3476,N_311);
and U5699 (N_5699,N_3919,N_1467);
nand U5700 (N_5700,N_304,N_1083);
nand U5701 (N_5701,N_4698,N_2132);
or U5702 (N_5702,N_4158,N_4841);
nand U5703 (N_5703,N_4723,N_2876);
nand U5704 (N_5704,N_4539,N_3905);
and U5705 (N_5705,N_4220,N_1356);
and U5706 (N_5706,N_4291,N_2848);
or U5707 (N_5707,N_2566,N_3080);
nor U5708 (N_5708,N_4135,N_2659);
and U5709 (N_5709,N_2314,N_2779);
xor U5710 (N_5710,N_4476,N_3334);
nor U5711 (N_5711,N_1700,N_4796);
and U5712 (N_5712,N_3938,N_3900);
nor U5713 (N_5713,N_718,N_1901);
nor U5714 (N_5714,N_2694,N_1620);
and U5715 (N_5715,N_3632,N_2740);
and U5716 (N_5716,N_1559,N_1112);
nor U5717 (N_5717,N_1203,N_2150);
nand U5718 (N_5718,N_1747,N_166);
and U5719 (N_5719,N_4179,N_887);
nand U5720 (N_5720,N_1166,N_1713);
or U5721 (N_5721,N_206,N_3024);
nand U5722 (N_5722,N_4014,N_2758);
nand U5723 (N_5723,N_282,N_2629);
nor U5724 (N_5724,N_1591,N_2985);
nor U5725 (N_5725,N_1868,N_660);
and U5726 (N_5726,N_1695,N_383);
nor U5727 (N_5727,N_537,N_151);
and U5728 (N_5728,N_4559,N_1409);
nor U5729 (N_5729,N_3441,N_4054);
nand U5730 (N_5730,N_4161,N_934);
and U5731 (N_5731,N_549,N_3255);
or U5732 (N_5732,N_1315,N_4350);
and U5733 (N_5733,N_1462,N_4787);
and U5734 (N_5734,N_4881,N_2119);
nand U5735 (N_5735,N_3037,N_2161);
or U5736 (N_5736,N_3412,N_1878);
nand U5737 (N_5737,N_3902,N_4072);
xor U5738 (N_5738,N_4522,N_4941);
or U5739 (N_5739,N_2722,N_1253);
or U5740 (N_5740,N_4813,N_274);
nand U5741 (N_5741,N_1153,N_1664);
nand U5742 (N_5742,N_257,N_3019);
and U5743 (N_5743,N_338,N_3100);
nand U5744 (N_5744,N_637,N_1346);
nand U5745 (N_5745,N_4511,N_4298);
xor U5746 (N_5746,N_2597,N_3004);
and U5747 (N_5747,N_4765,N_3056);
nand U5748 (N_5748,N_130,N_1959);
or U5749 (N_5749,N_4604,N_249);
nor U5750 (N_5750,N_1571,N_853);
xnor U5751 (N_5751,N_3987,N_3000);
and U5752 (N_5752,N_4989,N_3524);
and U5753 (N_5753,N_1802,N_3273);
nor U5754 (N_5754,N_3250,N_1690);
nand U5755 (N_5755,N_2468,N_4932);
or U5756 (N_5756,N_1414,N_4237);
xnor U5757 (N_5757,N_817,N_3427);
nand U5758 (N_5758,N_4109,N_2488);
and U5759 (N_5759,N_3985,N_622);
nand U5760 (N_5760,N_4519,N_950);
and U5761 (N_5761,N_2148,N_1569);
nor U5762 (N_5762,N_4060,N_815);
nor U5763 (N_5763,N_1935,N_396);
or U5764 (N_5764,N_859,N_34);
or U5765 (N_5765,N_1895,N_4425);
and U5766 (N_5766,N_4868,N_477);
nand U5767 (N_5767,N_1151,N_3409);
nand U5768 (N_5768,N_3033,N_3814);
or U5769 (N_5769,N_4146,N_2691);
nand U5770 (N_5770,N_4513,N_2223);
nand U5771 (N_5771,N_2501,N_3579);
or U5772 (N_5772,N_492,N_460);
nand U5773 (N_5773,N_3088,N_4532);
nand U5774 (N_5774,N_1880,N_2626);
nand U5775 (N_5775,N_4264,N_4890);
nor U5776 (N_5776,N_2201,N_1281);
nand U5777 (N_5777,N_715,N_3046);
and U5778 (N_5778,N_4922,N_4624);
and U5779 (N_5779,N_177,N_626);
or U5780 (N_5780,N_3118,N_3949);
or U5781 (N_5781,N_4208,N_2290);
and U5782 (N_5782,N_3010,N_2549);
or U5783 (N_5783,N_1844,N_1904);
nand U5784 (N_5784,N_3466,N_4730);
nand U5785 (N_5785,N_4701,N_4071);
and U5786 (N_5786,N_3069,N_4962);
nand U5787 (N_5787,N_2443,N_430);
nand U5788 (N_5788,N_3345,N_2510);
and U5789 (N_5789,N_334,N_4417);
xor U5790 (N_5790,N_3287,N_4040);
or U5791 (N_5791,N_360,N_4123);
nand U5792 (N_5792,N_2190,N_3477);
nor U5793 (N_5793,N_1428,N_3921);
and U5794 (N_5794,N_4223,N_1186);
or U5795 (N_5795,N_1397,N_2406);
nand U5796 (N_5796,N_3058,N_2377);
nand U5797 (N_5797,N_3203,N_1149);
nand U5798 (N_5798,N_4794,N_4880);
or U5799 (N_5799,N_126,N_4833);
nand U5800 (N_5800,N_468,N_1222);
or U5801 (N_5801,N_2492,N_1490);
or U5802 (N_5802,N_2239,N_2568);
nor U5803 (N_5803,N_3117,N_4127);
nand U5804 (N_5804,N_392,N_13);
nand U5805 (N_5805,N_2827,N_3654);
nand U5806 (N_5806,N_3130,N_4202);
or U5807 (N_5807,N_3574,N_176);
or U5808 (N_5808,N_1833,N_2695);
nand U5809 (N_5809,N_3337,N_878);
and U5810 (N_5810,N_972,N_1084);
nor U5811 (N_5811,N_4488,N_4911);
and U5812 (N_5812,N_3502,N_2591);
nand U5813 (N_5813,N_3396,N_66);
nand U5814 (N_5814,N_4682,N_435);
nor U5815 (N_5815,N_1613,N_2025);
nand U5816 (N_5816,N_777,N_3319);
nand U5817 (N_5817,N_2613,N_2027);
or U5818 (N_5818,N_162,N_2262);
nand U5819 (N_5819,N_1864,N_3556);
nor U5820 (N_5820,N_3658,N_3422);
nand U5821 (N_5821,N_574,N_2736);
or U5822 (N_5822,N_4785,N_3300);
and U5823 (N_5823,N_2575,N_552);
or U5824 (N_5824,N_2113,N_3888);
nand U5825 (N_5825,N_3293,N_1588);
nand U5826 (N_5826,N_3692,N_4225);
or U5827 (N_5827,N_1823,N_3001);
or U5828 (N_5828,N_4213,N_2927);
nand U5829 (N_5829,N_4937,N_3916);
or U5830 (N_5830,N_3532,N_4713);
or U5831 (N_5831,N_2493,N_1492);
and U5832 (N_5832,N_481,N_844);
and U5833 (N_5833,N_2885,N_1381);
or U5834 (N_5834,N_3045,N_1536);
nor U5835 (N_5835,N_3085,N_1791);
xor U5836 (N_5836,N_2580,N_996);
nor U5837 (N_5837,N_1518,N_2440);
nor U5838 (N_5838,N_2734,N_4337);
and U5839 (N_5839,N_2632,N_3779);
and U5840 (N_5840,N_2646,N_3503);
and U5841 (N_5841,N_2009,N_3210);
nand U5842 (N_5842,N_3123,N_793);
and U5843 (N_5843,N_2761,N_2188);
or U5844 (N_5844,N_1013,N_3922);
or U5845 (N_5845,N_577,N_4214);
nor U5846 (N_5846,N_2825,N_1499);
nor U5847 (N_5847,N_2031,N_1237);
and U5848 (N_5848,N_1174,N_3049);
and U5849 (N_5849,N_4003,N_1679);
nand U5850 (N_5850,N_3006,N_25);
nand U5851 (N_5851,N_4688,N_3460);
nand U5852 (N_5852,N_3490,N_1635);
nor U5853 (N_5853,N_3224,N_4838);
nor U5854 (N_5854,N_1705,N_3986);
nor U5855 (N_5855,N_3976,N_3122);
and U5856 (N_5856,N_150,N_2366);
or U5857 (N_5857,N_1905,N_1173);
or U5858 (N_5858,N_1734,N_3473);
or U5859 (N_5859,N_1067,N_2302);
or U5860 (N_5860,N_101,N_4720);
or U5861 (N_5861,N_575,N_1457);
or U5862 (N_5862,N_1491,N_102);
nand U5863 (N_5863,N_3843,N_677);
nand U5864 (N_5864,N_2601,N_4406);
and U5865 (N_5865,N_4260,N_1077);
nand U5866 (N_5866,N_1458,N_1072);
and U5867 (N_5867,N_2798,N_4473);
nand U5868 (N_5868,N_3639,N_2087);
nand U5869 (N_5869,N_615,N_708);
xnor U5870 (N_5870,N_3267,N_2677);
and U5871 (N_5871,N_2321,N_2533);
or U5872 (N_5872,N_4917,N_4000);
and U5873 (N_5873,N_2017,N_3648);
and U5874 (N_5874,N_4709,N_470);
and U5875 (N_5875,N_3305,N_3413);
and U5876 (N_5876,N_2146,N_1736);
nor U5877 (N_5877,N_3517,N_3791);
and U5878 (N_5878,N_1612,N_4342);
nor U5879 (N_5879,N_3407,N_510);
or U5880 (N_5880,N_2614,N_3030);
or U5881 (N_5881,N_353,N_2992);
and U5882 (N_5882,N_4884,N_673);
and U5883 (N_5883,N_3785,N_4600);
nor U5884 (N_5884,N_2362,N_3480);
xnor U5885 (N_5885,N_3047,N_2179);
nand U5886 (N_5886,N_3853,N_4460);
or U5887 (N_5887,N_1030,N_1343);
nor U5888 (N_5888,N_4863,N_2509);
and U5889 (N_5889,N_2189,N_77);
nor U5890 (N_5890,N_2442,N_2394);
nor U5891 (N_5891,N_509,N_3190);
and U5892 (N_5892,N_923,N_4370);
or U5893 (N_5893,N_1997,N_107);
nor U5894 (N_5894,N_3846,N_1429);
nand U5895 (N_5895,N_2970,N_1619);
nand U5896 (N_5896,N_4181,N_985);
nor U5897 (N_5897,N_1008,N_2766);
nand U5898 (N_5898,N_3930,N_35);
nor U5899 (N_5899,N_4535,N_436);
nor U5900 (N_5900,N_3297,N_1855);
nand U5901 (N_5901,N_82,N_4464);
and U5902 (N_5902,N_630,N_4082);
or U5903 (N_5903,N_3003,N_3227);
nor U5904 (N_5904,N_3332,N_4607);
and U5905 (N_5905,N_2244,N_2159);
or U5906 (N_5906,N_2893,N_1669);
nand U5907 (N_5907,N_4626,N_584);
or U5908 (N_5908,N_4498,N_4171);
xor U5909 (N_5909,N_540,N_2701);
nor U5910 (N_5910,N_2108,N_4722);
nand U5911 (N_5911,N_3180,N_493);
or U5912 (N_5912,N_4706,N_2222);
nor U5913 (N_5913,N_306,N_1917);
or U5914 (N_5914,N_2506,N_1972);
nand U5915 (N_5915,N_4066,N_1541);
or U5916 (N_5916,N_2803,N_1544);
xnor U5917 (N_5917,N_1944,N_2907);
nand U5918 (N_5918,N_3847,N_1129);
and U5919 (N_5919,N_831,N_606);
nor U5920 (N_5920,N_4455,N_31);
nor U5921 (N_5921,N_654,N_3257);
nand U5922 (N_5922,N_804,N_1865);
or U5923 (N_5923,N_2935,N_3678);
nand U5924 (N_5924,N_899,N_4151);
and U5925 (N_5925,N_132,N_3302);
nor U5926 (N_5926,N_3708,N_1255);
nor U5927 (N_5927,N_4851,N_3182);
xnor U5928 (N_5928,N_653,N_2295);
nand U5929 (N_5929,N_414,N_3848);
and U5930 (N_5930,N_959,N_1368);
nand U5931 (N_5931,N_2995,N_4557);
or U5932 (N_5932,N_1241,N_2078);
nor U5933 (N_5933,N_3638,N_2941);
nand U5934 (N_5934,N_801,N_220);
and U5935 (N_5935,N_930,N_2207);
and U5936 (N_5936,N_2843,N_4515);
xor U5937 (N_5937,N_111,N_2945);
nand U5938 (N_5938,N_2253,N_4166);
and U5939 (N_5939,N_4159,N_3998);
or U5940 (N_5940,N_4929,N_1137);
nand U5941 (N_5941,N_4226,N_1890);
or U5942 (N_5942,N_365,N_427);
nor U5943 (N_5943,N_3826,N_3547);
nand U5944 (N_5944,N_773,N_4286);
and U5945 (N_5945,N_2227,N_1826);
xnor U5946 (N_5946,N_3132,N_1858);
and U5947 (N_5947,N_403,N_2355);
nand U5948 (N_5948,N_1625,N_408);
or U5949 (N_5949,N_3882,N_4936);
nor U5950 (N_5950,N_24,N_2965);
nor U5951 (N_5951,N_3096,N_2590);
and U5952 (N_5952,N_3659,N_2186);
and U5953 (N_5953,N_4862,N_1662);
nor U5954 (N_5954,N_4028,N_2248);
nand U5955 (N_5955,N_4767,N_1339);
nand U5956 (N_5956,N_4281,N_2553);
nor U5957 (N_5957,N_2459,N_4318);
or U5958 (N_5958,N_4871,N_2678);
or U5959 (N_5959,N_2497,N_1431);
nand U5960 (N_5960,N_4852,N_669);
nand U5961 (N_5961,N_1856,N_53);
nand U5962 (N_5962,N_2853,N_4249);
and U5963 (N_5963,N_1638,N_4902);
or U5964 (N_5964,N_1383,N_1879);
xnor U5965 (N_5965,N_2745,N_1731);
or U5966 (N_5966,N_450,N_3496);
nand U5967 (N_5967,N_345,N_1313);
and U5968 (N_5968,N_3032,N_702);
or U5969 (N_5969,N_4200,N_3282);
nor U5970 (N_5970,N_4551,N_3592);
nor U5971 (N_5971,N_2055,N_4362);
nand U5972 (N_5972,N_2780,N_44);
nand U5973 (N_5973,N_3995,N_2183);
nand U5974 (N_5974,N_2541,N_2133);
and U5975 (N_5975,N_445,N_212);
nand U5976 (N_5976,N_2544,N_3799);
or U5977 (N_5977,N_229,N_1743);
nor U5978 (N_5978,N_2086,N_2844);
nand U5979 (N_5979,N_11,N_4255);
nor U5980 (N_5980,N_1338,N_2130);
nand U5981 (N_5981,N_4808,N_553);
nand U5982 (N_5982,N_193,N_3947);
and U5983 (N_5983,N_281,N_3469);
nand U5984 (N_5984,N_4572,N_3009);
and U5985 (N_5985,N_3200,N_3564);
or U5986 (N_5986,N_4346,N_2882);
or U5987 (N_5987,N_4422,N_4029);
and U5988 (N_5988,N_409,N_3689);
nand U5989 (N_5989,N_2320,N_1266);
nor U5990 (N_5990,N_2771,N_3650);
nor U5991 (N_5991,N_4059,N_2986);
or U5992 (N_5992,N_1163,N_1461);
or U5993 (N_5993,N_2361,N_3343);
or U5994 (N_5994,N_496,N_3471);
nand U5995 (N_5995,N_965,N_3405);
and U5996 (N_5996,N_4614,N_3956);
or U5997 (N_5997,N_3431,N_849);
and U5998 (N_5998,N_2743,N_4294);
nand U5999 (N_5999,N_511,N_2785);
xnor U6000 (N_6000,N_2666,N_4733);
nor U6001 (N_6001,N_4876,N_987);
nor U6002 (N_6002,N_213,N_3114);
nor U6003 (N_6003,N_2674,N_3454);
nand U6004 (N_6004,N_30,N_1410);
nand U6005 (N_6005,N_4957,N_3167);
or U6006 (N_6006,N_752,N_4008);
nor U6007 (N_6007,N_1813,N_1035);
or U6008 (N_6008,N_3197,N_1685);
and U6009 (N_6009,N_608,N_636);
or U6010 (N_6010,N_113,N_802);
and U6011 (N_6011,N_2485,N_417);
and U6012 (N_6012,N_983,N_3159);
nand U6013 (N_6013,N_2751,N_1770);
or U6014 (N_6014,N_967,N_3083);
or U6015 (N_6015,N_4222,N_1615);
and U6016 (N_6016,N_576,N_955);
nand U6017 (N_6017,N_4950,N_2987);
or U6018 (N_6018,N_1965,N_1325);
nand U6019 (N_6019,N_2371,N_1719);
and U6020 (N_6020,N_1036,N_1274);
and U6021 (N_6021,N_910,N_118);
nand U6022 (N_6022,N_3868,N_393);
and U6023 (N_6023,N_1815,N_4858);
or U6024 (N_6024,N_787,N_3721);
or U6025 (N_6025,N_1771,N_526);
nand U6026 (N_6026,N_1987,N_1348);
nor U6027 (N_6027,N_2683,N_519);
nand U6028 (N_6028,N_4509,N_3296);
nor U6029 (N_6029,N_20,N_2349);
nand U6030 (N_6030,N_918,N_2122);
nand U6031 (N_6031,N_3501,N_3402);
nand U6032 (N_6032,N_2528,N_4782);
and U6033 (N_6033,N_2778,N_1188);
and U6034 (N_6034,N_2919,N_1970);
or U6035 (N_6035,N_1352,N_1957);
nand U6036 (N_6036,N_3602,N_1440);
nand U6037 (N_6037,N_2368,N_2071);
nand U6038 (N_6038,N_4155,N_4925);
or U6039 (N_6039,N_1840,N_1586);
nor U6040 (N_6040,N_3775,N_1257);
nand U6041 (N_6041,N_2247,N_2194);
nor U6042 (N_6042,N_2102,N_1539);
and U6043 (N_6043,N_1517,N_1599);
or U6044 (N_6044,N_3696,N_1903);
nor U6045 (N_6045,N_3523,N_1279);
and U6046 (N_6046,N_686,N_3860);
and U6047 (N_6047,N_765,N_4170);
nor U6048 (N_6048,N_267,N_4412);
and U6049 (N_6049,N_390,N_635);
or U6050 (N_6050,N_2609,N_4697);
and U6051 (N_6051,N_3991,N_4799);
nand U6052 (N_6052,N_2034,N_1029);
nand U6053 (N_6053,N_2417,N_1057);
or U6054 (N_6054,N_4423,N_515);
or U6055 (N_6055,N_1191,N_837);
and U6056 (N_6056,N_324,N_2335);
and U6057 (N_6057,N_3363,N_2147);
nor U6058 (N_6058,N_3272,N_1349);
nor U6059 (N_6059,N_4038,N_2914);
or U6060 (N_6060,N_1676,N_895);
or U6061 (N_6061,N_4157,N_1764);
or U6062 (N_6062,N_2960,N_3674);
nor U6063 (N_6063,N_3862,N_4197);
xor U6064 (N_6064,N_4348,N_2806);
or U6065 (N_6065,N_3443,N_4587);
or U6066 (N_6066,N_800,N_4091);
or U6067 (N_6067,N_2003,N_3643);
and U6068 (N_6068,N_4313,N_581);
nor U6069 (N_6069,N_389,N_3700);
nand U6070 (N_6070,N_2438,N_2343);
xor U6071 (N_6071,N_2224,N_1933);
nand U6072 (N_6072,N_969,N_4047);
nand U6073 (N_6073,N_228,N_4489);
nand U6074 (N_6074,N_1389,N_4727);
or U6075 (N_6075,N_2044,N_3060);
nand U6076 (N_6076,N_4719,N_2966);
nand U6077 (N_6077,N_1714,N_2582);
or U6078 (N_6078,N_1377,N_2436);
nor U6079 (N_6079,N_1535,N_4674);
or U6080 (N_6080,N_1250,N_640);
and U6081 (N_6081,N_443,N_2171);
or U6082 (N_6082,N_3647,N_2158);
nand U6083 (N_6083,N_4629,N_1198);
and U6084 (N_6084,N_1322,N_2917);
nand U6085 (N_6085,N_3416,N_337);
nor U6086 (N_6086,N_1361,N_437);
or U6087 (N_6087,N_2638,N_4547);
or U6088 (N_6088,N_4441,N_3276);
nor U6089 (N_6089,N_1310,N_1994);
nand U6090 (N_6090,N_2947,N_971);
nand U6091 (N_6091,N_4041,N_799);
nand U6092 (N_6092,N_4268,N_2237);
nor U6093 (N_6093,N_4744,N_308);
or U6094 (N_6094,N_798,N_2412);
nand U6095 (N_6095,N_1523,N_1849);
or U6096 (N_6096,N_3400,N_180);
nor U6097 (N_6097,N_1911,N_2410);
nor U6098 (N_6098,N_4446,N_204);
nand U6099 (N_6099,N_763,N_1540);
and U6100 (N_6100,N_567,N_1787);
or U6101 (N_6101,N_682,N_2338);
nor U6102 (N_6102,N_687,N_993);
nand U6103 (N_6103,N_1557,N_2289);
xor U6104 (N_6104,N_3762,N_2521);
or U6105 (N_6105,N_4776,N_4692);
nand U6106 (N_6106,N_2856,N_3710);
or U6107 (N_6107,N_4195,N_4131);
nor U6108 (N_6108,N_4358,N_448);
or U6109 (N_6109,N_1943,N_795);
and U6110 (N_6110,N_744,N_2327);
nand U6111 (N_6111,N_2404,N_2035);
or U6112 (N_6112,N_1773,N_2835);
nand U6113 (N_6113,N_4296,N_173);
or U6114 (N_6114,N_1739,N_1703);
nand U6115 (N_6115,N_4892,N_3635);
nand U6116 (N_6116,N_4690,N_1775);
and U6117 (N_6117,N_4409,N_2311);
nor U6118 (N_6118,N_2050,N_3313);
nor U6119 (N_6119,N_1504,N_4491);
or U6120 (N_6120,N_4940,N_2692);
nor U6121 (N_6121,N_1196,N_3851);
nand U6122 (N_6122,N_1,N_4188);
nor U6123 (N_6123,N_4463,N_735);
nand U6124 (N_6124,N_2569,N_4372);
and U6125 (N_6125,N_4575,N_743);
or U6126 (N_6126,N_3198,N_3745);
nand U6127 (N_6127,N_1788,N_1847);
nand U6128 (N_6128,N_1019,N_610);
nor U6129 (N_6129,N_2534,N_4335);
nand U6130 (N_6130,N_2830,N_2554);
nand U6131 (N_6131,N_1759,N_867);
and U6132 (N_6132,N_1819,N_3268);
nor U6133 (N_6133,N_3684,N_3809);
nor U6134 (N_6134,N_1486,N_4282);
or U6135 (N_6135,N_651,N_415);
and U6136 (N_6136,N_2920,N_1148);
or U6137 (N_6137,N_2891,N_1355);
and U6138 (N_6138,N_1502,N_2573);
or U6139 (N_6139,N_2033,N_3885);
nor U6140 (N_6140,N_2578,N_2760);
nand U6141 (N_6141,N_2112,N_2932);
nand U6142 (N_6142,N_4846,N_3102);
or U6143 (N_6143,N_4070,N_3698);
nor U6144 (N_6144,N_3361,N_1390);
or U6145 (N_6145,N_2291,N_4396);
nand U6146 (N_6146,N_4154,N_2457);
nor U6147 (N_6147,N_1707,N_235);
nand U6148 (N_6148,N_892,N_1852);
or U6149 (N_6149,N_4861,N_3511);
and U6150 (N_6150,N_2134,N_4061);
nor U6151 (N_6151,N_2640,N_2039);
and U6152 (N_6152,N_1474,N_1229);
or U6153 (N_6153,N_2312,N_41);
xor U6154 (N_6154,N_948,N_341);
nand U6155 (N_6155,N_2905,N_1120);
and U6156 (N_6156,N_4343,N_3119);
or U6157 (N_6157,N_2283,N_1432);
nand U6158 (N_6158,N_2551,N_2260);
nor U6159 (N_6159,N_1983,N_280);
nand U6160 (N_6160,N_4985,N_4301);
or U6161 (N_6161,N_2791,N_359);
or U6162 (N_6162,N_4848,N_2978);
nor U6163 (N_6163,N_4315,N_7);
nand U6164 (N_6164,N_2414,N_4726);
and U6165 (N_6165,N_4134,N_4882);
and U6166 (N_6166,N_2382,N_4914);
or U6167 (N_6167,N_1121,N_1037);
or U6168 (N_6168,N_3463,N_1055);
and U6169 (N_6169,N_3589,N_896);
or U6170 (N_6170,N_336,N_3459);
nor U6171 (N_6171,N_4857,N_2979);
and U6172 (N_6172,N_2723,N_2606);
nand U6173 (N_6173,N_3299,N_3836);
nor U6174 (N_6174,N_3806,N_3211);
nand U6175 (N_6175,N_2874,N_2607);
and U6176 (N_6176,N_1633,N_851);
or U6177 (N_6177,N_2983,N_4453);
and U6178 (N_6178,N_727,N_2870);
or U6179 (N_6179,N_2564,N_3040);
and U6180 (N_6180,N_521,N_2085);
nor U6181 (N_6181,N_2931,N_1906);
or U6182 (N_6182,N_1452,N_4595);
nor U6183 (N_6183,N_1538,N_21);
and U6184 (N_6184,N_2063,N_712);
nand U6185 (N_6185,N_1582,N_4728);
xor U6186 (N_6186,N_3277,N_226);
xnor U6187 (N_6187,N_2345,N_942);
xnor U6188 (N_6188,N_2647,N_1555);
and U6189 (N_6189,N_2522,N_1277);
or U6190 (N_6190,N_1360,N_4608);
and U6191 (N_6191,N_1853,N_1485);
and U6192 (N_6192,N_186,N_2286);
nand U6193 (N_6193,N_1561,N_4429);
or U6194 (N_6194,N_4705,N_3661);
or U6195 (N_6195,N_3871,N_2399);
xnor U6196 (N_6196,N_4745,N_514);
and U6197 (N_6197,N_3421,N_534);
xor U6198 (N_6198,N_4681,N_4997);
nor U6199 (N_6199,N_1963,N_4445);
nor U6200 (N_6200,N_1071,N_73);
nand U6201 (N_6201,N_2127,N_659);
nor U6202 (N_6202,N_3087,N_1089);
nand U6203 (N_6203,N_4520,N_84);
and U6204 (N_6204,N_4541,N_429);
or U6205 (N_6205,N_2915,N_616);
or U6206 (N_6206,N_2478,N_729);
nand U6207 (N_6207,N_4883,N_4278);
nor U6208 (N_6208,N_2120,N_2757);
or U6209 (N_6209,N_4191,N_2511);
or U6210 (N_6210,N_4753,N_4926);
nand U6211 (N_6211,N_3590,N_3583);
nand U6212 (N_6212,N_1288,N_3913);
and U6213 (N_6213,N_2110,N_1040);
nand U6214 (N_6214,N_1039,N_2193);
or U6215 (N_6215,N_3804,N_4176);
and U6216 (N_6216,N_3565,N_1912);
nor U6217 (N_6217,N_424,N_3218);
nand U6218 (N_6218,N_405,N_3156);
and U6219 (N_6219,N_3121,N_1883);
nor U6220 (N_6220,N_3378,N_656);
or U6221 (N_6221,N_2768,N_2997);
and U6222 (N_6222,N_2696,N_2046);
and U6223 (N_6223,N_3845,N_3451);
and U6224 (N_6224,N_561,N_2184);
and U6225 (N_6225,N_4321,N_4140);
nor U6226 (N_6226,N_3777,N_3238);
nand U6227 (N_6227,N_3229,N_2860);
nor U6228 (N_6228,N_1553,N_4145);
nor U6229 (N_6229,N_3213,N_1754);
or U6230 (N_6230,N_1359,N_3487);
and U6231 (N_6231,N_1643,N_915);
and U6232 (N_6232,N_1340,N_768);
nand U6233 (N_6233,N_2282,N_3507);
nand U6234 (N_6234,N_2518,N_263);
and U6235 (N_6235,N_4063,N_2675);
nand U6236 (N_6236,N_1451,N_504);
and U6237 (N_6237,N_3145,N_674);
nand U6238 (N_6238,N_1524,N_873);
and U6239 (N_6239,N_1298,N_4431);
and U6240 (N_6240,N_1836,N_2116);
or U6241 (N_6241,N_3381,N_395);
and U6242 (N_6242,N_4531,N_1102);
and U6243 (N_6243,N_2445,N_4285);
and U6244 (N_6244,N_2057,N_2698);
or U6245 (N_6245,N_1704,N_3839);
and U6246 (N_6246,N_375,N_2977);
nand U6247 (N_6247,N_2536,N_4944);
nand U6248 (N_6248,N_1866,N_80);
nor U6249 (N_6249,N_3651,N_3944);
xor U6250 (N_6250,N_1167,N_1027);
and U6251 (N_6251,N_1358,N_3220);
and U6252 (N_6252,N_4707,N_1214);
and U6253 (N_6253,N_4259,N_1575);
and U6254 (N_6254,N_3856,N_3125);
nor U6255 (N_6255,N_3041,N_4167);
xor U6256 (N_6256,N_3834,N_1956);
nor U6257 (N_6257,N_3994,N_135);
nand U6258 (N_6258,N_775,N_4231);
nor U6259 (N_6259,N_4908,N_4812);
nor U6260 (N_6260,N_4699,N_1442);
or U6261 (N_6261,N_2323,N_1201);
nor U6262 (N_6262,N_1971,N_2048);
and U6263 (N_6263,N_1831,N_1636);
or U6264 (N_6264,N_2166,N_1835);
or U6265 (N_6265,N_3683,N_1761);
nand U6266 (N_6266,N_451,N_1934);
nor U6267 (N_6267,N_4136,N_4641);
nand U6268 (N_6268,N_903,N_3172);
and U6269 (N_6269,N_1294,N_4467);
and U6270 (N_6270,N_3141,N_4537);
and U6271 (N_6271,N_4274,N_1233);
nand U6272 (N_6272,N_4168,N_2650);
nand U6273 (N_6273,N_2018,N_4365);
nand U6274 (N_6274,N_4669,N_4203);
or U6275 (N_6275,N_3005,N_4527);
or U6276 (N_6276,N_2817,N_3025);
and U6277 (N_6277,N_3446,N_2630);
nor U6278 (N_6278,N_4994,N_2948);
or U6279 (N_6279,N_4480,N_3201);
or U6280 (N_6280,N_739,N_3746);
nor U6281 (N_6281,N_4499,N_4789);
xor U6282 (N_6282,N_4283,N_1108);
or U6283 (N_6283,N_1658,N_2022);
nor U6284 (N_6284,N_4786,N_4314);
nor U6285 (N_6285,N_3064,N_183);
or U6286 (N_6286,N_4577,N_749);
and U6287 (N_6287,N_741,N_3783);
or U6288 (N_6288,N_1926,N_3873);
and U6289 (N_6289,N_4948,N_4731);
nand U6290 (N_6290,N_2880,N_2337);
nand U6291 (N_6291,N_1476,N_4893);
nor U6292 (N_6292,N_1484,N_3474);
and U6293 (N_6293,N_4050,N_2124);
nand U6294 (N_6294,N_3640,N_1324);
nor U6295 (N_6295,N_1678,N_847);
nand U6296 (N_6296,N_3518,N_1141);
nor U6297 (N_6297,N_3555,N_4153);
and U6298 (N_6298,N_2308,N_726);
and U6299 (N_6299,N_4486,N_444);
nor U6300 (N_6300,N_3803,N_4625);
or U6301 (N_6301,N_251,N_3568);
and U6302 (N_6302,N_230,N_790);
nand U6303 (N_6303,N_4458,N_4732);
nand U6304 (N_6304,N_4571,N_2165);
or U6305 (N_6305,N_4634,N_3384);
and U6306 (N_6306,N_2339,N_4472);
or U6307 (N_6307,N_2045,N_376);
or U6308 (N_6308,N_3742,N_247);
nor U6309 (N_6309,N_2754,N_3147);
nand U6310 (N_6310,N_885,N_2191);
and U6311 (N_6311,N_4718,N_115);
and U6312 (N_6312,N_2111,N_4401);
nor U6313 (N_6313,N_2428,N_4495);
nand U6314 (N_6314,N_326,N_4174);
nand U6315 (N_6315,N_1469,N_217);
or U6316 (N_6316,N_3519,N_698);
or U6317 (N_6317,N_4916,N_4355);
or U6318 (N_6318,N_1081,N_1519);
xor U6319 (N_6319,N_2013,N_4101);
or U6320 (N_6320,N_3538,N_760);
nor U6321 (N_6321,N_3869,N_2097);
nand U6322 (N_6322,N_1408,N_891);
and U6323 (N_6323,N_4952,N_4258);
nand U6324 (N_6324,N_2731,N_2176);
or U6325 (N_6325,N_4482,N_966);
nand U6326 (N_6326,N_4738,N_3712);
or U6327 (N_6327,N_4434,N_1296);
nand U6328 (N_6328,N_2015,N_1817);
nor U6329 (N_6329,N_4904,N_2483);
and U6330 (N_6330,N_2820,N_3322);
and U6331 (N_6331,N_3665,N_3026);
nand U6332 (N_6332,N_426,N_1590);
or U6333 (N_6333,N_764,N_4975);
or U6334 (N_6334,N_1578,N_478);
nand U6335 (N_6335,N_2065,N_1362);
nand U6336 (N_6336,N_1069,N_348);
nor U6337 (N_6337,N_862,N_4609);
and U6338 (N_6338,N_2160,N_2697);
or U6339 (N_6339,N_1351,N_2737);
or U6340 (N_6340,N_1373,N_384);
and U6341 (N_6341,N_1095,N_2538);
or U6342 (N_6342,N_83,N_566);
xnor U6343 (N_6343,N_692,N_2610);
and U6344 (N_6344,N_194,N_2902);
or U6345 (N_6345,N_4415,N_23);
nor U6346 (N_6346,N_2886,N_1808);
and U6347 (N_6347,N_585,N_3335);
nand U6348 (N_6348,N_1828,N_3202);
or U6349 (N_6349,N_4332,N_1945);
nor U6350 (N_6350,N_4942,N_2341);
and U6351 (N_6351,N_1689,N_4169);
nor U6352 (N_6352,N_3750,N_88);
nand U6353 (N_6353,N_4501,N_2967);
nand U6354 (N_6354,N_4435,N_1779);
nor U6355 (N_6355,N_1839,N_3039);
and U6356 (N_6356,N_4380,N_3170);
and U6357 (N_6357,N_1218,N_1807);
and U6358 (N_6358,N_785,N_4534);
nor U6359 (N_6359,N_2911,N_2477);
and U6360 (N_6360,N_2386,N_940);
or U6361 (N_6361,N_2092,N_1631);
nand U6362 (N_6362,N_1283,N_3763);
nor U6363 (N_6363,N_3929,N_4288);
or U6364 (N_6364,N_2556,N_2702);
nor U6365 (N_6365,N_960,N_3181);
or U6366 (N_6366,N_1547,N_64);
and U6367 (N_6367,N_665,N_320);
nor U6368 (N_6368,N_1618,N_3622);
nand U6369 (N_6369,N_3606,N_59);
nor U6370 (N_6370,N_4927,N_1026);
nand U6371 (N_6371,N_377,N_536);
or U6372 (N_6372,N_679,N_2364);
or U6373 (N_6373,N_1913,N_4529);
or U6374 (N_6374,N_112,N_3978);
nand U6375 (N_6375,N_4400,N_2484);
nand U6376 (N_6376,N_2162,N_3438);
nand U6377 (N_6377,N_1600,N_54);
nor U6378 (N_6378,N_3625,N_4129);
and U6379 (N_6379,N_1595,N_2752);
nor U6380 (N_6380,N_214,N_3717);
nand U6381 (N_6381,N_4829,N_1259);
or U6382 (N_6382,N_2998,N_455);
nor U6383 (N_6383,N_4454,N_4303);
and U6384 (N_6384,N_3329,N_1316);
nand U6385 (N_6385,N_1181,N_2054);
nand U6386 (N_6386,N_2821,N_1111);
or U6387 (N_6387,N_4397,N_4784);
or U6388 (N_6388,N_4585,N_2685);
and U6389 (N_6389,N_1445,N_425);
or U6390 (N_6390,N_1090,N_3415);
and U6391 (N_6391,N_4737,N_4581);
nand U6392 (N_6392,N_995,N_1472);
and U6393 (N_6393,N_4960,N_4687);
or U6394 (N_6394,N_4646,N_1525);
nor U6395 (N_6395,N_634,N_2859);
nor U6396 (N_6396,N_1391,N_120);
or U6397 (N_6397,N_2304,N_1799);
xor U6398 (N_6398,N_4115,N_2644);
and U6399 (N_6399,N_4546,N_2463);
nor U6400 (N_6400,N_160,N_1859);
nor U6401 (N_6401,N_1042,N_4781);
or U6402 (N_6402,N_3491,N_691);
or U6403 (N_6403,N_4299,N_2479);
nor U6404 (N_6404,N_3977,N_422);
xor U6405 (N_6405,N_1532,N_4193);
and U6406 (N_6406,N_1772,N_2316);
and U6407 (N_6407,N_4836,N_1450);
or U6408 (N_6408,N_185,N_1740);
nand U6409 (N_6409,N_3223,N_4620);
nand U6410 (N_6410,N_1723,N_4678);
and U6411 (N_6411,N_4448,N_19);
nor U6412 (N_6412,N_3758,N_2049);
nand U6413 (N_6413,N_3614,N_932);
nor U6414 (N_6414,N_394,N_3144);
or U6415 (N_6415,N_327,N_1475);
or U6416 (N_6416,N_4031,N_1792);
nand U6417 (N_6417,N_4322,N_3688);
or U6418 (N_6418,N_3676,N_3878);
and U6419 (N_6419,N_140,N_3767);
nor U6420 (N_6420,N_1738,N_1667);
and U6421 (N_6421,N_2910,N_2812);
and U6422 (N_6422,N_2106,N_4643);
and U6423 (N_6423,N_3573,N_4915);
nand U6424 (N_6424,N_3727,N_4566);
or U6425 (N_6425,N_1710,N_2170);
and U6426 (N_6426,N_1318,N_2149);
nor U6427 (N_6427,N_284,N_218);
or U6428 (N_6428,N_3613,N_4685);
nor U6429 (N_6429,N_4582,N_821);
and U6430 (N_6430,N_591,N_4597);
and U6431 (N_6431,N_544,N_1496);
xor U6432 (N_6432,N_1902,N_3423);
or U6433 (N_6433,N_3786,N_1248);
nand U6434 (N_6434,N_3752,N_3191);
nand U6435 (N_6435,N_4084,N_2360);
nand U6436 (N_6436,N_4451,N_3768);
nand U6437 (N_6437,N_1182,N_4462);
xor U6438 (N_6438,N_4427,N_1435);
or U6439 (N_6439,N_29,N_1786);
nor U6440 (N_6440,N_4939,N_3832);
or U6441 (N_6441,N_2652,N_3788);
and U6442 (N_6442,N_1045,N_3854);
nand U6443 (N_6443,N_1607,N_2388);
or U6444 (N_6444,N_1673,N_4177);
nand U6445 (N_6445,N_4394,N_1939);
nor U6446 (N_6446,N_104,N_1372);
nor U6447 (N_6447,N_2100,N_4525);
nor U6448 (N_6448,N_3722,N_4043);
nor U6449 (N_6449,N_543,N_4126);
and U6450 (N_6450,N_2250,N_4704);
nor U6451 (N_6451,N_3755,N_1800);
and U6452 (N_6452,N_2181,N_33);
nand U6453 (N_6453,N_4433,N_2281);
and U6454 (N_6454,N_4033,N_623);
and U6455 (N_6455,N_278,N_2210);
or U6456 (N_6456,N_1725,N_3558);
and U6457 (N_6457,N_2007,N_1334);
and U6458 (N_6458,N_4324,N_1220);
or U6459 (N_6459,N_2448,N_442);
or U6460 (N_6460,N_1602,N_4055);
nor U6461 (N_6461,N_886,N_2660);
and U6462 (N_6462,N_3618,N_291);
and U6463 (N_6463,N_292,N_178);
xnor U6464 (N_6464,N_1896,N_401);
and U6465 (N_6465,N_4025,N_3252);
or U6466 (N_6466,N_1293,N_2828);
and U6467 (N_6467,N_1677,N_1114);
nand U6468 (N_6468,N_4373,N_3481);
nor U6469 (N_6469,N_4393,N_2255);
or U6470 (N_6470,N_260,N_2732);
nand U6471 (N_6471,N_2074,N_1378);
or U6472 (N_6472,N_3349,N_221);
and U6473 (N_6473,N_2883,N_551);
and U6474 (N_6474,N_1285,N_4421);
nor U6475 (N_6475,N_1691,N_2620);
nand U6476 (N_6476,N_1614,N_2139);
and U6477 (N_6477,N_2990,N_3936);
or U6478 (N_6478,N_4163,N_600);
or U6479 (N_6479,N_3893,N_3572);
and U6480 (N_6480,N_3074,N_1209);
nor U6481 (N_6481,N_3801,N_618);
or U6482 (N_6482,N_1076,N_2);
nor U6483 (N_6483,N_2274,N_152);
nand U6484 (N_6484,N_4724,N_3109);
nand U6485 (N_6485,N_3065,N_1834);
or U6486 (N_6486,N_379,N_78);
or U6487 (N_6487,N_502,N_67);
or U6488 (N_6488,N_4379,N_498);
nor U6489 (N_6489,N_3608,N_2137);
or U6490 (N_6490,N_952,N_4248);
nor U6491 (N_6491,N_3082,N_4958);
nand U6492 (N_6492,N_3811,N_3594);
and U6493 (N_6493,N_2411,N_2984);
nand U6494 (N_6494,N_2218,N_1821);
nand U6495 (N_6495,N_1062,N_90);
and U6496 (N_6496,N_1999,N_275);
nor U6497 (N_6497,N_4831,N_242);
and U6498 (N_6498,N_1441,N_287);
nand U6499 (N_6499,N_4524,N_1124);
or U6500 (N_6500,N_3339,N_1375);
nor U6501 (N_6501,N_3077,N_3630);
nor U6502 (N_6502,N_523,N_3597);
nand U6503 (N_6503,N_4356,N_3034);
xnor U6504 (N_6504,N_4468,N_3137);
nor U6505 (N_6505,N_2434,N_1860);
and U6506 (N_6506,N_3447,N_1001);
nand U6507 (N_6507,N_315,N_4592);
or U6508 (N_6508,N_1135,N_2547);
or U6509 (N_6509,N_411,N_1766);
nand U6510 (N_6510,N_423,N_354);
xor U6511 (N_6511,N_2464,N_2387);
nand U6512 (N_6512,N_2942,N_1718);
nand U6513 (N_6513,N_1830,N_1988);
or U6514 (N_6514,N_1846,N_2727);
nor U6515 (N_6515,N_4856,N_3531);
nand U6516 (N_6516,N_4439,N_4823);
nand U6517 (N_6517,N_4413,N_594);
or U6518 (N_6518,N_4437,N_1116);
nor U6519 (N_6519,N_3553,N_4987);
or U6520 (N_6520,N_1144,N_4764);
nand U6521 (N_6521,N_2762,N_2232);
nand U6522 (N_6522,N_1199,N_4325);
and U6523 (N_6523,N_809,N_3981);
nor U6524 (N_6524,N_1871,N_1543);
nor U6525 (N_6525,N_4992,N_1550);
nand U6526 (N_6526,N_300,N_364);
nand U6527 (N_6527,N_1498,N_2090);
or U6528 (N_6528,N_3584,N_4328);
and U6529 (N_6529,N_2152,N_4930);
and U6530 (N_6530,N_1079,N_4485);
nor U6531 (N_6531,N_597,N_2881);
nand U6532 (N_6532,N_4666,N_3235);
or U6533 (N_6533,N_1096,N_3963);
nand U6534 (N_6534,N_4262,N_412);
nor U6535 (N_6535,N_3356,N_824);
nand U6536 (N_6536,N_3566,N_3825);
and U6537 (N_6537,N_1597,N_4272);
nand U6538 (N_6538,N_753,N_3850);
nor U6539 (N_6539,N_1891,N_4046);
and U6540 (N_6540,N_1715,N_4584);
and U6541 (N_6541,N_2305,N_658);
nand U6542 (N_6542,N_159,N_2605);
nand U6543 (N_6543,N_2064,N_2974);
nor U6544 (N_6544,N_2144,N_74);
xor U6545 (N_6545,N_4352,N_4290);
or U6546 (N_6546,N_4357,N_3582);
xor U6547 (N_6547,N_1975,N_4340);
and U6548 (N_6548,N_607,N_1848);
nand U6549 (N_6549,N_3315,N_3336);
or U6550 (N_6550,N_4142,N_3013);
nand U6551 (N_6551,N_1142,N_4130);
or U6552 (N_6552,N_351,N_316);
nand U6553 (N_6553,N_89,N_3015);
or U6554 (N_6554,N_1460,N_3236);
and U6555 (N_6555,N_4652,N_224);
nor U6556 (N_6556,N_1692,N_262);
and U6557 (N_6557,N_4638,N_253);
and U6558 (N_6558,N_4689,N_72);
and U6559 (N_6559,N_747,N_4141);
nand U6560 (N_6560,N_4565,N_2572);
or U6561 (N_6561,N_2571,N_3734);
or U6562 (N_6562,N_4762,N_179);
nand U6563 (N_6563,N_2520,N_2243);
nor U6564 (N_6564,N_2153,N_3990);
or U6565 (N_6565,N_877,N_1893);
and U6566 (N_6566,N_1158,N_4068);
and U6567 (N_6567,N_3736,N_716);
nand U6568 (N_6568,N_3215,N_3135);
nand U6569 (N_6569,N_2336,N_2066);
or U6570 (N_6570,N_980,N_4099);
and U6571 (N_6571,N_4530,N_2023);
or U6572 (N_6572,N_1091,N_4680);
and U6573 (N_6573,N_4086,N_4506);
nor U6574 (N_6574,N_3894,N_2562);
nor U6575 (N_6575,N_4518,N_4769);
nand U6576 (N_6576,N_2135,N_946);
nor U6577 (N_6577,N_1405,N_2199);
and U6578 (N_6578,N_2892,N_4430);
nand U6579 (N_6579,N_652,N_3439);
and U6580 (N_6580,N_701,N_419);
or U6581 (N_6581,N_4659,N_2238);
nor U6582 (N_6582,N_2845,N_3093);
nor U6583 (N_6583,N_4341,N_3103);
nand U6584 (N_6584,N_590,N_1261);
nor U6585 (N_6585,N_133,N_1088);
and U6586 (N_6586,N_2994,N_1661);
or U6587 (N_6587,N_484,N_3178);
nand U6588 (N_6588,N_1130,N_462);
nand U6589 (N_6589,N_2636,N_170);
nand U6590 (N_6590,N_3702,N_1509);
nand U6591 (N_6591,N_4474,N_467);
or U6592 (N_6592,N_1172,N_1099);
and U6593 (N_6593,N_2851,N_2711);
nand U6594 (N_6594,N_1465,N_4676);
or U6595 (N_6595,N_4964,N_2855);
and U6596 (N_6596,N_1224,N_1683);
nand U6597 (N_6597,N_3575,N_3165);
or U6598 (N_6598,N_2098,N_4759);
nand U6599 (N_6599,N_2531,N_332);
nand U6600 (N_6600,N_4027,N_400);
nor U6601 (N_6601,N_3535,N_2865);
or U6602 (N_6602,N_1179,N_643);
and U6603 (N_6603,N_3569,N_2461);
nand U6604 (N_6604,N_4655,N_4175);
or U6605 (N_6605,N_2667,N_57);
and U6606 (N_6606,N_2709,N_2747);
or U6607 (N_6607,N_1488,N_4819);
nor U6608 (N_6608,N_774,N_4508);
nor U6609 (N_6609,N_3244,N_1317);
and U6610 (N_6610,N_3155,N_3957);
and U6611 (N_6611,N_1546,N_4550);
or U6612 (N_6612,N_4826,N_3028);
nand U6613 (N_6613,N_357,N_2266);
nand U6614 (N_6614,N_1570,N_4327);
nand U6615 (N_6615,N_3743,N_3323);
or U6616 (N_6616,N_1867,N_550);
or U6617 (N_6617,N_3230,N_517);
and U6618 (N_6618,N_724,N_1533);
and U6619 (N_6619,N_1208,N_1666);
and U6620 (N_6620,N_1107,N_4117);
and U6621 (N_6621,N_3194,N_3076);
nor U6622 (N_6622,N_3794,N_3699);
nor U6623 (N_6623,N_4228,N_1180);
or U6624 (N_6624,N_3780,N_3484);
nand U6625 (N_6625,N_4999,N_500);
or U6626 (N_6626,N_3222,N_4257);
nor U6627 (N_6627,N_1927,N_3457);
nand U6628 (N_6628,N_779,N_1735);
or U6629 (N_6629,N_3821,N_3149);
and U6630 (N_6630,N_4094,N_4502);
nor U6631 (N_6631,N_2884,N_2934);
or U6632 (N_6632,N_3321,N_3483);
and U6633 (N_6633,N_845,N_8);
or U6634 (N_6634,N_671,N_4757);
nand U6635 (N_6635,N_1242,N_3274);
or U6636 (N_6636,N_4853,N_2563);
nor U6637 (N_6637,N_4850,N_4330);
nand U6638 (N_6638,N_2352,N_571);
or U6639 (N_6639,N_2969,N_893);
nor U6640 (N_6640,N_4605,N_4037);
or U6641 (N_6641,N_3619,N_3312);
or U6642 (N_6642,N_1282,N_3909);
or U6643 (N_6643,N_466,N_4017);
nand U6644 (N_6644,N_3610,N_4105);
or U6645 (N_6645,N_266,N_3561);
nand U6646 (N_6646,N_2235,N_4825);
or U6647 (N_6647,N_2925,N_123);
or U6648 (N_6648,N_4563,N_1342);
nand U6649 (N_6649,N_3972,N_4479);
or U6650 (N_6650,N_2776,N_3587);
xnor U6651 (N_6651,N_85,N_1407);
or U6652 (N_6652,N_4190,N_1426);
xnor U6653 (N_6653,N_3150,N_175);
and U6654 (N_6654,N_165,N_398);
nand U6655 (N_6655,N_4395,N_1230);
nor U6656 (N_6656,N_1017,N_2868);
nand U6657 (N_6657,N_1531,N_4783);
nor U6658 (N_6658,N_1403,N_1760);
or U6659 (N_6659,N_3667,N_1565);
nor U6660 (N_6660,N_2405,N_810);
nand U6661 (N_6661,N_897,N_1216);
nor U6662 (N_6662,N_3095,N_1776);
xor U6663 (N_6663,N_2351,N_2814);
and U6664 (N_6664,N_4230,N_2195);
nand U6665 (N_6665,N_3512,N_3348);
and U6666 (N_6666,N_713,N_1178);
and U6667 (N_6667,N_483,N_1093);
and U6668 (N_6668,N_822,N_4209);
and U6669 (N_6669,N_4353,N_742);
nor U6670 (N_6670,N_936,N_1534);
nand U6671 (N_6671,N_737,N_4058);
and U6672 (N_6672,N_2375,N_4919);
or U6673 (N_6673,N_491,N_4963);
nor U6674 (N_6674,N_1205,N_3542);
or U6675 (N_6675,N_3485,N_1284);
and U6676 (N_6676,N_3241,N_1940);
and U6677 (N_6677,N_1022,N_238);
nand U6678 (N_6678,N_2084,N_2008);
or U6679 (N_6679,N_3425,N_3242);
nand U6680 (N_6680,N_961,N_144);
and U6681 (N_6681,N_3729,N_556);
and U6682 (N_6682,N_3383,N_45);
or U6683 (N_6683,N_1919,N_529);
nand U6684 (N_6684,N_47,N_2016);
xnor U6685 (N_6685,N_433,N_4806);
or U6686 (N_6686,N_3251,N_3818);
nand U6687 (N_6687,N_2777,N_3641);
or U6688 (N_6688,N_1985,N_2625);
and U6689 (N_6689,N_3148,N_4469);
and U6690 (N_6690,N_2525,N_1329);
nor U6691 (N_6691,N_4899,N_3666);
and U6692 (N_6692,N_4574,N_4233);
and U6693 (N_6693,N_3760,N_4227);
nor U6694 (N_6694,N_2435,N_198);
nor U6695 (N_6695,N_2373,N_312);
or U6696 (N_6696,N_4822,N_3646);
and U6697 (N_6697,N_3576,N_1824);
or U6698 (N_6698,N_700,N_2156);
nand U6699 (N_6699,N_4122,N_1264);
and U6700 (N_6700,N_4234,N_1327);
and U6701 (N_6701,N_546,N_4273);
or U6702 (N_6702,N_1308,N_3741);
nand U6703 (N_6703,N_908,N_1168);
and U6704 (N_6704,N_4633,N_3352);
nor U6705 (N_6705,N_2604,N_4578);
or U6706 (N_6706,N_1032,N_3106);
nor U6707 (N_6707,N_14,N_161);
nand U6708 (N_6708,N_4085,N_1306);
xor U6709 (N_6709,N_2258,N_4012);
xor U6710 (N_6710,N_256,N_3306);
and U6711 (N_6711,N_3861,N_4478);
and U6712 (N_6712,N_3759,N_1511);
and U6713 (N_6713,N_593,N_4271);
and U6714 (N_6714,N_4855,N_4810);
or U6715 (N_6715,N_4042,N_2317);
and U6716 (N_6716,N_541,N_4742);
nand U6717 (N_6717,N_2334,N_1651);
nor U6718 (N_6718,N_169,N_3773);
and U6719 (N_6719,N_3193,N_3917);
or U6720 (N_6720,N_3187,N_4165);
or U6721 (N_6721,N_2744,N_3374);
and U6722 (N_6722,N_2981,N_1478);
nand U6723 (N_6723,N_714,N_1455);
and U6724 (N_6724,N_95,N_3440);
or U6725 (N_6725,N_2913,N_507);
nor U6726 (N_6726,N_783,N_4715);
or U6727 (N_6727,N_3536,N_1002);
and U6728 (N_6728,N_1260,N_1545);
or U6729 (N_6729,N_2684,N_1136);
nor U6730 (N_6730,N_3347,N_4238);
and U6731 (N_6731,N_1964,N_2121);
nand U6732 (N_6732,N_4760,N_2552);
nand U6733 (N_6733,N_1556,N_1423);
and U6734 (N_6734,N_856,N_2026);
and U6735 (N_6735,N_3669,N_4149);
and U6736 (N_6736,N_3099,N_4552);
nand U6737 (N_6737,N_1119,N_641);
and U6738 (N_6738,N_890,N_3168);
nand U6739 (N_6739,N_1417,N_1741);
and U6740 (N_6740,N_586,N_3962);
nor U6741 (N_6741,N_2681,N_2866);
nand U6742 (N_6742,N_2515,N_2072);
nand U6743 (N_6743,N_3011,N_3020);
and U6744 (N_6744,N_3303,N_2369);
or U6745 (N_6745,N_3895,N_3774);
and U6746 (N_6746,N_3294,N_1827);
nand U6747 (N_6747,N_4801,N_4777);
nor U6748 (N_6748,N_3271,N_4654);
or U6749 (N_6749,N_270,N_3973);
nor U6750 (N_6750,N_3604,N_4013);
nor U6751 (N_6751,N_990,N_984);
nor U6752 (N_6752,N_3090,N_3456);
xnor U6753 (N_6753,N_4371,N_2356);
nor U6754 (N_6754,N_1297,N_4112);
nor U6755 (N_6755,N_2229,N_1537);
or U6756 (N_6756,N_129,N_3835);
nor U6757 (N_6757,N_709,N_4432);
nand U6758 (N_6758,N_1699,N_2594);
nand U6759 (N_6759,N_1206,N_103);
nor U6760 (N_6760,N_1246,N_2010);
nand U6761 (N_6761,N_4477,N_3209);
nor U6762 (N_6762,N_4164,N_16);
nand U6763 (N_6763,N_4102,N_1805);
and U6764 (N_6764,N_4289,N_1117);
and U6765 (N_6765,N_1862,N_4710);
nand U6766 (N_6766,N_3733,N_2621);
xor U6767 (N_6767,N_2400,N_3401);
or U6768 (N_6768,N_531,N_3373);
or U6769 (N_6769,N_3086,N_446);
nand U6770 (N_6770,N_2704,N_4903);
or U6771 (N_6771,N_4840,N_4934);
and U6772 (N_6772,N_1982,N_4775);
and U6773 (N_6773,N_149,N_92);
or U6774 (N_6774,N_1197,N_2233);
or U6775 (N_6775,N_55,N_2738);
xor U6776 (N_6776,N_2265,N_3185);
or U6777 (N_6777,N_3067,N_2912);
and U6778 (N_6778,N_4323,N_3289);
and U6779 (N_6779,N_277,N_3770);
nor U6780 (N_6780,N_2504,N_1980);
nand U6781 (N_6781,N_62,N_1733);
nor U6782 (N_6782,N_2513,N_319);
nor U6783 (N_6783,N_3631,N_4663);
nor U6784 (N_6784,N_154,N_1981);
and U6785 (N_6785,N_4734,N_3143);
nand U6786 (N_6786,N_3901,N_4658);
and U6787 (N_6787,N_592,N_4549);
and U6788 (N_6788,N_2367,N_4901);
or U6789 (N_6789,N_670,N_617);
nor U6790 (N_6790,N_4803,N_4526);
nor U6791 (N_6791,N_579,N_2292);
or U6792 (N_6792,N_647,N_2083);
nand U6793 (N_6793,N_3790,N_557);
nor U6794 (N_6794,N_4561,N_2211);
or U6795 (N_6795,N_2946,N_2996);
xor U6796 (N_6796,N_250,N_3838);
nor U6797 (N_6797,N_4593,N_240);
or U6798 (N_6798,N_1838,N_3228);
or U6799 (N_6799,N_3611,N_565);
and U6800 (N_6800,N_3450,N_4602);
xnor U6801 (N_6801,N_3935,N_1468);
nand U6802 (N_6802,N_2040,N_4457);
and U6803 (N_6803,N_792,N_4420);
nand U6804 (N_6804,N_675,N_346);
or U6805 (N_6805,N_1238,N_124);
nor U6806 (N_6806,N_819,N_1068);
or U6807 (N_6807,N_171,N_2167);
and U6808 (N_6808,N_1742,N_156);
nand U6809 (N_6809,N_3410,N_1592);
nand U6810 (N_6810,N_3993,N_1312);
nand U6811 (N_6811,N_488,N_2466);
or U6812 (N_6812,N_469,N_1020);
and U6813 (N_6813,N_4494,N_1908);
nor U6814 (N_6814,N_4399,N_3907);
nand U6815 (N_6815,N_2894,N_3560);
nor U6816 (N_6816,N_2726,N_1870);
nand U6817 (N_6817,N_871,N_4586);
xnor U6818 (N_6818,N_3304,N_865);
or U6819 (N_6819,N_1494,N_1784);
or U6820 (N_6820,N_2480,N_416);
nand U6821 (N_6821,N_2805,N_4405);
nor U6822 (N_6822,N_4067,N_2467);
nor U6823 (N_6823,N_828,N_1687);
or U6824 (N_6824,N_3896,N_2508);
nand U6825 (N_6825,N_1353,N_699);
and U6826 (N_6826,N_3820,N_917);
or U6827 (N_6827,N_520,N_516);
or U6828 (N_6828,N_1899,N_3465);
nand U6829 (N_6829,N_4694,N_4599);
and U6830 (N_6830,N_2904,N_1448);
nand U6831 (N_6831,N_4749,N_2561);
and U6832 (N_6832,N_3054,N_1463);
xnor U6833 (N_6833,N_4221,N_2205);
xor U6834 (N_6834,N_3744,N_3616);
and U6835 (N_6835,N_4627,N_2839);
and U6836 (N_6836,N_490,N_4968);
nand U6837 (N_6837,N_362,N_2956);
nor U6838 (N_6838,N_858,N_4339);
nand U6839 (N_6839,N_3586,N_3364);
or U6840 (N_6840,N_3549,N_3254);
nand U6841 (N_6841,N_1780,N_3146);
nand U6842 (N_6842,N_1887,N_4349);
or U6843 (N_6843,N_888,N_309);
nand U6844 (N_6844,N_1150,N_1006);
or U6845 (N_6845,N_4384,N_1046);
or U6846 (N_6846,N_2639,N_4408);
xor U6847 (N_6847,N_439,N_2117);
nand U6848 (N_6848,N_3551,N_2069);
and U6849 (N_6849,N_1782,N_906);
or U6850 (N_6850,N_2177,N_3506);
and U6851 (N_6851,N_3286,N_2576);
or U6852 (N_6852,N_4923,N_3246);
nor U6853 (N_6853,N_4830,N_882);
nor U6854 (N_6854,N_285,N_1907);
nand U6855 (N_6855,N_1558,N_4381);
or U6856 (N_6856,N_4928,N_864);
nand U6857 (N_6857,N_2999,N_4878);
nand U6858 (N_6858,N_1113,N_4452);
or U6859 (N_6859,N_457,N_3642);
and U6860 (N_6860,N_3318,N_4938);
and U6861 (N_6861,N_4695,N_937);
or U6862 (N_6862,N_4354,N_4180);
or U6863 (N_6863,N_1477,N_1946);
and U6864 (N_6864,N_4254,N_1123);
and U6865 (N_6865,N_3445,N_2280);
nor U6866 (N_6866,N_3585,N_110);
or U6867 (N_6867,N_621,N_1479);
and U6868 (N_6868,N_816,N_3281);
or U6869 (N_6869,N_369,N_1444);
nor U6870 (N_6870,N_2689,N_766);
or U6871 (N_6871,N_978,N_2833);
nor U6872 (N_6872,N_343,N_638);
nand U6873 (N_6873,N_43,N_2301);
or U6874 (N_6874,N_3662,N_2546);
xor U6875 (N_6875,N_3887,N_4199);
nand U6876 (N_6876,N_1816,N_1471);
or U6877 (N_6877,N_1909,N_1422);
and U6878 (N_6878,N_4821,N_3951);
and U6879 (N_6879,N_3173,N_1837);
or U6880 (N_6880,N_3104,N_4116);
nand U6881 (N_6881,N_3753,N_587);
nand U6882 (N_6882,N_1420,N_3050);
or U6883 (N_6883,N_4459,N_2476);
nor U6884 (N_6884,N_2788,N_909);
nand U6885 (N_6885,N_2671,N_1955);
or U6886 (N_6886,N_720,N_81);
and U6887 (N_6887,N_3939,N_4048);
nand U6888 (N_6888,N_1675,N_1175);
and U6889 (N_6889,N_3663,N_3042);
nand U6890 (N_6890,N_558,N_719);
and U6891 (N_6891,N_2673,N_2872);
nor U6892 (N_6892,N_1157,N_258);
nand U6893 (N_6893,N_3858,N_114);
nand U6894 (N_6894,N_1263,N_3837);
nand U6895 (N_6895,N_2548,N_3682);
nor U6896 (N_6896,N_1563,N_119);
nand U6897 (N_6897,N_497,N_4073);
nor U6898 (N_6898,N_3479,N_3735);
and U6899 (N_6899,N_2635,N_1268);
and U6900 (N_6900,N_3931,N_833);
or U6901 (N_6901,N_3376,N_4253);
nor U6902 (N_6902,N_3208,N_2080);
and U6903 (N_6903,N_3097,N_1004);
or U6904 (N_6904,N_870,N_2300);
or U6905 (N_6905,N_1336,N_2420);
nor U6906 (N_6906,N_2537,N_486);
or U6907 (N_6907,N_1931,N_2507);
or U6908 (N_6908,N_3781,N_3874);
and U6909 (N_6909,N_3634,N_195);
xnor U6910 (N_6910,N_302,N_254);
and U6911 (N_6911,N_3084,N_3436);
and U6912 (N_6912,N_1065,N_3824);
nor U6913 (N_6913,N_4712,N_3341);
nand U6914 (N_6914,N_96,N_938);
nand U6915 (N_6915,N_3908,N_2068);
and U6916 (N_6916,N_3344,N_431);
or U6917 (N_6917,N_4966,N_387);
nand U6918 (N_6918,N_2081,N_1466);
xnor U6919 (N_6919,N_4843,N_1923);
nor U6920 (N_6920,N_4906,N_3656);
nand U6921 (N_6921,N_3726,N_1986);
nand U6922 (N_6922,N_1634,N_874);
nor U6923 (N_6923,N_1010,N_904);
nor U6924 (N_6924,N_3945,N_1737);
nor U6925 (N_6925,N_3903,N_3612);
and U6926 (N_6926,N_3075,N_2680);
nor U6927 (N_6927,N_1295,N_535);
or U6928 (N_6928,N_404,N_2792);
or U6929 (N_6929,N_1152,N_3892);
nand U6930 (N_6930,N_4648,N_153);
nand U6931 (N_6931,N_1753,N_1567);
nor U6932 (N_6932,N_1767,N_3370);
or U6933 (N_6933,N_142,N_1984);
nor U6934 (N_6934,N_3174,N_3723);
or U6935 (N_6935,N_1749,N_2637);
or U6936 (N_6936,N_3486,N_2204);
or U6937 (N_6937,N_298,N_609);
nand U6938 (N_6938,N_1104,N_4879);
nor U6939 (N_6939,N_818,N_3442);
and U6940 (N_6940,N_4673,N_4143);
or U6941 (N_6941,N_1851,N_231);
or U6942 (N_6942,N_3161,N_2565);
nand U6943 (N_6943,N_63,N_3711);
nand U6944 (N_6944,N_2755,N_811);
nand U6945 (N_6945,N_2895,N_4750);
or U6946 (N_6946,N_3910,N_4889);
nor U6947 (N_6947,N_3690,N_476);
nor U6948 (N_6948,N_2126,N_1777);
nor U6949 (N_6949,N_3189,N_2487);
or U6950 (N_6950,N_684,N_1289);
nand U6951 (N_6951,N_939,N_1507);
nand U6952 (N_6952,N_1387,N_456);
nand U6953 (N_6953,N_1215,N_4317);
and U6954 (N_6954,N_3346,N_4751);
or U6955 (N_6955,N_2770,N_1746);
and U6956 (N_6956,N_4404,N_4128);
nor U6957 (N_6957,N_1803,N_1122);
xnor U6958 (N_6958,N_588,N_4766);
and U6959 (N_6959,N_632,N_2418);
nor U6960 (N_6960,N_3941,N_3265);
and U6961 (N_6961,N_3655,N_681);
or U6962 (N_6962,N_4402,N_4721);
nor U6963 (N_6963,N_368,N_4090);
and U6964 (N_6964,N_3881,N_957);
or U6965 (N_6965,N_158,N_628);
and U6966 (N_6966,N_1314,N_463);
or U6967 (N_6967,N_2324,N_2397);
or U6968 (N_6968,N_2430,N_2924);
nor U6969 (N_6969,N_2315,N_4205);
nor U6970 (N_6970,N_505,N_3514);
xnor U6971 (N_6971,N_3911,N_2719);
or U6972 (N_6972,N_1154,N_2656);
or U6973 (N_6973,N_1287,N_4201);
nand U6974 (N_6974,N_2208,N_1581);
nand U6975 (N_6975,N_4772,N_3668);
and U6976 (N_6976,N_1564,N_233);
nor U6977 (N_6977,N_3942,N_769);
nand U6978 (N_6978,N_1223,N_2073);
nand U6979 (N_6979,N_4224,N_4307);
nand U6980 (N_6980,N_1781,N_631);
nand U6981 (N_6981,N_4436,N_3637);
or U6982 (N_6982,N_27,N_3813);
nor U6983 (N_6983,N_3509,N_3657);
nor U6984 (N_6984,N_4211,N_3623);
and U6985 (N_6985,N_3390,N_2517);
or U6986 (N_6986,N_1080,N_1140);
or U6987 (N_6987,N_385,N_3636);
or U6988 (N_6988,N_4032,N_4120);
or U6989 (N_6989,N_3449,N_454);
and U6990 (N_6990,N_3175,N_1210);
or U6991 (N_6991,N_2574,N_1974);
nand U6992 (N_6992,N_1503,N_428);
and U6993 (N_6993,N_2359,N_3081);
or U6994 (N_6994,N_3233,N_863);
and U6995 (N_6995,N_4591,N_655);
and U6996 (N_6996,N_605,N_3926);
nand U6997 (N_6997,N_868,N_717);
nor U6998 (N_6998,N_261,N_1810);
or U6999 (N_6999,N_2968,N_881);
nor U7000 (N_7000,N_1483,N_3160);
nor U7001 (N_7001,N_3113,N_2593);
nand U7002 (N_7002,N_1419,N_3120);
nand U7003 (N_7003,N_4078,N_2765);
or U7004 (N_7004,N_2275,N_2365);
nor U7005 (N_7005,N_4657,N_4598);
and U7006 (N_7006,N_4119,N_3426);
nor U7007 (N_7007,N_1185,N_1587);
nor U7008 (N_7008,N_246,N_1094);
xnor U7009 (N_7009,N_2545,N_3411);
nand U7010 (N_7010,N_2850,N_1231);
and U7011 (N_7011,N_2287,N_3316);
xnor U7012 (N_7012,N_1243,N_4946);
and U7013 (N_7013,N_2789,N_595);
or U7014 (N_7014,N_532,N_108);
or U7015 (N_7015,N_381,N_1622);
nor U7016 (N_7016,N_805,N_555);
nor U7017 (N_7017,N_2076,N_1920);
and U7018 (N_7018,N_2197,N_3270);
and U7019 (N_7019,N_1882,N_3275);
nand U7020 (N_7020,N_4304,N_3388);
or U7021 (N_7021,N_639,N_4651);
nor U7022 (N_7022,N_2043,N_2532);
or U7023 (N_7023,N_4392,N_2570);
and U7024 (N_7024,N_3038,N_366);
nor U7025 (N_7025,N_3368,N_299);
or U7026 (N_7026,N_4912,N_68);
and U7027 (N_7027,N_4981,N_3324);
nand U7028 (N_7028,N_3675,N_3522);
and U7029 (N_7029,N_2374,N_234);
or U7030 (N_7030,N_1623,N_4138);
nor U7031 (N_7031,N_2958,N_1235);
nand U7032 (N_7032,N_1979,N_1843);
and U7033 (N_7033,N_4875,N_4218);
or U7034 (N_7034,N_10,N_1319);
or U7035 (N_7035,N_977,N_1369);
or U7036 (N_7036,N_1542,N_2735);
and U7037 (N_7037,N_269,N_796);
and U7038 (N_7038,N_1915,N_3855);
or U7039 (N_7039,N_317,N_680);
or U7040 (N_7040,N_3397,N_3151);
nor U7041 (N_7041,N_2972,N_1708);
or U7042 (N_7042,N_4735,N_2331);
and U7043 (N_7043,N_2164,N_2514);
or U7044 (N_7044,N_4945,N_3127);
or U7045 (N_7045,N_3946,N_272);
or U7046 (N_7046,N_4309,N_2519);
and U7047 (N_7047,N_1085,N_3626);
nand U7048 (N_7048,N_4714,N_1060);
and U7049 (N_7049,N_106,N_4716);
or U7050 (N_7050,N_4891,N_2172);
or U7051 (N_7051,N_4570,N_3533);
and U7052 (N_7052,N_2499,N_814);
or U7053 (N_7053,N_4514,N_4334);
nand U7054 (N_7054,N_981,N_861);
nand U7055 (N_7055,N_211,N_1572);
nand U7056 (N_7056,N_147,N_2823);
or U7057 (N_7057,N_494,N_840);
and U7058 (N_7058,N_17,N_1501);
and U7059 (N_7059,N_2456,N_4943);
or U7060 (N_7060,N_3823,N_3999);
nand U7061 (N_7061,N_318,N_4424);
nand U7062 (N_7062,N_2257,N_646);
or U7063 (N_7063,N_2313,N_927);
or U7064 (N_7064,N_3308,N_2676);
nor U7065 (N_7065,N_3964,N_3591);
or U7066 (N_7066,N_1724,N_3433);
or U7067 (N_7067,N_4886,N_781);
or U7068 (N_7068,N_2269,N_1726);
nor U7069 (N_7069,N_1244,N_3797);
nor U7070 (N_7070,N_3959,N_1604);
xnor U7071 (N_7071,N_4359,N_134);
nor U7072 (N_7072,N_1176,N_4847);
or U7073 (N_7073,N_3497,N_1105);
or U7074 (N_7074,N_2348,N_4990);
and U7075 (N_7075,N_4809,N_1783);
nor U7076 (N_7076,N_598,N_1320);
nor U7077 (N_7077,N_471,N_4015);
and U7078 (N_7078,N_578,N_3498);
nand U7079 (N_7079,N_2038,N_3815);
or U7080 (N_7080,N_842,N_3601);
and U7081 (N_7081,N_3867,N_1748);
and U7082 (N_7082,N_2353,N_3609);
and U7083 (N_7083,N_4982,N_1487);
nand U7084 (N_7084,N_650,N_1857);
nand U7085 (N_7085,N_3581,N_4311);
nor U7086 (N_7086,N_2115,N_1394);
nor U7087 (N_7087,N_1521,N_3338);
and U7088 (N_7088,N_3731,N_2841);
nand U7089 (N_7089,N_297,N_4887);
nor U7090 (N_7090,N_2733,N_4898);
xor U7091 (N_7091,N_3248,N_382);
or U7092 (N_7092,N_1012,N_2807);
nor U7093 (N_7093,N_3649,N_3124);
and U7094 (N_7094,N_2746,N_4267);
or U7095 (N_7095,N_1936,N_3351);
and U7096 (N_7096,N_2658,N_4444);
or U7097 (N_7097,N_1757,N_2665);
nand U7098 (N_7098,N_1804,N_1845);
nor U7099 (N_7099,N_2333,N_1183);
nor U7100 (N_7100,N_3707,N_4755);
nor U7101 (N_7101,N_1549,N_1937);
and U7102 (N_7102,N_3310,N_3404);
xor U7103 (N_7103,N_4331,N_954);
nand U7104 (N_7104,N_3891,N_499);
nor U7105 (N_7105,N_852,N_3570);
nor U7106 (N_7106,N_1953,N_695);
nor U7107 (N_7107,N_3134,N_3023);
and U7108 (N_7108,N_902,N_667);
nor U7109 (N_7109,N_3740,N_4144);
nand U7110 (N_7110,N_307,N_4684);
nand U7111 (N_7111,N_4725,N_189);
or U7112 (N_7112,N_2226,N_666);
nor U7113 (N_7113,N_3593,N_4302);
and U7114 (N_7114,N_693,N_438);
and U7115 (N_7115,N_1453,N_2142);
nor U7116 (N_7116,N_2567,N_2529);
or U7117 (N_7117,N_3730,N_991);
nand U7118 (N_7118,N_568,N_440);
or U7119 (N_7119,N_465,N_4007);
nand U7120 (N_7120,N_4368,N_664);
nor U7121 (N_7121,N_2729,N_1706);
nor U7122 (N_7122,N_2584,N_1436);
nand U7123 (N_7123,N_1132,N_2279);
nor U7124 (N_7124,N_1962,N_1366);
nor U7125 (N_7125,N_757,N_2653);
and U7126 (N_7126,N_1262,N_2491);
and U7127 (N_7127,N_3681,N_2816);
nor U7128 (N_7128,N_596,N_1007);
and U7129 (N_7129,N_2602,N_3588);
and U7130 (N_7130,N_4277,N_4006);
and U7131 (N_7131,N_4988,N_1745);
and U7132 (N_7132,N_449,N_2846);
nor U7133 (N_7133,N_4589,N_4310);
nand U7134 (N_7134,N_2496,N_199);
or U7135 (N_7135,N_1795,N_4814);
nor U7136 (N_7136,N_4124,N_2838);
nor U7137 (N_7137,N_1627,N_1028);
and U7138 (N_7138,N_1765,N_2991);
nor U7139 (N_7139,N_1978,N_2272);
or U7140 (N_7140,N_2973,N_4896);
or U7141 (N_7141,N_2019,N_4679);
or U7142 (N_7142,N_619,N_50);
or U7143 (N_7143,N_205,N_2446);
and U7144 (N_7144,N_3164,N_2786);
nand U7145 (N_7145,N_2668,N_3761);
and U7146 (N_7146,N_4148,N_3704);
or U7147 (N_7147,N_3128,N_4024);
and U7148 (N_7148,N_2332,N_3879);
and U7149 (N_7149,N_3482,N_3142);
or U7150 (N_7150,N_4740,N_3140);
nand U7151 (N_7151,N_1344,N_975);
or U7152 (N_7152,N_843,N_3961);
or U7153 (N_7153,N_2217,N_3495);
nand U7154 (N_7154,N_2140,N_1271);
and U7155 (N_7155,N_3232,N_4802);
and U7156 (N_7156,N_200,N_736);
and U7157 (N_7157,N_988,N_2423);
nor U7158 (N_7158,N_3212,N_1194);
nor U7159 (N_7159,N_4426,N_789);
and U7160 (N_7160,N_3955,N_884);
and U7161 (N_7161,N_2583,N_3554);
and U7162 (N_7162,N_2413,N_2686);
or U7163 (N_7163,N_2284,N_4077);
nand U7164 (N_7164,N_4185,N_1145);
nand U7165 (N_7165,N_2221,N_569);
nor U7166 (N_7166,N_953,N_2225);
nand U7167 (N_7167,N_2936,N_276);
or U7168 (N_7168,N_2390,N_2599);
or U7169 (N_7169,N_2460,N_1169);
or U7170 (N_7170,N_232,N_3327);
nor U7171 (N_7171,N_4069,N_2649);
nor U7172 (N_7172,N_2832,N_1396);
and U7173 (N_7173,N_1720,N_999);
or U7174 (N_7174,N_323,N_79);
or U7175 (N_7175,N_2109,N_3253);
nor U7176 (N_7176,N_662,N_931);
nand U7177 (N_7177,N_3578,N_1171);
nand U7178 (N_7178,N_1473,N_2811);
nand U7179 (N_7179,N_3071,N_1530);
nor U7180 (N_7180,N_3092,N_4820);
and U7181 (N_7181,N_3812,N_2294);
nand U7182 (N_7182,N_4920,N_4839);
nor U7183 (N_7183,N_3899,N_629);
nand U7184 (N_7184,N_2555,N_1384);
nor U7185 (N_7185,N_3513,N_2372);
nor U7186 (N_7186,N_1624,N_2212);
or U7187 (N_7187,N_2854,N_3687);
nand U7188 (N_7188,N_2131,N_56);
and U7189 (N_7189,N_2963,N_3259);
and U7190 (N_7190,N_2145,N_3430);
nor U7191 (N_7191,N_3508,N_2004);
nand U7192 (N_7192,N_399,N_2642);
and U7193 (N_7193,N_2389,N_3249);
and U7194 (N_7194,N_4743,N_745);
xor U7195 (N_7195,N_1585,N_1958);
and U7196 (N_7196,N_4308,N_1034);
and U7197 (N_7197,N_1272,N_4664);
and U7198 (N_7198,N_3530,N_314);
nor U7199 (N_7199,N_2793,N_4637);
nand U7200 (N_7200,N_1874,N_1526);
nor U7201 (N_7201,N_3489,N_3974);
nor U7202 (N_7202,N_1100,N_2213);
and U7203 (N_7203,N_2530,N_945);
nand U7204 (N_7204,N_239,N_2631);
and U7205 (N_7205,N_812,N_3298);
or U7206 (N_7206,N_2901,N_2849);
or U7207 (N_7207,N_2775,N_2808);
nor U7208 (N_7208,N_3243,N_964);
or U7209 (N_7209,N_2938,N_1560);
or U7210 (N_7210,N_371,N_929);
nand U7211 (N_7211,N_2982,N_2240);
nor U7212 (N_7212,N_2271,N_4931);
nand U7213 (N_7213,N_1960,N_3379);
and U7214 (N_7214,N_9,N_4347);
nand U7215 (N_7215,N_4198,N_4569);
xnor U7216 (N_7216,N_3725,N_1660);
nand U7217 (N_7217,N_2741,N_772);
and U7218 (N_7218,N_2342,N_4717);
and U7219 (N_7219,N_4961,N_4815);
or U7220 (N_7220,N_3810,N_227);
nor U7221 (N_7221,N_3802,N_4490);
nand U7222 (N_7222,N_2706,N_2169);
nor U7223 (N_7223,N_1024,N_672);
nand U7224 (N_7224,N_480,N_2214);
nor U7225 (N_7225,N_2542,N_4970);
and U7226 (N_7226,N_3672,N_4438);
nor U7227 (N_7227,N_1411,N_4564);
nor U7228 (N_7228,N_3898,N_1147);
nor U7229 (N_7229,N_1854,N_1628);
xnor U7230 (N_7230,N_225,N_288);
nor U7231 (N_7231,N_3157,N_4844);
nand U7232 (N_7232,N_441,N_91);
and U7233 (N_7233,N_3537,N_3044);
nor U7234 (N_7234,N_3139,N_4816);
nor U7235 (N_7235,N_4642,N_3766);
nand U7236 (N_7236,N_1789,N_2645);
nor U7237 (N_7237,N_4326,N_4702);
nor U7238 (N_7238,N_4016,N_728);
nor U7239 (N_7239,N_3395,N_1192);
and U7240 (N_7240,N_2075,N_2278);
nand U7241 (N_7241,N_1938,N_1115);
and U7242 (N_7242,N_219,N_3920);
or U7243 (N_7243,N_4533,N_3833);
or U7244 (N_7244,N_560,N_4576);
or U7245 (N_7245,N_2577,N_1814);
or U7246 (N_7246,N_2104,N_3406);
nor U7247 (N_7247,N_2473,N_2089);
nand U7248 (N_7248,N_941,N_2157);
nor U7249 (N_7249,N_4606,N_255);
and U7250 (N_7250,N_380,N_2708);
nand U7251 (N_7251,N_3645,N_4747);
or U7252 (N_7252,N_4622,N_2783);
nor U7253 (N_7253,N_704,N_4361);
or U7254 (N_7254,N_2718,N_4056);
or U7255 (N_7255,N_4383,N_4034);
nor U7256 (N_7256,N_3771,N_4009);
nor U7257 (N_7257,N_3234,N_4662);
nand U7258 (N_7258,N_2297,N_2012);
or U7259 (N_7259,N_1672,N_3552);
nand U7260 (N_7260,N_1134,N_2024);
nand U7261 (N_7261,N_1500,N_4305);
nand U7262 (N_7262,N_3152,N_2288);
or U7263 (N_7263,N_3192,N_2422);
or U7264 (N_7264,N_2155,N_3607);
and U7265 (N_7265,N_3470,N_4113);
and U7266 (N_7266,N_1709,N_294);
nor U7267 (N_7267,N_188,N_3600);
or U7268 (N_7268,N_943,N_2309);
or U7269 (N_7269,N_4345,N_4204);
and U7270 (N_7270,N_3937,N_1929);
or U7271 (N_7271,N_1047,N_562);
or U7272 (N_7272,N_4192,N_2769);
xor U7273 (N_7273,N_2787,N_1505);
nand U7274 (N_7274,N_1603,N_827);
nand U7275 (N_7275,N_4118,N_3863);
nor U7276 (N_7276,N_4300,N_4104);
nand U7277 (N_7277,N_1424,N_786);
nand U7278 (N_7278,N_1256,N_1236);
nor U7279 (N_7279,N_2474,N_2455);
nor U7280 (N_7280,N_4854,N_4805);
and U7281 (N_7281,N_1605,N_791);
or U7282 (N_7282,N_3108,N_4542);
and U7283 (N_7283,N_2037,N_1584);
and U7284 (N_7284,N_4266,N_3342);
or U7285 (N_7285,N_2376,N_168);
nor U7286 (N_7286,N_3266,N_12);
nor U7287 (N_7287,N_3392,N_1574);
and U7288 (N_7288,N_3499,N_3598);
or U7289 (N_7289,N_49,N_1888);
or U7290 (N_7290,N_613,N_1750);
or U7291 (N_7291,N_979,N_2857);
and U7292 (N_7292,N_1364,N_407);
and U7293 (N_7293,N_928,N_3177);
or U7294 (N_7294,N_4385,N_4763);
or U7295 (N_7295,N_2471,N_513);
nand U7296 (N_7296,N_2943,N_2900);
and U7297 (N_7297,N_3066,N_4245);
nand U7298 (N_7298,N_2688,N_2270);
and U7299 (N_7299,N_3073,N_3515);
or U7300 (N_7300,N_3176,N_4182);
and U7301 (N_7301,N_283,N_4251);
and U7302 (N_7302,N_3115,N_1721);
nor U7303 (N_7303,N_1050,N_3798);
nor U7304 (N_7304,N_3660,N_3394);
xor U7305 (N_7305,N_2869,N_3264);
or U7306 (N_7306,N_1139,N_3629);
nor U7307 (N_7307,N_3079,N_321);
nand U7308 (N_7308,N_2774,N_3311);
or U7309 (N_7309,N_703,N_1301);
nand U7310 (N_7310,N_3055,N_3914);
nor U7311 (N_7311,N_4567,N_2730);
nand U7312 (N_7312,N_3008,N_3101);
nor U7313 (N_7313,N_1053,N_2988);
or U7314 (N_7314,N_2705,N_4895);
and U7315 (N_7315,N_2273,N_2633);
and U7316 (N_7316,N_1437,N_2490);
nand U7317 (N_7317,N_1922,N_310);
nor U7318 (N_7318,N_4419,N_2928);
nand U7319 (N_7319,N_4556,N_2393);
nand U7320 (N_7320,N_36,N_331);
nand U7321 (N_7321,N_841,N_4771);
or U7322 (N_7322,N_2940,N_976);
nand U7323 (N_7323,N_4367,N_3186);
nand U7324 (N_7324,N_1016,N_3557);
and U7325 (N_7325,N_1952,N_970);
nor U7326 (N_7326,N_2847,N_620);
and U7327 (N_7327,N_3528,N_4631);
or U7328 (N_7328,N_3256,N_3714);
nor U7329 (N_7329,N_216,N_1323);
nor U7330 (N_7330,N_243,N_4064);
xor U7331 (N_7331,N_3857,N_2961);
nor U7332 (N_7332,N_1160,N_2699);
or U7333 (N_7333,N_4152,N_2840);
nand U7334 (N_7334,N_1155,N_4391);
or U7335 (N_7335,N_279,N_3382);
nand U7336 (N_7336,N_237,N_2764);
nor U7337 (N_7337,N_1763,N_1583);
nor U7338 (N_7338,N_3796,N_3133);
nand U7339 (N_7339,N_872,N_3563);
nor U7340 (N_7340,N_4984,N_1015);
and U7341 (N_7341,N_4918,N_2581);
and U7342 (N_7342,N_901,N_4797);
or U7343 (N_7343,N_2539,N_4955);
and U7344 (N_7344,N_1976,N_2143);
nor U7345 (N_7345,N_1376,N_4212);
or U7346 (N_7346,N_191,N_751);
nor U7347 (N_7347,N_4630,N_4870);
nand U7348 (N_7348,N_539,N_2242);
nand U7349 (N_7349,N_2560,N_2154);
or U7350 (N_7350,N_4700,N_1332);
nand U7351 (N_7351,N_4440,N_4083);
or U7352 (N_7352,N_4376,N_538);
and U7353 (N_7353,N_4618,N_4845);
nand U7354 (N_7354,N_2105,N_3527);
or U7355 (N_7355,N_1367,N_3012);
and U7356 (N_7356,N_3624,N_4110);
and U7357 (N_7357,N_1930,N_2608);
nor U7358 (N_7358,N_3052,N_1082);
or U7359 (N_7359,N_663,N_2059);
nor U7360 (N_7360,N_678,N_3627);
nor U7361 (N_7361,N_4683,N_3260);
or U7362 (N_7362,N_2871,N_4360);
nand U7363 (N_7363,N_3772,N_4246);
and U7364 (N_7364,N_3718,N_2954);
xnor U7365 (N_7365,N_661,N_1861);
and U7366 (N_7366,N_361,N_3559);
nand U7367 (N_7367,N_4410,N_2415);
or U7368 (N_7368,N_3500,N_4242);
nand U7369 (N_7369,N_2101,N_3247);
xnor U7370 (N_7370,N_2557,N_1118);
nand U7371 (N_7371,N_4635,N_3261);
nand U7372 (N_7372,N_1058,N_1033);
nor U7373 (N_7373,N_2759,N_1392);
and U7374 (N_7374,N_3679,N_3520);
or U7375 (N_7375,N_2794,N_2029);
and U7376 (N_7376,N_2185,N_293);
or U7377 (N_7377,N_2615,N_1433);
nand U7378 (N_7378,N_374,N_4108);
nand U7379 (N_7379,N_2585,N_1459);
nand U7380 (N_7380,N_1357,N_2200);
or U7381 (N_7381,N_3199,N_4114);
xor U7382 (N_7382,N_1061,N_2236);
or U7383 (N_7383,N_2523,N_3372);
and U7384 (N_7384,N_3331,N_4106);
nand U7385 (N_7385,N_1522,N_982);
nand U7386 (N_7386,N_2503,N_3621);
nand U7387 (N_7387,N_4035,N_2220);
nand U7388 (N_7388,N_2818,N_4947);
nor U7389 (N_7389,N_4885,N_93);
or U7390 (N_7390,N_4594,N_2182);
or U7391 (N_7391,N_690,N_4649);
nor U7392 (N_7392,N_2933,N_4336);
or U7393 (N_7393,N_1110,N_506);
xnor U7394 (N_7394,N_1048,N_1232);
nor U7395 (N_7395,N_1654,N_2937);
nor U7396 (N_7396,N_919,N_2136);
nand U7397 (N_7397,N_4596,N_4496);
and U7398 (N_7398,N_4670,N_1589);
nand U7399 (N_7399,N_2021,N_3890);
nor U7400 (N_7400,N_3059,N_935);
or U7401 (N_7401,N_4100,N_3021);
nand U7402 (N_7402,N_850,N_1200);
xnor U7403 (N_7403,N_4403,N_1876);
nand U7404 (N_7404,N_4186,N_734);
or U7405 (N_7405,N_2307,N_649);
nor U7406 (N_7406,N_4366,N_2749);
nor U7407 (N_7407,N_3782,N_370);
or U7408 (N_7408,N_3214,N_3680);
nand U7409 (N_7409,N_2370,N_2929);
and U7410 (N_7410,N_4512,N_3183);
nor U7411 (N_7411,N_3462,N_2067);
nor U7412 (N_7412,N_676,N_3290);
nand U7413 (N_7413,N_3789,N_26);
nor U7414 (N_7414,N_2955,N_611);
and U7415 (N_7415,N_2782,N_2047);
and U7416 (N_7416,N_1568,N_1439);
nand U7417 (N_7417,N_402,N_3925);
and U7418 (N_7418,N_2056,N_989);
nor U7419 (N_7419,N_2380,N_4758);
nor U7420 (N_7420,N_2796,N_1744);
nor U7421 (N_7421,N_4560,N_1280);
or U7422 (N_7422,N_1421,N_3859);
and U7423 (N_7423,N_4398,N_1170);
nor U7424 (N_7424,N_3280,N_4860);
and U7425 (N_7425,N_99,N_1948);
and U7426 (N_7426,N_1382,N_2898);
nor U7427 (N_7427,N_3216,N_373);
xnor U7428 (N_7428,N_4978,N_4053);
or U7429 (N_7429,N_4269,N_580);
and U7430 (N_7430,N_4677,N_3062);
or U7431 (N_7431,N_829,N_4312);
nor U7432 (N_7432,N_1616,N_1291);
and U7433 (N_7433,N_1829,N_4364);
nand U7434 (N_7434,N_4287,N_4244);
nand U7435 (N_7435,N_1044,N_1841);
xor U7436 (N_7436,N_3677,N_3933);
nor U7437 (N_7437,N_1790,N_4995);
or U7438 (N_7438,N_4568,N_750);
and U7439 (N_7439,N_1728,N_947);
and U7440 (N_7440,N_1446,N_4093);
nand U7441 (N_7441,N_3166,N_1516);
nand U7442 (N_7442,N_3864,N_1954);
or U7443 (N_7443,N_900,N_1640);
or U7444 (N_7444,N_3163,N_573);
nand U7445 (N_7445,N_1681,N_2192);
xor U7446 (N_7446,N_3756,N_542);
xnor U7447 (N_7447,N_754,N_4872);
and U7448 (N_7448,N_1626,N_4672);
nor U7449 (N_7449,N_820,N_3432);
nand U7450 (N_7450,N_4023,N_330);
and U7451 (N_7451,N_3417,N_770);
nand U7452 (N_7452,N_1884,N_4018);
nand U7453 (N_7453,N_2858,N_2431);
nor U7454 (N_7454,N_2246,N_2535);
or U7455 (N_7455,N_1193,N_3546);
or U7456 (N_7456,N_4965,N_4493);
or U7457 (N_7457,N_2310,N_3111);
and U7458 (N_7458,N_746,N_2896);
or U7459 (N_7459,N_4588,N_264);
nand U7460 (N_7460,N_3475,N_4236);
nor U7461 (N_7461,N_2944,N_2454);
or U7462 (N_7462,N_2498,N_4817);
nor U7463 (N_7463,N_2416,N_3153);
nand U7464 (N_7464,N_1146,N_1989);
or U7465 (N_7465,N_3787,N_2452);
or U7466 (N_7466,N_3043,N_3747);
nand U7467 (N_7467,N_1674,N_3158);
nor U7468 (N_7468,N_163,N_378);
and U7469 (N_7469,N_2826,N_3715);
nand U7470 (N_7470,N_3221,N_4983);
and U7471 (N_7471,N_3091,N_2095);
or U7472 (N_7472,N_4351,N_2252);
or U7473 (N_7473,N_4792,N_3285);
nor U7474 (N_7474,N_1576,N_522);
nand U7475 (N_7475,N_823,N_2679);
nand U7476 (N_7476,N_347,N_1228);
nor U7477 (N_7477,N_697,N_570);
and U7478 (N_7478,N_4521,N_1213);
xor U7479 (N_7479,N_1070,N_907);
nand U7480 (N_7480,N_3301,N_4675);
xor U7481 (N_7481,N_3154,N_4173);
or U7482 (N_7482,N_464,N_1610);
and U7483 (N_7483,N_3279,N_4121);
nor U7484 (N_7484,N_52,N_3195);
or U7485 (N_7485,N_4487,N_3795);
or U7486 (N_7486,N_241,N_1443);
and U7487 (N_7487,N_2042,N_4613);
or U7488 (N_7488,N_530,N_1023);
nor U7489 (N_7489,N_512,N_2249);
or U7490 (N_7490,N_3953,N_3359);
and U7491 (N_7491,N_2950,N_37);
nor U7492 (N_7492,N_2875,N_3870);
or U7493 (N_7493,N_3979,N_4252);
nor U7494 (N_7494,N_4503,N_3757);
nor U7495 (N_7495,N_916,N_4580);
nand U7496 (N_7496,N_210,N_4739);
nand U7497 (N_7497,N_3328,N_1697);
or U7498 (N_7498,N_4761,N_1401);
or U7499 (N_7499,N_1225,N_259);
nand U7500 (N_7500,N_4649,N_4992);
or U7501 (N_7501,N_2275,N_2021);
nor U7502 (N_7502,N_4384,N_4299);
nor U7503 (N_7503,N_3622,N_2005);
or U7504 (N_7504,N_946,N_1255);
nand U7505 (N_7505,N_2422,N_3041);
nand U7506 (N_7506,N_4026,N_3289);
nor U7507 (N_7507,N_1862,N_3604);
or U7508 (N_7508,N_3081,N_4115);
nor U7509 (N_7509,N_2033,N_1850);
and U7510 (N_7510,N_3660,N_3160);
or U7511 (N_7511,N_4591,N_4412);
and U7512 (N_7512,N_3138,N_3935);
xnor U7513 (N_7513,N_1566,N_2964);
nor U7514 (N_7514,N_221,N_3422);
and U7515 (N_7515,N_1202,N_4311);
and U7516 (N_7516,N_4666,N_4944);
and U7517 (N_7517,N_1765,N_3002);
or U7518 (N_7518,N_959,N_2398);
nor U7519 (N_7519,N_4779,N_1772);
or U7520 (N_7520,N_3575,N_345);
nand U7521 (N_7521,N_3971,N_1579);
nand U7522 (N_7522,N_4028,N_1504);
nor U7523 (N_7523,N_4422,N_4896);
or U7524 (N_7524,N_3519,N_2197);
or U7525 (N_7525,N_4188,N_3594);
or U7526 (N_7526,N_348,N_1258);
or U7527 (N_7527,N_1200,N_565);
nor U7528 (N_7528,N_365,N_95);
nor U7529 (N_7529,N_2156,N_1368);
nand U7530 (N_7530,N_1748,N_2121);
nand U7531 (N_7531,N_550,N_1556);
nor U7532 (N_7532,N_118,N_1088);
nor U7533 (N_7533,N_3665,N_4710);
or U7534 (N_7534,N_909,N_3374);
nor U7535 (N_7535,N_3523,N_4741);
and U7536 (N_7536,N_1623,N_195);
and U7537 (N_7537,N_4726,N_4820);
nor U7538 (N_7538,N_152,N_1086);
or U7539 (N_7539,N_2569,N_1969);
and U7540 (N_7540,N_1513,N_4375);
or U7541 (N_7541,N_152,N_1947);
and U7542 (N_7542,N_1205,N_4451);
and U7543 (N_7543,N_1157,N_4416);
nand U7544 (N_7544,N_3026,N_531);
nand U7545 (N_7545,N_4798,N_4763);
and U7546 (N_7546,N_499,N_277);
and U7547 (N_7547,N_1811,N_1512);
or U7548 (N_7548,N_2049,N_4149);
nor U7549 (N_7549,N_4712,N_3299);
nor U7550 (N_7550,N_2511,N_2053);
or U7551 (N_7551,N_829,N_3725);
nor U7552 (N_7552,N_619,N_4614);
nor U7553 (N_7553,N_4545,N_760);
nand U7554 (N_7554,N_4429,N_3835);
or U7555 (N_7555,N_1194,N_4509);
or U7556 (N_7556,N_3307,N_3472);
and U7557 (N_7557,N_2651,N_4366);
xnor U7558 (N_7558,N_4299,N_4065);
nor U7559 (N_7559,N_4154,N_162);
or U7560 (N_7560,N_3393,N_3333);
and U7561 (N_7561,N_1020,N_2135);
or U7562 (N_7562,N_3449,N_569);
xnor U7563 (N_7563,N_2832,N_154);
nand U7564 (N_7564,N_2408,N_1576);
nand U7565 (N_7565,N_727,N_2949);
and U7566 (N_7566,N_3312,N_3713);
and U7567 (N_7567,N_4613,N_1654);
and U7568 (N_7568,N_3778,N_1293);
nor U7569 (N_7569,N_4779,N_2341);
and U7570 (N_7570,N_4381,N_1704);
nor U7571 (N_7571,N_1367,N_3761);
and U7572 (N_7572,N_2789,N_354);
nor U7573 (N_7573,N_2812,N_2340);
nand U7574 (N_7574,N_941,N_1983);
or U7575 (N_7575,N_3086,N_915);
nor U7576 (N_7576,N_4584,N_2838);
nor U7577 (N_7577,N_3505,N_2042);
or U7578 (N_7578,N_218,N_1067);
or U7579 (N_7579,N_2618,N_3711);
nor U7580 (N_7580,N_3144,N_2133);
or U7581 (N_7581,N_2331,N_724);
nand U7582 (N_7582,N_2659,N_4122);
or U7583 (N_7583,N_237,N_2999);
nand U7584 (N_7584,N_3974,N_2815);
or U7585 (N_7585,N_1595,N_2501);
or U7586 (N_7586,N_679,N_2042);
and U7587 (N_7587,N_3098,N_4022);
nand U7588 (N_7588,N_1779,N_2198);
or U7589 (N_7589,N_4937,N_4923);
or U7590 (N_7590,N_2470,N_3140);
nand U7591 (N_7591,N_1271,N_4707);
nor U7592 (N_7592,N_1749,N_3180);
and U7593 (N_7593,N_3269,N_4327);
and U7594 (N_7594,N_3926,N_3214);
and U7595 (N_7595,N_3458,N_1763);
and U7596 (N_7596,N_3519,N_2107);
nand U7597 (N_7597,N_2619,N_4507);
or U7598 (N_7598,N_1701,N_2833);
nor U7599 (N_7599,N_4228,N_2468);
nor U7600 (N_7600,N_3164,N_2366);
nor U7601 (N_7601,N_3353,N_4351);
nor U7602 (N_7602,N_3988,N_776);
nand U7603 (N_7603,N_3495,N_2064);
or U7604 (N_7604,N_1404,N_3894);
nor U7605 (N_7605,N_1849,N_3869);
or U7606 (N_7606,N_1143,N_2557);
or U7607 (N_7607,N_2458,N_1491);
or U7608 (N_7608,N_4671,N_3386);
or U7609 (N_7609,N_4374,N_945);
nor U7610 (N_7610,N_1286,N_332);
nand U7611 (N_7611,N_4206,N_2765);
nand U7612 (N_7612,N_4756,N_1663);
nand U7613 (N_7613,N_2054,N_943);
and U7614 (N_7614,N_3726,N_3975);
or U7615 (N_7615,N_2356,N_2841);
and U7616 (N_7616,N_1869,N_2101);
nand U7617 (N_7617,N_4539,N_591);
and U7618 (N_7618,N_373,N_2859);
nor U7619 (N_7619,N_3459,N_2974);
or U7620 (N_7620,N_2179,N_3241);
nor U7621 (N_7621,N_3237,N_4172);
nand U7622 (N_7622,N_2755,N_1144);
nand U7623 (N_7623,N_1028,N_1284);
and U7624 (N_7624,N_4271,N_1772);
and U7625 (N_7625,N_542,N_2922);
nor U7626 (N_7626,N_4630,N_3938);
or U7627 (N_7627,N_1199,N_866);
nor U7628 (N_7628,N_4872,N_3400);
nor U7629 (N_7629,N_1410,N_3141);
and U7630 (N_7630,N_2841,N_1485);
or U7631 (N_7631,N_428,N_1337);
or U7632 (N_7632,N_596,N_458);
nor U7633 (N_7633,N_1422,N_4445);
nor U7634 (N_7634,N_1678,N_2039);
nand U7635 (N_7635,N_4517,N_3855);
and U7636 (N_7636,N_4516,N_4277);
or U7637 (N_7637,N_4181,N_4404);
nand U7638 (N_7638,N_1156,N_4561);
nor U7639 (N_7639,N_3611,N_1685);
and U7640 (N_7640,N_3642,N_1032);
nand U7641 (N_7641,N_3512,N_3096);
and U7642 (N_7642,N_796,N_3680);
and U7643 (N_7643,N_2820,N_4318);
or U7644 (N_7644,N_476,N_4927);
nand U7645 (N_7645,N_3947,N_3695);
and U7646 (N_7646,N_2824,N_2479);
nor U7647 (N_7647,N_829,N_4345);
and U7648 (N_7648,N_1034,N_1320);
nor U7649 (N_7649,N_1199,N_3525);
or U7650 (N_7650,N_4579,N_415);
and U7651 (N_7651,N_448,N_2006);
and U7652 (N_7652,N_2850,N_4827);
or U7653 (N_7653,N_1624,N_272);
nor U7654 (N_7654,N_3166,N_4705);
and U7655 (N_7655,N_360,N_3598);
xor U7656 (N_7656,N_4523,N_1248);
and U7657 (N_7657,N_661,N_147);
nor U7658 (N_7658,N_2385,N_1437);
and U7659 (N_7659,N_689,N_3958);
and U7660 (N_7660,N_4851,N_3312);
and U7661 (N_7661,N_141,N_4919);
nand U7662 (N_7662,N_4147,N_3129);
nand U7663 (N_7663,N_2372,N_1187);
nor U7664 (N_7664,N_2459,N_2523);
nor U7665 (N_7665,N_3991,N_2753);
nor U7666 (N_7666,N_4232,N_1008);
and U7667 (N_7667,N_3596,N_1850);
and U7668 (N_7668,N_4057,N_1098);
nand U7669 (N_7669,N_458,N_1185);
and U7670 (N_7670,N_4478,N_578);
nand U7671 (N_7671,N_733,N_4746);
nand U7672 (N_7672,N_2739,N_229);
and U7673 (N_7673,N_2372,N_2551);
nor U7674 (N_7674,N_1351,N_3857);
or U7675 (N_7675,N_499,N_2177);
xnor U7676 (N_7676,N_1572,N_1931);
nand U7677 (N_7677,N_3679,N_3667);
or U7678 (N_7678,N_4380,N_3557);
and U7679 (N_7679,N_2018,N_954);
nand U7680 (N_7680,N_2149,N_3613);
and U7681 (N_7681,N_3978,N_3141);
nor U7682 (N_7682,N_3535,N_404);
nor U7683 (N_7683,N_1743,N_1641);
or U7684 (N_7684,N_1815,N_2837);
and U7685 (N_7685,N_3202,N_4114);
and U7686 (N_7686,N_2796,N_84);
xor U7687 (N_7687,N_4112,N_3374);
nor U7688 (N_7688,N_1125,N_3615);
nor U7689 (N_7689,N_1671,N_4100);
nand U7690 (N_7690,N_673,N_1948);
nand U7691 (N_7691,N_2398,N_3568);
nor U7692 (N_7692,N_4727,N_3082);
or U7693 (N_7693,N_2895,N_4024);
nor U7694 (N_7694,N_1378,N_4465);
or U7695 (N_7695,N_2041,N_3266);
nand U7696 (N_7696,N_641,N_1097);
nand U7697 (N_7697,N_4440,N_3895);
or U7698 (N_7698,N_4940,N_2684);
or U7699 (N_7699,N_396,N_341);
nor U7700 (N_7700,N_2360,N_1299);
or U7701 (N_7701,N_3711,N_3520);
and U7702 (N_7702,N_920,N_2586);
nor U7703 (N_7703,N_2878,N_4285);
nand U7704 (N_7704,N_3980,N_317);
nand U7705 (N_7705,N_2525,N_2267);
and U7706 (N_7706,N_1292,N_661);
nand U7707 (N_7707,N_844,N_2269);
and U7708 (N_7708,N_3501,N_3803);
nand U7709 (N_7709,N_1979,N_2864);
or U7710 (N_7710,N_4205,N_3539);
nand U7711 (N_7711,N_4309,N_3106);
nor U7712 (N_7712,N_1656,N_3695);
nand U7713 (N_7713,N_2539,N_1777);
and U7714 (N_7714,N_2095,N_1137);
nand U7715 (N_7715,N_3756,N_4131);
nand U7716 (N_7716,N_4946,N_3093);
nor U7717 (N_7717,N_1059,N_4199);
and U7718 (N_7718,N_415,N_1108);
nand U7719 (N_7719,N_2219,N_3302);
and U7720 (N_7720,N_2113,N_3468);
nor U7721 (N_7721,N_2131,N_3874);
or U7722 (N_7722,N_1005,N_3312);
nand U7723 (N_7723,N_4873,N_2097);
and U7724 (N_7724,N_3661,N_4822);
or U7725 (N_7725,N_3804,N_1146);
or U7726 (N_7726,N_1236,N_4181);
nor U7727 (N_7727,N_3693,N_4456);
nand U7728 (N_7728,N_2571,N_1097);
nor U7729 (N_7729,N_2020,N_2683);
or U7730 (N_7730,N_3798,N_4147);
nor U7731 (N_7731,N_2150,N_4217);
and U7732 (N_7732,N_2648,N_2402);
nor U7733 (N_7733,N_3085,N_287);
and U7734 (N_7734,N_1215,N_1072);
nor U7735 (N_7735,N_3119,N_349);
or U7736 (N_7736,N_2048,N_1622);
nor U7737 (N_7737,N_1110,N_4633);
nand U7738 (N_7738,N_3681,N_1005);
nand U7739 (N_7739,N_4732,N_4673);
nand U7740 (N_7740,N_921,N_419);
and U7741 (N_7741,N_1173,N_4489);
and U7742 (N_7742,N_3339,N_1146);
or U7743 (N_7743,N_927,N_652);
nor U7744 (N_7744,N_3391,N_1346);
nor U7745 (N_7745,N_2721,N_1096);
or U7746 (N_7746,N_2006,N_2253);
or U7747 (N_7747,N_2867,N_1339);
nand U7748 (N_7748,N_1361,N_2165);
nand U7749 (N_7749,N_1865,N_2893);
nor U7750 (N_7750,N_1309,N_52);
xnor U7751 (N_7751,N_4302,N_3573);
or U7752 (N_7752,N_2619,N_742);
and U7753 (N_7753,N_1542,N_3289);
nor U7754 (N_7754,N_3996,N_2275);
nand U7755 (N_7755,N_3863,N_4652);
nor U7756 (N_7756,N_4309,N_49);
and U7757 (N_7757,N_3575,N_1475);
nand U7758 (N_7758,N_1905,N_1832);
and U7759 (N_7759,N_4753,N_3206);
or U7760 (N_7760,N_1388,N_3827);
nor U7761 (N_7761,N_2369,N_4699);
or U7762 (N_7762,N_760,N_442);
and U7763 (N_7763,N_1626,N_1231);
and U7764 (N_7764,N_4460,N_4070);
xnor U7765 (N_7765,N_537,N_930);
or U7766 (N_7766,N_1482,N_4994);
nand U7767 (N_7767,N_581,N_1956);
nor U7768 (N_7768,N_1085,N_4991);
and U7769 (N_7769,N_2247,N_776);
or U7770 (N_7770,N_1931,N_991);
or U7771 (N_7771,N_4916,N_4210);
and U7772 (N_7772,N_4619,N_2508);
nand U7773 (N_7773,N_2894,N_4337);
nand U7774 (N_7774,N_2088,N_3013);
nand U7775 (N_7775,N_3579,N_3853);
or U7776 (N_7776,N_307,N_2529);
and U7777 (N_7777,N_4157,N_2615);
xnor U7778 (N_7778,N_3889,N_565);
nand U7779 (N_7779,N_1620,N_3523);
nor U7780 (N_7780,N_1949,N_4747);
nand U7781 (N_7781,N_865,N_653);
and U7782 (N_7782,N_3634,N_2408);
nor U7783 (N_7783,N_2594,N_3048);
or U7784 (N_7784,N_2478,N_1754);
and U7785 (N_7785,N_4479,N_1755);
nor U7786 (N_7786,N_990,N_2036);
nor U7787 (N_7787,N_3866,N_1313);
nand U7788 (N_7788,N_269,N_3208);
nor U7789 (N_7789,N_4675,N_3609);
or U7790 (N_7790,N_3312,N_3958);
nand U7791 (N_7791,N_4944,N_499);
and U7792 (N_7792,N_3753,N_1232);
nand U7793 (N_7793,N_1364,N_2805);
or U7794 (N_7794,N_2027,N_4955);
nand U7795 (N_7795,N_3040,N_3959);
nand U7796 (N_7796,N_2460,N_997);
or U7797 (N_7797,N_4802,N_1871);
or U7798 (N_7798,N_2896,N_3883);
or U7799 (N_7799,N_2721,N_1032);
nand U7800 (N_7800,N_4978,N_510);
nand U7801 (N_7801,N_4547,N_2657);
nor U7802 (N_7802,N_3401,N_3944);
nand U7803 (N_7803,N_1213,N_1597);
nor U7804 (N_7804,N_4961,N_1055);
nor U7805 (N_7805,N_3812,N_1961);
and U7806 (N_7806,N_3444,N_3911);
nand U7807 (N_7807,N_2632,N_4837);
xnor U7808 (N_7808,N_151,N_4657);
or U7809 (N_7809,N_1149,N_2182);
nor U7810 (N_7810,N_2765,N_2198);
nor U7811 (N_7811,N_3026,N_655);
and U7812 (N_7812,N_4841,N_4568);
nand U7813 (N_7813,N_2727,N_3795);
nor U7814 (N_7814,N_4185,N_959);
and U7815 (N_7815,N_2144,N_2906);
or U7816 (N_7816,N_4766,N_3035);
xor U7817 (N_7817,N_1249,N_1417);
nand U7818 (N_7818,N_2783,N_330);
and U7819 (N_7819,N_3526,N_2096);
or U7820 (N_7820,N_501,N_2058);
or U7821 (N_7821,N_531,N_629);
and U7822 (N_7822,N_3012,N_127);
or U7823 (N_7823,N_4345,N_960);
or U7824 (N_7824,N_2902,N_193);
and U7825 (N_7825,N_3974,N_2010);
and U7826 (N_7826,N_1489,N_4033);
or U7827 (N_7827,N_903,N_1901);
or U7828 (N_7828,N_1415,N_1868);
and U7829 (N_7829,N_1342,N_1476);
nand U7830 (N_7830,N_525,N_4414);
nor U7831 (N_7831,N_3558,N_1784);
nand U7832 (N_7832,N_1480,N_3196);
nand U7833 (N_7833,N_2367,N_3173);
nand U7834 (N_7834,N_3991,N_374);
nand U7835 (N_7835,N_189,N_3482);
nand U7836 (N_7836,N_2015,N_3711);
nor U7837 (N_7837,N_4152,N_904);
or U7838 (N_7838,N_1003,N_1665);
and U7839 (N_7839,N_4611,N_4311);
nor U7840 (N_7840,N_3878,N_1483);
nand U7841 (N_7841,N_1098,N_350);
nand U7842 (N_7842,N_3121,N_2736);
and U7843 (N_7843,N_3380,N_1995);
nand U7844 (N_7844,N_1874,N_2754);
nand U7845 (N_7845,N_1685,N_3344);
or U7846 (N_7846,N_884,N_2572);
nand U7847 (N_7847,N_925,N_692);
or U7848 (N_7848,N_1278,N_3312);
xor U7849 (N_7849,N_4333,N_1407);
and U7850 (N_7850,N_2716,N_2489);
nand U7851 (N_7851,N_2742,N_3403);
or U7852 (N_7852,N_2987,N_3989);
nor U7853 (N_7853,N_955,N_4769);
nor U7854 (N_7854,N_3442,N_4133);
nor U7855 (N_7855,N_3153,N_4753);
or U7856 (N_7856,N_1395,N_3976);
nand U7857 (N_7857,N_1687,N_930);
and U7858 (N_7858,N_3268,N_3935);
nor U7859 (N_7859,N_897,N_1190);
nand U7860 (N_7860,N_1856,N_2602);
xor U7861 (N_7861,N_1643,N_2703);
nand U7862 (N_7862,N_1292,N_3815);
nor U7863 (N_7863,N_838,N_1775);
nand U7864 (N_7864,N_984,N_1174);
nand U7865 (N_7865,N_3040,N_2528);
xnor U7866 (N_7866,N_2410,N_569);
or U7867 (N_7867,N_899,N_2354);
nor U7868 (N_7868,N_690,N_3390);
nor U7869 (N_7869,N_3349,N_978);
or U7870 (N_7870,N_100,N_628);
or U7871 (N_7871,N_4628,N_2816);
or U7872 (N_7872,N_3228,N_3969);
nand U7873 (N_7873,N_3559,N_409);
and U7874 (N_7874,N_1612,N_2901);
and U7875 (N_7875,N_246,N_74);
nor U7876 (N_7876,N_2087,N_1443);
or U7877 (N_7877,N_3611,N_2177);
or U7878 (N_7878,N_4763,N_4196);
nor U7879 (N_7879,N_2950,N_4928);
nor U7880 (N_7880,N_3269,N_248);
nand U7881 (N_7881,N_657,N_1183);
nand U7882 (N_7882,N_3204,N_1301);
and U7883 (N_7883,N_967,N_1431);
nor U7884 (N_7884,N_1823,N_2226);
or U7885 (N_7885,N_2401,N_1751);
and U7886 (N_7886,N_1286,N_2088);
nor U7887 (N_7887,N_2779,N_3340);
nor U7888 (N_7888,N_3997,N_417);
nor U7889 (N_7889,N_2990,N_1195);
nand U7890 (N_7890,N_2316,N_4218);
or U7891 (N_7891,N_83,N_3926);
and U7892 (N_7892,N_2345,N_687);
or U7893 (N_7893,N_1679,N_568);
and U7894 (N_7894,N_1920,N_494);
nand U7895 (N_7895,N_4181,N_2997);
nor U7896 (N_7896,N_4952,N_2798);
nor U7897 (N_7897,N_2298,N_227);
nand U7898 (N_7898,N_4369,N_3668);
nand U7899 (N_7899,N_187,N_558);
nand U7900 (N_7900,N_2848,N_3561);
and U7901 (N_7901,N_980,N_3564);
nor U7902 (N_7902,N_1099,N_1586);
nand U7903 (N_7903,N_2110,N_2599);
and U7904 (N_7904,N_1855,N_3473);
nor U7905 (N_7905,N_1203,N_1575);
nor U7906 (N_7906,N_2576,N_2736);
nand U7907 (N_7907,N_6,N_427);
nor U7908 (N_7908,N_4869,N_4121);
or U7909 (N_7909,N_1109,N_4081);
or U7910 (N_7910,N_3942,N_820);
nor U7911 (N_7911,N_2731,N_674);
nor U7912 (N_7912,N_3145,N_4989);
nand U7913 (N_7913,N_3319,N_3978);
and U7914 (N_7914,N_2935,N_4064);
nand U7915 (N_7915,N_398,N_1017);
or U7916 (N_7916,N_115,N_1700);
nand U7917 (N_7917,N_312,N_863);
and U7918 (N_7918,N_2616,N_3061);
nor U7919 (N_7919,N_785,N_4669);
or U7920 (N_7920,N_1229,N_900);
nor U7921 (N_7921,N_3323,N_4484);
and U7922 (N_7922,N_2319,N_946);
or U7923 (N_7923,N_1467,N_1589);
nand U7924 (N_7924,N_3470,N_4308);
nand U7925 (N_7925,N_2013,N_1289);
nor U7926 (N_7926,N_1779,N_1541);
nor U7927 (N_7927,N_1040,N_1744);
xnor U7928 (N_7928,N_2885,N_2344);
or U7929 (N_7929,N_3197,N_188);
nor U7930 (N_7930,N_4978,N_4277);
nand U7931 (N_7931,N_2538,N_4106);
and U7932 (N_7932,N_3451,N_2682);
nand U7933 (N_7933,N_4851,N_175);
nand U7934 (N_7934,N_3778,N_2819);
nor U7935 (N_7935,N_3659,N_4178);
nor U7936 (N_7936,N_583,N_3334);
and U7937 (N_7937,N_1825,N_2078);
and U7938 (N_7938,N_2715,N_4480);
and U7939 (N_7939,N_4891,N_442);
or U7940 (N_7940,N_2659,N_817);
nor U7941 (N_7941,N_3177,N_4043);
and U7942 (N_7942,N_2816,N_468);
and U7943 (N_7943,N_3313,N_1441);
and U7944 (N_7944,N_2211,N_1357);
and U7945 (N_7945,N_1665,N_138);
nor U7946 (N_7946,N_4452,N_4795);
nor U7947 (N_7947,N_889,N_973);
or U7948 (N_7948,N_1291,N_3397);
nor U7949 (N_7949,N_4021,N_2055);
and U7950 (N_7950,N_4189,N_2303);
or U7951 (N_7951,N_1892,N_1698);
or U7952 (N_7952,N_774,N_4285);
or U7953 (N_7953,N_3875,N_1241);
nor U7954 (N_7954,N_1873,N_2820);
or U7955 (N_7955,N_2373,N_2050);
nand U7956 (N_7956,N_1303,N_148);
nand U7957 (N_7957,N_412,N_2370);
and U7958 (N_7958,N_598,N_3149);
nand U7959 (N_7959,N_4272,N_2875);
or U7960 (N_7960,N_1679,N_1396);
nand U7961 (N_7961,N_4314,N_2749);
nand U7962 (N_7962,N_2902,N_66);
nor U7963 (N_7963,N_4471,N_4170);
or U7964 (N_7964,N_685,N_1990);
nor U7965 (N_7965,N_555,N_709);
and U7966 (N_7966,N_4069,N_1901);
and U7967 (N_7967,N_1239,N_3939);
nor U7968 (N_7968,N_1432,N_2776);
or U7969 (N_7969,N_3688,N_2287);
nand U7970 (N_7970,N_2062,N_3480);
and U7971 (N_7971,N_2198,N_743);
or U7972 (N_7972,N_2092,N_3830);
nand U7973 (N_7973,N_3450,N_148);
and U7974 (N_7974,N_88,N_967);
or U7975 (N_7975,N_399,N_4966);
or U7976 (N_7976,N_1384,N_4341);
nand U7977 (N_7977,N_1033,N_3953);
or U7978 (N_7978,N_4138,N_4949);
and U7979 (N_7979,N_3385,N_2048);
nor U7980 (N_7980,N_4545,N_764);
or U7981 (N_7981,N_1072,N_2554);
and U7982 (N_7982,N_91,N_1813);
nor U7983 (N_7983,N_2668,N_3379);
nor U7984 (N_7984,N_4871,N_2811);
or U7985 (N_7985,N_2925,N_3664);
nand U7986 (N_7986,N_1478,N_3510);
nor U7987 (N_7987,N_3737,N_4744);
xnor U7988 (N_7988,N_694,N_3406);
and U7989 (N_7989,N_2305,N_4301);
nor U7990 (N_7990,N_4961,N_3547);
nand U7991 (N_7991,N_4124,N_301);
nor U7992 (N_7992,N_3561,N_2903);
nand U7993 (N_7993,N_4480,N_265);
nand U7994 (N_7994,N_1318,N_1897);
nor U7995 (N_7995,N_2925,N_1632);
or U7996 (N_7996,N_1075,N_250);
nand U7997 (N_7997,N_3640,N_1190);
and U7998 (N_7998,N_4904,N_4768);
nor U7999 (N_7999,N_4390,N_4167);
and U8000 (N_8000,N_4545,N_2597);
nor U8001 (N_8001,N_81,N_2004);
nand U8002 (N_8002,N_2260,N_3116);
nand U8003 (N_8003,N_2806,N_4123);
and U8004 (N_8004,N_1097,N_4190);
and U8005 (N_8005,N_635,N_3559);
nand U8006 (N_8006,N_2723,N_1723);
nor U8007 (N_8007,N_153,N_2662);
or U8008 (N_8008,N_2797,N_4814);
xnor U8009 (N_8009,N_4741,N_3079);
nor U8010 (N_8010,N_52,N_1171);
or U8011 (N_8011,N_308,N_1224);
or U8012 (N_8012,N_1128,N_4929);
nor U8013 (N_8013,N_1178,N_404);
or U8014 (N_8014,N_1506,N_1858);
and U8015 (N_8015,N_2540,N_1921);
nand U8016 (N_8016,N_2900,N_3471);
nand U8017 (N_8017,N_367,N_425);
and U8018 (N_8018,N_383,N_3340);
or U8019 (N_8019,N_292,N_3883);
nand U8020 (N_8020,N_1434,N_3029);
nor U8021 (N_8021,N_4544,N_1607);
nor U8022 (N_8022,N_4947,N_4442);
and U8023 (N_8023,N_787,N_1646);
or U8024 (N_8024,N_2863,N_2242);
or U8025 (N_8025,N_2930,N_620);
nor U8026 (N_8026,N_1735,N_1194);
and U8027 (N_8027,N_2426,N_181);
nor U8028 (N_8028,N_3638,N_4923);
or U8029 (N_8029,N_4858,N_3519);
or U8030 (N_8030,N_498,N_3568);
and U8031 (N_8031,N_1283,N_1503);
and U8032 (N_8032,N_2760,N_4396);
nand U8033 (N_8033,N_3893,N_4888);
nand U8034 (N_8034,N_1490,N_2294);
and U8035 (N_8035,N_2517,N_1594);
or U8036 (N_8036,N_2106,N_2477);
nor U8037 (N_8037,N_918,N_2588);
and U8038 (N_8038,N_421,N_4460);
nand U8039 (N_8039,N_2159,N_3608);
and U8040 (N_8040,N_4829,N_2883);
nor U8041 (N_8041,N_500,N_2276);
or U8042 (N_8042,N_2258,N_4396);
and U8043 (N_8043,N_2505,N_4060);
or U8044 (N_8044,N_4148,N_3039);
and U8045 (N_8045,N_3841,N_3337);
or U8046 (N_8046,N_3784,N_4783);
and U8047 (N_8047,N_3808,N_1892);
nand U8048 (N_8048,N_792,N_1584);
and U8049 (N_8049,N_558,N_626);
nor U8050 (N_8050,N_2508,N_3623);
or U8051 (N_8051,N_3315,N_3143);
and U8052 (N_8052,N_3933,N_3575);
nor U8053 (N_8053,N_1162,N_2084);
nor U8054 (N_8054,N_2991,N_3950);
nor U8055 (N_8055,N_2868,N_1333);
or U8056 (N_8056,N_4528,N_4185);
nor U8057 (N_8057,N_1550,N_1589);
nor U8058 (N_8058,N_2304,N_3216);
nand U8059 (N_8059,N_4657,N_3175);
and U8060 (N_8060,N_3978,N_3168);
nand U8061 (N_8061,N_3906,N_4196);
nand U8062 (N_8062,N_1039,N_2280);
nand U8063 (N_8063,N_3815,N_3755);
nand U8064 (N_8064,N_4579,N_236);
nand U8065 (N_8065,N_4323,N_2339);
and U8066 (N_8066,N_3529,N_2525);
and U8067 (N_8067,N_3961,N_144);
or U8068 (N_8068,N_405,N_647);
nand U8069 (N_8069,N_423,N_2045);
and U8070 (N_8070,N_4402,N_1087);
or U8071 (N_8071,N_1698,N_2244);
nand U8072 (N_8072,N_1192,N_2574);
and U8073 (N_8073,N_3060,N_1223);
nand U8074 (N_8074,N_3865,N_4495);
and U8075 (N_8075,N_1684,N_1738);
or U8076 (N_8076,N_1705,N_2100);
nand U8077 (N_8077,N_4038,N_2454);
or U8078 (N_8078,N_1295,N_3905);
nand U8079 (N_8079,N_135,N_4514);
and U8080 (N_8080,N_2571,N_2754);
nor U8081 (N_8081,N_586,N_2219);
nand U8082 (N_8082,N_426,N_4940);
nand U8083 (N_8083,N_3997,N_4189);
and U8084 (N_8084,N_3658,N_3718);
and U8085 (N_8085,N_2122,N_3336);
nor U8086 (N_8086,N_4256,N_4493);
nor U8087 (N_8087,N_4100,N_4274);
nand U8088 (N_8088,N_3748,N_3146);
and U8089 (N_8089,N_3473,N_3365);
nand U8090 (N_8090,N_3061,N_1206);
or U8091 (N_8091,N_3422,N_1828);
nand U8092 (N_8092,N_3320,N_656);
and U8093 (N_8093,N_3760,N_3631);
nor U8094 (N_8094,N_578,N_4503);
nor U8095 (N_8095,N_958,N_3529);
nand U8096 (N_8096,N_4909,N_2865);
nand U8097 (N_8097,N_4311,N_741);
nor U8098 (N_8098,N_2089,N_4089);
and U8099 (N_8099,N_4864,N_319);
and U8100 (N_8100,N_3811,N_935);
nor U8101 (N_8101,N_1922,N_126);
nand U8102 (N_8102,N_302,N_257);
and U8103 (N_8103,N_4905,N_3594);
nand U8104 (N_8104,N_45,N_306);
or U8105 (N_8105,N_2911,N_1855);
nor U8106 (N_8106,N_2987,N_3195);
and U8107 (N_8107,N_820,N_1019);
nor U8108 (N_8108,N_4924,N_462);
or U8109 (N_8109,N_2850,N_873);
nor U8110 (N_8110,N_3802,N_203);
nand U8111 (N_8111,N_3442,N_1551);
xnor U8112 (N_8112,N_3766,N_487);
and U8113 (N_8113,N_4269,N_2107);
or U8114 (N_8114,N_370,N_964);
nand U8115 (N_8115,N_2192,N_4747);
or U8116 (N_8116,N_3576,N_4481);
or U8117 (N_8117,N_4285,N_2485);
nand U8118 (N_8118,N_1566,N_2429);
nand U8119 (N_8119,N_553,N_4605);
nand U8120 (N_8120,N_3846,N_1999);
nand U8121 (N_8121,N_3989,N_2116);
nor U8122 (N_8122,N_3345,N_3340);
or U8123 (N_8123,N_3419,N_796);
or U8124 (N_8124,N_3735,N_2247);
or U8125 (N_8125,N_456,N_521);
and U8126 (N_8126,N_2151,N_4188);
and U8127 (N_8127,N_2889,N_3015);
nor U8128 (N_8128,N_4118,N_768);
and U8129 (N_8129,N_313,N_3160);
and U8130 (N_8130,N_4020,N_844);
and U8131 (N_8131,N_949,N_3048);
and U8132 (N_8132,N_472,N_202);
and U8133 (N_8133,N_3033,N_4586);
and U8134 (N_8134,N_1158,N_2298);
or U8135 (N_8135,N_3089,N_1009);
nor U8136 (N_8136,N_1645,N_1563);
nand U8137 (N_8137,N_3137,N_330);
and U8138 (N_8138,N_3764,N_1042);
and U8139 (N_8139,N_3581,N_1486);
and U8140 (N_8140,N_3531,N_4252);
or U8141 (N_8141,N_587,N_4614);
and U8142 (N_8142,N_4448,N_2898);
nand U8143 (N_8143,N_2639,N_3142);
nor U8144 (N_8144,N_3068,N_321);
and U8145 (N_8145,N_3336,N_285);
nand U8146 (N_8146,N_1260,N_3450);
or U8147 (N_8147,N_3482,N_1706);
and U8148 (N_8148,N_4480,N_4590);
nor U8149 (N_8149,N_1484,N_4399);
nor U8150 (N_8150,N_4490,N_1486);
or U8151 (N_8151,N_4232,N_4235);
and U8152 (N_8152,N_2650,N_4515);
and U8153 (N_8153,N_1506,N_3704);
nand U8154 (N_8154,N_357,N_4309);
nor U8155 (N_8155,N_1446,N_3822);
xor U8156 (N_8156,N_590,N_1128);
and U8157 (N_8157,N_3069,N_903);
nand U8158 (N_8158,N_2403,N_1464);
or U8159 (N_8159,N_2677,N_451);
nand U8160 (N_8160,N_3591,N_4979);
nor U8161 (N_8161,N_2631,N_684);
nor U8162 (N_8162,N_3179,N_3351);
or U8163 (N_8163,N_3045,N_1968);
nand U8164 (N_8164,N_1895,N_2867);
and U8165 (N_8165,N_4500,N_2437);
nor U8166 (N_8166,N_2302,N_2403);
and U8167 (N_8167,N_4605,N_365);
or U8168 (N_8168,N_2184,N_4380);
or U8169 (N_8169,N_2149,N_2085);
nand U8170 (N_8170,N_550,N_2349);
nor U8171 (N_8171,N_1596,N_735);
nand U8172 (N_8172,N_243,N_3434);
and U8173 (N_8173,N_2650,N_3520);
nor U8174 (N_8174,N_4229,N_2120);
nand U8175 (N_8175,N_3804,N_4496);
nor U8176 (N_8176,N_1063,N_4283);
nor U8177 (N_8177,N_4114,N_135);
and U8178 (N_8178,N_1003,N_4075);
xnor U8179 (N_8179,N_2111,N_1475);
nor U8180 (N_8180,N_1101,N_2345);
or U8181 (N_8181,N_724,N_1340);
and U8182 (N_8182,N_770,N_4292);
nor U8183 (N_8183,N_2620,N_4246);
nor U8184 (N_8184,N_3756,N_3022);
and U8185 (N_8185,N_4643,N_3964);
and U8186 (N_8186,N_4321,N_1995);
nor U8187 (N_8187,N_2493,N_4830);
nor U8188 (N_8188,N_1465,N_2331);
and U8189 (N_8189,N_2513,N_2444);
or U8190 (N_8190,N_1257,N_469);
or U8191 (N_8191,N_3021,N_3817);
and U8192 (N_8192,N_1075,N_1782);
nand U8193 (N_8193,N_1428,N_4025);
and U8194 (N_8194,N_2759,N_3104);
or U8195 (N_8195,N_2963,N_3337);
nor U8196 (N_8196,N_3698,N_544);
nand U8197 (N_8197,N_59,N_2393);
or U8198 (N_8198,N_1212,N_13);
nor U8199 (N_8199,N_3087,N_928);
and U8200 (N_8200,N_70,N_4079);
nor U8201 (N_8201,N_3328,N_3234);
or U8202 (N_8202,N_434,N_3751);
nor U8203 (N_8203,N_795,N_4536);
and U8204 (N_8204,N_1890,N_3663);
nor U8205 (N_8205,N_51,N_4571);
and U8206 (N_8206,N_429,N_337);
nand U8207 (N_8207,N_4715,N_4903);
nor U8208 (N_8208,N_3089,N_1407);
nor U8209 (N_8209,N_4789,N_1432);
xnor U8210 (N_8210,N_241,N_3734);
nor U8211 (N_8211,N_682,N_1690);
nor U8212 (N_8212,N_576,N_2940);
or U8213 (N_8213,N_1483,N_1925);
or U8214 (N_8214,N_930,N_4246);
and U8215 (N_8215,N_586,N_2178);
nand U8216 (N_8216,N_2025,N_1918);
nor U8217 (N_8217,N_1266,N_586);
or U8218 (N_8218,N_1777,N_3993);
and U8219 (N_8219,N_3704,N_4697);
or U8220 (N_8220,N_2979,N_1311);
nor U8221 (N_8221,N_4311,N_568);
nand U8222 (N_8222,N_3962,N_3151);
and U8223 (N_8223,N_3549,N_3344);
or U8224 (N_8224,N_2678,N_516);
nor U8225 (N_8225,N_1226,N_3460);
nand U8226 (N_8226,N_4788,N_438);
nand U8227 (N_8227,N_2806,N_1347);
nand U8228 (N_8228,N_3404,N_1390);
nor U8229 (N_8229,N_2954,N_2940);
nor U8230 (N_8230,N_251,N_2489);
and U8231 (N_8231,N_4123,N_2268);
nand U8232 (N_8232,N_1937,N_4221);
nor U8233 (N_8233,N_2177,N_457);
or U8234 (N_8234,N_1679,N_4058);
nor U8235 (N_8235,N_3135,N_3540);
nand U8236 (N_8236,N_1601,N_3077);
or U8237 (N_8237,N_525,N_994);
nand U8238 (N_8238,N_898,N_1406);
nand U8239 (N_8239,N_3174,N_2589);
nor U8240 (N_8240,N_4672,N_1466);
and U8241 (N_8241,N_926,N_3843);
nor U8242 (N_8242,N_4337,N_898);
nor U8243 (N_8243,N_38,N_1514);
and U8244 (N_8244,N_524,N_2632);
nor U8245 (N_8245,N_4969,N_4251);
and U8246 (N_8246,N_4523,N_2350);
and U8247 (N_8247,N_522,N_3506);
nand U8248 (N_8248,N_3238,N_2530);
and U8249 (N_8249,N_3893,N_910);
and U8250 (N_8250,N_1278,N_3783);
and U8251 (N_8251,N_2404,N_3955);
nand U8252 (N_8252,N_1523,N_2567);
nor U8253 (N_8253,N_1203,N_4988);
or U8254 (N_8254,N_1380,N_1138);
and U8255 (N_8255,N_4160,N_38);
and U8256 (N_8256,N_41,N_3605);
or U8257 (N_8257,N_275,N_4108);
nor U8258 (N_8258,N_4357,N_4599);
nand U8259 (N_8259,N_4427,N_2984);
and U8260 (N_8260,N_4643,N_3624);
or U8261 (N_8261,N_4724,N_1449);
nand U8262 (N_8262,N_2763,N_87);
nor U8263 (N_8263,N_928,N_2368);
nand U8264 (N_8264,N_3251,N_1859);
and U8265 (N_8265,N_97,N_67);
nor U8266 (N_8266,N_4773,N_345);
nand U8267 (N_8267,N_4698,N_4753);
nand U8268 (N_8268,N_578,N_957);
nor U8269 (N_8269,N_3707,N_1462);
nor U8270 (N_8270,N_2143,N_631);
or U8271 (N_8271,N_2638,N_1783);
nor U8272 (N_8272,N_1900,N_2317);
nor U8273 (N_8273,N_2812,N_595);
nor U8274 (N_8274,N_119,N_4168);
or U8275 (N_8275,N_4210,N_3585);
or U8276 (N_8276,N_1937,N_1668);
nand U8277 (N_8277,N_346,N_558);
nor U8278 (N_8278,N_1644,N_4769);
or U8279 (N_8279,N_1943,N_855);
xor U8280 (N_8280,N_2185,N_1219);
and U8281 (N_8281,N_1532,N_749);
nand U8282 (N_8282,N_559,N_4331);
and U8283 (N_8283,N_2253,N_1173);
nand U8284 (N_8284,N_1548,N_4544);
or U8285 (N_8285,N_122,N_858);
and U8286 (N_8286,N_1165,N_2178);
nor U8287 (N_8287,N_3814,N_801);
nand U8288 (N_8288,N_772,N_3847);
nor U8289 (N_8289,N_1101,N_3633);
nand U8290 (N_8290,N_2658,N_4978);
or U8291 (N_8291,N_189,N_4077);
xor U8292 (N_8292,N_3393,N_1257);
and U8293 (N_8293,N_4061,N_2354);
or U8294 (N_8294,N_3097,N_1078);
and U8295 (N_8295,N_880,N_4755);
nor U8296 (N_8296,N_1322,N_1840);
and U8297 (N_8297,N_1641,N_2785);
nor U8298 (N_8298,N_1840,N_3223);
nor U8299 (N_8299,N_1774,N_1749);
xor U8300 (N_8300,N_4890,N_3792);
nand U8301 (N_8301,N_1654,N_3690);
or U8302 (N_8302,N_3236,N_4311);
and U8303 (N_8303,N_1574,N_3064);
and U8304 (N_8304,N_4253,N_1954);
nand U8305 (N_8305,N_1026,N_1581);
and U8306 (N_8306,N_3405,N_1923);
and U8307 (N_8307,N_947,N_4776);
or U8308 (N_8308,N_4059,N_2534);
or U8309 (N_8309,N_2465,N_2136);
nor U8310 (N_8310,N_4721,N_4754);
nor U8311 (N_8311,N_719,N_3810);
nor U8312 (N_8312,N_338,N_2121);
and U8313 (N_8313,N_3784,N_3030);
nor U8314 (N_8314,N_1007,N_1574);
nor U8315 (N_8315,N_2870,N_2822);
or U8316 (N_8316,N_1226,N_4776);
or U8317 (N_8317,N_2752,N_2592);
or U8318 (N_8318,N_4342,N_4383);
nand U8319 (N_8319,N_207,N_1984);
nor U8320 (N_8320,N_4388,N_2589);
nor U8321 (N_8321,N_1552,N_908);
and U8322 (N_8322,N_2213,N_2994);
nor U8323 (N_8323,N_4643,N_1671);
nand U8324 (N_8324,N_4064,N_1135);
nor U8325 (N_8325,N_2074,N_2054);
nor U8326 (N_8326,N_1985,N_519);
nor U8327 (N_8327,N_1272,N_4166);
nand U8328 (N_8328,N_4052,N_52);
or U8329 (N_8329,N_1349,N_4749);
nand U8330 (N_8330,N_2960,N_495);
nand U8331 (N_8331,N_1448,N_4920);
nand U8332 (N_8332,N_4877,N_3772);
nand U8333 (N_8333,N_2346,N_1623);
and U8334 (N_8334,N_4575,N_4375);
nor U8335 (N_8335,N_1961,N_4970);
and U8336 (N_8336,N_1246,N_4797);
nand U8337 (N_8337,N_1375,N_2360);
nand U8338 (N_8338,N_2832,N_2660);
nor U8339 (N_8339,N_4137,N_1381);
or U8340 (N_8340,N_2383,N_4137);
and U8341 (N_8341,N_549,N_35);
nor U8342 (N_8342,N_2467,N_507);
and U8343 (N_8343,N_3813,N_1078);
nand U8344 (N_8344,N_4828,N_3692);
or U8345 (N_8345,N_3170,N_2100);
nand U8346 (N_8346,N_1883,N_228);
or U8347 (N_8347,N_270,N_479);
nor U8348 (N_8348,N_3659,N_3272);
nor U8349 (N_8349,N_1745,N_2485);
and U8350 (N_8350,N_4407,N_2605);
nand U8351 (N_8351,N_1659,N_1097);
nor U8352 (N_8352,N_1945,N_625);
or U8353 (N_8353,N_4012,N_4285);
nor U8354 (N_8354,N_1118,N_1939);
nand U8355 (N_8355,N_2215,N_4413);
nand U8356 (N_8356,N_3913,N_3054);
or U8357 (N_8357,N_880,N_2701);
or U8358 (N_8358,N_4617,N_1493);
and U8359 (N_8359,N_3371,N_819);
nand U8360 (N_8360,N_1097,N_907);
nor U8361 (N_8361,N_1184,N_2906);
or U8362 (N_8362,N_1031,N_1154);
nor U8363 (N_8363,N_2149,N_67);
and U8364 (N_8364,N_4867,N_3965);
or U8365 (N_8365,N_4594,N_2229);
and U8366 (N_8366,N_2651,N_2559);
nor U8367 (N_8367,N_3886,N_1206);
nand U8368 (N_8368,N_516,N_810);
nor U8369 (N_8369,N_2602,N_176);
nand U8370 (N_8370,N_939,N_3585);
or U8371 (N_8371,N_1745,N_3409);
nand U8372 (N_8372,N_4862,N_2558);
nand U8373 (N_8373,N_425,N_2005);
or U8374 (N_8374,N_1002,N_3117);
nand U8375 (N_8375,N_1210,N_2640);
nand U8376 (N_8376,N_1639,N_4941);
nor U8377 (N_8377,N_2907,N_258);
or U8378 (N_8378,N_4703,N_3876);
or U8379 (N_8379,N_1555,N_1942);
and U8380 (N_8380,N_3568,N_12);
and U8381 (N_8381,N_742,N_533);
or U8382 (N_8382,N_2291,N_3465);
and U8383 (N_8383,N_813,N_3985);
or U8384 (N_8384,N_4728,N_4573);
and U8385 (N_8385,N_4059,N_812);
nor U8386 (N_8386,N_3625,N_1137);
nand U8387 (N_8387,N_1602,N_4985);
or U8388 (N_8388,N_3485,N_2634);
nand U8389 (N_8389,N_3230,N_412);
and U8390 (N_8390,N_4062,N_1411);
and U8391 (N_8391,N_2095,N_347);
nor U8392 (N_8392,N_4283,N_3467);
and U8393 (N_8393,N_4759,N_3261);
nand U8394 (N_8394,N_114,N_1651);
or U8395 (N_8395,N_3338,N_1143);
nor U8396 (N_8396,N_2531,N_4302);
and U8397 (N_8397,N_2951,N_3255);
nand U8398 (N_8398,N_2650,N_1156);
nor U8399 (N_8399,N_3784,N_4827);
nor U8400 (N_8400,N_2249,N_799);
nor U8401 (N_8401,N_3656,N_3309);
or U8402 (N_8402,N_4072,N_4761);
nor U8403 (N_8403,N_3834,N_1960);
or U8404 (N_8404,N_2239,N_721);
nand U8405 (N_8405,N_20,N_924);
and U8406 (N_8406,N_4706,N_4926);
nand U8407 (N_8407,N_3610,N_1576);
and U8408 (N_8408,N_377,N_752);
nor U8409 (N_8409,N_529,N_4461);
or U8410 (N_8410,N_4114,N_4238);
and U8411 (N_8411,N_2255,N_4361);
or U8412 (N_8412,N_2279,N_397);
nor U8413 (N_8413,N_3710,N_3620);
nor U8414 (N_8414,N_2589,N_649);
nand U8415 (N_8415,N_1551,N_935);
xnor U8416 (N_8416,N_1324,N_2565);
nor U8417 (N_8417,N_2602,N_4388);
nand U8418 (N_8418,N_4938,N_753);
or U8419 (N_8419,N_2630,N_283);
nor U8420 (N_8420,N_1099,N_371);
and U8421 (N_8421,N_3664,N_2779);
and U8422 (N_8422,N_915,N_3418);
nand U8423 (N_8423,N_1443,N_4447);
nor U8424 (N_8424,N_3534,N_1347);
nand U8425 (N_8425,N_2861,N_2189);
or U8426 (N_8426,N_2038,N_210);
nand U8427 (N_8427,N_1668,N_1722);
or U8428 (N_8428,N_2465,N_1795);
and U8429 (N_8429,N_2625,N_1448);
and U8430 (N_8430,N_783,N_3055);
nor U8431 (N_8431,N_3475,N_2864);
nand U8432 (N_8432,N_2337,N_4582);
nor U8433 (N_8433,N_846,N_4281);
or U8434 (N_8434,N_4749,N_2182);
nand U8435 (N_8435,N_3128,N_819);
or U8436 (N_8436,N_1527,N_4208);
xnor U8437 (N_8437,N_4629,N_2945);
and U8438 (N_8438,N_4927,N_3211);
or U8439 (N_8439,N_128,N_550);
or U8440 (N_8440,N_4883,N_369);
nor U8441 (N_8441,N_1764,N_553);
and U8442 (N_8442,N_885,N_2967);
or U8443 (N_8443,N_813,N_4048);
nor U8444 (N_8444,N_114,N_2063);
nor U8445 (N_8445,N_4798,N_1763);
and U8446 (N_8446,N_2134,N_744);
nor U8447 (N_8447,N_3025,N_687);
or U8448 (N_8448,N_1926,N_3536);
nor U8449 (N_8449,N_4869,N_459);
and U8450 (N_8450,N_4075,N_930);
nor U8451 (N_8451,N_4137,N_1085);
nand U8452 (N_8452,N_4296,N_850);
nand U8453 (N_8453,N_3290,N_1638);
nor U8454 (N_8454,N_4089,N_2239);
or U8455 (N_8455,N_22,N_1614);
or U8456 (N_8456,N_2123,N_1560);
or U8457 (N_8457,N_1789,N_4462);
or U8458 (N_8458,N_1160,N_2116);
nor U8459 (N_8459,N_3132,N_943);
nor U8460 (N_8460,N_2933,N_570);
and U8461 (N_8461,N_3075,N_3099);
and U8462 (N_8462,N_2616,N_1902);
or U8463 (N_8463,N_38,N_2467);
or U8464 (N_8464,N_96,N_1794);
nand U8465 (N_8465,N_1863,N_1933);
and U8466 (N_8466,N_4039,N_1284);
or U8467 (N_8467,N_21,N_3182);
nor U8468 (N_8468,N_1489,N_3395);
and U8469 (N_8469,N_359,N_2074);
nor U8470 (N_8470,N_2584,N_1217);
or U8471 (N_8471,N_3934,N_120);
or U8472 (N_8472,N_3336,N_4257);
nor U8473 (N_8473,N_89,N_1376);
nor U8474 (N_8474,N_1772,N_384);
nand U8475 (N_8475,N_4619,N_4810);
nor U8476 (N_8476,N_63,N_788);
nor U8477 (N_8477,N_2987,N_4179);
nand U8478 (N_8478,N_655,N_3481);
nand U8479 (N_8479,N_1493,N_1391);
nand U8480 (N_8480,N_2170,N_3833);
nor U8481 (N_8481,N_3083,N_4452);
and U8482 (N_8482,N_4445,N_1602);
nand U8483 (N_8483,N_1363,N_3810);
nand U8484 (N_8484,N_2770,N_3443);
nand U8485 (N_8485,N_3635,N_4516);
nor U8486 (N_8486,N_4515,N_4562);
nand U8487 (N_8487,N_4985,N_3302);
nor U8488 (N_8488,N_391,N_3518);
or U8489 (N_8489,N_404,N_937);
and U8490 (N_8490,N_2039,N_4639);
or U8491 (N_8491,N_4375,N_876);
nor U8492 (N_8492,N_541,N_2443);
and U8493 (N_8493,N_2052,N_4768);
and U8494 (N_8494,N_1466,N_4889);
and U8495 (N_8495,N_561,N_847);
nor U8496 (N_8496,N_2186,N_4179);
and U8497 (N_8497,N_4457,N_3062);
xor U8498 (N_8498,N_529,N_365);
and U8499 (N_8499,N_4993,N_3674);
nand U8500 (N_8500,N_1491,N_2674);
nor U8501 (N_8501,N_2533,N_3183);
or U8502 (N_8502,N_821,N_2072);
nand U8503 (N_8503,N_2456,N_131);
nand U8504 (N_8504,N_3672,N_2941);
or U8505 (N_8505,N_725,N_3001);
nor U8506 (N_8506,N_3140,N_4133);
and U8507 (N_8507,N_4065,N_4041);
nor U8508 (N_8508,N_546,N_4505);
nand U8509 (N_8509,N_2156,N_3013);
and U8510 (N_8510,N_396,N_1349);
or U8511 (N_8511,N_2353,N_677);
nand U8512 (N_8512,N_4387,N_901);
nand U8513 (N_8513,N_2650,N_649);
nand U8514 (N_8514,N_586,N_4329);
nand U8515 (N_8515,N_3185,N_3067);
or U8516 (N_8516,N_3633,N_3578);
and U8517 (N_8517,N_4056,N_3487);
xnor U8518 (N_8518,N_3923,N_1655);
and U8519 (N_8519,N_3714,N_4760);
and U8520 (N_8520,N_1306,N_87);
nor U8521 (N_8521,N_759,N_4229);
and U8522 (N_8522,N_3335,N_2646);
nor U8523 (N_8523,N_1212,N_1142);
xor U8524 (N_8524,N_3379,N_1729);
or U8525 (N_8525,N_321,N_2172);
or U8526 (N_8526,N_1911,N_1992);
and U8527 (N_8527,N_3923,N_191);
and U8528 (N_8528,N_2146,N_2226);
or U8529 (N_8529,N_1881,N_2180);
or U8530 (N_8530,N_4316,N_4143);
or U8531 (N_8531,N_3574,N_3932);
and U8532 (N_8532,N_4573,N_2372);
or U8533 (N_8533,N_2592,N_3776);
nor U8534 (N_8534,N_125,N_3724);
nand U8535 (N_8535,N_1918,N_3287);
or U8536 (N_8536,N_3556,N_4427);
or U8537 (N_8537,N_2765,N_1015);
nor U8538 (N_8538,N_1746,N_2547);
nor U8539 (N_8539,N_3387,N_4551);
nand U8540 (N_8540,N_1155,N_1885);
and U8541 (N_8541,N_1464,N_4845);
or U8542 (N_8542,N_2738,N_1147);
nand U8543 (N_8543,N_4097,N_970);
nand U8544 (N_8544,N_3747,N_4077);
or U8545 (N_8545,N_644,N_1881);
and U8546 (N_8546,N_314,N_4023);
nor U8547 (N_8547,N_3251,N_3998);
nand U8548 (N_8548,N_1299,N_1827);
or U8549 (N_8549,N_4363,N_983);
nor U8550 (N_8550,N_2103,N_4242);
or U8551 (N_8551,N_3380,N_4105);
nor U8552 (N_8552,N_3734,N_3719);
nor U8553 (N_8553,N_3794,N_214);
and U8554 (N_8554,N_488,N_197);
nand U8555 (N_8555,N_2871,N_2970);
and U8556 (N_8556,N_1269,N_1483);
xnor U8557 (N_8557,N_763,N_1255);
nand U8558 (N_8558,N_887,N_39);
nand U8559 (N_8559,N_4020,N_4736);
nor U8560 (N_8560,N_3113,N_3590);
or U8561 (N_8561,N_4049,N_701);
nand U8562 (N_8562,N_2650,N_4555);
nand U8563 (N_8563,N_1122,N_4834);
and U8564 (N_8564,N_636,N_4687);
nand U8565 (N_8565,N_1122,N_848);
or U8566 (N_8566,N_3991,N_4644);
nand U8567 (N_8567,N_1793,N_4229);
nand U8568 (N_8568,N_94,N_1866);
nand U8569 (N_8569,N_4308,N_4610);
or U8570 (N_8570,N_1997,N_4416);
xor U8571 (N_8571,N_1395,N_1747);
nor U8572 (N_8572,N_1521,N_59);
and U8573 (N_8573,N_3006,N_384);
and U8574 (N_8574,N_2202,N_484);
nand U8575 (N_8575,N_61,N_3504);
and U8576 (N_8576,N_4717,N_1388);
nand U8577 (N_8577,N_822,N_1210);
and U8578 (N_8578,N_3748,N_1187);
nand U8579 (N_8579,N_654,N_2464);
or U8580 (N_8580,N_3553,N_2635);
or U8581 (N_8581,N_4155,N_2615);
or U8582 (N_8582,N_2066,N_941);
or U8583 (N_8583,N_396,N_1596);
and U8584 (N_8584,N_249,N_63);
and U8585 (N_8585,N_4687,N_3161);
nor U8586 (N_8586,N_1551,N_1888);
nor U8587 (N_8587,N_1250,N_2236);
and U8588 (N_8588,N_1790,N_2216);
nor U8589 (N_8589,N_4322,N_2184);
nor U8590 (N_8590,N_3955,N_3897);
nor U8591 (N_8591,N_4153,N_2486);
nand U8592 (N_8592,N_2561,N_934);
and U8593 (N_8593,N_2259,N_1038);
nor U8594 (N_8594,N_1267,N_1106);
nand U8595 (N_8595,N_1479,N_4265);
nand U8596 (N_8596,N_4378,N_521);
nor U8597 (N_8597,N_1306,N_3820);
nand U8598 (N_8598,N_3883,N_2469);
and U8599 (N_8599,N_4120,N_3868);
nand U8600 (N_8600,N_1466,N_3919);
xor U8601 (N_8601,N_1230,N_2984);
or U8602 (N_8602,N_4432,N_3340);
nand U8603 (N_8603,N_4070,N_1537);
or U8604 (N_8604,N_1789,N_1282);
and U8605 (N_8605,N_1796,N_4807);
nand U8606 (N_8606,N_2631,N_2149);
nor U8607 (N_8607,N_2691,N_4384);
nor U8608 (N_8608,N_2339,N_4579);
nor U8609 (N_8609,N_4218,N_924);
nand U8610 (N_8610,N_2724,N_4951);
nor U8611 (N_8611,N_3677,N_1910);
nand U8612 (N_8612,N_3333,N_1844);
or U8613 (N_8613,N_4870,N_2302);
nand U8614 (N_8614,N_2719,N_3231);
and U8615 (N_8615,N_4792,N_3707);
or U8616 (N_8616,N_3810,N_216);
or U8617 (N_8617,N_2139,N_5);
nor U8618 (N_8618,N_4845,N_551);
nor U8619 (N_8619,N_3934,N_2557);
nand U8620 (N_8620,N_4486,N_2051);
and U8621 (N_8621,N_3293,N_2480);
nand U8622 (N_8622,N_4807,N_2783);
or U8623 (N_8623,N_1620,N_254);
nor U8624 (N_8624,N_1370,N_3012);
or U8625 (N_8625,N_4219,N_2902);
nand U8626 (N_8626,N_4924,N_4115);
and U8627 (N_8627,N_3419,N_2835);
nor U8628 (N_8628,N_4794,N_4360);
nand U8629 (N_8629,N_3921,N_4534);
nor U8630 (N_8630,N_212,N_2535);
nor U8631 (N_8631,N_3900,N_2936);
nand U8632 (N_8632,N_1252,N_3559);
and U8633 (N_8633,N_4116,N_3204);
nand U8634 (N_8634,N_1839,N_4724);
nand U8635 (N_8635,N_4990,N_3256);
or U8636 (N_8636,N_1685,N_2614);
and U8637 (N_8637,N_2032,N_4631);
nand U8638 (N_8638,N_1036,N_1396);
nor U8639 (N_8639,N_4591,N_2814);
nand U8640 (N_8640,N_4970,N_1818);
and U8641 (N_8641,N_3639,N_2727);
nor U8642 (N_8642,N_2448,N_4238);
nor U8643 (N_8643,N_2553,N_1063);
and U8644 (N_8644,N_393,N_3052);
nand U8645 (N_8645,N_812,N_2739);
or U8646 (N_8646,N_2831,N_929);
or U8647 (N_8647,N_3932,N_2378);
or U8648 (N_8648,N_4843,N_2972);
and U8649 (N_8649,N_3264,N_2645);
nand U8650 (N_8650,N_4792,N_2856);
or U8651 (N_8651,N_1924,N_1791);
nand U8652 (N_8652,N_2625,N_4858);
xor U8653 (N_8653,N_3888,N_3321);
and U8654 (N_8654,N_730,N_1267);
nand U8655 (N_8655,N_4643,N_3308);
or U8656 (N_8656,N_2794,N_1957);
and U8657 (N_8657,N_226,N_1380);
nor U8658 (N_8658,N_3009,N_2484);
and U8659 (N_8659,N_825,N_4342);
nor U8660 (N_8660,N_1970,N_2882);
nand U8661 (N_8661,N_4243,N_2004);
and U8662 (N_8662,N_2337,N_2325);
or U8663 (N_8663,N_700,N_2119);
or U8664 (N_8664,N_1701,N_3784);
and U8665 (N_8665,N_4307,N_1603);
nor U8666 (N_8666,N_1850,N_2913);
and U8667 (N_8667,N_2689,N_4509);
nand U8668 (N_8668,N_3765,N_3488);
and U8669 (N_8669,N_2363,N_4129);
xor U8670 (N_8670,N_1801,N_3569);
and U8671 (N_8671,N_1094,N_733);
and U8672 (N_8672,N_1770,N_2075);
and U8673 (N_8673,N_199,N_4690);
nand U8674 (N_8674,N_691,N_4226);
nor U8675 (N_8675,N_3620,N_4212);
nand U8676 (N_8676,N_3961,N_513);
or U8677 (N_8677,N_3037,N_2855);
or U8678 (N_8678,N_3404,N_4066);
or U8679 (N_8679,N_3787,N_467);
or U8680 (N_8680,N_2368,N_3043);
nor U8681 (N_8681,N_3936,N_3651);
and U8682 (N_8682,N_1851,N_3107);
nand U8683 (N_8683,N_618,N_763);
nand U8684 (N_8684,N_4928,N_3303);
or U8685 (N_8685,N_76,N_2535);
and U8686 (N_8686,N_2845,N_5);
or U8687 (N_8687,N_938,N_4938);
and U8688 (N_8688,N_1701,N_1423);
or U8689 (N_8689,N_2639,N_3289);
and U8690 (N_8690,N_2216,N_125);
and U8691 (N_8691,N_741,N_4901);
nor U8692 (N_8692,N_969,N_3359);
xor U8693 (N_8693,N_4777,N_792);
and U8694 (N_8694,N_314,N_2753);
and U8695 (N_8695,N_3034,N_4116);
nand U8696 (N_8696,N_1083,N_1232);
and U8697 (N_8697,N_1519,N_1707);
and U8698 (N_8698,N_715,N_4743);
nand U8699 (N_8699,N_4070,N_3754);
nand U8700 (N_8700,N_2209,N_2715);
or U8701 (N_8701,N_4433,N_3325);
and U8702 (N_8702,N_4293,N_4379);
or U8703 (N_8703,N_2561,N_1893);
and U8704 (N_8704,N_1582,N_3352);
nor U8705 (N_8705,N_2622,N_4504);
and U8706 (N_8706,N_1722,N_3194);
and U8707 (N_8707,N_2174,N_59);
and U8708 (N_8708,N_2602,N_2015);
nor U8709 (N_8709,N_4812,N_2359);
or U8710 (N_8710,N_4181,N_3715);
nand U8711 (N_8711,N_1919,N_1812);
nand U8712 (N_8712,N_4832,N_473);
and U8713 (N_8713,N_3424,N_650);
or U8714 (N_8714,N_2796,N_799);
nor U8715 (N_8715,N_3108,N_684);
nor U8716 (N_8716,N_3117,N_2714);
and U8717 (N_8717,N_2902,N_1756);
or U8718 (N_8718,N_2001,N_2483);
and U8719 (N_8719,N_2559,N_3952);
nor U8720 (N_8720,N_2494,N_4398);
nor U8721 (N_8721,N_2237,N_513);
nor U8722 (N_8722,N_1791,N_2901);
and U8723 (N_8723,N_964,N_3555);
or U8724 (N_8724,N_203,N_1609);
and U8725 (N_8725,N_616,N_4128);
and U8726 (N_8726,N_737,N_2637);
and U8727 (N_8727,N_2116,N_2171);
or U8728 (N_8728,N_646,N_3921);
nor U8729 (N_8729,N_971,N_882);
nand U8730 (N_8730,N_3754,N_3294);
nand U8731 (N_8731,N_1387,N_3248);
or U8732 (N_8732,N_459,N_4785);
or U8733 (N_8733,N_976,N_3990);
nor U8734 (N_8734,N_253,N_2535);
nand U8735 (N_8735,N_1109,N_2119);
and U8736 (N_8736,N_3119,N_4302);
or U8737 (N_8737,N_4647,N_2371);
or U8738 (N_8738,N_3782,N_1529);
or U8739 (N_8739,N_1106,N_3934);
nand U8740 (N_8740,N_172,N_4975);
or U8741 (N_8741,N_4734,N_3652);
nand U8742 (N_8742,N_2028,N_3736);
nand U8743 (N_8743,N_913,N_2872);
nand U8744 (N_8744,N_4465,N_2205);
nor U8745 (N_8745,N_1141,N_2590);
and U8746 (N_8746,N_2750,N_3642);
and U8747 (N_8747,N_3806,N_57);
nor U8748 (N_8748,N_4476,N_4083);
nand U8749 (N_8749,N_569,N_918);
nand U8750 (N_8750,N_2345,N_3941);
nand U8751 (N_8751,N_524,N_1640);
or U8752 (N_8752,N_4710,N_2758);
nor U8753 (N_8753,N_4615,N_2151);
or U8754 (N_8754,N_4497,N_579);
nand U8755 (N_8755,N_1202,N_4112);
nand U8756 (N_8756,N_1936,N_2358);
nor U8757 (N_8757,N_2312,N_4858);
nand U8758 (N_8758,N_1954,N_759);
nand U8759 (N_8759,N_72,N_720);
and U8760 (N_8760,N_4543,N_4783);
or U8761 (N_8761,N_1236,N_1886);
and U8762 (N_8762,N_2840,N_2651);
or U8763 (N_8763,N_4332,N_621);
nor U8764 (N_8764,N_1517,N_2808);
nand U8765 (N_8765,N_1247,N_294);
or U8766 (N_8766,N_2162,N_2400);
nand U8767 (N_8767,N_4999,N_4927);
and U8768 (N_8768,N_4187,N_4219);
xnor U8769 (N_8769,N_1535,N_240);
nor U8770 (N_8770,N_4042,N_1750);
nor U8771 (N_8771,N_4676,N_3065);
or U8772 (N_8772,N_2755,N_3875);
nor U8773 (N_8773,N_664,N_1791);
nor U8774 (N_8774,N_632,N_1635);
nand U8775 (N_8775,N_485,N_3065);
nor U8776 (N_8776,N_3320,N_3504);
nand U8777 (N_8777,N_1421,N_4184);
and U8778 (N_8778,N_3712,N_4161);
and U8779 (N_8779,N_369,N_4159);
nor U8780 (N_8780,N_2537,N_4306);
and U8781 (N_8781,N_4455,N_3059);
and U8782 (N_8782,N_4877,N_1265);
nand U8783 (N_8783,N_4450,N_4221);
nand U8784 (N_8784,N_4172,N_1262);
or U8785 (N_8785,N_4469,N_3471);
or U8786 (N_8786,N_2645,N_4975);
or U8787 (N_8787,N_1900,N_2019);
or U8788 (N_8788,N_498,N_4124);
nor U8789 (N_8789,N_4613,N_4784);
or U8790 (N_8790,N_3324,N_3012);
nor U8791 (N_8791,N_1823,N_1512);
nand U8792 (N_8792,N_1298,N_2582);
nand U8793 (N_8793,N_1147,N_1855);
nor U8794 (N_8794,N_4402,N_42);
and U8795 (N_8795,N_3715,N_362);
nor U8796 (N_8796,N_2667,N_3625);
nand U8797 (N_8797,N_2662,N_4033);
nand U8798 (N_8798,N_4421,N_1486);
or U8799 (N_8799,N_1828,N_2130);
and U8800 (N_8800,N_3292,N_1974);
or U8801 (N_8801,N_4218,N_4096);
and U8802 (N_8802,N_505,N_4849);
and U8803 (N_8803,N_4059,N_4819);
or U8804 (N_8804,N_1855,N_1878);
nand U8805 (N_8805,N_3197,N_638);
nand U8806 (N_8806,N_103,N_1653);
nand U8807 (N_8807,N_467,N_2423);
nor U8808 (N_8808,N_2927,N_1170);
or U8809 (N_8809,N_499,N_1541);
nor U8810 (N_8810,N_3790,N_1607);
or U8811 (N_8811,N_2808,N_918);
and U8812 (N_8812,N_4871,N_280);
xnor U8813 (N_8813,N_4624,N_1440);
or U8814 (N_8814,N_1279,N_478);
nor U8815 (N_8815,N_845,N_4007);
nand U8816 (N_8816,N_656,N_1305);
nand U8817 (N_8817,N_346,N_4019);
nor U8818 (N_8818,N_607,N_1813);
or U8819 (N_8819,N_660,N_500);
nor U8820 (N_8820,N_3289,N_1741);
nand U8821 (N_8821,N_681,N_2936);
nor U8822 (N_8822,N_4613,N_4008);
or U8823 (N_8823,N_1181,N_3145);
or U8824 (N_8824,N_4493,N_3097);
and U8825 (N_8825,N_396,N_1762);
nor U8826 (N_8826,N_65,N_3926);
nand U8827 (N_8827,N_3140,N_1459);
nor U8828 (N_8828,N_3327,N_1049);
or U8829 (N_8829,N_911,N_356);
and U8830 (N_8830,N_240,N_425);
or U8831 (N_8831,N_2509,N_3775);
or U8832 (N_8832,N_2092,N_4133);
nor U8833 (N_8833,N_4038,N_3184);
or U8834 (N_8834,N_4694,N_1314);
nor U8835 (N_8835,N_3686,N_687);
and U8836 (N_8836,N_1818,N_2229);
nand U8837 (N_8837,N_1041,N_389);
nand U8838 (N_8838,N_1708,N_727);
nand U8839 (N_8839,N_1581,N_3519);
and U8840 (N_8840,N_2093,N_1578);
nor U8841 (N_8841,N_2310,N_111);
or U8842 (N_8842,N_2471,N_2115);
nand U8843 (N_8843,N_160,N_4369);
nand U8844 (N_8844,N_2110,N_2589);
nor U8845 (N_8845,N_3428,N_3012);
or U8846 (N_8846,N_4303,N_1858);
or U8847 (N_8847,N_3716,N_1819);
nor U8848 (N_8848,N_3268,N_3774);
nor U8849 (N_8849,N_1915,N_2952);
or U8850 (N_8850,N_4673,N_100);
or U8851 (N_8851,N_3254,N_3939);
and U8852 (N_8852,N_3622,N_1543);
nor U8853 (N_8853,N_1436,N_52);
nor U8854 (N_8854,N_2122,N_4238);
nor U8855 (N_8855,N_3968,N_607);
and U8856 (N_8856,N_4369,N_1966);
and U8857 (N_8857,N_2142,N_2396);
or U8858 (N_8858,N_4671,N_4724);
nor U8859 (N_8859,N_1780,N_4695);
nor U8860 (N_8860,N_4464,N_3501);
nor U8861 (N_8861,N_4751,N_3601);
or U8862 (N_8862,N_1452,N_1265);
nor U8863 (N_8863,N_1654,N_2125);
and U8864 (N_8864,N_4451,N_442);
and U8865 (N_8865,N_34,N_1395);
nand U8866 (N_8866,N_809,N_813);
or U8867 (N_8867,N_1114,N_3144);
and U8868 (N_8868,N_1390,N_1407);
nand U8869 (N_8869,N_4515,N_3936);
nor U8870 (N_8870,N_791,N_4061);
nand U8871 (N_8871,N_279,N_4152);
nand U8872 (N_8872,N_4944,N_302);
nor U8873 (N_8873,N_2873,N_613);
and U8874 (N_8874,N_1058,N_1442);
nor U8875 (N_8875,N_2096,N_3129);
nand U8876 (N_8876,N_4130,N_2344);
nand U8877 (N_8877,N_1955,N_1925);
and U8878 (N_8878,N_4466,N_3452);
nor U8879 (N_8879,N_1754,N_1110);
nor U8880 (N_8880,N_2119,N_2620);
nand U8881 (N_8881,N_3117,N_4553);
or U8882 (N_8882,N_422,N_4886);
xnor U8883 (N_8883,N_3229,N_4524);
and U8884 (N_8884,N_2030,N_650);
or U8885 (N_8885,N_590,N_1133);
nor U8886 (N_8886,N_3419,N_1057);
nand U8887 (N_8887,N_4811,N_1913);
and U8888 (N_8888,N_3047,N_3748);
nand U8889 (N_8889,N_3105,N_1257);
nand U8890 (N_8890,N_872,N_3630);
nand U8891 (N_8891,N_1414,N_1933);
nor U8892 (N_8892,N_294,N_4812);
or U8893 (N_8893,N_3155,N_951);
or U8894 (N_8894,N_3842,N_1479);
nor U8895 (N_8895,N_774,N_938);
xor U8896 (N_8896,N_1382,N_75);
nor U8897 (N_8897,N_2753,N_3942);
nor U8898 (N_8898,N_1250,N_2772);
nor U8899 (N_8899,N_1159,N_2621);
or U8900 (N_8900,N_1595,N_2272);
nor U8901 (N_8901,N_2459,N_1720);
nor U8902 (N_8902,N_4825,N_1495);
or U8903 (N_8903,N_4729,N_4057);
and U8904 (N_8904,N_2212,N_536);
nand U8905 (N_8905,N_4884,N_4626);
nor U8906 (N_8906,N_531,N_2058);
nor U8907 (N_8907,N_2399,N_4200);
or U8908 (N_8908,N_2193,N_3072);
nor U8909 (N_8909,N_3706,N_3468);
and U8910 (N_8910,N_4009,N_3400);
or U8911 (N_8911,N_685,N_25);
or U8912 (N_8912,N_4741,N_1209);
and U8913 (N_8913,N_2617,N_2802);
nand U8914 (N_8914,N_4487,N_1470);
or U8915 (N_8915,N_3701,N_931);
and U8916 (N_8916,N_4265,N_4770);
nand U8917 (N_8917,N_3186,N_3168);
and U8918 (N_8918,N_1827,N_3594);
nor U8919 (N_8919,N_830,N_3211);
nor U8920 (N_8920,N_4107,N_4833);
nor U8921 (N_8921,N_2177,N_1030);
nor U8922 (N_8922,N_4810,N_3394);
or U8923 (N_8923,N_2,N_1547);
nor U8924 (N_8924,N_4378,N_2947);
nor U8925 (N_8925,N_4891,N_337);
and U8926 (N_8926,N_3093,N_2296);
and U8927 (N_8927,N_712,N_1899);
or U8928 (N_8928,N_4265,N_907);
nand U8929 (N_8929,N_2397,N_672);
nor U8930 (N_8930,N_3960,N_4849);
nor U8931 (N_8931,N_4670,N_2573);
nand U8932 (N_8932,N_3645,N_4268);
nand U8933 (N_8933,N_4073,N_733);
or U8934 (N_8934,N_1945,N_2829);
nor U8935 (N_8935,N_2344,N_2896);
and U8936 (N_8936,N_683,N_758);
or U8937 (N_8937,N_4333,N_1546);
nor U8938 (N_8938,N_3402,N_3937);
or U8939 (N_8939,N_971,N_1233);
and U8940 (N_8940,N_286,N_4667);
nand U8941 (N_8941,N_613,N_1722);
nor U8942 (N_8942,N_2141,N_3288);
or U8943 (N_8943,N_4135,N_2017);
nor U8944 (N_8944,N_4511,N_2182);
or U8945 (N_8945,N_2074,N_1628);
nand U8946 (N_8946,N_1529,N_4770);
nor U8947 (N_8947,N_1313,N_1785);
nand U8948 (N_8948,N_2123,N_817);
or U8949 (N_8949,N_3255,N_3146);
nand U8950 (N_8950,N_873,N_4030);
nand U8951 (N_8951,N_1872,N_1114);
nand U8952 (N_8952,N_2985,N_1784);
or U8953 (N_8953,N_4846,N_4657);
or U8954 (N_8954,N_1702,N_2968);
nand U8955 (N_8955,N_657,N_1652);
nor U8956 (N_8956,N_2547,N_2078);
and U8957 (N_8957,N_3269,N_822);
nor U8958 (N_8958,N_3808,N_761);
nand U8959 (N_8959,N_1578,N_192);
or U8960 (N_8960,N_4786,N_4896);
nand U8961 (N_8961,N_2651,N_316);
and U8962 (N_8962,N_1003,N_884);
nand U8963 (N_8963,N_4185,N_2771);
nor U8964 (N_8964,N_3587,N_1203);
xor U8965 (N_8965,N_2350,N_1036);
or U8966 (N_8966,N_1194,N_3041);
or U8967 (N_8967,N_2844,N_462);
and U8968 (N_8968,N_4217,N_4049);
and U8969 (N_8969,N_3792,N_1496);
and U8970 (N_8970,N_4610,N_3483);
and U8971 (N_8971,N_2997,N_1073);
or U8972 (N_8972,N_1129,N_73);
nand U8973 (N_8973,N_4250,N_1120);
and U8974 (N_8974,N_4460,N_3699);
nor U8975 (N_8975,N_1402,N_4214);
and U8976 (N_8976,N_1502,N_4491);
or U8977 (N_8977,N_1686,N_435);
nand U8978 (N_8978,N_4845,N_824);
nor U8979 (N_8979,N_2128,N_1328);
or U8980 (N_8980,N_283,N_2660);
and U8981 (N_8981,N_894,N_2232);
nor U8982 (N_8982,N_4368,N_4538);
or U8983 (N_8983,N_4869,N_3512);
or U8984 (N_8984,N_3425,N_4800);
and U8985 (N_8985,N_770,N_2630);
and U8986 (N_8986,N_2826,N_3055);
nand U8987 (N_8987,N_518,N_4569);
nor U8988 (N_8988,N_2685,N_4487);
nor U8989 (N_8989,N_1320,N_2961);
and U8990 (N_8990,N_2795,N_46);
or U8991 (N_8991,N_736,N_4484);
or U8992 (N_8992,N_1259,N_388);
nand U8993 (N_8993,N_3391,N_4253);
or U8994 (N_8994,N_4364,N_1532);
nand U8995 (N_8995,N_1467,N_3788);
nor U8996 (N_8996,N_124,N_4764);
nand U8997 (N_8997,N_3818,N_4200);
or U8998 (N_8998,N_2692,N_3227);
xor U8999 (N_8999,N_1309,N_1628);
or U9000 (N_9000,N_2433,N_588);
and U9001 (N_9001,N_2765,N_3754);
nor U9002 (N_9002,N_60,N_1907);
or U9003 (N_9003,N_1824,N_4329);
nor U9004 (N_9004,N_2220,N_3642);
and U9005 (N_9005,N_1595,N_613);
nand U9006 (N_9006,N_2561,N_4358);
or U9007 (N_9007,N_3788,N_4812);
or U9008 (N_9008,N_3032,N_1148);
nand U9009 (N_9009,N_4564,N_581);
nand U9010 (N_9010,N_1659,N_3469);
or U9011 (N_9011,N_1658,N_3491);
nor U9012 (N_9012,N_4323,N_1136);
nor U9013 (N_9013,N_2462,N_3171);
nor U9014 (N_9014,N_3167,N_4600);
xor U9015 (N_9015,N_1472,N_1695);
or U9016 (N_9016,N_1388,N_3068);
nand U9017 (N_9017,N_2318,N_587);
and U9018 (N_9018,N_4210,N_3224);
and U9019 (N_9019,N_2401,N_1882);
or U9020 (N_9020,N_2474,N_363);
and U9021 (N_9021,N_1144,N_3061);
nor U9022 (N_9022,N_747,N_1045);
nand U9023 (N_9023,N_3926,N_805);
or U9024 (N_9024,N_657,N_3908);
or U9025 (N_9025,N_3120,N_2421);
and U9026 (N_9026,N_4568,N_1358);
nor U9027 (N_9027,N_4586,N_4065);
nor U9028 (N_9028,N_4947,N_3716);
or U9029 (N_9029,N_3064,N_849);
and U9030 (N_9030,N_4689,N_1429);
and U9031 (N_9031,N_731,N_3732);
nand U9032 (N_9032,N_3233,N_4080);
nand U9033 (N_9033,N_2318,N_3243);
or U9034 (N_9034,N_2008,N_391);
and U9035 (N_9035,N_4339,N_1798);
nand U9036 (N_9036,N_3924,N_4170);
or U9037 (N_9037,N_886,N_2798);
nand U9038 (N_9038,N_2878,N_2558);
or U9039 (N_9039,N_432,N_2730);
and U9040 (N_9040,N_447,N_630);
and U9041 (N_9041,N_4268,N_4541);
nor U9042 (N_9042,N_441,N_3324);
nand U9043 (N_9043,N_2693,N_1743);
and U9044 (N_9044,N_354,N_489);
nand U9045 (N_9045,N_4290,N_2388);
or U9046 (N_9046,N_1240,N_4259);
nor U9047 (N_9047,N_1879,N_641);
or U9048 (N_9048,N_3727,N_747);
nor U9049 (N_9049,N_3027,N_1583);
nand U9050 (N_9050,N_859,N_2151);
nor U9051 (N_9051,N_97,N_1791);
or U9052 (N_9052,N_1964,N_1201);
or U9053 (N_9053,N_4652,N_354);
or U9054 (N_9054,N_2914,N_1585);
or U9055 (N_9055,N_3828,N_4872);
and U9056 (N_9056,N_103,N_2624);
nand U9057 (N_9057,N_1471,N_3913);
and U9058 (N_9058,N_4884,N_3422);
and U9059 (N_9059,N_1448,N_737);
nor U9060 (N_9060,N_2376,N_1427);
nor U9061 (N_9061,N_3986,N_2344);
nor U9062 (N_9062,N_679,N_3422);
nand U9063 (N_9063,N_394,N_404);
nor U9064 (N_9064,N_4685,N_1123);
and U9065 (N_9065,N_1957,N_2601);
or U9066 (N_9066,N_3375,N_3135);
nand U9067 (N_9067,N_4378,N_414);
nor U9068 (N_9068,N_4123,N_1898);
nand U9069 (N_9069,N_1149,N_953);
nor U9070 (N_9070,N_4985,N_2578);
xnor U9071 (N_9071,N_1455,N_103);
nor U9072 (N_9072,N_1980,N_4487);
nor U9073 (N_9073,N_4293,N_1219);
nor U9074 (N_9074,N_925,N_952);
or U9075 (N_9075,N_2654,N_4049);
nand U9076 (N_9076,N_150,N_4689);
and U9077 (N_9077,N_3934,N_2742);
or U9078 (N_9078,N_826,N_665);
and U9079 (N_9079,N_1180,N_448);
nor U9080 (N_9080,N_2319,N_3360);
or U9081 (N_9081,N_1315,N_2981);
and U9082 (N_9082,N_209,N_2218);
and U9083 (N_9083,N_154,N_1930);
nor U9084 (N_9084,N_2636,N_91);
nand U9085 (N_9085,N_4691,N_2614);
or U9086 (N_9086,N_1550,N_2971);
xnor U9087 (N_9087,N_4364,N_4290);
nand U9088 (N_9088,N_1680,N_3474);
nand U9089 (N_9089,N_131,N_3185);
and U9090 (N_9090,N_4771,N_2301);
and U9091 (N_9091,N_2489,N_4962);
and U9092 (N_9092,N_1575,N_2950);
nand U9093 (N_9093,N_839,N_2444);
and U9094 (N_9094,N_1280,N_771);
and U9095 (N_9095,N_3101,N_1705);
and U9096 (N_9096,N_2876,N_2185);
or U9097 (N_9097,N_4047,N_2206);
nand U9098 (N_9098,N_4043,N_1437);
nand U9099 (N_9099,N_1337,N_4704);
nand U9100 (N_9100,N_1246,N_262);
and U9101 (N_9101,N_1376,N_4036);
and U9102 (N_9102,N_664,N_4355);
nand U9103 (N_9103,N_2250,N_4716);
and U9104 (N_9104,N_1918,N_4901);
nor U9105 (N_9105,N_3621,N_1286);
nor U9106 (N_9106,N_75,N_2842);
nor U9107 (N_9107,N_2434,N_4899);
nand U9108 (N_9108,N_784,N_329);
nand U9109 (N_9109,N_4208,N_1335);
nand U9110 (N_9110,N_2824,N_1328);
nand U9111 (N_9111,N_1060,N_3404);
nand U9112 (N_9112,N_2054,N_1677);
or U9113 (N_9113,N_1510,N_40);
or U9114 (N_9114,N_2113,N_3147);
or U9115 (N_9115,N_834,N_2215);
or U9116 (N_9116,N_3486,N_1682);
nor U9117 (N_9117,N_2055,N_3733);
or U9118 (N_9118,N_1848,N_4650);
nor U9119 (N_9119,N_3700,N_2905);
nor U9120 (N_9120,N_2550,N_2180);
nand U9121 (N_9121,N_3671,N_2318);
or U9122 (N_9122,N_3695,N_3339);
and U9123 (N_9123,N_521,N_1643);
or U9124 (N_9124,N_2188,N_1571);
and U9125 (N_9125,N_1879,N_670);
or U9126 (N_9126,N_3190,N_2693);
and U9127 (N_9127,N_4443,N_1015);
and U9128 (N_9128,N_3248,N_3210);
or U9129 (N_9129,N_1427,N_4985);
nor U9130 (N_9130,N_3772,N_1483);
nand U9131 (N_9131,N_2335,N_4199);
and U9132 (N_9132,N_1174,N_3340);
nand U9133 (N_9133,N_4640,N_1081);
or U9134 (N_9134,N_4698,N_352);
and U9135 (N_9135,N_2059,N_439);
and U9136 (N_9136,N_3339,N_1778);
nand U9137 (N_9137,N_2898,N_3336);
and U9138 (N_9138,N_4443,N_170);
nor U9139 (N_9139,N_309,N_4749);
nand U9140 (N_9140,N_3456,N_2874);
and U9141 (N_9141,N_1212,N_4975);
or U9142 (N_9142,N_2333,N_2831);
and U9143 (N_9143,N_723,N_2268);
or U9144 (N_9144,N_2075,N_1581);
or U9145 (N_9145,N_3379,N_3022);
and U9146 (N_9146,N_3836,N_1607);
nor U9147 (N_9147,N_241,N_1749);
nand U9148 (N_9148,N_2071,N_1370);
nand U9149 (N_9149,N_2725,N_4806);
nand U9150 (N_9150,N_3517,N_4826);
nor U9151 (N_9151,N_3548,N_1441);
nor U9152 (N_9152,N_3565,N_1614);
and U9153 (N_9153,N_1510,N_269);
or U9154 (N_9154,N_166,N_784);
nor U9155 (N_9155,N_4873,N_2964);
nand U9156 (N_9156,N_2184,N_1960);
or U9157 (N_9157,N_3881,N_1948);
or U9158 (N_9158,N_1112,N_3997);
and U9159 (N_9159,N_414,N_184);
and U9160 (N_9160,N_177,N_4836);
nand U9161 (N_9161,N_550,N_2856);
or U9162 (N_9162,N_15,N_4850);
nand U9163 (N_9163,N_968,N_2036);
nor U9164 (N_9164,N_559,N_2597);
or U9165 (N_9165,N_849,N_1826);
and U9166 (N_9166,N_3120,N_2355);
nand U9167 (N_9167,N_3440,N_1463);
or U9168 (N_9168,N_4365,N_862);
and U9169 (N_9169,N_4081,N_2102);
or U9170 (N_9170,N_1050,N_1892);
nor U9171 (N_9171,N_1648,N_4886);
or U9172 (N_9172,N_3315,N_3910);
nor U9173 (N_9173,N_2799,N_2662);
nor U9174 (N_9174,N_106,N_3895);
or U9175 (N_9175,N_4749,N_3836);
and U9176 (N_9176,N_868,N_772);
nand U9177 (N_9177,N_4142,N_4258);
or U9178 (N_9178,N_4402,N_2103);
nand U9179 (N_9179,N_3169,N_1154);
and U9180 (N_9180,N_256,N_1092);
nor U9181 (N_9181,N_4873,N_2838);
or U9182 (N_9182,N_1209,N_1816);
nor U9183 (N_9183,N_4166,N_1518);
nand U9184 (N_9184,N_3864,N_77);
nand U9185 (N_9185,N_952,N_1792);
nand U9186 (N_9186,N_1874,N_247);
nor U9187 (N_9187,N_1070,N_543);
nor U9188 (N_9188,N_4281,N_3769);
or U9189 (N_9189,N_467,N_1633);
nand U9190 (N_9190,N_976,N_1480);
nor U9191 (N_9191,N_2389,N_2962);
and U9192 (N_9192,N_3410,N_2221);
and U9193 (N_9193,N_812,N_4152);
or U9194 (N_9194,N_4681,N_457);
nor U9195 (N_9195,N_3298,N_3935);
and U9196 (N_9196,N_4056,N_4603);
nor U9197 (N_9197,N_73,N_4274);
or U9198 (N_9198,N_2145,N_4237);
or U9199 (N_9199,N_3331,N_1443);
and U9200 (N_9200,N_2634,N_3498);
or U9201 (N_9201,N_361,N_4835);
nor U9202 (N_9202,N_4435,N_3469);
and U9203 (N_9203,N_78,N_1741);
nand U9204 (N_9204,N_2300,N_4384);
or U9205 (N_9205,N_2533,N_3462);
or U9206 (N_9206,N_3871,N_3696);
or U9207 (N_9207,N_4572,N_1289);
xnor U9208 (N_9208,N_3679,N_913);
xnor U9209 (N_9209,N_1735,N_1720);
and U9210 (N_9210,N_3500,N_1477);
and U9211 (N_9211,N_2171,N_498);
or U9212 (N_9212,N_1744,N_676);
or U9213 (N_9213,N_4171,N_3204);
nor U9214 (N_9214,N_3913,N_1292);
or U9215 (N_9215,N_3030,N_2570);
and U9216 (N_9216,N_729,N_3385);
nor U9217 (N_9217,N_379,N_3005);
nor U9218 (N_9218,N_508,N_1232);
nor U9219 (N_9219,N_18,N_4993);
nand U9220 (N_9220,N_1999,N_3609);
nand U9221 (N_9221,N_857,N_2579);
nor U9222 (N_9222,N_1524,N_1978);
or U9223 (N_9223,N_3128,N_771);
and U9224 (N_9224,N_1644,N_2755);
nand U9225 (N_9225,N_1024,N_2867);
or U9226 (N_9226,N_4487,N_3504);
xnor U9227 (N_9227,N_4205,N_1239);
or U9228 (N_9228,N_2872,N_4480);
or U9229 (N_9229,N_4571,N_4890);
or U9230 (N_9230,N_2235,N_2908);
xor U9231 (N_9231,N_1926,N_2);
or U9232 (N_9232,N_41,N_3171);
and U9233 (N_9233,N_1518,N_3731);
nand U9234 (N_9234,N_2135,N_2675);
nor U9235 (N_9235,N_2839,N_813);
nor U9236 (N_9236,N_4453,N_4620);
and U9237 (N_9237,N_2390,N_2118);
or U9238 (N_9238,N_3513,N_3376);
nor U9239 (N_9239,N_2757,N_4932);
nor U9240 (N_9240,N_3995,N_3418);
nand U9241 (N_9241,N_2484,N_372);
nand U9242 (N_9242,N_2428,N_3611);
or U9243 (N_9243,N_3754,N_479);
nand U9244 (N_9244,N_2074,N_3019);
nor U9245 (N_9245,N_4302,N_2707);
nand U9246 (N_9246,N_45,N_2173);
nand U9247 (N_9247,N_2397,N_4471);
nand U9248 (N_9248,N_2716,N_3602);
nor U9249 (N_9249,N_438,N_2303);
and U9250 (N_9250,N_4952,N_3483);
nor U9251 (N_9251,N_4326,N_1144);
or U9252 (N_9252,N_296,N_4872);
or U9253 (N_9253,N_1257,N_3249);
or U9254 (N_9254,N_3903,N_3191);
or U9255 (N_9255,N_3070,N_2017);
nor U9256 (N_9256,N_1878,N_4733);
nand U9257 (N_9257,N_2770,N_4172);
nand U9258 (N_9258,N_2760,N_2931);
nor U9259 (N_9259,N_1650,N_1278);
or U9260 (N_9260,N_3581,N_4474);
nor U9261 (N_9261,N_1183,N_2056);
nand U9262 (N_9262,N_3006,N_1001);
nand U9263 (N_9263,N_2505,N_4986);
nand U9264 (N_9264,N_3028,N_2016);
and U9265 (N_9265,N_3666,N_2380);
nand U9266 (N_9266,N_1311,N_1280);
nor U9267 (N_9267,N_1911,N_1484);
and U9268 (N_9268,N_1092,N_1193);
and U9269 (N_9269,N_2008,N_1939);
or U9270 (N_9270,N_988,N_2766);
nor U9271 (N_9271,N_4242,N_1322);
nor U9272 (N_9272,N_2529,N_3112);
or U9273 (N_9273,N_3959,N_702);
nor U9274 (N_9274,N_3812,N_3601);
or U9275 (N_9275,N_3428,N_3974);
and U9276 (N_9276,N_2847,N_2334);
and U9277 (N_9277,N_600,N_4470);
nor U9278 (N_9278,N_1830,N_1070);
nand U9279 (N_9279,N_2184,N_4856);
xnor U9280 (N_9280,N_124,N_4822);
nand U9281 (N_9281,N_3199,N_4365);
and U9282 (N_9282,N_2915,N_4489);
nor U9283 (N_9283,N_4244,N_3790);
and U9284 (N_9284,N_4664,N_4364);
nor U9285 (N_9285,N_3311,N_3843);
and U9286 (N_9286,N_4990,N_3634);
and U9287 (N_9287,N_2465,N_2237);
or U9288 (N_9288,N_2626,N_2799);
nor U9289 (N_9289,N_2553,N_3723);
or U9290 (N_9290,N_3914,N_3014);
and U9291 (N_9291,N_4949,N_967);
or U9292 (N_9292,N_4183,N_2344);
nand U9293 (N_9293,N_483,N_2954);
nand U9294 (N_9294,N_669,N_814);
nor U9295 (N_9295,N_2045,N_2933);
and U9296 (N_9296,N_4219,N_3159);
nand U9297 (N_9297,N_4816,N_3154);
nand U9298 (N_9298,N_34,N_4758);
nand U9299 (N_9299,N_4315,N_3584);
nand U9300 (N_9300,N_4322,N_1340);
nand U9301 (N_9301,N_3748,N_3949);
and U9302 (N_9302,N_210,N_696);
nor U9303 (N_9303,N_1696,N_4465);
nor U9304 (N_9304,N_303,N_1218);
and U9305 (N_9305,N_4690,N_2951);
nand U9306 (N_9306,N_4969,N_2835);
nor U9307 (N_9307,N_1515,N_176);
nor U9308 (N_9308,N_3665,N_4928);
nor U9309 (N_9309,N_2543,N_459);
and U9310 (N_9310,N_4907,N_4304);
and U9311 (N_9311,N_1110,N_1135);
or U9312 (N_9312,N_1524,N_723);
nor U9313 (N_9313,N_4868,N_583);
or U9314 (N_9314,N_440,N_2319);
nand U9315 (N_9315,N_4784,N_15);
and U9316 (N_9316,N_4169,N_553);
xor U9317 (N_9317,N_510,N_105);
nand U9318 (N_9318,N_1197,N_908);
nand U9319 (N_9319,N_3721,N_4185);
nand U9320 (N_9320,N_2750,N_75);
nor U9321 (N_9321,N_2334,N_1246);
nand U9322 (N_9322,N_897,N_4838);
nor U9323 (N_9323,N_1086,N_138);
nand U9324 (N_9324,N_2804,N_1397);
nor U9325 (N_9325,N_2905,N_861);
or U9326 (N_9326,N_4782,N_4333);
or U9327 (N_9327,N_1073,N_4453);
nor U9328 (N_9328,N_1164,N_3412);
or U9329 (N_9329,N_566,N_1950);
nand U9330 (N_9330,N_498,N_1755);
or U9331 (N_9331,N_4126,N_2197);
and U9332 (N_9332,N_3004,N_1582);
nor U9333 (N_9333,N_780,N_2803);
nand U9334 (N_9334,N_4668,N_1346);
or U9335 (N_9335,N_1515,N_2452);
nand U9336 (N_9336,N_351,N_1272);
or U9337 (N_9337,N_1603,N_1874);
xor U9338 (N_9338,N_1958,N_1911);
nor U9339 (N_9339,N_3382,N_1628);
or U9340 (N_9340,N_4829,N_1998);
and U9341 (N_9341,N_3359,N_313);
xnor U9342 (N_9342,N_514,N_223);
or U9343 (N_9343,N_1949,N_3422);
or U9344 (N_9344,N_2077,N_4168);
or U9345 (N_9345,N_2202,N_1584);
nor U9346 (N_9346,N_4472,N_4267);
or U9347 (N_9347,N_276,N_3673);
nand U9348 (N_9348,N_1631,N_4778);
or U9349 (N_9349,N_2958,N_4717);
and U9350 (N_9350,N_1012,N_2644);
and U9351 (N_9351,N_1893,N_1561);
nand U9352 (N_9352,N_4400,N_1820);
or U9353 (N_9353,N_1444,N_4470);
or U9354 (N_9354,N_4223,N_553);
nand U9355 (N_9355,N_1281,N_4953);
nand U9356 (N_9356,N_928,N_4159);
nor U9357 (N_9357,N_4858,N_1356);
and U9358 (N_9358,N_3487,N_4929);
nor U9359 (N_9359,N_933,N_3390);
and U9360 (N_9360,N_1107,N_2006);
nor U9361 (N_9361,N_706,N_2023);
nor U9362 (N_9362,N_1598,N_42);
nor U9363 (N_9363,N_601,N_3505);
nor U9364 (N_9364,N_704,N_945);
and U9365 (N_9365,N_3634,N_2781);
and U9366 (N_9366,N_2221,N_762);
or U9367 (N_9367,N_4018,N_4041);
and U9368 (N_9368,N_2341,N_922);
and U9369 (N_9369,N_691,N_3093);
nand U9370 (N_9370,N_4155,N_523);
nand U9371 (N_9371,N_2434,N_653);
nand U9372 (N_9372,N_4992,N_2366);
and U9373 (N_9373,N_1616,N_4687);
nor U9374 (N_9374,N_2064,N_3525);
nor U9375 (N_9375,N_3376,N_672);
or U9376 (N_9376,N_4174,N_3527);
and U9377 (N_9377,N_387,N_4977);
nor U9378 (N_9378,N_3789,N_84);
and U9379 (N_9379,N_426,N_4337);
nand U9380 (N_9380,N_4399,N_1720);
nor U9381 (N_9381,N_1062,N_436);
nand U9382 (N_9382,N_4596,N_988);
nand U9383 (N_9383,N_4654,N_1239);
and U9384 (N_9384,N_942,N_3450);
or U9385 (N_9385,N_3707,N_4741);
and U9386 (N_9386,N_903,N_340);
nor U9387 (N_9387,N_2979,N_2817);
and U9388 (N_9388,N_4347,N_2541);
and U9389 (N_9389,N_174,N_4374);
nand U9390 (N_9390,N_4186,N_1212);
nand U9391 (N_9391,N_3361,N_1824);
nor U9392 (N_9392,N_303,N_3843);
and U9393 (N_9393,N_3768,N_3677);
or U9394 (N_9394,N_4590,N_1581);
or U9395 (N_9395,N_4107,N_3041);
nor U9396 (N_9396,N_3184,N_2343);
xor U9397 (N_9397,N_3733,N_3104);
or U9398 (N_9398,N_1126,N_1418);
nor U9399 (N_9399,N_660,N_2366);
and U9400 (N_9400,N_4730,N_71);
nor U9401 (N_9401,N_3829,N_2566);
and U9402 (N_9402,N_1683,N_4065);
or U9403 (N_9403,N_2022,N_2527);
or U9404 (N_9404,N_2636,N_3666);
and U9405 (N_9405,N_3441,N_3300);
nor U9406 (N_9406,N_3402,N_2252);
and U9407 (N_9407,N_3211,N_4596);
nand U9408 (N_9408,N_3805,N_3678);
and U9409 (N_9409,N_3129,N_3525);
nand U9410 (N_9410,N_1821,N_583);
nor U9411 (N_9411,N_751,N_1331);
or U9412 (N_9412,N_3777,N_3535);
or U9413 (N_9413,N_4390,N_1533);
or U9414 (N_9414,N_4717,N_2462);
nand U9415 (N_9415,N_3923,N_900);
xor U9416 (N_9416,N_225,N_1115);
nand U9417 (N_9417,N_4335,N_135);
nor U9418 (N_9418,N_3278,N_2810);
and U9419 (N_9419,N_3002,N_1860);
xor U9420 (N_9420,N_3014,N_4630);
nor U9421 (N_9421,N_692,N_666);
nor U9422 (N_9422,N_1769,N_1687);
nand U9423 (N_9423,N_4433,N_521);
and U9424 (N_9424,N_3910,N_4272);
and U9425 (N_9425,N_1172,N_1534);
xor U9426 (N_9426,N_2042,N_1469);
and U9427 (N_9427,N_2636,N_3622);
and U9428 (N_9428,N_2680,N_4059);
and U9429 (N_9429,N_1096,N_4536);
or U9430 (N_9430,N_256,N_2551);
and U9431 (N_9431,N_2809,N_1214);
and U9432 (N_9432,N_1965,N_1525);
or U9433 (N_9433,N_3371,N_387);
nor U9434 (N_9434,N_3376,N_3132);
and U9435 (N_9435,N_947,N_4433);
and U9436 (N_9436,N_1226,N_1707);
nand U9437 (N_9437,N_2964,N_2909);
nand U9438 (N_9438,N_2234,N_3840);
nor U9439 (N_9439,N_3554,N_2684);
or U9440 (N_9440,N_2256,N_4428);
or U9441 (N_9441,N_3735,N_1192);
and U9442 (N_9442,N_2503,N_4172);
or U9443 (N_9443,N_4238,N_3828);
nor U9444 (N_9444,N_3388,N_3238);
nor U9445 (N_9445,N_4634,N_4881);
xor U9446 (N_9446,N_149,N_1472);
nor U9447 (N_9447,N_4454,N_371);
and U9448 (N_9448,N_2599,N_3068);
and U9449 (N_9449,N_545,N_1713);
nor U9450 (N_9450,N_2987,N_3657);
nor U9451 (N_9451,N_4575,N_1901);
nor U9452 (N_9452,N_1410,N_1347);
and U9453 (N_9453,N_449,N_2436);
and U9454 (N_9454,N_3165,N_664);
nor U9455 (N_9455,N_3638,N_2630);
nand U9456 (N_9456,N_86,N_2376);
nor U9457 (N_9457,N_4340,N_2646);
or U9458 (N_9458,N_3621,N_76);
nor U9459 (N_9459,N_2465,N_767);
nand U9460 (N_9460,N_1135,N_4779);
or U9461 (N_9461,N_4807,N_2614);
and U9462 (N_9462,N_3611,N_2325);
and U9463 (N_9463,N_1200,N_647);
nor U9464 (N_9464,N_3259,N_1097);
or U9465 (N_9465,N_108,N_3650);
and U9466 (N_9466,N_1126,N_1955);
and U9467 (N_9467,N_4686,N_2090);
nand U9468 (N_9468,N_4191,N_4241);
nor U9469 (N_9469,N_2330,N_1555);
nor U9470 (N_9470,N_1741,N_4013);
nand U9471 (N_9471,N_4914,N_2364);
nor U9472 (N_9472,N_2695,N_4511);
nor U9473 (N_9473,N_8,N_3465);
nor U9474 (N_9474,N_1517,N_1027);
nor U9475 (N_9475,N_2430,N_4238);
nand U9476 (N_9476,N_3828,N_4288);
nand U9477 (N_9477,N_3890,N_4827);
or U9478 (N_9478,N_4912,N_3333);
nor U9479 (N_9479,N_4088,N_4443);
nand U9480 (N_9480,N_2206,N_4100);
and U9481 (N_9481,N_4669,N_3579);
nor U9482 (N_9482,N_1751,N_3436);
and U9483 (N_9483,N_1506,N_496);
or U9484 (N_9484,N_1817,N_2033);
nand U9485 (N_9485,N_3968,N_4816);
or U9486 (N_9486,N_4161,N_3918);
or U9487 (N_9487,N_861,N_4878);
or U9488 (N_9488,N_3970,N_927);
and U9489 (N_9489,N_4309,N_3627);
nor U9490 (N_9490,N_2003,N_2387);
nor U9491 (N_9491,N_515,N_3729);
nor U9492 (N_9492,N_1636,N_80);
or U9493 (N_9493,N_640,N_2338);
and U9494 (N_9494,N_2421,N_2336);
nand U9495 (N_9495,N_1895,N_1732);
and U9496 (N_9496,N_2838,N_1596);
or U9497 (N_9497,N_3838,N_3819);
nor U9498 (N_9498,N_1594,N_745);
nand U9499 (N_9499,N_2130,N_1781);
nand U9500 (N_9500,N_2125,N_4668);
xnor U9501 (N_9501,N_986,N_1571);
nand U9502 (N_9502,N_2633,N_4601);
nand U9503 (N_9503,N_2062,N_2712);
nand U9504 (N_9504,N_3532,N_372);
and U9505 (N_9505,N_4159,N_3843);
nor U9506 (N_9506,N_916,N_134);
and U9507 (N_9507,N_1380,N_4253);
nor U9508 (N_9508,N_585,N_2021);
nand U9509 (N_9509,N_1018,N_1242);
and U9510 (N_9510,N_1974,N_2765);
or U9511 (N_9511,N_1040,N_506);
or U9512 (N_9512,N_994,N_3276);
or U9513 (N_9513,N_3944,N_3083);
nor U9514 (N_9514,N_1438,N_3010);
or U9515 (N_9515,N_934,N_1968);
nand U9516 (N_9516,N_2439,N_2510);
and U9517 (N_9517,N_2732,N_461);
nor U9518 (N_9518,N_2491,N_1968);
nand U9519 (N_9519,N_4483,N_1522);
nor U9520 (N_9520,N_3017,N_4177);
nor U9521 (N_9521,N_1321,N_2573);
nand U9522 (N_9522,N_4896,N_1900);
nor U9523 (N_9523,N_1819,N_4652);
nor U9524 (N_9524,N_4177,N_2659);
and U9525 (N_9525,N_849,N_4395);
nor U9526 (N_9526,N_3139,N_4902);
and U9527 (N_9527,N_278,N_2688);
nor U9528 (N_9528,N_1784,N_4428);
nand U9529 (N_9529,N_1390,N_3571);
nand U9530 (N_9530,N_1533,N_1742);
and U9531 (N_9531,N_3361,N_347);
nor U9532 (N_9532,N_1466,N_4944);
and U9533 (N_9533,N_2160,N_1469);
and U9534 (N_9534,N_3999,N_872);
and U9535 (N_9535,N_256,N_4455);
nor U9536 (N_9536,N_4852,N_3259);
nor U9537 (N_9537,N_2077,N_4241);
nor U9538 (N_9538,N_1106,N_4498);
nor U9539 (N_9539,N_3792,N_1393);
or U9540 (N_9540,N_3111,N_3312);
or U9541 (N_9541,N_2723,N_1418);
nor U9542 (N_9542,N_2493,N_2891);
nor U9543 (N_9543,N_3941,N_3458);
and U9544 (N_9544,N_512,N_4790);
or U9545 (N_9545,N_955,N_1721);
or U9546 (N_9546,N_173,N_767);
nand U9547 (N_9547,N_4392,N_2105);
or U9548 (N_9548,N_2360,N_1544);
and U9549 (N_9549,N_2070,N_2014);
or U9550 (N_9550,N_2289,N_231);
nand U9551 (N_9551,N_4867,N_3119);
and U9552 (N_9552,N_1091,N_4636);
nor U9553 (N_9553,N_3198,N_1295);
nor U9554 (N_9554,N_1156,N_4539);
nor U9555 (N_9555,N_1419,N_2095);
nor U9556 (N_9556,N_4674,N_4481);
and U9557 (N_9557,N_4920,N_831);
nor U9558 (N_9558,N_4901,N_3016);
nand U9559 (N_9559,N_1556,N_696);
or U9560 (N_9560,N_2441,N_2380);
and U9561 (N_9561,N_3825,N_4744);
and U9562 (N_9562,N_3226,N_1307);
and U9563 (N_9563,N_3035,N_4554);
nor U9564 (N_9564,N_4387,N_239);
and U9565 (N_9565,N_1491,N_4401);
nor U9566 (N_9566,N_3618,N_1407);
or U9567 (N_9567,N_1109,N_4141);
or U9568 (N_9568,N_353,N_212);
or U9569 (N_9569,N_1516,N_4219);
nor U9570 (N_9570,N_1701,N_250);
nor U9571 (N_9571,N_3920,N_4312);
nand U9572 (N_9572,N_4086,N_3933);
nand U9573 (N_9573,N_3173,N_4997);
nor U9574 (N_9574,N_2494,N_3645);
or U9575 (N_9575,N_3494,N_2758);
and U9576 (N_9576,N_2836,N_665);
nor U9577 (N_9577,N_1722,N_1609);
nor U9578 (N_9578,N_2745,N_96);
nand U9579 (N_9579,N_2744,N_3442);
nand U9580 (N_9580,N_1713,N_3044);
or U9581 (N_9581,N_1604,N_3877);
nor U9582 (N_9582,N_557,N_2093);
nand U9583 (N_9583,N_3911,N_818);
nand U9584 (N_9584,N_914,N_3156);
nor U9585 (N_9585,N_913,N_1059);
nor U9586 (N_9586,N_3582,N_1691);
nand U9587 (N_9587,N_3577,N_2258);
or U9588 (N_9588,N_3499,N_1453);
nor U9589 (N_9589,N_1418,N_998);
nand U9590 (N_9590,N_3415,N_2892);
nand U9591 (N_9591,N_2590,N_1799);
or U9592 (N_9592,N_4545,N_3836);
nand U9593 (N_9593,N_3624,N_4730);
nor U9594 (N_9594,N_2123,N_3196);
and U9595 (N_9595,N_1563,N_3249);
or U9596 (N_9596,N_361,N_3549);
nor U9597 (N_9597,N_4973,N_3456);
nand U9598 (N_9598,N_1690,N_4315);
and U9599 (N_9599,N_1599,N_3007);
nor U9600 (N_9600,N_1541,N_3161);
and U9601 (N_9601,N_31,N_791);
nand U9602 (N_9602,N_717,N_1994);
nor U9603 (N_9603,N_2686,N_4085);
nor U9604 (N_9604,N_2853,N_780);
nand U9605 (N_9605,N_3470,N_2126);
and U9606 (N_9606,N_1758,N_2393);
nand U9607 (N_9607,N_1931,N_4973);
and U9608 (N_9608,N_1199,N_3550);
nor U9609 (N_9609,N_1821,N_3615);
and U9610 (N_9610,N_3317,N_3378);
nand U9611 (N_9611,N_3287,N_2578);
and U9612 (N_9612,N_2756,N_4559);
nor U9613 (N_9613,N_1795,N_332);
nand U9614 (N_9614,N_4615,N_685);
or U9615 (N_9615,N_3279,N_1800);
and U9616 (N_9616,N_1465,N_1882);
or U9617 (N_9617,N_1399,N_4475);
and U9618 (N_9618,N_124,N_4471);
and U9619 (N_9619,N_1660,N_316);
nand U9620 (N_9620,N_1950,N_3496);
or U9621 (N_9621,N_2846,N_3219);
nand U9622 (N_9622,N_3682,N_4898);
and U9623 (N_9623,N_3953,N_3426);
nor U9624 (N_9624,N_3298,N_705);
and U9625 (N_9625,N_4722,N_4117);
nand U9626 (N_9626,N_1039,N_323);
or U9627 (N_9627,N_4718,N_3958);
or U9628 (N_9628,N_4288,N_3223);
nor U9629 (N_9629,N_2711,N_4476);
nor U9630 (N_9630,N_181,N_3038);
and U9631 (N_9631,N_3368,N_4575);
nor U9632 (N_9632,N_2430,N_4909);
or U9633 (N_9633,N_2438,N_543);
nand U9634 (N_9634,N_4435,N_2984);
nand U9635 (N_9635,N_1437,N_196);
xor U9636 (N_9636,N_1114,N_2344);
and U9637 (N_9637,N_4176,N_2060);
or U9638 (N_9638,N_3439,N_4206);
and U9639 (N_9639,N_1,N_562);
and U9640 (N_9640,N_3918,N_1780);
or U9641 (N_9641,N_1480,N_4892);
nor U9642 (N_9642,N_564,N_342);
nor U9643 (N_9643,N_2281,N_4526);
or U9644 (N_9644,N_2932,N_254);
and U9645 (N_9645,N_1939,N_1293);
nor U9646 (N_9646,N_3868,N_808);
nand U9647 (N_9647,N_33,N_43);
nor U9648 (N_9648,N_4799,N_4325);
and U9649 (N_9649,N_3393,N_3059);
xnor U9650 (N_9650,N_4833,N_1581);
and U9651 (N_9651,N_2800,N_626);
nor U9652 (N_9652,N_1720,N_2390);
or U9653 (N_9653,N_107,N_1083);
nor U9654 (N_9654,N_2263,N_1658);
and U9655 (N_9655,N_1507,N_1588);
nor U9656 (N_9656,N_4439,N_2536);
nand U9657 (N_9657,N_1876,N_2692);
nand U9658 (N_9658,N_2339,N_44);
and U9659 (N_9659,N_805,N_4957);
nand U9660 (N_9660,N_3049,N_1463);
and U9661 (N_9661,N_2002,N_3799);
nor U9662 (N_9662,N_3984,N_4683);
nand U9663 (N_9663,N_1222,N_1832);
nand U9664 (N_9664,N_1215,N_2302);
nor U9665 (N_9665,N_3499,N_3429);
xor U9666 (N_9666,N_3586,N_2039);
xnor U9667 (N_9667,N_819,N_4762);
nor U9668 (N_9668,N_2104,N_4304);
or U9669 (N_9669,N_3229,N_2097);
and U9670 (N_9670,N_802,N_4334);
or U9671 (N_9671,N_3737,N_966);
and U9672 (N_9672,N_3684,N_1531);
and U9673 (N_9673,N_2304,N_3017);
nor U9674 (N_9674,N_4779,N_2066);
nand U9675 (N_9675,N_1640,N_1617);
or U9676 (N_9676,N_3521,N_4643);
or U9677 (N_9677,N_1963,N_245);
or U9678 (N_9678,N_1801,N_4335);
or U9679 (N_9679,N_2837,N_2442);
and U9680 (N_9680,N_319,N_3530);
nor U9681 (N_9681,N_231,N_1499);
nor U9682 (N_9682,N_2685,N_2585);
and U9683 (N_9683,N_2205,N_1929);
or U9684 (N_9684,N_3406,N_430);
and U9685 (N_9685,N_1662,N_2903);
or U9686 (N_9686,N_2182,N_1230);
and U9687 (N_9687,N_4252,N_514);
xnor U9688 (N_9688,N_2596,N_4633);
or U9689 (N_9689,N_2515,N_2425);
or U9690 (N_9690,N_1271,N_4076);
or U9691 (N_9691,N_1505,N_213);
and U9692 (N_9692,N_4823,N_12);
and U9693 (N_9693,N_147,N_4226);
nand U9694 (N_9694,N_783,N_3084);
and U9695 (N_9695,N_1245,N_301);
or U9696 (N_9696,N_2106,N_3841);
nor U9697 (N_9697,N_2913,N_729);
or U9698 (N_9698,N_4716,N_237);
nor U9699 (N_9699,N_1438,N_1495);
and U9700 (N_9700,N_3606,N_895);
nand U9701 (N_9701,N_184,N_4860);
nand U9702 (N_9702,N_4297,N_1293);
and U9703 (N_9703,N_1289,N_2729);
nor U9704 (N_9704,N_2671,N_791);
nor U9705 (N_9705,N_1131,N_1962);
and U9706 (N_9706,N_2268,N_4156);
and U9707 (N_9707,N_334,N_636);
nand U9708 (N_9708,N_237,N_2637);
nor U9709 (N_9709,N_4293,N_1783);
and U9710 (N_9710,N_2983,N_439);
and U9711 (N_9711,N_2630,N_181);
and U9712 (N_9712,N_735,N_2662);
nor U9713 (N_9713,N_3003,N_1315);
nor U9714 (N_9714,N_4726,N_2161);
or U9715 (N_9715,N_136,N_757);
and U9716 (N_9716,N_739,N_3792);
or U9717 (N_9717,N_4019,N_3027);
nor U9718 (N_9718,N_1888,N_3);
and U9719 (N_9719,N_1869,N_3817);
and U9720 (N_9720,N_4569,N_3675);
or U9721 (N_9721,N_850,N_4706);
nand U9722 (N_9722,N_2367,N_3990);
and U9723 (N_9723,N_3531,N_1851);
and U9724 (N_9724,N_2513,N_2610);
nor U9725 (N_9725,N_1823,N_2355);
nand U9726 (N_9726,N_1641,N_3450);
or U9727 (N_9727,N_3249,N_4928);
nor U9728 (N_9728,N_4524,N_659);
xor U9729 (N_9729,N_941,N_4977);
and U9730 (N_9730,N_2796,N_2197);
nand U9731 (N_9731,N_2484,N_235);
or U9732 (N_9732,N_4628,N_4060);
nand U9733 (N_9733,N_4690,N_1332);
or U9734 (N_9734,N_2379,N_4141);
or U9735 (N_9735,N_469,N_4157);
and U9736 (N_9736,N_3841,N_4872);
nor U9737 (N_9737,N_1163,N_1287);
nor U9738 (N_9738,N_2962,N_743);
and U9739 (N_9739,N_2105,N_1523);
or U9740 (N_9740,N_4913,N_4071);
nand U9741 (N_9741,N_949,N_2143);
and U9742 (N_9742,N_3205,N_1515);
nand U9743 (N_9743,N_3504,N_4507);
or U9744 (N_9744,N_2564,N_380);
nand U9745 (N_9745,N_721,N_1555);
and U9746 (N_9746,N_3833,N_3345);
nor U9747 (N_9747,N_2005,N_1565);
nand U9748 (N_9748,N_1972,N_2327);
xnor U9749 (N_9749,N_3494,N_4779);
and U9750 (N_9750,N_1293,N_555);
nand U9751 (N_9751,N_882,N_2467);
nand U9752 (N_9752,N_3946,N_2433);
nand U9753 (N_9753,N_3867,N_2934);
nor U9754 (N_9754,N_3299,N_827);
or U9755 (N_9755,N_1823,N_971);
and U9756 (N_9756,N_3699,N_62);
nand U9757 (N_9757,N_3613,N_1990);
or U9758 (N_9758,N_4917,N_1543);
or U9759 (N_9759,N_1416,N_4789);
or U9760 (N_9760,N_4353,N_2848);
nand U9761 (N_9761,N_1522,N_1347);
and U9762 (N_9762,N_2941,N_3318);
and U9763 (N_9763,N_640,N_2180);
nor U9764 (N_9764,N_3936,N_31);
and U9765 (N_9765,N_1854,N_4294);
nor U9766 (N_9766,N_366,N_3651);
xor U9767 (N_9767,N_2439,N_3978);
or U9768 (N_9768,N_4896,N_3104);
or U9769 (N_9769,N_2141,N_1312);
or U9770 (N_9770,N_2944,N_1126);
nand U9771 (N_9771,N_439,N_978);
and U9772 (N_9772,N_2521,N_2176);
and U9773 (N_9773,N_3887,N_2162);
or U9774 (N_9774,N_1586,N_1261);
or U9775 (N_9775,N_333,N_3648);
nand U9776 (N_9776,N_642,N_9);
and U9777 (N_9777,N_3980,N_3573);
and U9778 (N_9778,N_4055,N_526);
and U9779 (N_9779,N_2761,N_4967);
nor U9780 (N_9780,N_4760,N_3313);
nand U9781 (N_9781,N_3696,N_1378);
or U9782 (N_9782,N_1214,N_3334);
or U9783 (N_9783,N_1483,N_3890);
nand U9784 (N_9784,N_559,N_2575);
nand U9785 (N_9785,N_1446,N_1474);
nand U9786 (N_9786,N_4768,N_1998);
nand U9787 (N_9787,N_1572,N_181);
nor U9788 (N_9788,N_4273,N_1071);
nor U9789 (N_9789,N_854,N_1140);
and U9790 (N_9790,N_2701,N_3240);
or U9791 (N_9791,N_410,N_4536);
nand U9792 (N_9792,N_4056,N_973);
and U9793 (N_9793,N_116,N_2616);
nor U9794 (N_9794,N_2573,N_945);
or U9795 (N_9795,N_4150,N_3975);
and U9796 (N_9796,N_1024,N_2418);
nor U9797 (N_9797,N_4211,N_675);
nand U9798 (N_9798,N_103,N_4143);
nand U9799 (N_9799,N_2938,N_2680);
nor U9800 (N_9800,N_285,N_4394);
nor U9801 (N_9801,N_3679,N_2427);
and U9802 (N_9802,N_232,N_2339);
nand U9803 (N_9803,N_3678,N_1801);
or U9804 (N_9804,N_3807,N_116);
and U9805 (N_9805,N_2745,N_1368);
and U9806 (N_9806,N_3094,N_944);
nand U9807 (N_9807,N_203,N_1772);
and U9808 (N_9808,N_1509,N_31);
xor U9809 (N_9809,N_4994,N_984);
and U9810 (N_9810,N_581,N_4861);
nand U9811 (N_9811,N_460,N_2837);
or U9812 (N_9812,N_277,N_3397);
and U9813 (N_9813,N_1070,N_3982);
nor U9814 (N_9814,N_3420,N_1376);
nor U9815 (N_9815,N_3947,N_592);
and U9816 (N_9816,N_2576,N_2673);
nor U9817 (N_9817,N_1495,N_3402);
nor U9818 (N_9818,N_2005,N_2342);
nor U9819 (N_9819,N_3648,N_689);
nand U9820 (N_9820,N_678,N_1997);
and U9821 (N_9821,N_1156,N_2947);
nand U9822 (N_9822,N_3277,N_3335);
nand U9823 (N_9823,N_206,N_2869);
nor U9824 (N_9824,N_4270,N_4722);
or U9825 (N_9825,N_3808,N_3843);
xnor U9826 (N_9826,N_735,N_1695);
nor U9827 (N_9827,N_248,N_2156);
or U9828 (N_9828,N_1860,N_129);
nor U9829 (N_9829,N_4390,N_4852);
nand U9830 (N_9830,N_2075,N_4065);
nor U9831 (N_9831,N_4869,N_1350);
nor U9832 (N_9832,N_375,N_1495);
nor U9833 (N_9833,N_1678,N_2885);
or U9834 (N_9834,N_4621,N_4738);
nand U9835 (N_9835,N_25,N_2913);
or U9836 (N_9836,N_2147,N_4761);
nor U9837 (N_9837,N_3178,N_1264);
nand U9838 (N_9838,N_4905,N_2603);
nor U9839 (N_9839,N_4887,N_2015);
or U9840 (N_9840,N_489,N_643);
and U9841 (N_9841,N_550,N_3294);
nand U9842 (N_9842,N_4812,N_4739);
nor U9843 (N_9843,N_2062,N_1300);
nor U9844 (N_9844,N_188,N_321);
nand U9845 (N_9845,N_456,N_172);
nor U9846 (N_9846,N_2975,N_3287);
nand U9847 (N_9847,N_1900,N_4903);
nand U9848 (N_9848,N_335,N_1562);
nor U9849 (N_9849,N_564,N_3562);
or U9850 (N_9850,N_294,N_1282);
or U9851 (N_9851,N_2320,N_833);
nand U9852 (N_9852,N_3383,N_3033);
nand U9853 (N_9853,N_205,N_859);
and U9854 (N_9854,N_3822,N_4780);
nor U9855 (N_9855,N_2045,N_2367);
and U9856 (N_9856,N_2275,N_4969);
nand U9857 (N_9857,N_1687,N_209);
and U9858 (N_9858,N_3707,N_4547);
nor U9859 (N_9859,N_979,N_3864);
nor U9860 (N_9860,N_2650,N_4809);
nand U9861 (N_9861,N_2005,N_1707);
nor U9862 (N_9862,N_127,N_4964);
xnor U9863 (N_9863,N_1196,N_1244);
nor U9864 (N_9864,N_4169,N_3403);
nor U9865 (N_9865,N_2928,N_3850);
nor U9866 (N_9866,N_3852,N_3499);
and U9867 (N_9867,N_2236,N_4824);
nor U9868 (N_9868,N_3532,N_4300);
nor U9869 (N_9869,N_2592,N_473);
and U9870 (N_9870,N_256,N_3507);
and U9871 (N_9871,N_2227,N_4015);
nor U9872 (N_9872,N_3509,N_4696);
nand U9873 (N_9873,N_3179,N_3945);
nor U9874 (N_9874,N_4991,N_4726);
and U9875 (N_9875,N_3517,N_3513);
or U9876 (N_9876,N_3091,N_2767);
and U9877 (N_9877,N_2045,N_2593);
and U9878 (N_9878,N_2679,N_2348);
and U9879 (N_9879,N_2846,N_699);
and U9880 (N_9880,N_2418,N_4226);
nand U9881 (N_9881,N_1854,N_2779);
nand U9882 (N_9882,N_745,N_2306);
nand U9883 (N_9883,N_1997,N_4223);
or U9884 (N_9884,N_4482,N_3250);
or U9885 (N_9885,N_4315,N_3282);
nand U9886 (N_9886,N_558,N_1787);
or U9887 (N_9887,N_415,N_3117);
nor U9888 (N_9888,N_4842,N_596);
or U9889 (N_9889,N_1584,N_2973);
and U9890 (N_9890,N_3370,N_2676);
or U9891 (N_9891,N_4505,N_106);
nand U9892 (N_9892,N_1966,N_3878);
xor U9893 (N_9893,N_2384,N_2893);
and U9894 (N_9894,N_853,N_513);
and U9895 (N_9895,N_2234,N_2937);
nand U9896 (N_9896,N_2965,N_1937);
and U9897 (N_9897,N_2802,N_3898);
nor U9898 (N_9898,N_3013,N_2085);
nor U9899 (N_9899,N_3250,N_626);
and U9900 (N_9900,N_742,N_2010);
nand U9901 (N_9901,N_1859,N_1527);
and U9902 (N_9902,N_4790,N_4078);
nand U9903 (N_9903,N_4610,N_971);
or U9904 (N_9904,N_97,N_3347);
or U9905 (N_9905,N_1589,N_1913);
nand U9906 (N_9906,N_3208,N_588);
or U9907 (N_9907,N_1495,N_1445);
nand U9908 (N_9908,N_2136,N_3206);
or U9909 (N_9909,N_76,N_1226);
and U9910 (N_9910,N_3983,N_1081);
nand U9911 (N_9911,N_2030,N_3798);
nor U9912 (N_9912,N_2538,N_2442);
nand U9913 (N_9913,N_2934,N_4763);
nor U9914 (N_9914,N_1027,N_3575);
or U9915 (N_9915,N_2810,N_3900);
and U9916 (N_9916,N_171,N_4754);
or U9917 (N_9917,N_3794,N_1115);
or U9918 (N_9918,N_514,N_4607);
or U9919 (N_9919,N_4028,N_4862);
and U9920 (N_9920,N_2809,N_4663);
nand U9921 (N_9921,N_3886,N_959);
nor U9922 (N_9922,N_1043,N_2739);
nor U9923 (N_9923,N_2348,N_318);
nand U9924 (N_9924,N_2944,N_3180);
or U9925 (N_9925,N_681,N_1034);
nor U9926 (N_9926,N_4902,N_4912);
or U9927 (N_9927,N_4624,N_1778);
nor U9928 (N_9928,N_1570,N_3739);
xnor U9929 (N_9929,N_1649,N_146);
nor U9930 (N_9930,N_2991,N_4284);
and U9931 (N_9931,N_2448,N_1151);
and U9932 (N_9932,N_2550,N_2673);
nand U9933 (N_9933,N_3775,N_17);
or U9934 (N_9934,N_4096,N_4996);
nor U9935 (N_9935,N_4041,N_4680);
or U9936 (N_9936,N_947,N_1457);
nor U9937 (N_9937,N_3033,N_3498);
and U9938 (N_9938,N_4162,N_500);
nand U9939 (N_9939,N_3467,N_1316);
nand U9940 (N_9940,N_808,N_2106);
or U9941 (N_9941,N_4133,N_1950);
nand U9942 (N_9942,N_2006,N_3789);
or U9943 (N_9943,N_4027,N_3763);
nand U9944 (N_9944,N_4802,N_4861);
nand U9945 (N_9945,N_1292,N_1958);
nand U9946 (N_9946,N_3750,N_1708);
and U9947 (N_9947,N_4251,N_1805);
nand U9948 (N_9948,N_2268,N_3019);
nor U9949 (N_9949,N_2495,N_82);
or U9950 (N_9950,N_4923,N_1940);
nor U9951 (N_9951,N_2520,N_3534);
nor U9952 (N_9952,N_699,N_514);
nand U9953 (N_9953,N_1013,N_3509);
and U9954 (N_9954,N_4393,N_3727);
nand U9955 (N_9955,N_675,N_0);
nand U9956 (N_9956,N_997,N_3599);
or U9957 (N_9957,N_279,N_564);
nor U9958 (N_9958,N_223,N_463);
nand U9959 (N_9959,N_4889,N_2996);
nor U9960 (N_9960,N_1936,N_3451);
and U9961 (N_9961,N_4560,N_4072);
nand U9962 (N_9962,N_4535,N_2698);
or U9963 (N_9963,N_1942,N_4193);
nand U9964 (N_9964,N_2082,N_3034);
or U9965 (N_9965,N_4780,N_3720);
nand U9966 (N_9966,N_4802,N_484);
nor U9967 (N_9967,N_4448,N_3833);
and U9968 (N_9968,N_817,N_3972);
nor U9969 (N_9969,N_3791,N_4119);
nand U9970 (N_9970,N_4819,N_4071);
nor U9971 (N_9971,N_3880,N_403);
xor U9972 (N_9972,N_2307,N_1485);
and U9973 (N_9973,N_2127,N_1153);
and U9974 (N_9974,N_1549,N_71);
or U9975 (N_9975,N_964,N_2594);
xor U9976 (N_9976,N_3053,N_688);
or U9977 (N_9977,N_1016,N_4024);
nor U9978 (N_9978,N_872,N_2545);
or U9979 (N_9979,N_2395,N_1559);
nand U9980 (N_9980,N_3436,N_4934);
nor U9981 (N_9981,N_3466,N_1634);
nand U9982 (N_9982,N_4794,N_1025);
nor U9983 (N_9983,N_2383,N_4533);
or U9984 (N_9984,N_531,N_3068);
and U9985 (N_9985,N_3196,N_2333);
nor U9986 (N_9986,N_4664,N_2634);
nand U9987 (N_9987,N_1028,N_1739);
and U9988 (N_9988,N_4273,N_1776);
nor U9989 (N_9989,N_1663,N_4093);
and U9990 (N_9990,N_1062,N_1781);
nor U9991 (N_9991,N_2538,N_692);
nor U9992 (N_9992,N_1119,N_1967);
and U9993 (N_9993,N_2719,N_432);
nor U9994 (N_9994,N_3108,N_2843);
and U9995 (N_9995,N_4471,N_756);
nor U9996 (N_9996,N_784,N_1625);
nor U9997 (N_9997,N_2672,N_1226);
nand U9998 (N_9998,N_4145,N_4167);
nor U9999 (N_9999,N_3016,N_494);
xnor U10000 (N_10000,N_9449,N_7659);
or U10001 (N_10001,N_8138,N_5520);
xor U10002 (N_10002,N_6494,N_7220);
nor U10003 (N_10003,N_9152,N_9170);
nor U10004 (N_10004,N_7988,N_9600);
nand U10005 (N_10005,N_8856,N_5625);
or U10006 (N_10006,N_7528,N_7827);
nand U10007 (N_10007,N_8376,N_7752);
xnor U10008 (N_10008,N_6285,N_6347);
nand U10009 (N_10009,N_5858,N_5422);
nor U10010 (N_10010,N_6114,N_8105);
nor U10011 (N_10011,N_9958,N_9935);
or U10012 (N_10012,N_5577,N_8194);
nand U10013 (N_10013,N_7694,N_5897);
and U10014 (N_10014,N_5549,N_6062);
and U10015 (N_10015,N_5782,N_9862);
and U10016 (N_10016,N_5586,N_8555);
or U10017 (N_10017,N_5256,N_9256);
or U10018 (N_10018,N_5127,N_7262);
nand U10019 (N_10019,N_8979,N_7840);
and U10020 (N_10020,N_9881,N_7045);
nor U10021 (N_10021,N_5132,N_8364);
nor U10022 (N_10022,N_8304,N_7065);
nand U10023 (N_10023,N_9114,N_5995);
and U10024 (N_10024,N_5458,N_9988);
or U10025 (N_10025,N_6903,N_5922);
nand U10026 (N_10026,N_8295,N_6230);
nand U10027 (N_10027,N_8183,N_8581);
nor U10028 (N_10028,N_8539,N_8523);
nand U10029 (N_10029,N_9052,N_5450);
and U10030 (N_10030,N_8245,N_9489);
and U10031 (N_10031,N_9482,N_5065);
xnor U10032 (N_10032,N_9488,N_6605);
nor U10033 (N_10033,N_9897,N_7655);
or U10034 (N_10034,N_9984,N_8877);
and U10035 (N_10035,N_8641,N_6514);
nand U10036 (N_10036,N_9300,N_5423);
nand U10037 (N_10037,N_9993,N_8862);
or U10038 (N_10038,N_5654,N_9512);
or U10039 (N_10039,N_6104,N_6243);
and U10040 (N_10040,N_9978,N_8493);
nor U10041 (N_10041,N_5184,N_5864);
and U10042 (N_10042,N_5105,N_5221);
nand U10043 (N_10043,N_5944,N_5424);
xor U10044 (N_10044,N_7669,N_5509);
nor U10045 (N_10045,N_6739,N_6756);
or U10046 (N_10046,N_8779,N_9670);
nand U10047 (N_10047,N_6536,N_6065);
nor U10048 (N_10048,N_5372,N_7200);
or U10049 (N_10049,N_5506,N_9153);
and U10050 (N_10050,N_9606,N_6659);
nand U10051 (N_10051,N_9530,N_7182);
or U10052 (N_10052,N_6164,N_7632);
nor U10053 (N_10053,N_6124,N_7380);
nor U10054 (N_10054,N_6591,N_8071);
nor U10055 (N_10055,N_7617,N_8323);
or U10056 (N_10056,N_9090,N_7496);
nor U10057 (N_10057,N_7545,N_8838);
and U10058 (N_10058,N_6220,N_5725);
or U10059 (N_10059,N_7502,N_7644);
nor U10060 (N_10060,N_6918,N_8525);
nor U10061 (N_10061,N_8811,N_6460);
nand U10062 (N_10062,N_5350,N_7124);
xnor U10063 (N_10063,N_5501,N_9507);
nand U10064 (N_10064,N_5730,N_6951);
and U10065 (N_10065,N_5879,N_8154);
nor U10066 (N_10066,N_8265,N_7587);
or U10067 (N_10067,N_8644,N_5718);
nor U10068 (N_10068,N_6806,N_7571);
nor U10069 (N_10069,N_9046,N_8760);
or U10070 (N_10070,N_8799,N_6170);
or U10071 (N_10071,N_7719,N_9183);
nand U10072 (N_10072,N_7133,N_5125);
or U10073 (N_10073,N_5592,N_9991);
and U10074 (N_10074,N_9027,N_6556);
or U10075 (N_10075,N_5845,N_6141);
nand U10076 (N_10076,N_9119,N_9207);
or U10077 (N_10077,N_9000,N_7607);
or U10078 (N_10078,N_7347,N_6288);
nor U10079 (N_10079,N_6775,N_6781);
or U10080 (N_10080,N_6575,N_6505);
nand U10081 (N_10081,N_9062,N_7148);
nand U10082 (N_10082,N_8787,N_5305);
or U10083 (N_10083,N_5134,N_7432);
and U10084 (N_10084,N_8035,N_7900);
and U10085 (N_10085,N_8516,N_7964);
nand U10086 (N_10086,N_7915,N_7491);
or U10087 (N_10087,N_8828,N_9615);
nor U10088 (N_10088,N_5167,N_7848);
or U10089 (N_10089,N_8094,N_8600);
nor U10090 (N_10090,N_9217,N_8701);
nand U10091 (N_10091,N_6673,N_7076);
and U10092 (N_10092,N_9731,N_9011);
nor U10093 (N_10093,N_6593,N_8906);
nor U10094 (N_10094,N_8778,N_8583);
nand U10095 (N_10095,N_6510,N_7335);
nor U10096 (N_10096,N_9882,N_8240);
nor U10097 (N_10097,N_8266,N_9225);
xor U10098 (N_10098,N_5407,N_5449);
nand U10099 (N_10099,N_5175,N_5201);
and U10100 (N_10100,N_5417,N_5445);
or U10101 (N_10101,N_7880,N_5243);
and U10102 (N_10102,N_7501,N_7938);
nand U10103 (N_10103,N_7961,N_9117);
nand U10104 (N_10104,N_5789,N_6725);
and U10105 (N_10105,N_5135,N_7864);
or U10106 (N_10106,N_9084,N_9920);
and U10107 (N_10107,N_8844,N_7277);
nand U10108 (N_10108,N_6327,N_9852);
and U10109 (N_10109,N_5024,N_6737);
nor U10110 (N_10110,N_6043,N_6297);
nand U10111 (N_10111,N_5629,N_8260);
or U10112 (N_10112,N_6216,N_7140);
and U10113 (N_10113,N_6315,N_5164);
or U10114 (N_10114,N_7305,N_7459);
and U10115 (N_10115,N_7542,N_7497);
nor U10116 (N_10116,N_6910,N_5825);
and U10117 (N_10117,N_7025,N_8820);
nand U10118 (N_10118,N_7803,N_5042);
nor U10119 (N_10119,N_5670,N_5652);
or U10120 (N_10120,N_8785,N_6430);
nor U10121 (N_10121,N_7831,N_7532);
nand U10122 (N_10122,N_9927,N_7167);
nand U10123 (N_10123,N_5368,N_8716);
nor U10124 (N_10124,N_9483,N_7372);
and U10125 (N_10125,N_9146,N_9222);
nand U10126 (N_10126,N_6862,N_8872);
nor U10127 (N_10127,N_9083,N_5640);
nor U10128 (N_10128,N_8226,N_7169);
nor U10129 (N_10129,N_6222,N_7663);
and U10130 (N_10130,N_5067,N_8440);
nand U10131 (N_10131,N_6018,N_6416);
nor U10132 (N_10132,N_7135,N_9470);
and U10133 (N_10133,N_5514,N_8141);
nand U10134 (N_10134,N_7780,N_9880);
and U10135 (N_10135,N_8394,N_9548);
or U10136 (N_10136,N_7260,N_9742);
and U10137 (N_10137,N_9209,N_9924);
or U10138 (N_10138,N_6610,N_6056);
or U10139 (N_10139,N_9894,N_9841);
nor U10140 (N_10140,N_9294,N_9045);
and U10141 (N_10141,N_8291,N_5028);
nand U10142 (N_10142,N_8434,N_7294);
nand U10143 (N_10143,N_8252,N_9120);
or U10144 (N_10144,N_8224,N_8300);
and U10145 (N_10145,N_8788,N_5385);
and U10146 (N_10146,N_7885,N_9901);
nor U10147 (N_10147,N_5542,N_5456);
or U10148 (N_10148,N_9667,N_7709);
and U10149 (N_10149,N_8978,N_5881);
nand U10150 (N_10150,N_5531,N_5307);
and U10151 (N_10151,N_5357,N_7868);
and U10152 (N_10152,N_5814,N_7410);
nand U10153 (N_10153,N_6326,N_9908);
nand U10154 (N_10154,N_5851,N_8248);
or U10155 (N_10155,N_8682,N_5714);
or U10156 (N_10156,N_5204,N_6837);
nand U10157 (N_10157,N_8253,N_9680);
xnor U10158 (N_10158,N_6695,N_5062);
xor U10159 (N_10159,N_6271,N_8160);
and U10160 (N_10160,N_9356,N_7495);
nor U10161 (N_10161,N_9234,N_8993);
or U10162 (N_10162,N_7082,N_8810);
nor U10163 (N_10163,N_8042,N_6176);
or U10164 (N_10164,N_9337,N_8798);
nand U10165 (N_10165,N_8743,N_6606);
or U10166 (N_10166,N_9434,N_6313);
or U10167 (N_10167,N_9768,N_9258);
nand U10168 (N_10168,N_7996,N_9017);
nand U10169 (N_10169,N_7834,N_5268);
or U10170 (N_10170,N_5587,N_5381);
and U10171 (N_10171,N_9568,N_6988);
xor U10172 (N_10172,N_9203,N_6014);
or U10173 (N_10173,N_7143,N_7474);
or U10174 (N_10174,N_7877,N_5802);
nor U10175 (N_10175,N_7762,N_9231);
and U10176 (N_10176,N_7117,N_5055);
and U10177 (N_10177,N_8262,N_6708);
nor U10178 (N_10178,N_5994,N_9812);
nand U10179 (N_10179,N_6492,N_7947);
and U10180 (N_10180,N_9412,N_6645);
and U10181 (N_10181,N_8986,N_8378);
nand U10182 (N_10182,N_8825,N_7763);
xnor U10183 (N_10183,N_9306,N_9279);
and U10184 (N_10184,N_9896,N_7521);
nand U10185 (N_10185,N_6560,N_8665);
nand U10186 (N_10186,N_7091,N_8786);
and U10187 (N_10187,N_7552,N_5760);
or U10188 (N_10188,N_5533,N_7952);
nor U10189 (N_10189,N_6516,N_8009);
and U10190 (N_10190,N_5959,N_8954);
nor U10191 (N_10191,N_9613,N_9747);
and U10192 (N_10192,N_6394,N_9029);
or U10193 (N_10193,N_8696,N_5137);
nand U10194 (N_10194,N_9953,N_9527);
nand U10195 (N_10195,N_9298,N_9939);
nor U10196 (N_10196,N_6880,N_8025);
and U10197 (N_10197,N_8081,N_9148);
or U10198 (N_10198,N_7873,N_6827);
xor U10199 (N_10199,N_6330,N_8168);
or U10200 (N_10200,N_7767,N_8128);
nor U10201 (N_10201,N_6960,N_9113);
or U10202 (N_10202,N_7022,N_8623);
and U10203 (N_10203,N_9506,N_9807);
nor U10204 (N_10204,N_7478,N_8853);
nand U10205 (N_10205,N_6522,N_6142);
and U10206 (N_10206,N_9601,N_5643);
nand U10207 (N_10207,N_6668,N_8393);
xnor U10208 (N_10208,N_9278,N_5997);
and U10209 (N_10209,N_5658,N_9289);
and U10210 (N_10210,N_6929,N_7995);
nor U10211 (N_10211,N_8187,N_9677);
nand U10212 (N_10212,N_7578,N_5130);
nor U10213 (N_10213,N_9473,N_9674);
nor U10214 (N_10214,N_7470,N_7218);
or U10215 (N_10215,N_8340,N_9824);
or U10216 (N_10216,N_6228,N_9849);
and U10217 (N_10217,N_9031,N_6799);
or U10218 (N_10218,N_9210,N_5702);
and U10219 (N_10219,N_9701,N_7725);
nor U10220 (N_10220,N_8792,N_5401);
and U10221 (N_10221,N_8246,N_8919);
nor U10222 (N_10222,N_6692,N_6419);
nand U10223 (N_10223,N_6199,N_7860);
nor U10224 (N_10224,N_6848,N_5279);
nor U10225 (N_10225,N_9697,N_5064);
nor U10226 (N_10226,N_6789,N_5242);
or U10227 (N_10227,N_5092,N_6221);
and U10228 (N_10228,N_5724,N_7040);
and U10229 (N_10229,N_8230,N_5508);
or U10230 (N_10230,N_5388,N_6295);
or U10231 (N_10231,N_6426,N_7906);
xor U10232 (N_10232,N_6537,N_9163);
nand U10233 (N_10233,N_7703,N_8011);
and U10234 (N_10234,N_8733,N_8088);
nor U10235 (N_10235,N_5053,N_9886);
and U10236 (N_10236,N_8851,N_5202);
nand U10237 (N_10237,N_5143,N_7603);
xor U10238 (N_10238,N_5193,N_7358);
nand U10239 (N_10239,N_6549,N_8180);
or U10240 (N_10240,N_6783,N_5673);
or U10241 (N_10241,N_8878,N_6025);
nor U10242 (N_10242,N_5521,N_7816);
and U10243 (N_10243,N_9887,N_8683);
nand U10244 (N_10244,N_8585,N_7329);
and U10245 (N_10245,N_7458,N_9583);
or U10246 (N_10246,N_8713,N_5320);
nand U10247 (N_10247,N_5219,N_9254);
and U10248 (N_10248,N_6404,N_9546);
and U10249 (N_10249,N_6248,N_5768);
or U10250 (N_10250,N_5122,N_9273);
and U10251 (N_10251,N_7454,N_5044);
nand U10252 (N_10252,N_8790,N_5603);
or U10253 (N_10253,N_6178,N_6380);
nand U10254 (N_10254,N_7484,N_9429);
and U10255 (N_10255,N_7321,N_9302);
and U10256 (N_10256,N_5133,N_6672);
or U10257 (N_10257,N_9539,N_9270);
nor U10258 (N_10258,N_6085,N_8761);
nand U10259 (N_10259,N_9476,N_5084);
and U10260 (N_10260,N_9989,N_8604);
nor U10261 (N_10261,N_9964,N_7685);
and U10262 (N_10262,N_5174,N_9373);
or U10263 (N_10263,N_7047,N_9474);
nor U10264 (N_10264,N_8946,N_9475);
or U10265 (N_10265,N_7238,N_8972);
nor U10266 (N_10266,N_9538,N_5970);
nor U10267 (N_10267,N_5834,N_7159);
nand U10268 (N_10268,N_7773,N_9172);
or U10269 (N_10269,N_5181,N_7345);
and U10270 (N_10270,N_6697,N_9004);
or U10271 (N_10271,N_6869,N_8655);
nand U10272 (N_10272,N_6156,N_7258);
nor U10273 (N_10273,N_6874,N_5274);
or U10274 (N_10274,N_8095,N_6499);
and U10275 (N_10275,N_7754,N_7798);
or U10276 (N_10276,N_6282,N_6107);
or U10277 (N_10277,N_5941,N_7727);
nand U10278 (N_10278,N_8568,N_9664);
and U10279 (N_10279,N_8537,N_6603);
nor U10280 (N_10280,N_8868,N_9353);
and U10281 (N_10281,N_6508,N_7581);
nand U10282 (N_10282,N_9968,N_6845);
or U10283 (N_10283,N_5615,N_5910);
or U10284 (N_10284,N_9411,N_8331);
nor U10285 (N_10285,N_6831,N_9969);
nand U10286 (N_10286,N_8554,N_7211);
nand U10287 (N_10287,N_9537,N_9907);
nand U10288 (N_10288,N_7292,N_6979);
or U10289 (N_10289,N_7978,N_7979);
nand U10290 (N_10290,N_9040,N_8529);
or U10291 (N_10291,N_9039,N_9695);
or U10292 (N_10292,N_7660,N_7067);
xor U10293 (N_10293,N_7867,N_8392);
nor U10294 (N_10294,N_5329,N_5148);
nand U10295 (N_10295,N_5917,N_8111);
nand U10296 (N_10296,N_6227,N_9779);
and U10297 (N_10297,N_5698,N_6238);
nand U10298 (N_10298,N_6009,N_8812);
and U10299 (N_10299,N_5735,N_6320);
nor U10300 (N_10300,N_6515,N_9202);
nand U10301 (N_10301,N_6876,N_8857);
or U10302 (N_10302,N_6046,N_7287);
nor U10303 (N_10303,N_7696,N_7422);
nand U10304 (N_10304,N_5573,N_8358);
nor U10305 (N_10305,N_7077,N_7477);
or U10306 (N_10306,N_9092,N_8515);
and U10307 (N_10307,N_9136,N_8254);
or U10308 (N_10308,N_6663,N_8902);
nor U10309 (N_10309,N_9446,N_8867);
nor U10310 (N_10310,N_5228,N_8957);
or U10311 (N_10311,N_9357,N_8460);
nor U10312 (N_10312,N_7138,N_8741);
or U10313 (N_10313,N_7369,N_6595);
and U10314 (N_10314,N_8387,N_8669);
nand U10315 (N_10315,N_7317,N_8158);
or U10316 (N_10316,N_7086,N_8150);
and U10317 (N_10317,N_7766,N_8191);
nor U10318 (N_10318,N_8730,N_8890);
nand U10319 (N_10319,N_6276,N_9574);
and U10320 (N_10320,N_7393,N_7215);
nand U10321 (N_10321,N_7375,N_9350);
and U10322 (N_10322,N_7958,N_6078);
or U10323 (N_10323,N_7895,N_8702);
nand U10324 (N_10324,N_7433,N_8821);
or U10325 (N_10325,N_7569,N_5877);
nand U10326 (N_10326,N_5938,N_6209);
or U10327 (N_10327,N_6179,N_9728);
nand U10328 (N_10328,N_6965,N_5630);
nor U10329 (N_10329,N_7453,N_6932);
and U10330 (N_10330,N_7080,N_7673);
nor U10331 (N_10331,N_8606,N_9063);
and U10332 (N_10332,N_7267,N_5162);
and U10333 (N_10333,N_6760,N_5186);
or U10334 (N_10334,N_5505,N_9757);
or U10335 (N_10335,N_9095,N_5319);
or U10336 (N_10336,N_7889,N_7268);
nor U10337 (N_10337,N_6759,N_9525);
nor U10338 (N_10338,N_9056,N_8524);
or U10339 (N_10339,N_6250,N_5593);
or U10340 (N_10340,N_5237,N_5738);
or U10341 (N_10341,N_6474,N_7602);
nand U10342 (N_10342,N_6642,N_5614);
or U10343 (N_10343,N_8848,N_8735);
nand U10344 (N_10344,N_6011,N_5010);
nand U10345 (N_10345,N_7541,N_8155);
and U10346 (N_10346,N_5774,N_8936);
and U10347 (N_10347,N_5906,N_7739);
nand U10348 (N_10348,N_9866,N_7352);
or U10349 (N_10349,N_6149,N_9741);
and U10350 (N_10350,N_5019,N_6213);
and U10351 (N_10351,N_5389,N_7249);
and U10352 (N_10352,N_8391,N_7708);
and U10353 (N_10353,N_9992,N_9058);
and U10354 (N_10354,N_9957,N_6709);
nor U10355 (N_10355,N_8829,N_8127);
nor U10356 (N_10356,N_9874,N_8658);
nand U10357 (N_10357,N_5559,N_9218);
nand U10358 (N_10358,N_5599,N_7046);
nor U10359 (N_10359,N_6626,N_8998);
nand U10360 (N_10360,N_8797,N_5840);
or U10361 (N_10361,N_9245,N_9421);
nor U10362 (N_10362,N_5847,N_8461);
nor U10363 (N_10363,N_7801,N_5567);
nor U10364 (N_10364,N_5618,N_5142);
or U10365 (N_10365,N_8384,N_7024);
and U10366 (N_10366,N_6402,N_5912);
nand U10367 (N_10367,N_9732,N_6195);
and U10368 (N_10368,N_5656,N_9775);
nand U10369 (N_10369,N_7679,N_8306);
nor U10370 (N_10370,N_7450,N_7590);
and U10371 (N_10371,N_7993,N_6844);
and U10372 (N_10372,N_5518,N_5058);
nor U10373 (N_10373,N_8162,N_5620);
nand U10374 (N_10374,N_5411,N_5563);
xnor U10375 (N_10375,N_8079,N_8126);
nand U10376 (N_10376,N_9834,N_5611);
nor U10377 (N_10377,N_7424,N_6449);
or U10378 (N_10378,N_7311,N_5442);
nor U10379 (N_10379,N_6005,N_7483);
nor U10380 (N_10380,N_8603,N_7235);
and U10381 (N_10381,N_9154,N_7370);
nand U10382 (N_10382,N_5409,N_6289);
or U10383 (N_10383,N_9923,N_6552);
or U10384 (N_10384,N_8459,N_6722);
or U10385 (N_10385,N_9790,N_8030);
and U10386 (N_10386,N_9961,N_5172);
and U10387 (N_10387,N_9904,N_9929);
xnor U10388 (N_10388,N_5266,N_9888);
and U10389 (N_10389,N_7991,N_6007);
nand U10390 (N_10390,N_9648,N_6718);
nor U10391 (N_10391,N_8744,N_6808);
or U10392 (N_10392,N_5781,N_5267);
and U10393 (N_10393,N_5257,N_7851);
and U10394 (N_10394,N_5470,N_5886);
nand U10395 (N_10395,N_5537,N_5500);
and U10396 (N_10396,N_8439,N_6128);
nor U10397 (N_10397,N_9778,N_8144);
nand U10398 (N_10398,N_7536,N_6888);
or U10399 (N_10399,N_6071,N_8835);
or U10400 (N_10400,N_9481,N_9550);
nand U10401 (N_10401,N_5188,N_6809);
nand U10402 (N_10402,N_6738,N_5207);
nor U10403 (N_10403,N_7884,N_8342);
xnor U10404 (N_10404,N_6118,N_5855);
and U10405 (N_10405,N_6318,N_5867);
and U10406 (N_10406,N_8133,N_6643);
or U10407 (N_10407,N_9611,N_8947);
nor U10408 (N_10408,N_8272,N_7180);
nand U10409 (N_10409,N_6414,N_8146);
or U10410 (N_10410,N_5465,N_6959);
xor U10411 (N_10411,N_6632,N_5185);
nor U10412 (N_10412,N_7547,N_6480);
or U10413 (N_10413,N_5375,N_7427);
nand U10414 (N_10414,N_9660,N_7517);
xor U10415 (N_10415,N_6064,N_5649);
and U10416 (N_10416,N_9526,N_8667);
or U10417 (N_10417,N_6561,N_7652);
nor U10418 (N_10418,N_5655,N_8953);
nor U10419 (N_10419,N_9067,N_8448);
and U10420 (N_10420,N_7028,N_9575);
or U10421 (N_10421,N_7334,N_5050);
or U10422 (N_10422,N_5336,N_8468);
or U10423 (N_10423,N_8766,N_7426);
or U10424 (N_10424,N_7378,N_8015);
nand U10425 (N_10425,N_6052,N_9577);
nand U10426 (N_10426,N_6518,N_6524);
xor U10427 (N_10427,N_9573,N_7934);
and U10428 (N_10428,N_5119,N_5993);
nor U10429 (N_10429,N_5366,N_9232);
and U10430 (N_10430,N_5787,N_9689);
and U10431 (N_10431,N_6915,N_6165);
or U10432 (N_10432,N_8031,N_8940);
or U10433 (N_10433,N_9521,N_8620);
nand U10434 (N_10434,N_8420,N_7810);
nand U10435 (N_10435,N_7626,N_9342);
nor U10436 (N_10436,N_7481,N_6362);
and U10437 (N_10437,N_7339,N_6779);
nor U10438 (N_10438,N_9025,N_8474);
or U10439 (N_10439,N_9293,N_6667);
and U10440 (N_10440,N_8311,N_6028);
nand U10441 (N_10441,N_9903,N_5195);
nand U10442 (N_10442,N_7912,N_8653);
nand U10443 (N_10443,N_6386,N_5078);
nand U10444 (N_10444,N_8039,N_9338);
and U10445 (N_10445,N_8619,N_6554);
nand U10446 (N_10446,N_6323,N_9637);
nand U10447 (N_10447,N_6528,N_9739);
and U10448 (N_10448,N_9804,N_8463);
and U10449 (N_10449,N_5008,N_7073);
and U10450 (N_10450,N_9774,N_6937);
or U10451 (N_10451,N_7638,N_9043);
nand U10452 (N_10452,N_6923,N_8319);
nand U10453 (N_10453,N_8199,N_5346);
and U10454 (N_10454,N_7300,N_5933);
or U10455 (N_10455,N_6433,N_8136);
and U10456 (N_10456,N_9023,N_8822);
and U10457 (N_10457,N_6173,N_5680);
or U10458 (N_10458,N_8710,N_5613);
and U10459 (N_10459,N_9361,N_6080);
xor U10460 (N_10460,N_8281,N_6100);
nand U10461 (N_10461,N_5081,N_6675);
or U10462 (N_10462,N_6770,N_7109);
and U10463 (N_10463,N_6558,N_6720);
and U10464 (N_10464,N_8666,N_6598);
and U10465 (N_10465,N_5973,N_5792);
nor U10466 (N_10466,N_5747,N_8973);
nor U10467 (N_10467,N_8115,N_8377);
nor U10468 (N_10468,N_5491,N_9515);
and U10469 (N_10469,N_9347,N_9443);
or U10470 (N_10470,N_7353,N_9427);
nor U10471 (N_10471,N_9239,N_5636);
or U10472 (N_10472,N_7172,N_6828);
or U10473 (N_10473,N_7302,N_7676);
and U10474 (N_10474,N_6013,N_5244);
nand U10475 (N_10475,N_5525,N_7017);
and U10476 (N_10476,N_6802,N_5069);
nor U10477 (N_10477,N_6553,N_6378);
or U10478 (N_10478,N_6385,N_9524);
or U10479 (N_10479,N_9578,N_7994);
or U10480 (N_10480,N_8558,N_9944);
and U10481 (N_10481,N_6217,N_8408);
or U10482 (N_10482,N_7844,N_6990);
nor U10483 (N_10483,N_9703,N_7093);
nand U10484 (N_10484,N_6249,N_8024);
nand U10485 (N_10485,N_8037,N_7373);
and U10486 (N_10486,N_9788,N_7823);
and U10487 (N_10487,N_7534,N_7515);
or U10488 (N_10488,N_5926,N_7746);
nor U10489 (N_10489,N_7634,N_8477);
and U10490 (N_10490,N_7349,N_8630);
nor U10491 (N_10491,N_7630,N_7207);
nand U10492 (N_10492,N_6422,N_6944);
nand U10493 (N_10493,N_7695,N_5331);
or U10494 (N_10494,N_7883,N_5771);
or U10495 (N_10495,N_5685,N_7014);
nor U10496 (N_10496,N_8104,N_5080);
nand U10497 (N_10497,N_9545,N_8225);
and U10498 (N_10498,N_9382,N_5918);
and U10499 (N_10499,N_7544,N_6963);
and U10500 (N_10500,N_7058,N_6572);
nor U10501 (N_10501,N_6345,N_9709);
or U10502 (N_10502,N_5475,N_8131);
nand U10503 (N_10503,N_9301,N_5335);
nand U10504 (N_10504,N_7817,N_7113);
nor U10505 (N_10505,N_7461,N_7406);
xor U10506 (N_10506,N_8292,N_5566);
or U10507 (N_10507,N_8123,N_8027);
nand U10508 (N_10508,N_8654,N_5369);
nand U10509 (N_10509,N_6300,N_6146);
xnor U10510 (N_10510,N_9921,N_9590);
nand U10511 (N_10511,N_6233,N_8269);
and U10512 (N_10512,N_8330,N_7941);
nor U10513 (N_10513,N_8103,N_6872);
and U10514 (N_10514,N_6342,N_9922);
or U10515 (N_10515,N_6203,N_8969);
nor U10516 (N_10516,N_7494,N_5005);
or U10517 (N_10517,N_6657,N_5015);
xnor U10518 (N_10518,N_5355,N_6198);
nor U10519 (N_10519,N_8925,N_5996);
nor U10520 (N_10520,N_9815,N_7063);
and U10521 (N_10521,N_9171,N_8019);
and U10522 (N_10522,N_5303,N_9074);
and U10523 (N_10523,N_6223,N_7723);
and U10524 (N_10524,N_5211,N_9628);
nand U10525 (N_10525,N_6636,N_9817);
nor U10526 (N_10526,N_7184,N_6177);
nor U10527 (N_10527,N_9686,N_7956);
nand U10528 (N_10528,N_5441,N_9818);
or U10529 (N_10529,N_9426,N_9793);
and U10530 (N_10530,N_9299,N_9325);
nand U10531 (N_10531,N_6791,N_5651);
nand U10532 (N_10532,N_9178,N_8373);
or U10533 (N_10533,N_9752,N_5088);
and U10534 (N_10534,N_9432,N_5887);
and U10535 (N_10535,N_9111,N_6439);
nand U10536 (N_10536,N_9167,N_9895);
nor U10537 (N_10537,N_9592,N_7130);
nand U10538 (N_10538,N_7691,N_8561);
nor U10539 (N_10539,N_5889,N_6035);
nand U10540 (N_10540,N_9876,N_5568);
and U10541 (N_10541,N_5756,N_8227);
nor U10542 (N_10542,N_8368,N_6048);
or U10543 (N_10543,N_9118,N_7508);
and U10544 (N_10544,N_5301,N_6940);
nand U10545 (N_10545,N_5440,N_9200);
and U10546 (N_10546,N_7570,N_8694);
or U10547 (N_10547,N_5095,N_5607);
and U10548 (N_10548,N_8411,N_5545);
and U10549 (N_10549,N_7683,N_5283);
nor U10550 (N_10550,N_8322,N_6771);
nor U10551 (N_10551,N_9838,N_6162);
nand U10552 (N_10552,N_5102,N_8204);
and U10553 (N_10553,N_9206,N_8495);
xnor U10554 (N_10554,N_9806,N_8189);
nand U10555 (N_10555,N_5594,N_6985);
and U10556 (N_10556,N_7472,N_8072);
xnor U10557 (N_10557,N_7151,N_6621);
nand U10558 (N_10558,N_9771,N_7601);
nor U10559 (N_10559,N_5576,N_6049);
and U10560 (N_10560,N_8503,N_9900);
or U10561 (N_10561,N_9684,N_7713);
nand U10562 (N_10562,N_5057,N_9496);
nand U10563 (N_10563,N_6088,N_5793);
and U10564 (N_10564,N_9566,N_7548);
and U10565 (N_10565,N_5965,N_9341);
nor U10566 (N_10566,N_6109,N_8006);
and U10567 (N_10567,N_5830,N_6185);
nor U10568 (N_10568,N_7301,N_9123);
nand U10569 (N_10569,N_6817,N_7419);
nor U10570 (N_10570,N_5018,N_9861);
nand U10571 (N_10571,N_9714,N_5298);
nand U10572 (N_10572,N_7185,N_9365);
nand U10573 (N_10573,N_8379,N_5530);
nor U10574 (N_10574,N_6302,N_6479);
xor U10575 (N_10575,N_8794,N_8628);
nand U10576 (N_10576,N_7778,N_6527);
and U10577 (N_10577,N_9144,N_8490);
xor U10578 (N_10578,N_6542,N_7059);
and U10579 (N_10579,N_6401,N_8264);
nor U10580 (N_10580,N_7838,N_9141);
nor U10581 (N_10581,N_5100,N_5173);
and U10582 (N_10582,N_9199,N_5216);
nand U10583 (N_10583,N_6333,N_6658);
nand U10584 (N_10584,N_6682,N_8886);
nor U10585 (N_10585,N_7635,N_7872);
nand U10586 (N_10586,N_8971,N_6856);
xor U10587 (N_10587,N_8413,N_8426);
or U10588 (N_10588,N_5302,N_5126);
nand U10589 (N_10589,N_9950,N_9013);
xnor U10590 (N_10590,N_5308,N_6649);
or U10591 (N_10591,N_8289,N_6472);
nand U10592 (N_10592,N_8370,N_8674);
or U10593 (N_10593,N_7954,N_8780);
and U10594 (N_10594,N_7257,N_5273);
or U10595 (N_10595,N_6105,N_6531);
nand U10596 (N_10596,N_6390,N_9564);
or U10597 (N_10597,N_5418,N_5001);
and U10598 (N_10598,N_6382,N_7136);
and U10599 (N_10599,N_7214,N_5891);
and U10600 (N_10600,N_5954,N_9976);
nor U10601 (N_10601,N_9938,N_8372);
nand U10602 (N_10602,N_7753,N_8482);
or U10603 (N_10603,N_6911,N_9066);
or U10604 (N_10604,N_9612,N_8805);
and U10605 (N_10605,N_9324,N_8206);
nand U10606 (N_10606,N_7835,N_9458);
nor U10607 (N_10607,N_9942,N_9467);
or U10608 (N_10608,N_5098,N_7814);
and U10609 (N_10609,N_5271,N_5663);
nand U10610 (N_10610,N_5515,N_6359);
nand U10611 (N_10611,N_6724,N_7156);
nand U10612 (N_10612,N_7749,N_6360);
and U10613 (N_10613,N_7960,N_5161);
nor U10614 (N_10614,N_7068,N_8018);
and U10615 (N_10615,N_7748,N_6106);
xnor U10616 (N_10616,N_8065,N_5803);
nor U10617 (N_10617,N_8649,N_6920);
or U10618 (N_10618,N_5554,N_9050);
nor U10619 (N_10619,N_9719,N_6752);
or U10620 (N_10620,N_7771,N_8684);
nor U10621 (N_10621,N_6010,N_5985);
nor U10622 (N_10622,N_6646,N_6324);
nand U10623 (N_10623,N_8726,N_8773);
or U10624 (N_10624,N_5478,N_9563);
nor U10625 (N_10625,N_9451,N_7882);
nor U10626 (N_10626,N_5532,N_7743);
and U10627 (N_10627,N_9661,N_8803);
xor U10628 (N_10628,N_9645,N_7111);
nand U10629 (N_10629,N_9425,N_6652);
or U10630 (N_10630,N_5408,N_9396);
nand U10631 (N_10631,N_8592,N_6769);
and U10632 (N_10632,N_7057,N_7079);
nor U10633 (N_10633,N_6081,N_8924);
nor U10634 (N_10634,N_6171,N_7628);
nand U10635 (N_10635,N_8897,N_9974);
nand U10636 (N_10636,N_9070,N_8406);
nor U10637 (N_10637,N_8318,N_8301);
nand U10638 (N_10638,N_7383,N_5448);
nor U10639 (N_10639,N_6096,N_7197);
and U10640 (N_10640,N_9819,N_5106);
nand U10641 (N_10641,N_6943,N_8855);
or U10642 (N_10642,N_8479,N_5068);
nand U10643 (N_10643,N_7562,N_5197);
and U10644 (N_10644,N_8888,N_5248);
or U10645 (N_10645,N_8933,N_7208);
nand U10646 (N_10646,N_6135,N_8497);
nand U10647 (N_10647,N_9945,N_9280);
nor U10648 (N_10648,N_7283,N_6008);
or U10649 (N_10649,N_5874,N_5490);
or U10650 (N_10650,N_8257,N_9175);
nor U10651 (N_10651,N_5731,N_8419);
nor U10652 (N_10652,N_5928,N_5497);
or U10653 (N_10653,N_8675,N_6437);
nor U10654 (N_10654,N_8488,N_9952);
nor U10655 (N_10655,N_7127,N_8807);
and U10656 (N_10656,N_9264,N_9155);
and U10657 (N_10657,N_9917,N_8673);
or U10658 (N_10658,N_5484,N_6777);
nand U10659 (N_10659,N_6202,N_5118);
and U10660 (N_10660,N_5966,N_7852);
nor U10661 (N_10661,N_6666,N_5245);
or U10662 (N_10662,N_7648,N_5317);
or U10663 (N_10663,N_7285,N_6373);
nor U10664 (N_10664,N_6906,N_8091);
nor U10665 (N_10665,N_9101,N_5662);
nor U10666 (N_10666,N_5940,N_6857);
nand U10667 (N_10667,N_6154,N_6053);
or U10668 (N_10668,N_5565,N_5386);
or U10669 (N_10669,N_7161,N_6967);
nor U10670 (N_10670,N_7384,N_6982);
and U10671 (N_10671,N_8708,N_5734);
nand U10672 (N_10672,N_7064,N_7613);
nand U10673 (N_10673,N_6519,N_5550);
or U10674 (N_10674,N_7913,N_7449);
nand U10675 (N_10675,N_5226,N_5347);
and U10676 (N_10676,N_7103,N_6671);
nor U10677 (N_10677,N_8992,N_8995);
nand U10678 (N_10678,N_8532,N_7671);
and U10679 (N_10679,N_8632,N_8703);
nor U10680 (N_10680,N_5805,N_5895);
nand U10681 (N_10681,N_8586,N_6066);
and U10682 (N_10682,N_6506,N_9556);
nor U10683 (N_10683,N_5280,N_5727);
nand U10684 (N_10684,N_7916,N_9138);
and U10685 (N_10685,N_5677,N_8637);
nor U10686 (N_10686,N_5513,N_8442);
nor U10687 (N_10687,N_5000,N_9266);
nor U10688 (N_10688,N_5956,N_9794);
and U10689 (N_10689,N_5524,N_7651);
or U10690 (N_10690,N_6786,N_5536);
nand U10691 (N_10691,N_7413,N_6866);
nor U10692 (N_10692,N_5110,N_6033);
or U10693 (N_10693,N_5998,N_5314);
or U10694 (N_10694,N_5949,N_5498);
and U10695 (N_10695,N_9305,N_8704);
or U10696 (N_10696,N_5645,N_6099);
nor U10697 (N_10697,N_6533,N_8443);
nor U10698 (N_10698,N_8549,N_8309);
nand U10699 (N_10699,N_8861,N_7036);
and U10700 (N_10700,N_7239,N_6917);
nand U10701 (N_10701,N_5541,N_8903);
or U10702 (N_10702,N_7750,N_6121);
nor U10703 (N_10703,N_7710,N_9509);
nor U10704 (N_10704,N_7187,N_6237);
nand U10705 (N_10705,N_5399,N_9786);
nand U10706 (N_10706,N_5968,N_6520);
nand U10707 (N_10707,N_8983,N_6966);
nand U10708 (N_10708,N_5121,N_8698);
or U10709 (N_10709,N_5619,N_7273);
nand U10710 (N_10710,N_8038,N_9351);
nand U10711 (N_10711,N_8371,N_6614);
nand U10712 (N_10712,N_8588,N_5412);
nand U10713 (N_10713,N_8560,N_7667);
and U10714 (N_10714,N_9792,N_8002);
or U10715 (N_10715,N_5077,N_9098);
and U10716 (N_10716,N_6891,N_9189);
nor U10717 (N_10717,N_9898,N_7861);
nand U10718 (N_10718,N_8353,N_5166);
or U10719 (N_10719,N_9216,N_8101);
or U10720 (N_10720,N_7356,N_7071);
xnor U10721 (N_10721,N_5047,N_9899);
nand U10722 (N_10722,N_6859,N_9871);
nand U10723 (N_10723,N_5581,N_9364);
and U10724 (N_10724,N_9692,N_9623);
nor U10725 (N_10725,N_5964,N_7764);
and U10726 (N_10726,N_5231,N_9149);
and U10727 (N_10727,N_7395,N_5073);
or U10728 (N_10728,N_6137,N_8022);
and U10729 (N_10729,N_9261,N_8066);
nand U10730 (N_10730,N_7940,N_6215);
nor U10731 (N_10731,N_7409,N_7654);
nand U10732 (N_10732,N_8976,N_7811);
and U10733 (N_10733,N_7085,N_6332);
or U10734 (N_10734,N_5743,N_5623);
or U10735 (N_10735,N_6564,N_6517);
nand U10736 (N_10736,N_6578,N_9493);
and U10737 (N_10737,N_9561,N_8845);
nor U10738 (N_10738,N_6307,N_8677);
or U10739 (N_10739,N_5626,N_9681);
nand U10740 (N_10740,N_5608,N_5076);
and U10741 (N_10741,N_5721,N_7969);
xor U10742 (N_10742,N_9269,N_9014);
or U10743 (N_10743,N_5494,N_7318);
nand U10744 (N_10744,N_8913,N_8955);
and U10745 (N_10745,N_8396,N_8166);
or U10746 (N_10746,N_5153,N_5155);
or U10747 (N_10747,N_9333,N_7048);
and U10748 (N_10748,N_6408,N_6157);
and U10749 (N_10749,N_8207,N_8048);
nor U10750 (N_10750,N_7251,N_9041);
nand U10751 (N_10751,N_9442,N_8157);
or U10752 (N_10752,N_7417,N_5711);
nor U10753 (N_10753,N_8706,N_5312);
nand U10754 (N_10754,N_8436,N_6229);
nor U10755 (N_10755,N_7271,N_6545);
or U10756 (N_10756,N_9230,N_7275);
nor U10757 (N_10757,N_9419,N_9941);
nor U10758 (N_10758,N_9007,N_9139);
and U10759 (N_10759,N_6393,N_8132);
or U10760 (N_10760,N_7876,N_5165);
nor U10761 (N_10761,N_5713,N_7145);
nor U10762 (N_10762,N_5706,N_5029);
and U10763 (N_10763,N_8333,N_7003);
and U10764 (N_10764,N_7286,N_6267);
nand U10765 (N_10765,N_9089,N_8912);
nor U10766 (N_10766,N_5060,N_7647);
and U10767 (N_10767,N_6079,N_9237);
and U10768 (N_10768,N_9916,N_7737);
nor U10769 (N_10769,N_9502,N_5665);
or U10770 (N_10770,N_9832,N_5701);
and U10771 (N_10771,N_6245,N_5975);
or U10772 (N_10772,N_6892,N_7052);
nor U10773 (N_10773,N_6115,N_9450);
nand U10774 (N_10774,N_8341,N_8952);
xnor U10775 (N_10775,N_5590,N_9885);
nand U10776 (N_10776,N_7514,N_5653);
or U10777 (N_10777,N_8757,N_7711);
and U10778 (N_10778,N_5913,N_6551);
nor U10779 (N_10779,N_7712,N_8917);
nor U10780 (N_10780,N_7414,N_9477);
nor U10781 (N_10781,N_6306,N_8179);
nor U10782 (N_10782,N_6730,N_8582);
or U10783 (N_10783,N_7016,N_8445);
and U10784 (N_10784,N_5218,N_6395);
nor U10785 (N_10785,N_5880,N_8945);
nor U10786 (N_10786,N_8748,N_5376);
nor U10787 (N_10787,N_5775,N_6734);
and U10788 (N_10788,N_9049,N_6810);
nand U10789 (N_10789,N_9401,N_5728);
nor U10790 (N_10790,N_7102,N_6694);
nor U10791 (N_10791,N_6933,N_8458);
or U10792 (N_10792,N_8599,N_8563);
and U10793 (N_10793,N_5429,N_7879);
xnor U10794 (N_10794,N_8846,N_8602);
and U10795 (N_10795,N_9706,N_7756);
nor U10796 (N_10796,N_6681,N_5430);
and U10797 (N_10797,N_5227,N_6021);
and U10798 (N_10798,N_9156,N_7376);
or U10799 (N_10799,N_8324,N_5754);
or U10800 (N_10800,N_5987,N_8535);
or U10801 (N_10801,N_8749,N_6885);
and U10802 (N_10802,N_5394,N_5006);
and U10803 (N_10803,N_5779,N_6798);
or U10804 (N_10804,N_9857,N_5304);
nand U10805 (N_10805,N_5642,N_9311);
or U10806 (N_10806,N_8086,N_8056);
and U10807 (N_10807,N_9388,N_6811);
nand U10808 (N_10808,N_6889,N_9914);
nand U10809 (N_10809,N_5093,N_9847);
nor U10810 (N_10810,N_9122,N_6192);
nand U10811 (N_10811,N_5083,N_9789);
or U10812 (N_10812,N_9808,N_8464);
nor U10813 (N_10813,N_6927,N_7284);
nor U10814 (N_10814,N_7962,N_7357);
and U10815 (N_10815,N_5794,N_6314);
and U10816 (N_10816,N_5061,N_5025);
or U10817 (N_10817,N_7758,N_6772);
nor U10818 (N_10818,N_5539,N_8329);
nor U10819 (N_10819,N_6867,N_6921);
or U10820 (N_10820,N_5354,N_6523);
and U10821 (N_10821,N_8429,N_8720);
or U10822 (N_10822,N_8007,N_9855);
nand U10823 (N_10823,N_9186,N_7808);
and U10824 (N_10824,N_6148,N_8310);
nor U10825 (N_10825,N_9195,N_6980);
nor U10826 (N_10826,N_8591,N_5250);
and U10827 (N_10827,N_5258,N_6341);
nor U10828 (N_10828,N_7825,N_8645);
and U10829 (N_10829,N_5671,N_8467);
and U10830 (N_10830,N_8562,N_8944);
and U10831 (N_10831,N_5923,N_7027);
or U10832 (N_10832,N_5544,N_8093);
nand U10833 (N_10833,N_6134,N_6044);
nand U10834 (N_10834,N_6942,N_6839);
xnor U10835 (N_10835,N_5502,N_6648);
nand U10836 (N_10836,N_7599,N_6555);
nand U10837 (N_10837,N_6299,N_8188);
nor U10838 (N_10838,N_8352,N_6319);
nor U10839 (N_10839,N_9559,N_7785);
xor U10840 (N_10840,N_8217,N_8125);
nand U10841 (N_10841,N_8738,N_5485);
nor U10842 (N_10842,N_7568,N_6374);
or U10843 (N_10843,N_7039,N_8354);
or U10844 (N_10844,N_5962,N_6358);
and U10845 (N_10845,N_7035,N_6543);
nor U10846 (N_10846,N_6204,N_8580);
and U10847 (N_10847,N_8700,N_6761);
or U10848 (N_10848,N_7760,N_9549);
and U10849 (N_10849,N_8553,N_6015);
nand U10850 (N_10850,N_7788,N_7875);
or U10851 (N_10851,N_9936,N_8609);
or U10852 (N_10852,N_5548,N_9374);
nand U10853 (N_10853,N_7557,N_8435);
nand U10854 (N_10854,N_6583,N_5538);
nand U10855 (N_10855,N_6997,N_7686);
nand U10856 (N_10856,N_8893,N_5991);
nand U10857 (N_10857,N_9919,N_8680);
or U10858 (N_10858,N_6883,N_5829);
and U10859 (N_10859,N_9219,N_7465);
and U10860 (N_10860,N_9313,N_9813);
and U10861 (N_10861,N_5832,N_9406);
nor U10862 (N_10862,N_8386,N_5764);
and U10863 (N_10863,N_5294,N_5748);
nor U10864 (N_10864,N_6047,N_5841);
xnor U10865 (N_10865,N_6887,N_7745);
nand U10866 (N_10866,N_9363,N_6214);
nor U10867 (N_10867,N_7800,N_7404);
or U10868 (N_10868,N_6001,N_9383);
and U10869 (N_10869,N_5588,N_9068);
nand U10870 (N_10870,N_8507,N_9652);
nor U10871 (N_10871,N_8693,N_7108);
nor U10872 (N_10872,N_8053,N_8965);
or U10873 (N_10873,N_6424,N_7105);
or U10874 (N_10874,N_9377,N_5739);
nor U10875 (N_10875,N_9635,N_7219);
or U10876 (N_10876,N_6745,N_9690);
or U10877 (N_10877,N_9630,N_9312);
nand U10878 (N_10878,N_7442,N_6383);
nand U10879 (N_10879,N_7699,N_9019);
and U10880 (N_10880,N_5633,N_8608);
or U10881 (N_10881,N_9868,N_8899);
and U10882 (N_10882,N_7856,N_8293);
nand U10883 (N_10883,N_9933,N_7421);
nand U10884 (N_10884,N_9236,N_8232);
nor U10885 (N_10885,N_9740,N_7684);
or U10886 (N_10886,N_5624,N_6113);
nand U10887 (N_10887,N_8948,N_7240);
nand U10888 (N_10888,N_5939,N_6956);
nand U10889 (N_10889,N_9842,N_5943);
or U10890 (N_10890,N_9962,N_7869);
or U10891 (N_10891,N_9986,N_7430);
nor U10892 (N_10892,N_5109,N_8263);
and U10893 (N_10893,N_9878,N_6283);
nor U10894 (N_10894,N_5843,N_5937);
nor U10895 (N_10895,N_5733,N_8196);
nor U10896 (N_10896,N_6814,N_8784);
and U10897 (N_10897,N_6987,N_8455);
or U10898 (N_10898,N_5487,N_7192);
nand U10899 (N_10899,N_9024,N_7476);
nand U10900 (N_10900,N_8348,N_6503);
nand U10901 (N_10901,N_6594,N_9696);
or U10902 (N_10902,N_6754,N_9143);
and U10903 (N_10903,N_7083,N_9713);
nor U10904 (N_10904,N_8597,N_7485);
nor U10905 (N_10905,N_5223,N_8100);
nor U10906 (N_10906,N_6698,N_8999);
or U10907 (N_10907,N_9892,N_8219);
or U10908 (N_10908,N_9391,N_5560);
nor U10909 (N_10909,N_7115,N_8622);
nand U10910 (N_10910,N_5678,N_6983);
nor U10911 (N_10911,N_9469,N_8332);
nand U10912 (N_10912,N_9725,N_8437);
nand U10913 (N_10913,N_5639,N_9282);
nand U10914 (N_10914,N_8116,N_7397);
or U10915 (N_10915,N_5920,N_5351);
nor U10916 (N_10916,N_6586,N_8192);
nand U10917 (N_10917,N_5571,N_8988);
nor U10918 (N_10918,N_5447,N_9816);
nor U10919 (N_10919,N_8167,N_8729);
nor U10920 (N_10920,N_6678,N_8594);
and U10921 (N_10921,N_8498,N_6338);
nand U10922 (N_10922,N_7500,N_8222);
nand U10923 (N_10923,N_7030,N_7572);
nor U10924 (N_10924,N_6155,N_8615);
nand U10925 (N_10925,N_8577,N_6117);
or U10926 (N_10926,N_5349,N_7303);
or U10927 (N_10927,N_6526,N_8462);
nand U10928 (N_10928,N_6930,N_9208);
nor U10929 (N_10929,N_7526,N_7662);
nand U10930 (N_10930,N_8108,N_6559);
nand U10931 (N_10931,N_7820,N_6029);
or U10932 (N_10932,N_6881,N_9290);
nor U10933 (N_10933,N_5289,N_5556);
nand U10934 (N_10934,N_5585,N_5045);
nor U10935 (N_10935,N_7160,N_5974);
nor U10936 (N_10936,N_8578,N_7698);
nor U10937 (N_10937,N_5648,N_6656);
and U10938 (N_10938,N_9749,N_9720);
and U10939 (N_10939,N_9766,N_6909);
or U10940 (N_10940,N_8470,N_8326);
xnor U10941 (N_10941,N_6051,N_6969);
or U10942 (N_10942,N_6580,N_5726);
or U10943 (N_10943,N_6024,N_7716);
and U10944 (N_10944,N_7836,N_9587);
or U10945 (N_10945,N_9554,N_6726);
or U10946 (N_10946,N_9994,N_9099);
or U10947 (N_10947,N_9259,N_8005);
or U10948 (N_10948,N_7226,N_6262);
nor U10949 (N_10949,N_6616,N_5292);
nor U10950 (N_10950,N_9780,N_7056);
nand U10951 (N_10951,N_6447,N_9598);
and U10952 (N_10952,N_9850,N_7248);
and U10953 (N_10953,N_9093,N_9159);
xnor U10954 (N_10954,N_7809,N_7731);
nand U10955 (N_10955,N_5309,N_8885);
and U10956 (N_10956,N_8685,N_5627);
or U10957 (N_10957,N_9034,N_5517);
and U10958 (N_10958,N_8642,N_9044);
and U10959 (N_10959,N_8181,N_7272);
and U10960 (N_10960,N_5746,N_6618);
or U10961 (N_10961,N_7415,N_7295);
or U10962 (N_10962,N_7902,N_5238);
and U10963 (N_10963,N_5572,N_7361);
and U10964 (N_10964,N_5225,N_7344);
or U10965 (N_10965,N_7050,N_9708);
or U10966 (N_10966,N_7288,N_8273);
nand U10967 (N_10967,N_9787,N_9286);
or U10968 (N_10968,N_7924,N_6257);
nor U10969 (N_10969,N_7933,N_8883);
and U10970 (N_10970,N_7637,N_5027);
and U10971 (N_10971,N_9244,N_5745);
nand U10972 (N_10972,N_7641,N_7486);
nand U10973 (N_10973,N_9856,N_6423);
nand U10974 (N_10974,N_5866,N_9355);
and U10975 (N_10975,N_7591,N_7870);
nand U10976 (N_10976,N_5034,N_5562);
nor U10977 (N_10977,N_7247,N_8633);
or U10978 (N_10978,N_9268,N_9959);
or U10979 (N_10979,N_6138,N_6241);
nand U10980 (N_10980,N_7738,N_5382);
nor U10981 (N_10981,N_8528,N_5934);
nand U10982 (N_10982,N_5286,N_8513);
nand U10983 (N_10983,N_6896,N_8026);
nand U10984 (N_10984,N_9743,N_8013);
nand U10985 (N_10985,N_9776,N_6569);
nand U10986 (N_10986,N_6328,N_5091);
nand U10987 (N_10987,N_9934,N_5160);
nand U10988 (N_10988,N_9188,N_5288);
nor U10989 (N_10989,N_8664,N_9867);
or U10990 (N_10990,N_6784,N_8176);
nand U10991 (N_10991,N_6231,N_6042);
or U10992 (N_10992,N_9272,N_8826);
and U10993 (N_10993,N_5836,N_8008);
nand U10994 (N_10994,N_8137,N_9700);
nor U10995 (N_10995,N_9826,N_9540);
or U10996 (N_10996,N_5591,N_8107);
nor U10997 (N_10997,N_5650,N_5561);
or U10998 (N_10998,N_5661,N_7546);
or U10999 (N_10999,N_5911,N_8721);
or U11000 (N_11000,N_7855,N_5674);
nand U11001 (N_11001,N_5217,N_7034);
nor U11002 (N_11002,N_9597,N_9649);
or U11003 (N_11003,N_6097,N_8911);
and U11004 (N_11004,N_6946,N_5466);
nand U11005 (N_11005,N_7575,N_6187);
or U11006 (N_11006,N_5387,N_7619);
nand U11007 (N_11007,N_8453,N_8901);
nor U11008 (N_11008,N_5758,N_7953);
and U11009 (N_11009,N_6258,N_7298);
nand U11010 (N_11010,N_7092,N_8357);
nor U11011 (N_11011,N_7717,N_8084);
nand U11012 (N_11012,N_6699,N_7537);
or U11013 (N_11013,N_5334,N_5321);
or U11014 (N_11014,N_8889,N_7821);
and U11015 (N_11015,N_9699,N_9722);
nor U11016 (N_11016,N_8449,N_9781);
nand U11017 (N_11017,N_7693,N_7975);
nor U11018 (N_11018,N_8557,N_7832);
nor U11019 (N_11019,N_5232,N_5344);
nand U11020 (N_11020,N_5888,N_9346);
nor U11021 (N_11021,N_7139,N_7791);
or U11022 (N_11022,N_7527,N_9065);
or U11023 (N_11023,N_6941,N_8489);
and U11024 (N_11024,N_6145,N_9012);
nand U11025 (N_11025,N_9928,N_5859);
nor U11026 (N_11026,N_7614,N_9369);
nand U11027 (N_11027,N_5333,N_5717);
or U11028 (N_11028,N_5511,N_7558);
nor U11029 (N_11029,N_7350,N_5154);
and U11030 (N_11030,N_6490,N_5051);
or U11031 (N_11031,N_7585,N_7011);
or U11032 (N_11032,N_9491,N_9166);
nor U11033 (N_11033,N_8118,N_7976);
and U11034 (N_11034,N_6717,N_7650);
or U11035 (N_11035,N_6870,N_7701);
nor U11036 (N_11036,N_6130,N_5916);
nor U11037 (N_11037,N_7308,N_6077);
nor U11038 (N_11038,N_7444,N_9800);
and U11039 (N_11039,N_7306,N_7420);
and U11040 (N_11040,N_5059,N_5751);
nor U11041 (N_11041,N_8492,N_7090);
xor U11042 (N_11042,N_9036,N_6922);
or U11043 (N_11043,N_8317,N_5410);
nor U11044 (N_11044,N_7653,N_7516);
or U11045 (N_11045,N_5715,N_6820);
and U11046 (N_11046,N_5168,N_8520);
or U11047 (N_11047,N_7310,N_6371);
and U11048 (N_11048,N_7700,N_6829);
nand U11049 (N_11049,N_9360,N_6976);
nor U11050 (N_11050,N_8381,N_6644);
or U11051 (N_11051,N_6226,N_5762);
nand U11052 (N_11052,N_5686,N_8709);
and U11053 (N_11053,N_8681,N_6303);
or U11054 (N_11054,N_8407,N_9215);
and U11055 (N_11055,N_8556,N_7625);
or U11056 (N_11056,N_7278,N_5380);
and U11057 (N_11057,N_5817,N_7070);
nand U11058 (N_11058,N_9683,N_9879);
nor U11059 (N_11059,N_5753,N_9097);
nor U11060 (N_11060,N_6640,N_9054);
and U11061 (N_11061,N_6721,N_5284);
and U11062 (N_11062,N_8831,N_8932);
nand U11063 (N_11063,N_5114,N_9315);
or U11064 (N_11064,N_5791,N_6797);
and U11065 (N_11065,N_9654,N_9500);
or U11066 (N_11066,N_7053,N_5617);
nand U11067 (N_11067,N_6592,N_9381);
or U11068 (N_11068,N_6435,N_6702);
and U11069 (N_11069,N_6006,N_7623);
and U11070 (N_11070,N_8177,N_5026);
and U11071 (N_11071,N_7742,N_6468);
nand U11072 (N_11072,N_8061,N_5597);
nor U11073 (N_11073,N_7721,N_6174);
and U11074 (N_11074,N_7589,N_5900);
or U11075 (N_11075,N_6741,N_8892);
or U11076 (N_11076,N_7440,N_5831);
and U11077 (N_11077,N_6676,N_9410);
or U11078 (N_11078,N_6563,N_9340);
and U11079 (N_11079,N_7747,N_8697);
nor U11080 (N_11080,N_5149,N_5096);
nor U11081 (N_11081,N_9658,N_9263);
nand U11082 (N_11082,N_7319,N_8815);
and U11083 (N_11083,N_9755,N_9077);
or U11084 (N_11084,N_7245,N_7179);
xor U11085 (N_11085,N_6886,N_6821);
nor U11086 (N_11086,N_8349,N_6425);
nand U11087 (N_11087,N_5330,N_6344);
nand U11088 (N_11088,N_7932,N_5326);
and U11089 (N_11089,N_5595,N_6637);
and U11090 (N_11090,N_9091,N_7966);
nand U11091 (N_11091,N_6381,N_6851);
nor U11092 (N_11092,N_5929,N_7456);
or U11093 (N_11093,N_6654,N_7371);
or U11094 (N_11094,N_9753,N_7914);
and U11095 (N_11095,N_8220,N_9193);
and U11096 (N_11096,N_6758,N_7131);
and U11097 (N_11097,N_8968,N_8873);
nand U11098 (N_11098,N_5800,N_7364);
or U11099 (N_11099,N_5693,N_9717);
or U11100 (N_11100,N_5761,N_6660);
and U11101 (N_11101,N_9126,N_9552);
or U11102 (N_11102,N_5894,N_9797);
and U11103 (N_11103,N_5784,N_9307);
nor U11104 (N_11104,N_6205,N_9943);
and U11105 (N_11105,N_5037,N_9308);
or U11106 (N_11106,N_5609,N_8097);
or U11107 (N_11107,N_7937,N_8611);
nor U11108 (N_11108,N_7533,N_8951);
or U11109 (N_11109,N_6836,N_9764);
or U11110 (N_11110,N_9336,N_6865);
nand U11111 (N_11111,N_5931,N_5453);
and U11112 (N_11112,N_8139,N_8939);
nand U11113 (N_11113,N_5463,N_5275);
nand U11114 (N_11114,N_7943,N_6647);
nand U11115 (N_11115,N_7909,N_5159);
nand U11116 (N_11116,N_5822,N_8500);
or U11117 (N_11117,N_7463,N_8699);
nor U11118 (N_11118,N_5295,N_7770);
nor U11119 (N_11119,N_8064,N_6436);
and U11120 (N_11120,N_7198,N_7777);
and U11121 (N_11121,N_5117,N_5942);
nor U11122 (N_11122,N_8981,N_9327);
and U11123 (N_11123,N_6619,N_5842);
and U11124 (N_11124,N_8380,N_9636);
nand U11125 (N_11125,N_8090,N_5086);
nand U11126 (N_11126,N_5338,N_9729);
or U11127 (N_11127,N_6317,N_7524);
nor U11128 (N_11128,N_5902,N_9128);
xnor U11129 (N_11129,N_9174,N_8544);
nand U11130 (N_11130,N_7985,N_5534);
and U11131 (N_11131,N_7577,N_9185);
nand U11132 (N_11132,N_8943,N_8687);
and U11133 (N_11133,N_6650,N_9932);
nor U11134 (N_11134,N_8970,N_9571);
nand U11135 (N_11135,N_9931,N_6949);
nand U11136 (N_11136,N_8417,N_6387);
nand U11137 (N_11137,N_6625,N_8750);
nand U11138 (N_11138,N_5432,N_8336);
nor U11139 (N_11139,N_9499,N_7858);
and U11140 (N_11140,N_5236,N_6486);
nor U11141 (N_11141,N_5291,N_8171);
nor U11142 (N_11142,N_5850,N_9663);
nand U11143 (N_11143,N_7579,N_7468);
nand U11144 (N_11144,N_9629,N_9711);
or U11145 (N_11145,N_8480,N_6651);
nor U11146 (N_11146,N_6535,N_6060);
nor U11147 (N_11147,N_5704,N_6566);
or U11148 (N_11148,N_5492,N_9734);
or U11149 (N_11149,N_7367,N_8617);
and U11150 (N_11150,N_5578,N_8036);
or U11151 (N_11151,N_9304,N_9368);
nand U11152 (N_11152,N_5467,N_5816);
and U11153 (N_11153,N_8692,N_7460);
and U11154 (N_11154,N_7612,N_6521);
nor U11155 (N_11155,N_5264,N_5322);
and U11156 (N_11156,N_6613,N_7903);
or U11157 (N_11157,N_7757,N_5664);
and U11158 (N_11158,N_7818,N_8284);
and U11159 (N_11159,N_7464,N_9121);
xnor U11160 (N_11160,N_7447,N_8776);
and U11161 (N_11161,N_5921,N_6349);
or U11162 (N_11162,N_5398,N_9758);
or U11163 (N_11163,N_5031,N_6443);
nor U11164 (N_11164,N_8210,N_6268);
nor U11165 (N_11165,N_7202,N_9021);
nor U11166 (N_11166,N_6665,N_5002);
and U11167 (N_11167,N_6785,N_9710);
and U11168 (N_11168,N_9281,N_7326);
and U11169 (N_11169,N_8099,N_9241);
or U11170 (N_11170,N_7963,N_9194);
or U11171 (N_11171,N_7000,N_6890);
nand U11172 (N_11172,N_5446,N_5116);
xnor U11173 (N_11173,N_5905,N_7436);
and U11174 (N_11174,N_7792,N_7898);
nand U11175 (N_11175,N_6159,N_5584);
nor U11176 (N_11176,N_7664,N_8430);
nor U11177 (N_11177,N_8367,N_9309);
nor U11178 (N_11178,N_8276,N_9445);
nand U11179 (N_11179,N_7538,N_6763);
nand U11180 (N_11180,N_9756,N_5054);
and U11181 (N_11181,N_5370,N_7123);
nor U11182 (N_11182,N_6068,N_8032);
xor U11183 (N_11183,N_6507,N_8521);
or U11184 (N_11184,N_9557,N_5870);
nor U11185 (N_11185,N_7797,N_7919);
xor U11186 (N_11186,N_9413,N_9594);
or U11187 (N_11187,N_5799,N_7871);
nor U11188 (N_11188,N_8441,N_5512);
nor U11189 (N_11189,N_7776,N_6585);
and U11190 (N_11190,N_5437,N_7106);
or U11191 (N_11191,N_7164,N_9142);
nor U11192 (N_11192,N_9693,N_6971);
or U11193 (N_11193,N_6484,N_7847);
nand U11194 (N_11194,N_9803,N_5689);
nand U11195 (N_11195,N_8650,N_7555);
nor U11196 (N_11196,N_5697,N_8896);
nor U11197 (N_11197,N_8159,N_7315);
and U11198 (N_11198,N_5925,N_6003);
nor U11199 (N_11199,N_8982,N_5032);
nand U11200 (N_11200,N_8149,N_9513);
and U11201 (N_11201,N_8190,N_6912);
nand U11202 (N_11202,N_9822,N_6475);
or U11203 (N_11203,N_5371,N_8559);
nor U11204 (N_11204,N_5393,N_6111);
or U11205 (N_11205,N_7512,N_8174);
or U11206 (N_11206,N_8010,N_9452);
and U11207 (N_11207,N_5757,N_7918);
xnor U11208 (N_11208,N_5809,N_5801);
or U11209 (N_11209,N_8345,N_7980);
xor U11210 (N_11210,N_8670,N_5646);
nand U11211 (N_11211,N_5259,N_8915);
or U11212 (N_11212,N_8610,N_9643);
or U11213 (N_11213,N_9147,N_6955);
or U11214 (N_11214,N_6445,N_7930);
nor U11215 (N_11215,N_6110,N_9769);
nand U11216 (N_11216,N_5785,N_8153);
or U11217 (N_11217,N_6455,N_9977);
xor U11218 (N_11218,N_9726,N_5846);
or U11219 (N_11219,N_5413,N_6895);
or U11220 (N_11220,N_7972,N_6950);
nor U11221 (N_11221,N_8625,N_7974);
or U11222 (N_11222,N_9490,N_5176);
nor U11223 (N_11223,N_7722,N_6992);
and U11224 (N_11224,N_9431,N_5213);
and U11225 (N_11225,N_5206,N_5790);
nand U11226 (N_11226,N_6945,N_6150);
xor U11227 (N_11227,N_8806,N_6841);
or U11228 (N_11228,N_7010,N_5892);
nand U11229 (N_11229,N_8017,N_7178);
and U11230 (N_11230,N_9520,N_8135);
nand U11231 (N_11231,N_9257,N_6928);
and U11232 (N_11232,N_8472,N_6370);
nand U11233 (N_11233,N_7323,N_5496);
and U11234 (N_11234,N_9164,N_6782);
nor U11235 (N_11235,N_6465,N_8085);
or U11236 (N_11236,N_6167,N_8651);
and U11237 (N_11237,N_7565,N_8335);
xor U11238 (N_11238,N_8898,N_9846);
nand U11239 (N_11239,N_6166,N_7282);
or U11240 (N_11240,N_5616,N_8950);
nor U11241 (N_11241,N_9579,N_9980);
and U11242 (N_11242,N_8961,N_7291);
or U11243 (N_11243,N_7633,N_6207);
or U11244 (N_11244,N_7793,N_7209);
nor U11245 (N_11245,N_7402,N_7265);
or U11246 (N_11246,N_5443,N_6417);
nor U11247 (N_11247,N_8548,N_9486);
or U11248 (N_11248,N_7687,N_5666);
nor U11249 (N_11249,N_9517,N_9965);
or U11250 (N_11250,N_7244,N_6279);
nor U11251 (N_11251,N_9588,N_5337);
or U11252 (N_11252,N_7498,N_9678);
nand U11253 (N_11253,N_9026,N_5479);
or U11254 (N_11254,N_9212,N_7859);
nor U11255 (N_11255,N_9478,N_6073);
xnor U11256 (N_11256,N_5003,N_7232);
and U11257 (N_11257,N_7346,N_8616);
nor U11258 (N_11258,N_9129,N_5087);
nor U11259 (N_11259,N_7072,N_9983);
and U11260 (N_11260,N_6312,N_6925);
nand U11261 (N_11261,N_7324,N_9028);
nand U11262 (N_11262,N_7718,N_9140);
or U11263 (N_11263,N_8451,N_8958);
or U11264 (N_11264,N_9379,N_8974);
or U11265 (N_11265,N_6418,N_9669);
nand U11266 (N_11266,N_5839,N_5365);
or U11267 (N_11267,N_7690,N_5978);
nor U11268 (N_11268,N_9243,N_5210);
nor U11269 (N_11269,N_7992,N_8213);
nand U11270 (N_11270,N_7038,N_8382);
or U11271 (N_11271,N_8977,N_7948);
nand U11272 (N_11272,N_7330,N_8569);
or U11273 (N_11273,N_6612,N_7443);
xor U11274 (N_11274,N_6058,N_9872);
and U11275 (N_11275,N_8120,N_6310);
nand U11276 (N_11276,N_9430,N_9069);
nand U11277 (N_11277,N_9137,N_5952);
and U11278 (N_11278,N_5777,N_5035);
nor U11279 (N_11279,N_6120,N_6089);
nand U11280 (N_11280,N_8092,N_8657);
or U11281 (N_11281,N_9998,N_7049);
xnor U11282 (N_11282,N_8671,N_5844);
nor U11283 (N_11283,N_5345,N_5403);
nand U11284 (N_11284,N_9662,N_7551);
nand U11285 (N_11285,N_7563,N_6624);
or U11286 (N_11286,N_5056,N_5838);
and U11287 (N_11287,N_8347,N_9814);
nand U11288 (N_11288,N_8639,N_6453);
or U11289 (N_11289,N_5857,N_9930);
nand U11290 (N_11290,N_8029,N_6482);
nor U11291 (N_11291,N_8298,N_7874);
and U11292 (N_11292,N_8050,N_8819);
or U11293 (N_11293,N_9724,N_6750);
nor U11294 (N_11294,N_6587,N_7407);
and U11295 (N_11295,N_8938,N_5111);
xor U11296 (N_11296,N_9248,N_8456);
and U11297 (N_11297,N_7939,N_8574);
nand U11298 (N_11298,N_8789,N_5278);
nand U11299 (N_11299,N_9676,N_8102);
nor U11300 (N_11300,N_7865,N_9891);
or U11301 (N_11301,N_6853,N_7488);
or U11302 (N_11302,N_7596,N_5094);
nor U11303 (N_11303,N_6131,N_5315);
xnor U11304 (N_11304,N_5967,N_6934);
or U11305 (N_11305,N_7112,N_8362);
nor U11306 (N_11306,N_8875,N_5720);
and U11307 (N_11307,N_6818,N_8476);
nand U11308 (N_11308,N_5930,N_8830);
or U11309 (N_11309,N_9314,N_8067);
nor U11310 (N_11310,N_9595,N_6388);
nor U11311 (N_11311,N_5397,N_7377);
nor U11312 (N_11312,N_9150,N_8791);
and U11313 (N_11313,N_6061,N_5695);
or U11314 (N_11314,N_5835,N_5980);
and U11315 (N_11315,N_6067,N_9275);
nor U11316 (N_11316,N_6266,N_8736);
and U11317 (N_11317,N_8000,N_8547);
nand U11318 (N_11318,N_8446,N_9224);
nand U11319 (N_11319,N_7084,N_8077);
and U11320 (N_11320,N_7724,N_9733);
or U11321 (N_11321,N_9030,N_7195);
nand U11322 (N_11322,N_7887,N_7230);
and U11323 (N_11323,N_6457,N_7807);
nand U11324 (N_11324,N_8063,N_5299);
or U11325 (N_11325,N_6083,N_7411);
or U11326 (N_11326,N_9799,N_9673);
nand U11327 (N_11327,N_9323,N_8388);
nand U11328 (N_11328,N_5454,N_8652);
nand U11329 (N_11329,N_9632,N_9840);
or U11330 (N_11330,N_5737,N_8865);
or U11331 (N_11331,N_9607,N_9179);
or U11332 (N_11332,N_5682,N_8747);
and U11333 (N_11333,N_7735,N_8080);
nand U11334 (N_11334,N_6169,N_6403);
nor U11335 (N_11335,N_8715,N_8540);
and U11336 (N_11336,N_6847,N_6101);
or U11337 (N_11337,N_7381,N_6749);
nand U11338 (N_11338,N_7714,N_5815);
nor U11339 (N_11339,N_8575,N_8598);
and U11340 (N_11340,N_6034,N_8308);
and U11341 (N_11341,N_8869,N_5631);
or U11342 (N_11342,N_6242,N_7507);
and U11343 (N_11343,N_5723,N_5885);
and U11344 (N_11344,N_9322,N_8404);
nand U11345 (N_11345,N_9345,N_8305);
and U11346 (N_11346,N_8607,N_5763);
nand U11347 (N_11347,N_6322,N_7556);
nor U11348 (N_11348,N_5457,N_9420);
or U11349 (N_11349,N_8711,N_9462);
nor U11350 (N_11350,N_6270,N_7388);
or U11351 (N_11351,N_6529,N_7549);
nor U11352 (N_11352,N_5958,N_6017);
and U11353 (N_11353,N_6757,N_5191);
or U11354 (N_11354,N_6907,N_9626);
and U11355 (N_11355,N_8506,N_5837);
nor U11356 (N_11356,N_8839,N_8679);
and U11357 (N_11357,N_8661,N_5659);
nand U11358 (N_11358,N_6476,N_6019);
nand U11359 (N_11359,N_7586,N_7009);
nand U11360 (N_11360,N_5989,N_6350);
and U11361 (N_11361,N_9329,N_8285);
nor U11362 (N_11362,N_6812,N_9103);
and U11363 (N_11363,N_9071,N_9086);
nor U11364 (N_11364,N_8130,N_7604);
nor U11365 (N_11365,N_7550,N_7849);
and U11366 (N_11366,N_7055,N_8864);
nor U11367 (N_11367,N_9604,N_6834);
and U11368 (N_11368,N_6023,N_8186);
nor U11369 (N_11369,N_9181,N_9589);
nand U11370 (N_11370,N_8876,N_7366);
or U11371 (N_11371,N_6239,N_5736);
nor U11372 (N_11372,N_9416,N_9999);
or U11373 (N_11373,N_6440,N_7142);
and U11374 (N_11374,N_8268,N_9085);
nor U11375 (N_11375,N_5547,N_6264);
and U11376 (N_11376,N_5192,N_8491);
nand U11377 (N_11377,N_8478,N_6501);
nand U11378 (N_11378,N_7193,N_8870);
nand U11379 (N_11379,N_9395,N_7584);
xnor U11380 (N_11380,N_5969,N_8584);
nand U11381 (N_11381,N_8215,N_8200);
nor U11382 (N_11382,N_7863,N_8545);
nand U11383 (N_11383,N_7908,N_8020);
xor U11384 (N_11384,N_8228,N_7854);
and U11385 (N_11385,N_7429,N_8327);
and U11386 (N_11386,N_7236,N_5414);
and U11387 (N_11387,N_5390,N_7983);
or U11388 (N_11388,N_9100,N_8211);
nor U11389 (N_11389,N_8956,N_7893);
nor U11390 (N_11390,N_6188,N_6376);
nor U11391 (N_11391,N_5971,N_7670);
nor U11392 (N_11392,N_5011,N_8275);
nor U11393 (N_11393,N_6139,N_9905);
nand U11394 (N_11394,N_5570,N_9390);
and U11395 (N_11395,N_5362,N_6337);
nor U11396 (N_11396,N_8197,N_5621);
nand U11397 (N_11397,N_8923,N_9682);
nor U11398 (N_11398,N_6849,N_6152);
and U11399 (N_11399,N_8546,N_7539);
and U11400 (N_11400,N_5657,N_8412);
nand U11401 (N_11401,N_9081,N_8238);
nand U11402 (N_11402,N_8350,N_7266);
and U11403 (N_11403,N_7624,N_6252);
nor U11404 (N_11404,N_7078,N_6805);
or U11405 (N_11405,N_5529,N_9973);
or U11406 (N_11406,N_5963,N_9405);
or U11407 (N_11407,N_8203,N_5392);
nor U11408 (N_11408,N_8937,N_5546);
xor U11409 (N_11409,N_5036,N_8337);
nand U11410 (N_11410,N_9398,N_9460);
and U11411 (N_11411,N_7929,N_8647);
or U11412 (N_11412,N_7165,N_5074);
or U11413 (N_11413,N_8113,N_6497);
nand U11414 (N_11414,N_5138,N_5601);
or U11415 (N_11415,N_9553,N_5898);
and U11416 (N_11416,N_6059,N_8287);
and U11417 (N_11417,N_9783,N_5200);
nor U11418 (N_11418,N_5810,N_9785);
or U11419 (N_11419,N_5807,N_9288);
nand U11420 (N_11420,N_6842,N_7768);
nand U11421 (N_11421,N_7951,N_9204);
and U11422 (N_11422,N_6129,N_7782);
or U11423 (N_11423,N_9820,N_7379);
nor U11424 (N_11424,N_5269,N_8542);
and U11425 (N_11425,N_9542,N_5598);
nor U11426 (N_11426,N_8987,N_9918);
and U11427 (N_11427,N_9707,N_6952);
and U11428 (N_11428,N_9376,N_5600);
and U11429 (N_11429,N_9184,N_6206);
or U11430 (N_11430,N_5523,N_6855);
or U11431 (N_11431,N_9702,N_8216);
or U11432 (N_11432,N_9655,N_5909);
nor U11433 (N_11433,N_7896,N_7269);
nor U11434 (N_11434,N_7060,N_9213);
or U11435 (N_11435,N_8935,N_9182);
nor U11436 (N_11436,N_8078,N_9809);
and U11437 (N_11437,N_9267,N_6329);
nand U11438 (N_11438,N_6825,N_8813);
nor U11439 (N_11439,N_7333,N_8074);
or U11440 (N_11440,N_6576,N_7362);
or U11441 (N_11441,N_8454,N_6629);
nor U11442 (N_11442,N_7229,N_8573);
or U11443 (N_11443,N_9825,N_9531);
nand U11444 (N_11444,N_6762,N_9471);
nor U11445 (N_11445,N_6680,N_7252);
nor U11446 (N_11446,N_7982,N_9889);
and U11447 (N_11447,N_8638,N_9448);
or U11448 (N_11448,N_7041,N_5214);
and U11449 (N_11449,N_7741,N_7795);
and U11450 (N_11450,N_5869,N_7928);
nor U11451 (N_11451,N_8718,N_8175);
or U11452 (N_11452,N_8596,N_5205);
nor U11453 (N_11453,N_8576,N_8841);
nand U11454 (N_11454,N_6473,N_9242);
or U11455 (N_11455,N_7222,N_8049);
and U11456 (N_11456,N_6112,N_5786);
and U11457 (N_11457,N_6894,N_5811);
xor U11458 (N_11458,N_8934,N_6608);
nor U11459 (N_11459,N_6127,N_6711);
and U11460 (N_11460,N_7765,N_6409);
xnor U11461 (N_11461,N_8021,N_7881);
nor U11462 (N_11462,N_9387,N_7643);
and U11463 (N_11463,N_5516,N_7365);
and U11464 (N_11464,N_7892,N_9037);
nand U11465 (N_11465,N_5007,N_9187);
nor U11466 (N_11466,N_5233,N_9657);
nor U11467 (N_11467,N_5675,N_8178);
nand U11468 (N_11468,N_5290,N_9622);
nand U11469 (N_11469,N_9777,N_9191);
and U11470 (N_11470,N_8746,N_6133);
and U11471 (N_11471,N_6351,N_9459);
or U11472 (N_11472,N_8705,N_7018);
nor U11473 (N_11473,N_9453,N_5316);
nand U11474 (N_11474,N_7399,N_7824);
nor U11475 (N_11475,N_7337,N_9773);
and U11476 (N_11476,N_8098,N_5434);
and U11477 (N_11477,N_9616,N_6843);
and U11478 (N_11478,N_7480,N_9173);
xnor U11479 (N_11479,N_5384,N_6074);
and U11480 (N_11480,N_6500,N_7566);
and U11481 (N_11481,N_6796,N_6379);
or U11482 (N_11482,N_6574,N_6615);
nor U11483 (N_11483,N_8631,N_7580);
nand U11484 (N_11484,N_6389,N_5893);
nor U11485 (N_11485,N_6200,N_6653);
nand U11486 (N_11486,N_8920,N_6261);
or U11487 (N_11487,N_6428,N_5983);
nand U11488 (N_11488,N_9631,N_6875);
and U11489 (N_11489,N_6538,N_7471);
and U11490 (N_11490,N_9937,N_8241);
or U11491 (N_11491,N_5488,N_6816);
xor U11492 (N_11492,N_7276,N_7790);
nor U11493 (N_11493,N_7582,N_5241);
and U11494 (N_11494,N_9492,N_7905);
or U11495 (N_11495,N_7560,N_8076);
and U11496 (N_11496,N_6630,N_7237);
and U11497 (N_11497,N_6244,N_7327);
or U11498 (N_11498,N_8866,N_8884);
nand U11499 (N_11499,N_5014,N_9022);
or U11500 (N_11500,N_9996,N_5012);
or U11501 (N_11501,N_7878,N_9284);
nor U11502 (N_11502,N_6463,N_8363);
nand U11503 (N_11503,N_8942,N_8296);
nor U11504 (N_11504,N_9830,N_9354);
or U11505 (N_11505,N_6190,N_9498);
nand U11506 (N_11506,N_6893,N_7325);
or U11507 (N_11507,N_7990,N_9745);
and U11508 (N_11508,N_5948,N_9821);
nand U11509 (N_11509,N_8403,N_7203);
nor U11510 (N_11510,N_7110,N_6075);
and U11511 (N_11511,N_7666,N_8214);
nor U11512 (N_11512,N_5480,N_8234);
xor U11513 (N_11513,N_6132,N_5374);
or U11514 (N_11514,N_9096,N_7846);
nand U11515 (N_11515,N_6860,N_7243);
or U11516 (N_11516,N_9529,N_7588);
nand U11517 (N_11517,N_8566,N_6406);
and U11518 (N_11518,N_5048,N_6631);
nor U11519 (N_11519,N_5255,N_8165);
nor U11520 (N_11520,N_7600,N_6454);
and U11521 (N_11521,N_7736,N_9893);
xor U11522 (N_11522,N_7576,N_6747);
or U11523 (N_11523,N_8205,N_7210);
or U11524 (N_11524,N_8414,N_8034);
or U11525 (N_11525,N_6459,N_8534);
or U11526 (N_11526,N_7204,N_6931);
nor U11527 (N_11527,N_9875,N_6550);
or U11528 (N_11528,N_9196,N_6163);
nand U11529 (N_11529,N_8148,N_8237);
nor U11530 (N_11530,N_7188,N_6792);
nand U11531 (N_11531,N_6776,N_5070);
nand U11532 (N_11532,N_6301,N_6707);
nor U11533 (N_11533,N_7819,N_8572);
nor U11534 (N_11534,N_6161,N_7862);
nand U11535 (N_11535,N_7259,N_6367);
or U11536 (N_11536,N_5144,N_6298);
nand U11537 (N_11537,N_7987,N_9802);
or U11538 (N_11538,N_5356,N_8447);
nor U11539 (N_11539,N_5856,N_7274);
nor U11540 (N_11540,N_6063,N_8567);
or U11541 (N_11541,N_9765,N_8212);
and U11542 (N_11542,N_8475,N_9603);
nand U11543 (N_11543,N_7689,N_7120);
nand U11544 (N_11544,N_8962,N_7530);
and U11545 (N_11545,N_5672,N_6512);
nand U11546 (N_11546,N_7636,N_8054);
nand U11547 (N_11547,N_5873,N_5788);
or U11548 (N_11548,N_7196,N_5139);
nand U11549 (N_11549,N_8605,N_9003);
nor U11550 (N_11550,N_7128,N_6568);
nor U11551 (N_11551,N_7121,N_9320);
and U11552 (N_11552,N_7089,N_6787);
xnor U11553 (N_11553,N_7787,N_7423);
nor U11554 (N_11554,N_6072,N_6086);
nand U11555 (N_11555,N_5632,N_7263);
nand U11556 (N_11556,N_8909,N_5528);
and U11557 (N_11557,N_8106,N_5220);
nand U11558 (N_11558,N_8247,N_7452);
nor U11559 (N_11559,N_9441,N_7646);
nor U11560 (N_11560,N_9610,N_6265);
nor U11561 (N_11561,N_5824,N_7416);
and U11562 (N_11562,N_5433,N_5419);
nor U11563 (N_11563,N_8041,N_8223);
xor U11564 (N_11564,N_5703,N_7051);
nand U11565 (N_11565,N_6027,N_5285);
nand U11566 (N_11566,N_5579,N_5240);
and U11567 (N_11567,N_7418,N_7772);
or U11568 (N_11568,N_6354,N_9160);
nand U11569 (N_11569,N_9247,N_6710);
or U11570 (N_11570,N_6122,N_9865);
and U11571 (N_11571,N_6412,N_8930);
or U11572 (N_11572,N_9331,N_7967);
and U11573 (N_11573,N_6835,N_9602);
nand U11574 (N_11574,N_9853,N_8343);
nor U11575 (N_11575,N_8089,N_8564);
nand U11576 (N_11576,N_8768,N_7225);
and U11577 (N_11577,N_9487,N_6819);
or U11578 (N_11578,N_7706,N_7755);
or U11579 (N_11579,N_5797,N_6815);
or U11580 (N_11580,N_8908,N_9392);
nand U11581 (N_11581,N_6196,N_8552);
nand U11582 (N_11582,N_8321,N_9371);
nor U11583 (N_11583,N_8283,N_9238);
nand U11584 (N_11584,N_7279,N_5552);
nor U11585 (N_11585,N_5179,N_6916);
nor U11586 (N_11586,N_8758,N_9503);
nand U11587 (N_11587,N_6336,N_5171);
nand U11588 (N_11588,N_8959,N_7904);
nand U11589 (N_11589,N_7075,N_9763);
and U11590 (N_11590,N_7163,N_7649);
nor U11591 (N_11591,N_5358,N_7168);
and U11592 (N_11592,N_5158,N_6116);
nor U11593 (N_11593,N_9439,N_6036);
nand U11594 (N_11594,N_9979,N_7314);
or U11595 (N_11595,N_8960,N_8926);
and U11596 (N_11596,N_6235,N_7312);
and U11597 (N_11597,N_7241,N_9687);
and U11598 (N_11598,N_8997,N_6090);
and U11599 (N_11599,N_7509,N_6984);
or U11600 (N_11600,N_8075,N_8991);
and U11601 (N_11601,N_5364,N_9251);
nor U11602 (N_11602,N_8771,N_7152);
or U11603 (N_11603,N_8334,N_9581);
nor U11604 (N_11604,N_7511,N_8259);
nor U11605 (N_11605,N_5596,N_5459);
nand U11606 (N_11606,N_6696,N_5612);
nor U11607 (N_11607,N_8487,N_5981);
nand U11608 (N_11608,N_6852,N_9484);
xor U11609 (N_11609,N_5253,N_6456);
nor U11610 (N_11610,N_8802,N_6091);
and U11611 (N_11611,N_8244,N_5400);
and U11612 (N_11612,N_9409,N_5438);
nor U11613 (N_11613,N_8565,N_6125);
and U11614 (N_11614,N_9465,N_8678);
nor U11615 (N_11615,N_7264,N_9399);
nor U11616 (N_11616,N_8023,N_7162);
and U11617 (N_11617,N_7412,N_8929);
and U11618 (N_11618,N_6487,N_5352);
and U11619 (N_11619,N_6826,N_6824);
nor U11620 (N_11620,N_8356,N_5427);
and U11621 (N_11621,N_7144,N_8635);
and U11622 (N_11622,N_6182,N_7403);
nor U11623 (N_11623,N_6822,N_6291);
nor U11624 (N_11624,N_9015,N_5976);
and U11625 (N_11625,N_7181,N_7032);
nand U11626 (N_11626,N_6823,N_7595);
nand U11627 (N_11627,N_9059,N_9082);
or U11628 (N_11628,N_8881,N_9104);
or U11629 (N_11629,N_7434,N_7338);
or U11630 (N_11630,N_5460,N_8964);
nand U11631 (N_11631,N_6325,N_8469);
nor U11632 (N_11632,N_8119,N_6936);
xnor U11633 (N_11633,N_8543,N_5444);
or U11634 (N_11634,N_7833,N_7658);
nand U11635 (N_11635,N_6400,N_6596);
nand U11636 (N_11636,N_8833,N_6778);
nand U11637 (N_11637,N_6511,N_9260);
or U11638 (N_11638,N_9330,N_8243);
nand U11639 (N_11639,N_7621,N_7857);
nand U11640 (N_11640,N_6597,N_9380);
nor U11641 (N_11641,N_7320,N_9370);
or U11642 (N_11642,N_7261,N_7891);
or U11643 (N_11643,N_5230,N_8727);
xnor U11644 (N_11644,N_8843,N_8112);
or U11645 (N_11645,N_9960,N_6691);
nand U11646 (N_11646,N_6638,N_7081);
or U11647 (N_11647,N_6938,N_8152);
nand U11648 (N_11648,N_5341,N_9858);
nor U11649 (N_11649,N_8646,N_7359);
nor U11650 (N_11650,N_7100,N_7007);
or U11651 (N_11651,N_5272,N_6639);
nand U11652 (N_11652,N_6366,N_5575);
nand U11653 (N_11653,N_8634,N_5688);
nand U11654 (N_11654,N_9249,N_6153);
nand U11655 (N_11655,N_5796,N_7242);
nor U11656 (N_11656,N_8847,N_6633);
nand U11657 (N_11657,N_6355,N_7391);
nor U11658 (N_11658,N_7231,N_8834);
and U11659 (N_11659,N_8452,N_7564);
and U11660 (N_11660,N_8060,N_7171);
and U11661 (N_11661,N_6742,N_8781);
nor U11662 (N_11662,N_7385,N_5038);
nor U11663 (N_11663,N_7888,N_8541);
and U11664 (N_11664,N_9447,N_9608);
nand U11665 (N_11665,N_7026,N_9712);
nor U11666 (N_11666,N_9650,N_8428);
or U11667 (N_11667,N_9415,N_9586);
xnor U11668 (N_11668,N_7605,N_8473);
nor U11669 (N_11669,N_7629,N_6968);
or U11670 (N_11670,N_9444,N_7781);
nor U11671 (N_11671,N_5472,N_5765);
nor U11672 (N_11672,N_7166,N_8895);
nand U11673 (N_11673,N_8255,N_7680);
nor U11674 (N_11674,N_9738,N_5719);
and U11675 (N_11675,N_6361,N_7194);
nor U11676 (N_11676,N_6972,N_9131);
nand U11677 (N_11677,N_9271,N_9494);
or U11678 (N_11678,N_9599,N_9956);
or U11679 (N_11679,N_5431,N_7598);
nand U11680 (N_11680,N_7732,N_7492);
nor U11681 (N_11681,N_8415,N_5023);
and U11682 (N_11682,N_6947,N_5022);
and U11683 (N_11683,N_5543,N_6037);
or U11684 (N_11684,N_9252,N_5798);
or U11685 (N_11685,N_7098,N_8201);
and U11686 (N_11686,N_6804,N_5136);
and U11687 (N_11687,N_9417,N_6641);
and U11688 (N_11688,N_5115,N_8505);
nand U11689 (N_11689,N_9197,N_9190);
or U11690 (N_11690,N_9902,N_8014);
nand U11691 (N_11691,N_8688,N_7804);
xnor U11692 (N_11692,N_7213,N_7519);
and U11693 (N_11693,N_9339,N_5147);
nor U11694 (N_11694,N_6136,N_9675);
nand U11695 (N_11695,N_9859,N_6493);
nor U11696 (N_11696,N_5676,N_8431);
or U11697 (N_11697,N_7096,N_6873);
or U11698 (N_11698,N_7922,N_5140);
nor U11699 (N_11699,N_9497,N_6183);
and U11700 (N_11700,N_9805,N_7805);
xnor U11701 (N_11701,N_7597,N_7729);
nor U11702 (N_11702,N_8728,N_8122);
nor U11703 (N_11703,N_6534,N_5605);
nand U11704 (N_11704,N_9954,N_7290);
nor U11705 (N_11705,N_5982,N_6031);
nor U11706 (N_11706,N_6168,N_9127);
nand U11707 (N_11707,N_5828,N_6087);
nand U11708 (N_11708,N_8231,N_7620);
and U11709 (N_11709,N_7998,N_8587);
and U11710 (N_11710,N_8140,N_9547);
nor U11711 (N_11711,N_7224,N_5986);
and U11712 (N_11712,N_5282,N_7054);
xor U11713 (N_11713,N_8405,N_8164);
or U11714 (N_11714,N_9328,N_7529);
nand U11715 (N_11715,N_5972,N_9073);
nor U11716 (N_11716,N_6411,N_5890);
nor U11717 (N_11717,N_7608,N_7688);
or U11718 (N_11718,N_6478,N_6012);
nand U11719 (N_11719,N_9018,N_6000);
or U11720 (N_11720,N_9134,N_9228);
nor U11721 (N_11721,N_9835,N_7336);
nor U11722 (N_11722,N_7487,N_5353);
and U11723 (N_11723,N_9335,N_5510);
and U11724 (N_11724,N_5246,N_8751);
nand U11725 (N_11725,N_6731,N_9836);
or U11726 (N_11726,N_7250,N_8239);
and U11727 (N_11727,N_9283,N_7681);
nor U11728 (N_11728,N_8424,N_5908);
or U11729 (N_11729,N_6259,N_8536);
nand U11730 (N_11730,N_6914,N_5854);
nand U11731 (N_11731,N_9438,N_6604);
nor U11732 (N_11732,N_6995,N_8325);
and U11733 (N_11733,N_9480,N_5198);
or U11734 (N_11734,N_5190,N_5157);
nor U11735 (N_11735,N_6348,N_5131);
nor U11736 (N_11736,N_6151,N_7389);
or U11737 (N_11737,N_5783,N_8202);
nor U11738 (N_11738,N_6579,N_9397);
nand U11739 (N_11739,N_9744,N_8967);
nand U11740 (N_11740,N_5262,N_9366);
nand U11741 (N_11741,N_7839,N_5767);
nand U11742 (N_11742,N_9514,N_5766);
and U11743 (N_11743,N_6470,N_9522);
nand U11744 (N_11744,N_8589,N_9951);
nand U11745 (N_11745,N_5610,N_6040);
and U11746 (N_11746,N_7574,N_6530);
or U11747 (N_11747,N_6703,N_7946);
or U11748 (N_11748,N_8629,N_6977);
or U11749 (N_11749,N_9132,N_6296);
nor U11750 (N_11750,N_5474,N_7074);
nor U11751 (N_11751,N_7583,N_7920);
and U11752 (N_11752,N_6346,N_8047);
and U11753 (N_11753,N_6041,N_7837);
and U11754 (N_11754,N_8501,N_8648);
nand U11755 (N_11755,N_8184,N_5992);
nand U11756 (N_11756,N_5260,N_5462);
nor U11757 (N_11757,N_7567,N_5104);
or U11758 (N_11758,N_6466,N_9220);
nand U11759 (N_11759,N_5428,N_7137);
or U11760 (N_11760,N_9107,N_7307);
or U11761 (N_11761,N_6986,N_5097);
nand U11762 (N_11762,N_5574,N_9177);
nor U11763 (N_11763,N_9870,N_8161);
nand U11764 (N_11764,N_5904,N_6704);
nand U11765 (N_11765,N_6057,N_6331);
nor U11766 (N_11766,N_8399,N_8278);
and U11767 (N_11767,N_6864,N_9133);
or U11768 (N_11768,N_8502,N_6356);
nor U11769 (N_11769,N_8832,N_7786);
nand U11770 (N_11770,N_7457,N_8512);
or U11771 (N_11771,N_9384,N_6410);
nand U11772 (N_11772,N_5229,N_5953);
nand U11773 (N_11773,N_5277,N_7986);
and U11774 (N_11774,N_6140,N_5852);
nor U11775 (N_11775,N_6353,N_8739);
nand U11776 (N_11776,N_5378,N_6398);
nand U11777 (N_11777,N_9511,N_6774);
and U11778 (N_11778,N_5770,N_6794);
nand U11779 (N_11779,N_5564,N_5589);
and U11780 (N_11780,N_6924,N_7970);
nor U11781 (N_11781,N_6340,N_6970);
and U11782 (N_11782,N_5436,N_6197);
nand U11783 (N_11783,N_9585,N_7122);
or U11784 (N_11784,N_9625,N_7390);
nor U11785 (N_11785,N_6452,N_7949);
nand U11786 (N_11786,N_7815,N_5348);
nor U11787 (N_11787,N_5884,N_8314);
and U11788 (N_11788,N_8745,N_7799);
nor U11789 (N_11789,N_7789,N_8533);
and U11790 (N_11790,N_9591,N_6286);
nor U11791 (N_11791,N_5452,N_5861);
nor U11792 (N_11792,N_5741,N_6444);
and U11793 (N_11793,N_8659,N_9211);
nor U11794 (N_11794,N_7610,N_6687);
or U11795 (N_11795,N_8422,N_7829);
nand U11796 (N_11796,N_6962,N_7173);
or U11797 (N_11797,N_5896,N_9115);
and U11798 (N_11798,N_9079,N_8531);
or U11799 (N_11799,N_9233,N_5391);
nor U11800 (N_11800,N_9735,N_6693);
nor U11801 (N_11801,N_6727,N_6246);
or U11802 (N_11802,N_7126,N_8369);
nand U11803 (N_11803,N_9464,N_9214);
or U11804 (N_11804,N_5323,N_8769);
nor U11805 (N_11805,N_8522,N_6126);
nor U11806 (N_11806,N_6438,N_8621);
nor U11807 (N_11807,N_8307,N_7466);
and U11808 (N_11808,N_7355,N_8299);
nor U11809 (N_11809,N_8096,N_9523);
nand U11810 (N_11810,N_7901,N_8509);
and U11811 (N_11811,N_8640,N_6413);
or U11812 (N_11812,N_9873,N_9572);
and U11813 (N_11813,N_8775,N_7066);
nand U11814 (N_11814,N_9982,N_9078);
or U11815 (N_11815,N_6570,N_6974);
nand U11816 (N_11816,N_7186,N_7021);
nand U11817 (N_11817,N_5853,N_5415);
or U11818 (N_11818,N_9617,N_6684);
nor U11819 (N_11819,N_7400,N_7146);
or U11820 (N_11820,N_9596,N_6256);
nand U11821 (N_11821,N_9326,N_8359);
or U11822 (N_11822,N_6957,N_6502);
and U11823 (N_11823,N_9265,N_6541);
xor U11824 (N_11824,N_5129,N_5039);
and U11825 (N_11825,N_9698,N_8062);
nor U11826 (N_11826,N_9424,N_7490);
or U11827 (N_11827,N_9672,N_6076);
or U11828 (N_11828,N_8809,N_6685);
nor U11829 (N_11829,N_5020,N_8672);
nor U11830 (N_11830,N_6343,N_5170);
or U11831 (N_11831,N_8725,N_6180);
xor U11832 (N_11832,N_7360,N_6838);
and U11833 (N_11833,N_6365,N_7008);
or U11834 (N_11834,N_5882,N_6397);
and U11835 (N_11835,N_6050,N_7280);
or U11836 (N_11836,N_5914,N_5749);
nand U11837 (N_11837,N_5208,N_5021);
nor U11838 (N_11838,N_9076,N_6807);
nand U11839 (N_11839,N_9915,N_6369);
nand U11840 (N_11840,N_9754,N_6172);
nor U11841 (N_11841,N_5325,N_6432);
nand U11842 (N_11842,N_6119,N_7343);
or U11843 (N_11843,N_6958,N_9831);
and U11844 (N_11844,N_6790,N_9829);
nor U11845 (N_11845,N_9038,N_8538);
and U11846 (N_11846,N_5961,N_5634);
nor U11847 (N_11847,N_5582,N_9285);
nand U11848 (N_11848,N_7611,N_7559);
or U11849 (N_11849,N_8261,N_9372);
or U11850 (N_11850,N_9295,N_9221);
nand U11851 (N_11851,N_7304,N_8496);
or U11852 (N_11852,N_8984,N_6601);
and U11853 (N_11853,N_9087,N_7328);
nor U11854 (N_11854,N_9641,N_5827);
and U11855 (N_11855,N_5212,N_6546);
or U11856 (N_11856,N_8040,N_6184);
nand U11857 (N_11857,N_7191,N_9544);
and U11858 (N_11858,N_9378,N_6281);
and U11859 (N_11859,N_9198,N_6363);
and U11860 (N_11860,N_6082,N_7640);
or U11861 (N_11861,N_6868,N_5692);
or U11862 (N_11862,N_6448,N_9761);
or U11863 (N_11863,N_6218,N_5558);
nand U11864 (N_11864,N_5951,N_9784);
nor U11865 (N_11865,N_5339,N_5251);
nor U11866 (N_11866,N_5744,N_9772);
nor U11867 (N_11867,N_8783,N_7830);
nor U11868 (N_11868,N_6767,N_5955);
or U11869 (N_11869,N_9402,N_7448);
or U11870 (N_11870,N_9913,N_8863);
and U11871 (N_11871,N_5235,N_5527);
nor U11872 (N_11872,N_7467,N_8907);
or U11873 (N_11873,N_7535,N_9721);
xnor U11874 (N_11874,N_6208,N_8921);
nand U11875 (N_11875,N_9505,N_8267);
and U11876 (N_11876,N_9436,N_5780);
nand U11877 (N_11877,N_5222,N_7850);
and U11878 (N_11878,N_7518,N_6147);
or U11879 (N_11879,N_9440,N_8057);
nor U11880 (N_11880,N_5960,N_5252);
nor U11881 (N_11881,N_6384,N_5604);
or U11882 (N_11882,N_5628,N_7439);
or U11883 (N_11883,N_5049,N_7945);
or U11884 (N_11884,N_8854,N_8383);
or U11885 (N_11885,N_7037,N_7890);
nand U11886 (N_11886,N_5367,N_9292);
xnor U11887 (N_11887,N_9562,N_6123);
or U11888 (N_11888,N_9504,N_5141);
and U11889 (N_11889,N_5082,N_8519);
nand U11890 (N_11890,N_6498,N_7013);
and U11891 (N_11891,N_7927,N_9250);
or U11892 (N_11892,N_9495,N_5668);
and U11893 (N_11893,N_6488,N_8466);
or U11894 (N_11894,N_8073,N_7473);
or U11895 (N_11895,N_6251,N_7897);
nand U11896 (N_11896,N_7794,N_7955);
nor U11897 (N_11897,N_9287,N_6588);
nor U11898 (N_11898,N_9456,N_5328);
xor U11899 (N_11899,N_9389,N_5526);
nand U11900 (N_11900,N_6833,N_7540);
or U11901 (N_11901,N_5482,N_9348);
nand U11902 (N_11902,N_5163,N_6540);
or U11903 (N_11903,N_6998,N_6442);
or U11904 (N_11904,N_9723,N_7479);
and U11905 (N_11905,N_9106,N_6978);
xnor U11906 (N_11906,N_9176,N_6525);
or U11907 (N_11907,N_8762,N_9001);
xor U11908 (N_11908,N_9910,N_9094);
nand U11909 (N_11909,N_9042,N_9109);
and U11910 (N_11910,N_5927,N_9319);
and U11911 (N_11911,N_8271,N_9485);
nor U11912 (N_11912,N_7438,N_7129);
nand U11913 (N_11913,N_6274,N_9408);
xnor U11914 (N_11914,N_5489,N_5476);
or U11915 (N_11915,N_6272,N_6908);
or U11916 (N_11916,N_8045,N_7672);
nor U11917 (N_11917,N_5755,N_9461);
or U11918 (N_11918,N_7004,N_7730);
and U11919 (N_11919,N_6292,N_8366);
or U11920 (N_11920,N_9276,N_8858);
and U11921 (N_11921,N_7639,N_5752);
and U11922 (N_11922,N_6464,N_5455);
nand U11923 (N_11923,N_7775,N_9344);
or U11924 (N_11924,N_5405,N_6309);
nand U11925 (N_11925,N_5004,N_5016);
or U11926 (N_11926,N_7437,N_6277);
xor U11927 (N_11927,N_5009,N_5287);
and U11928 (N_11928,N_7001,N_8990);
nand U11929 (N_11929,N_9533,N_6253);
nand U11930 (N_11930,N_8156,N_6095);
and U11931 (N_11931,N_5690,N_9125);
nor U11932 (N_11932,N_5471,N_5085);
nand U11933 (N_11933,N_6793,N_6902);
and U11934 (N_11934,N_5833,N_9791);
nor U11935 (N_11935,N_7627,N_9884);
nor U11936 (N_11936,N_6471,N_9640);
nor U11937 (N_11937,N_7907,N_7675);
nand U11938 (N_11938,N_5046,N_6232);
nand U11939 (N_11939,N_5177,N_8859);
nor U11940 (N_11940,N_8770,N_5813);
nand U11941 (N_11941,N_8484,N_7029);
nor U11942 (N_11942,N_5935,N_7642);
nor U11943 (N_11943,N_6532,N_6919);
or U11944 (N_11944,N_8551,N_7917);
nor U11945 (N_11945,N_6926,N_8499);
or U11946 (N_11946,N_6334,N_7158);
or U11947 (N_11947,N_5128,N_8849);
or U11948 (N_11948,N_5947,N_8274);
or U11949 (N_11949,N_9032,N_9737);
and U11950 (N_11950,N_7309,N_9075);
nand U11951 (N_11951,N_5907,N_9694);
and U11952 (N_11952,N_8355,N_7759);
and U11953 (N_11953,N_8966,N_7087);
nand U11954 (N_11954,N_7606,N_5946);
or U11955 (N_11955,N_9827,N_7977);
and U11956 (N_11956,N_6765,N_7095);
nor U11957 (N_11957,N_8385,N_9851);
nor U11958 (N_11958,N_7843,N_6743);
nand U11959 (N_11959,N_9169,N_7183);
or U11960 (N_11960,N_7505,N_6620);
nor U11961 (N_11961,N_8808,N_8882);
or U11962 (N_11962,N_5306,N_8016);
or U11963 (N_11963,N_6108,N_6377);
or U11964 (N_11964,N_7322,N_6175);
nor U11965 (N_11965,N_5863,N_7374);
or U11966 (N_11966,N_9277,N_8767);
nand U11967 (N_11967,N_6450,N_9064);
nor U11968 (N_11968,N_5679,N_8795);
nand U11969 (N_11969,N_6263,N_6674);
nand U11970 (N_11970,N_8351,N_6565);
xor U11971 (N_11971,N_9666,N_6800);
and U11972 (N_11972,N_5435,N_5821);
or U11973 (N_11973,N_7520,N_6688);
nor U11974 (N_11974,N_7899,N_9620);
or U11975 (N_11975,N_5883,N_8827);
or U11976 (N_11976,N_9621,N_6623);
nor U11977 (N_11977,N_5705,N_6420);
and U11978 (N_11978,N_9229,N_6813);
nand U11979 (N_11979,N_7217,N_7697);
or U11980 (N_11980,N_9543,N_8614);
nor U11981 (N_11981,N_7475,N_5013);
nor U11982 (N_11982,N_8916,N_8836);
or U11983 (N_11983,N_5421,N_5261);
nand U11984 (N_11984,N_8400,N_6462);
nand U11985 (N_11985,N_6562,N_8668);
and U11986 (N_11986,N_7469,N_9016);
and U11987 (N_11987,N_8402,N_7997);
nand U11988 (N_11988,N_8504,N_9535);
or U11989 (N_11989,N_8033,N_8361);
or U11990 (N_11990,N_9609,N_9055);
and U11991 (N_11991,N_5772,N_5324);
nand U11992 (N_11992,N_6898,N_9565);
xor U11993 (N_11993,N_5150,N_8686);
and U11994 (N_11994,N_6999,N_6964);
nand U11995 (N_11995,N_9201,N_6513);
xor U11996 (N_11996,N_9869,N_5239);
and U11997 (N_11997,N_8927,N_6421);
nand U11998 (N_11998,N_8714,N_6504);
nand U11999 (N_11999,N_8742,N_5691);
nor U12000 (N_12000,N_5120,N_5707);
and U12001 (N_12001,N_9972,N_5812);
nor U12002 (N_12002,N_8360,N_5075);
and U12003 (N_12003,N_9303,N_5950);
or U12004 (N_12004,N_5265,N_6748);
nand U12005 (N_12005,N_6247,N_5862);
nand U12006 (N_12006,N_5079,N_6294);
nand U12007 (N_12007,N_7926,N_7704);
and U12008 (N_12008,N_5209,N_8527);
nand U12009 (N_12009,N_9837,N_7692);
and U12010 (N_12010,N_6599,N_8229);
or U12011 (N_12011,N_9668,N_6045);
or U12012 (N_12012,N_6670,N_5030);
nand U12013 (N_12013,N_5687,N_7523);
nand U12014 (N_12014,N_6939,N_8910);
nand U12015 (N_12015,N_5710,N_8800);
or U12016 (N_12016,N_7020,N_9161);
or U12017 (N_12017,N_5699,N_5052);
or U12018 (N_12018,N_5495,N_8816);
nand U12019 (N_12019,N_5876,N_8879);
nand U12020 (N_12020,N_8723,N_8012);
and U12021 (N_12021,N_8494,N_5145);
nand U12022 (N_12022,N_7233,N_7921);
and U12023 (N_12023,N_9005,N_6311);
nand U12024 (N_12024,N_7733,N_6308);
nor U12025 (N_12025,N_9691,N_6225);
nor U12026 (N_12026,N_5103,N_9088);
nand U12027 (N_12027,N_8860,N_9414);
and U12028 (N_12028,N_7503,N_8880);
or U12029 (N_12029,N_8028,N_9437);
and U12030 (N_12030,N_8124,N_7177);
or U12031 (N_12031,N_8290,N_6339);
nand U12032 (N_12032,N_8185,N_5569);
and U12033 (N_12033,N_5868,N_6729);
nor U12034 (N_12034,N_5396,N_8270);
nor U12035 (N_12035,N_9833,N_8438);
nand U12036 (N_12036,N_7866,N_5957);
and U12037 (N_12037,N_7206,N_6547);
nor U12038 (N_12038,N_6948,N_6441);
or U12039 (N_12039,N_6211,N_8570);
nor U12040 (N_12040,N_5383,N_9519);
or U12041 (N_12041,N_6539,N_8624);
nand U12042 (N_12042,N_6335,N_8288);
and U12043 (N_12043,N_9501,N_8251);
nand U12044 (N_12044,N_6407,N_5311);
or U12045 (N_12045,N_9404,N_6677);
nand U12046 (N_12046,N_6901,N_5395);
and U12047 (N_12047,N_9318,N_5903);
and U12048 (N_12048,N_9385,N_9909);
nor U12049 (N_12049,N_5729,N_7656);
nor U12050 (N_12050,N_7677,N_9877);
nor U12051 (N_12051,N_8001,N_8221);
or U12052 (N_12052,N_9006,N_5090);
nor U12053 (N_12053,N_8905,N_9060);
nand U12054 (N_12054,N_8209,N_5063);
nand U12055 (N_12055,N_6600,N_8110);
nand U12056 (N_12056,N_7253,N_9715);
or U12057 (N_12057,N_6458,N_8724);
nor U12058 (N_12058,N_5804,N_9848);
or U12059 (N_12059,N_7382,N_5247);
or U12060 (N_12060,N_9061,N_5199);
nor U12061 (N_12061,N_8801,N_6994);
nor U12062 (N_12062,N_5750,N_6590);
nor U12063 (N_12063,N_7553,N_6219);
nand U12064 (N_12064,N_6788,N_9987);
xor U12065 (N_12065,N_7989,N_6451);
and U12066 (N_12066,N_5878,N_9158);
and U12067 (N_12067,N_9002,N_7149);
and U12068 (N_12068,N_9995,N_8871);
xnor U12069 (N_12069,N_8320,N_8250);
or U12070 (N_12070,N_7622,N_6201);
or U12071 (N_12071,N_9393,N_7506);
nand U12072 (N_12072,N_9679,N_6193);
xnor U12073 (N_12073,N_7822,N_8425);
nand U12074 (N_12074,N_6733,N_8070);
or U12075 (N_12075,N_6989,N_9151);
nor U12076 (N_12076,N_9736,N_6701);
and U12077 (N_12077,N_9227,N_5420);
nor U12078 (N_12078,N_6038,N_7665);
nor U12079 (N_12079,N_9053,N_6861);
and U12080 (N_12080,N_9367,N_8691);
or U12081 (N_12081,N_9843,N_5439);
nor U12082 (N_12082,N_6212,N_8145);
nor U12083 (N_12083,N_8627,N_6481);
or U12084 (N_12084,N_5773,N_7387);
nor U12085 (N_12085,N_5112,N_6755);
nor U12086 (N_12086,N_5297,N_9685);
nand U12087 (N_12087,N_7199,N_5196);
and U12088 (N_12088,N_8900,N_9343);
nor U12089 (N_12089,N_5234,N_5194);
nor U12090 (N_12090,N_7682,N_6700);
and U12091 (N_12091,N_7812,N_7645);
nor U12092 (N_12092,N_8759,N_5776);
nand U12093 (N_12093,N_7761,N_8550);
nand U12094 (N_12094,N_9906,N_6705);
xor U12095 (N_12095,N_6863,N_7398);
nor U12096 (N_12096,N_7774,N_7674);
and U12097 (N_12097,N_9639,N_6260);
nor U12098 (N_12098,N_9750,N_5865);
nand U12099 (N_12099,N_6723,N_7999);
nor U12100 (N_12100,N_7489,N_7154);
nand U12101 (N_12101,N_8365,N_7616);
xnor U12102 (N_12102,N_9105,N_9911);
nor U12103 (N_12103,N_7981,N_8793);
and U12104 (N_12104,N_9165,N_5915);
nand U12105 (N_12105,N_9472,N_9845);
and U12106 (N_12106,N_6732,N_8279);
and U12107 (N_12107,N_6321,N_9730);
nor U12108 (N_12108,N_7270,N_5769);
nand U12109 (N_12109,N_8198,N_5169);
or U12110 (N_12110,N_8571,N_8142);
or U12111 (N_12111,N_5151,N_5379);
nor U12112 (N_12112,N_7227,N_9168);
or U12113 (N_12113,N_8753,N_8852);
and U12114 (N_12114,N_8409,N_8931);
and U12115 (N_12115,N_9110,N_6364);
nor U12116 (N_12116,N_9386,N_6399);
nand U12117 (N_12117,N_7678,N_6092);
or U12118 (N_12118,N_5108,N_7061);
or U12119 (N_12119,N_9534,N_8663);
nor U12120 (N_12120,N_7720,N_8517);
nor U12121 (N_12121,N_5732,N_5932);
xor U12122 (N_12122,N_9454,N_5901);
and U12123 (N_12123,N_9718,N_6961);
nor U12124 (N_12124,N_6900,N_6584);
or U12125 (N_12125,N_5359,N_6273);
nand U12126 (N_12126,N_5683,N_9782);
and U12127 (N_12127,N_6392,N_9116);
or U12128 (N_12128,N_6904,N_5806);
nor U12129 (N_12129,N_8280,N_6004);
nand U12130 (N_12130,N_9033,N_5426);
nand U12131 (N_12131,N_8837,N_6746);
nand U12132 (N_12132,N_7482,N_5361);
nor U12133 (N_12133,N_5469,N_5493);
or U12134 (N_12134,N_9508,N_9124);
or U12135 (N_12135,N_5468,N_8151);
nand U12136 (N_12136,N_9963,N_7221);
or U12137 (N_12137,N_7228,N_5709);
or U12138 (N_12138,N_9828,N_6803);
or U12139 (N_12139,N_7525,N_8416);
nor U12140 (N_12140,N_9510,N_9375);
nand U12141 (N_12141,N_8874,N_8764);
and U12142 (N_12142,N_6234,N_7157);
or U12143 (N_12143,N_7332,N_9358);
and U12144 (N_12144,N_5113,N_8418);
nor U12145 (N_12145,N_7368,N_5360);
and U12146 (N_12146,N_8526,N_7499);
nor U12147 (N_12147,N_5183,N_8689);
nor U12148 (N_12148,N_7935,N_7348);
nor U12149 (N_12149,N_5740,N_8595);
nor U12150 (N_12150,N_6496,N_7002);
and U12151 (N_12151,N_8236,N_7522);
nor U12152 (N_12152,N_9570,N_6427);
or U12153 (N_12153,N_8636,N_6485);
nand U12154 (N_12154,N_7734,N_8055);
nand U12155 (N_12155,N_8765,N_7401);
and U12156 (N_12156,N_9704,N_5296);
nand U12157 (N_12157,N_6280,N_6495);
or U12158 (N_12158,N_9746,N_6975);
nor U12159 (N_12159,N_9297,N_7615);
or U12160 (N_12160,N_5899,N_7313);
and U12161 (N_12161,N_8850,N_7006);
nor U12162 (N_12162,N_7657,N_6602);
or U12163 (N_12163,N_7094,N_9321);
xnor U12164 (N_12164,N_6981,N_8134);
or U12165 (N_12165,N_7101,N_9423);
nand U12166 (N_12166,N_6094,N_7431);
nor U12167 (N_12167,N_9349,N_9997);
xnor U12168 (N_12168,N_7740,N_7043);
nor U12169 (N_12169,N_5519,N_9716);
and U12170 (N_12170,N_7965,N_6158);
or U12171 (N_12171,N_9048,N_7150);
xor U12172 (N_12172,N_6830,N_6973);
nor U12173 (N_12173,N_6489,N_7104);
or U12174 (N_12174,N_7316,N_6773);
nor U12175 (N_12175,N_6144,N_9926);
or U12176 (N_12176,N_6854,N_9466);
nor U12177 (N_12177,N_5700,N_8817);
and U12178 (N_12178,N_6611,N_7234);
nand U12179 (N_12179,N_5696,N_8486);
nand U12180 (N_12180,N_8450,N_8481);
nand U12181 (N_12181,N_6795,N_8129);
nor U12182 (N_12182,N_8508,N_5041);
or U12183 (N_12183,N_5363,N_6316);
xnor U12184 (N_12184,N_9795,N_8752);
nand U12185 (N_12185,N_8737,N_5404);
nand U12186 (N_12186,N_9940,N_5180);
nand U12187 (N_12187,N_6662,N_9463);
and U12188 (N_12188,N_9394,N_5481);
or U12189 (N_12189,N_9890,N_6634);
and U12190 (N_12190,N_7826,N_8069);
nor U12191 (N_12191,N_6897,N_9008);
nor U12192 (N_12192,N_5332,N_9948);
nand U12193 (N_12193,N_7668,N_5716);
nand U12194 (N_12194,N_6224,N_5402);
nor U12195 (N_12195,N_5373,N_8172);
nor U12196 (N_12196,N_6991,N_8511);
nand U12197 (N_12197,N_6669,N_7959);
and U12198 (N_12198,N_8193,N_7062);
or U12199 (N_12199,N_5270,N_9274);
nor U12200 (N_12200,N_6084,N_7592);
or U12201 (N_12201,N_5203,N_7455);
nand U12202 (N_12202,N_9751,N_6740);
and U12203 (N_12203,N_8824,N_7097);
or U12204 (N_12204,N_6093,N_7175);
nor U12205 (N_12205,N_6143,N_6655);
nand U12206 (N_12206,N_6544,N_9422);
and U12207 (N_12207,N_6679,N_6305);
nor U12208 (N_12208,N_9967,N_9633);
and U12209 (N_12209,N_7341,N_8722);
nand U12210 (N_12210,N_6446,N_9653);
nor U12211 (N_12211,N_8043,N_7973);
nor U12212 (N_12212,N_8695,N_7702);
nand U12213 (N_12213,N_8052,N_9659);
and U12214 (N_12214,N_6573,N_7132);
and U12215 (N_12215,N_8242,N_8432);
nor U12216 (N_12216,N_5622,N_9205);
or U12217 (N_12217,N_6589,N_6607);
nor U12218 (N_12218,N_6706,N_6287);
xor U12219 (N_12219,N_8046,N_8249);
xor U12220 (N_12220,N_5249,N_7408);
and U12221 (N_12221,N_5535,N_5637);
nor U12222 (N_12222,N_7968,N_8068);
or U12223 (N_12223,N_8814,N_5647);
and U12224 (N_12224,N_8823,N_8316);
nor U12225 (N_12225,N_9656,N_7116);
nor U12226 (N_12226,N_6858,N_8818);
or U12227 (N_12227,N_6054,N_9727);
nor U12228 (N_12228,N_5043,N_5778);
nand U12229 (N_12229,N_6467,N_8465);
nor U12230 (N_12230,N_5849,N_7779);
or U12231 (N_12231,N_8755,N_5499);
nand U12232 (N_12232,N_7769,N_5602);
or U12233 (N_12233,N_9760,N_9112);
and U12234 (N_12234,N_7950,N_7705);
nor U12235 (N_12235,N_7813,N_8277);
or U12236 (N_12236,N_6030,N_8051);
nor U12237 (N_12237,N_7281,N_7504);
or U12238 (N_12238,N_9518,N_9291);
and U12239 (N_12239,N_7033,N_8302);
and U12240 (N_12240,N_9798,N_8410);
and U12241 (N_12241,N_8339,N_8346);
and U12242 (N_12242,N_6850,N_6582);
nand U12243 (N_12243,N_5263,N_8612);
nor U12244 (N_12244,N_8170,N_8163);
nand U12245 (N_12245,N_9407,N_9316);
and U12246 (N_12246,N_9253,N_8763);
nand U12247 (N_12247,N_6840,N_8530);
and U12248 (N_12248,N_8218,N_7957);
and U12249 (N_12249,N_8510,N_9102);
and U12250 (N_12250,N_6627,N_6661);
and U12251 (N_12251,N_8117,N_6871);
nand U12252 (N_12252,N_9949,N_5977);
or U12253 (N_12253,N_8774,N_9108);
or U12254 (N_12254,N_8294,N_5988);
or U12255 (N_12255,N_9010,N_6477);
and U12256 (N_12256,N_8433,N_6275);
nor U12257 (N_12257,N_5504,N_9532);
and U12258 (N_12258,N_7088,N_9981);
or U12259 (N_12259,N_7925,N_5606);
xor U12260 (N_12260,N_9558,N_9332);
xor U12261 (N_12261,N_6055,N_8732);
nand U12262 (N_12262,N_7216,N_7513);
and U12263 (N_12263,N_5872,N_6728);
nand U12264 (N_12264,N_7707,N_6571);
or U12265 (N_12265,N_8949,N_6002);
or U12266 (N_12266,N_5644,N_6415);
and U12267 (N_12267,N_8044,N_7784);
nor U12268 (N_12268,N_6686,N_5040);
or U12269 (N_12269,N_8395,N_6548);
nand U12270 (N_12270,N_5461,N_5669);
nand U12271 (N_12271,N_5984,N_5178);
nor U12272 (N_12272,N_5072,N_5660);
or U12273 (N_12273,N_9811,N_6434);
and U12274 (N_12274,N_7446,N_6628);
or U12275 (N_12275,N_5722,N_8344);
or U12276 (N_12276,N_9770,N_6352);
nor U12277 (N_12277,N_9883,N_7069);
and U12278 (N_12278,N_9576,N_9844);
nor U12279 (N_12279,N_9569,N_5406);
nand U12280 (N_12280,N_7853,N_7728);
and U12281 (N_12281,N_6683,N_8303);
and U12282 (N_12282,N_9536,N_9418);
and U12283 (N_12283,N_9223,N_6780);
or U12284 (N_12284,N_9516,N_5820);
nand U12285 (N_12285,N_9162,N_7015);
nor U12286 (N_12286,N_9970,N_7255);
or U12287 (N_12287,N_8796,N_7451);
nand U12288 (N_12288,N_8717,N_8918);
and U12289 (N_12289,N_5694,N_8312);
and U12290 (N_12290,N_5017,N_5503);
or U12291 (N_12291,N_5293,N_9145);
nor U12292 (N_12292,N_9334,N_7396);
and U12293 (N_12293,N_9580,N_6405);
and U12294 (N_12294,N_5823,N_5425);
nand U12295 (N_12295,N_7942,N_6491);
or U12296 (N_12296,N_9130,N_5187);
or U12297 (N_12297,N_9975,N_8121);
or U12298 (N_12298,N_6877,N_7119);
or U12299 (N_12299,N_6899,N_6290);
nor U12300 (N_12300,N_8922,N_6846);
nor U12301 (N_12301,N_5708,N_8989);
nand U12302 (N_12302,N_7842,N_6609);
nand U12303 (N_12303,N_9762,N_7354);
or U12304 (N_12304,N_5667,N_6160);
and U12305 (N_12305,N_5681,N_8656);
nor U12306 (N_12306,N_9192,N_7561);
nor U12307 (N_12307,N_8328,N_7910);
nand U12308 (N_12308,N_5742,N_8985);
or U12309 (N_12309,N_8390,N_5522);
and U12310 (N_12310,N_9362,N_9823);
or U12311 (N_12311,N_5580,N_7428);
nand U12312 (N_12312,N_6954,N_5712);
xor U12313 (N_12313,N_7190,N_6483);
and U12314 (N_12314,N_7176,N_8397);
nand U12315 (N_12315,N_7531,N_8423);
and U12316 (N_12316,N_7331,N_9642);
and U12317 (N_12317,N_8286,N_6194);
nor U12318 (N_12318,N_9035,N_6429);
nor U12319 (N_12319,N_9759,N_5152);
nand U12320 (N_12320,N_8003,N_7256);
nor U12321 (N_12321,N_8282,N_9255);
nor U12322 (N_12322,N_5281,N_9618);
and U12323 (N_12323,N_5795,N_6372);
or U12324 (N_12324,N_9240,N_6617);
or U12325 (N_12325,N_5189,N_6368);
and U12326 (N_12326,N_7894,N_6712);
and U12327 (N_12327,N_8941,N_5826);
nand U12328 (N_12328,N_9644,N_9009);
and U12329 (N_12329,N_5089,N_5464);
nand U12330 (N_12330,N_7462,N_9925);
or U12331 (N_12331,N_7012,N_8058);
nand U12332 (N_12332,N_6039,N_5477);
or U12333 (N_12333,N_6735,N_9646);
nor U12334 (N_12334,N_7212,N_9955);
and U12335 (N_12335,N_5343,N_6210);
and U12336 (N_12336,N_8772,N_6020);
nand U12337 (N_12337,N_6269,N_6098);
nand U12338 (N_12338,N_5327,N_8579);
xor U12339 (N_12339,N_8235,N_9226);
nand U12340 (N_12340,N_6461,N_8514);
and U12341 (N_12341,N_6278,N_5635);
or U12342 (N_12342,N_7114,N_7783);
and U12343 (N_12343,N_5276,N_6069);
nand U12344 (N_12344,N_6905,N_6736);
nand U12345 (N_12345,N_5990,N_7363);
and U12346 (N_12346,N_6714,N_7107);
and U12347 (N_12347,N_6913,N_9080);
nor U12348 (N_12348,N_6189,N_9317);
or U12349 (N_12349,N_8208,N_8338);
nand U12350 (N_12350,N_8313,N_8427);
nand U12351 (N_12351,N_9400,N_5507);
nand U12352 (N_12352,N_7019,N_9403);
or U12353 (N_12353,N_6236,N_6935);
xnor U12354 (N_12354,N_5638,N_5945);
nand U12355 (N_12355,N_9157,N_7044);
nor U12356 (N_12356,N_8894,N_7984);
and U12357 (N_12357,N_6070,N_7405);
or U12358 (N_12358,N_6635,N_8618);
or U12359 (N_12359,N_5099,N_7031);
and U12360 (N_12360,N_8143,N_8928);
and U12361 (N_12361,N_9627,N_5033);
nand U12362 (N_12362,N_9605,N_8613);
or U12363 (N_12363,N_7510,N_6022);
or U12364 (N_12364,N_7342,N_6764);
nor U12365 (N_12365,N_8590,N_7125);
or U12366 (N_12366,N_8457,N_6396);
and U12367 (N_12367,N_9072,N_6431);
and U12368 (N_12368,N_5101,N_7299);
or U12369 (N_12369,N_7394,N_9262);
nor U12370 (N_12370,N_5071,N_5483);
or U12371 (N_12371,N_6993,N_5924);
nor U12372 (N_12372,N_6751,N_7289);
and U12373 (N_12373,N_5156,N_6240);
nand U12374 (N_12374,N_8975,N_5808);
and U12375 (N_12375,N_7618,N_8719);
or U12376 (N_12376,N_6293,N_8114);
nor U12377 (N_12377,N_8963,N_9863);
nand U12378 (N_12378,N_7944,N_7189);
nor U12379 (N_12379,N_6690,N_6391);
nand U12380 (N_12380,N_7351,N_5557);
or U12381 (N_12381,N_9296,N_8754);
nand U12382 (N_12382,N_9614,N_7806);
and U12383 (N_12383,N_8980,N_7751);
and U12384 (N_12384,N_8389,N_9796);
and U12385 (N_12385,N_8258,N_5875);
and U12386 (N_12386,N_6016,N_9479);
nand U12387 (N_12387,N_9748,N_7174);
nor U12388 (N_12388,N_8601,N_6622);
nor U12389 (N_12389,N_7936,N_8375);
nor U12390 (N_12390,N_5871,N_8734);
nor U12391 (N_12391,N_9810,N_8690);
xor U12392 (N_12392,N_9310,N_9567);
and U12393 (N_12393,N_5340,N_7340);
and U12394 (N_12394,N_9593,N_7841);
xor U12395 (N_12395,N_6716,N_6882);
and U12396 (N_12396,N_7153,N_5066);
and U12397 (N_12397,N_5254,N_7594);
or U12398 (N_12398,N_9705,N_6186);
nor U12399 (N_12399,N_8173,N_9971);
nand U12400 (N_12400,N_7134,N_5123);
nor U12401 (N_12401,N_6884,N_8315);
nor U12402 (N_12402,N_5224,N_9912);
or U12403 (N_12403,N_7296,N_8782);
and U12404 (N_12404,N_9801,N_8109);
or U12405 (N_12405,N_8471,N_6766);
or U12406 (N_12406,N_8518,N_8676);
nor U12407 (N_12407,N_8169,N_7042);
or U12408 (N_12408,N_5215,N_6557);
nor U12409 (N_12409,N_6469,N_7828);
nor U12410 (N_12410,N_6953,N_9860);
and U12411 (N_12411,N_8087,N_5182);
and U12412 (N_12412,N_6102,N_5342);
nand U12413 (N_12413,N_8421,N_8887);
or U12414 (N_12414,N_7845,N_7293);
nand U12415 (N_12415,N_6254,N_7246);
or U12416 (N_12416,N_9624,N_5999);
or U12417 (N_12417,N_7297,N_6181);
and U12418 (N_12418,N_9246,N_6357);
or U12419 (N_12419,N_7802,N_6879);
nor U12420 (N_12420,N_8914,N_8662);
nor U12421 (N_12421,N_9651,N_8996);
nand U12422 (N_12422,N_7931,N_5318);
nand U12423 (N_12423,N_7923,N_6713);
and U12424 (N_12424,N_9020,N_7099);
and U12425 (N_12425,N_9947,N_6689);
and U12426 (N_12426,N_5416,N_7661);
xnor U12427 (N_12427,N_7118,N_9560);
and U12428 (N_12428,N_8182,N_9057);
or U12429 (N_12429,N_7005,N_9433);
or U12430 (N_12430,N_5848,N_7445);
nor U12431 (N_12431,N_6375,N_8083);
and U12432 (N_12432,N_7425,N_9647);
and U12433 (N_12433,N_7223,N_7726);
nand U12434 (N_12434,N_5759,N_6719);
nor U12435 (N_12435,N_9990,N_7715);
or U12436 (N_12436,N_7170,N_9528);
and U12437 (N_12437,N_7796,N_7155);
or U12438 (N_12438,N_9555,N_5684);
and U12439 (N_12439,N_5107,N_7886);
or U12440 (N_12440,N_7493,N_6026);
nor U12441 (N_12441,N_7435,N_8233);
nor U12442 (N_12442,N_9688,N_8660);
or U12443 (N_12443,N_9985,N_6581);
nor U12444 (N_12444,N_8994,N_9541);
nor U12445 (N_12445,N_8842,N_8777);
and U12446 (N_12446,N_6768,N_7593);
nand U12447 (N_12447,N_9966,N_8904);
or U12448 (N_12448,N_8082,N_8731);
nand U12449 (N_12449,N_9854,N_5979);
nand U12450 (N_12450,N_5377,N_8483);
or U12451 (N_12451,N_8643,N_9671);
nand U12452 (N_12452,N_9235,N_6744);
or U12453 (N_12453,N_8195,N_5124);
and U12454 (N_12454,N_9839,N_8059);
or U12455 (N_12455,N_9665,N_6103);
and U12456 (N_12456,N_9457,N_9455);
nand U12457 (N_12457,N_5860,N_6032);
and U12458 (N_12458,N_5553,N_9551);
and U12459 (N_12459,N_5819,N_6255);
and U12460 (N_12460,N_8444,N_6878);
and U12461 (N_12461,N_6715,N_7205);
and U12462 (N_12462,N_7971,N_5555);
or U12463 (N_12463,N_5551,N_9584);
and U12464 (N_12464,N_5313,N_6191);
and U12465 (N_12465,N_8840,N_5310);
or U12466 (N_12466,N_8485,N_5540);
or U12467 (N_12467,N_7441,N_9435);
xnor U12468 (N_12468,N_8401,N_6304);
and U12469 (N_12469,N_5818,N_9352);
and U12470 (N_12470,N_6664,N_8398);
nor U12471 (N_12471,N_6567,N_8374);
or U12472 (N_12472,N_7392,N_5486);
or U12473 (N_12473,N_8804,N_5919);
and U12474 (N_12474,N_5936,N_7554);
nor U12475 (N_12475,N_8297,N_6753);
nor U12476 (N_12476,N_8593,N_9864);
nand U12477 (N_12477,N_5146,N_6996);
nand U12478 (N_12478,N_6577,N_9634);
or U12479 (N_12479,N_9051,N_5473);
nor U12480 (N_12480,N_7911,N_7201);
xnor U12481 (N_12481,N_8756,N_7254);
nand U12482 (N_12482,N_8626,N_9468);
or U12483 (N_12483,N_8707,N_9180);
nor U12484 (N_12484,N_9638,N_6832);
nor U12485 (N_12485,N_8004,N_7543);
xnor U12486 (N_12486,N_8256,N_8147);
nand U12487 (N_12487,N_5641,N_9047);
nor U12488 (N_12488,N_8891,N_8712);
or U12489 (N_12489,N_8740,N_5300);
nand U12490 (N_12490,N_7744,N_7573);
or U12491 (N_12491,N_9359,N_7609);
or U12492 (N_12492,N_7147,N_9428);
nand U12493 (N_12493,N_6284,N_6509);
nand U12494 (N_12494,N_5451,N_7023);
or U12495 (N_12495,N_9946,N_9582);
nand U12496 (N_12496,N_9767,N_9619);
nand U12497 (N_12497,N_5583,N_7141);
nand U12498 (N_12498,N_9135,N_6801);
or U12499 (N_12499,N_7386,N_7631);
nor U12500 (N_12500,N_6375,N_9325);
nand U12501 (N_12501,N_8595,N_8804);
nor U12502 (N_12502,N_5624,N_5667);
nor U12503 (N_12503,N_8815,N_6098);
nand U12504 (N_12504,N_5381,N_7721);
or U12505 (N_12505,N_8053,N_7521);
nand U12506 (N_12506,N_7843,N_7963);
nor U12507 (N_12507,N_7928,N_7900);
nand U12508 (N_12508,N_6895,N_5443);
nand U12509 (N_12509,N_6614,N_9726);
nand U12510 (N_12510,N_5650,N_5955);
nor U12511 (N_12511,N_8872,N_7392);
and U12512 (N_12512,N_8871,N_5013);
or U12513 (N_12513,N_7101,N_8599);
nand U12514 (N_12514,N_7810,N_6084);
or U12515 (N_12515,N_9383,N_7313);
and U12516 (N_12516,N_7167,N_6366);
nand U12517 (N_12517,N_8858,N_7039);
nand U12518 (N_12518,N_7019,N_5982);
nor U12519 (N_12519,N_5336,N_8415);
nor U12520 (N_12520,N_5546,N_6301);
or U12521 (N_12521,N_9828,N_6107);
nand U12522 (N_12522,N_8339,N_9995);
nor U12523 (N_12523,N_6878,N_9172);
or U12524 (N_12524,N_5570,N_5299);
nand U12525 (N_12525,N_6038,N_5181);
nand U12526 (N_12526,N_5735,N_7836);
and U12527 (N_12527,N_9345,N_7191);
nor U12528 (N_12528,N_5025,N_7133);
or U12529 (N_12529,N_7795,N_7475);
and U12530 (N_12530,N_9963,N_8823);
or U12531 (N_12531,N_8181,N_5764);
xnor U12532 (N_12532,N_7753,N_6964);
nand U12533 (N_12533,N_5721,N_9804);
nand U12534 (N_12534,N_7160,N_7667);
nand U12535 (N_12535,N_5701,N_8404);
nor U12536 (N_12536,N_7756,N_5103);
or U12537 (N_12537,N_9027,N_8162);
xor U12538 (N_12538,N_6361,N_5812);
and U12539 (N_12539,N_8155,N_7484);
and U12540 (N_12540,N_7850,N_5373);
nor U12541 (N_12541,N_5522,N_9020);
nor U12542 (N_12542,N_6064,N_6249);
nand U12543 (N_12543,N_6949,N_7027);
or U12544 (N_12544,N_8306,N_6642);
and U12545 (N_12545,N_6553,N_9512);
nand U12546 (N_12546,N_6493,N_7774);
or U12547 (N_12547,N_6861,N_6364);
or U12548 (N_12548,N_8163,N_6060);
nand U12549 (N_12549,N_8321,N_9190);
nor U12550 (N_12550,N_8362,N_7836);
nand U12551 (N_12551,N_9937,N_9723);
and U12552 (N_12552,N_9183,N_7651);
or U12553 (N_12553,N_9141,N_7440);
and U12554 (N_12554,N_6245,N_6058);
or U12555 (N_12555,N_7422,N_6212);
nor U12556 (N_12556,N_7835,N_9706);
and U12557 (N_12557,N_5243,N_6996);
and U12558 (N_12558,N_8784,N_5650);
or U12559 (N_12559,N_9854,N_7907);
or U12560 (N_12560,N_5501,N_5159);
and U12561 (N_12561,N_8806,N_9739);
nor U12562 (N_12562,N_5278,N_5969);
nor U12563 (N_12563,N_9037,N_9556);
or U12564 (N_12564,N_6613,N_5989);
and U12565 (N_12565,N_7148,N_7715);
or U12566 (N_12566,N_6028,N_7744);
or U12567 (N_12567,N_7850,N_6093);
and U12568 (N_12568,N_9337,N_5660);
and U12569 (N_12569,N_5559,N_5270);
or U12570 (N_12570,N_6812,N_6864);
nor U12571 (N_12571,N_7998,N_9740);
nor U12572 (N_12572,N_6245,N_5480);
nand U12573 (N_12573,N_9508,N_9226);
and U12574 (N_12574,N_6230,N_6842);
nand U12575 (N_12575,N_5111,N_6846);
and U12576 (N_12576,N_7324,N_8365);
nand U12577 (N_12577,N_5782,N_7474);
nand U12578 (N_12578,N_6371,N_6939);
nand U12579 (N_12579,N_9011,N_6545);
and U12580 (N_12580,N_9877,N_9929);
nand U12581 (N_12581,N_8462,N_5097);
nor U12582 (N_12582,N_7640,N_9680);
and U12583 (N_12583,N_8211,N_8941);
or U12584 (N_12584,N_8793,N_7506);
nor U12585 (N_12585,N_8263,N_7168);
nor U12586 (N_12586,N_5657,N_5556);
or U12587 (N_12587,N_6340,N_6543);
or U12588 (N_12588,N_5082,N_6700);
nand U12589 (N_12589,N_9339,N_8934);
or U12590 (N_12590,N_9202,N_5618);
and U12591 (N_12591,N_9862,N_6900);
and U12592 (N_12592,N_7010,N_5667);
and U12593 (N_12593,N_8628,N_5238);
nand U12594 (N_12594,N_5176,N_6506);
nand U12595 (N_12595,N_6718,N_7864);
or U12596 (N_12596,N_8351,N_6405);
or U12597 (N_12597,N_6273,N_6076);
or U12598 (N_12598,N_6032,N_9238);
nand U12599 (N_12599,N_9840,N_9684);
and U12600 (N_12600,N_7204,N_8363);
or U12601 (N_12601,N_9684,N_5489);
or U12602 (N_12602,N_5898,N_7822);
and U12603 (N_12603,N_7848,N_7043);
nor U12604 (N_12604,N_8148,N_9006);
or U12605 (N_12605,N_9447,N_7683);
or U12606 (N_12606,N_7709,N_8820);
nand U12607 (N_12607,N_8397,N_7331);
nand U12608 (N_12608,N_9537,N_6805);
and U12609 (N_12609,N_7489,N_8890);
xor U12610 (N_12610,N_8143,N_5821);
or U12611 (N_12611,N_6039,N_5491);
and U12612 (N_12612,N_9789,N_7035);
or U12613 (N_12613,N_7675,N_8533);
nor U12614 (N_12614,N_8182,N_8050);
and U12615 (N_12615,N_5017,N_9707);
xnor U12616 (N_12616,N_7376,N_8506);
or U12617 (N_12617,N_5601,N_9353);
or U12618 (N_12618,N_8143,N_6734);
nor U12619 (N_12619,N_9451,N_5531);
nor U12620 (N_12620,N_6959,N_8734);
nand U12621 (N_12621,N_5217,N_8747);
nor U12622 (N_12622,N_9268,N_9695);
nor U12623 (N_12623,N_6192,N_8403);
or U12624 (N_12624,N_7663,N_7624);
nor U12625 (N_12625,N_8108,N_8019);
and U12626 (N_12626,N_9708,N_7348);
nand U12627 (N_12627,N_8495,N_8200);
and U12628 (N_12628,N_6941,N_6274);
and U12629 (N_12629,N_9039,N_9542);
nor U12630 (N_12630,N_5047,N_7801);
nand U12631 (N_12631,N_8302,N_8644);
and U12632 (N_12632,N_7539,N_9365);
nor U12633 (N_12633,N_7346,N_7861);
nor U12634 (N_12634,N_6910,N_8806);
nor U12635 (N_12635,N_7312,N_5711);
nor U12636 (N_12636,N_8407,N_5281);
and U12637 (N_12637,N_9428,N_8233);
nor U12638 (N_12638,N_7113,N_8423);
or U12639 (N_12639,N_8307,N_5928);
or U12640 (N_12640,N_9540,N_7562);
and U12641 (N_12641,N_7497,N_5491);
and U12642 (N_12642,N_8918,N_6479);
nor U12643 (N_12643,N_7228,N_6051);
or U12644 (N_12644,N_7839,N_9384);
and U12645 (N_12645,N_9401,N_8324);
nor U12646 (N_12646,N_7321,N_5396);
and U12647 (N_12647,N_5696,N_9237);
nand U12648 (N_12648,N_6911,N_9549);
and U12649 (N_12649,N_5129,N_5012);
xnor U12650 (N_12650,N_8394,N_8439);
and U12651 (N_12651,N_5530,N_8669);
nor U12652 (N_12652,N_8852,N_5102);
and U12653 (N_12653,N_7624,N_7263);
and U12654 (N_12654,N_9992,N_8834);
and U12655 (N_12655,N_8341,N_9385);
nand U12656 (N_12656,N_6474,N_6455);
nand U12657 (N_12657,N_5015,N_9742);
nor U12658 (N_12658,N_8829,N_7701);
or U12659 (N_12659,N_7174,N_9832);
and U12660 (N_12660,N_6021,N_5983);
nand U12661 (N_12661,N_8882,N_7644);
or U12662 (N_12662,N_5089,N_6179);
or U12663 (N_12663,N_7011,N_5639);
or U12664 (N_12664,N_9368,N_7773);
nor U12665 (N_12665,N_5457,N_5965);
or U12666 (N_12666,N_7033,N_7660);
and U12667 (N_12667,N_6345,N_7001);
nor U12668 (N_12668,N_9337,N_9152);
nand U12669 (N_12669,N_8728,N_5546);
nor U12670 (N_12670,N_6814,N_9826);
or U12671 (N_12671,N_6266,N_9090);
nand U12672 (N_12672,N_6812,N_5933);
and U12673 (N_12673,N_5645,N_5879);
and U12674 (N_12674,N_7891,N_9567);
and U12675 (N_12675,N_5454,N_8715);
and U12676 (N_12676,N_7265,N_5943);
and U12677 (N_12677,N_7193,N_8545);
nor U12678 (N_12678,N_6896,N_7798);
nand U12679 (N_12679,N_5535,N_9811);
nor U12680 (N_12680,N_9680,N_9135);
and U12681 (N_12681,N_6510,N_5327);
nand U12682 (N_12682,N_8976,N_7922);
or U12683 (N_12683,N_7278,N_9592);
nand U12684 (N_12684,N_8845,N_9552);
nor U12685 (N_12685,N_5895,N_6766);
and U12686 (N_12686,N_7460,N_6452);
nor U12687 (N_12687,N_5809,N_7940);
and U12688 (N_12688,N_9563,N_9843);
nand U12689 (N_12689,N_5796,N_7872);
xnor U12690 (N_12690,N_6391,N_8235);
or U12691 (N_12691,N_5182,N_8309);
nor U12692 (N_12692,N_5895,N_6572);
nand U12693 (N_12693,N_6864,N_8498);
nand U12694 (N_12694,N_6152,N_9679);
or U12695 (N_12695,N_7879,N_5092);
nor U12696 (N_12696,N_6399,N_7379);
and U12697 (N_12697,N_8961,N_9417);
nand U12698 (N_12698,N_5816,N_9136);
or U12699 (N_12699,N_7157,N_9588);
and U12700 (N_12700,N_6553,N_6789);
or U12701 (N_12701,N_7499,N_9671);
or U12702 (N_12702,N_9786,N_7984);
nor U12703 (N_12703,N_7668,N_6477);
nand U12704 (N_12704,N_5246,N_8172);
xor U12705 (N_12705,N_9915,N_6997);
xor U12706 (N_12706,N_5289,N_5370);
nand U12707 (N_12707,N_7352,N_5766);
or U12708 (N_12708,N_8006,N_9216);
nor U12709 (N_12709,N_6384,N_8086);
or U12710 (N_12710,N_8498,N_6042);
and U12711 (N_12711,N_5314,N_7980);
nor U12712 (N_12712,N_8366,N_9210);
and U12713 (N_12713,N_6802,N_7876);
nor U12714 (N_12714,N_8327,N_9717);
nor U12715 (N_12715,N_5048,N_6232);
and U12716 (N_12716,N_6603,N_7053);
nor U12717 (N_12717,N_8762,N_7924);
or U12718 (N_12718,N_5946,N_5587);
nand U12719 (N_12719,N_9568,N_8697);
nand U12720 (N_12720,N_7273,N_6435);
and U12721 (N_12721,N_7811,N_6873);
or U12722 (N_12722,N_7308,N_8684);
nor U12723 (N_12723,N_8257,N_6063);
nand U12724 (N_12724,N_5321,N_5931);
nand U12725 (N_12725,N_9847,N_8548);
or U12726 (N_12726,N_7781,N_9754);
or U12727 (N_12727,N_9685,N_9422);
nor U12728 (N_12728,N_5785,N_8760);
and U12729 (N_12729,N_9331,N_8241);
or U12730 (N_12730,N_8037,N_6786);
nand U12731 (N_12731,N_8229,N_9273);
or U12732 (N_12732,N_8717,N_9651);
and U12733 (N_12733,N_5069,N_8114);
and U12734 (N_12734,N_8748,N_7703);
nor U12735 (N_12735,N_5058,N_7175);
or U12736 (N_12736,N_8933,N_9717);
or U12737 (N_12737,N_8406,N_9850);
nor U12738 (N_12738,N_8740,N_8871);
and U12739 (N_12739,N_5045,N_6903);
or U12740 (N_12740,N_9482,N_7545);
or U12741 (N_12741,N_5273,N_7181);
and U12742 (N_12742,N_5898,N_6852);
and U12743 (N_12743,N_7673,N_5606);
nand U12744 (N_12744,N_5301,N_5504);
nor U12745 (N_12745,N_5017,N_9290);
and U12746 (N_12746,N_8999,N_7704);
nand U12747 (N_12747,N_8770,N_6204);
and U12748 (N_12748,N_6558,N_5470);
and U12749 (N_12749,N_7565,N_6055);
nor U12750 (N_12750,N_5400,N_9286);
nand U12751 (N_12751,N_7484,N_9023);
or U12752 (N_12752,N_8499,N_6798);
or U12753 (N_12753,N_9416,N_8382);
and U12754 (N_12754,N_5595,N_5223);
nor U12755 (N_12755,N_8513,N_8142);
or U12756 (N_12756,N_7359,N_8652);
or U12757 (N_12757,N_6745,N_9889);
and U12758 (N_12758,N_7808,N_8410);
and U12759 (N_12759,N_8728,N_5995);
and U12760 (N_12760,N_5759,N_9420);
nor U12761 (N_12761,N_6092,N_7928);
or U12762 (N_12762,N_5445,N_5777);
and U12763 (N_12763,N_7115,N_9660);
nand U12764 (N_12764,N_7963,N_8372);
and U12765 (N_12765,N_9981,N_7369);
or U12766 (N_12766,N_5339,N_5568);
xnor U12767 (N_12767,N_9727,N_7600);
nor U12768 (N_12768,N_7673,N_7858);
and U12769 (N_12769,N_7862,N_8697);
nor U12770 (N_12770,N_8565,N_5240);
and U12771 (N_12771,N_5646,N_7965);
and U12772 (N_12772,N_9351,N_7715);
nand U12773 (N_12773,N_7592,N_7952);
nor U12774 (N_12774,N_5793,N_7444);
and U12775 (N_12775,N_7461,N_8201);
and U12776 (N_12776,N_6107,N_5402);
or U12777 (N_12777,N_5724,N_7226);
nand U12778 (N_12778,N_5222,N_8790);
nor U12779 (N_12779,N_6137,N_5877);
or U12780 (N_12780,N_6463,N_6748);
and U12781 (N_12781,N_9909,N_6440);
and U12782 (N_12782,N_8871,N_5115);
and U12783 (N_12783,N_9305,N_5821);
and U12784 (N_12784,N_7499,N_9916);
nand U12785 (N_12785,N_5028,N_9143);
nor U12786 (N_12786,N_7318,N_9402);
or U12787 (N_12787,N_7240,N_5763);
nor U12788 (N_12788,N_7704,N_5434);
and U12789 (N_12789,N_8848,N_5024);
nand U12790 (N_12790,N_8866,N_7418);
or U12791 (N_12791,N_8576,N_8136);
nand U12792 (N_12792,N_5550,N_6056);
nand U12793 (N_12793,N_8415,N_9240);
and U12794 (N_12794,N_7436,N_9904);
nand U12795 (N_12795,N_7425,N_6586);
nand U12796 (N_12796,N_9181,N_9959);
and U12797 (N_12797,N_8024,N_6160);
nor U12798 (N_12798,N_8626,N_8047);
or U12799 (N_12799,N_8848,N_8414);
or U12800 (N_12800,N_8063,N_9552);
and U12801 (N_12801,N_8353,N_8676);
or U12802 (N_12802,N_5778,N_6498);
and U12803 (N_12803,N_9770,N_6780);
or U12804 (N_12804,N_8738,N_6895);
or U12805 (N_12805,N_9490,N_7984);
nand U12806 (N_12806,N_9274,N_8915);
and U12807 (N_12807,N_5849,N_6118);
nor U12808 (N_12808,N_6832,N_6044);
and U12809 (N_12809,N_5628,N_5026);
nand U12810 (N_12810,N_5233,N_7655);
or U12811 (N_12811,N_8673,N_8934);
or U12812 (N_12812,N_8058,N_6034);
or U12813 (N_12813,N_9350,N_5641);
and U12814 (N_12814,N_5154,N_5792);
or U12815 (N_12815,N_9109,N_8118);
and U12816 (N_12816,N_9454,N_7803);
nor U12817 (N_12817,N_8136,N_8311);
and U12818 (N_12818,N_9150,N_7882);
or U12819 (N_12819,N_5304,N_6560);
or U12820 (N_12820,N_8578,N_5286);
and U12821 (N_12821,N_8547,N_6793);
nor U12822 (N_12822,N_7422,N_6174);
or U12823 (N_12823,N_9524,N_8762);
or U12824 (N_12824,N_5861,N_5325);
or U12825 (N_12825,N_8379,N_6049);
and U12826 (N_12826,N_6998,N_6382);
and U12827 (N_12827,N_8459,N_5993);
nor U12828 (N_12828,N_9385,N_9531);
nor U12829 (N_12829,N_9014,N_8031);
nand U12830 (N_12830,N_6928,N_8026);
nand U12831 (N_12831,N_6539,N_6538);
and U12832 (N_12832,N_7898,N_7022);
nand U12833 (N_12833,N_6079,N_5588);
and U12834 (N_12834,N_8124,N_6698);
and U12835 (N_12835,N_7303,N_9703);
nor U12836 (N_12836,N_9555,N_7531);
xnor U12837 (N_12837,N_7267,N_7889);
nor U12838 (N_12838,N_6832,N_5898);
nand U12839 (N_12839,N_5886,N_7550);
nor U12840 (N_12840,N_6119,N_7968);
or U12841 (N_12841,N_9159,N_6325);
and U12842 (N_12842,N_6040,N_7150);
nor U12843 (N_12843,N_6624,N_6947);
xnor U12844 (N_12844,N_5610,N_6597);
xor U12845 (N_12845,N_9121,N_7503);
or U12846 (N_12846,N_7328,N_5780);
nand U12847 (N_12847,N_9534,N_6016);
and U12848 (N_12848,N_9723,N_5645);
xor U12849 (N_12849,N_5816,N_8430);
or U12850 (N_12850,N_9534,N_6272);
nor U12851 (N_12851,N_5288,N_5850);
nor U12852 (N_12852,N_8367,N_8481);
nor U12853 (N_12853,N_5274,N_8890);
and U12854 (N_12854,N_9977,N_8796);
nor U12855 (N_12855,N_5732,N_6930);
nor U12856 (N_12856,N_6249,N_6354);
and U12857 (N_12857,N_6277,N_8000);
and U12858 (N_12858,N_9101,N_8177);
or U12859 (N_12859,N_5428,N_9841);
and U12860 (N_12860,N_8204,N_9619);
nor U12861 (N_12861,N_9858,N_8092);
nor U12862 (N_12862,N_6720,N_7350);
xor U12863 (N_12863,N_6736,N_7147);
or U12864 (N_12864,N_6353,N_9689);
or U12865 (N_12865,N_7557,N_9072);
nand U12866 (N_12866,N_7038,N_9462);
or U12867 (N_12867,N_5626,N_5039);
and U12868 (N_12868,N_5706,N_5377);
or U12869 (N_12869,N_7513,N_7151);
and U12870 (N_12870,N_8857,N_7645);
nand U12871 (N_12871,N_9126,N_9384);
or U12872 (N_12872,N_5737,N_9444);
nand U12873 (N_12873,N_5275,N_8752);
nand U12874 (N_12874,N_8912,N_8117);
nor U12875 (N_12875,N_8099,N_6626);
and U12876 (N_12876,N_8643,N_7841);
or U12877 (N_12877,N_7893,N_8582);
nand U12878 (N_12878,N_6025,N_6873);
nand U12879 (N_12879,N_7713,N_9397);
nor U12880 (N_12880,N_8122,N_5829);
nand U12881 (N_12881,N_5804,N_7410);
nor U12882 (N_12882,N_6402,N_5221);
nand U12883 (N_12883,N_5707,N_6621);
and U12884 (N_12884,N_6768,N_5024);
and U12885 (N_12885,N_6360,N_8205);
nand U12886 (N_12886,N_5434,N_7638);
or U12887 (N_12887,N_7547,N_7882);
and U12888 (N_12888,N_9756,N_8156);
and U12889 (N_12889,N_9599,N_9308);
and U12890 (N_12890,N_6258,N_5126);
or U12891 (N_12891,N_9399,N_9659);
nor U12892 (N_12892,N_6231,N_5250);
nor U12893 (N_12893,N_6093,N_8829);
and U12894 (N_12894,N_9293,N_8165);
or U12895 (N_12895,N_7539,N_7478);
nand U12896 (N_12896,N_8500,N_5666);
nand U12897 (N_12897,N_8367,N_5998);
or U12898 (N_12898,N_8252,N_9890);
nor U12899 (N_12899,N_5764,N_8336);
xor U12900 (N_12900,N_5882,N_6722);
and U12901 (N_12901,N_5901,N_9746);
or U12902 (N_12902,N_6125,N_7389);
or U12903 (N_12903,N_9144,N_7414);
nor U12904 (N_12904,N_5803,N_7029);
nor U12905 (N_12905,N_6263,N_7375);
nand U12906 (N_12906,N_9326,N_5595);
and U12907 (N_12907,N_7003,N_9608);
nor U12908 (N_12908,N_8718,N_9637);
and U12909 (N_12909,N_5154,N_8342);
nor U12910 (N_12910,N_5564,N_9931);
or U12911 (N_12911,N_9810,N_8816);
and U12912 (N_12912,N_6484,N_9476);
nor U12913 (N_12913,N_6508,N_5594);
nand U12914 (N_12914,N_7259,N_6643);
or U12915 (N_12915,N_8987,N_8535);
nor U12916 (N_12916,N_5195,N_6431);
nor U12917 (N_12917,N_7693,N_9668);
or U12918 (N_12918,N_9179,N_9683);
and U12919 (N_12919,N_7692,N_6288);
nand U12920 (N_12920,N_6348,N_9518);
nand U12921 (N_12921,N_9008,N_8181);
and U12922 (N_12922,N_8983,N_8709);
or U12923 (N_12923,N_6104,N_7417);
nor U12924 (N_12924,N_8545,N_9225);
nand U12925 (N_12925,N_6973,N_5729);
or U12926 (N_12926,N_6719,N_9884);
and U12927 (N_12927,N_6861,N_9561);
and U12928 (N_12928,N_5310,N_7806);
nor U12929 (N_12929,N_9986,N_5872);
and U12930 (N_12930,N_9847,N_5981);
and U12931 (N_12931,N_7480,N_8121);
nand U12932 (N_12932,N_6988,N_9850);
nor U12933 (N_12933,N_9000,N_5004);
and U12934 (N_12934,N_9613,N_7526);
or U12935 (N_12935,N_5569,N_8269);
nand U12936 (N_12936,N_8702,N_8476);
or U12937 (N_12937,N_8840,N_8465);
nor U12938 (N_12938,N_8955,N_9705);
or U12939 (N_12939,N_8668,N_8141);
or U12940 (N_12940,N_8567,N_8728);
nor U12941 (N_12941,N_6963,N_7042);
or U12942 (N_12942,N_6668,N_9596);
and U12943 (N_12943,N_7305,N_5976);
or U12944 (N_12944,N_6062,N_8433);
nor U12945 (N_12945,N_9624,N_9993);
and U12946 (N_12946,N_8600,N_9636);
or U12947 (N_12947,N_8922,N_5685);
nand U12948 (N_12948,N_8553,N_8305);
nor U12949 (N_12949,N_8118,N_8327);
nor U12950 (N_12950,N_8649,N_8223);
nand U12951 (N_12951,N_9389,N_5750);
and U12952 (N_12952,N_8552,N_9924);
or U12953 (N_12953,N_5643,N_5813);
nand U12954 (N_12954,N_8801,N_5450);
nor U12955 (N_12955,N_9094,N_7170);
nand U12956 (N_12956,N_7840,N_6839);
nor U12957 (N_12957,N_7276,N_5115);
nand U12958 (N_12958,N_7785,N_5611);
and U12959 (N_12959,N_7938,N_9754);
xor U12960 (N_12960,N_9732,N_5273);
nand U12961 (N_12961,N_6962,N_8270);
nand U12962 (N_12962,N_9787,N_9395);
xor U12963 (N_12963,N_8533,N_6458);
nand U12964 (N_12964,N_7883,N_8594);
xnor U12965 (N_12965,N_9311,N_8342);
or U12966 (N_12966,N_7775,N_9400);
nor U12967 (N_12967,N_7119,N_9603);
nand U12968 (N_12968,N_6699,N_6787);
or U12969 (N_12969,N_5324,N_6503);
xor U12970 (N_12970,N_5262,N_7126);
nor U12971 (N_12971,N_9748,N_7055);
nor U12972 (N_12972,N_7466,N_9381);
nand U12973 (N_12973,N_6500,N_6647);
nand U12974 (N_12974,N_7642,N_8770);
and U12975 (N_12975,N_9541,N_8937);
nor U12976 (N_12976,N_6515,N_6296);
xor U12977 (N_12977,N_5689,N_7981);
nand U12978 (N_12978,N_6577,N_6138);
nand U12979 (N_12979,N_7870,N_6300);
and U12980 (N_12980,N_5079,N_9518);
nand U12981 (N_12981,N_5632,N_9074);
xnor U12982 (N_12982,N_8077,N_9726);
nor U12983 (N_12983,N_8620,N_9192);
nand U12984 (N_12984,N_5138,N_9356);
nand U12985 (N_12985,N_8815,N_6949);
nor U12986 (N_12986,N_6706,N_8787);
and U12987 (N_12987,N_7283,N_8761);
nor U12988 (N_12988,N_6292,N_7580);
nor U12989 (N_12989,N_6337,N_6905);
and U12990 (N_12990,N_5577,N_5975);
nor U12991 (N_12991,N_8762,N_5669);
and U12992 (N_12992,N_6516,N_7826);
nor U12993 (N_12993,N_6096,N_9133);
nand U12994 (N_12994,N_8897,N_9779);
and U12995 (N_12995,N_6121,N_9982);
and U12996 (N_12996,N_9617,N_8012);
and U12997 (N_12997,N_6427,N_9131);
and U12998 (N_12998,N_7645,N_6111);
nor U12999 (N_12999,N_5550,N_6599);
and U13000 (N_13000,N_8130,N_8354);
nor U13001 (N_13001,N_5811,N_7237);
and U13002 (N_13002,N_9767,N_8298);
and U13003 (N_13003,N_5818,N_7075);
or U13004 (N_13004,N_6696,N_9893);
nor U13005 (N_13005,N_9243,N_6449);
nor U13006 (N_13006,N_6432,N_6590);
and U13007 (N_13007,N_5978,N_5028);
and U13008 (N_13008,N_9227,N_8760);
nand U13009 (N_13009,N_9039,N_9380);
and U13010 (N_13010,N_8579,N_7707);
nor U13011 (N_13011,N_5152,N_7079);
nand U13012 (N_13012,N_6283,N_9865);
and U13013 (N_13013,N_5731,N_5172);
nand U13014 (N_13014,N_9226,N_9081);
or U13015 (N_13015,N_8993,N_9467);
and U13016 (N_13016,N_7408,N_5494);
and U13017 (N_13017,N_7104,N_6732);
nor U13018 (N_13018,N_8240,N_7716);
and U13019 (N_13019,N_6135,N_9110);
nor U13020 (N_13020,N_8339,N_9531);
nor U13021 (N_13021,N_8940,N_9128);
nand U13022 (N_13022,N_9958,N_7987);
nor U13023 (N_13023,N_8540,N_9213);
and U13024 (N_13024,N_7814,N_5774);
and U13025 (N_13025,N_9864,N_6390);
and U13026 (N_13026,N_6033,N_6410);
nor U13027 (N_13027,N_7755,N_5553);
and U13028 (N_13028,N_6729,N_9040);
nor U13029 (N_13029,N_7512,N_8556);
or U13030 (N_13030,N_7159,N_9860);
nand U13031 (N_13031,N_5127,N_9716);
nor U13032 (N_13032,N_5363,N_7225);
nor U13033 (N_13033,N_6152,N_6310);
nor U13034 (N_13034,N_7780,N_6129);
nor U13035 (N_13035,N_9787,N_8405);
nor U13036 (N_13036,N_7040,N_7543);
nor U13037 (N_13037,N_7239,N_6503);
or U13038 (N_13038,N_7683,N_7294);
or U13039 (N_13039,N_8862,N_7756);
xnor U13040 (N_13040,N_5330,N_7148);
or U13041 (N_13041,N_6168,N_7161);
nor U13042 (N_13042,N_5034,N_8558);
or U13043 (N_13043,N_6261,N_5767);
nor U13044 (N_13044,N_5303,N_9139);
and U13045 (N_13045,N_9267,N_6964);
and U13046 (N_13046,N_5872,N_7256);
or U13047 (N_13047,N_5366,N_9441);
or U13048 (N_13048,N_8935,N_7348);
nor U13049 (N_13049,N_7561,N_8723);
and U13050 (N_13050,N_5730,N_7585);
nand U13051 (N_13051,N_9919,N_7467);
or U13052 (N_13052,N_6804,N_8331);
nand U13053 (N_13053,N_8801,N_9583);
or U13054 (N_13054,N_8299,N_5319);
nand U13055 (N_13055,N_7598,N_8111);
nor U13056 (N_13056,N_9810,N_8934);
or U13057 (N_13057,N_8814,N_9835);
nand U13058 (N_13058,N_8456,N_5902);
or U13059 (N_13059,N_9207,N_9244);
nand U13060 (N_13060,N_9920,N_7372);
and U13061 (N_13061,N_5907,N_9871);
nand U13062 (N_13062,N_5111,N_6266);
and U13063 (N_13063,N_6906,N_6655);
nor U13064 (N_13064,N_6368,N_5814);
or U13065 (N_13065,N_6569,N_7248);
or U13066 (N_13066,N_6520,N_7026);
or U13067 (N_13067,N_8629,N_5667);
or U13068 (N_13068,N_6719,N_5681);
and U13069 (N_13069,N_5993,N_5133);
or U13070 (N_13070,N_6006,N_5862);
nand U13071 (N_13071,N_8271,N_9360);
and U13072 (N_13072,N_6542,N_5733);
nor U13073 (N_13073,N_7389,N_7743);
nand U13074 (N_13074,N_6471,N_6103);
nor U13075 (N_13075,N_8674,N_9290);
nor U13076 (N_13076,N_9709,N_7208);
or U13077 (N_13077,N_7663,N_7489);
and U13078 (N_13078,N_9157,N_6123);
and U13079 (N_13079,N_7692,N_5437);
or U13080 (N_13080,N_6929,N_8675);
nor U13081 (N_13081,N_9915,N_7960);
and U13082 (N_13082,N_9971,N_5148);
or U13083 (N_13083,N_9692,N_6179);
nor U13084 (N_13084,N_5852,N_7980);
or U13085 (N_13085,N_8944,N_5309);
nor U13086 (N_13086,N_7210,N_5023);
nand U13087 (N_13087,N_7076,N_9531);
or U13088 (N_13088,N_6722,N_6778);
nand U13089 (N_13089,N_9123,N_6997);
nor U13090 (N_13090,N_8377,N_7967);
and U13091 (N_13091,N_6938,N_7500);
and U13092 (N_13092,N_8016,N_6520);
nand U13093 (N_13093,N_9626,N_7471);
nand U13094 (N_13094,N_8532,N_8947);
or U13095 (N_13095,N_6814,N_7910);
nand U13096 (N_13096,N_8498,N_9112);
xor U13097 (N_13097,N_9080,N_6230);
xnor U13098 (N_13098,N_9335,N_5214);
or U13099 (N_13099,N_6912,N_9537);
or U13100 (N_13100,N_9078,N_9911);
or U13101 (N_13101,N_6020,N_5539);
nand U13102 (N_13102,N_5359,N_5483);
nor U13103 (N_13103,N_9381,N_9072);
and U13104 (N_13104,N_7831,N_7539);
and U13105 (N_13105,N_8332,N_5195);
nand U13106 (N_13106,N_5083,N_7046);
or U13107 (N_13107,N_5003,N_8424);
nor U13108 (N_13108,N_6190,N_5730);
nor U13109 (N_13109,N_6912,N_6065);
and U13110 (N_13110,N_6739,N_7917);
or U13111 (N_13111,N_6680,N_7061);
and U13112 (N_13112,N_6276,N_7073);
nor U13113 (N_13113,N_5808,N_7084);
nand U13114 (N_13114,N_6830,N_9920);
and U13115 (N_13115,N_5081,N_7649);
and U13116 (N_13116,N_8236,N_9954);
and U13117 (N_13117,N_9110,N_5912);
nand U13118 (N_13118,N_7276,N_6250);
and U13119 (N_13119,N_5941,N_9596);
or U13120 (N_13120,N_9649,N_7770);
nand U13121 (N_13121,N_5859,N_9671);
nand U13122 (N_13122,N_8129,N_5362);
and U13123 (N_13123,N_9871,N_9845);
nand U13124 (N_13124,N_8322,N_8335);
and U13125 (N_13125,N_6282,N_5391);
nand U13126 (N_13126,N_9997,N_6047);
and U13127 (N_13127,N_9079,N_8588);
or U13128 (N_13128,N_5955,N_8281);
or U13129 (N_13129,N_6604,N_6125);
nand U13130 (N_13130,N_9154,N_8941);
or U13131 (N_13131,N_9003,N_9514);
and U13132 (N_13132,N_5016,N_7010);
nand U13133 (N_13133,N_8910,N_6817);
nor U13134 (N_13134,N_5654,N_6071);
xor U13135 (N_13135,N_6495,N_7965);
or U13136 (N_13136,N_6802,N_9421);
or U13137 (N_13137,N_5290,N_7383);
and U13138 (N_13138,N_5393,N_7018);
nand U13139 (N_13139,N_7121,N_5541);
and U13140 (N_13140,N_9824,N_8447);
nand U13141 (N_13141,N_8320,N_5696);
nand U13142 (N_13142,N_6756,N_6893);
and U13143 (N_13143,N_9251,N_9044);
nor U13144 (N_13144,N_8873,N_8316);
nor U13145 (N_13145,N_8364,N_9289);
nor U13146 (N_13146,N_8225,N_7443);
nand U13147 (N_13147,N_5903,N_9620);
and U13148 (N_13148,N_8472,N_9620);
or U13149 (N_13149,N_7593,N_5540);
and U13150 (N_13150,N_7775,N_8847);
nor U13151 (N_13151,N_9664,N_5069);
nor U13152 (N_13152,N_5165,N_6819);
and U13153 (N_13153,N_5874,N_5102);
or U13154 (N_13154,N_6655,N_8002);
and U13155 (N_13155,N_9889,N_5164);
and U13156 (N_13156,N_8288,N_9535);
and U13157 (N_13157,N_7797,N_6106);
or U13158 (N_13158,N_6057,N_7611);
or U13159 (N_13159,N_5178,N_5111);
nand U13160 (N_13160,N_7316,N_7441);
nor U13161 (N_13161,N_9334,N_6452);
nand U13162 (N_13162,N_5492,N_8352);
or U13163 (N_13163,N_9438,N_7790);
nand U13164 (N_13164,N_8114,N_9553);
nand U13165 (N_13165,N_9738,N_7863);
and U13166 (N_13166,N_5683,N_7782);
and U13167 (N_13167,N_5851,N_5827);
nor U13168 (N_13168,N_9993,N_6493);
nand U13169 (N_13169,N_7244,N_6483);
and U13170 (N_13170,N_8357,N_9030);
nand U13171 (N_13171,N_6302,N_5564);
or U13172 (N_13172,N_8142,N_6889);
nand U13173 (N_13173,N_7337,N_6845);
nand U13174 (N_13174,N_7534,N_7032);
nor U13175 (N_13175,N_7081,N_5699);
nor U13176 (N_13176,N_5918,N_6177);
and U13177 (N_13177,N_5648,N_5866);
or U13178 (N_13178,N_7012,N_9715);
nand U13179 (N_13179,N_9424,N_6975);
nor U13180 (N_13180,N_5695,N_9195);
nand U13181 (N_13181,N_9614,N_7638);
and U13182 (N_13182,N_8770,N_7609);
nor U13183 (N_13183,N_9746,N_9432);
or U13184 (N_13184,N_9355,N_8100);
or U13185 (N_13185,N_9256,N_7673);
nand U13186 (N_13186,N_9741,N_5537);
nor U13187 (N_13187,N_8951,N_7328);
and U13188 (N_13188,N_5806,N_7474);
nand U13189 (N_13189,N_8410,N_6035);
nand U13190 (N_13190,N_6216,N_5978);
and U13191 (N_13191,N_9488,N_8394);
xnor U13192 (N_13192,N_6940,N_8084);
nand U13193 (N_13193,N_6353,N_9023);
nand U13194 (N_13194,N_9267,N_6340);
nor U13195 (N_13195,N_9912,N_8107);
nor U13196 (N_13196,N_8311,N_7221);
or U13197 (N_13197,N_8130,N_5429);
nand U13198 (N_13198,N_8467,N_6226);
nand U13199 (N_13199,N_6733,N_9394);
and U13200 (N_13200,N_8662,N_7014);
or U13201 (N_13201,N_8882,N_9419);
or U13202 (N_13202,N_7242,N_8366);
nor U13203 (N_13203,N_8969,N_7889);
and U13204 (N_13204,N_6437,N_5778);
or U13205 (N_13205,N_6465,N_9861);
or U13206 (N_13206,N_7624,N_9480);
nor U13207 (N_13207,N_8921,N_7416);
and U13208 (N_13208,N_8033,N_5084);
nor U13209 (N_13209,N_5652,N_9139);
nor U13210 (N_13210,N_6698,N_8478);
nand U13211 (N_13211,N_5514,N_6536);
nand U13212 (N_13212,N_6942,N_6715);
or U13213 (N_13213,N_5399,N_9309);
or U13214 (N_13214,N_6768,N_8237);
or U13215 (N_13215,N_6691,N_9391);
and U13216 (N_13216,N_5899,N_8706);
and U13217 (N_13217,N_8427,N_6226);
or U13218 (N_13218,N_7425,N_8452);
or U13219 (N_13219,N_9960,N_6523);
or U13220 (N_13220,N_7465,N_9564);
or U13221 (N_13221,N_7412,N_5854);
and U13222 (N_13222,N_6084,N_8182);
and U13223 (N_13223,N_7931,N_9260);
nand U13224 (N_13224,N_7605,N_6527);
xnor U13225 (N_13225,N_5898,N_6507);
nor U13226 (N_13226,N_6517,N_7548);
nor U13227 (N_13227,N_8600,N_7172);
or U13228 (N_13228,N_8301,N_7669);
or U13229 (N_13229,N_7819,N_6087);
nor U13230 (N_13230,N_9710,N_5455);
nor U13231 (N_13231,N_8542,N_9696);
and U13232 (N_13232,N_8684,N_6232);
nor U13233 (N_13233,N_8773,N_9842);
nor U13234 (N_13234,N_6903,N_9270);
nand U13235 (N_13235,N_7850,N_7899);
nand U13236 (N_13236,N_6351,N_6406);
and U13237 (N_13237,N_8738,N_8138);
or U13238 (N_13238,N_8051,N_5567);
nand U13239 (N_13239,N_8837,N_6227);
xor U13240 (N_13240,N_9988,N_5447);
or U13241 (N_13241,N_5556,N_7253);
or U13242 (N_13242,N_7968,N_9199);
or U13243 (N_13243,N_8666,N_6731);
or U13244 (N_13244,N_5055,N_6821);
xnor U13245 (N_13245,N_5010,N_5711);
nor U13246 (N_13246,N_8707,N_6042);
and U13247 (N_13247,N_6171,N_8570);
or U13248 (N_13248,N_8144,N_8968);
nor U13249 (N_13249,N_5196,N_6451);
nor U13250 (N_13250,N_9900,N_9521);
and U13251 (N_13251,N_6227,N_6964);
nand U13252 (N_13252,N_7214,N_6330);
nor U13253 (N_13253,N_7567,N_8566);
and U13254 (N_13254,N_9536,N_8625);
or U13255 (N_13255,N_7216,N_6540);
or U13256 (N_13256,N_5548,N_8567);
or U13257 (N_13257,N_5785,N_7555);
nand U13258 (N_13258,N_5568,N_6274);
nand U13259 (N_13259,N_7720,N_6348);
and U13260 (N_13260,N_9424,N_5991);
or U13261 (N_13261,N_5549,N_6694);
nor U13262 (N_13262,N_7685,N_9393);
and U13263 (N_13263,N_8211,N_7009);
or U13264 (N_13264,N_9351,N_9603);
or U13265 (N_13265,N_7610,N_8242);
nand U13266 (N_13266,N_5883,N_9174);
nand U13267 (N_13267,N_6450,N_6659);
nor U13268 (N_13268,N_5710,N_6249);
or U13269 (N_13269,N_7006,N_6107);
nor U13270 (N_13270,N_6312,N_6398);
or U13271 (N_13271,N_8854,N_5891);
or U13272 (N_13272,N_9643,N_9321);
or U13273 (N_13273,N_8299,N_9113);
nor U13274 (N_13274,N_8091,N_5335);
or U13275 (N_13275,N_5736,N_6250);
or U13276 (N_13276,N_8553,N_6996);
nand U13277 (N_13277,N_6831,N_8270);
or U13278 (N_13278,N_6783,N_8555);
nor U13279 (N_13279,N_8699,N_7736);
xor U13280 (N_13280,N_7883,N_5790);
or U13281 (N_13281,N_6911,N_9439);
or U13282 (N_13282,N_8288,N_5559);
or U13283 (N_13283,N_9193,N_9076);
and U13284 (N_13284,N_9422,N_7027);
and U13285 (N_13285,N_9956,N_7611);
and U13286 (N_13286,N_7686,N_5050);
or U13287 (N_13287,N_9894,N_9353);
nor U13288 (N_13288,N_6967,N_6139);
or U13289 (N_13289,N_8289,N_7641);
nor U13290 (N_13290,N_8830,N_7112);
and U13291 (N_13291,N_5018,N_7299);
and U13292 (N_13292,N_6202,N_7346);
nor U13293 (N_13293,N_9548,N_5152);
or U13294 (N_13294,N_5274,N_5110);
or U13295 (N_13295,N_7655,N_5853);
nor U13296 (N_13296,N_7045,N_9305);
and U13297 (N_13297,N_9422,N_9942);
nor U13298 (N_13298,N_8102,N_8481);
nor U13299 (N_13299,N_9289,N_9522);
nor U13300 (N_13300,N_9460,N_9092);
and U13301 (N_13301,N_6687,N_9378);
or U13302 (N_13302,N_7591,N_6224);
or U13303 (N_13303,N_7539,N_8548);
or U13304 (N_13304,N_6650,N_7954);
and U13305 (N_13305,N_8727,N_9834);
nand U13306 (N_13306,N_7923,N_7634);
or U13307 (N_13307,N_5350,N_6629);
and U13308 (N_13308,N_5180,N_7991);
and U13309 (N_13309,N_7476,N_7842);
xor U13310 (N_13310,N_5825,N_7836);
or U13311 (N_13311,N_9669,N_5355);
and U13312 (N_13312,N_8580,N_6930);
nor U13313 (N_13313,N_6212,N_5274);
nand U13314 (N_13314,N_8086,N_6227);
or U13315 (N_13315,N_5598,N_9356);
nand U13316 (N_13316,N_6631,N_7752);
and U13317 (N_13317,N_6486,N_7641);
or U13318 (N_13318,N_5847,N_7800);
or U13319 (N_13319,N_8504,N_6097);
and U13320 (N_13320,N_8810,N_6514);
nand U13321 (N_13321,N_5389,N_8009);
and U13322 (N_13322,N_9305,N_7105);
nand U13323 (N_13323,N_5759,N_5543);
or U13324 (N_13324,N_6463,N_5911);
and U13325 (N_13325,N_7013,N_7164);
or U13326 (N_13326,N_7832,N_5302);
nand U13327 (N_13327,N_8306,N_9719);
or U13328 (N_13328,N_7481,N_9831);
and U13329 (N_13329,N_9140,N_7359);
and U13330 (N_13330,N_9510,N_6821);
nand U13331 (N_13331,N_9199,N_5178);
and U13332 (N_13332,N_5424,N_6458);
nand U13333 (N_13333,N_6460,N_5044);
nand U13334 (N_13334,N_8880,N_6957);
nor U13335 (N_13335,N_8938,N_9040);
nand U13336 (N_13336,N_5866,N_8988);
nand U13337 (N_13337,N_5579,N_7886);
nor U13338 (N_13338,N_5311,N_9636);
and U13339 (N_13339,N_7953,N_5902);
nand U13340 (N_13340,N_6811,N_6910);
or U13341 (N_13341,N_6949,N_7201);
and U13342 (N_13342,N_6278,N_8149);
nand U13343 (N_13343,N_9092,N_9642);
nand U13344 (N_13344,N_9017,N_6517);
and U13345 (N_13345,N_7084,N_9487);
nor U13346 (N_13346,N_7785,N_7158);
nand U13347 (N_13347,N_7634,N_5549);
nor U13348 (N_13348,N_9658,N_9932);
nand U13349 (N_13349,N_8109,N_5916);
and U13350 (N_13350,N_8246,N_8706);
and U13351 (N_13351,N_8853,N_7685);
and U13352 (N_13352,N_9564,N_9123);
nor U13353 (N_13353,N_8888,N_8849);
or U13354 (N_13354,N_6201,N_8489);
nor U13355 (N_13355,N_8303,N_5935);
xor U13356 (N_13356,N_6008,N_9079);
nor U13357 (N_13357,N_6781,N_5281);
or U13358 (N_13358,N_9987,N_8034);
and U13359 (N_13359,N_8285,N_8636);
and U13360 (N_13360,N_8154,N_9883);
nor U13361 (N_13361,N_7087,N_6494);
nand U13362 (N_13362,N_7742,N_6153);
or U13363 (N_13363,N_8943,N_9103);
or U13364 (N_13364,N_5301,N_7865);
xor U13365 (N_13365,N_8476,N_8000);
and U13366 (N_13366,N_7564,N_7088);
nor U13367 (N_13367,N_5222,N_5904);
nand U13368 (N_13368,N_5231,N_5204);
nand U13369 (N_13369,N_6368,N_7774);
and U13370 (N_13370,N_7247,N_9181);
nor U13371 (N_13371,N_5735,N_9631);
nor U13372 (N_13372,N_8713,N_7488);
nand U13373 (N_13373,N_9982,N_5724);
and U13374 (N_13374,N_6661,N_6012);
or U13375 (N_13375,N_5119,N_9685);
and U13376 (N_13376,N_7665,N_6197);
nand U13377 (N_13377,N_6963,N_6262);
xnor U13378 (N_13378,N_7544,N_7342);
xnor U13379 (N_13379,N_5799,N_7948);
nand U13380 (N_13380,N_9568,N_8038);
nor U13381 (N_13381,N_6524,N_6245);
and U13382 (N_13382,N_8596,N_5138);
nand U13383 (N_13383,N_6792,N_6008);
nand U13384 (N_13384,N_5594,N_5867);
nor U13385 (N_13385,N_9962,N_7938);
nor U13386 (N_13386,N_8213,N_7515);
and U13387 (N_13387,N_7621,N_5717);
nand U13388 (N_13388,N_6959,N_9951);
nand U13389 (N_13389,N_9316,N_9558);
and U13390 (N_13390,N_8141,N_8944);
or U13391 (N_13391,N_5821,N_5994);
nand U13392 (N_13392,N_8804,N_9422);
or U13393 (N_13393,N_8814,N_9681);
nand U13394 (N_13394,N_9029,N_5981);
nor U13395 (N_13395,N_7713,N_8551);
and U13396 (N_13396,N_6421,N_9101);
nor U13397 (N_13397,N_7323,N_9218);
or U13398 (N_13398,N_8626,N_9033);
and U13399 (N_13399,N_5367,N_6182);
or U13400 (N_13400,N_6404,N_6617);
nor U13401 (N_13401,N_8322,N_8659);
nand U13402 (N_13402,N_9170,N_7400);
nor U13403 (N_13403,N_9322,N_5904);
and U13404 (N_13404,N_5415,N_7510);
or U13405 (N_13405,N_9161,N_9516);
nor U13406 (N_13406,N_5214,N_7972);
nand U13407 (N_13407,N_5406,N_5133);
and U13408 (N_13408,N_8231,N_8413);
nand U13409 (N_13409,N_5847,N_5150);
and U13410 (N_13410,N_6789,N_6283);
nand U13411 (N_13411,N_8338,N_8308);
or U13412 (N_13412,N_7927,N_9805);
or U13413 (N_13413,N_5778,N_5450);
nor U13414 (N_13414,N_7421,N_8651);
or U13415 (N_13415,N_7263,N_6033);
nor U13416 (N_13416,N_8170,N_7820);
or U13417 (N_13417,N_5108,N_7795);
or U13418 (N_13418,N_5564,N_7618);
nor U13419 (N_13419,N_6115,N_8787);
or U13420 (N_13420,N_5817,N_9871);
and U13421 (N_13421,N_7416,N_5515);
and U13422 (N_13422,N_7346,N_8492);
nand U13423 (N_13423,N_8163,N_8146);
nand U13424 (N_13424,N_8007,N_8077);
or U13425 (N_13425,N_7995,N_9249);
nand U13426 (N_13426,N_8548,N_7620);
and U13427 (N_13427,N_9819,N_8547);
nor U13428 (N_13428,N_5692,N_8382);
nand U13429 (N_13429,N_9780,N_5535);
nand U13430 (N_13430,N_5821,N_8424);
or U13431 (N_13431,N_9955,N_8542);
or U13432 (N_13432,N_9934,N_5372);
or U13433 (N_13433,N_6812,N_6368);
or U13434 (N_13434,N_8631,N_5884);
and U13435 (N_13435,N_5147,N_7843);
nor U13436 (N_13436,N_5155,N_5512);
or U13437 (N_13437,N_7390,N_8552);
and U13438 (N_13438,N_5646,N_9423);
xor U13439 (N_13439,N_5595,N_7533);
and U13440 (N_13440,N_5709,N_6286);
or U13441 (N_13441,N_5088,N_5443);
nand U13442 (N_13442,N_8071,N_8352);
and U13443 (N_13443,N_7107,N_7297);
and U13444 (N_13444,N_9849,N_9837);
nand U13445 (N_13445,N_8047,N_5587);
nand U13446 (N_13446,N_8414,N_6526);
and U13447 (N_13447,N_5463,N_8196);
nand U13448 (N_13448,N_7979,N_8570);
nand U13449 (N_13449,N_7785,N_9020);
nand U13450 (N_13450,N_8340,N_8712);
and U13451 (N_13451,N_7552,N_6345);
or U13452 (N_13452,N_9736,N_7148);
nand U13453 (N_13453,N_5256,N_7164);
and U13454 (N_13454,N_9746,N_7486);
nand U13455 (N_13455,N_8604,N_8091);
and U13456 (N_13456,N_9955,N_7226);
xnor U13457 (N_13457,N_7210,N_6769);
nor U13458 (N_13458,N_5740,N_6157);
or U13459 (N_13459,N_5009,N_9977);
and U13460 (N_13460,N_7853,N_8124);
or U13461 (N_13461,N_6864,N_6637);
nand U13462 (N_13462,N_7892,N_7346);
xnor U13463 (N_13463,N_8625,N_8587);
or U13464 (N_13464,N_6568,N_7555);
and U13465 (N_13465,N_5358,N_7354);
nor U13466 (N_13466,N_8440,N_9330);
or U13467 (N_13467,N_6888,N_6025);
or U13468 (N_13468,N_8984,N_9129);
nor U13469 (N_13469,N_9480,N_8960);
nor U13470 (N_13470,N_8852,N_7052);
or U13471 (N_13471,N_9476,N_6305);
nand U13472 (N_13472,N_9343,N_7654);
or U13473 (N_13473,N_6092,N_7348);
nand U13474 (N_13474,N_6485,N_8933);
nand U13475 (N_13475,N_6509,N_5065);
nand U13476 (N_13476,N_8059,N_5078);
or U13477 (N_13477,N_5678,N_9754);
nor U13478 (N_13478,N_6499,N_5809);
xnor U13479 (N_13479,N_8168,N_6076);
nor U13480 (N_13480,N_5662,N_8526);
and U13481 (N_13481,N_5855,N_9418);
nor U13482 (N_13482,N_5445,N_8931);
and U13483 (N_13483,N_5093,N_6354);
and U13484 (N_13484,N_8006,N_6787);
or U13485 (N_13485,N_5791,N_5188);
or U13486 (N_13486,N_7714,N_8881);
nand U13487 (N_13487,N_5019,N_9442);
nor U13488 (N_13488,N_6186,N_6235);
or U13489 (N_13489,N_5839,N_6910);
xnor U13490 (N_13490,N_6795,N_7194);
nor U13491 (N_13491,N_7759,N_7166);
or U13492 (N_13492,N_9888,N_9739);
nor U13493 (N_13493,N_8779,N_7664);
and U13494 (N_13494,N_7507,N_7161);
and U13495 (N_13495,N_9902,N_5057);
and U13496 (N_13496,N_5051,N_9811);
and U13497 (N_13497,N_5593,N_7120);
nor U13498 (N_13498,N_7213,N_8681);
or U13499 (N_13499,N_9618,N_8907);
nand U13500 (N_13500,N_7270,N_8899);
or U13501 (N_13501,N_9096,N_6095);
nand U13502 (N_13502,N_9911,N_7535);
and U13503 (N_13503,N_5734,N_7155);
nor U13504 (N_13504,N_9489,N_6578);
nor U13505 (N_13505,N_9825,N_8035);
or U13506 (N_13506,N_7944,N_5760);
or U13507 (N_13507,N_6046,N_5605);
nor U13508 (N_13508,N_8532,N_7740);
and U13509 (N_13509,N_7739,N_8867);
and U13510 (N_13510,N_8163,N_7919);
and U13511 (N_13511,N_9734,N_6357);
nand U13512 (N_13512,N_7268,N_9828);
nand U13513 (N_13513,N_5672,N_9290);
and U13514 (N_13514,N_5771,N_8925);
nand U13515 (N_13515,N_6502,N_9228);
or U13516 (N_13516,N_9875,N_9745);
and U13517 (N_13517,N_9165,N_8114);
nor U13518 (N_13518,N_5307,N_6080);
or U13519 (N_13519,N_8031,N_7787);
and U13520 (N_13520,N_7985,N_5284);
and U13521 (N_13521,N_8168,N_5918);
nor U13522 (N_13522,N_6936,N_6497);
or U13523 (N_13523,N_6943,N_7157);
nor U13524 (N_13524,N_8436,N_6770);
nand U13525 (N_13525,N_8568,N_6269);
or U13526 (N_13526,N_8558,N_9017);
nand U13527 (N_13527,N_7757,N_5586);
or U13528 (N_13528,N_9437,N_6019);
nand U13529 (N_13529,N_5550,N_6449);
nor U13530 (N_13530,N_5744,N_6909);
or U13531 (N_13531,N_7398,N_8167);
nor U13532 (N_13532,N_9594,N_6105);
and U13533 (N_13533,N_6969,N_5702);
and U13534 (N_13534,N_6897,N_7576);
nand U13535 (N_13535,N_9395,N_5697);
nor U13536 (N_13536,N_7633,N_5991);
nor U13537 (N_13537,N_9639,N_8443);
nand U13538 (N_13538,N_9633,N_8812);
or U13539 (N_13539,N_5579,N_6291);
nand U13540 (N_13540,N_8051,N_7037);
or U13541 (N_13541,N_9685,N_9841);
or U13542 (N_13542,N_7638,N_6836);
and U13543 (N_13543,N_9165,N_7309);
nor U13544 (N_13544,N_6647,N_9020);
and U13545 (N_13545,N_6310,N_9259);
or U13546 (N_13546,N_8700,N_7065);
nand U13547 (N_13547,N_8460,N_9596);
nand U13548 (N_13548,N_7041,N_9271);
nand U13549 (N_13549,N_6648,N_8793);
or U13550 (N_13550,N_6907,N_6234);
or U13551 (N_13551,N_6428,N_7811);
or U13552 (N_13552,N_5973,N_5955);
nand U13553 (N_13553,N_7345,N_5353);
nand U13554 (N_13554,N_6601,N_6381);
and U13555 (N_13555,N_5539,N_5235);
or U13556 (N_13556,N_5489,N_9518);
or U13557 (N_13557,N_6320,N_5205);
or U13558 (N_13558,N_8370,N_9608);
nand U13559 (N_13559,N_7333,N_9513);
or U13560 (N_13560,N_9833,N_8469);
or U13561 (N_13561,N_7932,N_9437);
nor U13562 (N_13562,N_9415,N_9657);
nor U13563 (N_13563,N_9902,N_6672);
and U13564 (N_13564,N_9905,N_6492);
nand U13565 (N_13565,N_7213,N_8919);
nand U13566 (N_13566,N_7809,N_5659);
or U13567 (N_13567,N_9461,N_9380);
nor U13568 (N_13568,N_8573,N_7597);
or U13569 (N_13569,N_5744,N_6849);
and U13570 (N_13570,N_6590,N_6888);
nor U13571 (N_13571,N_6173,N_5881);
and U13572 (N_13572,N_9625,N_8706);
nor U13573 (N_13573,N_6344,N_6858);
and U13574 (N_13574,N_5883,N_7054);
nand U13575 (N_13575,N_6934,N_7382);
and U13576 (N_13576,N_9847,N_8760);
or U13577 (N_13577,N_7778,N_8401);
or U13578 (N_13578,N_7567,N_8950);
or U13579 (N_13579,N_8268,N_8981);
nand U13580 (N_13580,N_8643,N_9111);
nand U13581 (N_13581,N_5728,N_8247);
nand U13582 (N_13582,N_7891,N_5078);
nand U13583 (N_13583,N_5655,N_9689);
nor U13584 (N_13584,N_9481,N_7672);
and U13585 (N_13585,N_7192,N_5998);
or U13586 (N_13586,N_6973,N_5707);
and U13587 (N_13587,N_9357,N_6469);
xnor U13588 (N_13588,N_9490,N_6460);
and U13589 (N_13589,N_9670,N_9344);
nor U13590 (N_13590,N_6367,N_6286);
or U13591 (N_13591,N_9619,N_5890);
nor U13592 (N_13592,N_5549,N_9602);
nand U13593 (N_13593,N_5964,N_5908);
and U13594 (N_13594,N_5934,N_9098);
or U13595 (N_13595,N_7644,N_5794);
nand U13596 (N_13596,N_7373,N_7809);
nor U13597 (N_13597,N_9843,N_6572);
nand U13598 (N_13598,N_8291,N_7175);
or U13599 (N_13599,N_8122,N_8276);
nor U13600 (N_13600,N_9764,N_6730);
or U13601 (N_13601,N_9892,N_8540);
or U13602 (N_13602,N_5728,N_8279);
or U13603 (N_13603,N_6520,N_7215);
and U13604 (N_13604,N_7906,N_8745);
and U13605 (N_13605,N_8894,N_5293);
nor U13606 (N_13606,N_7169,N_9109);
or U13607 (N_13607,N_7968,N_6044);
nor U13608 (N_13608,N_8953,N_7941);
nand U13609 (N_13609,N_9516,N_8050);
or U13610 (N_13610,N_6823,N_7975);
nand U13611 (N_13611,N_8147,N_9018);
nor U13612 (N_13612,N_8464,N_6544);
and U13613 (N_13613,N_5121,N_8777);
nor U13614 (N_13614,N_9334,N_7247);
or U13615 (N_13615,N_5977,N_9737);
nor U13616 (N_13616,N_5725,N_5359);
and U13617 (N_13617,N_6825,N_5889);
and U13618 (N_13618,N_7182,N_8444);
nand U13619 (N_13619,N_7995,N_6580);
nor U13620 (N_13620,N_5230,N_5131);
nor U13621 (N_13621,N_7437,N_6505);
nand U13622 (N_13622,N_5049,N_6624);
and U13623 (N_13623,N_5969,N_8751);
nand U13624 (N_13624,N_9731,N_8537);
nor U13625 (N_13625,N_9967,N_6336);
or U13626 (N_13626,N_9952,N_8276);
or U13627 (N_13627,N_9590,N_6822);
nor U13628 (N_13628,N_9476,N_9523);
nor U13629 (N_13629,N_9995,N_5274);
nand U13630 (N_13630,N_7679,N_9554);
nor U13631 (N_13631,N_6728,N_9087);
and U13632 (N_13632,N_7070,N_5223);
nor U13633 (N_13633,N_5929,N_7123);
or U13634 (N_13634,N_6642,N_6049);
and U13635 (N_13635,N_7492,N_6614);
and U13636 (N_13636,N_7756,N_6211);
nand U13637 (N_13637,N_6799,N_5231);
nand U13638 (N_13638,N_8675,N_7649);
nor U13639 (N_13639,N_7535,N_7959);
nor U13640 (N_13640,N_8142,N_8710);
nand U13641 (N_13641,N_7011,N_6689);
nand U13642 (N_13642,N_9015,N_9757);
or U13643 (N_13643,N_6195,N_6298);
nand U13644 (N_13644,N_8547,N_5570);
and U13645 (N_13645,N_5486,N_6199);
or U13646 (N_13646,N_6308,N_7216);
and U13647 (N_13647,N_6439,N_6032);
xor U13648 (N_13648,N_5133,N_7201);
nor U13649 (N_13649,N_7094,N_7597);
nand U13650 (N_13650,N_6097,N_6662);
nor U13651 (N_13651,N_6832,N_8390);
or U13652 (N_13652,N_9289,N_5095);
and U13653 (N_13653,N_7838,N_8546);
or U13654 (N_13654,N_9449,N_6465);
and U13655 (N_13655,N_8780,N_9241);
nor U13656 (N_13656,N_5566,N_6039);
or U13657 (N_13657,N_6320,N_7722);
nor U13658 (N_13658,N_6491,N_5867);
nand U13659 (N_13659,N_5868,N_9923);
and U13660 (N_13660,N_7058,N_9090);
or U13661 (N_13661,N_8447,N_7925);
nor U13662 (N_13662,N_8825,N_6397);
nand U13663 (N_13663,N_8506,N_9106);
nor U13664 (N_13664,N_5765,N_5071);
nor U13665 (N_13665,N_7754,N_5394);
xnor U13666 (N_13666,N_7726,N_7016);
or U13667 (N_13667,N_9048,N_5180);
nor U13668 (N_13668,N_8962,N_7699);
or U13669 (N_13669,N_7447,N_8723);
or U13670 (N_13670,N_8751,N_5863);
nor U13671 (N_13671,N_8443,N_7713);
nand U13672 (N_13672,N_6927,N_6976);
nor U13673 (N_13673,N_7533,N_6413);
and U13674 (N_13674,N_8430,N_6692);
nor U13675 (N_13675,N_8808,N_8957);
or U13676 (N_13676,N_7231,N_7763);
or U13677 (N_13677,N_7621,N_6243);
and U13678 (N_13678,N_7987,N_8742);
and U13679 (N_13679,N_6158,N_6909);
and U13680 (N_13680,N_8792,N_8625);
nor U13681 (N_13681,N_7251,N_5420);
nor U13682 (N_13682,N_5867,N_9424);
nor U13683 (N_13683,N_7840,N_8419);
nand U13684 (N_13684,N_9509,N_8818);
xnor U13685 (N_13685,N_8332,N_7450);
or U13686 (N_13686,N_9929,N_9205);
nor U13687 (N_13687,N_5462,N_8432);
and U13688 (N_13688,N_6379,N_6867);
nor U13689 (N_13689,N_8895,N_7221);
or U13690 (N_13690,N_5920,N_9352);
nor U13691 (N_13691,N_9622,N_9844);
nand U13692 (N_13692,N_6493,N_9087);
nor U13693 (N_13693,N_5880,N_6300);
nand U13694 (N_13694,N_9466,N_8692);
nor U13695 (N_13695,N_8758,N_7149);
and U13696 (N_13696,N_5570,N_6799);
nor U13697 (N_13697,N_9261,N_8890);
nand U13698 (N_13698,N_7202,N_7586);
nand U13699 (N_13699,N_5029,N_5507);
and U13700 (N_13700,N_7840,N_5274);
nand U13701 (N_13701,N_7466,N_5310);
or U13702 (N_13702,N_5364,N_8361);
nor U13703 (N_13703,N_8283,N_9848);
nor U13704 (N_13704,N_6149,N_5488);
xnor U13705 (N_13705,N_6398,N_7783);
nor U13706 (N_13706,N_9621,N_8177);
nor U13707 (N_13707,N_9968,N_8515);
nor U13708 (N_13708,N_6729,N_5407);
nor U13709 (N_13709,N_9159,N_7134);
or U13710 (N_13710,N_6334,N_5623);
nor U13711 (N_13711,N_7057,N_5694);
or U13712 (N_13712,N_9943,N_5040);
nor U13713 (N_13713,N_6761,N_7993);
or U13714 (N_13714,N_9979,N_8700);
nor U13715 (N_13715,N_6408,N_7627);
and U13716 (N_13716,N_9716,N_9204);
nor U13717 (N_13717,N_8533,N_6782);
and U13718 (N_13718,N_6565,N_9661);
nor U13719 (N_13719,N_8271,N_5561);
nor U13720 (N_13720,N_6198,N_8790);
and U13721 (N_13721,N_6516,N_5625);
nand U13722 (N_13722,N_7364,N_6387);
or U13723 (N_13723,N_5370,N_5012);
and U13724 (N_13724,N_9686,N_6114);
and U13725 (N_13725,N_8753,N_5963);
nor U13726 (N_13726,N_6870,N_5647);
nand U13727 (N_13727,N_9506,N_8551);
or U13728 (N_13728,N_9034,N_7731);
and U13729 (N_13729,N_7409,N_9974);
or U13730 (N_13730,N_6963,N_7036);
or U13731 (N_13731,N_7003,N_9696);
nor U13732 (N_13732,N_6343,N_7009);
nor U13733 (N_13733,N_6118,N_8043);
and U13734 (N_13734,N_7287,N_9849);
nor U13735 (N_13735,N_5263,N_7009);
nor U13736 (N_13736,N_5184,N_7139);
nor U13737 (N_13737,N_5997,N_5189);
and U13738 (N_13738,N_9555,N_8793);
or U13739 (N_13739,N_9656,N_7546);
or U13740 (N_13740,N_6011,N_6808);
nand U13741 (N_13741,N_5392,N_8524);
or U13742 (N_13742,N_5172,N_5610);
nor U13743 (N_13743,N_9339,N_6523);
nand U13744 (N_13744,N_9078,N_7842);
nor U13745 (N_13745,N_8994,N_6214);
or U13746 (N_13746,N_7915,N_8835);
and U13747 (N_13747,N_7797,N_9161);
or U13748 (N_13748,N_7201,N_7014);
nor U13749 (N_13749,N_7990,N_6952);
and U13750 (N_13750,N_7916,N_8690);
and U13751 (N_13751,N_7714,N_9888);
nor U13752 (N_13752,N_6163,N_8970);
or U13753 (N_13753,N_9038,N_9696);
or U13754 (N_13754,N_8551,N_6112);
nor U13755 (N_13755,N_7505,N_7440);
nand U13756 (N_13756,N_6728,N_5847);
or U13757 (N_13757,N_6063,N_8078);
and U13758 (N_13758,N_6106,N_6296);
nor U13759 (N_13759,N_9067,N_6407);
xnor U13760 (N_13760,N_5521,N_6304);
nand U13761 (N_13761,N_8809,N_5673);
nand U13762 (N_13762,N_6322,N_6958);
or U13763 (N_13763,N_7940,N_5293);
nand U13764 (N_13764,N_9762,N_7462);
and U13765 (N_13765,N_8342,N_6305);
xnor U13766 (N_13766,N_9960,N_8257);
nand U13767 (N_13767,N_8279,N_9516);
nor U13768 (N_13768,N_8933,N_6076);
nor U13769 (N_13769,N_8640,N_8174);
or U13770 (N_13770,N_6205,N_5609);
or U13771 (N_13771,N_9821,N_9315);
nand U13772 (N_13772,N_8561,N_6103);
nand U13773 (N_13773,N_9353,N_8812);
nand U13774 (N_13774,N_8020,N_6469);
nand U13775 (N_13775,N_6540,N_7301);
nand U13776 (N_13776,N_8961,N_7008);
nand U13777 (N_13777,N_7220,N_8189);
or U13778 (N_13778,N_7323,N_5198);
nand U13779 (N_13779,N_6860,N_7442);
nand U13780 (N_13780,N_9824,N_9510);
nand U13781 (N_13781,N_7111,N_9537);
nor U13782 (N_13782,N_6917,N_7208);
nand U13783 (N_13783,N_9288,N_5891);
nor U13784 (N_13784,N_7855,N_7033);
xnor U13785 (N_13785,N_7499,N_6146);
nand U13786 (N_13786,N_7594,N_8827);
nand U13787 (N_13787,N_7372,N_6561);
and U13788 (N_13788,N_7841,N_7332);
or U13789 (N_13789,N_6307,N_9137);
nand U13790 (N_13790,N_9455,N_6483);
or U13791 (N_13791,N_9189,N_9477);
or U13792 (N_13792,N_7614,N_5427);
or U13793 (N_13793,N_6430,N_7561);
nand U13794 (N_13794,N_7659,N_8932);
nand U13795 (N_13795,N_5701,N_9621);
and U13796 (N_13796,N_8464,N_7255);
or U13797 (N_13797,N_7486,N_6737);
nor U13798 (N_13798,N_8082,N_8370);
nor U13799 (N_13799,N_6293,N_7233);
or U13800 (N_13800,N_9417,N_9724);
nor U13801 (N_13801,N_9526,N_8137);
or U13802 (N_13802,N_8635,N_8224);
or U13803 (N_13803,N_5705,N_6227);
nand U13804 (N_13804,N_7317,N_5605);
or U13805 (N_13805,N_9802,N_5323);
nor U13806 (N_13806,N_8011,N_6139);
nor U13807 (N_13807,N_6198,N_6173);
and U13808 (N_13808,N_5427,N_7872);
or U13809 (N_13809,N_7093,N_5326);
or U13810 (N_13810,N_7388,N_8190);
xnor U13811 (N_13811,N_5249,N_7084);
or U13812 (N_13812,N_9357,N_8056);
nand U13813 (N_13813,N_6092,N_8062);
and U13814 (N_13814,N_8152,N_8130);
and U13815 (N_13815,N_7223,N_5491);
nor U13816 (N_13816,N_5840,N_6225);
nand U13817 (N_13817,N_9294,N_8857);
nor U13818 (N_13818,N_6577,N_7125);
nor U13819 (N_13819,N_9379,N_8508);
nor U13820 (N_13820,N_6970,N_7099);
xor U13821 (N_13821,N_6029,N_9322);
and U13822 (N_13822,N_9634,N_9970);
nand U13823 (N_13823,N_6505,N_9357);
nand U13824 (N_13824,N_8074,N_8721);
or U13825 (N_13825,N_9301,N_6450);
or U13826 (N_13826,N_7942,N_5489);
nor U13827 (N_13827,N_5996,N_6685);
nand U13828 (N_13828,N_8887,N_6149);
nand U13829 (N_13829,N_7701,N_9653);
and U13830 (N_13830,N_9918,N_8715);
and U13831 (N_13831,N_5835,N_8652);
nand U13832 (N_13832,N_8200,N_5220);
nand U13833 (N_13833,N_7664,N_6037);
nand U13834 (N_13834,N_7379,N_6537);
and U13835 (N_13835,N_9426,N_5267);
or U13836 (N_13836,N_7910,N_5860);
and U13837 (N_13837,N_7273,N_7851);
nor U13838 (N_13838,N_8549,N_9163);
nand U13839 (N_13839,N_9345,N_9372);
nor U13840 (N_13840,N_7510,N_6686);
and U13841 (N_13841,N_9126,N_7001);
or U13842 (N_13842,N_6309,N_9172);
or U13843 (N_13843,N_9263,N_8947);
or U13844 (N_13844,N_9824,N_8396);
and U13845 (N_13845,N_7801,N_8091);
nor U13846 (N_13846,N_9440,N_8123);
nand U13847 (N_13847,N_6535,N_6120);
nor U13848 (N_13848,N_5767,N_5290);
and U13849 (N_13849,N_5859,N_7494);
and U13850 (N_13850,N_9796,N_5589);
and U13851 (N_13851,N_5272,N_6857);
xor U13852 (N_13852,N_7564,N_7205);
or U13853 (N_13853,N_6231,N_8285);
nor U13854 (N_13854,N_6748,N_8635);
and U13855 (N_13855,N_7946,N_7387);
nor U13856 (N_13856,N_6607,N_7766);
and U13857 (N_13857,N_6727,N_9020);
nor U13858 (N_13858,N_6351,N_7123);
and U13859 (N_13859,N_8487,N_6153);
and U13860 (N_13860,N_7809,N_8145);
and U13861 (N_13861,N_5951,N_6789);
nor U13862 (N_13862,N_9901,N_6040);
or U13863 (N_13863,N_6185,N_8969);
and U13864 (N_13864,N_7108,N_9788);
nand U13865 (N_13865,N_5943,N_9972);
and U13866 (N_13866,N_9634,N_9218);
nand U13867 (N_13867,N_8058,N_5095);
nor U13868 (N_13868,N_7463,N_9691);
and U13869 (N_13869,N_7652,N_6250);
and U13870 (N_13870,N_5725,N_9768);
nand U13871 (N_13871,N_7830,N_9297);
nand U13872 (N_13872,N_7529,N_8565);
xor U13873 (N_13873,N_5992,N_6678);
or U13874 (N_13874,N_8403,N_8702);
nor U13875 (N_13875,N_8803,N_7520);
and U13876 (N_13876,N_7520,N_9474);
nor U13877 (N_13877,N_6022,N_7772);
nand U13878 (N_13878,N_5163,N_5959);
nor U13879 (N_13879,N_9679,N_5491);
nand U13880 (N_13880,N_6939,N_6986);
nor U13881 (N_13881,N_9063,N_9007);
and U13882 (N_13882,N_5116,N_8898);
nor U13883 (N_13883,N_9186,N_9098);
nand U13884 (N_13884,N_9365,N_7006);
nor U13885 (N_13885,N_7222,N_6574);
nand U13886 (N_13886,N_8202,N_9514);
or U13887 (N_13887,N_5622,N_7765);
or U13888 (N_13888,N_6438,N_9419);
and U13889 (N_13889,N_5144,N_8501);
or U13890 (N_13890,N_9410,N_6299);
and U13891 (N_13891,N_9142,N_9033);
and U13892 (N_13892,N_5935,N_8809);
and U13893 (N_13893,N_9305,N_8681);
or U13894 (N_13894,N_6391,N_6756);
nand U13895 (N_13895,N_5039,N_9733);
nor U13896 (N_13896,N_6884,N_9722);
or U13897 (N_13897,N_5842,N_6689);
nor U13898 (N_13898,N_8230,N_7487);
nand U13899 (N_13899,N_9503,N_5091);
and U13900 (N_13900,N_9311,N_6969);
and U13901 (N_13901,N_8016,N_8780);
nand U13902 (N_13902,N_5192,N_7689);
and U13903 (N_13903,N_6079,N_5278);
or U13904 (N_13904,N_9560,N_5887);
nand U13905 (N_13905,N_6638,N_6017);
nand U13906 (N_13906,N_7795,N_8952);
or U13907 (N_13907,N_8013,N_7188);
and U13908 (N_13908,N_9773,N_9011);
or U13909 (N_13909,N_5570,N_8025);
or U13910 (N_13910,N_9032,N_6465);
nor U13911 (N_13911,N_7378,N_7281);
and U13912 (N_13912,N_5690,N_9886);
and U13913 (N_13913,N_6660,N_6716);
nand U13914 (N_13914,N_5247,N_6967);
nand U13915 (N_13915,N_6941,N_7185);
or U13916 (N_13916,N_6847,N_5263);
nor U13917 (N_13917,N_8116,N_9963);
and U13918 (N_13918,N_9521,N_7913);
nand U13919 (N_13919,N_9872,N_9540);
nand U13920 (N_13920,N_8427,N_5564);
and U13921 (N_13921,N_8462,N_5083);
nand U13922 (N_13922,N_9054,N_7536);
and U13923 (N_13923,N_5782,N_5472);
nor U13924 (N_13924,N_5928,N_9939);
nand U13925 (N_13925,N_7901,N_8174);
or U13926 (N_13926,N_5809,N_6726);
nor U13927 (N_13927,N_8302,N_5484);
and U13928 (N_13928,N_5940,N_7703);
or U13929 (N_13929,N_7532,N_5601);
and U13930 (N_13930,N_7915,N_6156);
and U13931 (N_13931,N_8386,N_9275);
nand U13932 (N_13932,N_6114,N_5819);
nand U13933 (N_13933,N_8698,N_9000);
nand U13934 (N_13934,N_9960,N_5049);
or U13935 (N_13935,N_5442,N_7111);
or U13936 (N_13936,N_5267,N_5283);
nor U13937 (N_13937,N_8417,N_6897);
nand U13938 (N_13938,N_9400,N_5729);
and U13939 (N_13939,N_5241,N_5636);
nor U13940 (N_13940,N_6670,N_8136);
nor U13941 (N_13941,N_9733,N_7210);
or U13942 (N_13942,N_5348,N_7651);
or U13943 (N_13943,N_9617,N_5147);
nor U13944 (N_13944,N_6311,N_6580);
nand U13945 (N_13945,N_7502,N_7820);
nand U13946 (N_13946,N_9010,N_9515);
or U13947 (N_13947,N_5468,N_9650);
or U13948 (N_13948,N_7447,N_6469);
and U13949 (N_13949,N_9115,N_9423);
and U13950 (N_13950,N_9867,N_9712);
or U13951 (N_13951,N_5444,N_9057);
and U13952 (N_13952,N_6881,N_7307);
nand U13953 (N_13953,N_9483,N_6476);
or U13954 (N_13954,N_6847,N_6935);
or U13955 (N_13955,N_7119,N_7852);
and U13956 (N_13956,N_5947,N_8953);
nor U13957 (N_13957,N_9793,N_8440);
and U13958 (N_13958,N_8021,N_7491);
or U13959 (N_13959,N_5347,N_7403);
and U13960 (N_13960,N_5407,N_5037);
nand U13961 (N_13961,N_5611,N_9708);
or U13962 (N_13962,N_6036,N_8067);
xor U13963 (N_13963,N_8129,N_9868);
and U13964 (N_13964,N_8660,N_5764);
nor U13965 (N_13965,N_5530,N_7465);
or U13966 (N_13966,N_6433,N_6813);
nor U13967 (N_13967,N_5284,N_7531);
nor U13968 (N_13968,N_9616,N_8968);
or U13969 (N_13969,N_6317,N_9153);
nand U13970 (N_13970,N_5243,N_9016);
nand U13971 (N_13971,N_5766,N_5497);
xor U13972 (N_13972,N_6202,N_5823);
or U13973 (N_13973,N_6583,N_8452);
nand U13974 (N_13974,N_8281,N_5296);
and U13975 (N_13975,N_5225,N_7092);
nand U13976 (N_13976,N_6067,N_6286);
nor U13977 (N_13977,N_6239,N_9223);
or U13978 (N_13978,N_7003,N_5112);
or U13979 (N_13979,N_5643,N_8261);
and U13980 (N_13980,N_6259,N_8062);
nand U13981 (N_13981,N_8814,N_7667);
nand U13982 (N_13982,N_8587,N_9747);
nand U13983 (N_13983,N_6178,N_6797);
and U13984 (N_13984,N_9560,N_6371);
nand U13985 (N_13985,N_9976,N_7658);
xor U13986 (N_13986,N_5782,N_5415);
and U13987 (N_13987,N_7345,N_5333);
and U13988 (N_13988,N_9473,N_9776);
or U13989 (N_13989,N_6988,N_9240);
or U13990 (N_13990,N_8109,N_9751);
or U13991 (N_13991,N_5733,N_6328);
or U13992 (N_13992,N_8869,N_7093);
or U13993 (N_13993,N_9554,N_9730);
nand U13994 (N_13994,N_7588,N_5696);
and U13995 (N_13995,N_9013,N_8203);
nor U13996 (N_13996,N_6533,N_5504);
nor U13997 (N_13997,N_8508,N_9413);
nand U13998 (N_13998,N_8086,N_7135);
nand U13999 (N_13999,N_7589,N_6800);
nand U14000 (N_14000,N_7438,N_9353);
and U14001 (N_14001,N_6760,N_7177);
or U14002 (N_14002,N_6220,N_9541);
or U14003 (N_14003,N_6556,N_6458);
or U14004 (N_14004,N_8348,N_7546);
xor U14005 (N_14005,N_5626,N_7997);
or U14006 (N_14006,N_6381,N_6352);
xor U14007 (N_14007,N_7422,N_9694);
nand U14008 (N_14008,N_9571,N_6042);
and U14009 (N_14009,N_8480,N_7799);
nand U14010 (N_14010,N_7052,N_9586);
nor U14011 (N_14011,N_8196,N_8752);
nor U14012 (N_14012,N_9824,N_8169);
or U14013 (N_14013,N_9820,N_9893);
or U14014 (N_14014,N_9732,N_9041);
and U14015 (N_14015,N_8262,N_8802);
nand U14016 (N_14016,N_7379,N_9611);
and U14017 (N_14017,N_7141,N_7905);
and U14018 (N_14018,N_7059,N_8768);
nor U14019 (N_14019,N_9882,N_7215);
or U14020 (N_14020,N_7886,N_6678);
or U14021 (N_14021,N_5218,N_7804);
nor U14022 (N_14022,N_5842,N_5832);
or U14023 (N_14023,N_8671,N_7080);
nand U14024 (N_14024,N_6528,N_9039);
nand U14025 (N_14025,N_5647,N_6722);
or U14026 (N_14026,N_6171,N_8622);
and U14027 (N_14027,N_7919,N_5189);
nor U14028 (N_14028,N_9524,N_9319);
and U14029 (N_14029,N_7894,N_8297);
nor U14030 (N_14030,N_9190,N_7608);
nand U14031 (N_14031,N_9248,N_9307);
or U14032 (N_14032,N_7188,N_5285);
nor U14033 (N_14033,N_9698,N_6523);
nand U14034 (N_14034,N_6526,N_8397);
and U14035 (N_14035,N_9390,N_9130);
nand U14036 (N_14036,N_6885,N_9943);
or U14037 (N_14037,N_5958,N_5016);
nor U14038 (N_14038,N_8288,N_6198);
nor U14039 (N_14039,N_7046,N_8078);
and U14040 (N_14040,N_7974,N_7793);
and U14041 (N_14041,N_7327,N_6329);
nand U14042 (N_14042,N_8014,N_9966);
xor U14043 (N_14043,N_7996,N_8505);
nor U14044 (N_14044,N_6312,N_7307);
nor U14045 (N_14045,N_7208,N_9348);
nand U14046 (N_14046,N_5143,N_6976);
or U14047 (N_14047,N_7122,N_5078);
and U14048 (N_14048,N_7752,N_6901);
nor U14049 (N_14049,N_5587,N_6800);
nand U14050 (N_14050,N_7151,N_6059);
or U14051 (N_14051,N_7929,N_8250);
nand U14052 (N_14052,N_9713,N_6900);
and U14053 (N_14053,N_8843,N_6169);
nor U14054 (N_14054,N_5808,N_8792);
nor U14055 (N_14055,N_7644,N_6698);
nor U14056 (N_14056,N_5738,N_6291);
or U14057 (N_14057,N_9123,N_5108);
nand U14058 (N_14058,N_5730,N_8125);
or U14059 (N_14059,N_6355,N_6090);
or U14060 (N_14060,N_7104,N_7216);
or U14061 (N_14061,N_8931,N_9539);
nand U14062 (N_14062,N_7897,N_8451);
and U14063 (N_14063,N_9061,N_6918);
nand U14064 (N_14064,N_6657,N_8119);
nand U14065 (N_14065,N_9238,N_6038);
nand U14066 (N_14066,N_6175,N_5734);
xnor U14067 (N_14067,N_6080,N_8504);
and U14068 (N_14068,N_9384,N_6380);
nand U14069 (N_14069,N_8424,N_8029);
and U14070 (N_14070,N_7860,N_5797);
nand U14071 (N_14071,N_5800,N_5905);
xnor U14072 (N_14072,N_5031,N_8572);
nor U14073 (N_14073,N_5544,N_7336);
and U14074 (N_14074,N_9894,N_6857);
and U14075 (N_14075,N_9627,N_6367);
and U14076 (N_14076,N_7296,N_5141);
nor U14077 (N_14077,N_6746,N_7566);
or U14078 (N_14078,N_7412,N_6190);
nand U14079 (N_14079,N_9242,N_7620);
nand U14080 (N_14080,N_7375,N_8253);
and U14081 (N_14081,N_5976,N_5038);
or U14082 (N_14082,N_9418,N_6339);
nand U14083 (N_14083,N_7869,N_9842);
and U14084 (N_14084,N_8602,N_6234);
nor U14085 (N_14085,N_8857,N_5418);
or U14086 (N_14086,N_6586,N_7586);
nand U14087 (N_14087,N_6088,N_8093);
and U14088 (N_14088,N_6059,N_5967);
or U14089 (N_14089,N_9143,N_8406);
nor U14090 (N_14090,N_7778,N_7035);
or U14091 (N_14091,N_7658,N_8269);
nand U14092 (N_14092,N_9584,N_5259);
or U14093 (N_14093,N_6885,N_7280);
xor U14094 (N_14094,N_8496,N_7474);
and U14095 (N_14095,N_9125,N_9527);
and U14096 (N_14096,N_5034,N_6519);
nor U14097 (N_14097,N_7300,N_5773);
and U14098 (N_14098,N_5510,N_5759);
nor U14099 (N_14099,N_9934,N_7554);
and U14100 (N_14100,N_7538,N_6011);
and U14101 (N_14101,N_9694,N_9089);
nor U14102 (N_14102,N_9244,N_5682);
or U14103 (N_14103,N_6848,N_6946);
and U14104 (N_14104,N_6411,N_8722);
or U14105 (N_14105,N_7050,N_6369);
and U14106 (N_14106,N_9009,N_8363);
nor U14107 (N_14107,N_7700,N_8853);
and U14108 (N_14108,N_5481,N_9189);
or U14109 (N_14109,N_8806,N_6104);
nand U14110 (N_14110,N_9145,N_6451);
nand U14111 (N_14111,N_9269,N_8298);
nand U14112 (N_14112,N_6303,N_7868);
nand U14113 (N_14113,N_7450,N_8330);
or U14114 (N_14114,N_8412,N_7219);
nand U14115 (N_14115,N_7022,N_7070);
nor U14116 (N_14116,N_5877,N_8612);
or U14117 (N_14117,N_6514,N_8683);
nand U14118 (N_14118,N_8880,N_8596);
or U14119 (N_14119,N_9964,N_8893);
and U14120 (N_14120,N_6670,N_7327);
nand U14121 (N_14121,N_5788,N_8457);
nor U14122 (N_14122,N_9566,N_6603);
nand U14123 (N_14123,N_8588,N_8402);
nor U14124 (N_14124,N_7575,N_8108);
nor U14125 (N_14125,N_5721,N_5416);
and U14126 (N_14126,N_5048,N_7011);
and U14127 (N_14127,N_8064,N_8458);
nand U14128 (N_14128,N_6464,N_8775);
and U14129 (N_14129,N_9739,N_6146);
and U14130 (N_14130,N_7572,N_6757);
or U14131 (N_14131,N_8571,N_8132);
nor U14132 (N_14132,N_8690,N_9391);
or U14133 (N_14133,N_7161,N_7749);
and U14134 (N_14134,N_7817,N_5483);
or U14135 (N_14135,N_5660,N_7073);
nand U14136 (N_14136,N_7181,N_9087);
or U14137 (N_14137,N_5195,N_6640);
xnor U14138 (N_14138,N_7676,N_9467);
and U14139 (N_14139,N_8302,N_7946);
or U14140 (N_14140,N_6815,N_5997);
and U14141 (N_14141,N_5006,N_7479);
or U14142 (N_14142,N_9394,N_8217);
nor U14143 (N_14143,N_8517,N_7512);
and U14144 (N_14144,N_8534,N_9678);
nor U14145 (N_14145,N_7468,N_9895);
nand U14146 (N_14146,N_9519,N_6885);
xnor U14147 (N_14147,N_6379,N_6894);
or U14148 (N_14148,N_9334,N_8706);
and U14149 (N_14149,N_6421,N_6307);
nand U14150 (N_14150,N_5385,N_8748);
and U14151 (N_14151,N_6977,N_9596);
nor U14152 (N_14152,N_7848,N_7023);
or U14153 (N_14153,N_7870,N_5239);
and U14154 (N_14154,N_7648,N_9926);
nand U14155 (N_14155,N_5976,N_6093);
or U14156 (N_14156,N_7657,N_9372);
xnor U14157 (N_14157,N_6282,N_6236);
nor U14158 (N_14158,N_7477,N_5795);
nand U14159 (N_14159,N_7901,N_5101);
and U14160 (N_14160,N_9514,N_7514);
nand U14161 (N_14161,N_9986,N_7304);
nor U14162 (N_14162,N_6348,N_5628);
or U14163 (N_14163,N_8295,N_6560);
or U14164 (N_14164,N_6781,N_7666);
and U14165 (N_14165,N_9785,N_9920);
nand U14166 (N_14166,N_9154,N_8904);
nand U14167 (N_14167,N_7253,N_8035);
nor U14168 (N_14168,N_6472,N_7701);
nand U14169 (N_14169,N_9462,N_8929);
nor U14170 (N_14170,N_8465,N_5087);
or U14171 (N_14171,N_6275,N_7106);
or U14172 (N_14172,N_9929,N_9828);
nor U14173 (N_14173,N_8243,N_9209);
nor U14174 (N_14174,N_9013,N_7893);
nor U14175 (N_14175,N_9376,N_5316);
nand U14176 (N_14176,N_9642,N_6797);
nand U14177 (N_14177,N_6985,N_7819);
and U14178 (N_14178,N_7012,N_5995);
or U14179 (N_14179,N_5659,N_7594);
nand U14180 (N_14180,N_8639,N_5867);
or U14181 (N_14181,N_8673,N_8045);
nor U14182 (N_14182,N_8561,N_5145);
and U14183 (N_14183,N_7651,N_5009);
nor U14184 (N_14184,N_9019,N_6229);
and U14185 (N_14185,N_8630,N_7930);
nand U14186 (N_14186,N_9294,N_9414);
nor U14187 (N_14187,N_7387,N_8990);
and U14188 (N_14188,N_8955,N_5997);
or U14189 (N_14189,N_8627,N_8194);
nand U14190 (N_14190,N_8415,N_9962);
nand U14191 (N_14191,N_7603,N_7133);
and U14192 (N_14192,N_8580,N_5759);
nor U14193 (N_14193,N_8138,N_7990);
nor U14194 (N_14194,N_5340,N_9022);
or U14195 (N_14195,N_8001,N_6574);
nand U14196 (N_14196,N_7790,N_9743);
nand U14197 (N_14197,N_7788,N_9205);
nand U14198 (N_14198,N_5937,N_5665);
xnor U14199 (N_14199,N_7229,N_9720);
or U14200 (N_14200,N_9196,N_5423);
and U14201 (N_14201,N_6755,N_8255);
or U14202 (N_14202,N_5807,N_6921);
nand U14203 (N_14203,N_5557,N_8719);
and U14204 (N_14204,N_6674,N_7361);
and U14205 (N_14205,N_5069,N_5674);
xor U14206 (N_14206,N_8773,N_8784);
and U14207 (N_14207,N_6792,N_7183);
or U14208 (N_14208,N_6428,N_8090);
or U14209 (N_14209,N_8125,N_6680);
and U14210 (N_14210,N_9637,N_5983);
and U14211 (N_14211,N_9454,N_6681);
nand U14212 (N_14212,N_5771,N_8069);
nor U14213 (N_14213,N_7116,N_7788);
nor U14214 (N_14214,N_9516,N_6109);
nand U14215 (N_14215,N_8293,N_6815);
nor U14216 (N_14216,N_5430,N_8114);
or U14217 (N_14217,N_7563,N_7499);
nand U14218 (N_14218,N_6562,N_8535);
nor U14219 (N_14219,N_8813,N_7182);
nor U14220 (N_14220,N_8528,N_5848);
or U14221 (N_14221,N_5712,N_9629);
nor U14222 (N_14222,N_7448,N_5663);
nor U14223 (N_14223,N_5916,N_6267);
or U14224 (N_14224,N_8341,N_5137);
nor U14225 (N_14225,N_8194,N_7653);
xnor U14226 (N_14226,N_8188,N_8439);
nor U14227 (N_14227,N_6052,N_7624);
nor U14228 (N_14228,N_5708,N_8389);
nand U14229 (N_14229,N_9778,N_8779);
nor U14230 (N_14230,N_7541,N_9207);
nor U14231 (N_14231,N_9319,N_5233);
or U14232 (N_14232,N_9890,N_6830);
and U14233 (N_14233,N_7381,N_8491);
nor U14234 (N_14234,N_8070,N_7069);
and U14235 (N_14235,N_6451,N_7355);
and U14236 (N_14236,N_6367,N_8928);
nand U14237 (N_14237,N_5833,N_9112);
and U14238 (N_14238,N_9169,N_5462);
and U14239 (N_14239,N_9469,N_6943);
or U14240 (N_14240,N_6955,N_6526);
or U14241 (N_14241,N_5632,N_5025);
nor U14242 (N_14242,N_9309,N_9038);
and U14243 (N_14243,N_7040,N_6532);
nor U14244 (N_14244,N_8420,N_9209);
nor U14245 (N_14245,N_6630,N_5649);
and U14246 (N_14246,N_7976,N_7942);
and U14247 (N_14247,N_5625,N_5415);
or U14248 (N_14248,N_7110,N_9445);
nor U14249 (N_14249,N_9872,N_7628);
or U14250 (N_14250,N_8886,N_9747);
and U14251 (N_14251,N_5632,N_5200);
nor U14252 (N_14252,N_9374,N_8328);
nand U14253 (N_14253,N_8506,N_5456);
nor U14254 (N_14254,N_9314,N_7009);
nor U14255 (N_14255,N_5212,N_6422);
nand U14256 (N_14256,N_7954,N_9283);
and U14257 (N_14257,N_8044,N_8675);
or U14258 (N_14258,N_7150,N_8633);
nor U14259 (N_14259,N_8617,N_6991);
nand U14260 (N_14260,N_8920,N_7559);
and U14261 (N_14261,N_8316,N_6139);
and U14262 (N_14262,N_9090,N_6574);
nor U14263 (N_14263,N_6979,N_6408);
nand U14264 (N_14264,N_7377,N_9473);
or U14265 (N_14265,N_7951,N_9634);
nand U14266 (N_14266,N_8419,N_7928);
xor U14267 (N_14267,N_8687,N_7225);
and U14268 (N_14268,N_5311,N_8419);
nor U14269 (N_14269,N_8440,N_9325);
and U14270 (N_14270,N_5007,N_8739);
or U14271 (N_14271,N_7061,N_5062);
nand U14272 (N_14272,N_7124,N_5897);
or U14273 (N_14273,N_5884,N_5799);
or U14274 (N_14274,N_6808,N_6452);
or U14275 (N_14275,N_6054,N_7964);
nand U14276 (N_14276,N_5128,N_6260);
or U14277 (N_14277,N_5032,N_6491);
or U14278 (N_14278,N_9336,N_6174);
and U14279 (N_14279,N_5569,N_5129);
xor U14280 (N_14280,N_6006,N_5825);
nand U14281 (N_14281,N_6264,N_6046);
and U14282 (N_14282,N_6568,N_8269);
or U14283 (N_14283,N_5698,N_6204);
nand U14284 (N_14284,N_5550,N_7599);
or U14285 (N_14285,N_5103,N_8034);
and U14286 (N_14286,N_8155,N_9571);
nand U14287 (N_14287,N_7405,N_9292);
nand U14288 (N_14288,N_7234,N_9089);
nand U14289 (N_14289,N_8201,N_7963);
or U14290 (N_14290,N_8568,N_6870);
or U14291 (N_14291,N_5209,N_5338);
nand U14292 (N_14292,N_7444,N_5826);
nor U14293 (N_14293,N_9379,N_8016);
and U14294 (N_14294,N_6294,N_6809);
nand U14295 (N_14295,N_9071,N_5107);
nor U14296 (N_14296,N_7672,N_5329);
and U14297 (N_14297,N_5348,N_5337);
nor U14298 (N_14298,N_6758,N_9321);
nand U14299 (N_14299,N_9393,N_7379);
and U14300 (N_14300,N_7323,N_6657);
nand U14301 (N_14301,N_5068,N_7297);
or U14302 (N_14302,N_7713,N_5709);
nor U14303 (N_14303,N_5489,N_8369);
and U14304 (N_14304,N_7720,N_8007);
and U14305 (N_14305,N_6390,N_8900);
nand U14306 (N_14306,N_7253,N_6923);
or U14307 (N_14307,N_8607,N_5821);
and U14308 (N_14308,N_6399,N_7086);
or U14309 (N_14309,N_6507,N_8852);
and U14310 (N_14310,N_5555,N_7046);
and U14311 (N_14311,N_5237,N_6955);
nand U14312 (N_14312,N_7071,N_7441);
nand U14313 (N_14313,N_9320,N_7387);
nor U14314 (N_14314,N_8341,N_8510);
and U14315 (N_14315,N_5309,N_5171);
or U14316 (N_14316,N_9389,N_5339);
and U14317 (N_14317,N_9139,N_7317);
nand U14318 (N_14318,N_6858,N_9614);
or U14319 (N_14319,N_5021,N_6589);
and U14320 (N_14320,N_6541,N_8504);
and U14321 (N_14321,N_9782,N_9158);
xor U14322 (N_14322,N_8645,N_5055);
or U14323 (N_14323,N_8007,N_7342);
nand U14324 (N_14324,N_5470,N_9070);
or U14325 (N_14325,N_8247,N_8695);
nor U14326 (N_14326,N_5554,N_9789);
or U14327 (N_14327,N_9154,N_5867);
or U14328 (N_14328,N_5352,N_5126);
and U14329 (N_14329,N_5793,N_6856);
nand U14330 (N_14330,N_6605,N_9681);
and U14331 (N_14331,N_6128,N_7377);
or U14332 (N_14332,N_5292,N_9145);
nand U14333 (N_14333,N_6911,N_7036);
or U14334 (N_14334,N_9506,N_9389);
nor U14335 (N_14335,N_8843,N_7466);
nor U14336 (N_14336,N_8871,N_5448);
nor U14337 (N_14337,N_6850,N_7145);
nand U14338 (N_14338,N_6855,N_7980);
and U14339 (N_14339,N_8776,N_6222);
or U14340 (N_14340,N_5736,N_9276);
nand U14341 (N_14341,N_5976,N_7232);
nand U14342 (N_14342,N_5690,N_5890);
or U14343 (N_14343,N_6062,N_9218);
nor U14344 (N_14344,N_6043,N_6541);
and U14345 (N_14345,N_5538,N_9880);
or U14346 (N_14346,N_8464,N_6282);
nor U14347 (N_14347,N_5034,N_5493);
xor U14348 (N_14348,N_6524,N_9019);
nor U14349 (N_14349,N_8705,N_7221);
and U14350 (N_14350,N_9813,N_7445);
nor U14351 (N_14351,N_5170,N_6761);
nor U14352 (N_14352,N_8580,N_7332);
xor U14353 (N_14353,N_5115,N_8985);
and U14354 (N_14354,N_8216,N_8023);
nand U14355 (N_14355,N_8039,N_6238);
and U14356 (N_14356,N_9926,N_6906);
nand U14357 (N_14357,N_6995,N_9050);
and U14358 (N_14358,N_6224,N_7587);
nor U14359 (N_14359,N_7493,N_6938);
nand U14360 (N_14360,N_6037,N_9094);
or U14361 (N_14361,N_6060,N_8339);
nand U14362 (N_14362,N_9333,N_6811);
nor U14363 (N_14363,N_9994,N_5132);
nand U14364 (N_14364,N_9342,N_7019);
nor U14365 (N_14365,N_9937,N_6923);
nor U14366 (N_14366,N_7511,N_7229);
nor U14367 (N_14367,N_6843,N_5965);
nand U14368 (N_14368,N_5172,N_6071);
nor U14369 (N_14369,N_6889,N_5198);
and U14370 (N_14370,N_6130,N_8252);
nor U14371 (N_14371,N_5589,N_9549);
and U14372 (N_14372,N_9252,N_9841);
and U14373 (N_14373,N_8203,N_8826);
and U14374 (N_14374,N_9807,N_9751);
nand U14375 (N_14375,N_9947,N_9662);
nand U14376 (N_14376,N_7479,N_9173);
nand U14377 (N_14377,N_8790,N_7769);
and U14378 (N_14378,N_5960,N_6389);
nand U14379 (N_14379,N_6756,N_7301);
or U14380 (N_14380,N_7837,N_8868);
and U14381 (N_14381,N_9345,N_6779);
or U14382 (N_14382,N_5797,N_5128);
nor U14383 (N_14383,N_6472,N_5890);
and U14384 (N_14384,N_8325,N_6344);
nand U14385 (N_14385,N_6315,N_6035);
nor U14386 (N_14386,N_6963,N_6769);
nand U14387 (N_14387,N_6214,N_8463);
nor U14388 (N_14388,N_8935,N_7897);
nor U14389 (N_14389,N_6500,N_6842);
nor U14390 (N_14390,N_8122,N_7054);
nor U14391 (N_14391,N_5718,N_9676);
or U14392 (N_14392,N_9847,N_8110);
nor U14393 (N_14393,N_7127,N_8507);
and U14394 (N_14394,N_5867,N_6546);
and U14395 (N_14395,N_5058,N_5698);
nand U14396 (N_14396,N_7553,N_9775);
and U14397 (N_14397,N_9116,N_9404);
nor U14398 (N_14398,N_9055,N_9433);
nand U14399 (N_14399,N_7815,N_8436);
or U14400 (N_14400,N_7990,N_7693);
and U14401 (N_14401,N_5490,N_9389);
nor U14402 (N_14402,N_7778,N_5876);
and U14403 (N_14403,N_9296,N_8067);
xnor U14404 (N_14404,N_9033,N_5215);
and U14405 (N_14405,N_6662,N_6292);
and U14406 (N_14406,N_7690,N_8320);
and U14407 (N_14407,N_8094,N_7144);
and U14408 (N_14408,N_6005,N_7187);
and U14409 (N_14409,N_5923,N_7445);
nor U14410 (N_14410,N_6030,N_8639);
nand U14411 (N_14411,N_6237,N_7690);
nand U14412 (N_14412,N_6042,N_5101);
and U14413 (N_14413,N_9825,N_6696);
and U14414 (N_14414,N_7534,N_7374);
or U14415 (N_14415,N_5485,N_8439);
or U14416 (N_14416,N_8090,N_6976);
and U14417 (N_14417,N_8372,N_9217);
nor U14418 (N_14418,N_6832,N_7808);
nand U14419 (N_14419,N_5961,N_7988);
and U14420 (N_14420,N_7744,N_7772);
nand U14421 (N_14421,N_6413,N_6547);
xnor U14422 (N_14422,N_6419,N_7492);
or U14423 (N_14423,N_7490,N_9544);
or U14424 (N_14424,N_5159,N_6478);
or U14425 (N_14425,N_8519,N_8965);
nand U14426 (N_14426,N_9775,N_6477);
nand U14427 (N_14427,N_6440,N_9095);
nand U14428 (N_14428,N_7972,N_7713);
xnor U14429 (N_14429,N_6704,N_7278);
or U14430 (N_14430,N_7139,N_8109);
nand U14431 (N_14431,N_5065,N_8483);
nor U14432 (N_14432,N_8548,N_8688);
nand U14433 (N_14433,N_9246,N_8019);
and U14434 (N_14434,N_6778,N_8791);
or U14435 (N_14435,N_7587,N_7692);
and U14436 (N_14436,N_6938,N_5471);
nand U14437 (N_14437,N_7321,N_5934);
nand U14438 (N_14438,N_7204,N_8577);
and U14439 (N_14439,N_6108,N_5242);
xor U14440 (N_14440,N_7512,N_5122);
and U14441 (N_14441,N_5802,N_7476);
and U14442 (N_14442,N_7297,N_6038);
nor U14443 (N_14443,N_8346,N_5000);
nand U14444 (N_14444,N_6422,N_7236);
nand U14445 (N_14445,N_7305,N_9493);
nand U14446 (N_14446,N_9995,N_7163);
and U14447 (N_14447,N_7067,N_9822);
or U14448 (N_14448,N_6429,N_7809);
nor U14449 (N_14449,N_7988,N_6070);
and U14450 (N_14450,N_5219,N_8158);
or U14451 (N_14451,N_7040,N_7218);
and U14452 (N_14452,N_7379,N_6131);
nand U14453 (N_14453,N_9936,N_5927);
or U14454 (N_14454,N_7398,N_5104);
nand U14455 (N_14455,N_5146,N_5236);
and U14456 (N_14456,N_5781,N_5761);
and U14457 (N_14457,N_6450,N_8204);
or U14458 (N_14458,N_6317,N_9261);
nand U14459 (N_14459,N_8528,N_7810);
and U14460 (N_14460,N_5591,N_7588);
nor U14461 (N_14461,N_6913,N_5349);
nor U14462 (N_14462,N_5396,N_7516);
nor U14463 (N_14463,N_6060,N_9667);
and U14464 (N_14464,N_6494,N_5993);
nor U14465 (N_14465,N_9215,N_8972);
nor U14466 (N_14466,N_8173,N_8447);
and U14467 (N_14467,N_7578,N_5883);
nor U14468 (N_14468,N_7488,N_8298);
and U14469 (N_14469,N_8351,N_5648);
xnor U14470 (N_14470,N_8044,N_9986);
and U14471 (N_14471,N_9050,N_7539);
nand U14472 (N_14472,N_9776,N_7881);
nor U14473 (N_14473,N_7845,N_7107);
nor U14474 (N_14474,N_9487,N_9253);
or U14475 (N_14475,N_6806,N_5095);
nand U14476 (N_14476,N_9994,N_8802);
or U14477 (N_14477,N_7941,N_9352);
nor U14478 (N_14478,N_9757,N_7038);
nand U14479 (N_14479,N_5336,N_6814);
nand U14480 (N_14480,N_7849,N_8920);
nand U14481 (N_14481,N_8779,N_7572);
nor U14482 (N_14482,N_9341,N_7384);
nor U14483 (N_14483,N_6807,N_5899);
or U14484 (N_14484,N_9383,N_7967);
or U14485 (N_14485,N_6231,N_9344);
and U14486 (N_14486,N_6074,N_9149);
xnor U14487 (N_14487,N_8748,N_8039);
nor U14488 (N_14488,N_5822,N_6776);
xnor U14489 (N_14489,N_9547,N_7153);
and U14490 (N_14490,N_9307,N_5747);
and U14491 (N_14491,N_5632,N_8654);
nand U14492 (N_14492,N_7113,N_5760);
and U14493 (N_14493,N_6656,N_9396);
nand U14494 (N_14494,N_6800,N_8890);
nand U14495 (N_14495,N_8770,N_5729);
nand U14496 (N_14496,N_6176,N_8191);
nor U14497 (N_14497,N_7116,N_7010);
nor U14498 (N_14498,N_9367,N_6525);
nor U14499 (N_14499,N_6515,N_8887);
or U14500 (N_14500,N_7097,N_8479);
nand U14501 (N_14501,N_8531,N_7490);
nor U14502 (N_14502,N_5967,N_5531);
nor U14503 (N_14503,N_5462,N_7612);
nand U14504 (N_14504,N_8012,N_6669);
and U14505 (N_14505,N_9092,N_5505);
and U14506 (N_14506,N_7229,N_8516);
nor U14507 (N_14507,N_6461,N_6482);
nand U14508 (N_14508,N_5115,N_8424);
and U14509 (N_14509,N_9511,N_9553);
xor U14510 (N_14510,N_9837,N_9243);
and U14511 (N_14511,N_9648,N_8539);
nor U14512 (N_14512,N_5020,N_6396);
or U14513 (N_14513,N_8338,N_8245);
nor U14514 (N_14514,N_6098,N_8581);
or U14515 (N_14515,N_6947,N_8738);
nand U14516 (N_14516,N_7816,N_6746);
nor U14517 (N_14517,N_8195,N_8769);
or U14518 (N_14518,N_9358,N_6569);
nand U14519 (N_14519,N_6332,N_9685);
and U14520 (N_14520,N_8903,N_6439);
and U14521 (N_14521,N_7317,N_8078);
nand U14522 (N_14522,N_5998,N_8137);
nor U14523 (N_14523,N_9199,N_9208);
nor U14524 (N_14524,N_5054,N_9324);
and U14525 (N_14525,N_5724,N_6873);
nor U14526 (N_14526,N_5611,N_5739);
nand U14527 (N_14527,N_7650,N_6840);
nor U14528 (N_14528,N_5385,N_6782);
or U14529 (N_14529,N_5705,N_5709);
and U14530 (N_14530,N_7168,N_6992);
and U14531 (N_14531,N_8347,N_6263);
nor U14532 (N_14532,N_9650,N_7482);
xor U14533 (N_14533,N_9189,N_8208);
or U14534 (N_14534,N_7127,N_7313);
or U14535 (N_14535,N_7866,N_9909);
nand U14536 (N_14536,N_9099,N_9884);
or U14537 (N_14537,N_9074,N_9729);
nor U14538 (N_14538,N_9174,N_6179);
and U14539 (N_14539,N_5200,N_9163);
and U14540 (N_14540,N_5893,N_5772);
or U14541 (N_14541,N_5316,N_8232);
nand U14542 (N_14542,N_9710,N_6404);
and U14543 (N_14543,N_9704,N_5500);
nor U14544 (N_14544,N_7251,N_7066);
nand U14545 (N_14545,N_6665,N_9499);
or U14546 (N_14546,N_5973,N_6644);
nand U14547 (N_14547,N_7255,N_7834);
and U14548 (N_14548,N_7319,N_5761);
and U14549 (N_14549,N_9343,N_6225);
and U14550 (N_14550,N_6245,N_5233);
or U14551 (N_14551,N_7756,N_6430);
or U14552 (N_14552,N_5010,N_5297);
or U14553 (N_14553,N_5102,N_6453);
nor U14554 (N_14554,N_8922,N_6693);
nor U14555 (N_14555,N_6788,N_7851);
and U14556 (N_14556,N_9537,N_9470);
nor U14557 (N_14557,N_7216,N_6969);
and U14558 (N_14558,N_6622,N_7924);
nor U14559 (N_14559,N_9640,N_5859);
or U14560 (N_14560,N_9795,N_9215);
nand U14561 (N_14561,N_6002,N_7352);
nor U14562 (N_14562,N_7653,N_7317);
or U14563 (N_14563,N_6175,N_9862);
nand U14564 (N_14564,N_6077,N_7630);
and U14565 (N_14565,N_6593,N_7429);
or U14566 (N_14566,N_8082,N_8764);
nor U14567 (N_14567,N_7645,N_5210);
and U14568 (N_14568,N_9392,N_8332);
and U14569 (N_14569,N_6686,N_8930);
nand U14570 (N_14570,N_7091,N_5421);
or U14571 (N_14571,N_6570,N_6831);
nand U14572 (N_14572,N_5285,N_6860);
and U14573 (N_14573,N_9705,N_6593);
and U14574 (N_14574,N_7670,N_7614);
nor U14575 (N_14575,N_7681,N_9544);
or U14576 (N_14576,N_7888,N_5551);
nand U14577 (N_14577,N_5911,N_9536);
or U14578 (N_14578,N_5176,N_8128);
and U14579 (N_14579,N_9170,N_8408);
nor U14580 (N_14580,N_5297,N_6109);
nand U14581 (N_14581,N_9729,N_9748);
nor U14582 (N_14582,N_6880,N_7981);
nand U14583 (N_14583,N_6283,N_5259);
or U14584 (N_14584,N_6358,N_6294);
or U14585 (N_14585,N_6739,N_5185);
and U14586 (N_14586,N_9795,N_8210);
nor U14587 (N_14587,N_5933,N_9744);
nor U14588 (N_14588,N_8936,N_5849);
and U14589 (N_14589,N_8555,N_6304);
and U14590 (N_14590,N_6556,N_6433);
and U14591 (N_14591,N_9138,N_6096);
nand U14592 (N_14592,N_9532,N_9024);
or U14593 (N_14593,N_9785,N_8049);
nand U14594 (N_14594,N_8994,N_9273);
nor U14595 (N_14595,N_7467,N_5517);
or U14596 (N_14596,N_9000,N_6503);
or U14597 (N_14597,N_6339,N_7982);
or U14598 (N_14598,N_9756,N_6188);
or U14599 (N_14599,N_6417,N_9804);
nand U14600 (N_14600,N_8328,N_5803);
or U14601 (N_14601,N_8371,N_8128);
nand U14602 (N_14602,N_8848,N_8591);
nand U14603 (N_14603,N_7628,N_5133);
and U14604 (N_14604,N_5198,N_5332);
and U14605 (N_14605,N_9687,N_9542);
nand U14606 (N_14606,N_8482,N_8134);
or U14607 (N_14607,N_6202,N_9519);
or U14608 (N_14608,N_5069,N_8320);
nand U14609 (N_14609,N_8163,N_5120);
nor U14610 (N_14610,N_7320,N_6383);
nor U14611 (N_14611,N_5812,N_5805);
or U14612 (N_14612,N_5898,N_8857);
nand U14613 (N_14613,N_7293,N_7996);
nand U14614 (N_14614,N_6610,N_5854);
and U14615 (N_14615,N_5167,N_8082);
nor U14616 (N_14616,N_8127,N_6080);
nor U14617 (N_14617,N_5182,N_7074);
xor U14618 (N_14618,N_7300,N_6389);
nor U14619 (N_14619,N_7595,N_7079);
nand U14620 (N_14620,N_7485,N_8655);
and U14621 (N_14621,N_8101,N_9538);
and U14622 (N_14622,N_8236,N_9759);
or U14623 (N_14623,N_8001,N_9060);
nand U14624 (N_14624,N_5596,N_5079);
nand U14625 (N_14625,N_5110,N_8802);
xnor U14626 (N_14626,N_6276,N_6927);
nor U14627 (N_14627,N_7151,N_6533);
and U14628 (N_14628,N_6195,N_5021);
or U14629 (N_14629,N_7985,N_6524);
and U14630 (N_14630,N_5864,N_7998);
xor U14631 (N_14631,N_6878,N_7046);
nor U14632 (N_14632,N_9002,N_7830);
xor U14633 (N_14633,N_9405,N_6130);
nor U14634 (N_14634,N_9024,N_7305);
nand U14635 (N_14635,N_9614,N_7493);
and U14636 (N_14636,N_8090,N_7728);
or U14637 (N_14637,N_5747,N_5868);
or U14638 (N_14638,N_7268,N_6632);
and U14639 (N_14639,N_5808,N_8051);
nand U14640 (N_14640,N_8042,N_7473);
and U14641 (N_14641,N_6608,N_8624);
nor U14642 (N_14642,N_9305,N_8214);
or U14643 (N_14643,N_6029,N_8210);
nor U14644 (N_14644,N_8925,N_6208);
or U14645 (N_14645,N_9734,N_7918);
nor U14646 (N_14646,N_7521,N_6822);
and U14647 (N_14647,N_8468,N_5188);
nor U14648 (N_14648,N_6984,N_6747);
and U14649 (N_14649,N_7379,N_5040);
or U14650 (N_14650,N_7954,N_7702);
xor U14651 (N_14651,N_7464,N_6054);
and U14652 (N_14652,N_9575,N_8969);
and U14653 (N_14653,N_7267,N_9053);
nand U14654 (N_14654,N_5702,N_7200);
and U14655 (N_14655,N_5579,N_6169);
and U14656 (N_14656,N_5972,N_5499);
or U14657 (N_14657,N_7080,N_5092);
and U14658 (N_14658,N_8547,N_7733);
nor U14659 (N_14659,N_9656,N_6266);
xor U14660 (N_14660,N_7767,N_5940);
and U14661 (N_14661,N_8676,N_9774);
nand U14662 (N_14662,N_6497,N_9578);
nand U14663 (N_14663,N_8367,N_5495);
and U14664 (N_14664,N_5284,N_8748);
nor U14665 (N_14665,N_9872,N_7368);
and U14666 (N_14666,N_7718,N_8161);
nor U14667 (N_14667,N_8908,N_5021);
nor U14668 (N_14668,N_5999,N_9807);
and U14669 (N_14669,N_6594,N_6656);
or U14670 (N_14670,N_5389,N_6735);
or U14671 (N_14671,N_5686,N_6686);
and U14672 (N_14672,N_6182,N_8766);
and U14673 (N_14673,N_9035,N_6866);
nor U14674 (N_14674,N_6860,N_5089);
nor U14675 (N_14675,N_5558,N_7592);
nand U14676 (N_14676,N_6351,N_8142);
or U14677 (N_14677,N_9310,N_8752);
nor U14678 (N_14678,N_9574,N_8930);
and U14679 (N_14679,N_9140,N_7851);
nor U14680 (N_14680,N_9013,N_5697);
and U14681 (N_14681,N_8723,N_9219);
nand U14682 (N_14682,N_6581,N_8015);
or U14683 (N_14683,N_9718,N_9536);
or U14684 (N_14684,N_6249,N_5031);
nor U14685 (N_14685,N_7582,N_6154);
nand U14686 (N_14686,N_6604,N_8013);
and U14687 (N_14687,N_6198,N_7073);
or U14688 (N_14688,N_7053,N_5230);
or U14689 (N_14689,N_6487,N_7481);
or U14690 (N_14690,N_5524,N_7291);
and U14691 (N_14691,N_6477,N_5756);
and U14692 (N_14692,N_8828,N_6946);
and U14693 (N_14693,N_9270,N_6209);
or U14694 (N_14694,N_9403,N_8931);
or U14695 (N_14695,N_6518,N_8374);
or U14696 (N_14696,N_9743,N_7496);
nor U14697 (N_14697,N_7832,N_6384);
and U14698 (N_14698,N_5413,N_7115);
or U14699 (N_14699,N_9314,N_9471);
nand U14700 (N_14700,N_8931,N_8999);
and U14701 (N_14701,N_8635,N_6868);
nand U14702 (N_14702,N_7493,N_8593);
nor U14703 (N_14703,N_7479,N_9777);
nand U14704 (N_14704,N_6063,N_7480);
or U14705 (N_14705,N_5590,N_7892);
nand U14706 (N_14706,N_6529,N_8526);
and U14707 (N_14707,N_5229,N_7034);
xnor U14708 (N_14708,N_8267,N_5661);
nand U14709 (N_14709,N_5357,N_6252);
and U14710 (N_14710,N_7904,N_6411);
nor U14711 (N_14711,N_7136,N_9571);
nand U14712 (N_14712,N_5753,N_9483);
and U14713 (N_14713,N_8214,N_6906);
nor U14714 (N_14714,N_6878,N_5528);
nand U14715 (N_14715,N_5525,N_5302);
or U14716 (N_14716,N_8191,N_9445);
nor U14717 (N_14717,N_7405,N_6009);
and U14718 (N_14718,N_5594,N_5827);
and U14719 (N_14719,N_5722,N_7598);
nor U14720 (N_14720,N_7089,N_6854);
nand U14721 (N_14721,N_6556,N_6235);
nand U14722 (N_14722,N_9711,N_7975);
nor U14723 (N_14723,N_6832,N_7984);
nor U14724 (N_14724,N_6126,N_5811);
nor U14725 (N_14725,N_6676,N_7414);
nand U14726 (N_14726,N_9610,N_7693);
or U14727 (N_14727,N_7917,N_8293);
and U14728 (N_14728,N_8703,N_9771);
and U14729 (N_14729,N_7583,N_6988);
and U14730 (N_14730,N_9430,N_7744);
and U14731 (N_14731,N_8727,N_8535);
nor U14732 (N_14732,N_9615,N_7010);
nor U14733 (N_14733,N_9933,N_7051);
nand U14734 (N_14734,N_9797,N_8322);
and U14735 (N_14735,N_9917,N_7540);
nand U14736 (N_14736,N_9406,N_8221);
and U14737 (N_14737,N_8716,N_9923);
or U14738 (N_14738,N_6412,N_8885);
nand U14739 (N_14739,N_5734,N_5685);
nand U14740 (N_14740,N_7916,N_9706);
nand U14741 (N_14741,N_9980,N_9973);
or U14742 (N_14742,N_9016,N_8540);
nor U14743 (N_14743,N_6787,N_5063);
nand U14744 (N_14744,N_6769,N_5932);
or U14745 (N_14745,N_9440,N_6136);
nand U14746 (N_14746,N_7845,N_6734);
or U14747 (N_14747,N_6241,N_7428);
nor U14748 (N_14748,N_8472,N_7927);
and U14749 (N_14749,N_9509,N_8195);
nor U14750 (N_14750,N_5347,N_5443);
nand U14751 (N_14751,N_6541,N_9028);
nand U14752 (N_14752,N_6925,N_7340);
nor U14753 (N_14753,N_6550,N_9042);
and U14754 (N_14754,N_9067,N_8226);
nand U14755 (N_14755,N_5488,N_6961);
nor U14756 (N_14756,N_5406,N_8452);
nor U14757 (N_14757,N_8499,N_5893);
or U14758 (N_14758,N_6124,N_6966);
xnor U14759 (N_14759,N_7480,N_8100);
nor U14760 (N_14760,N_6057,N_6088);
and U14761 (N_14761,N_6875,N_5082);
nor U14762 (N_14762,N_9146,N_5882);
nor U14763 (N_14763,N_5754,N_7754);
and U14764 (N_14764,N_6136,N_5410);
and U14765 (N_14765,N_9476,N_5010);
or U14766 (N_14766,N_9333,N_9484);
or U14767 (N_14767,N_8449,N_7527);
nor U14768 (N_14768,N_9218,N_7063);
or U14769 (N_14769,N_8038,N_5124);
xnor U14770 (N_14770,N_6869,N_5085);
or U14771 (N_14771,N_6989,N_6416);
nand U14772 (N_14772,N_7620,N_8981);
nand U14773 (N_14773,N_6285,N_6266);
nand U14774 (N_14774,N_7954,N_8109);
or U14775 (N_14775,N_7357,N_9172);
and U14776 (N_14776,N_5752,N_8316);
and U14777 (N_14777,N_7551,N_5278);
nand U14778 (N_14778,N_6342,N_8489);
nand U14779 (N_14779,N_6191,N_9626);
or U14780 (N_14780,N_6561,N_6693);
or U14781 (N_14781,N_5602,N_8264);
or U14782 (N_14782,N_8414,N_9909);
nand U14783 (N_14783,N_9766,N_5620);
nor U14784 (N_14784,N_6941,N_6079);
or U14785 (N_14785,N_6621,N_8363);
and U14786 (N_14786,N_6078,N_5141);
nand U14787 (N_14787,N_6057,N_6547);
or U14788 (N_14788,N_8273,N_5627);
nor U14789 (N_14789,N_5738,N_5226);
nand U14790 (N_14790,N_8891,N_9208);
or U14791 (N_14791,N_8257,N_9814);
and U14792 (N_14792,N_9659,N_7295);
nand U14793 (N_14793,N_7946,N_7242);
nand U14794 (N_14794,N_6574,N_5870);
and U14795 (N_14795,N_6728,N_8971);
nor U14796 (N_14796,N_8503,N_9022);
nand U14797 (N_14797,N_8513,N_7208);
nor U14798 (N_14798,N_8453,N_9247);
and U14799 (N_14799,N_9477,N_5818);
and U14800 (N_14800,N_7006,N_7313);
nor U14801 (N_14801,N_6924,N_9915);
and U14802 (N_14802,N_5258,N_5335);
nand U14803 (N_14803,N_5253,N_9528);
and U14804 (N_14804,N_5124,N_5462);
nand U14805 (N_14805,N_7571,N_8447);
nand U14806 (N_14806,N_5795,N_8968);
nand U14807 (N_14807,N_6966,N_5236);
nand U14808 (N_14808,N_9178,N_6057);
or U14809 (N_14809,N_7620,N_6770);
and U14810 (N_14810,N_8052,N_7757);
nand U14811 (N_14811,N_8147,N_9794);
or U14812 (N_14812,N_5133,N_7460);
nand U14813 (N_14813,N_8158,N_8272);
nand U14814 (N_14814,N_9142,N_7885);
or U14815 (N_14815,N_5039,N_5638);
nand U14816 (N_14816,N_6126,N_9451);
nand U14817 (N_14817,N_6579,N_8535);
nand U14818 (N_14818,N_8310,N_6220);
or U14819 (N_14819,N_6296,N_5704);
xnor U14820 (N_14820,N_8691,N_5368);
and U14821 (N_14821,N_8436,N_7154);
nor U14822 (N_14822,N_6171,N_5975);
nand U14823 (N_14823,N_8335,N_6772);
and U14824 (N_14824,N_5778,N_8543);
nor U14825 (N_14825,N_7189,N_7989);
nor U14826 (N_14826,N_6533,N_6867);
or U14827 (N_14827,N_7647,N_9921);
or U14828 (N_14828,N_5685,N_8821);
or U14829 (N_14829,N_7525,N_6773);
xnor U14830 (N_14830,N_6904,N_8427);
and U14831 (N_14831,N_7322,N_7210);
nor U14832 (N_14832,N_6079,N_9945);
nand U14833 (N_14833,N_7947,N_5544);
or U14834 (N_14834,N_7383,N_6526);
nand U14835 (N_14835,N_8139,N_8296);
or U14836 (N_14836,N_6067,N_9100);
and U14837 (N_14837,N_8914,N_7156);
nand U14838 (N_14838,N_8302,N_8994);
and U14839 (N_14839,N_9347,N_5835);
and U14840 (N_14840,N_5663,N_6645);
and U14841 (N_14841,N_9095,N_5472);
nand U14842 (N_14842,N_6184,N_6796);
nor U14843 (N_14843,N_9715,N_9025);
and U14844 (N_14844,N_7222,N_7332);
or U14845 (N_14845,N_6022,N_8496);
nor U14846 (N_14846,N_5947,N_6544);
and U14847 (N_14847,N_7327,N_9017);
nand U14848 (N_14848,N_5114,N_5469);
or U14849 (N_14849,N_6428,N_5181);
nor U14850 (N_14850,N_6710,N_5951);
nor U14851 (N_14851,N_8090,N_5696);
or U14852 (N_14852,N_7294,N_7766);
or U14853 (N_14853,N_8708,N_8166);
or U14854 (N_14854,N_6753,N_5933);
nor U14855 (N_14855,N_5781,N_9424);
and U14856 (N_14856,N_5793,N_7949);
and U14857 (N_14857,N_9789,N_7083);
xor U14858 (N_14858,N_8374,N_5213);
and U14859 (N_14859,N_6764,N_5665);
or U14860 (N_14860,N_8230,N_7942);
nand U14861 (N_14861,N_8416,N_6103);
nor U14862 (N_14862,N_5887,N_7423);
or U14863 (N_14863,N_5814,N_9981);
nand U14864 (N_14864,N_8433,N_5621);
or U14865 (N_14865,N_5537,N_5077);
and U14866 (N_14866,N_8289,N_7577);
or U14867 (N_14867,N_8973,N_7370);
and U14868 (N_14868,N_7278,N_7661);
nor U14869 (N_14869,N_7568,N_8434);
nand U14870 (N_14870,N_8191,N_9966);
nor U14871 (N_14871,N_6836,N_6288);
nor U14872 (N_14872,N_9129,N_9194);
and U14873 (N_14873,N_9450,N_9654);
nand U14874 (N_14874,N_8976,N_7596);
or U14875 (N_14875,N_8907,N_7908);
nand U14876 (N_14876,N_9144,N_9243);
and U14877 (N_14877,N_8415,N_8372);
and U14878 (N_14878,N_6129,N_9312);
or U14879 (N_14879,N_8237,N_5837);
nand U14880 (N_14880,N_7847,N_5092);
nor U14881 (N_14881,N_6316,N_7854);
or U14882 (N_14882,N_9521,N_6544);
nor U14883 (N_14883,N_5550,N_5369);
or U14884 (N_14884,N_9512,N_5129);
nand U14885 (N_14885,N_6984,N_8189);
or U14886 (N_14886,N_8846,N_8921);
nor U14887 (N_14887,N_5971,N_8285);
nand U14888 (N_14888,N_7462,N_5489);
or U14889 (N_14889,N_6874,N_9175);
nor U14890 (N_14890,N_8112,N_7799);
and U14891 (N_14891,N_5336,N_7804);
xnor U14892 (N_14892,N_6996,N_8425);
and U14893 (N_14893,N_9005,N_8980);
nor U14894 (N_14894,N_6041,N_9325);
or U14895 (N_14895,N_8782,N_8911);
nor U14896 (N_14896,N_9727,N_6683);
nand U14897 (N_14897,N_6519,N_9011);
xor U14898 (N_14898,N_8542,N_5899);
and U14899 (N_14899,N_8618,N_5014);
nor U14900 (N_14900,N_9901,N_8534);
nor U14901 (N_14901,N_9126,N_7284);
nor U14902 (N_14902,N_7143,N_8385);
nand U14903 (N_14903,N_6319,N_9053);
nand U14904 (N_14904,N_9720,N_9029);
and U14905 (N_14905,N_7096,N_7931);
and U14906 (N_14906,N_9702,N_7042);
nand U14907 (N_14907,N_8963,N_5430);
nor U14908 (N_14908,N_8191,N_6154);
and U14909 (N_14909,N_5014,N_8678);
or U14910 (N_14910,N_9913,N_6789);
nor U14911 (N_14911,N_8728,N_9235);
and U14912 (N_14912,N_8208,N_8561);
or U14913 (N_14913,N_6139,N_7111);
nand U14914 (N_14914,N_5091,N_9404);
nand U14915 (N_14915,N_9343,N_5212);
nor U14916 (N_14916,N_9495,N_8160);
and U14917 (N_14917,N_9104,N_8335);
nand U14918 (N_14918,N_6167,N_7797);
nand U14919 (N_14919,N_9594,N_5886);
or U14920 (N_14920,N_5592,N_7261);
and U14921 (N_14921,N_7950,N_6770);
nand U14922 (N_14922,N_8021,N_9974);
or U14923 (N_14923,N_6564,N_6194);
or U14924 (N_14924,N_8328,N_8597);
and U14925 (N_14925,N_9721,N_9481);
and U14926 (N_14926,N_5536,N_9020);
nand U14927 (N_14927,N_7155,N_6484);
or U14928 (N_14928,N_7920,N_8305);
or U14929 (N_14929,N_8925,N_8859);
and U14930 (N_14930,N_8728,N_9484);
nand U14931 (N_14931,N_9801,N_9905);
nor U14932 (N_14932,N_6458,N_7110);
or U14933 (N_14933,N_6364,N_8179);
and U14934 (N_14934,N_6164,N_9537);
nor U14935 (N_14935,N_9245,N_7408);
and U14936 (N_14936,N_6824,N_5557);
and U14937 (N_14937,N_7097,N_5738);
nand U14938 (N_14938,N_8948,N_9786);
nor U14939 (N_14939,N_8880,N_9915);
and U14940 (N_14940,N_5750,N_8273);
or U14941 (N_14941,N_5915,N_8886);
or U14942 (N_14942,N_6000,N_7037);
and U14943 (N_14943,N_6241,N_8362);
or U14944 (N_14944,N_6943,N_8260);
nand U14945 (N_14945,N_8273,N_6701);
nand U14946 (N_14946,N_9894,N_5126);
and U14947 (N_14947,N_8561,N_5517);
or U14948 (N_14948,N_7970,N_7139);
or U14949 (N_14949,N_9979,N_7893);
and U14950 (N_14950,N_8606,N_5582);
or U14951 (N_14951,N_9989,N_8237);
nor U14952 (N_14952,N_8692,N_6482);
nor U14953 (N_14953,N_8305,N_6361);
nand U14954 (N_14954,N_6351,N_9505);
and U14955 (N_14955,N_6375,N_7240);
nor U14956 (N_14956,N_9084,N_5170);
nor U14957 (N_14957,N_6902,N_7261);
and U14958 (N_14958,N_9918,N_9349);
and U14959 (N_14959,N_9894,N_9759);
nor U14960 (N_14960,N_6501,N_5048);
or U14961 (N_14961,N_7862,N_8563);
and U14962 (N_14962,N_9023,N_6594);
xor U14963 (N_14963,N_6177,N_6775);
and U14964 (N_14964,N_8576,N_7875);
and U14965 (N_14965,N_6892,N_8407);
nor U14966 (N_14966,N_7338,N_8380);
and U14967 (N_14967,N_6630,N_6859);
or U14968 (N_14968,N_7714,N_9315);
nor U14969 (N_14969,N_5187,N_6268);
or U14970 (N_14970,N_8417,N_5683);
and U14971 (N_14971,N_9130,N_7136);
or U14972 (N_14972,N_8183,N_9240);
and U14973 (N_14973,N_5370,N_7739);
or U14974 (N_14974,N_6458,N_5209);
nor U14975 (N_14975,N_5422,N_9899);
nor U14976 (N_14976,N_6128,N_7562);
nor U14977 (N_14977,N_6821,N_7564);
nand U14978 (N_14978,N_9053,N_7629);
nand U14979 (N_14979,N_5411,N_6851);
nand U14980 (N_14980,N_8684,N_9326);
nor U14981 (N_14981,N_5646,N_9556);
nor U14982 (N_14982,N_7426,N_5234);
or U14983 (N_14983,N_9068,N_6194);
nor U14984 (N_14984,N_6448,N_8238);
or U14985 (N_14985,N_6194,N_8942);
or U14986 (N_14986,N_8877,N_7852);
and U14987 (N_14987,N_7624,N_9586);
nand U14988 (N_14988,N_6161,N_8524);
or U14989 (N_14989,N_8939,N_9357);
nor U14990 (N_14990,N_8085,N_8695);
nand U14991 (N_14991,N_7580,N_9452);
and U14992 (N_14992,N_7826,N_6730);
or U14993 (N_14993,N_8667,N_5344);
nand U14994 (N_14994,N_5443,N_9867);
and U14995 (N_14995,N_6641,N_7615);
nor U14996 (N_14996,N_7198,N_8201);
and U14997 (N_14997,N_6478,N_7576);
or U14998 (N_14998,N_8433,N_6241);
nand U14999 (N_14999,N_8974,N_7182);
nand U15000 (N_15000,N_12635,N_10026);
nand U15001 (N_15001,N_12092,N_12249);
xor U15002 (N_15002,N_10937,N_14547);
and U15003 (N_15003,N_10404,N_13268);
nor U15004 (N_15004,N_12382,N_11839);
nor U15005 (N_15005,N_11474,N_12825);
nor U15006 (N_15006,N_14789,N_10706);
nor U15007 (N_15007,N_10731,N_14209);
nand U15008 (N_15008,N_10364,N_10194);
and U15009 (N_15009,N_10532,N_14368);
and U15010 (N_15010,N_11284,N_11954);
and U15011 (N_15011,N_12811,N_10492);
nor U15012 (N_15012,N_10565,N_13709);
nand U15013 (N_15013,N_12498,N_10462);
or U15014 (N_15014,N_10338,N_13938);
and U15015 (N_15015,N_13075,N_14298);
nand U15016 (N_15016,N_12908,N_13808);
and U15017 (N_15017,N_10711,N_14441);
nand U15018 (N_15018,N_14664,N_12844);
nand U15019 (N_15019,N_10129,N_10155);
nor U15020 (N_15020,N_10389,N_13291);
and U15021 (N_15021,N_12982,N_10999);
and U15022 (N_15022,N_12898,N_13362);
or U15023 (N_15023,N_13302,N_13880);
and U15024 (N_15024,N_14573,N_14217);
nor U15025 (N_15025,N_12333,N_14267);
nand U15026 (N_15026,N_14606,N_10045);
nor U15027 (N_15027,N_10961,N_11554);
nor U15028 (N_15028,N_12262,N_10967);
nand U15029 (N_15029,N_14629,N_11236);
nand U15030 (N_15030,N_10454,N_14948);
and U15031 (N_15031,N_11462,N_12461);
nor U15032 (N_15032,N_10801,N_10883);
and U15033 (N_15033,N_10333,N_13231);
nand U15034 (N_15034,N_13345,N_11705);
and U15035 (N_15035,N_12253,N_11750);
and U15036 (N_15036,N_13108,N_12732);
nor U15037 (N_15037,N_12667,N_11257);
and U15038 (N_15038,N_10366,N_14266);
or U15039 (N_15039,N_12234,N_10311);
nand U15040 (N_15040,N_11953,N_13083);
nand U15041 (N_15041,N_13181,N_14875);
nand U15042 (N_15042,N_10931,N_13884);
and U15043 (N_15043,N_12912,N_13007);
and U15044 (N_15044,N_12703,N_10522);
or U15045 (N_15045,N_11487,N_10924);
nand U15046 (N_15046,N_12455,N_10715);
and U15047 (N_15047,N_13626,N_13816);
or U15048 (N_15048,N_10166,N_13650);
or U15049 (N_15049,N_14213,N_13629);
nor U15050 (N_15050,N_14846,N_13276);
nand U15051 (N_15051,N_10187,N_10641);
and U15052 (N_15052,N_14869,N_14491);
and U15053 (N_15053,N_13900,N_10341);
xnor U15054 (N_15054,N_12040,N_14968);
nand U15055 (N_15055,N_14139,N_11547);
or U15056 (N_15056,N_12583,N_14633);
nor U15057 (N_15057,N_10470,N_11024);
nor U15058 (N_15058,N_11090,N_11282);
nand U15059 (N_15059,N_13842,N_12189);
nand U15060 (N_15060,N_10132,N_14103);
or U15061 (N_15061,N_12311,N_12185);
nor U15062 (N_15062,N_11218,N_14147);
nor U15063 (N_15063,N_13397,N_12926);
nand U15064 (N_15064,N_13682,N_13811);
and U15065 (N_15065,N_14660,N_14177);
and U15066 (N_15066,N_11849,N_13680);
or U15067 (N_15067,N_12218,N_13801);
nand U15068 (N_15068,N_14541,N_14167);
or U15069 (N_15069,N_14513,N_14277);
nand U15070 (N_15070,N_11845,N_14210);
or U15071 (N_15071,N_12839,N_12107);
nand U15072 (N_15072,N_13215,N_12959);
and U15073 (N_15073,N_12695,N_12188);
nand U15074 (N_15074,N_10870,N_12889);
or U15075 (N_15075,N_13175,N_10727);
or U15076 (N_15076,N_11007,N_10951);
or U15077 (N_15077,N_14165,N_12699);
nand U15078 (N_15078,N_11737,N_11773);
or U15079 (N_15079,N_11740,N_11144);
or U15080 (N_15080,N_14745,N_10992);
and U15081 (N_15081,N_12822,N_12377);
or U15082 (N_15082,N_12213,N_12660);
xor U15083 (N_15083,N_13935,N_13590);
nor U15084 (N_15084,N_11341,N_13122);
and U15085 (N_15085,N_12832,N_14042);
or U15086 (N_15086,N_12404,N_11334);
or U15087 (N_15087,N_12722,N_11729);
and U15088 (N_15088,N_14688,N_12228);
or U15089 (N_15089,N_12401,N_13723);
and U15090 (N_15090,N_13343,N_10893);
and U15091 (N_15091,N_13594,N_12038);
nand U15092 (N_15092,N_13352,N_13470);
or U15093 (N_15093,N_13167,N_14215);
or U15094 (N_15094,N_13687,N_11806);
or U15095 (N_15095,N_12309,N_11053);
nor U15096 (N_15096,N_11030,N_11461);
or U15097 (N_15097,N_11939,N_12584);
and U15098 (N_15098,N_14507,N_13125);
nor U15099 (N_15099,N_12998,N_12101);
and U15100 (N_15100,N_10230,N_13556);
or U15101 (N_15101,N_13263,N_13545);
nand U15102 (N_15102,N_11891,N_13966);
and U15103 (N_15103,N_13156,N_14456);
nand U15104 (N_15104,N_13320,N_10013);
xor U15105 (N_15105,N_12108,N_10545);
or U15106 (N_15106,N_14559,N_10971);
nand U15107 (N_15107,N_14062,N_14918);
nand U15108 (N_15108,N_14889,N_12577);
and U15109 (N_15109,N_11320,N_10347);
nor U15110 (N_15110,N_10424,N_10786);
nor U15111 (N_15111,N_12638,N_12353);
nor U15112 (N_15112,N_11790,N_13241);
or U15113 (N_15113,N_10472,N_14973);
nor U15114 (N_15114,N_14160,N_14767);
or U15115 (N_15115,N_11924,N_13359);
or U15116 (N_15116,N_12741,N_13867);
nor U15117 (N_15117,N_13930,N_11751);
or U15118 (N_15118,N_14785,N_11615);
or U15119 (N_15119,N_12184,N_10344);
and U15120 (N_15120,N_13432,N_10688);
nor U15121 (N_15121,N_12385,N_10741);
nand U15122 (N_15122,N_14098,N_14954);
or U15123 (N_15123,N_11078,N_12015);
nand U15124 (N_15124,N_14976,N_11039);
nand U15125 (N_15125,N_13897,N_10824);
nor U15126 (N_15126,N_11532,N_10509);
nand U15127 (N_15127,N_10131,N_10853);
or U15128 (N_15128,N_11361,N_14627);
and U15129 (N_15129,N_13465,N_11522);
nor U15130 (N_15130,N_10310,N_13149);
or U15131 (N_15131,N_11324,N_11048);
and U15132 (N_15132,N_10676,N_11111);
nand U15133 (N_15133,N_11108,N_12677);
and U15134 (N_15134,N_11811,N_13737);
nand U15135 (N_15135,N_14933,N_12933);
nand U15136 (N_15136,N_10257,N_12486);
and U15137 (N_15137,N_12663,N_13858);
nor U15138 (N_15138,N_14342,N_14109);
or U15139 (N_15139,N_13982,N_12025);
or U15140 (N_15140,N_13970,N_10038);
nand U15141 (N_15141,N_10319,N_12984);
nor U15142 (N_15142,N_14190,N_13610);
and U15143 (N_15143,N_14157,N_10001);
or U15144 (N_15144,N_10839,N_13441);
and U15145 (N_15145,N_10516,N_11372);
and U15146 (N_15146,N_11204,N_13752);
nor U15147 (N_15147,N_12975,N_14930);
or U15148 (N_15148,N_13730,N_11465);
nor U15149 (N_15149,N_10638,N_12049);
or U15150 (N_15150,N_10667,N_13036);
nand U15151 (N_15151,N_14646,N_14991);
nor U15152 (N_15152,N_10467,N_13177);
or U15153 (N_15153,N_10864,N_13163);
nor U15154 (N_15154,N_14877,N_13492);
and U15155 (N_15155,N_12402,N_14686);
and U15156 (N_15156,N_14383,N_13455);
or U15157 (N_15157,N_12095,N_11906);
or U15158 (N_15158,N_13541,N_11416);
or U15159 (N_15159,N_10655,N_11092);
nand U15160 (N_15160,N_10037,N_13836);
and U15161 (N_15161,N_11645,N_12626);
and U15162 (N_15162,N_10499,N_13666);
nand U15163 (N_15163,N_10498,N_13478);
or U15164 (N_15164,N_13503,N_12182);
and U15165 (N_15165,N_11943,N_13032);
and U15166 (N_15166,N_11743,N_13479);
nor U15167 (N_15167,N_12103,N_11096);
or U15168 (N_15168,N_13734,N_10019);
nor U15169 (N_15169,N_10184,N_12211);
nor U15170 (N_15170,N_14700,N_11023);
nand U15171 (N_15171,N_11703,N_13347);
and U15172 (N_15172,N_10790,N_10325);
xnor U15173 (N_15173,N_14706,N_11022);
nor U15174 (N_15174,N_14926,N_10416);
or U15175 (N_15175,N_10584,N_13293);
nor U15176 (N_15176,N_14450,N_11802);
and U15177 (N_15177,N_14347,N_12750);
nor U15178 (N_15178,N_14561,N_12821);
nor U15179 (N_15179,N_14415,N_13823);
and U15180 (N_15180,N_10530,N_13550);
nand U15181 (N_15181,N_13238,N_13950);
nor U15182 (N_15182,N_13513,N_13846);
or U15183 (N_15183,N_12160,N_11499);
nand U15184 (N_15184,N_13148,N_12089);
nand U15185 (N_15185,N_11033,N_11794);
or U15186 (N_15186,N_11951,N_10866);
and U15187 (N_15187,N_14044,N_12227);
or U15188 (N_15188,N_14678,N_14421);
nor U15189 (N_15189,N_14356,N_14416);
nor U15190 (N_15190,N_14986,N_12425);
or U15191 (N_15191,N_11398,N_11647);
and U15192 (N_15192,N_12481,N_13374);
nand U15193 (N_15193,N_10585,N_11037);
nor U15194 (N_15194,N_13979,N_13851);
nand U15195 (N_15195,N_13059,N_13250);
nand U15196 (N_15196,N_14278,N_11159);
and U15197 (N_15197,N_10703,N_14281);
nor U15198 (N_15198,N_12444,N_14265);
nand U15199 (N_15199,N_10953,N_13143);
and U15200 (N_15200,N_14680,N_11337);
or U15201 (N_15201,N_13439,N_14837);
or U15202 (N_15202,N_12911,N_10996);
and U15203 (N_15203,N_12603,N_13894);
and U15204 (N_15204,N_11259,N_11103);
or U15205 (N_15205,N_13121,N_13365);
nor U15206 (N_15206,N_11805,N_12562);
nor U15207 (N_15207,N_11525,N_12712);
and U15208 (N_15208,N_12494,N_11363);
nor U15209 (N_15209,N_12701,N_13022);
xor U15210 (N_15210,N_13314,N_10009);
or U15211 (N_15211,N_12893,N_13693);
and U15212 (N_15212,N_12798,N_13297);
or U15213 (N_15213,N_10494,N_10557);
nor U15214 (N_15214,N_14114,N_14064);
nand U15215 (N_15215,N_10978,N_14398);
nand U15216 (N_15216,N_12717,N_14835);
and U15217 (N_15217,N_10117,N_10141);
nor U15218 (N_15218,N_12022,N_13614);
or U15219 (N_15219,N_14553,N_10308);
nand U15220 (N_15220,N_10253,N_10966);
nand U15221 (N_15221,N_11399,N_10005);
nand U15222 (N_15222,N_12432,N_11911);
nor U15223 (N_15223,N_14304,N_11779);
nand U15224 (N_15224,N_10980,N_13561);
and U15225 (N_15225,N_11829,N_13778);
or U15226 (N_15226,N_10204,N_12743);
nand U15227 (N_15227,N_14740,N_14539);
or U15228 (N_15228,N_11093,N_12295);
nor U15229 (N_15229,N_14748,N_13791);
nor U15230 (N_15230,N_10597,N_12187);
or U15231 (N_15231,N_10634,N_12058);
or U15232 (N_15232,N_13945,N_12968);
nor U15233 (N_15233,N_11539,N_10767);
or U15234 (N_15234,N_12068,N_14104);
or U15235 (N_15235,N_13404,N_10172);
or U15236 (N_15236,N_10779,N_13068);
nand U15237 (N_15237,N_14498,N_12413);
or U15238 (N_15238,N_11675,N_11313);
or U15239 (N_15239,N_12541,N_10578);
and U15240 (N_15240,N_13909,N_13976);
nand U15241 (N_15241,N_10900,N_12772);
nor U15242 (N_15242,N_11219,N_11898);
nand U15243 (N_15243,N_14549,N_10456);
or U15244 (N_15244,N_14023,N_10888);
and U15245 (N_15245,N_13637,N_12597);
or U15246 (N_15246,N_14838,N_14000);
nor U15247 (N_15247,N_12097,N_13208);
and U15248 (N_15248,N_13228,N_10107);
or U15249 (N_15249,N_14999,N_10195);
nand U15250 (N_15250,N_11255,N_12043);
nor U15251 (N_15251,N_14754,N_11874);
and U15252 (N_15252,N_11860,N_13393);
and U15253 (N_15253,N_11294,N_12179);
or U15254 (N_15254,N_10081,N_11047);
or U15255 (N_15255,N_13173,N_13398);
or U15256 (N_15256,N_11784,N_13401);
nor U15257 (N_15257,N_13048,N_14176);
or U15258 (N_15258,N_11803,N_13538);
or U15259 (N_15259,N_13989,N_12305);
nor U15260 (N_15260,N_12980,N_13678);
and U15261 (N_15261,N_10549,N_14118);
nand U15262 (N_15262,N_12676,N_14094);
or U15263 (N_15263,N_13763,N_12810);
nor U15264 (N_15264,N_11858,N_12247);
nor U15265 (N_15265,N_14753,N_12350);
or U15266 (N_15266,N_11269,N_11001);
nand U15267 (N_15267,N_12742,N_11360);
nand U15268 (N_15268,N_14119,N_10068);
or U15269 (N_15269,N_14855,N_10702);
nor U15270 (N_15270,N_13179,N_12707);
and U15271 (N_15271,N_10283,N_14797);
and U15272 (N_15272,N_14331,N_11419);
nand U15273 (N_15273,N_10007,N_14418);
and U15274 (N_15274,N_13045,N_14598);
or U15275 (N_15275,N_13187,N_14648);
xnor U15276 (N_15276,N_12320,N_13453);
nand U15277 (N_15277,N_13275,N_12060);
nor U15278 (N_15278,N_14865,N_12005);
or U15279 (N_15279,N_10481,N_10636);
and U15280 (N_15280,N_11814,N_14741);
nand U15281 (N_15281,N_14358,N_11748);
nor U15282 (N_15282,N_11343,N_10923);
nand U15283 (N_15283,N_10692,N_13572);
or U15284 (N_15284,N_13206,N_13917);
or U15285 (N_15285,N_11908,N_10465);
or U15286 (N_15286,N_14107,N_12949);
or U15287 (N_15287,N_10859,N_10848);
and U15288 (N_15288,N_14497,N_10533);
nand U15289 (N_15289,N_13684,N_13613);
nor U15290 (N_15290,N_10750,N_12548);
or U15291 (N_15291,N_12493,N_14381);
or U15292 (N_15292,N_10624,N_11440);
or U15293 (N_15293,N_12899,N_12591);
nand U15294 (N_15294,N_12273,N_13110);
or U15295 (N_15295,N_14113,N_14258);
or U15296 (N_15296,N_11202,N_13688);
or U15297 (N_15297,N_11327,N_10328);
nor U15298 (N_15298,N_13606,N_14622);
nor U15299 (N_15299,N_11622,N_10814);
and U15300 (N_15300,N_13409,N_10393);
nor U15301 (N_15301,N_10738,N_14617);
and U15302 (N_15302,N_12071,N_13558);
or U15303 (N_15303,N_10455,N_13705);
or U15304 (N_15304,N_13956,N_11339);
nor U15305 (N_15305,N_12467,N_10103);
and U15306 (N_15306,N_12930,N_14071);
nand U15307 (N_15307,N_13138,N_11604);
nor U15308 (N_15308,N_14562,N_14022);
xnor U15309 (N_15309,N_13588,N_11590);
and U15310 (N_15310,N_11610,N_14153);
nand U15311 (N_15311,N_13849,N_12123);
nor U15312 (N_15312,N_12348,N_11634);
or U15313 (N_15313,N_13212,N_12199);
and U15314 (N_15314,N_12549,N_14159);
nand U15315 (N_15315,N_10278,N_12730);
or U15316 (N_15316,N_10029,N_10617);
and U15317 (N_15317,N_10548,N_14942);
or U15318 (N_15318,N_14938,N_12624);
and U15319 (N_15319,N_10766,N_14024);
or U15320 (N_15320,N_13951,N_14290);
nor U15321 (N_15321,N_13973,N_12149);
or U15322 (N_15322,N_13218,N_10477);
or U15323 (N_15323,N_10247,N_13563);
nand U15324 (N_15324,N_13109,N_14626);
nor U15325 (N_15325,N_11964,N_11588);
nor U15326 (N_15326,N_12414,N_10326);
and U15327 (N_15327,N_11373,N_12323);
nor U15328 (N_15328,N_11382,N_11544);
and U15329 (N_15329,N_12617,N_11384);
and U15330 (N_15330,N_12483,N_13226);
nand U15331 (N_15331,N_10649,N_11716);
and U15332 (N_15332,N_12315,N_13805);
and U15333 (N_15333,N_10072,N_10713);
nand U15334 (N_15334,N_10595,N_10563);
and U15335 (N_15335,N_10569,N_12601);
nor U15336 (N_15336,N_12692,N_12511);
or U15337 (N_15337,N_12275,N_11707);
or U15338 (N_15338,N_12989,N_11905);
nand U15339 (N_15339,N_12298,N_13621);
nor U15340 (N_15340,N_14971,N_11808);
nand U15341 (N_15341,N_14033,N_13460);
or U15342 (N_15342,N_13411,N_12940);
nand U15343 (N_15343,N_11594,N_14886);
or U15344 (N_15344,N_13354,N_13616);
and U15345 (N_15345,N_12851,N_10066);
nand U15346 (N_15346,N_12937,N_10955);
nand U15347 (N_15347,N_13160,N_12112);
and U15348 (N_15348,N_11686,N_14735);
or U15349 (N_15349,N_12371,N_12879);
and U15350 (N_15350,N_14836,N_13391);
or U15351 (N_15351,N_13259,N_10273);
and U15352 (N_15352,N_11541,N_13262);
nand U15353 (N_15353,N_12849,N_14673);
nor U15354 (N_15354,N_14355,N_10046);
nor U15355 (N_15355,N_10886,N_13476);
and U15356 (N_15356,N_13718,N_12927);
and U15357 (N_15357,N_12981,N_13754);
nor U15358 (N_15358,N_11226,N_12961);
nand U15359 (N_15359,N_12592,N_10163);
and U15360 (N_15360,N_14485,N_13102);
or U15361 (N_15361,N_11081,N_14079);
nor U15362 (N_15362,N_13812,N_13278);
or U15363 (N_15363,N_10293,N_12872);
and U15364 (N_15364,N_12888,N_12173);
and U15365 (N_15365,N_12858,N_11721);
or U15366 (N_15366,N_13920,N_12560);
nor U15367 (N_15367,N_14600,N_14394);
or U15368 (N_15368,N_14443,N_13491);
nor U15369 (N_15369,N_14870,N_12770);
nand U15370 (N_15370,N_14295,N_14263);
nor U15371 (N_15371,N_13346,N_10447);
and U15372 (N_15372,N_13017,N_11689);
nand U15373 (N_15373,N_13013,N_14864);
or U15374 (N_15374,N_13433,N_14682);
or U15375 (N_15375,N_12914,N_11064);
nand U15376 (N_15376,N_14470,N_10758);
nor U15377 (N_15377,N_12010,N_14546);
or U15378 (N_15378,N_10699,N_10832);
or U15379 (N_15379,N_12115,N_14316);
and U15380 (N_15380,N_10259,N_11841);
and U15381 (N_15381,N_14229,N_11584);
nand U15382 (N_15382,N_12124,N_14582);
and U15383 (N_15383,N_14074,N_10755);
or U15384 (N_15384,N_11290,N_11975);
nand U15385 (N_15385,N_12869,N_14077);
and U15386 (N_15386,N_12609,N_10830);
nor U15387 (N_15387,N_10196,N_12782);
nor U15388 (N_15388,N_10950,N_14008);
nor U15389 (N_15389,N_13609,N_13328);
or U15390 (N_15390,N_14140,N_12113);
nand U15391 (N_15391,N_10280,N_14173);
and U15392 (N_15392,N_12081,N_10241);
and U15393 (N_15393,N_14337,N_13062);
nand U15394 (N_15394,N_13086,N_11231);
nand U15395 (N_15395,N_12126,N_14459);
nand U15396 (N_15396,N_12098,N_10802);
or U15397 (N_15397,N_10302,N_11217);
and U15398 (N_15398,N_13198,N_12718);
or U15399 (N_15399,N_11529,N_10600);
and U15400 (N_15400,N_11295,N_12535);
nand U15401 (N_15401,N_10906,N_10431);
and U15402 (N_15402,N_12485,N_13234);
xnor U15403 (N_15403,N_14427,N_10764);
nand U15404 (N_15404,N_14280,N_10907);
nor U15405 (N_15405,N_12006,N_14908);
or U15406 (N_15406,N_13366,N_10593);
xnor U15407 (N_15407,N_10317,N_13225);
or U15408 (N_15408,N_13111,N_13990);
and U15409 (N_15409,N_10486,N_10002);
or U15410 (N_15410,N_11215,N_13926);
nand U15411 (N_15411,N_10101,N_10450);
and U15412 (N_15412,N_12289,N_10240);
nand U15413 (N_15413,N_10915,N_11044);
xnor U15414 (N_15414,N_11432,N_13843);
and U15415 (N_15415,N_12367,N_12443);
nor U15416 (N_15416,N_13578,N_11301);
nand U15417 (N_15417,N_11851,N_11006);
nand U15418 (N_15418,N_14207,N_12574);
nor U15419 (N_15419,N_10523,N_13012);
nand U15420 (N_15420,N_11763,N_14414);
and U15421 (N_15421,N_12607,N_12128);
or U15422 (N_15422,N_14218,N_12430);
and U15423 (N_15423,N_13793,N_12448);
nand U15424 (N_15424,N_12856,N_10503);
nor U15425 (N_15425,N_13041,N_10423);
nand U15426 (N_15426,N_14013,N_10871);
and U15427 (N_15427,N_10397,N_12543);
nor U15428 (N_15428,N_13499,N_11965);
and U15429 (N_15429,N_13813,N_12161);
nor U15430 (N_15430,N_12542,N_10232);
nor U15431 (N_15431,N_13874,N_14108);
and U15432 (N_15432,N_14637,N_13270);
nand U15433 (N_15433,N_11349,N_14504);
and U15434 (N_15434,N_11635,N_13169);
nor U15435 (N_15435,N_11983,N_11606);
or U15436 (N_15436,N_12285,N_14847);
xor U15437 (N_15437,N_10861,N_14699);
nor U15438 (N_15438,N_11317,N_12423);
and U15439 (N_15439,N_14041,N_12748);
nor U15440 (N_15440,N_14211,N_12666);
nand U15441 (N_15441,N_11676,N_10130);
and U15442 (N_15442,N_11124,N_14468);
or U15443 (N_15443,N_11245,N_12649);
and U15444 (N_15444,N_13765,N_14988);
and U15445 (N_15445,N_14810,N_13430);
or U15446 (N_15446,N_14493,N_13959);
or U15447 (N_15447,N_14089,N_13285);
or U15448 (N_15448,N_11611,N_11727);
nand U15449 (N_15449,N_10990,N_10047);
or U15450 (N_15450,N_11310,N_11830);
or U15451 (N_15451,N_14242,N_11035);
nand U15452 (N_15452,N_12008,N_10579);
nor U15453 (N_15453,N_14841,N_14088);
nor U15454 (N_15454,N_14274,N_10314);
or U15455 (N_15455,N_12883,N_12988);
and U15456 (N_15456,N_13420,N_14638);
and U15457 (N_15457,N_14453,N_13204);
and U15458 (N_15458,N_12977,N_10260);
nor U15459 (N_15459,N_13091,N_11960);
nor U15460 (N_15460,N_14320,N_13468);
and U15461 (N_15461,N_13652,N_13073);
nand U15462 (N_15462,N_14532,N_14698);
and U15463 (N_15463,N_10717,N_12616);
nor U15464 (N_15464,N_13337,N_10508);
nor U15465 (N_15465,N_11671,N_14444);
or U15466 (N_15466,N_14155,N_10581);
or U15467 (N_15467,N_11577,N_11684);
nor U15468 (N_15468,N_11870,N_12056);
and U15469 (N_15469,N_12023,N_12990);
nor U15470 (N_15470,N_10723,N_14769);
and U15471 (N_15471,N_11937,N_12226);
and U15472 (N_15472,N_14795,N_14206);
and U15473 (N_15473,N_10025,N_11277);
and U15474 (N_15474,N_13353,N_11145);
nor U15475 (N_15475,N_12066,N_12263);
and U15476 (N_15476,N_12558,N_10178);
nor U15477 (N_15477,N_14028,N_11105);
nand U15478 (N_15478,N_10628,N_11162);
nand U15479 (N_15479,N_11074,N_10272);
nand U15480 (N_15480,N_13780,N_13787);
and U15481 (N_15481,N_10176,N_11782);
xnor U15482 (N_15482,N_11823,N_10388);
nor U15483 (N_15483,N_11429,N_13146);
nand U15484 (N_15484,N_14996,N_14105);
nand U15485 (N_15485,N_11552,N_13510);
nand U15486 (N_15486,N_10223,N_12523);
nor U15487 (N_15487,N_12499,N_10177);
nor U15488 (N_15488,N_10518,N_14346);
nand U15489 (N_15489,N_14471,N_10964);
nor U15490 (N_15490,N_10975,N_14812);
nand U15491 (N_15491,N_14625,N_13819);
nor U15492 (N_15492,N_14472,N_14844);
nand U15493 (N_15493,N_10793,N_13830);
nor U15494 (N_15494,N_14371,N_10645);
nor U15495 (N_15495,N_12487,N_13769);
and U15496 (N_15496,N_12806,N_14352);
xnor U15497 (N_15497,N_12809,N_14856);
nor U15498 (N_15498,N_12803,N_12318);
or U15499 (N_15499,N_10457,N_12841);
and U15500 (N_15500,N_10190,N_12779);
or U15501 (N_15501,N_13651,N_11401);
and U15502 (N_15502,N_11271,N_14396);
nor U15503 (N_15503,N_13057,N_11207);
and U15504 (N_15504,N_11358,N_14876);
nor U15505 (N_15505,N_13954,N_11287);
nor U15506 (N_15506,N_10076,N_13050);
nor U15507 (N_15507,N_12261,N_12357);
nor U15508 (N_15508,N_11167,N_13131);
nor U15509 (N_15509,N_13176,N_11475);
and U15510 (N_15510,N_12713,N_14958);
nor U15511 (N_15511,N_13100,N_14923);
nor U15512 (N_15512,N_12488,N_11002);
nor U15513 (N_15513,N_12427,N_12027);
and U15514 (N_15514,N_10705,N_10564);
or U15515 (N_15515,N_13786,N_14796);
or U15516 (N_15516,N_12303,N_11738);
nand U15517 (N_15517,N_12230,N_13521);
and U15518 (N_15518,N_14827,N_13037);
and U15519 (N_15519,N_14983,N_10090);
and U15520 (N_15520,N_10773,N_12970);
or U15521 (N_15521,N_14708,N_10540);
nand U15522 (N_15522,N_13417,N_13788);
nand U15523 (N_15523,N_14565,N_12167);
and U15524 (N_15524,N_12737,N_10179);
and U15525 (N_15525,N_12892,N_14463);
or U15526 (N_15526,N_10877,N_13281);
or U15527 (N_15527,N_14150,N_13674);
or U15528 (N_15528,N_11104,N_10445);
nand U15529 (N_15529,N_10042,N_14061);
and U15530 (N_15530,N_12891,N_13698);
and U15531 (N_15531,N_13498,N_12689);
nand U15532 (N_15532,N_14940,N_14842);
nor U15533 (N_15533,N_14243,N_13865);
and U15534 (N_15534,N_11853,N_11755);
nor U15535 (N_15535,N_11025,N_10693);
nand U15536 (N_15536,N_14017,N_14249);
nor U15537 (N_15537,N_12902,N_11146);
nand U15538 (N_15538,N_10057,N_11362);
nor U15539 (N_15539,N_14422,N_14193);
nand U15540 (N_15540,N_12783,N_11042);
or U15541 (N_15541,N_11917,N_13180);
or U15542 (N_15542,N_10039,N_14607);
and U15543 (N_15543,N_10213,N_12551);
nor U15544 (N_15544,N_12327,N_12531);
nand U15545 (N_15545,N_14100,N_10170);
nor U15546 (N_15546,N_14725,N_12153);
nor U15547 (N_15547,N_14481,N_14730);
nand U15548 (N_15548,N_12484,N_12156);
nor U15549 (N_15549,N_14765,N_12999);
and U15550 (N_15550,N_10080,N_13134);
nand U15551 (N_15551,N_14674,N_12322);
nand U15552 (N_15552,N_13416,N_11079);
nor U15553 (N_15553,N_13540,N_10226);
or U15554 (N_15554,N_12386,N_14613);
nor U15555 (N_15555,N_12284,N_13746);
and U15556 (N_15556,N_14333,N_10561);
nor U15557 (N_15557,N_11507,N_10753);
and U15558 (N_15558,N_14499,N_14798);
nand U15559 (N_15559,N_13821,N_14161);
nand U15560 (N_15560,N_14198,N_12046);
and U15561 (N_15561,N_12140,N_13634);
or U15562 (N_15562,N_10938,N_14768);
or U15563 (N_15563,N_14816,N_13915);
nand U15564 (N_15564,N_12768,N_12447);
nor U15565 (N_15565,N_10485,N_14457);
nor U15566 (N_15566,N_12169,N_13236);
nand U15567 (N_15567,N_10719,N_13969);
nand U15568 (N_15568,N_13360,N_10903);
nor U15569 (N_15569,N_14382,N_10282);
xor U15570 (N_15570,N_14431,N_11471);
nand U15571 (N_15571,N_12192,N_11062);
or U15572 (N_15572,N_10074,N_13931);
nand U15573 (N_15573,N_11354,N_10372);
nor U15574 (N_15574,N_14260,N_11789);
nand U15575 (N_15575,N_14492,N_13593);
nand U15576 (N_15576,N_11220,N_12727);
nor U15577 (N_15577,N_14184,N_11601);
or U15578 (N_15578,N_14204,N_11378);
or U15579 (N_15579,N_14405,N_13369);
nor U15580 (N_15580,N_10909,N_13952);
xnor U15581 (N_15581,N_10048,N_10199);
nor U15582 (N_15582,N_14345,N_10200);
nand U15583 (N_15583,N_11768,N_10437);
nor U15584 (N_15584,N_13818,N_14148);
nor U15585 (N_15585,N_12438,N_12733);
or U15586 (N_15586,N_12675,N_13611);
or U15587 (N_15587,N_12072,N_10784);
or U15588 (N_15588,N_10288,N_13511);
nor U15589 (N_15589,N_10432,N_13484);
nand U15590 (N_15590,N_11316,N_13654);
nor U15591 (N_15591,N_13248,N_11813);
xnor U15592 (N_15592,N_13341,N_14757);
and U15593 (N_15593,N_14909,N_11297);
or U15594 (N_15594,N_13798,N_13458);
nand U15595 (N_15595,N_12186,N_11582);
nand U15596 (N_15596,N_10586,N_12258);
or U15597 (N_15597,N_14657,N_10988);
or U15598 (N_15598,N_12079,N_10946);
and U15599 (N_15599,N_12142,N_10365);
and U15600 (N_15600,N_14447,N_11229);
or U15601 (N_15601,N_10127,N_13577);
nor U15602 (N_15602,N_11375,N_13189);
nor U15603 (N_15603,N_11161,N_10464);
nor U15604 (N_15604,N_10577,N_14892);
nor U15605 (N_15605,N_12435,N_13116);
nor U15606 (N_15606,N_10730,N_11928);
and U15607 (N_15607,N_14002,N_14336);
nand U15608 (N_15608,N_11519,N_10721);
nand U15609 (N_15609,N_10405,N_11609);
nand U15610 (N_15610,N_11649,N_11907);
or U15611 (N_15611,N_12561,N_10474);
and U15612 (N_15612,N_10419,N_12264);
and U15613 (N_15613,N_14883,N_13700);
or U15614 (N_15614,N_14922,N_12157);
nor U15615 (N_15615,N_12996,N_11321);
or U15616 (N_15616,N_13361,N_11213);
nand U15617 (N_15617,N_12409,N_10828);
or U15618 (N_15618,N_12684,N_13300);
or U15619 (N_15619,N_10850,N_13853);
nor U15620 (N_15620,N_14830,N_12691);
and U15621 (N_15621,N_11589,N_10069);
nor U15622 (N_15622,N_10088,N_14531);
or U15623 (N_15623,N_13993,N_11617);
or U15624 (N_15624,N_11396,N_11850);
nand U15625 (N_15625,N_11197,N_14848);
nand U15626 (N_15626,N_10440,N_14712);
nand U15627 (N_15627,N_14244,N_14567);
nand U15628 (N_15628,N_14653,N_10292);
nor U15629 (N_15629,N_13331,N_14540);
or U15630 (N_15630,N_13683,N_14641);
and U15631 (N_15631,N_10571,N_11921);
and U15632 (N_15632,N_11307,N_10997);
nand U15633 (N_15633,N_12934,N_12411);
nand U15634 (N_15634,N_13771,N_10686);
and U15635 (N_15635,N_12784,N_11679);
or U15636 (N_15636,N_14934,N_13202);
and U15637 (N_15637,N_12514,N_11412);
nor U15638 (N_15638,N_13847,N_14484);
and U15639 (N_15639,N_13633,N_11469);
and U15640 (N_15640,N_11902,N_13351);
and U15641 (N_15641,N_13392,N_14144);
or U15642 (N_15642,N_13583,N_11179);
nand U15643 (N_15643,N_12137,N_12132);
nor U15644 (N_15644,N_12871,N_11710);
nor U15645 (N_15645,N_12517,N_10387);
nand U15646 (N_15646,N_14987,N_12001);
and U15647 (N_15647,N_14927,N_14952);
or U15648 (N_15648,N_10145,N_11949);
nor U15649 (N_15649,N_14401,N_12236);
and U15650 (N_15650,N_11450,N_13309);
nor U15651 (N_15651,N_11693,N_10852);
and U15652 (N_15652,N_14820,N_13789);
nand U15653 (N_15653,N_13355,N_14777);
or U15654 (N_15654,N_11776,N_14262);
or U15655 (N_15655,N_10471,N_10782);
or U15656 (N_15656,N_12652,N_13635);
nor U15657 (N_15657,N_12242,N_10104);
nor U15658 (N_15658,N_11800,N_12191);
or U15659 (N_15659,N_11463,N_13519);
nand U15660 (N_15660,N_13323,N_14379);
and U15661 (N_15661,N_14083,N_13269);
nor U15662 (N_15662,N_12439,N_14252);
or U15663 (N_15663,N_11430,N_10202);
or U15664 (N_15664,N_14972,N_14049);
nand U15665 (N_15665,N_13701,N_10373);
nand U15666 (N_15666,N_12938,N_12415);
nor U15667 (N_15667,N_11828,N_10949);
and U15668 (N_15668,N_14296,N_10211);
nand U15669 (N_15669,N_12291,N_10301);
nor U15670 (N_15670,N_10459,N_14529);
or U15671 (N_15671,N_10528,N_10740);
nand U15672 (N_15672,N_12599,N_13516);
and U15673 (N_15673,N_11318,N_12176);
and U15674 (N_15674,N_11664,N_13716);
xor U15675 (N_15675,N_14250,N_14543);
and U15676 (N_15676,N_14821,N_12830);
nand U15677 (N_15677,N_12065,N_12328);
nand U15678 (N_15678,N_10835,N_10882);
and U15679 (N_15679,N_14270,N_12602);
nand U15680 (N_15680,N_11873,N_14102);
nand U15681 (N_15681,N_14949,N_14221);
nor U15682 (N_15682,N_13055,N_12513);
xnor U15683 (N_15683,N_11786,N_13533);
xor U15684 (N_15684,N_12644,N_10116);
or U15685 (N_15685,N_12876,N_11099);
nor U15686 (N_15686,N_10185,N_14537);
nor U15687 (N_15687,N_13372,N_13255);
xor U15688 (N_15688,N_12556,N_11699);
and U15689 (N_15689,N_12820,N_12063);
and U15690 (N_15690,N_13645,N_14301);
and U15691 (N_15691,N_10065,N_12947);
and U15692 (N_15692,N_12529,N_13394);
nand U15693 (N_15693,N_13580,N_13962);
nand U15694 (N_15694,N_12818,N_11551);
or U15695 (N_15695,N_12611,N_10547);
or U15696 (N_15696,N_14424,N_13912);
or U15697 (N_15697,N_11164,N_12894);
nand U15698 (N_15698,N_11054,N_11868);
and U15699 (N_15699,N_10466,N_11646);
and U15700 (N_15700,N_13852,N_13141);
xnor U15701 (N_15701,N_13719,N_10084);
nand U15702 (N_15702,N_13065,N_10295);
or U15703 (N_15703,N_14761,N_13299);
and U15704 (N_15704,N_12518,N_10816);
or U15705 (N_15705,N_10112,N_12394);
or U15706 (N_15706,N_12210,N_10233);
and U15707 (N_15707,N_10880,N_11043);
and U15708 (N_15708,N_14462,N_11968);
or U15709 (N_15709,N_14257,N_13066);
xnor U15710 (N_15710,N_14719,N_10031);
nor U15711 (N_15711,N_14906,N_12051);
nand U15712 (N_15712,N_13704,N_12222);
or U15713 (N_15713,N_11503,N_12292);
nand U15714 (N_15714,N_10193,N_10126);
nor U15715 (N_15715,N_12509,N_13462);
and U15716 (N_15716,N_10865,N_13560);
nor U15717 (N_15717,N_12753,N_10148);
nand U15718 (N_15718,N_14399,N_12593);
nand U15719 (N_15719,N_11974,N_12654);
nor U15720 (N_15720,N_12159,N_14326);
and U15721 (N_15721,N_13338,N_13342);
nand U15722 (N_15722,N_12708,N_10605);
or U15723 (N_15723,N_13747,N_10385);
or U15724 (N_15724,N_12002,N_14325);
nor U15725 (N_15725,N_11553,N_12771);
nand U15726 (N_15726,N_12102,N_13348);
nor U15727 (N_15727,N_10299,N_13575);
nand U15728 (N_15728,N_10441,N_11837);
and U15729 (N_15729,N_13972,N_11488);
and U15730 (N_15730,N_14729,N_13697);
or U15731 (N_15731,N_10654,N_11540);
and U15732 (N_15732,N_13795,N_10425);
or U15733 (N_15733,N_11896,N_10098);
or U15734 (N_15734,N_11195,N_11073);
nand U15735 (N_15735,N_14738,N_11565);
nor U15736 (N_15736,N_12547,N_13905);
or U15737 (N_15737,N_14808,N_13375);
nand U15738 (N_15738,N_11767,N_10161);
or U15739 (N_15739,N_11656,N_13627);
or U15740 (N_15740,N_14324,N_11460);
and U15741 (N_15741,N_12288,N_14873);
nand U15742 (N_15742,N_13378,N_10191);
and U15743 (N_15743,N_13672,N_12628);
nor U15744 (N_15744,N_12709,N_14759);
nor U15745 (N_15745,N_11189,N_12763);
nand U15746 (N_15746,N_12106,N_11410);
nand U15747 (N_15747,N_13090,N_11842);
or U15748 (N_15748,N_12639,N_10920);
nor U15749 (N_15749,N_12757,N_11797);
or U15750 (N_15750,N_12269,N_11756);
nand U15751 (N_15751,N_13828,N_14406);
and U15752 (N_15752,N_14087,N_13607);
or U15753 (N_15753,N_14974,N_10020);
nand U15754 (N_15754,N_14964,N_14039);
or U15755 (N_15755,N_11046,N_11116);
nor U15756 (N_15756,N_14048,N_12834);
and U15757 (N_15757,N_14634,N_11935);
xnor U15758 (N_15758,N_10630,N_14461);
and U15759 (N_15759,N_12794,N_10330);
nand U15760 (N_15760,N_12790,N_13026);
or U15761 (N_15761,N_11618,N_14880);
nand U15762 (N_15762,N_10994,N_11406);
nor U15763 (N_15763,N_14476,N_13023);
and U15764 (N_15764,N_14718,N_10701);
nor U15765 (N_15765,N_13063,N_13310);
and U15766 (N_15766,N_12613,N_12445);
and U15767 (N_15767,N_14794,N_14254);
or U15768 (N_15768,N_14477,N_13598);
and U15769 (N_15769,N_13046,N_11227);
or U15770 (N_15770,N_11381,N_12373);
nand U15771 (N_15771,N_14175,N_14589);
or U15772 (N_15772,N_13646,N_12502);
and U15773 (N_15773,N_10544,N_14654);
nand U15774 (N_15774,N_10378,N_12870);
nand U15775 (N_15775,N_14750,N_14512);
nor U15776 (N_15776,N_11370,N_13093);
nor U15777 (N_15777,N_10897,N_12890);
nor U15778 (N_15778,N_11329,N_12278);
nor U15779 (N_15779,N_13658,N_13356);
nor U15780 (N_15780,N_13617,N_13128);
or U15781 (N_15781,N_14662,N_10327);
xnor U15782 (N_15782,N_11182,N_10407);
nor U15783 (N_15783,N_13004,N_11443);
nand U15784 (N_15784,N_13834,N_10763);
and U15785 (N_15785,N_13214,N_10162);
nand U15786 (N_15786,N_14216,N_13423);
nor U15787 (N_15787,N_12969,N_14781);
and U15788 (N_15788,N_13205,N_11088);
and U15789 (N_15789,N_11942,N_12875);
nor U15790 (N_15790,N_10096,N_14602);
or U15791 (N_15791,N_12728,N_10556);
and U15792 (N_15792,N_11796,N_11456);
or U15793 (N_15793,N_12860,N_14084);
or U15794 (N_15794,N_12680,N_11494);
or U15795 (N_15795,N_10857,N_14055);
nand U15796 (N_15796,N_13171,N_14378);
nand U15797 (N_15797,N_10677,N_11702);
nor U15798 (N_15798,N_11660,N_10224);
nor U15799 (N_15799,N_13525,N_12216);
nor U15800 (N_15800,N_13772,N_11843);
and U15801 (N_15801,N_12950,N_13892);
nor U15802 (N_15802,N_12736,N_14410);
nor U15803 (N_15803,N_12789,N_12466);
or U15804 (N_15804,N_13657,N_12668);
or U15805 (N_15805,N_10082,N_11212);
nand U15806 (N_15806,N_13287,N_14291);
nor U15807 (N_15807,N_12074,N_11293);
nand U15808 (N_15808,N_13257,N_14985);
or U15809 (N_15809,N_13243,N_14318);
nand U15810 (N_15810,N_14950,N_11575);
and U15811 (N_15811,N_11408,N_13070);
or U15812 (N_15812,N_14756,N_13288);
or U15813 (N_15813,N_14921,N_10972);
nand U15814 (N_15814,N_14849,N_10943);
nor U15815 (N_15815,N_12850,N_11157);
and U15816 (N_15816,N_10480,N_13822);
nor U15817 (N_15817,N_10914,N_12585);
nor U15818 (N_15818,N_10977,N_11864);
nor U15819 (N_15819,N_13483,N_12345);
and U15820 (N_15820,N_12265,N_12133);
nor U15821 (N_15821,N_12942,N_10089);
nor U15822 (N_15822,N_10334,N_11423);
nor U15823 (N_15823,N_10438,N_10948);
and U15824 (N_15824,N_11657,N_13298);
nor U15825 (N_15825,N_12441,N_11379);
and U15826 (N_15826,N_12237,N_14435);
and U15827 (N_15827,N_10216,N_13245);
nand U15828 (N_15828,N_12566,N_14685);
nand U15829 (N_15829,N_10136,N_11573);
or U15830 (N_15830,N_11045,N_12648);
or U15831 (N_15831,N_14124,N_14315);
nand U15832 (N_15832,N_10133,N_11059);
nor U15833 (N_15833,N_12032,N_14858);
nand U15834 (N_15834,N_11286,N_12594);
nand U15835 (N_15835,N_13481,N_11049);
nand U15836 (N_15836,N_14959,N_11484);
and U15837 (N_15837,N_14713,N_14021);
and U15838 (N_15838,N_10777,N_10488);
and U15839 (N_15839,N_12501,N_13442);
or U15840 (N_15840,N_13507,N_12240);
and U15841 (N_15841,N_12637,N_11391);
nand U15842 (N_15842,N_11694,N_14692);
and U15843 (N_15843,N_11091,N_14806);
nand U15844 (N_15844,N_12045,N_12735);
or U15845 (N_15845,N_11600,N_11347);
or U15846 (N_15846,N_14389,N_14046);
or U15847 (N_15847,N_12012,N_12147);
or U15848 (N_15848,N_10298,N_10968);
and U15849 (N_15849,N_11308,N_13145);
nor U15850 (N_15850,N_12340,N_12144);
and U15851 (N_15851,N_14650,N_12267);
nand U15852 (N_15852,N_11852,N_11535);
nand U15853 (N_15853,N_14658,N_12901);
nand U15854 (N_15854,N_12033,N_11235);
nand U15855 (N_15855,N_11969,N_10236);
nor U15856 (N_15856,N_13703,N_10826);
or U15857 (N_15857,N_10408,N_11504);
and U15858 (N_15858,N_13220,N_14191);
nor U15859 (N_15859,N_14478,N_14335);
or U15860 (N_15860,N_14068,N_12055);
or U15861 (N_15861,N_13902,N_11880);
and U15862 (N_15862,N_13466,N_14495);
or U15863 (N_15863,N_10446,N_14018);
nor U15864 (N_15864,N_13564,N_14825);
and U15865 (N_15865,N_10479,N_11254);
or U15866 (N_15866,N_11148,N_11950);
nor U15867 (N_15867,N_10219,N_10050);
or U15868 (N_15868,N_12376,N_10908);
nand U15869 (N_15869,N_13127,N_11991);
nand U15870 (N_15870,N_13410,N_13628);
nand U15871 (N_15871,N_13783,N_11593);
and U15872 (N_15872,N_11725,N_12388);
nor U15873 (N_15873,N_12598,N_11201);
and U15874 (N_15874,N_10627,N_13732);
and U15875 (N_15875,N_14132,N_12030);
or U15876 (N_15876,N_10124,N_10840);
nor U15877 (N_15877,N_13946,N_14436);
or U15878 (N_15878,N_12983,N_14642);
or U15879 (N_15879,N_12831,N_12122);
nor U15880 (N_15880,N_10674,N_12910);
and U15881 (N_15881,N_14570,N_10403);
and U15882 (N_15882,N_10904,N_12516);
nand U15883 (N_15883,N_11747,N_11749);
nor U15884 (N_15884,N_13162,N_13965);
nor U15885 (N_15885,N_13870,N_12166);
and U15886 (N_15886,N_12868,N_12164);
and U15887 (N_15887,N_11149,N_11652);
and U15888 (N_15888,N_13151,N_13164);
nand U15889 (N_15889,N_13928,N_10381);
or U15890 (N_15890,N_12151,N_14672);
and U15891 (N_15891,N_13869,N_13724);
nor U15892 (N_15892,N_11409,N_10214);
nor U15893 (N_15893,N_10121,N_10973);
nor U15894 (N_15894,N_14183,N_12795);
nor U15895 (N_15895,N_10439,N_14995);
or U15896 (N_15896,N_11275,N_14833);
nor U15897 (N_15897,N_14566,N_11889);
xnor U15898 (N_15898,N_14980,N_12482);
nor U15899 (N_15899,N_10336,N_12778);
nor U15900 (N_15900,N_11840,N_11166);
and U15901 (N_15901,N_13251,N_14121);
xnor U15902 (N_15902,N_14935,N_12141);
and U15903 (N_15903,N_13207,N_12948);
or U15904 (N_15904,N_14905,N_11192);
and U15905 (N_15905,N_14516,N_10607);
nand U15906 (N_15906,N_13358,N_10933);
or U15907 (N_15907,N_10028,N_10058);
nor U15908 (N_15908,N_12685,N_11625);
and U15909 (N_15909,N_13717,N_12084);
nand U15910 (N_15910,N_11132,N_10234);
or U15911 (N_15911,N_10837,N_12175);
nor U15912 (N_15912,N_11639,N_10970);
and U15913 (N_15913,N_11390,N_14241);
nand U15914 (N_15914,N_12319,N_10324);
nor U15915 (N_15915,N_14978,N_12392);
nor U15916 (N_15916,N_11138,N_10683);
nand U15917 (N_15917,N_12724,N_14845);
or U15918 (N_15918,N_12671,N_10159);
nand U15919 (N_15919,N_10855,N_14067);
nand U15920 (N_15920,N_11422,N_13602);
or U15921 (N_15921,N_10192,N_13743);
nor U15922 (N_15922,N_10489,N_11506);
or U15923 (N_15923,N_10061,N_10063);
and U15924 (N_15924,N_13888,N_11792);
and U15925 (N_15925,N_11933,N_14370);
nand U15926 (N_15926,N_14112,N_12744);
nor U15927 (N_15927,N_12150,N_12546);
nor U15928 (N_15928,N_11838,N_12406);
nor U15929 (N_15929,N_14238,N_11296);
or U15930 (N_15930,N_11448,N_14255);
nor U15931 (N_15931,N_13367,N_11562);
or U15932 (N_15932,N_11017,N_10413);
nand U15933 (N_15933,N_12195,N_10567);
and U15934 (N_15934,N_12673,N_14720);
nor U15935 (N_15935,N_14955,N_11783);
and U15936 (N_15936,N_13085,N_10105);
nand U15937 (N_15937,N_13759,N_14752);
nor U15938 (N_15938,N_13486,N_12579);
nor U15939 (N_15939,N_13168,N_11453);
nand U15940 (N_15940,N_14360,N_12955);
or U15941 (N_15941,N_13604,N_13940);
and U15942 (N_15942,N_14060,N_12979);
nor U15943 (N_15943,N_10426,N_10143);
or U15944 (N_15944,N_11915,N_13887);
xnor U15945 (N_15945,N_12131,N_13408);
and U15946 (N_15946,N_10335,N_13589);
or U15947 (N_15947,N_11542,N_11437);
and U15948 (N_15948,N_10979,N_10697);
and U15949 (N_15949,N_10809,N_10598);
or U15950 (N_15950,N_13106,N_10783);
nand U15951 (N_15951,N_10604,N_11861);
or U15952 (N_15952,N_13612,N_12370);
nand U15953 (N_15953,N_13286,N_11242);
and U15954 (N_15954,N_14030,N_14902);
or U15955 (N_15955,N_14145,N_12252);
nand U15956 (N_15956,N_13461,N_12928);
or U15957 (N_15957,N_13447,N_12154);
nor U15958 (N_15958,N_10235,N_10349);
and U15959 (N_15959,N_11879,N_13067);
or U15960 (N_15960,N_14989,N_13427);
nor U15961 (N_15961,N_10374,N_14853);
and U15962 (N_15962,N_11129,N_13124);
xor U15963 (N_15963,N_14885,N_14611);
nor U15964 (N_15964,N_11181,N_12244);
nand U15965 (N_15965,N_10660,N_14224);
nand U15966 (N_15966,N_13051,N_14623);
and U15967 (N_15967,N_12307,N_13690);
nand U15968 (N_15968,N_14027,N_11335);
or U15969 (N_15969,N_13573,N_12973);
and U15970 (N_15970,N_13882,N_14248);
and U15971 (N_15971,N_11400,N_11258);
and U15972 (N_15972,N_13707,N_14116);
nor U15973 (N_15973,N_10342,N_12760);
nor U15974 (N_15974,N_11583,N_14605);
or U15975 (N_15975,N_11728,N_12009);
and U15976 (N_15976,N_14802,N_12456);
nor U15977 (N_15977,N_10167,N_12408);
nand U15978 (N_15978,N_10836,N_10303);
and U15979 (N_15979,N_13223,N_14494);
or U15980 (N_15980,N_12279,N_14322);
or U15981 (N_15981,N_14580,N_13244);
nand U15982 (N_15982,N_12463,N_14956);
nor U15983 (N_15983,N_13591,N_12669);
and U15984 (N_15984,N_11438,N_13335);
and U15985 (N_15985,N_14188,N_11230);
and U15986 (N_15986,N_14051,N_14851);
and U15987 (N_15987,N_13922,N_10573);
or U15988 (N_15988,N_14563,N_11486);
or U15989 (N_15989,N_13968,N_12326);
and U15990 (N_15990,N_12389,N_12824);
and U15991 (N_15991,N_14004,N_14866);
nor U15992 (N_15992,N_11680,N_10844);
nand U15993 (N_15993,N_14586,N_12232);
nor U15994 (N_15994,N_11040,N_10345);
nand U15995 (N_15995,N_14945,N_12576);
or U15996 (N_15996,N_14413,N_14548);
and U15997 (N_15997,N_14994,N_10810);
and U15998 (N_15998,N_11764,N_13557);
and U15999 (N_15999,N_14703,N_14701);
or U16000 (N_16000,N_14696,N_14551);
or U16001 (N_16001,N_11780,N_11510);
or U16002 (N_16002,N_10490,N_14621);
nor U16003 (N_16003,N_12245,N_14505);
nand U16004 (N_16004,N_11788,N_13562);
nor U16005 (N_16005,N_11619,N_10500);
or U16006 (N_16006,N_12044,N_13382);
or U16007 (N_16007,N_13978,N_10010);
nor U16008 (N_16008,N_14366,N_14603);
and U16009 (N_16009,N_12088,N_12886);
and U16010 (N_16010,N_11280,N_14714);
and U16011 (N_16011,N_11524,N_12925);
and U16012 (N_16012,N_14631,N_11775);
nand U16013 (N_16013,N_12864,N_11630);
and U16014 (N_16014,N_10661,N_11996);
nor U16015 (N_16015,N_11351,N_10174);
or U16016 (N_16016,N_10289,N_14234);
or U16017 (N_16017,N_14944,N_10789);
nand U16018 (N_16018,N_12537,N_12715);
or U16019 (N_16019,N_12087,N_14604);
and U16020 (N_16020,N_14737,N_10493);
and U16021 (N_16021,N_12459,N_12152);
nor U16022 (N_16022,N_10945,N_12995);
nand U16023 (N_16023,N_11566,N_10304);
or U16024 (N_16024,N_11012,N_12339);
nand U16025 (N_16025,N_14879,N_13103);
nor U16026 (N_16026,N_14171,N_10537);
or U16027 (N_16027,N_13166,N_12110);
and U16028 (N_16028,N_12476,N_13883);
and U16029 (N_16029,N_10478,N_13261);
nand U16030 (N_16030,N_11052,N_14651);
or U16031 (N_16031,N_10262,N_10733);
nor U16032 (N_16032,N_11214,N_11836);
nor U16033 (N_16033,N_13303,N_11696);
nor U16034 (N_16034,N_10243,N_11517);
nand U16035 (N_16035,N_13290,N_14760);
or U16036 (N_16036,N_11570,N_13844);
and U16037 (N_16037,N_14454,N_12207);
or U16038 (N_16038,N_10912,N_14465);
or U16039 (N_16039,N_12878,N_12916);
nor U16040 (N_16040,N_12335,N_12917);
or U16041 (N_16041,N_10515,N_13195);
nand U16042 (N_16042,N_14506,N_10944);
nand U16043 (N_16043,N_13040,N_13890);
nor U16044 (N_16044,N_14095,N_13581);
or U16045 (N_16045,N_14309,N_12799);
or U16046 (N_16046,N_14388,N_10205);
nor U16047 (N_16047,N_12077,N_11246);
or U16048 (N_16048,N_10443,N_10751);
and U16049 (N_16049,N_10222,N_14572);
and U16050 (N_16050,N_11638,N_12922);
or U16051 (N_16051,N_11496,N_12325);
nor U16052 (N_16052,N_11385,N_10274);
nor U16053 (N_16053,N_10401,N_10694);
nand U16054 (N_16054,N_13587,N_13820);
or U16055 (N_16055,N_11706,N_10140);
or U16056 (N_16056,N_10662,N_11556);
nand U16057 (N_16057,N_10512,N_12997);
nor U16058 (N_16058,N_14149,N_10412);
xor U16059 (N_16059,N_12904,N_14237);
nor U16060 (N_16060,N_10780,N_12492);
or U16061 (N_16061,N_13665,N_14393);
or U16062 (N_16062,N_10884,N_11793);
nand U16063 (N_16063,N_12780,N_13089);
or U16064 (N_16064,N_10941,N_10505);
or U16065 (N_16065,N_13895,N_12379);
nand U16066 (N_16066,N_10086,N_14420);
or U16067 (N_16067,N_11596,N_14045);
and U16068 (N_16068,N_11176,N_12418);
and U16069 (N_16069,N_12573,N_12867);
nor U16070 (N_16070,N_12952,N_12880);
and U16071 (N_16071,N_10761,N_10380);
nand U16072 (N_16072,N_11520,N_14912);
nand U16073 (N_16073,N_13619,N_14981);
or U16074 (N_16074,N_11094,N_12390);
nor U16075 (N_16075,N_11807,N_13222);
nand U16076 (N_16076,N_10064,N_14058);
and U16077 (N_16077,N_14612,N_14659);
or U16078 (N_16078,N_10363,N_12631);
nor U16079 (N_16079,N_11692,N_10969);
nor U16080 (N_16080,N_10246,N_12522);
nor U16081 (N_16081,N_12193,N_12075);
or U16082 (N_16082,N_13555,N_11993);
and U16083 (N_16083,N_12212,N_14426);
nand U16084 (N_16084,N_11955,N_11264);
nor U16085 (N_16085,N_11387,N_10294);
and U16086 (N_16086,N_13866,N_14306);
and U16087 (N_16087,N_14508,N_10264);
and U16088 (N_16088,N_11158,N_14488);
nor U16089 (N_16089,N_14578,N_12767);
xnor U16090 (N_16090,N_10083,N_14805);
xnor U16091 (N_16091,N_10918,N_14233);
or U16092 (N_16092,N_14734,N_13804);
or U16093 (N_16093,N_11199,N_11178);
and U16094 (N_16094,N_10144,N_10538);
or U16095 (N_16095,N_10475,N_10436);
and U16096 (N_16096,N_12725,N_14928);
and U16097 (N_16097,N_11821,N_12478);
nor U16098 (N_16098,N_12374,N_11244);
and U16099 (N_16099,N_11534,N_13914);
or U16100 (N_16100,N_11404,N_13446);
nor U16101 (N_16101,N_12035,N_10553);
or U16102 (N_16102,N_12181,N_14429);
or U16103 (N_16103,N_13273,N_14727);
and U16104 (N_16104,N_14913,N_11627);
or U16105 (N_16105,N_11513,N_13474);
nor U16106 (N_16106,N_11603,N_13623);
and U16107 (N_16107,N_10792,N_11458);
or U16108 (N_16108,N_10566,N_11140);
and U16109 (N_16109,N_14130,N_13240);
nor U16110 (N_16110,N_14009,N_11063);
and U16111 (N_16111,N_10960,N_12595);
nand U16112 (N_16112,N_12436,N_10114);
or U16113 (N_16113,N_13910,N_11744);
and U16114 (N_16114,N_11172,N_14179);
or U16115 (N_16115,N_12208,N_10115);
nor U16116 (N_16116,N_14619,N_12197);
nand U16117 (N_16117,N_11887,N_13477);
nor U16118 (N_16118,N_10689,N_11492);
and U16119 (N_16119,N_12203,N_12939);
and U16120 (N_16120,N_10982,N_12656);
and U16121 (N_16121,N_13373,N_12125);
and U16122 (N_16122,N_10878,N_12440);
or U16123 (N_16123,N_12007,N_14437);
nor U16124 (N_16124,N_12085,N_13005);
and U16125 (N_16125,N_13864,N_12552);
nand U16126 (N_16126,N_12257,N_12580);
nor U16127 (N_16127,N_11894,N_13508);
and U16128 (N_16128,N_11032,N_10188);
nor U16129 (N_16129,N_12272,N_10119);
or U16130 (N_16130,N_12862,N_12568);
and U16131 (N_16131,N_14588,N_14667);
and U16132 (N_16132,N_13677,N_13773);
nor U16133 (N_16133,N_10663,N_12881);
or U16134 (N_16134,N_11086,N_14666);
and U16135 (N_16135,N_10635,N_12873);
and U16136 (N_16136,N_12861,N_10639);
or U16137 (N_16137,N_13316,N_11567);
nor U16138 (N_16138,N_12665,N_12365);
or U16139 (N_16139,N_11169,N_12243);
and U16140 (N_16140,N_13796,N_10829);
xnor U16141 (N_16141,N_10642,N_12882);
xor U16142 (N_16142,N_11735,N_12437);
nor U16143 (N_16143,N_11724,N_11923);
and U16144 (N_16144,N_11723,N_12194);
nor U16145 (N_16145,N_12773,N_11405);
xor U16146 (N_16146,N_12480,N_11759);
xnor U16147 (N_16147,N_11833,N_12037);
nand U16148 (N_16148,N_14967,N_13029);
or U16149 (N_16149,N_13376,N_10012);
nand U16150 (N_16150,N_11824,N_12816);
and U16151 (N_16151,N_11546,N_14063);
nand U16152 (N_16152,N_14583,N_12286);
nor U16153 (N_16153,N_11478,N_10225);
and U16154 (N_16154,N_10678,N_12704);
nand U16155 (N_16155,N_13001,N_10514);
nor U16156 (N_16156,N_13024,N_13881);
and U16157 (N_16157,N_12630,N_10510);
nor U16158 (N_16158,N_14595,N_12229);
and U16159 (N_16159,N_10963,N_13794);
xor U16160 (N_16160,N_11516,N_10125);
and U16161 (N_16161,N_11106,N_12457);
nor U16162 (N_16162,N_13764,N_13201);
nand U16163 (N_16163,N_12683,N_14758);
nand U16164 (N_16164,N_10173,N_10995);
xnor U16165 (N_16165,N_10266,N_13407);
and U16166 (N_16166,N_11123,N_10079);
and U16167 (N_16167,N_11353,N_10670);
nand U16168 (N_16168,N_13981,N_11427);
nor U16169 (N_16169,N_10519,N_12530);
nand U16170 (N_16170,N_12014,N_14723);
and U16171 (N_16171,N_14644,N_14675);
nor U16172 (N_16172,N_14832,N_10774);
xor U16173 (N_16173,N_11681,N_14732);
and U16174 (N_16174,N_13839,N_13235);
or U16175 (N_16175,N_11731,N_12111);
or U16176 (N_16176,N_12354,N_13246);
or U16177 (N_16177,N_12536,N_11417);
and U16178 (N_16178,N_13641,N_10543);
nand U16179 (N_16179,N_10846,N_13463);
or U16180 (N_16180,N_13165,N_11098);
and U16181 (N_16181,N_13247,N_12036);
or U16182 (N_16182,N_13554,N_11498);
or U16183 (N_16183,N_12521,N_11160);
nor U16184 (N_16184,N_14181,N_12473);
xnor U16185 (N_16185,N_11644,N_13501);
nand U16186 (N_16186,N_14576,N_11305);
nand U16187 (N_16187,N_14446,N_13333);
and U16188 (N_16188,N_11717,N_11075);
and U16189 (N_16189,N_11457,N_10520);
xnor U16190 (N_16190,N_10182,N_14312);
or U16191 (N_16191,N_14090,N_11690);
and U16192 (N_16192,N_10276,N_11134);
nand U16193 (N_16193,N_14771,N_14791);
nor U16194 (N_16194,N_13076,N_10629);
nor U16195 (N_16195,N_12512,N_13872);
nand U16196 (N_16196,N_11279,N_13137);
and U16197 (N_16197,N_13659,N_10650);
or U16198 (N_16198,N_11881,N_10414);
or U16199 (N_16199,N_14430,N_13548);
and U16200 (N_16200,N_10501,N_14814);
nand U16201 (N_16201,N_11712,N_14867);
or U16202 (N_16202,N_13568,N_11459);
nor U16203 (N_16203,N_13332,N_14134);
nand U16204 (N_16204,N_14724,N_11994);
nor U16205 (N_16205,N_11101,N_12465);
nand U16206 (N_16206,N_11934,N_10018);
or U16207 (N_16207,N_12813,N_11021);
or U16208 (N_16208,N_14014,N_10067);
or U16209 (N_16209,N_13042,N_10321);
xor U16210 (N_16210,N_13193,N_13676);
or U16211 (N_16211,N_13006,N_14860);
xor U16212 (N_16212,N_13445,N_10546);
nor U16213 (N_16213,N_14500,N_11198);
nor U16214 (N_16214,N_10576,N_11726);
or U16215 (N_16215,N_12758,N_10868);
nand U16216 (N_16216,N_10059,N_10122);
and U16217 (N_16217,N_12446,N_10271);
nand U16218 (N_16218,N_11451,N_10833);
and U16219 (N_16219,N_14440,N_11633);
nor U16220 (N_16220,N_12178,N_12442);
or U16221 (N_16221,N_11900,N_14636);
nor U16222 (N_16222,N_13473,N_12936);
and U16223 (N_16223,N_14158,N_10929);
nor U16224 (N_16224,N_13105,N_11122);
and U16225 (N_16225,N_11407,N_10208);
and U16226 (N_16226,N_11938,N_11121);
and U16227 (N_16227,N_13726,N_10398);
nand U16228 (N_16228,N_10000,N_14710);
nand U16229 (N_16229,N_13664,N_13758);
nand U16230 (N_16230,N_11832,N_10197);
or U16231 (N_16231,N_14522,N_12608);
and U16232 (N_16232,N_10017,N_14807);
or U16233 (N_16233,N_11368,N_14910);
or U16234 (N_16234,N_12606,N_14557);
or U16235 (N_16235,N_11932,N_14040);
or U16236 (N_16236,N_10361,N_12505);
nand U16237 (N_16237,N_14891,N_12061);
nor U16238 (N_16238,N_11956,N_14330);
and U16239 (N_16239,N_14904,N_12745);
and U16240 (N_16240,N_11439,N_10872);
and U16241 (N_16241,N_10421,N_10621);
and U16242 (N_16242,N_14790,N_12064);
and U16243 (N_16243,N_11411,N_14711);
nor U16244 (N_16244,N_14226,N_12605);
or U16245 (N_16245,N_13504,N_14208);
nor U16246 (N_16246,N_13727,N_14328);
or U16247 (N_16247,N_10806,N_12696);
nand U16248 (N_16248,N_12506,N_14610);
or U16249 (N_16249,N_11827,N_12082);
and U16250 (N_16250,N_11509,N_14645);
nor U16251 (N_16251,N_13751,N_14340);
nand U16252 (N_16252,N_13694,N_14115);
and U16253 (N_16253,N_13840,N_12016);
and U16254 (N_16254,N_11927,N_10601);
or U16255 (N_16255,N_12924,N_12711);
nand U16256 (N_16256,N_13903,N_10053);
or U16257 (N_16257,N_13908,N_13766);
nor U16258 (N_16258,N_13826,N_10504);
xor U16259 (N_16259,N_11574,N_14823);
or U16260 (N_16260,N_12764,N_13308);
or U16261 (N_16261,N_13861,N_13415);
nor U16262 (N_16262,N_14661,N_13469);
nand U16263 (N_16263,N_12557,N_14200);
and U16264 (N_16264,N_10673,N_10137);
nor U16265 (N_16265,N_12135,N_14556);
or U16266 (N_16266,N_10418,N_13158);
or U16267 (N_16267,N_11338,N_10807);
nor U16268 (N_16268,N_14029,N_11865);
nor U16269 (N_16269,N_14809,N_11163);
or U16270 (N_16270,N_11491,N_11985);
and U16271 (N_16271,N_10656,N_14594);
nand U16272 (N_16272,N_11330,N_13918);
nor U16273 (N_16273,N_12587,N_10596);
and U16274 (N_16274,N_11322,N_14240);
and U16275 (N_16275,N_12380,N_12391);
nand U16276 (N_16276,N_10611,N_13078);
nor U16277 (N_16277,N_11714,N_10221);
nand U16278 (N_16278,N_12047,N_13464);
or U16279 (N_16279,N_11135,N_13161);
and U16280 (N_16280,N_14560,N_14411);
nor U16281 (N_16281,N_12700,N_13282);
or U16282 (N_16282,N_12148,N_10430);
nor U16283 (N_16283,N_11068,N_11558);
nand U16284 (N_16284,N_14169,N_11877);
nand U16285 (N_16285,N_11173,N_14194);
nand U16286 (N_16286,N_14483,N_13924);
nor U16287 (N_16287,N_12746,N_12460);
and U16288 (N_16288,N_13371,N_10375);
or U16289 (N_16289,N_13249,N_13860);
nand U16290 (N_16290,N_13536,N_10668);
nand U16291 (N_16291,N_10290,N_14283);
or U16292 (N_16292,N_12747,N_14163);
nand U16293 (N_16293,N_11599,N_11683);
nor U16294 (N_16294,N_13457,N_14341);
and U16295 (N_16295,N_13322,N_10149);
or U16296 (N_16296,N_10215,N_12221);
or U16297 (N_16297,N_11990,N_10591);
nor U16298 (N_16298,N_12053,N_13792);
and U16299 (N_16299,N_11753,N_13728);
or U16300 (N_16300,N_14228,N_10608);
and U16301 (N_16301,N_13567,N_10879);
and U16302 (N_16302,N_11183,N_10394);
and U16303 (N_16303,N_13252,N_12426);
and U16304 (N_16304,N_13668,N_14293);
nand U16305 (N_16305,N_13934,N_10632);
and U16306 (N_16306,N_14174,N_11926);
nor U16307 (N_16307,N_12256,N_11674);
and U16308 (N_16308,N_14894,N_11580);
nand U16309 (N_16309,N_11331,N_12863);
and U16310 (N_16310,N_14599,N_10123);
nand U16311 (N_16311,N_13280,N_11654);
or U16312 (N_16312,N_10746,N_13761);
nand U16313 (N_16313,N_12859,N_11420);
or U16314 (N_16314,N_12421,N_14408);
or U16315 (N_16315,N_13797,N_12570);
nand U16316 (N_16316,N_10795,N_12238);
or U16317 (N_16317,N_11425,N_11119);
and U16318 (N_16318,N_10171,N_14831);
or U16319 (N_16319,N_10590,N_13997);
and U16320 (N_16320,N_12479,N_12682);
and U16321 (N_16321,N_11340,N_11778);
or U16322 (N_16322,N_10449,N_13047);
nor U16323 (N_16323,N_12674,N_12721);
nand U16324 (N_16324,N_14085,N_14689);
nor U16325 (N_16325,N_14372,N_10320);
nand U16326 (N_16326,N_14609,N_11597);
and U16327 (N_16327,N_13618,N_13901);
and U16328 (N_16328,N_13283,N_14279);
nor U16329 (N_16329,N_14473,N_12845);
or U16330 (N_16330,N_14475,N_11559);
or U16331 (N_16331,N_13925,N_13025);
or U16332 (N_16332,N_12360,N_13803);
nand U16333 (N_16333,N_13876,N_14815);
or U16334 (N_16334,N_10337,N_10613);
nand U16335 (N_16335,N_14192,N_12731);
or U16336 (N_16336,N_12575,N_11701);
nand U16337 (N_16337,N_10297,N_14223);
and U16338 (N_16338,N_12833,N_11914);
nor U16339 (N_16339,N_12612,N_10351);
and U16340 (N_16340,N_14859,N_13271);
or U16341 (N_16341,N_13454,N_13077);
or U16342 (N_16342,N_12564,N_12837);
nand U16343 (N_16343,N_10917,N_14050);
and U16344 (N_16344,N_14434,N_13802);
nor U16345 (N_16345,N_14893,N_14970);
nand U16346 (N_16346,N_11421,N_12266);
or U16347 (N_16347,N_10700,N_14632);
nand U16348 (N_16348,N_12734,N_10269);
nor U16349 (N_16349,N_12381,N_12078);
and U16350 (N_16350,N_11153,N_14628);
and U16351 (N_16351,N_13192,N_11076);
or U16352 (N_16352,N_14545,N_13731);
nor U16353 (N_16353,N_12337,N_11261);
and U16354 (N_16354,N_10169,N_11325);
nor U16355 (N_16355,N_13537,N_13123);
nor U16356 (N_16356,N_14202,N_14489);
nand U16357 (N_16357,N_11367,N_13152);
or U16358 (N_16358,N_11581,N_12281);
nor U16359 (N_16359,N_12434,N_14364);
or U16360 (N_16360,N_11154,N_10887);
nor U16361 (N_16361,N_10648,N_13725);
nand U16362 (N_16362,N_14533,N_14946);
nor U16363 (N_16363,N_13517,N_12633);
or U16364 (N_16364,N_13566,N_12618);
or U16365 (N_16365,N_14969,N_11058);
nand U16366 (N_16366,N_10834,N_13753);
or U16367 (N_16367,N_11233,N_10362);
or U16368 (N_16368,N_12070,N_12739);
nand U16369 (N_16369,N_14136,N_14878);
nor U16370 (N_16370,N_14196,N_12474);
xnor U16371 (N_16371,N_11464,N_11031);
and U16372 (N_16372,N_14936,N_12393);
nor U16373 (N_16373,N_13824,N_10984);
nor U16374 (N_16374,N_12991,N_12749);
nor U16375 (N_16375,N_13186,N_13631);
nand U16376 (N_16376,N_14438,N_14253);
and U16377 (N_16377,N_11777,N_14093);
nand U16378 (N_16378,N_14110,N_12846);
or U16379 (N_16379,N_14289,N_13576);
or U16380 (N_16380,N_12219,N_13000);
nor U16381 (N_16381,N_10285,N_10644);
or U16382 (N_16382,N_11626,N_14480);
nor U16383 (N_16383,N_10716,N_14073);
nand U16384 (N_16384,N_12259,N_13178);
and U16385 (N_16385,N_12270,N_13986);
nand U16386 (N_16386,N_10743,N_10390);
nand U16387 (N_16387,N_12048,N_13784);
nand U16388 (N_16388,N_11355,N_13671);
nor U16389 (N_16389,N_14742,N_13307);
xor U16390 (N_16390,N_14482,N_14178);
and U16391 (N_16391,N_12976,N_13052);
or U16392 (N_16392,N_13662,N_11403);
and U16393 (N_16393,N_13692,N_11249);
or U16394 (N_16394,N_14639,N_12449);
nor U16395 (N_16395,N_11165,N_13814);
nand U16396 (N_16396,N_12643,N_10799);
or U16397 (N_16397,N_11027,N_12826);
nand U16398 (N_16398,N_14903,N_13640);
or U16399 (N_16399,N_13854,N_13349);
and U16400 (N_16400,N_14026,N_11376);
nand U16401 (N_16401,N_14466,N_10902);
nor U16402 (N_16402,N_10106,N_11065);
xor U16403 (N_16403,N_11659,N_13913);
xnor U16404 (N_16404,N_10843,N_13472);
nor U16405 (N_16405,N_11518,N_14133);
nand U16406 (N_16406,N_12797,N_13932);
and U16407 (N_16407,N_13790,N_14317);
xnor U16408 (N_16408,N_11992,N_13035);
or U16409 (N_16409,N_11677,N_11016);
or U16410 (N_16410,N_11118,N_12283);
or U16411 (N_16411,N_14264,N_14693);
xnor U16412 (N_16412,N_13140,N_10100);
nor U16413 (N_16413,N_13644,N_14643);
nand U16414 (N_16414,N_11395,N_12913);
nand U16415 (N_16415,N_14069,N_14681);
or U16416 (N_16416,N_13531,N_12396);
nor U16417 (N_16417,N_12201,N_12729);
and U16418 (N_16418,N_10062,N_10535);
nand U16419 (N_16419,N_12765,N_10369);
or U16420 (N_16420,N_13425,N_11958);
or U16421 (N_16421,N_10796,N_11598);
xor U16422 (N_16422,N_10360,N_13984);
xor U16423 (N_16423,N_10823,N_14915);
or U16424 (N_16424,N_10417,N_11607);
nor U16425 (N_16425,N_11237,N_10312);
nand U16426 (N_16426,N_11348,N_13711);
or U16427 (N_16427,N_11278,N_13856);
xor U16428 (N_16428,N_10860,N_11913);
or U16429 (N_16429,N_13911,N_12346);
nor U16430 (N_16430,N_13183,N_14385);
nand U16431 (N_16431,N_14524,N_13528);
or U16432 (N_16432,N_13043,N_10643);
nor U16433 (N_16433,N_10402,N_11009);
and U16434 (N_16434,N_14214,N_12756);
and U16435 (N_16435,N_11493,N_12866);
nor U16436 (N_16436,N_11669,N_14025);
nand U16437 (N_16437,N_14172,N_13767);
or U16438 (N_16438,N_14726,N_12422);
nor U16439 (N_16439,N_11505,N_12324);
and U16440 (N_16440,N_10710,N_11114);
or U16441 (N_16441,N_10874,N_11959);
or U16442 (N_16442,N_13608,N_13809);
and U16443 (N_16443,N_14687,N_12755);
nand U16444 (N_16444,N_10300,N_11109);
or U16445 (N_16445,N_13500,N_13139);
and U16446 (N_16446,N_12857,N_13147);
and U16447 (N_16447,N_10913,N_12255);
or U16448 (N_16448,N_11151,N_10646);
nand U16449 (N_16449,N_14054,N_14369);
nand U16450 (N_16450,N_10869,N_12960);
or U16451 (N_16451,N_12828,N_11871);
nand U16452 (N_16452,N_13886,N_11862);
nand U16453 (N_16453,N_12777,N_12504);
and U16454 (N_16454,N_10704,N_13295);
nand U16455 (N_16455,N_14647,N_11886);
or U16456 (N_16456,N_11578,N_11283);
and U16457 (N_16457,N_11944,N_11281);
or U16458 (N_16458,N_12627,N_12366);
and U16459 (N_16459,N_10318,N_12090);
or U16460 (N_16460,N_10954,N_12321);
xnor U16461 (N_16461,N_11999,N_14751);
nand U16462 (N_16462,N_14861,N_10410);
or U16463 (N_16463,N_11256,N_13967);
nor U16464 (N_16464,N_12796,N_13848);
nor U16465 (N_16465,N_14977,N_10664);
nand U16466 (N_16466,N_11480,N_10329);
nor U16467 (N_16467,N_14236,N_14212);
nor U16468 (N_16468,N_11415,N_14691);
nand U16469 (N_16469,N_14577,N_14452);
or U16470 (N_16470,N_13998,N_14314);
nor U16471 (N_16471,N_11981,N_14313);
or U16472 (N_16472,N_14819,N_14189);
nor U16473 (N_16473,N_11483,N_11561);
nand U16474 (N_16474,N_10183,N_14308);
nor U16475 (N_16475,N_11136,N_14490);
and U16476 (N_16476,N_13209,N_11855);
nand U16477 (N_16477,N_10041,N_13115);
nand U16478 (N_16478,N_10181,N_10739);
nor U16479 (N_16479,N_13673,N_10875);
or U16480 (N_16480,N_10296,N_11899);
nor U16481 (N_16481,N_13437,N_14261);
or U16482 (N_16482,N_11650,N_11292);
nor U16483 (N_16483,N_11263,N_10637);
nor U16484 (N_16484,N_10078,N_11185);
or U16485 (N_16485,N_10529,N_13768);
nor U16486 (N_16486,N_14428,N_11248);
nand U16487 (N_16487,N_10682,N_10147);
and U16488 (N_16488,N_11302,N_12716);
and U16489 (N_16489,N_14788,N_11739);
nor U16490 (N_16490,N_12250,N_12966);
or U16491 (N_16491,N_11713,N_12031);
and U16492 (N_16492,N_13949,N_10818);
or U16493 (N_16493,N_10348,N_10685);
or U16494 (N_16494,N_12539,N_14593);
and U16495 (N_16495,N_11393,N_13113);
nor U16496 (N_16496,N_12819,N_12300);
and U16497 (N_16497,N_12225,N_13044);
nor U16498 (N_16498,N_14271,N_10905);
or U16499 (N_16499,N_10759,N_13871);
and U16500 (N_16500,N_12163,N_11209);
nor U16501 (N_16501,N_13509,N_10442);
or U16502 (N_16502,N_12469,N_13995);
or U16503 (N_16503,N_10757,N_13549);
nor U16504 (N_16504,N_13014,N_14899);
and U16505 (N_16505,N_14284,N_11512);
or U16506 (N_16506,N_11196,N_12358);
nor U16507 (N_16507,N_12920,N_10258);
nor U16508 (N_16508,N_12655,N_11125);
nor U16509 (N_16509,N_14141,N_13885);
xor U16510 (N_16510,N_12944,N_14733);
nand U16511 (N_16511,N_10356,N_12372);
or U16512 (N_16512,N_13799,N_13256);
nand U16513 (N_16513,N_12294,N_12581);
and U16514 (N_16514,N_11414,N_11605);
and U16515 (N_16515,N_11771,N_11766);
nor U16516 (N_16516,N_11055,N_11799);
or U16517 (N_16517,N_14282,N_12774);
or U16518 (N_16518,N_11080,N_11511);
and U16519 (N_16519,N_13553,N_14332);
nor U16520 (N_16520,N_11141,N_10517);
or U16521 (N_16521,N_10108,N_13010);
nand U16522 (N_16522,N_11946,N_12840);
nor U16523 (N_16523,N_12931,N_11050);
and U16524 (N_16524,N_11761,N_12641);
nand U16525 (N_16525,N_11863,N_11791);
or U16526 (N_16526,N_10962,N_13233);
nor U16527 (N_16527,N_13857,N_11015);
nand U16528 (N_16528,N_12139,N_10724);
or U16529 (N_16529,N_12622,N_10696);
or U16530 (N_16530,N_12571,N_12314);
nand U16531 (N_16531,N_11187,N_10153);
nor U16532 (N_16532,N_11434,N_11815);
or U16533 (N_16533,N_10916,N_11919);
nand U16534 (N_16534,N_11147,N_10368);
nand U16535 (N_16535,N_12495,N_11636);
nor U16536 (N_16536,N_13739,N_10987);
or U16537 (N_16537,N_12342,N_10157);
and U16538 (N_16538,N_14047,N_12958);
nand U16539 (N_16539,N_10008,N_13203);
nor U16540 (N_16540,N_11084,N_10056);
nand U16541 (N_16541,N_12623,N_14728);
or U16542 (N_16542,N_10099,N_14705);
nor U16543 (N_16543,N_14739,N_11945);
nand U16544 (N_16544,N_13565,N_13084);
or U16545 (N_16545,N_13681,N_14235);
or U16546 (N_16546,N_11357,N_14395);
or U16547 (N_16547,N_14086,N_14778);
or U16548 (N_16548,N_10928,N_12276);
xnor U16549 (N_16549,N_11971,N_13776);
or U16550 (N_16550,N_14300,N_12233);
nand U16551 (N_16551,N_12503,N_10382);
nor U16552 (N_16552,N_10926,N_10542);
xnor U16553 (N_16553,N_10574,N_11941);
nand U16554 (N_16554,N_11620,N_11691);
or U16555 (N_16555,N_10952,N_10332);
nor U16556 (N_16556,N_14684,N_13841);
nand U16557 (N_16557,N_12136,N_14517);
and U16558 (N_16558,N_13064,N_11311);
and U16559 (N_16559,N_14536,N_12093);
nor U16560 (N_16560,N_12852,N_12788);
nand U16561 (N_16561,N_13330,N_14433);
xnor U16562 (N_16562,N_10684,N_13625);
nand U16563 (N_16563,N_12681,N_13190);
nand U16564 (N_16564,N_10524,N_13729);
or U16565 (N_16565,N_12274,N_10052);
and U16566 (N_16566,N_12349,N_10734);
or U16567 (N_16567,N_10035,N_12198);
nor U16568 (N_16568,N_11722,N_10395);
nor U16569 (N_16569,N_13495,N_14694);
or U16570 (N_16570,N_13574,N_10138);
and U16571 (N_16571,N_11175,N_11515);
and U16572 (N_16572,N_13258,N_10238);
or U16573 (N_16573,N_14367,N_11531);
nor U16574 (N_16574,N_12200,N_14709);
nand U16575 (N_16575,N_14979,N_14762);
nor U16576 (N_16576,N_13605,N_12231);
nand U16577 (N_16577,N_11688,N_13757);
or U16578 (N_16578,N_11901,N_11857);
and U16579 (N_16579,N_11497,N_12287);
and U16580 (N_16580,N_13735,N_11651);
or U16581 (N_16581,N_13157,N_12338);
nor U16582 (N_16582,N_13120,N_10384);
or U16583 (N_16583,N_14135,N_10956);
xor U16584 (N_16584,N_11097,N_10594);
nor U16585 (N_16585,N_11931,N_10092);
nor U16586 (N_16586,N_13515,N_10323);
and U16587 (N_16587,N_13774,N_11500);
and U16588 (N_16588,N_12004,N_14525);
and U16589 (N_16589,N_14351,N_13669);
or U16590 (N_16590,N_14019,N_10139);
or U16591 (N_16591,N_14746,N_10672);
nand U16592 (N_16592,N_13891,N_10735);
nor U16593 (N_16593,N_13994,N_14929);
or U16594 (N_16594,N_11859,N_10811);
nand U16595 (N_16595,N_13061,N_14736);
nand U16596 (N_16596,N_12634,N_13559);
or U16597 (N_16597,N_11454,N_11435);
or U16598 (N_16598,N_10732,N_12836);
or U16599 (N_16599,N_12759,N_14501);
and U16600 (N_16600,N_14012,N_12378);
xor U16601 (N_16601,N_13522,N_10736);
or U16602 (N_16602,N_10085,N_14334);
or U16603 (N_16603,N_14156,N_13386);
xor U16604 (N_16604,N_12524,N_10043);
and U16605 (N_16605,N_14943,N_10800);
and U16606 (N_16606,N_10468,N_12395);
and U16607 (N_16607,N_10775,N_13639);
nor U16608 (N_16608,N_14558,N_10618);
nor U16609 (N_16609,N_11624,N_14286);
and U16610 (N_16610,N_11051,N_10895);
and U16611 (N_16611,N_11071,N_11377);
or U16612 (N_16612,N_11477,N_10896);
nand U16613 (N_16613,N_10728,N_10525);
or U16614 (N_16614,N_11120,N_13873);
or U16615 (N_16615,N_12336,N_13118);
and U16616 (N_16616,N_11332,N_13080);
or U16617 (N_16617,N_11595,N_11388);
or U16618 (N_16618,N_12895,N_11642);
nor U16619 (N_16619,N_11243,N_10151);
and U16620 (N_16620,N_12808,N_13530);
and U16621 (N_16621,N_13714,N_11102);
and U16622 (N_16622,N_13632,N_10287);
or U16623 (N_16623,N_14128,N_13104);
nand U16624 (N_16624,N_11110,N_12905);
nor U16625 (N_16625,N_10712,N_10679);
nor U16626 (N_16626,N_14020,N_12650);
and U16627 (N_16627,N_14035,N_12306);
nor U16628 (N_16628,N_13756,N_12919);
or U16629 (N_16629,N_11087,N_14901);
or U16630 (N_16630,N_11077,N_10460);
and U16631 (N_16631,N_12471,N_13069);
nand U16632 (N_16632,N_12351,N_14391);
and U16633 (N_16633,N_12280,N_13142);
nor U16634 (N_16634,N_13712,N_14839);
nor U16635 (N_16635,N_14151,N_10614);
and U16636 (N_16636,N_11260,N_12590);
nor U16637 (N_16637,N_14775,N_14359);
xor U16638 (N_16638,N_11306,N_13363);
nor U16639 (N_16639,N_11067,N_13748);
or U16640 (N_16640,N_10935,N_14834);
nor U16641 (N_16641,N_10346,N_11895);
or U16642 (N_16642,N_11034,N_11602);
nor U16643 (N_16643,N_10858,N_12884);
and U16644 (N_16644,N_13306,N_11346);
or U16645 (N_16645,N_13101,N_14671);
nand U16646 (N_16646,N_11653,N_12714);
nor U16647 (N_16647,N_10666,N_13906);
nor U16648 (N_16648,N_10458,N_12489);
nand U16649 (N_16649,N_14400,N_14824);
and U16650 (N_16650,N_13480,N_12686);
nor U16651 (N_16651,N_11835,N_10768);
or U16652 (N_16652,N_13422,N_12578);
nor U16653 (N_16653,N_14122,N_14704);
nand U16654 (N_16654,N_13806,N_13296);
nand U16655 (N_16655,N_11228,N_13653);
or U16656 (N_16656,N_11977,N_12659);
xor U16657 (N_16657,N_10006,N_13196);
nand U16658 (N_16658,N_10227,N_10527);
nor U16659 (N_16659,N_13009,N_11131);
and U16660 (N_16660,N_14993,N_13546);
nand U16661 (N_16661,N_12205,N_12678);
nor U16662 (N_16662,N_11916,N_13039);
nor U16663 (N_16663,N_13569,N_14294);
or U16664 (N_16664,N_13097,N_13224);
nand U16665 (N_16665,N_10709,N_11180);
nor U16666 (N_16666,N_13318,N_14997);
nand U16667 (N_16667,N_11061,N_14348);
nor U16668 (N_16668,N_14652,N_12407);
and U16669 (N_16669,N_13749,N_13159);
nand U16670 (N_16670,N_10771,N_12096);
nand U16671 (N_16671,N_10551,N_10444);
nand U16672 (N_16672,N_10263,N_11018);
xnor U16673 (N_16673,N_11345,N_10094);
and U16674 (N_16674,N_14683,N_12054);
or U16675 (N_16675,N_11402,N_10863);
or U16676 (N_16676,N_10027,N_13879);
and U16677 (N_16677,N_14362,N_10203);
nor U16678 (N_16678,N_13327,N_13958);
or U16679 (N_16679,N_12762,N_14170);
or U16680 (N_16680,N_12491,N_14620);
nor U16681 (N_16681,N_10856,N_14817);
xnor U16682 (N_16682,N_11270,N_13155);
and U16683 (N_16683,N_13154,N_13031);
or U16684 (N_16684,N_10255,N_14375);
nor U16685 (N_16685,N_10651,N_12086);
nand U16686 (N_16686,N_11225,N_11661);
and U16687 (N_16687,N_13136,N_13523);
nor U16688 (N_16688,N_11637,N_14220);
and U16689 (N_16689,N_13927,N_10890);
nor U16690 (N_16690,N_13896,N_11190);
and U16691 (N_16691,N_11904,N_12034);
nor U16692 (N_16692,N_12215,N_10652);
and U16693 (N_16693,N_13490,N_12317);
and U16694 (N_16694,N_10491,N_13648);
or U16695 (N_16695,N_14862,N_12282);
and U16696 (N_16696,N_11142,N_12235);
or U16697 (N_16697,N_13095,N_10788);
or U16698 (N_16698,N_14591,N_13953);
nor U16699 (N_16699,N_12672,N_10610);
or U16700 (N_16700,N_12220,N_12640);
and U16701 (N_16701,N_10239,N_12290);
or U16702 (N_16702,N_12308,N_12416);
or U16703 (N_16703,N_12563,N_13971);
nand U16704 (N_16704,N_12941,N_12645);
nand U16705 (N_16705,N_14256,N_11514);
or U16706 (N_16706,N_11262,N_13364);
or U16707 (N_16707,N_12815,N_11878);
nor U16708 (N_16708,N_11665,N_11394);
nand U16709 (N_16709,N_12143,N_12246);
or U16710 (N_16710,N_10156,N_12965);
or U16711 (N_16711,N_13475,N_11888);
and U16712 (N_16712,N_14800,N_11720);
xor U16713 (N_16713,N_10150,N_11495);
nand U16714 (N_16714,N_12954,N_14793);
and U16715 (N_16715,N_13685,N_10014);
or U16716 (N_16716,N_14697,N_13699);
nand U16717 (N_16717,N_13405,N_14829);
or U16718 (N_16718,N_10256,N_14779);
nand U16719 (N_16719,N_11801,N_10291);
or U16720 (N_16720,N_11369,N_11587);
or U16721 (N_16721,N_11397,N_14852);
nand U16722 (N_16722,N_14951,N_11251);
and U16723 (N_16723,N_13960,N_13292);
and U16724 (N_16724,N_10111,N_13112);
nand U16725 (N_16725,N_13324,N_11741);
nor U16726 (N_16726,N_12720,N_11083);
nor U16727 (N_16727,N_12929,N_11890);
nand U16728 (N_16728,N_11276,N_11700);
nand U16729 (N_16729,N_11986,N_10339);
nand U16730 (N_16730,N_14338,N_14199);
nand U16731 (N_16731,N_14460,N_14520);
or U16732 (N_16732,N_14407,N_14259);
nand U16733 (N_16733,N_13643,N_11299);
nor U16734 (N_16734,N_11973,N_14828);
or U16735 (N_16735,N_13532,N_12155);
or U16736 (N_16736,N_13775,N_14881);
or U16737 (N_16737,N_13921,N_14527);
nand U16738 (N_16738,N_13596,N_13585);
and U16739 (N_16739,N_10281,N_11616);
nor U16740 (N_16740,N_13336,N_10409);
and U16741 (N_16741,N_14919,N_13649);
or U16742 (N_16742,N_11742,N_10989);
and U16743 (N_16743,N_14774,N_10898);
nand U16744 (N_16744,N_13992,N_10894);
or U16745 (N_16745,N_10495,N_14528);
or U16746 (N_16746,N_11300,N_12410);
nor U16747 (N_16747,N_14702,N_14099);
and U16748 (N_16748,N_11020,N_14402);
and U16749 (N_16749,N_14380,N_11952);
or U16750 (N_16750,N_11563,N_10665);
nor U16751 (N_16751,N_10484,N_13265);
or U16752 (N_16752,N_11708,N_10626);
nand U16753 (N_16753,N_11333,N_10228);
or U16754 (N_16754,N_14412,N_13188);
or U16755 (N_16755,N_14896,N_11987);
and U16756 (N_16756,N_11847,N_12428);
nor U16757 (N_16757,N_11356,N_10831);
and U16758 (N_16758,N_12100,N_13319);
and U16759 (N_16759,N_14868,N_12214);
nand U16760 (N_16760,N_13862,N_13049);
nor U16761 (N_16761,N_13402,N_13135);
nand U16762 (N_16762,N_13720,N_13092);
and U16763 (N_16763,N_12052,N_14925);
nor U16764 (N_16764,N_12041,N_13388);
xnor U16765 (N_16765,N_11127,N_13305);
or U16766 (N_16766,N_13194,N_13452);
nand U16767 (N_16767,N_10930,N_12906);
and U16768 (N_16768,N_10570,N_11312);
or U16769 (N_16769,N_12363,N_12310);
and U16770 (N_16770,N_13744,N_10631);
and U16771 (N_16771,N_14542,N_11929);
nand U16772 (N_16772,N_14941,N_14911);
nand U16773 (N_16773,N_10974,N_13444);
and U16774 (N_16774,N_14916,N_10707);
nand U16775 (N_16775,N_11424,N_14307);
nor U16776 (N_16776,N_13389,N_14990);
nand U16777 (N_16777,N_12896,N_11117);
nor U16778 (N_16778,N_11978,N_10268);
and U16779 (N_16779,N_13016,N_14590);
and U16780 (N_16780,N_14272,N_14245);
and U16781 (N_16781,N_11685,N_14804);
nand U16782 (N_16782,N_13957,N_10377);
and U16783 (N_16783,N_12985,N_10469);
and U16784 (N_16784,N_13385,N_14251);
or U16785 (N_16785,N_11232,N_14822);
and U16786 (N_16786,N_11732,N_11579);
nor U16787 (N_16787,N_10815,N_10036);
nor U16788 (N_16788,N_12387,N_11772);
nor U16789 (N_16789,N_10765,N_10580);
and U16790 (N_16790,N_13227,N_10502);
nand U16791 (N_16791,N_12003,N_14960);
nand U16792 (N_16792,N_13387,N_14690);
and U16793 (N_16793,N_10420,N_10658);
and U16794 (N_16794,N_11253,N_11328);
nor U16795 (N_16795,N_13898,N_13421);
and U16796 (N_16796,N_10675,N_11787);
or U16797 (N_16797,N_12946,N_13964);
nor U16798 (N_16798,N_13199,N_13599);
and U16799 (N_16799,N_12855,N_12223);
and U16800 (N_16800,N_13087,N_13524);
and U16801 (N_16801,N_12752,N_13807);
or U16802 (N_16802,N_14467,N_11557);
nor U16803 (N_16803,N_11643,N_11011);
or U16804 (N_16804,N_13242,N_13267);
nand U16805 (N_16805,N_10051,N_14092);
nand U16806 (N_16806,N_10881,N_13907);
and U16807 (N_16807,N_10218,N_13294);
and U16808 (N_16808,N_14770,N_13675);
and U16809 (N_16809,N_13592,N_11272);
or U16810 (N_16810,N_14914,N_14496);
nand U16811 (N_16811,N_14743,N_13899);
and U16812 (N_16812,N_11571,N_10776);
and U16813 (N_16813,N_13601,N_14518);
nor U16814 (N_16814,N_13390,N_11760);
nor U16815 (N_16815,N_13451,N_12915);
nor U16816 (N_16816,N_13622,N_11266);
or U16817 (N_16817,N_10587,N_12301);
and U16818 (N_16818,N_12843,N_13686);
and U16819 (N_16819,N_11666,N_11538);
nand U16820 (N_16820,N_10134,N_10841);
nand U16821 (N_16821,N_14782,N_14656);
or U16822 (N_16822,N_12900,N_11326);
nand U16823 (N_16823,N_13875,N_11537);
or U16824 (N_16824,N_12589,N_13301);
nor U16825 (N_16825,N_10720,N_10231);
or U16826 (N_16826,N_11026,N_14126);
and U16827 (N_16827,N_11490,N_12647);
nor U16828 (N_16828,N_14523,N_11530);
nand U16829 (N_16829,N_13443,N_12804);
or U16830 (N_16830,N_11150,N_12105);
or U16831 (N_16831,N_10885,N_11502);
nor U16832 (N_16832,N_10354,N_12963);
and U16833 (N_16833,N_10168,N_10957);
nand U16834 (N_16834,N_12600,N_12313);
nand U16835 (N_16835,N_14571,N_13831);
nand U16836 (N_16836,N_13655,N_12477);
and U16837 (N_16837,N_11005,N_14924);
nor U16838 (N_16838,N_10554,N_12497);
nand U16839 (N_16839,N_12073,N_13595);
xnor U16840 (N_16840,N_11222,N_12341);
nand U16841 (N_16841,N_10680,N_12738);
nand U16842 (N_16842,N_12355,N_14106);
or U16843 (N_16843,N_12368,N_13019);
xor U16844 (N_16844,N_14669,N_14592);
nand U16845 (N_16845,N_10120,N_11100);
nand U16846 (N_16846,N_11746,N_14432);
and U16847 (N_16847,N_11628,N_14125);
or U16848 (N_16848,N_10687,N_11133);
and U16849 (N_16849,N_11113,N_14569);
nor U16850 (N_16850,N_12026,N_13429);
or U16851 (N_16851,N_13424,N_12361);
or U16852 (N_16852,N_10249,N_10075);
or U16853 (N_16853,N_11447,N_11614);
nor U16854 (N_16854,N_10033,N_11112);
nor U16855 (N_16855,N_11170,N_13661);
nor U16856 (N_16856,N_10357,N_14003);
nand U16857 (N_16857,N_13539,N_12569);
nor U16858 (N_16858,N_13304,N_11107);
or U16859 (N_16859,N_12698,N_11631);
or U16860 (N_16860,N_12204,N_10690);
nand U16861 (N_16861,N_14630,N_11736);
or U16862 (N_16862,N_11730,N_13750);
nor U16863 (N_16863,N_14747,N_12651);
and U16864 (N_16864,N_12451,N_11762);
or U16865 (N_16865,N_14070,N_13961);
and U16866 (N_16866,N_14564,N_14766);
nor U16867 (N_16867,N_11922,N_11903);
and U16868 (N_16868,N_11171,N_14451);
xnor U16869 (N_16869,N_11240,N_10911);
nand U16870 (N_16870,N_10087,N_14152);
nor U16871 (N_16871,N_12299,N_13518);
nor U16872 (N_16872,N_13132,N_11298);
nor U16873 (N_16873,N_12853,N_13438);
or U16874 (N_16874,N_13829,N_11089);
or U16875 (N_16875,N_14445,N_10160);
nand U16876 (N_16876,N_14585,N_13733);
nor U16877 (N_16877,N_13395,N_10021);
and U16878 (N_16878,N_13838,N_11672);
nor U16879 (N_16879,N_12297,N_10034);
nand U16880 (N_16880,N_14874,N_12134);
nor U16881 (N_16881,N_14232,N_14225);
nand U16882 (N_16882,N_10340,N_11930);
nor U16883 (N_16883,N_13431,N_10154);
or U16884 (N_16884,N_10376,N_12662);
nor U16885 (N_16885,N_10922,N_13893);
nand U16886 (N_16886,N_11314,N_12545);
and U16887 (N_16887,N_12935,N_10383);
nor U16888 (N_16888,N_13184,N_10854);
and U16889 (N_16889,N_14526,N_14897);
xnor U16890 (N_16890,N_10392,N_14357);
and U16891 (N_16891,N_13339,N_14511);
nand U16892 (N_16892,N_13130,N_12419);
or U16893 (N_16893,N_14574,N_10539);
or U16894 (N_16894,N_14329,N_10726);
nand U16895 (N_16895,N_12642,N_11066);
and U16896 (N_16896,N_12165,N_11371);
or U16897 (N_16897,N_13944,N_13542);
or U16898 (N_16898,N_11980,N_14584);
or U16899 (N_16899,N_13413,N_13506);
nor U16900 (N_16900,N_10286,N_10109);
or U16901 (N_16901,N_12751,N_14297);
nor U16902 (N_16902,N_10583,N_14015);
nand U16903 (N_16903,N_14390,N_11013);
nor U16904 (N_16904,N_12344,N_14166);
nand U16905 (N_16905,N_10175,N_12224);
nand U16906 (N_16906,N_11224,N_11014);
or U16907 (N_16907,N_13033,N_11038);
nor U16908 (N_16908,N_11572,N_14744);
or U16909 (N_16909,N_12974,N_11998);
or U16910 (N_16910,N_14550,N_11304);
nor U16911 (N_16911,N_10891,N_10589);
and U16912 (N_16912,N_13815,N_14305);
nor U16913 (N_16913,N_12775,N_10371);
and U16914 (N_16914,N_14349,N_11056);
nor U16915 (N_16915,N_13534,N_14423);
nand U16916 (N_16916,N_10754,N_10657);
nand U16917 (N_16917,N_13738,N_10976);
and U16918 (N_16918,N_11359,N_11433);
or U16919 (N_16919,N_13647,N_11194);
nor U16920 (N_16920,N_10400,N_14486);
nor U16921 (N_16921,N_12400,N_11029);
nand U16922 (N_16922,N_13350,N_13603);
nand U16923 (N_16923,N_10422,N_10016);
and U16924 (N_16924,N_11466,N_10932);
nand U16925 (N_16925,N_10821,N_12956);
nand U16926 (N_16926,N_12076,N_10552);
nand U16927 (N_16927,N_11809,N_11947);
and U16928 (N_16928,N_12706,N_13488);
or U16929 (N_16929,N_11818,N_10993);
and U16930 (N_16930,N_14992,N_11137);
or U16931 (N_16931,N_12020,N_11875);
nand U16932 (N_16932,N_14937,N_11010);
nor U16933 (N_16933,N_12332,N_13514);
or U16934 (N_16934,N_12433,N_14679);
nor U16935 (N_16935,N_12369,N_12129);
nand U16936 (N_16936,N_11629,N_13544);
and U16937 (N_16937,N_10315,N_12170);
nor U16938 (N_16938,N_14884,N_13221);
nor U16939 (N_16939,N_13977,N_10819);
and U16940 (N_16940,N_14799,N_12842);
nand U16941 (N_16941,N_10947,N_12726);
nand U16942 (N_16942,N_13800,N_12397);
and U16943 (N_16943,N_11130,N_11482);
and U16944 (N_16944,N_14920,N_11918);
or U16945 (N_16945,N_12661,N_12847);
nand U16946 (N_16946,N_11526,N_11536);
nor U16947 (N_16947,N_12740,N_12520);
nand U16948 (N_16948,N_11844,N_12792);
xnor U16949 (N_16949,N_13600,N_14544);
and U16950 (N_16950,N_13315,N_12829);
or U16951 (N_16951,N_11216,N_13426);
or U16952 (N_16952,N_14755,N_12398);
nand U16953 (N_16953,N_11452,N_10307);
or U16954 (N_16954,N_10011,N_11640);
or U16955 (N_16955,N_10189,N_10511);
and U16956 (N_16956,N_12117,N_14203);
and U16957 (N_16957,N_12687,N_11234);
or U16958 (N_16958,N_14510,N_10428);
or U16959 (N_16959,N_12776,N_13679);
or U16960 (N_16960,N_12121,N_12183);
nand U16961 (N_16961,N_10506,N_11757);
nand U16962 (N_16962,N_10803,N_11795);
and U16963 (N_16963,N_10049,N_11072);
nor U16964 (N_16964,N_12992,N_11303);
nand U16965 (N_16965,N_11274,N_14053);
nor U16966 (N_16966,N_11586,N_11936);
or U16967 (N_16967,N_14502,N_11188);
or U16968 (N_16968,N_10433,N_13713);
nor U16969 (N_16969,N_12619,N_12399);
nor U16970 (N_16970,N_10244,N_13740);
or U16971 (N_16971,N_14882,N_11967);
or U16972 (N_16972,N_11754,N_13975);
nor U16973 (N_16973,N_14717,N_13239);
nand U16974 (N_16974,N_10770,N_14065);
nand U16975 (N_16975,N_10778,N_12761);
nand U16976 (N_16976,N_11364,N_12029);
or U16977 (N_16977,N_11288,N_10616);
or U16978 (N_16978,N_10343,N_13060);
nor U16979 (N_16979,N_13434,N_13200);
and U16980 (N_16980,N_13991,N_11995);
nor U16981 (N_16981,N_12793,N_10998);
and U16982 (N_16982,N_13710,N_12251);
or U16983 (N_16983,N_14663,N_14137);
nand U16984 (N_16984,N_13191,N_13570);
xor U16985 (N_16985,N_14818,N_10113);
nand U16986 (N_16986,N_13942,N_14618);
and U16987 (N_16987,N_10575,N_11208);
and U16988 (N_16988,N_10714,N_10093);
nand U16989 (N_16989,N_13923,N_14907);
and U16990 (N_16990,N_14552,N_11961);
or U16991 (N_16991,N_14801,N_10434);
nor U16992 (N_16992,N_11920,N_12330);
and U16993 (N_16993,N_13502,N_11057);
nand U16994 (N_16994,N_12646,N_14900);
nand U16995 (N_16995,N_10708,N_12174);
and U16996 (N_16996,N_11608,N_13999);
or U16997 (N_16997,N_12688,N_11883);
or U16998 (N_16998,N_13983,N_14509);
nand U16999 (N_16999,N_12359,N_10252);
and U17000 (N_17000,N_13436,N_11695);
nand U17001 (N_17001,N_14327,N_10772);
or U17002 (N_17002,N_11521,N_13660);
xor U17003 (N_17003,N_12540,N_13850);
nand U17004 (N_17004,N_14966,N_11822);
nand U17005 (N_17005,N_14162,N_12271);
nand U17006 (N_17006,N_14888,N_11455);
nor U17007 (N_17007,N_10427,N_12146);
or U17008 (N_17008,N_10633,N_13114);
nand U17009 (N_17009,N_11569,N_14665);
nor U17010 (N_17010,N_11856,N_13642);
and U17011 (N_17011,N_10838,N_10851);
nand U17012 (N_17012,N_10640,N_14640);
and U17013 (N_17013,N_11997,N_10070);
or U17014 (N_17014,N_13459,N_13947);
nand U17015 (N_17015,N_14792,N_14503);
and U17016 (N_17016,N_13963,N_13038);
nand U17017 (N_17017,N_10582,N_14455);
nor U17018 (N_17018,N_10146,N_10808);
nor U17019 (N_17019,N_14205,N_10695);
nand U17020 (N_17020,N_11291,N_12420);
and U17021 (N_17021,N_10749,N_11872);
or U17022 (N_17022,N_13237,N_13119);
nand U17023 (N_17023,N_10927,N_13440);
or U17024 (N_17024,N_13493,N_14780);
or U17025 (N_17025,N_12475,N_10745);
or U17026 (N_17026,N_13702,N_11765);
or U17027 (N_17027,N_12582,N_13099);
nor U17028 (N_17028,N_12586,N_14514);
and U17029 (N_17029,N_10055,N_12470);
and U17030 (N_17030,N_11758,N_11069);
or U17031 (N_17031,N_13210,N_10513);
nor U17032 (N_17032,N_12312,N_11386);
or U17033 (N_17033,N_13497,N_12116);
and U17034 (N_17034,N_13584,N_11380);
or U17035 (N_17035,N_13696,N_10873);
and U17036 (N_17036,N_13745,N_14363);
and U17037 (N_17037,N_14487,N_11128);
and U17038 (N_17038,N_13313,N_12119);
or U17039 (N_17039,N_13133,N_11848);
or U17040 (N_17040,N_13219,N_10451);
nor U17041 (N_17041,N_10991,N_14377);
or U17042 (N_17042,N_13762,N_12887);
and U17043 (N_17043,N_13150,N_14448);
nor U17044 (N_17044,N_12127,N_10237);
and U17045 (N_17045,N_12302,N_10609);
nand U17046 (N_17046,N_14078,N_12923);
nor U17047 (N_17047,N_12957,N_10024);
nor U17048 (N_17048,N_11820,N_14568);
and U17049 (N_17049,N_12525,N_11028);
and U17050 (N_17050,N_13579,N_11115);
or U17051 (N_17051,N_11568,N_11413);
and U17052 (N_17052,N_10316,N_12697);
and U17053 (N_17053,N_10435,N_13071);
or U17054 (N_17054,N_13929,N_12331);
or U17055 (N_17055,N_12316,N_13505);
nand U17056 (N_17056,N_10791,N_12011);
nor U17057 (N_17057,N_13312,N_14180);
nor U17058 (N_17058,N_11250,N_11155);
nand U17059 (N_17059,N_12632,N_14957);
and U17060 (N_17060,N_14321,N_12145);
nand U17061 (N_17061,N_12785,N_12304);
and U17062 (N_17062,N_12490,N_13526);
or U17063 (N_17063,N_10876,N_14474);
nand U17064 (N_17064,N_11548,N_13636);
or U17065 (N_17065,N_14555,N_11252);
xor U17066 (N_17066,N_13742,N_10396);
or U17067 (N_17067,N_14392,N_12042);
and U17068 (N_17068,N_11203,N_12710);
nor U17069 (N_17069,N_14469,N_14154);
and U17070 (N_17070,N_14129,N_14239);
nor U17071 (N_17071,N_12719,N_11940);
nand U17072 (N_17072,N_10560,N_14962);
nand U17073 (N_17073,N_13471,N_11752);
nand U17074 (N_17074,N_11019,N_12555);
and U17075 (N_17075,N_11989,N_10797);
nand U17076 (N_17076,N_10379,N_11247);
and U17077 (N_17077,N_14097,N_12062);
or U17078 (N_17078,N_10986,N_10725);
or U17079 (N_17079,N_11925,N_14895);
nand U17080 (N_17080,N_14749,N_14530);
and U17081 (N_17081,N_13449,N_12383);
nand U17082 (N_17082,N_13996,N_12472);
xor U17083 (N_17083,N_13074,N_13419);
or U17084 (N_17084,N_10306,N_14080);
and U17085 (N_17085,N_12059,N_10186);
and U17086 (N_17086,N_11126,N_13003);
and U17087 (N_17087,N_11468,N_10265);
xnor U17088 (N_17088,N_13002,N_10820);
nand U17089 (N_17089,N_13722,N_14898);
and U17090 (N_17090,N_10198,N_11621);
and U17091 (N_17091,N_10619,N_12817);
or U17092 (N_17092,N_12039,N_11206);
and U17093 (N_17093,N_13878,N_11186);
or U17094 (N_17094,N_14464,N_11682);
nand U17095 (N_17095,N_10313,N_10867);
nor U17096 (N_17096,N_14230,N_14676);
or U17097 (N_17097,N_12532,N_13284);
xnor U17098 (N_17098,N_10207,N_11060);
and U17099 (N_17099,N_10558,N_11826);
or U17100 (N_17100,N_10521,N_13779);
or U17101 (N_17101,N_10206,N_13782);
nand U17102 (N_17102,N_13311,N_10534);
or U17103 (N_17103,N_13230,N_14857);
or U17104 (N_17104,N_13216,N_10279);
nand U17105 (N_17105,N_10804,N_14386);
or U17106 (N_17106,N_12823,N_14783);
nand U17107 (N_17107,N_10568,N_10752);
or U17108 (N_17108,N_12454,N_10077);
or U17109 (N_17109,N_13859,N_11655);
nor U17110 (N_17110,N_10748,N_12190);
nor U17111 (N_17111,N_12362,N_11428);
nand U17112 (N_17112,N_12588,N_11591);
nor U17113 (N_17113,N_13520,N_13817);
nor U17114 (N_17114,N_11528,N_13939);
and U17115 (N_17115,N_12972,N_14287);
nor U17116 (N_17116,N_11912,N_14201);
or U17117 (N_17117,N_14521,N_14168);
or U17118 (N_17118,N_11323,N_10722);
and U17119 (N_17119,N_12723,N_13987);
nor U17120 (N_17120,N_14773,N_12453);
or U17121 (N_17121,N_13008,N_14776);
or U17122 (N_17122,N_13232,N_12114);
or U17123 (N_17123,N_14310,N_10606);
xor U17124 (N_17124,N_13980,N_11564);
and U17125 (N_17125,N_11082,N_11070);
nor U17126 (N_17126,N_12554,N_13380);
and U17127 (N_17127,N_11550,N_11698);
and U17128 (N_17128,N_14344,N_10599);
xnor U17129 (N_17129,N_11445,N_12854);
or U17130 (N_17130,N_12781,N_13082);
nand U17131 (N_17131,N_11663,N_11885);
nand U17132 (N_17132,N_14917,N_14187);
nor U17133 (N_17133,N_14138,N_14649);
and U17134 (N_17134,N_13096,N_10355);
nand U17135 (N_17135,N_14091,N_13985);
nor U17136 (N_17136,N_11798,N_13334);
or U17137 (N_17137,N_11184,N_11817);
nand U17138 (N_17138,N_11205,N_10251);
nor U17139 (N_17139,N_11854,N_10322);
nand U17140 (N_17140,N_11910,N_12814);
or U17141 (N_17141,N_11309,N_11592);
and U17142 (N_17142,N_11972,N_12943);
and U17143 (N_17143,N_11442,N_14931);
nor U17144 (N_17144,N_13670,N_11632);
nand U17145 (N_17145,N_12172,N_12013);
xnor U17146 (N_17146,N_14554,N_11352);
nor U17147 (N_17147,N_11446,N_10785);
nand U17148 (N_17148,N_10305,N_11613);
nor U17149 (N_17149,N_12177,N_11392);
nand U17150 (N_17150,N_14614,N_12019);
nand U17151 (N_17151,N_14037,N_11549);
nand U17152 (N_17152,N_10901,N_11350);
nor U17153 (N_17153,N_13889,N_12986);
nand U17154 (N_17154,N_12464,N_13695);
nand U17155 (N_17155,N_13904,N_10003);
nor U17156 (N_17156,N_13948,N_12109);
and U17157 (N_17157,N_11819,N_12429);
nor U17158 (N_17158,N_13863,N_10476);
nand U17159 (N_17159,N_13837,N_10217);
nor U17160 (N_17160,N_13254,N_14587);
and U17161 (N_17161,N_11715,N_10353);
nor U17162 (N_17162,N_12657,N_12987);
nor U17163 (N_17163,N_12526,N_11174);
nor U17164 (N_17164,N_12967,N_12559);
nor U17165 (N_17165,N_10889,N_12171);
or U17166 (N_17166,N_10275,N_12024);
nand U17167 (N_17167,N_13018,N_14032);
xor U17168 (N_17168,N_11976,N_10350);
nand U17169 (N_17169,N_13448,N_14624);
nand U17170 (N_17170,N_12384,N_10615);
nand U17171 (N_17171,N_13020,N_12118);
nor U17172 (N_17172,N_12615,N_11436);
and U17173 (N_17173,N_14409,N_10787);
or U17174 (N_17174,N_14677,N_14227);
nor U17175 (N_17175,N_10729,N_10983);
and U17176 (N_17176,N_10985,N_12452);
or U17177 (N_17177,N_14811,N_10681);
nand U17178 (N_17178,N_14772,N_13217);
and U17179 (N_17179,N_12527,N_12807);
and U17180 (N_17180,N_13496,N_12217);
nand U17181 (N_17181,N_11004,N_13264);
nor U17182 (N_17182,N_14222,N_13736);
and U17183 (N_17183,N_12508,N_12596);
nand U17184 (N_17184,N_12921,N_12538);
nand U17185 (N_17185,N_12690,N_11383);
nand U17186 (N_17186,N_14111,N_12067);
nor U17187 (N_17187,N_11501,N_13571);
or U17188 (N_17188,N_13153,N_14052);
nor U17189 (N_17189,N_12412,N_11957);
or U17190 (N_17190,N_14670,N_13721);
and U17191 (N_17191,N_14101,N_14146);
nor U17192 (N_17192,N_11948,N_14374);
or U17193 (N_17193,N_12202,N_12964);
and U17194 (N_17194,N_10958,N_11003);
nand U17195 (N_17195,N_13260,N_14247);
and U17196 (N_17196,N_10030,N_10603);
or U17197 (N_17197,N_11623,N_14072);
or U17198 (N_17198,N_11812,N_11988);
nor U17199 (N_17199,N_14721,N_14963);
nand U17200 (N_17200,N_10559,N_14219);
or U17201 (N_17201,N_14299,N_14731);
or U17202 (N_17202,N_14840,N_10653);
xor U17203 (N_17203,N_13213,N_10939);
nand U17204 (N_17204,N_13547,N_10180);
and U17205 (N_17205,N_14197,N_10429);
and U17206 (N_17206,N_11687,N_11963);
nor U17207 (N_17207,N_11273,N_13211);
and U17208 (N_17208,N_10461,N_14373);
or U17209 (N_17209,N_13689,N_12679);
nor U17210 (N_17210,N_13877,N_13833);
xor U17211 (N_17211,N_13428,N_12104);
nor U17212 (N_17212,N_12951,N_11238);
nand U17213 (N_17213,N_10220,N_10284);
and U17214 (N_17214,N_12766,N_12565);
or U17215 (N_17215,N_14354,N_14616);
or U17216 (N_17216,N_13317,N_12352);
nand U17217 (N_17217,N_13081,N_11745);
nand U17218 (N_17218,N_12099,N_14803);
and U17219 (N_17219,N_11576,N_11221);
nand U17220 (N_17220,N_13015,N_12021);
and U17221 (N_17221,N_11267,N_14707);
nor U17222 (N_17222,N_10805,N_11662);
nand U17223 (N_17223,N_11523,N_11882);
or U17224 (N_17224,N_11897,N_14005);
and U17225 (N_17225,N_13868,N_13988);
nand U17226 (N_17226,N_12827,N_10242);
nor U17227 (N_17227,N_13126,N_14763);
nor U17228 (N_17228,N_10526,N_12614);
or U17229 (N_17229,N_10473,N_11555);
nor U17230 (N_17230,N_12206,N_10892);
and U17231 (N_17231,N_14534,N_13810);
nand U17232 (N_17232,N_11982,N_14273);
nand U17233 (N_17233,N_13715,N_10352);
nor U17234 (N_17234,N_10588,N_14419);
and U17235 (N_17235,N_14854,N_10277);
and U17236 (N_17236,N_12018,N_10073);
and U17237 (N_17237,N_11979,N_12993);
xor U17238 (N_17238,N_12787,N_10659);
nand U17239 (N_17239,N_12162,N_10245);
and U17240 (N_17240,N_11673,N_10044);
or U17241 (N_17241,N_10842,N_10718);
or U17242 (N_17242,N_13667,N_14034);
and U17243 (N_17243,N_12971,N_10164);
nor U17244 (N_17244,N_11867,N_13741);
xor U17245 (N_17245,N_12801,N_14057);
or U17246 (N_17246,N_14863,N_10781);
or U17247 (N_17247,N_12610,N_12621);
and U17248 (N_17248,N_14947,N_10095);
and U17249 (N_17249,N_11825,N_13325);
nor U17250 (N_17250,N_13597,N_14449);
and U17251 (N_17251,N_11884,N_10965);
or U17252 (N_17252,N_12636,N_14404);
and U17253 (N_17253,N_10128,N_10849);
nand U17254 (N_17254,N_10248,N_10015);
and U17255 (N_17255,N_14597,N_14871);
or U17256 (N_17256,N_12028,N_14384);
and U17257 (N_17257,N_12885,N_14786);
nand U17258 (N_17258,N_12907,N_12180);
and U17259 (N_17259,N_12567,N_12754);
and U17260 (N_17260,N_10497,N_12334);
xnor U17261 (N_17261,N_13053,N_14339);
nor U17262 (N_17262,N_10555,N_10358);
and U17263 (N_17263,N_14579,N_13974);
nor U17264 (N_17264,N_10934,N_13630);
and U17265 (N_17265,N_14953,N_12865);
and U17266 (N_17266,N_10862,N_12069);
nand U17267 (N_17267,N_11481,N_10562);
and U17268 (N_17268,N_10691,N_12168);
nor U17269 (N_17269,N_12260,N_14787);
or U17270 (N_17270,N_10919,N_14581);
and U17271 (N_17271,N_14575,N_11733);
nor U17272 (N_17272,N_14365,N_13021);
xnor U17273 (N_17273,N_12507,N_13272);
or U17274 (N_17274,N_13414,N_13418);
nor U17275 (N_17275,N_12604,N_10102);
nor U17276 (N_17276,N_13845,N_10210);
nand U17277 (N_17277,N_14120,N_14397);
and U17278 (N_17278,N_10391,N_10756);
and U17279 (N_17279,N_10209,N_11485);
or U17280 (N_17280,N_13058,N_14635);
nand U17281 (N_17281,N_13072,N_11365);
or U17282 (N_17282,N_10250,N_11476);
or U17283 (N_17283,N_12553,N_14998);
nor U17284 (N_17284,N_11769,N_12620);
or U17285 (N_17285,N_14056,N_13129);
nor U17286 (N_17286,N_10022,N_12424);
and U17287 (N_17287,N_13955,N_12017);
nor U17288 (N_17288,N_13172,N_10669);
or U17289 (N_17289,N_11418,N_10910);
or U17290 (N_17290,N_12528,N_14695);
and U17291 (N_17291,N_10921,N_14850);
and U17292 (N_17292,N_10415,N_12356);
or U17293 (N_17293,N_14601,N_10625);
nor U17294 (N_17294,N_11036,N_11816);
or U17295 (N_17295,N_14813,N_12769);
nor U17296 (N_17296,N_13941,N_11984);
or U17297 (N_17297,N_10825,N_14195);
or U17298 (N_17298,N_10496,N_13399);
nor U17299 (N_17299,N_11426,N_12239);
nand U17300 (N_17300,N_10698,N_14081);
nor U17301 (N_17301,N_10406,N_13340);
nor U17302 (N_17302,N_10647,N_13916);
or U17303 (N_17303,N_11612,N_12625);
or U17304 (N_17304,N_13943,N_11719);
or U17305 (N_17305,N_12835,N_10487);
or U17306 (N_17306,N_11527,N_10671);
and U17307 (N_17307,N_14319,N_12057);
or U17308 (N_17308,N_11966,N_11876);
or U17309 (N_17309,N_10812,N_14036);
nand U17310 (N_17310,N_11641,N_10023);
or U17311 (N_17311,N_14417,N_11734);
nand U17312 (N_17312,N_10822,N_14764);
and U17313 (N_17313,N_12544,N_14076);
xor U17314 (N_17314,N_12658,N_11711);
nand U17315 (N_17315,N_13527,N_14292);
nand U17316 (N_17316,N_10737,N_10004);
or U17317 (N_17317,N_11697,N_10032);
or U17318 (N_17318,N_10142,N_13760);
and U17319 (N_17319,N_14323,N_14066);
nor U17320 (N_17320,N_13512,N_10845);
nand U17321 (N_17321,N_10942,N_13266);
nand U17322 (N_17322,N_14479,N_12405);
and U17323 (N_17323,N_13289,N_13552);
or U17324 (N_17324,N_13529,N_12138);
nand U17325 (N_17325,N_12791,N_10744);
nor U17326 (N_17326,N_12978,N_10453);
nand U17327 (N_17327,N_11008,N_14269);
nand U17328 (N_17328,N_11441,N_11444);
and U17329 (N_17329,N_14143,N_12945);
or U17330 (N_17330,N_13777,N_11658);
nor U17331 (N_17331,N_10229,N_12918);
nand U17332 (N_17332,N_10399,N_10152);
and U17333 (N_17333,N_14096,N_14932);
and U17334 (N_17334,N_13551,N_14082);
nor U17335 (N_17335,N_14843,N_14016);
and U17336 (N_17336,N_10359,N_12468);
and U17337 (N_17337,N_13620,N_12254);
nor U17338 (N_17338,N_12533,N_14031);
nand U17339 (N_17339,N_14185,N_13825);
and U17340 (N_17340,N_14872,N_14887);
and U17341 (N_17341,N_14716,N_11239);
nor U17342 (N_17342,N_12664,N_11804);
xor U17343 (N_17343,N_13855,N_12158);
nand U17344 (N_17344,N_11191,N_13182);
and U17345 (N_17345,N_11193,N_11893);
and U17346 (N_17346,N_14715,N_12693);
nor U17347 (N_17347,N_10622,N_11431);
and U17348 (N_17348,N_13450,N_14608);
nand U17349 (N_17349,N_14127,N_10054);
and U17350 (N_17350,N_14288,N_11810);
nand U17351 (N_17351,N_14142,N_11336);
nand U17352 (N_17352,N_10760,N_13377);
nand U17353 (N_17353,N_13034,N_13706);
nor U17354 (N_17354,N_10536,N_12050);
nand U17355 (N_17355,N_13094,N_10620);
nand U17356 (N_17356,N_12629,N_12296);
or U17357 (N_17357,N_14276,N_10261);
nor U17358 (N_17358,N_11866,N_12848);
nand U17359 (N_17359,N_14131,N_12953);
nand U17360 (N_17360,N_12403,N_12670);
or U17361 (N_17361,N_12080,N_12802);
and U17362 (N_17362,N_13028,N_10212);
nor U17363 (N_17363,N_12572,N_10386);
nand U17364 (N_17364,N_10463,N_14006);
nor U17365 (N_17365,N_11344,N_13384);
nand U17366 (N_17366,N_10531,N_14425);
or U17367 (N_17367,N_13403,N_13936);
or U17368 (N_17368,N_10936,N_13485);
and U17369 (N_17369,N_14311,N_13624);
nand U17370 (N_17370,N_14303,N_12450);
or U17371 (N_17371,N_10769,N_11472);
nand U17372 (N_17372,N_11152,N_11285);
and U17373 (N_17373,N_14231,N_10541);
and U17374 (N_17374,N_11366,N_10899);
or U17375 (N_17375,N_13919,N_13098);
and U17376 (N_17376,N_14982,N_13174);
nand U17377 (N_17377,N_14007,N_13107);
or U17378 (N_17378,N_13383,N_10091);
nand U17379 (N_17379,N_11449,N_12120);
or U17380 (N_17380,N_12083,N_13456);
or U17381 (N_17381,N_10959,N_10813);
and U17382 (N_17382,N_14538,N_10482);
nor U17383 (N_17383,N_11962,N_13277);
and U17384 (N_17384,N_12874,N_14075);
nor U17385 (N_17385,N_14668,N_11709);
xnor U17386 (N_17386,N_10135,N_13586);
nand U17387 (N_17387,N_13253,N_13933);
nand U17388 (N_17388,N_10110,N_10097);
nor U17389 (N_17389,N_10507,N_12496);
or U17390 (N_17390,N_11268,N_13827);
nand U17391 (N_17391,N_14275,N_11560);
nor U17392 (N_17392,N_13326,N_13011);
nand U17393 (N_17393,N_13543,N_14302);
or U17394 (N_17394,N_10254,N_12838);
nor U17395 (N_17395,N_12241,N_14535);
nand U17396 (N_17396,N_11085,N_13117);
nor U17397 (N_17397,N_10201,N_10071);
or U17398 (N_17398,N_11704,N_13088);
or U17399 (N_17399,N_11774,N_13467);
or U17400 (N_17400,N_11342,N_14519);
or U17401 (N_17401,N_14655,N_12702);
or U17402 (N_17402,N_12550,N_12877);
nand U17403 (N_17403,N_11869,N_11909);
or U17404 (N_17404,N_12510,N_13079);
nand U17405 (N_17405,N_14596,N_10270);
nor U17406 (N_17406,N_14285,N_10370);
and U17407 (N_17407,N_10448,N_10118);
nor U17408 (N_17408,N_11374,N_12500);
nand U17409 (N_17409,N_12000,N_10165);
nor U17410 (N_17410,N_13368,N_13144);
xnor U17411 (N_17411,N_11467,N_13321);
nand U17412 (N_17412,N_10762,N_10817);
or U17413 (N_17413,N_11095,N_12343);
nand U17414 (N_17414,N_11668,N_11533);
nor U17415 (N_17415,N_14001,N_13785);
nor U17416 (N_17416,N_12534,N_13396);
or U17417 (N_17417,N_13663,N_14615);
xor U17418 (N_17418,N_13487,N_11473);
nand U17419 (N_17419,N_11156,N_10158);
and U17420 (N_17420,N_13489,N_10367);
or U17421 (N_17421,N_13030,N_11970);
nand U17422 (N_17422,N_11241,N_11470);
and U17423 (N_17423,N_14961,N_13027);
nor U17424 (N_17424,N_12694,N_13329);
nor U17425 (N_17425,N_10411,N_13638);
xor U17426 (N_17426,N_12812,N_11585);
and U17427 (N_17427,N_10827,N_13370);
nand U17428 (N_17428,N_11389,N_12897);
and U17429 (N_17429,N_13656,N_11770);
nand U17430 (N_17430,N_12130,N_12519);
nand U17431 (N_17431,N_11210,N_10040);
and U17432 (N_17432,N_13170,N_12431);
and U17433 (N_17433,N_13279,N_11718);
nand U17434 (N_17434,N_14984,N_14439);
and U17435 (N_17435,N_11785,N_14784);
nor U17436 (N_17436,N_12458,N_13400);
nand U17437 (N_17437,N_14182,N_12347);
nor U17438 (N_17438,N_12705,N_10060);
xor U17439 (N_17439,N_10452,N_10925);
and U17440 (N_17440,N_14350,N_11177);
nor U17441 (N_17441,N_13379,N_13406);
nor U17442 (N_17442,N_11543,N_14965);
nand U17443 (N_17443,N_11211,N_12196);
nor U17444 (N_17444,N_12248,N_13708);
nand U17445 (N_17445,N_13832,N_13615);
or U17446 (N_17446,N_12962,N_12903);
nand U17447 (N_17447,N_10794,N_12094);
or U17448 (N_17448,N_11667,N_14043);
and U17449 (N_17449,N_13357,N_13835);
nand U17450 (N_17450,N_11892,N_10592);
nand U17451 (N_17451,N_13344,N_10550);
or U17452 (N_17452,N_11265,N_11489);
or U17453 (N_17453,N_14975,N_13381);
and U17454 (N_17454,N_12994,N_11223);
or U17455 (N_17455,N_13274,N_14038);
nor U17456 (N_17456,N_12091,N_11648);
or U17457 (N_17457,N_10747,N_14186);
or U17458 (N_17458,N_13755,N_13494);
nand U17459 (N_17459,N_10572,N_12209);
or U17460 (N_17460,N_11315,N_11041);
nor U17461 (N_17461,N_13482,N_10483);
nor U17462 (N_17462,N_12786,N_11846);
and U17463 (N_17463,N_12375,N_10331);
xor U17464 (N_17464,N_12293,N_12268);
nand U17465 (N_17465,N_14164,N_14458);
nor U17466 (N_17466,N_14246,N_14722);
and U17467 (N_17467,N_14059,N_14890);
xor U17468 (N_17468,N_14010,N_13229);
nor U17469 (N_17469,N_11289,N_11200);
xnor U17470 (N_17470,N_11479,N_10940);
or U17471 (N_17471,N_11545,N_12909);
and U17472 (N_17472,N_10612,N_13054);
xor U17473 (N_17473,N_13582,N_12417);
and U17474 (N_17474,N_10623,N_14361);
and U17475 (N_17475,N_12329,N_10981);
nor U17476 (N_17476,N_10309,N_13535);
and U17477 (N_17477,N_14117,N_13185);
or U17478 (N_17478,N_10267,N_11670);
nand U17479 (N_17479,N_13435,N_12364);
and U17480 (N_17480,N_10602,N_11143);
and U17481 (N_17481,N_11781,N_11834);
or U17482 (N_17482,N_13781,N_14353);
nor U17483 (N_17483,N_10742,N_12805);
nor U17484 (N_17484,N_12515,N_12653);
or U17485 (N_17485,N_12277,N_10798);
nor U17486 (N_17486,N_11139,N_14515);
xor U17487 (N_17487,N_11000,N_12932);
and U17488 (N_17488,N_14011,N_14268);
or U17489 (N_17489,N_13937,N_11319);
nand U17490 (N_17490,N_14403,N_10847);
nor U17491 (N_17491,N_13412,N_13770);
and U17492 (N_17492,N_11831,N_14123);
and U17493 (N_17493,N_14387,N_14826);
xnor U17494 (N_17494,N_14939,N_14442);
nor U17495 (N_17495,N_13691,N_13056);
nand U17496 (N_17496,N_11508,N_11168);
and U17497 (N_17497,N_14343,N_12800);
and U17498 (N_17498,N_12462,N_11678);
and U17499 (N_17499,N_13197,N_14376);
nand U17500 (N_17500,N_10893,N_14447);
nand U17501 (N_17501,N_11332,N_10058);
or U17502 (N_17502,N_12405,N_14656);
and U17503 (N_17503,N_11948,N_11836);
and U17504 (N_17504,N_13635,N_10341);
nand U17505 (N_17505,N_11409,N_11939);
xnor U17506 (N_17506,N_13224,N_10405);
or U17507 (N_17507,N_14228,N_11230);
or U17508 (N_17508,N_12155,N_10733);
or U17509 (N_17509,N_13991,N_12729);
or U17510 (N_17510,N_14358,N_10160);
and U17511 (N_17511,N_10312,N_10949);
and U17512 (N_17512,N_12435,N_14881);
or U17513 (N_17513,N_14311,N_10915);
nand U17514 (N_17514,N_10482,N_13194);
and U17515 (N_17515,N_11356,N_14322);
nor U17516 (N_17516,N_11459,N_11894);
and U17517 (N_17517,N_12385,N_11304);
and U17518 (N_17518,N_11007,N_12074);
and U17519 (N_17519,N_13835,N_12078);
or U17520 (N_17520,N_11079,N_12010);
nand U17521 (N_17521,N_14779,N_12334);
nor U17522 (N_17522,N_14893,N_14415);
nor U17523 (N_17523,N_13422,N_10040);
nand U17524 (N_17524,N_14360,N_10153);
and U17525 (N_17525,N_11061,N_10621);
or U17526 (N_17526,N_13693,N_10615);
or U17527 (N_17527,N_14320,N_12753);
and U17528 (N_17528,N_14676,N_11062);
and U17529 (N_17529,N_11157,N_12658);
nand U17530 (N_17530,N_13809,N_10860);
nand U17531 (N_17531,N_11358,N_12184);
nor U17532 (N_17532,N_12402,N_11153);
or U17533 (N_17533,N_10141,N_13182);
nand U17534 (N_17534,N_13165,N_12315);
or U17535 (N_17535,N_11491,N_11587);
nand U17536 (N_17536,N_13411,N_10560);
or U17537 (N_17537,N_14353,N_13292);
nor U17538 (N_17538,N_13399,N_14421);
nor U17539 (N_17539,N_13427,N_11248);
nor U17540 (N_17540,N_11515,N_10366);
and U17541 (N_17541,N_10904,N_14648);
or U17542 (N_17542,N_13546,N_13130);
nor U17543 (N_17543,N_11725,N_12165);
nand U17544 (N_17544,N_12208,N_14721);
nand U17545 (N_17545,N_10087,N_11312);
nor U17546 (N_17546,N_11006,N_14699);
nand U17547 (N_17547,N_13754,N_12739);
or U17548 (N_17548,N_12714,N_13986);
nand U17549 (N_17549,N_14359,N_12697);
nor U17550 (N_17550,N_11693,N_14641);
nand U17551 (N_17551,N_14302,N_11839);
and U17552 (N_17552,N_10302,N_12388);
nand U17553 (N_17553,N_14154,N_12444);
nor U17554 (N_17554,N_11477,N_13829);
nand U17555 (N_17555,N_12864,N_10041);
or U17556 (N_17556,N_13873,N_11113);
nor U17557 (N_17557,N_13511,N_11164);
or U17558 (N_17558,N_11347,N_12197);
nand U17559 (N_17559,N_12775,N_10892);
nand U17560 (N_17560,N_14177,N_11969);
nor U17561 (N_17561,N_11938,N_11515);
xnor U17562 (N_17562,N_14303,N_13541);
nor U17563 (N_17563,N_11418,N_14456);
or U17564 (N_17564,N_10916,N_13320);
nor U17565 (N_17565,N_13218,N_14923);
and U17566 (N_17566,N_14157,N_14365);
or U17567 (N_17567,N_10438,N_12468);
and U17568 (N_17568,N_11540,N_10984);
nand U17569 (N_17569,N_14399,N_12589);
or U17570 (N_17570,N_10119,N_14475);
nor U17571 (N_17571,N_12216,N_10883);
nor U17572 (N_17572,N_13047,N_11030);
and U17573 (N_17573,N_13137,N_11450);
and U17574 (N_17574,N_12793,N_14650);
xor U17575 (N_17575,N_14142,N_14161);
nor U17576 (N_17576,N_11129,N_14959);
and U17577 (N_17577,N_10628,N_12844);
or U17578 (N_17578,N_12086,N_11060);
or U17579 (N_17579,N_13410,N_14647);
and U17580 (N_17580,N_10729,N_14741);
nor U17581 (N_17581,N_12710,N_10707);
nand U17582 (N_17582,N_10439,N_12089);
nand U17583 (N_17583,N_14910,N_12226);
or U17584 (N_17584,N_14111,N_10472);
and U17585 (N_17585,N_14673,N_12740);
and U17586 (N_17586,N_10997,N_11233);
nor U17587 (N_17587,N_11906,N_14865);
or U17588 (N_17588,N_13869,N_13859);
nand U17589 (N_17589,N_13886,N_12820);
nand U17590 (N_17590,N_14199,N_10439);
or U17591 (N_17591,N_14343,N_12343);
and U17592 (N_17592,N_10851,N_11196);
and U17593 (N_17593,N_11181,N_13426);
or U17594 (N_17594,N_14339,N_14587);
or U17595 (N_17595,N_12899,N_13697);
nand U17596 (N_17596,N_10482,N_13538);
nand U17597 (N_17597,N_12891,N_14228);
xnor U17598 (N_17598,N_14055,N_11282);
or U17599 (N_17599,N_11989,N_10001);
and U17600 (N_17600,N_13301,N_10422);
and U17601 (N_17601,N_13382,N_14248);
nor U17602 (N_17602,N_11797,N_12626);
or U17603 (N_17603,N_10128,N_14640);
or U17604 (N_17604,N_14657,N_10619);
nor U17605 (N_17605,N_14982,N_10195);
and U17606 (N_17606,N_11651,N_12434);
or U17607 (N_17607,N_11915,N_13970);
and U17608 (N_17608,N_10797,N_11045);
and U17609 (N_17609,N_10693,N_12581);
or U17610 (N_17610,N_10177,N_14900);
or U17611 (N_17611,N_14550,N_13707);
or U17612 (N_17612,N_14637,N_12555);
and U17613 (N_17613,N_10387,N_11744);
nor U17614 (N_17614,N_10642,N_10294);
or U17615 (N_17615,N_12963,N_11405);
xor U17616 (N_17616,N_12546,N_10152);
and U17617 (N_17617,N_14635,N_12196);
and U17618 (N_17618,N_11942,N_11192);
and U17619 (N_17619,N_10661,N_11504);
or U17620 (N_17620,N_13858,N_12689);
or U17621 (N_17621,N_14118,N_10959);
or U17622 (N_17622,N_13182,N_13819);
nand U17623 (N_17623,N_13174,N_12123);
or U17624 (N_17624,N_12418,N_13651);
nand U17625 (N_17625,N_11942,N_12211);
and U17626 (N_17626,N_12200,N_12720);
nand U17627 (N_17627,N_13621,N_11296);
and U17628 (N_17628,N_13135,N_13694);
and U17629 (N_17629,N_11493,N_14353);
nor U17630 (N_17630,N_11835,N_11993);
or U17631 (N_17631,N_10023,N_12798);
xnor U17632 (N_17632,N_12827,N_13704);
or U17633 (N_17633,N_10412,N_13007);
or U17634 (N_17634,N_13470,N_11342);
nor U17635 (N_17635,N_14903,N_11167);
nand U17636 (N_17636,N_14748,N_10724);
or U17637 (N_17637,N_13008,N_11630);
xor U17638 (N_17638,N_13385,N_11736);
nor U17639 (N_17639,N_10032,N_13992);
nand U17640 (N_17640,N_11517,N_13742);
nor U17641 (N_17641,N_14065,N_13905);
nor U17642 (N_17642,N_10264,N_11093);
nor U17643 (N_17643,N_14692,N_12229);
or U17644 (N_17644,N_14091,N_12491);
nand U17645 (N_17645,N_14357,N_13836);
and U17646 (N_17646,N_13841,N_12735);
xor U17647 (N_17647,N_10749,N_10447);
and U17648 (N_17648,N_10118,N_11347);
or U17649 (N_17649,N_14900,N_11274);
and U17650 (N_17650,N_12734,N_13852);
or U17651 (N_17651,N_11228,N_10326);
nor U17652 (N_17652,N_12274,N_10404);
or U17653 (N_17653,N_12929,N_13987);
nor U17654 (N_17654,N_13143,N_12424);
nor U17655 (N_17655,N_11494,N_14934);
nor U17656 (N_17656,N_10410,N_10223);
and U17657 (N_17657,N_12418,N_13312);
and U17658 (N_17658,N_12646,N_10149);
or U17659 (N_17659,N_14688,N_11549);
nor U17660 (N_17660,N_12965,N_14299);
nand U17661 (N_17661,N_13373,N_10967);
xnor U17662 (N_17662,N_12599,N_12000);
nor U17663 (N_17663,N_13740,N_13996);
or U17664 (N_17664,N_11743,N_11280);
or U17665 (N_17665,N_10710,N_14962);
nor U17666 (N_17666,N_10818,N_13635);
or U17667 (N_17667,N_12999,N_10040);
nand U17668 (N_17668,N_10713,N_11766);
nand U17669 (N_17669,N_11418,N_14699);
nand U17670 (N_17670,N_14956,N_11193);
and U17671 (N_17671,N_12757,N_13024);
or U17672 (N_17672,N_10332,N_13325);
nor U17673 (N_17673,N_10846,N_13052);
and U17674 (N_17674,N_12916,N_10346);
or U17675 (N_17675,N_10232,N_11750);
or U17676 (N_17676,N_10964,N_14989);
nand U17677 (N_17677,N_14865,N_14256);
and U17678 (N_17678,N_12574,N_13601);
nand U17679 (N_17679,N_10184,N_10295);
nor U17680 (N_17680,N_12325,N_14355);
nand U17681 (N_17681,N_11158,N_13411);
nor U17682 (N_17682,N_11529,N_12755);
nand U17683 (N_17683,N_12761,N_14982);
nor U17684 (N_17684,N_14735,N_14243);
and U17685 (N_17685,N_12861,N_11516);
or U17686 (N_17686,N_11916,N_14951);
nand U17687 (N_17687,N_11763,N_13374);
nand U17688 (N_17688,N_11858,N_14405);
nor U17689 (N_17689,N_12535,N_11042);
nand U17690 (N_17690,N_11173,N_12481);
or U17691 (N_17691,N_13212,N_14558);
and U17692 (N_17692,N_13310,N_13071);
nor U17693 (N_17693,N_12611,N_11487);
nand U17694 (N_17694,N_10015,N_10461);
nand U17695 (N_17695,N_13937,N_10298);
and U17696 (N_17696,N_13317,N_13254);
nand U17697 (N_17697,N_12150,N_11365);
nor U17698 (N_17698,N_10883,N_10717);
nand U17699 (N_17699,N_13355,N_14557);
or U17700 (N_17700,N_12881,N_12182);
nor U17701 (N_17701,N_11421,N_10886);
nor U17702 (N_17702,N_14315,N_10436);
nand U17703 (N_17703,N_14141,N_13569);
and U17704 (N_17704,N_14864,N_13365);
or U17705 (N_17705,N_13059,N_13930);
nand U17706 (N_17706,N_10931,N_10964);
nor U17707 (N_17707,N_14552,N_12158);
or U17708 (N_17708,N_12791,N_11817);
nand U17709 (N_17709,N_12468,N_10973);
nor U17710 (N_17710,N_12802,N_12308);
nand U17711 (N_17711,N_14839,N_12547);
or U17712 (N_17712,N_11270,N_11515);
and U17713 (N_17713,N_10283,N_12187);
or U17714 (N_17714,N_13422,N_10517);
nand U17715 (N_17715,N_11209,N_13434);
and U17716 (N_17716,N_10156,N_10894);
or U17717 (N_17717,N_13713,N_13912);
nand U17718 (N_17718,N_12575,N_13859);
nand U17719 (N_17719,N_10702,N_11859);
nand U17720 (N_17720,N_11891,N_11769);
nand U17721 (N_17721,N_13609,N_13838);
nand U17722 (N_17722,N_12119,N_11565);
nand U17723 (N_17723,N_14810,N_11243);
xor U17724 (N_17724,N_13868,N_13216);
and U17725 (N_17725,N_13697,N_12943);
nand U17726 (N_17726,N_11556,N_10642);
nand U17727 (N_17727,N_10628,N_11236);
or U17728 (N_17728,N_11324,N_13230);
and U17729 (N_17729,N_12880,N_10538);
or U17730 (N_17730,N_13528,N_14172);
xnor U17731 (N_17731,N_13472,N_14858);
nor U17732 (N_17732,N_12314,N_12165);
nor U17733 (N_17733,N_12384,N_10251);
and U17734 (N_17734,N_14549,N_14972);
and U17735 (N_17735,N_14113,N_10451);
nor U17736 (N_17736,N_11514,N_13827);
nor U17737 (N_17737,N_11149,N_14286);
nand U17738 (N_17738,N_13294,N_13183);
and U17739 (N_17739,N_12789,N_14579);
nand U17740 (N_17740,N_14833,N_10954);
or U17741 (N_17741,N_10809,N_13092);
or U17742 (N_17742,N_12747,N_14294);
and U17743 (N_17743,N_14081,N_13926);
nor U17744 (N_17744,N_13089,N_12958);
nor U17745 (N_17745,N_12086,N_13897);
nand U17746 (N_17746,N_12429,N_14948);
nand U17747 (N_17747,N_13141,N_10675);
nor U17748 (N_17748,N_13380,N_10428);
and U17749 (N_17749,N_14984,N_13016);
nor U17750 (N_17750,N_14248,N_11278);
and U17751 (N_17751,N_12508,N_13165);
and U17752 (N_17752,N_12410,N_10556);
and U17753 (N_17753,N_13516,N_11383);
nor U17754 (N_17754,N_11335,N_13755);
nand U17755 (N_17755,N_12006,N_14849);
or U17756 (N_17756,N_13087,N_12571);
nand U17757 (N_17757,N_12319,N_12681);
and U17758 (N_17758,N_14906,N_10560);
nor U17759 (N_17759,N_13337,N_10016);
nand U17760 (N_17760,N_14782,N_10513);
nand U17761 (N_17761,N_11070,N_10752);
nor U17762 (N_17762,N_10687,N_11648);
or U17763 (N_17763,N_13993,N_11883);
nand U17764 (N_17764,N_11865,N_10937);
and U17765 (N_17765,N_12819,N_10457);
nor U17766 (N_17766,N_13654,N_11100);
or U17767 (N_17767,N_10092,N_11086);
and U17768 (N_17768,N_12916,N_11597);
nand U17769 (N_17769,N_10291,N_10279);
nand U17770 (N_17770,N_10741,N_10328);
and U17771 (N_17771,N_14167,N_14317);
and U17772 (N_17772,N_12539,N_14863);
nand U17773 (N_17773,N_13920,N_13449);
nand U17774 (N_17774,N_11018,N_14326);
and U17775 (N_17775,N_11600,N_12877);
nand U17776 (N_17776,N_12100,N_11974);
nor U17777 (N_17777,N_10978,N_12308);
or U17778 (N_17778,N_14720,N_13100);
or U17779 (N_17779,N_13903,N_10844);
or U17780 (N_17780,N_12352,N_11635);
and U17781 (N_17781,N_13569,N_13625);
nor U17782 (N_17782,N_11237,N_10337);
nand U17783 (N_17783,N_12183,N_13206);
nand U17784 (N_17784,N_11324,N_12956);
or U17785 (N_17785,N_13684,N_12024);
nor U17786 (N_17786,N_11322,N_14995);
nand U17787 (N_17787,N_13304,N_13018);
nor U17788 (N_17788,N_13420,N_13002);
and U17789 (N_17789,N_13690,N_13508);
and U17790 (N_17790,N_10748,N_11967);
nor U17791 (N_17791,N_14857,N_14519);
or U17792 (N_17792,N_12733,N_10379);
nand U17793 (N_17793,N_10519,N_12492);
nand U17794 (N_17794,N_12273,N_10604);
nand U17795 (N_17795,N_13597,N_10028);
and U17796 (N_17796,N_12961,N_10967);
nor U17797 (N_17797,N_10671,N_14348);
and U17798 (N_17798,N_14210,N_12070);
or U17799 (N_17799,N_13605,N_11968);
nor U17800 (N_17800,N_12197,N_12760);
and U17801 (N_17801,N_13071,N_11031);
or U17802 (N_17802,N_10172,N_12752);
nand U17803 (N_17803,N_14403,N_12092);
and U17804 (N_17804,N_14823,N_13000);
nand U17805 (N_17805,N_13689,N_11670);
or U17806 (N_17806,N_12022,N_14020);
xor U17807 (N_17807,N_12238,N_10439);
xnor U17808 (N_17808,N_13016,N_13858);
nand U17809 (N_17809,N_11519,N_14823);
nand U17810 (N_17810,N_10973,N_11613);
nor U17811 (N_17811,N_10109,N_10099);
nor U17812 (N_17812,N_10270,N_10870);
and U17813 (N_17813,N_13184,N_14735);
and U17814 (N_17814,N_10318,N_11345);
nor U17815 (N_17815,N_10263,N_13256);
nand U17816 (N_17816,N_13316,N_13555);
or U17817 (N_17817,N_13114,N_11621);
nand U17818 (N_17818,N_10262,N_10326);
and U17819 (N_17819,N_11273,N_14175);
nor U17820 (N_17820,N_11328,N_11559);
nand U17821 (N_17821,N_10478,N_10474);
nor U17822 (N_17822,N_11175,N_11362);
nand U17823 (N_17823,N_11317,N_13943);
nor U17824 (N_17824,N_11544,N_10025);
nor U17825 (N_17825,N_14735,N_13177);
nand U17826 (N_17826,N_10322,N_12451);
xnor U17827 (N_17827,N_13325,N_13124);
or U17828 (N_17828,N_11007,N_14476);
nor U17829 (N_17829,N_12184,N_13135);
or U17830 (N_17830,N_12240,N_10744);
nor U17831 (N_17831,N_11390,N_10415);
nand U17832 (N_17832,N_12779,N_11902);
nand U17833 (N_17833,N_13370,N_10964);
nor U17834 (N_17834,N_11625,N_11734);
nor U17835 (N_17835,N_11590,N_13778);
nand U17836 (N_17836,N_13674,N_11996);
or U17837 (N_17837,N_11957,N_14775);
or U17838 (N_17838,N_13586,N_12240);
nor U17839 (N_17839,N_10447,N_11031);
or U17840 (N_17840,N_13953,N_11718);
nor U17841 (N_17841,N_10107,N_10844);
nand U17842 (N_17842,N_14368,N_13061);
and U17843 (N_17843,N_12898,N_11303);
and U17844 (N_17844,N_13146,N_13802);
and U17845 (N_17845,N_14110,N_14804);
and U17846 (N_17846,N_10429,N_13557);
nand U17847 (N_17847,N_13682,N_13446);
and U17848 (N_17848,N_12150,N_12847);
or U17849 (N_17849,N_13382,N_11725);
nor U17850 (N_17850,N_11606,N_12449);
or U17851 (N_17851,N_11778,N_10380);
nor U17852 (N_17852,N_13771,N_13368);
and U17853 (N_17853,N_11979,N_10415);
nor U17854 (N_17854,N_11479,N_14427);
nor U17855 (N_17855,N_13144,N_13370);
or U17856 (N_17856,N_14543,N_10636);
nand U17857 (N_17857,N_13648,N_10885);
and U17858 (N_17858,N_13372,N_12015);
and U17859 (N_17859,N_11836,N_10146);
or U17860 (N_17860,N_11722,N_14389);
and U17861 (N_17861,N_12628,N_13804);
or U17862 (N_17862,N_11960,N_14276);
or U17863 (N_17863,N_12029,N_10864);
and U17864 (N_17864,N_10833,N_10533);
and U17865 (N_17865,N_14020,N_12208);
nor U17866 (N_17866,N_14375,N_11775);
or U17867 (N_17867,N_13215,N_12857);
or U17868 (N_17868,N_14234,N_14349);
nor U17869 (N_17869,N_14126,N_10175);
or U17870 (N_17870,N_10028,N_10280);
xnor U17871 (N_17871,N_12978,N_12818);
and U17872 (N_17872,N_10440,N_11469);
nor U17873 (N_17873,N_11979,N_12966);
nor U17874 (N_17874,N_11532,N_10353);
and U17875 (N_17875,N_13946,N_14891);
or U17876 (N_17876,N_14001,N_14231);
and U17877 (N_17877,N_10371,N_13928);
nor U17878 (N_17878,N_11944,N_12774);
and U17879 (N_17879,N_13370,N_11720);
nand U17880 (N_17880,N_10963,N_11818);
nor U17881 (N_17881,N_10537,N_11390);
nor U17882 (N_17882,N_10109,N_11105);
nand U17883 (N_17883,N_14949,N_12523);
nor U17884 (N_17884,N_12841,N_10093);
nor U17885 (N_17885,N_11379,N_14259);
nor U17886 (N_17886,N_10662,N_13245);
or U17887 (N_17887,N_13595,N_12805);
xnor U17888 (N_17888,N_11110,N_14792);
or U17889 (N_17889,N_11278,N_10967);
or U17890 (N_17890,N_14660,N_14623);
and U17891 (N_17891,N_13885,N_11704);
nand U17892 (N_17892,N_14251,N_14073);
or U17893 (N_17893,N_11531,N_12069);
nand U17894 (N_17894,N_10993,N_11458);
and U17895 (N_17895,N_13969,N_12866);
nand U17896 (N_17896,N_10812,N_12900);
nand U17897 (N_17897,N_13345,N_12474);
and U17898 (N_17898,N_12543,N_14262);
nor U17899 (N_17899,N_11998,N_13111);
and U17900 (N_17900,N_13783,N_10715);
or U17901 (N_17901,N_11962,N_11931);
or U17902 (N_17902,N_10514,N_11605);
nand U17903 (N_17903,N_13047,N_14121);
or U17904 (N_17904,N_14206,N_10638);
nand U17905 (N_17905,N_13077,N_13353);
nand U17906 (N_17906,N_10247,N_12854);
nor U17907 (N_17907,N_12523,N_13378);
nor U17908 (N_17908,N_10581,N_11372);
or U17909 (N_17909,N_10383,N_11105);
and U17910 (N_17910,N_13520,N_14715);
or U17911 (N_17911,N_14442,N_14834);
nor U17912 (N_17912,N_12645,N_13653);
or U17913 (N_17913,N_11400,N_10946);
nor U17914 (N_17914,N_13899,N_11886);
or U17915 (N_17915,N_13101,N_10264);
nor U17916 (N_17916,N_14624,N_14871);
and U17917 (N_17917,N_13369,N_13146);
and U17918 (N_17918,N_11358,N_10035);
nand U17919 (N_17919,N_12067,N_10542);
or U17920 (N_17920,N_14622,N_12332);
nand U17921 (N_17921,N_11420,N_10240);
nor U17922 (N_17922,N_10088,N_10789);
or U17923 (N_17923,N_12551,N_13744);
nand U17924 (N_17924,N_13662,N_14469);
nand U17925 (N_17925,N_14159,N_10918);
and U17926 (N_17926,N_10532,N_10132);
nor U17927 (N_17927,N_13387,N_13367);
and U17928 (N_17928,N_13907,N_13411);
xor U17929 (N_17929,N_12866,N_10931);
and U17930 (N_17930,N_10746,N_12943);
and U17931 (N_17931,N_10052,N_14794);
nor U17932 (N_17932,N_10278,N_10544);
nor U17933 (N_17933,N_14331,N_11819);
nor U17934 (N_17934,N_11871,N_14506);
nor U17935 (N_17935,N_10369,N_10156);
nand U17936 (N_17936,N_12634,N_10367);
nand U17937 (N_17937,N_10509,N_10531);
and U17938 (N_17938,N_11845,N_12115);
nor U17939 (N_17939,N_14935,N_13266);
nor U17940 (N_17940,N_12303,N_10546);
nand U17941 (N_17941,N_12026,N_11547);
nor U17942 (N_17942,N_10513,N_13896);
nand U17943 (N_17943,N_14943,N_14612);
nand U17944 (N_17944,N_12872,N_12398);
and U17945 (N_17945,N_13899,N_13631);
nor U17946 (N_17946,N_10412,N_14466);
nor U17947 (N_17947,N_12221,N_14753);
xnor U17948 (N_17948,N_13605,N_10042);
and U17949 (N_17949,N_12349,N_10816);
or U17950 (N_17950,N_11740,N_10045);
or U17951 (N_17951,N_10565,N_14172);
or U17952 (N_17952,N_12357,N_12336);
nand U17953 (N_17953,N_10546,N_11817);
or U17954 (N_17954,N_13591,N_11336);
nand U17955 (N_17955,N_13085,N_10067);
and U17956 (N_17956,N_13312,N_10040);
or U17957 (N_17957,N_10462,N_11025);
or U17958 (N_17958,N_10900,N_10072);
nand U17959 (N_17959,N_10209,N_14137);
or U17960 (N_17960,N_10723,N_14476);
nand U17961 (N_17961,N_10805,N_13238);
and U17962 (N_17962,N_14656,N_12758);
or U17963 (N_17963,N_12847,N_13854);
nand U17964 (N_17964,N_13483,N_10980);
nand U17965 (N_17965,N_10988,N_14809);
nand U17966 (N_17966,N_14594,N_11889);
nand U17967 (N_17967,N_11233,N_11940);
nor U17968 (N_17968,N_10823,N_11658);
nor U17969 (N_17969,N_13197,N_10958);
and U17970 (N_17970,N_12427,N_12794);
nor U17971 (N_17971,N_13107,N_14230);
nand U17972 (N_17972,N_11594,N_13054);
nand U17973 (N_17973,N_14962,N_14882);
xor U17974 (N_17974,N_12905,N_12027);
nand U17975 (N_17975,N_14902,N_14322);
nor U17976 (N_17976,N_13865,N_11989);
nand U17977 (N_17977,N_11301,N_12962);
or U17978 (N_17978,N_12581,N_14308);
or U17979 (N_17979,N_11551,N_14730);
and U17980 (N_17980,N_11531,N_13563);
and U17981 (N_17981,N_10585,N_11436);
nor U17982 (N_17982,N_14483,N_11929);
or U17983 (N_17983,N_11220,N_14368);
nor U17984 (N_17984,N_14745,N_14597);
or U17985 (N_17985,N_11473,N_13246);
or U17986 (N_17986,N_13589,N_12973);
nor U17987 (N_17987,N_12078,N_12199);
or U17988 (N_17988,N_14165,N_12959);
xor U17989 (N_17989,N_11754,N_13905);
nand U17990 (N_17990,N_10265,N_14670);
and U17991 (N_17991,N_12168,N_11768);
nand U17992 (N_17992,N_11966,N_10264);
and U17993 (N_17993,N_11320,N_13603);
and U17994 (N_17994,N_11325,N_14088);
xor U17995 (N_17995,N_12450,N_14911);
and U17996 (N_17996,N_12590,N_12156);
or U17997 (N_17997,N_14007,N_13440);
or U17998 (N_17998,N_13425,N_14538);
or U17999 (N_17999,N_11702,N_10655);
and U18000 (N_18000,N_13793,N_11653);
nor U18001 (N_18001,N_10678,N_13522);
and U18002 (N_18002,N_11424,N_10325);
nand U18003 (N_18003,N_10997,N_11671);
nor U18004 (N_18004,N_11209,N_10747);
or U18005 (N_18005,N_14448,N_12045);
and U18006 (N_18006,N_14125,N_13776);
or U18007 (N_18007,N_14158,N_14974);
or U18008 (N_18008,N_10507,N_14402);
nor U18009 (N_18009,N_12423,N_13701);
nand U18010 (N_18010,N_13590,N_13764);
nand U18011 (N_18011,N_13369,N_12092);
and U18012 (N_18012,N_11974,N_14538);
nand U18013 (N_18013,N_14980,N_11017);
or U18014 (N_18014,N_14438,N_14543);
or U18015 (N_18015,N_14169,N_11022);
or U18016 (N_18016,N_12716,N_12725);
xnor U18017 (N_18017,N_11180,N_12964);
or U18018 (N_18018,N_10757,N_14008);
nand U18019 (N_18019,N_11656,N_12328);
or U18020 (N_18020,N_11542,N_14274);
or U18021 (N_18021,N_14435,N_10421);
nor U18022 (N_18022,N_13613,N_12086);
or U18023 (N_18023,N_11725,N_12520);
and U18024 (N_18024,N_10448,N_13015);
nor U18025 (N_18025,N_11509,N_14533);
nor U18026 (N_18026,N_11347,N_12030);
nor U18027 (N_18027,N_12169,N_13288);
and U18028 (N_18028,N_13775,N_12079);
nand U18029 (N_18029,N_12380,N_10148);
nand U18030 (N_18030,N_10369,N_10571);
or U18031 (N_18031,N_12282,N_10452);
nor U18032 (N_18032,N_11367,N_11642);
nand U18033 (N_18033,N_12076,N_12939);
nor U18034 (N_18034,N_10154,N_12656);
nor U18035 (N_18035,N_11145,N_10499);
nor U18036 (N_18036,N_14542,N_14430);
nand U18037 (N_18037,N_12179,N_11092);
or U18038 (N_18038,N_13894,N_13494);
nand U18039 (N_18039,N_14788,N_11017);
nand U18040 (N_18040,N_10763,N_11085);
nand U18041 (N_18041,N_14944,N_12857);
or U18042 (N_18042,N_14601,N_14489);
nor U18043 (N_18043,N_11696,N_13295);
or U18044 (N_18044,N_11045,N_14685);
nand U18045 (N_18045,N_14946,N_12901);
and U18046 (N_18046,N_13673,N_14833);
and U18047 (N_18047,N_12995,N_12571);
and U18048 (N_18048,N_11462,N_12540);
or U18049 (N_18049,N_12953,N_10555);
and U18050 (N_18050,N_14537,N_10356);
or U18051 (N_18051,N_11751,N_10770);
nor U18052 (N_18052,N_14541,N_14882);
or U18053 (N_18053,N_11394,N_11174);
nor U18054 (N_18054,N_13447,N_14982);
or U18055 (N_18055,N_10961,N_10618);
nor U18056 (N_18056,N_14916,N_14181);
nor U18057 (N_18057,N_10307,N_12803);
and U18058 (N_18058,N_12684,N_13311);
or U18059 (N_18059,N_13116,N_11792);
and U18060 (N_18060,N_13211,N_10078);
or U18061 (N_18061,N_13607,N_10733);
and U18062 (N_18062,N_14063,N_12491);
nand U18063 (N_18063,N_12527,N_14933);
nor U18064 (N_18064,N_12491,N_14427);
nand U18065 (N_18065,N_11494,N_13125);
nand U18066 (N_18066,N_11552,N_14464);
nor U18067 (N_18067,N_10877,N_10650);
nand U18068 (N_18068,N_14856,N_13319);
and U18069 (N_18069,N_11149,N_12774);
nor U18070 (N_18070,N_12721,N_11163);
nor U18071 (N_18071,N_11094,N_14609);
nand U18072 (N_18072,N_13745,N_13662);
nor U18073 (N_18073,N_11661,N_13965);
and U18074 (N_18074,N_14446,N_14086);
and U18075 (N_18075,N_11420,N_11504);
nand U18076 (N_18076,N_12636,N_11326);
nand U18077 (N_18077,N_13790,N_10005);
nand U18078 (N_18078,N_11784,N_10825);
nand U18079 (N_18079,N_11809,N_12020);
or U18080 (N_18080,N_12657,N_12434);
or U18081 (N_18081,N_13827,N_14412);
nor U18082 (N_18082,N_13467,N_14762);
xor U18083 (N_18083,N_12876,N_13718);
or U18084 (N_18084,N_14125,N_10105);
nor U18085 (N_18085,N_12272,N_11984);
or U18086 (N_18086,N_14655,N_13845);
nand U18087 (N_18087,N_14896,N_13205);
nand U18088 (N_18088,N_11659,N_14897);
or U18089 (N_18089,N_13314,N_14437);
nor U18090 (N_18090,N_11743,N_14303);
nor U18091 (N_18091,N_12953,N_12451);
nand U18092 (N_18092,N_13946,N_14243);
nand U18093 (N_18093,N_11120,N_10376);
nor U18094 (N_18094,N_14628,N_10416);
and U18095 (N_18095,N_13478,N_10453);
nand U18096 (N_18096,N_11609,N_14915);
xnor U18097 (N_18097,N_11525,N_14957);
or U18098 (N_18098,N_13526,N_13282);
and U18099 (N_18099,N_14801,N_14826);
nand U18100 (N_18100,N_10176,N_14006);
or U18101 (N_18101,N_13912,N_12049);
nor U18102 (N_18102,N_10138,N_11298);
nor U18103 (N_18103,N_11887,N_11503);
nor U18104 (N_18104,N_10795,N_14513);
nor U18105 (N_18105,N_12731,N_14008);
nand U18106 (N_18106,N_13254,N_12263);
nor U18107 (N_18107,N_14937,N_14625);
nand U18108 (N_18108,N_11127,N_10584);
nand U18109 (N_18109,N_12978,N_14296);
or U18110 (N_18110,N_11568,N_12283);
and U18111 (N_18111,N_11263,N_11441);
or U18112 (N_18112,N_14491,N_12894);
nor U18113 (N_18113,N_11192,N_12309);
nand U18114 (N_18114,N_14945,N_12196);
nand U18115 (N_18115,N_11394,N_10271);
or U18116 (N_18116,N_10415,N_13963);
nor U18117 (N_18117,N_11393,N_14245);
nand U18118 (N_18118,N_12735,N_11426);
and U18119 (N_18119,N_12555,N_13222);
or U18120 (N_18120,N_12365,N_12186);
nand U18121 (N_18121,N_10098,N_13933);
xor U18122 (N_18122,N_11025,N_14096);
or U18123 (N_18123,N_13973,N_13591);
nor U18124 (N_18124,N_14008,N_13134);
and U18125 (N_18125,N_13942,N_13154);
or U18126 (N_18126,N_12791,N_13506);
nor U18127 (N_18127,N_12647,N_12352);
nand U18128 (N_18128,N_13802,N_11531);
and U18129 (N_18129,N_14244,N_13725);
nor U18130 (N_18130,N_11967,N_10185);
nor U18131 (N_18131,N_14392,N_14679);
and U18132 (N_18132,N_10228,N_11856);
nand U18133 (N_18133,N_11223,N_11133);
or U18134 (N_18134,N_14503,N_11785);
nor U18135 (N_18135,N_14213,N_10557);
nand U18136 (N_18136,N_10959,N_14331);
or U18137 (N_18137,N_12730,N_10852);
and U18138 (N_18138,N_14659,N_11883);
nor U18139 (N_18139,N_13039,N_12113);
or U18140 (N_18140,N_10657,N_12974);
nand U18141 (N_18141,N_13541,N_13950);
or U18142 (N_18142,N_13374,N_14846);
and U18143 (N_18143,N_14382,N_12217);
nand U18144 (N_18144,N_14234,N_10937);
and U18145 (N_18145,N_13517,N_11384);
and U18146 (N_18146,N_12916,N_11395);
or U18147 (N_18147,N_10200,N_11037);
nor U18148 (N_18148,N_14044,N_11191);
xor U18149 (N_18149,N_12645,N_11342);
nor U18150 (N_18150,N_12842,N_14427);
nand U18151 (N_18151,N_14299,N_14204);
or U18152 (N_18152,N_14960,N_10214);
nand U18153 (N_18153,N_13036,N_14904);
and U18154 (N_18154,N_10498,N_13261);
nand U18155 (N_18155,N_13268,N_12279);
nor U18156 (N_18156,N_10808,N_11049);
nand U18157 (N_18157,N_11768,N_13796);
and U18158 (N_18158,N_13395,N_14051);
or U18159 (N_18159,N_13364,N_12061);
nor U18160 (N_18160,N_12552,N_10851);
nor U18161 (N_18161,N_11325,N_12745);
xor U18162 (N_18162,N_12622,N_11482);
nor U18163 (N_18163,N_11412,N_13851);
nand U18164 (N_18164,N_11986,N_11109);
or U18165 (N_18165,N_14493,N_13996);
and U18166 (N_18166,N_12815,N_14696);
nand U18167 (N_18167,N_12321,N_13180);
nor U18168 (N_18168,N_14784,N_14121);
and U18169 (N_18169,N_12376,N_14980);
xor U18170 (N_18170,N_13450,N_12912);
nand U18171 (N_18171,N_11839,N_11985);
and U18172 (N_18172,N_14382,N_10194);
nor U18173 (N_18173,N_14868,N_11017);
or U18174 (N_18174,N_14702,N_10206);
nand U18175 (N_18175,N_14285,N_11143);
nor U18176 (N_18176,N_14168,N_12940);
nand U18177 (N_18177,N_11686,N_11330);
or U18178 (N_18178,N_11491,N_10620);
nand U18179 (N_18179,N_12658,N_13703);
nor U18180 (N_18180,N_14452,N_10607);
nand U18181 (N_18181,N_11180,N_14806);
or U18182 (N_18182,N_11467,N_12481);
and U18183 (N_18183,N_12764,N_13860);
nand U18184 (N_18184,N_12108,N_13309);
nor U18185 (N_18185,N_10646,N_11848);
and U18186 (N_18186,N_13982,N_10754);
nand U18187 (N_18187,N_13552,N_12015);
or U18188 (N_18188,N_10493,N_12788);
nand U18189 (N_18189,N_11441,N_10509);
xor U18190 (N_18190,N_12542,N_13060);
and U18191 (N_18191,N_13102,N_11457);
and U18192 (N_18192,N_12122,N_14163);
nand U18193 (N_18193,N_12889,N_11490);
nor U18194 (N_18194,N_12305,N_11575);
and U18195 (N_18195,N_13595,N_14524);
nand U18196 (N_18196,N_14305,N_13288);
or U18197 (N_18197,N_10678,N_11751);
and U18198 (N_18198,N_10185,N_13095);
nor U18199 (N_18199,N_13115,N_13331);
nor U18200 (N_18200,N_13890,N_11021);
xnor U18201 (N_18201,N_12773,N_13152);
and U18202 (N_18202,N_12396,N_12763);
nand U18203 (N_18203,N_10693,N_13979);
or U18204 (N_18204,N_10017,N_13192);
nor U18205 (N_18205,N_13876,N_10794);
or U18206 (N_18206,N_10705,N_13169);
nor U18207 (N_18207,N_14427,N_10613);
or U18208 (N_18208,N_14184,N_10701);
or U18209 (N_18209,N_13269,N_10052);
or U18210 (N_18210,N_13391,N_13756);
and U18211 (N_18211,N_13803,N_12775);
and U18212 (N_18212,N_14419,N_14489);
nor U18213 (N_18213,N_12477,N_12717);
nor U18214 (N_18214,N_12089,N_14860);
or U18215 (N_18215,N_10911,N_14110);
and U18216 (N_18216,N_13574,N_11054);
and U18217 (N_18217,N_13800,N_12362);
nor U18218 (N_18218,N_12201,N_11297);
nor U18219 (N_18219,N_11037,N_10453);
or U18220 (N_18220,N_12354,N_11817);
nor U18221 (N_18221,N_14725,N_11344);
nand U18222 (N_18222,N_14989,N_14534);
or U18223 (N_18223,N_11468,N_12859);
and U18224 (N_18224,N_13563,N_14331);
or U18225 (N_18225,N_12360,N_14726);
or U18226 (N_18226,N_12753,N_14087);
nor U18227 (N_18227,N_12282,N_10803);
nor U18228 (N_18228,N_11658,N_14159);
or U18229 (N_18229,N_13755,N_10313);
nand U18230 (N_18230,N_13671,N_13988);
nand U18231 (N_18231,N_10077,N_12168);
nor U18232 (N_18232,N_10522,N_10384);
nand U18233 (N_18233,N_14196,N_11405);
and U18234 (N_18234,N_14875,N_10482);
xor U18235 (N_18235,N_14356,N_14854);
nand U18236 (N_18236,N_11731,N_14663);
or U18237 (N_18237,N_11048,N_14739);
and U18238 (N_18238,N_13751,N_13202);
or U18239 (N_18239,N_10947,N_13160);
and U18240 (N_18240,N_10886,N_13424);
nand U18241 (N_18241,N_12682,N_11027);
nor U18242 (N_18242,N_11821,N_13687);
nand U18243 (N_18243,N_12773,N_13383);
or U18244 (N_18244,N_11712,N_10371);
or U18245 (N_18245,N_10659,N_12457);
and U18246 (N_18246,N_12765,N_13601);
nand U18247 (N_18247,N_12984,N_13480);
or U18248 (N_18248,N_13318,N_13965);
nand U18249 (N_18249,N_12185,N_12132);
and U18250 (N_18250,N_12812,N_14050);
and U18251 (N_18251,N_12286,N_13706);
nand U18252 (N_18252,N_10032,N_14002);
nor U18253 (N_18253,N_10632,N_14192);
and U18254 (N_18254,N_11458,N_14097);
or U18255 (N_18255,N_10280,N_13825);
and U18256 (N_18256,N_10309,N_11379);
and U18257 (N_18257,N_13534,N_13704);
xnor U18258 (N_18258,N_10183,N_12750);
xor U18259 (N_18259,N_10111,N_12494);
nor U18260 (N_18260,N_12464,N_12386);
and U18261 (N_18261,N_13915,N_13562);
nor U18262 (N_18262,N_12532,N_10946);
nand U18263 (N_18263,N_12668,N_14051);
nor U18264 (N_18264,N_13383,N_10452);
nor U18265 (N_18265,N_11154,N_12010);
and U18266 (N_18266,N_13966,N_11488);
or U18267 (N_18267,N_10126,N_13732);
nand U18268 (N_18268,N_11724,N_14706);
and U18269 (N_18269,N_12925,N_13656);
nor U18270 (N_18270,N_12784,N_13822);
and U18271 (N_18271,N_14427,N_14198);
nand U18272 (N_18272,N_12328,N_10255);
or U18273 (N_18273,N_14242,N_12530);
nand U18274 (N_18274,N_14802,N_13639);
nand U18275 (N_18275,N_11615,N_13215);
nor U18276 (N_18276,N_13747,N_13748);
or U18277 (N_18277,N_11755,N_14029);
and U18278 (N_18278,N_10111,N_13794);
nor U18279 (N_18279,N_13476,N_11106);
nor U18280 (N_18280,N_14543,N_12457);
nor U18281 (N_18281,N_14128,N_12687);
and U18282 (N_18282,N_10315,N_13902);
and U18283 (N_18283,N_14599,N_14790);
or U18284 (N_18284,N_11339,N_13554);
or U18285 (N_18285,N_10161,N_10493);
or U18286 (N_18286,N_11133,N_13111);
or U18287 (N_18287,N_14457,N_14155);
nor U18288 (N_18288,N_14443,N_11834);
nor U18289 (N_18289,N_10269,N_11066);
and U18290 (N_18290,N_14641,N_12122);
and U18291 (N_18291,N_14060,N_10060);
nand U18292 (N_18292,N_10182,N_14687);
and U18293 (N_18293,N_10602,N_10302);
nand U18294 (N_18294,N_12935,N_12621);
or U18295 (N_18295,N_11322,N_14614);
xnor U18296 (N_18296,N_14962,N_14218);
and U18297 (N_18297,N_14980,N_12902);
or U18298 (N_18298,N_11680,N_14793);
nand U18299 (N_18299,N_13290,N_13603);
nor U18300 (N_18300,N_13622,N_13949);
or U18301 (N_18301,N_11178,N_11964);
and U18302 (N_18302,N_14089,N_12022);
nor U18303 (N_18303,N_14263,N_11865);
nand U18304 (N_18304,N_13603,N_12450);
nor U18305 (N_18305,N_12674,N_11337);
nor U18306 (N_18306,N_13803,N_14003);
nand U18307 (N_18307,N_11764,N_11179);
and U18308 (N_18308,N_11949,N_12627);
nand U18309 (N_18309,N_11034,N_12246);
nand U18310 (N_18310,N_12422,N_13564);
or U18311 (N_18311,N_12257,N_13291);
and U18312 (N_18312,N_10592,N_12945);
nand U18313 (N_18313,N_10747,N_10193);
and U18314 (N_18314,N_12475,N_10321);
or U18315 (N_18315,N_10403,N_11645);
nand U18316 (N_18316,N_10909,N_11527);
xor U18317 (N_18317,N_14832,N_10432);
or U18318 (N_18318,N_11428,N_14821);
nand U18319 (N_18319,N_10853,N_11836);
or U18320 (N_18320,N_14888,N_11519);
and U18321 (N_18321,N_14626,N_11697);
nor U18322 (N_18322,N_14548,N_13928);
nor U18323 (N_18323,N_12569,N_12898);
nand U18324 (N_18324,N_12481,N_10452);
nand U18325 (N_18325,N_12363,N_13430);
and U18326 (N_18326,N_14389,N_11042);
and U18327 (N_18327,N_11866,N_10048);
and U18328 (N_18328,N_11180,N_13884);
nand U18329 (N_18329,N_12453,N_13535);
nand U18330 (N_18330,N_14282,N_14376);
nand U18331 (N_18331,N_14487,N_13590);
nor U18332 (N_18332,N_12071,N_12896);
and U18333 (N_18333,N_13444,N_14949);
and U18334 (N_18334,N_12401,N_11150);
nand U18335 (N_18335,N_14789,N_12835);
nor U18336 (N_18336,N_14681,N_11996);
nor U18337 (N_18337,N_12456,N_14841);
nand U18338 (N_18338,N_11301,N_13612);
nor U18339 (N_18339,N_13189,N_14589);
or U18340 (N_18340,N_10001,N_10035);
nand U18341 (N_18341,N_13038,N_10580);
and U18342 (N_18342,N_12829,N_12880);
and U18343 (N_18343,N_14478,N_13143);
nand U18344 (N_18344,N_10814,N_12668);
nor U18345 (N_18345,N_13745,N_14308);
nor U18346 (N_18346,N_10218,N_12723);
or U18347 (N_18347,N_12158,N_14891);
or U18348 (N_18348,N_11756,N_13475);
and U18349 (N_18349,N_12458,N_14205);
nand U18350 (N_18350,N_13062,N_13180);
and U18351 (N_18351,N_12402,N_10063);
and U18352 (N_18352,N_11722,N_14428);
or U18353 (N_18353,N_14324,N_11087);
nand U18354 (N_18354,N_13502,N_13465);
nand U18355 (N_18355,N_14926,N_14555);
or U18356 (N_18356,N_11119,N_12501);
or U18357 (N_18357,N_10852,N_10295);
and U18358 (N_18358,N_14482,N_13685);
nor U18359 (N_18359,N_10932,N_14138);
nor U18360 (N_18360,N_11119,N_10040);
nor U18361 (N_18361,N_12002,N_10536);
nand U18362 (N_18362,N_10116,N_10232);
and U18363 (N_18363,N_12833,N_12793);
nand U18364 (N_18364,N_12043,N_12445);
nand U18365 (N_18365,N_13649,N_13864);
nor U18366 (N_18366,N_12995,N_11027);
and U18367 (N_18367,N_12491,N_10162);
or U18368 (N_18368,N_10769,N_10853);
nand U18369 (N_18369,N_10663,N_10391);
nor U18370 (N_18370,N_11210,N_10281);
nor U18371 (N_18371,N_14179,N_10062);
nor U18372 (N_18372,N_11178,N_13932);
nor U18373 (N_18373,N_13149,N_12180);
or U18374 (N_18374,N_14605,N_13671);
or U18375 (N_18375,N_10368,N_14794);
or U18376 (N_18376,N_14522,N_12031);
and U18377 (N_18377,N_14242,N_11588);
or U18378 (N_18378,N_10617,N_13832);
and U18379 (N_18379,N_11771,N_13453);
or U18380 (N_18380,N_12259,N_11040);
or U18381 (N_18381,N_14121,N_12986);
xnor U18382 (N_18382,N_11515,N_10402);
nand U18383 (N_18383,N_14571,N_11942);
or U18384 (N_18384,N_13077,N_12918);
nor U18385 (N_18385,N_11505,N_12101);
nand U18386 (N_18386,N_13707,N_14712);
nor U18387 (N_18387,N_10377,N_13635);
nor U18388 (N_18388,N_11440,N_14223);
nor U18389 (N_18389,N_13590,N_13467);
or U18390 (N_18390,N_12077,N_14816);
and U18391 (N_18391,N_14518,N_11795);
and U18392 (N_18392,N_12698,N_10554);
nand U18393 (N_18393,N_10587,N_10173);
nor U18394 (N_18394,N_13616,N_11813);
nand U18395 (N_18395,N_10087,N_14359);
nor U18396 (N_18396,N_12692,N_10389);
and U18397 (N_18397,N_11283,N_10023);
or U18398 (N_18398,N_13920,N_14987);
and U18399 (N_18399,N_14345,N_13265);
nand U18400 (N_18400,N_14830,N_14838);
or U18401 (N_18401,N_14403,N_13620);
or U18402 (N_18402,N_10439,N_13070);
nor U18403 (N_18403,N_14027,N_13121);
or U18404 (N_18404,N_11076,N_11907);
or U18405 (N_18405,N_13265,N_12883);
and U18406 (N_18406,N_10058,N_11905);
nand U18407 (N_18407,N_12441,N_13970);
xnor U18408 (N_18408,N_11880,N_14998);
nor U18409 (N_18409,N_14965,N_10168);
nand U18410 (N_18410,N_13659,N_11137);
nor U18411 (N_18411,N_13671,N_10265);
or U18412 (N_18412,N_14684,N_11725);
and U18413 (N_18413,N_10873,N_14005);
xor U18414 (N_18414,N_11848,N_12129);
xor U18415 (N_18415,N_10862,N_14098);
nand U18416 (N_18416,N_10416,N_13002);
nand U18417 (N_18417,N_11517,N_13938);
nor U18418 (N_18418,N_14358,N_11197);
nand U18419 (N_18419,N_10209,N_11471);
nand U18420 (N_18420,N_10841,N_14562);
and U18421 (N_18421,N_12103,N_13426);
or U18422 (N_18422,N_12761,N_13355);
nor U18423 (N_18423,N_14852,N_14797);
and U18424 (N_18424,N_12793,N_11126);
nor U18425 (N_18425,N_11888,N_10254);
nor U18426 (N_18426,N_12943,N_13560);
and U18427 (N_18427,N_12700,N_13092);
nand U18428 (N_18428,N_11581,N_10860);
or U18429 (N_18429,N_10102,N_10974);
or U18430 (N_18430,N_12910,N_14064);
and U18431 (N_18431,N_12324,N_10900);
and U18432 (N_18432,N_14822,N_14433);
nand U18433 (N_18433,N_13972,N_13050);
or U18434 (N_18434,N_12354,N_11253);
nor U18435 (N_18435,N_11650,N_14247);
nor U18436 (N_18436,N_10383,N_13470);
nor U18437 (N_18437,N_10485,N_12067);
nor U18438 (N_18438,N_13286,N_12296);
nor U18439 (N_18439,N_14941,N_10542);
nand U18440 (N_18440,N_13740,N_12181);
nor U18441 (N_18441,N_10741,N_10140);
nor U18442 (N_18442,N_12817,N_10567);
nand U18443 (N_18443,N_14409,N_14482);
nor U18444 (N_18444,N_10040,N_12644);
nand U18445 (N_18445,N_13910,N_11159);
nor U18446 (N_18446,N_14657,N_10656);
xor U18447 (N_18447,N_14172,N_14452);
nor U18448 (N_18448,N_12690,N_12742);
or U18449 (N_18449,N_13881,N_13082);
nor U18450 (N_18450,N_11695,N_12717);
nand U18451 (N_18451,N_14679,N_14918);
nand U18452 (N_18452,N_13208,N_10463);
and U18453 (N_18453,N_12977,N_11575);
nor U18454 (N_18454,N_13999,N_11650);
or U18455 (N_18455,N_10880,N_11152);
nand U18456 (N_18456,N_13762,N_13313);
and U18457 (N_18457,N_11786,N_12537);
and U18458 (N_18458,N_14267,N_10702);
or U18459 (N_18459,N_12907,N_10906);
nand U18460 (N_18460,N_14571,N_12373);
or U18461 (N_18461,N_13600,N_10941);
nand U18462 (N_18462,N_13376,N_10710);
nor U18463 (N_18463,N_14774,N_14838);
and U18464 (N_18464,N_10628,N_10303);
xnor U18465 (N_18465,N_14162,N_10088);
or U18466 (N_18466,N_11561,N_13971);
and U18467 (N_18467,N_14709,N_12790);
nor U18468 (N_18468,N_10975,N_12452);
nand U18469 (N_18469,N_14082,N_11228);
and U18470 (N_18470,N_14124,N_11292);
or U18471 (N_18471,N_11631,N_11601);
nand U18472 (N_18472,N_11579,N_14849);
nand U18473 (N_18473,N_13191,N_13084);
nor U18474 (N_18474,N_10990,N_12794);
or U18475 (N_18475,N_12307,N_14392);
and U18476 (N_18476,N_14264,N_11969);
and U18477 (N_18477,N_12996,N_11429);
and U18478 (N_18478,N_11552,N_13005);
and U18479 (N_18479,N_13912,N_10950);
and U18480 (N_18480,N_13265,N_11618);
nand U18481 (N_18481,N_12403,N_10697);
nand U18482 (N_18482,N_14771,N_10183);
nand U18483 (N_18483,N_14041,N_13032);
and U18484 (N_18484,N_11800,N_11240);
xor U18485 (N_18485,N_10428,N_11431);
and U18486 (N_18486,N_13812,N_14791);
and U18487 (N_18487,N_13547,N_13553);
and U18488 (N_18488,N_10068,N_13980);
or U18489 (N_18489,N_13712,N_13890);
and U18490 (N_18490,N_12776,N_10275);
and U18491 (N_18491,N_11282,N_11939);
nor U18492 (N_18492,N_11583,N_12430);
xnor U18493 (N_18493,N_10299,N_11269);
nand U18494 (N_18494,N_12272,N_11132);
nor U18495 (N_18495,N_12543,N_13151);
and U18496 (N_18496,N_12244,N_13248);
and U18497 (N_18497,N_14613,N_11624);
nor U18498 (N_18498,N_12294,N_13276);
nor U18499 (N_18499,N_14842,N_10422);
or U18500 (N_18500,N_10767,N_11709);
nand U18501 (N_18501,N_10832,N_14187);
nand U18502 (N_18502,N_12679,N_11009);
nand U18503 (N_18503,N_13725,N_14828);
and U18504 (N_18504,N_13376,N_11761);
nand U18505 (N_18505,N_13278,N_13966);
and U18506 (N_18506,N_14588,N_11865);
and U18507 (N_18507,N_13470,N_12658);
nor U18508 (N_18508,N_14780,N_12970);
and U18509 (N_18509,N_13553,N_13739);
or U18510 (N_18510,N_14946,N_13008);
nand U18511 (N_18511,N_13601,N_11195);
nand U18512 (N_18512,N_12437,N_14818);
xnor U18513 (N_18513,N_12867,N_13092);
nor U18514 (N_18514,N_14841,N_12830);
and U18515 (N_18515,N_14510,N_13726);
or U18516 (N_18516,N_10914,N_12295);
or U18517 (N_18517,N_11558,N_11166);
and U18518 (N_18518,N_10129,N_10654);
or U18519 (N_18519,N_13026,N_11919);
and U18520 (N_18520,N_10022,N_10331);
nand U18521 (N_18521,N_11163,N_14825);
nand U18522 (N_18522,N_11694,N_12768);
nand U18523 (N_18523,N_10222,N_10230);
nand U18524 (N_18524,N_13601,N_14122);
and U18525 (N_18525,N_14008,N_11960);
or U18526 (N_18526,N_13606,N_10122);
and U18527 (N_18527,N_13523,N_13878);
nand U18528 (N_18528,N_12047,N_12983);
nor U18529 (N_18529,N_12207,N_11036);
nand U18530 (N_18530,N_11272,N_10832);
or U18531 (N_18531,N_11278,N_14894);
nor U18532 (N_18532,N_12572,N_12133);
nand U18533 (N_18533,N_14104,N_12336);
nand U18534 (N_18534,N_14090,N_10032);
and U18535 (N_18535,N_14215,N_11220);
and U18536 (N_18536,N_12151,N_13908);
nand U18537 (N_18537,N_11113,N_13214);
nand U18538 (N_18538,N_11302,N_14021);
nor U18539 (N_18539,N_12770,N_12882);
nor U18540 (N_18540,N_12905,N_10126);
or U18541 (N_18541,N_11013,N_10032);
nand U18542 (N_18542,N_10994,N_10252);
nand U18543 (N_18543,N_14770,N_12792);
nand U18544 (N_18544,N_12035,N_13571);
and U18545 (N_18545,N_10243,N_12328);
nand U18546 (N_18546,N_11483,N_10650);
or U18547 (N_18547,N_11108,N_10308);
or U18548 (N_18548,N_12516,N_10135);
and U18549 (N_18549,N_12070,N_12854);
or U18550 (N_18550,N_14406,N_11992);
or U18551 (N_18551,N_12579,N_13567);
nor U18552 (N_18552,N_11505,N_13344);
and U18553 (N_18553,N_12386,N_11606);
and U18554 (N_18554,N_10971,N_12182);
nand U18555 (N_18555,N_14952,N_10942);
nor U18556 (N_18556,N_13189,N_14039);
or U18557 (N_18557,N_12208,N_13145);
nand U18558 (N_18558,N_14033,N_10292);
nor U18559 (N_18559,N_14323,N_13335);
or U18560 (N_18560,N_10956,N_13274);
nor U18561 (N_18561,N_10529,N_14748);
nand U18562 (N_18562,N_11797,N_14303);
xnor U18563 (N_18563,N_12860,N_13070);
nor U18564 (N_18564,N_13793,N_12191);
nand U18565 (N_18565,N_12006,N_14477);
or U18566 (N_18566,N_10626,N_14935);
or U18567 (N_18567,N_13904,N_12872);
or U18568 (N_18568,N_11801,N_11968);
nand U18569 (N_18569,N_14179,N_12665);
and U18570 (N_18570,N_12225,N_11367);
and U18571 (N_18571,N_10162,N_11833);
and U18572 (N_18572,N_10204,N_14666);
nor U18573 (N_18573,N_11103,N_14612);
or U18574 (N_18574,N_12545,N_10645);
or U18575 (N_18575,N_13718,N_12853);
or U18576 (N_18576,N_14572,N_11117);
nand U18577 (N_18577,N_13627,N_12626);
nor U18578 (N_18578,N_10060,N_12812);
nor U18579 (N_18579,N_14321,N_13547);
nor U18580 (N_18580,N_10609,N_10035);
or U18581 (N_18581,N_10545,N_12671);
nor U18582 (N_18582,N_13533,N_13028);
nand U18583 (N_18583,N_11927,N_14168);
nand U18584 (N_18584,N_14945,N_11267);
nand U18585 (N_18585,N_14183,N_12019);
and U18586 (N_18586,N_14602,N_13014);
nand U18587 (N_18587,N_12130,N_10484);
and U18588 (N_18588,N_12095,N_10669);
and U18589 (N_18589,N_13429,N_10026);
or U18590 (N_18590,N_14774,N_11534);
nor U18591 (N_18591,N_14433,N_11297);
or U18592 (N_18592,N_12292,N_14637);
or U18593 (N_18593,N_11873,N_14389);
nand U18594 (N_18594,N_10697,N_10938);
and U18595 (N_18595,N_10947,N_12362);
and U18596 (N_18596,N_12895,N_10491);
nor U18597 (N_18597,N_11757,N_10438);
or U18598 (N_18598,N_10122,N_11391);
and U18599 (N_18599,N_13759,N_12715);
or U18600 (N_18600,N_12182,N_11878);
and U18601 (N_18601,N_14405,N_10232);
or U18602 (N_18602,N_11364,N_10811);
and U18603 (N_18603,N_10853,N_11758);
or U18604 (N_18604,N_12501,N_11699);
and U18605 (N_18605,N_10667,N_11863);
and U18606 (N_18606,N_13685,N_10589);
nor U18607 (N_18607,N_10977,N_13162);
nand U18608 (N_18608,N_12355,N_11156);
and U18609 (N_18609,N_10341,N_12019);
nand U18610 (N_18610,N_10368,N_11385);
xor U18611 (N_18611,N_14076,N_14686);
and U18612 (N_18612,N_10061,N_12113);
nand U18613 (N_18613,N_12754,N_13542);
nor U18614 (N_18614,N_12892,N_14726);
nor U18615 (N_18615,N_11224,N_13168);
nand U18616 (N_18616,N_10669,N_13139);
and U18617 (N_18617,N_14685,N_11312);
and U18618 (N_18618,N_11086,N_12791);
and U18619 (N_18619,N_13641,N_11969);
and U18620 (N_18620,N_12170,N_13757);
nand U18621 (N_18621,N_14146,N_10212);
nor U18622 (N_18622,N_12720,N_10809);
nand U18623 (N_18623,N_12495,N_11697);
or U18624 (N_18624,N_12282,N_14822);
or U18625 (N_18625,N_14281,N_11665);
nand U18626 (N_18626,N_10803,N_12232);
and U18627 (N_18627,N_13789,N_10484);
and U18628 (N_18628,N_13973,N_11726);
nand U18629 (N_18629,N_14498,N_10720);
nor U18630 (N_18630,N_11524,N_13719);
nand U18631 (N_18631,N_10160,N_11252);
and U18632 (N_18632,N_14443,N_12774);
nor U18633 (N_18633,N_11878,N_13284);
and U18634 (N_18634,N_13741,N_14437);
nand U18635 (N_18635,N_11976,N_11474);
or U18636 (N_18636,N_10895,N_10769);
nor U18637 (N_18637,N_12920,N_11518);
and U18638 (N_18638,N_12440,N_14288);
or U18639 (N_18639,N_13200,N_11737);
or U18640 (N_18640,N_12093,N_12916);
and U18641 (N_18641,N_11220,N_10172);
nor U18642 (N_18642,N_11767,N_11736);
nand U18643 (N_18643,N_12196,N_10540);
nand U18644 (N_18644,N_13417,N_12804);
or U18645 (N_18645,N_11327,N_13526);
nand U18646 (N_18646,N_14018,N_14951);
nor U18647 (N_18647,N_11832,N_12060);
nor U18648 (N_18648,N_11895,N_14305);
or U18649 (N_18649,N_13778,N_10840);
or U18650 (N_18650,N_14121,N_13676);
and U18651 (N_18651,N_10919,N_14618);
nand U18652 (N_18652,N_11344,N_11336);
nand U18653 (N_18653,N_11174,N_10292);
and U18654 (N_18654,N_13502,N_14403);
and U18655 (N_18655,N_10121,N_12989);
nand U18656 (N_18656,N_13246,N_11566);
or U18657 (N_18657,N_12557,N_14090);
nor U18658 (N_18658,N_14624,N_14986);
or U18659 (N_18659,N_13651,N_14855);
xnor U18660 (N_18660,N_13664,N_10042);
or U18661 (N_18661,N_10486,N_12606);
nor U18662 (N_18662,N_11315,N_11967);
or U18663 (N_18663,N_14018,N_12738);
or U18664 (N_18664,N_12661,N_13965);
nor U18665 (N_18665,N_13689,N_14452);
or U18666 (N_18666,N_14656,N_12141);
and U18667 (N_18667,N_10501,N_14305);
and U18668 (N_18668,N_10910,N_13081);
or U18669 (N_18669,N_11195,N_13837);
nor U18670 (N_18670,N_10526,N_12505);
nand U18671 (N_18671,N_12863,N_12474);
and U18672 (N_18672,N_13963,N_12457);
xor U18673 (N_18673,N_10668,N_11346);
or U18674 (N_18674,N_13620,N_14515);
nor U18675 (N_18675,N_10818,N_10947);
nand U18676 (N_18676,N_13469,N_14266);
or U18677 (N_18677,N_10248,N_14384);
nand U18678 (N_18678,N_13555,N_10179);
and U18679 (N_18679,N_11383,N_13797);
or U18680 (N_18680,N_10259,N_11096);
xnor U18681 (N_18681,N_14127,N_14512);
and U18682 (N_18682,N_12993,N_10459);
nand U18683 (N_18683,N_13043,N_13954);
and U18684 (N_18684,N_13092,N_11391);
nor U18685 (N_18685,N_12610,N_14377);
and U18686 (N_18686,N_10635,N_10480);
or U18687 (N_18687,N_11105,N_13527);
or U18688 (N_18688,N_10481,N_11781);
and U18689 (N_18689,N_12530,N_12453);
xor U18690 (N_18690,N_12418,N_11673);
or U18691 (N_18691,N_12023,N_12667);
or U18692 (N_18692,N_13100,N_14856);
nor U18693 (N_18693,N_10285,N_10286);
nand U18694 (N_18694,N_14159,N_13356);
and U18695 (N_18695,N_10573,N_14421);
nand U18696 (N_18696,N_11930,N_14686);
and U18697 (N_18697,N_10379,N_10675);
and U18698 (N_18698,N_11133,N_11194);
xnor U18699 (N_18699,N_14491,N_12597);
or U18700 (N_18700,N_12554,N_12922);
or U18701 (N_18701,N_10038,N_13463);
or U18702 (N_18702,N_12779,N_12034);
or U18703 (N_18703,N_12699,N_14023);
and U18704 (N_18704,N_10838,N_14999);
and U18705 (N_18705,N_13784,N_12506);
nor U18706 (N_18706,N_13864,N_11799);
and U18707 (N_18707,N_10183,N_11066);
nor U18708 (N_18708,N_12711,N_10612);
or U18709 (N_18709,N_11977,N_12040);
and U18710 (N_18710,N_14857,N_14907);
nand U18711 (N_18711,N_12063,N_11390);
nand U18712 (N_18712,N_14861,N_13533);
nor U18713 (N_18713,N_13484,N_13379);
nand U18714 (N_18714,N_13470,N_13185);
and U18715 (N_18715,N_10298,N_13331);
and U18716 (N_18716,N_14586,N_12790);
xnor U18717 (N_18717,N_14811,N_13628);
nand U18718 (N_18718,N_13109,N_12875);
nand U18719 (N_18719,N_12444,N_12861);
and U18720 (N_18720,N_14111,N_13071);
or U18721 (N_18721,N_11985,N_14176);
and U18722 (N_18722,N_10084,N_10231);
or U18723 (N_18723,N_14862,N_14059);
nand U18724 (N_18724,N_11373,N_14272);
nor U18725 (N_18725,N_11980,N_14152);
nor U18726 (N_18726,N_11478,N_12122);
xnor U18727 (N_18727,N_14901,N_10816);
xor U18728 (N_18728,N_14077,N_13194);
nand U18729 (N_18729,N_13388,N_14688);
and U18730 (N_18730,N_14762,N_12924);
nand U18731 (N_18731,N_10813,N_14680);
nand U18732 (N_18732,N_11308,N_10083);
nand U18733 (N_18733,N_12035,N_13127);
or U18734 (N_18734,N_12611,N_10956);
nand U18735 (N_18735,N_14688,N_14741);
or U18736 (N_18736,N_13658,N_13290);
and U18737 (N_18737,N_13620,N_14309);
xor U18738 (N_18738,N_14715,N_13799);
nand U18739 (N_18739,N_14376,N_11713);
or U18740 (N_18740,N_10262,N_11752);
nor U18741 (N_18741,N_13443,N_10560);
and U18742 (N_18742,N_11566,N_14308);
or U18743 (N_18743,N_10772,N_12043);
and U18744 (N_18744,N_11809,N_13041);
nand U18745 (N_18745,N_11922,N_11513);
and U18746 (N_18746,N_14054,N_10291);
nand U18747 (N_18747,N_10930,N_11026);
or U18748 (N_18748,N_13552,N_10355);
and U18749 (N_18749,N_14386,N_12725);
or U18750 (N_18750,N_11319,N_12375);
nor U18751 (N_18751,N_12868,N_11487);
nand U18752 (N_18752,N_13611,N_10687);
or U18753 (N_18753,N_13247,N_14091);
or U18754 (N_18754,N_14747,N_14752);
nand U18755 (N_18755,N_10974,N_13062);
nor U18756 (N_18756,N_14326,N_12841);
or U18757 (N_18757,N_11437,N_12269);
nor U18758 (N_18758,N_14244,N_12104);
nor U18759 (N_18759,N_14683,N_14848);
or U18760 (N_18760,N_14840,N_13751);
nor U18761 (N_18761,N_14962,N_11954);
or U18762 (N_18762,N_12935,N_12217);
or U18763 (N_18763,N_10869,N_12645);
nand U18764 (N_18764,N_13902,N_10795);
nand U18765 (N_18765,N_14625,N_12117);
and U18766 (N_18766,N_10165,N_12549);
or U18767 (N_18767,N_14719,N_14622);
and U18768 (N_18768,N_13307,N_10731);
nor U18769 (N_18769,N_10303,N_14287);
and U18770 (N_18770,N_13609,N_13257);
nor U18771 (N_18771,N_11905,N_13868);
nor U18772 (N_18772,N_11935,N_11760);
nor U18773 (N_18773,N_10118,N_13370);
nand U18774 (N_18774,N_11182,N_13186);
xor U18775 (N_18775,N_12084,N_12584);
and U18776 (N_18776,N_12272,N_10317);
xor U18777 (N_18777,N_10641,N_14483);
or U18778 (N_18778,N_10247,N_10774);
and U18779 (N_18779,N_14514,N_14430);
and U18780 (N_18780,N_12490,N_13158);
nand U18781 (N_18781,N_13716,N_14516);
or U18782 (N_18782,N_11859,N_13353);
nor U18783 (N_18783,N_12225,N_11009);
or U18784 (N_18784,N_14421,N_14941);
and U18785 (N_18785,N_11160,N_14571);
nand U18786 (N_18786,N_13586,N_13475);
xor U18787 (N_18787,N_13883,N_10751);
nor U18788 (N_18788,N_14502,N_10697);
and U18789 (N_18789,N_11585,N_12956);
nand U18790 (N_18790,N_11815,N_12020);
or U18791 (N_18791,N_13085,N_10884);
or U18792 (N_18792,N_10205,N_13742);
nand U18793 (N_18793,N_10627,N_11731);
nand U18794 (N_18794,N_12936,N_12128);
nor U18795 (N_18795,N_13924,N_11117);
or U18796 (N_18796,N_14974,N_10585);
or U18797 (N_18797,N_13642,N_12895);
nor U18798 (N_18798,N_13070,N_12330);
nand U18799 (N_18799,N_13095,N_13553);
or U18800 (N_18800,N_10208,N_11829);
nand U18801 (N_18801,N_11916,N_12507);
nor U18802 (N_18802,N_12328,N_11798);
or U18803 (N_18803,N_13955,N_14114);
nor U18804 (N_18804,N_14365,N_13193);
or U18805 (N_18805,N_14586,N_14727);
nand U18806 (N_18806,N_13230,N_11019);
nor U18807 (N_18807,N_10218,N_10891);
nor U18808 (N_18808,N_10346,N_13206);
nor U18809 (N_18809,N_10208,N_14329);
or U18810 (N_18810,N_11964,N_10740);
nor U18811 (N_18811,N_14314,N_10770);
nor U18812 (N_18812,N_10286,N_10199);
and U18813 (N_18813,N_13688,N_14255);
or U18814 (N_18814,N_11230,N_12527);
and U18815 (N_18815,N_13044,N_10508);
or U18816 (N_18816,N_12653,N_13023);
or U18817 (N_18817,N_14950,N_11310);
and U18818 (N_18818,N_11332,N_11896);
and U18819 (N_18819,N_12550,N_12447);
nor U18820 (N_18820,N_14052,N_11164);
nand U18821 (N_18821,N_14254,N_10675);
and U18822 (N_18822,N_14130,N_13338);
nor U18823 (N_18823,N_14114,N_14231);
or U18824 (N_18824,N_12695,N_13647);
and U18825 (N_18825,N_11166,N_11235);
nand U18826 (N_18826,N_11362,N_10370);
nor U18827 (N_18827,N_14577,N_10072);
nor U18828 (N_18828,N_13033,N_11874);
and U18829 (N_18829,N_11176,N_14122);
or U18830 (N_18830,N_10162,N_11430);
or U18831 (N_18831,N_10973,N_10139);
nor U18832 (N_18832,N_10737,N_14487);
xor U18833 (N_18833,N_10065,N_14950);
nand U18834 (N_18834,N_13090,N_10125);
nand U18835 (N_18835,N_10661,N_14852);
nor U18836 (N_18836,N_11211,N_11940);
nor U18837 (N_18837,N_10599,N_12346);
nand U18838 (N_18838,N_14453,N_10815);
nand U18839 (N_18839,N_14008,N_13570);
and U18840 (N_18840,N_12325,N_10478);
or U18841 (N_18841,N_14942,N_14842);
xor U18842 (N_18842,N_11758,N_11036);
nor U18843 (N_18843,N_11250,N_10276);
and U18844 (N_18844,N_11805,N_10659);
nand U18845 (N_18845,N_14008,N_14566);
or U18846 (N_18846,N_10059,N_14139);
and U18847 (N_18847,N_12429,N_14225);
nor U18848 (N_18848,N_13107,N_14448);
xnor U18849 (N_18849,N_10119,N_10066);
nand U18850 (N_18850,N_14772,N_10016);
nand U18851 (N_18851,N_14273,N_13512);
nand U18852 (N_18852,N_12395,N_12690);
nand U18853 (N_18853,N_11793,N_11106);
nand U18854 (N_18854,N_11702,N_13205);
and U18855 (N_18855,N_10252,N_13425);
and U18856 (N_18856,N_14388,N_14048);
and U18857 (N_18857,N_12912,N_11389);
nand U18858 (N_18858,N_14792,N_14222);
nor U18859 (N_18859,N_12132,N_12171);
nor U18860 (N_18860,N_11068,N_14091);
or U18861 (N_18861,N_13872,N_10175);
nor U18862 (N_18862,N_11495,N_14878);
and U18863 (N_18863,N_13589,N_14350);
or U18864 (N_18864,N_10871,N_12660);
nand U18865 (N_18865,N_11491,N_12757);
nor U18866 (N_18866,N_11500,N_10676);
xnor U18867 (N_18867,N_10148,N_13036);
nor U18868 (N_18868,N_11342,N_10574);
and U18869 (N_18869,N_14272,N_11621);
nor U18870 (N_18870,N_13346,N_10191);
nand U18871 (N_18871,N_10504,N_11172);
nand U18872 (N_18872,N_12553,N_14996);
and U18873 (N_18873,N_12764,N_10005);
and U18874 (N_18874,N_12008,N_12029);
or U18875 (N_18875,N_10747,N_10041);
and U18876 (N_18876,N_10849,N_11165);
or U18877 (N_18877,N_12686,N_12652);
nand U18878 (N_18878,N_10588,N_11995);
or U18879 (N_18879,N_14486,N_13421);
nor U18880 (N_18880,N_13294,N_14754);
xnor U18881 (N_18881,N_13062,N_13296);
nand U18882 (N_18882,N_13015,N_11699);
and U18883 (N_18883,N_12538,N_11254);
and U18884 (N_18884,N_11553,N_13100);
and U18885 (N_18885,N_11725,N_10810);
nand U18886 (N_18886,N_12308,N_12411);
nor U18887 (N_18887,N_13752,N_10101);
nor U18888 (N_18888,N_10967,N_12637);
or U18889 (N_18889,N_11987,N_12874);
and U18890 (N_18890,N_14162,N_12789);
and U18891 (N_18891,N_11607,N_14373);
nor U18892 (N_18892,N_10669,N_11270);
nand U18893 (N_18893,N_13071,N_12573);
nand U18894 (N_18894,N_13709,N_13467);
nand U18895 (N_18895,N_10590,N_12801);
nand U18896 (N_18896,N_12488,N_10899);
and U18897 (N_18897,N_14170,N_13000);
or U18898 (N_18898,N_12434,N_10888);
nand U18899 (N_18899,N_12011,N_11649);
and U18900 (N_18900,N_11623,N_13392);
nor U18901 (N_18901,N_13268,N_10428);
nand U18902 (N_18902,N_10145,N_12635);
nor U18903 (N_18903,N_11531,N_10509);
or U18904 (N_18904,N_13447,N_10427);
nor U18905 (N_18905,N_11885,N_13666);
nand U18906 (N_18906,N_12080,N_10395);
nor U18907 (N_18907,N_10145,N_10374);
nor U18908 (N_18908,N_11009,N_11381);
and U18909 (N_18909,N_13896,N_12549);
xnor U18910 (N_18910,N_10573,N_11510);
nor U18911 (N_18911,N_14279,N_13384);
nand U18912 (N_18912,N_13267,N_13460);
nand U18913 (N_18913,N_12465,N_10788);
or U18914 (N_18914,N_11942,N_10329);
nand U18915 (N_18915,N_10621,N_14877);
nand U18916 (N_18916,N_14968,N_12995);
nor U18917 (N_18917,N_12665,N_10486);
nand U18918 (N_18918,N_12403,N_13901);
or U18919 (N_18919,N_13940,N_11626);
or U18920 (N_18920,N_11091,N_11790);
nor U18921 (N_18921,N_14828,N_11394);
or U18922 (N_18922,N_10690,N_14987);
nor U18923 (N_18923,N_12617,N_14267);
and U18924 (N_18924,N_10923,N_11576);
nor U18925 (N_18925,N_14539,N_12576);
nand U18926 (N_18926,N_12065,N_11581);
or U18927 (N_18927,N_13965,N_10516);
nand U18928 (N_18928,N_10652,N_11328);
nor U18929 (N_18929,N_11069,N_12069);
or U18930 (N_18930,N_10996,N_13261);
or U18931 (N_18931,N_10964,N_14407);
and U18932 (N_18932,N_12112,N_10037);
or U18933 (N_18933,N_12673,N_12107);
nor U18934 (N_18934,N_13832,N_14221);
nand U18935 (N_18935,N_10689,N_11106);
nand U18936 (N_18936,N_11196,N_10343);
nand U18937 (N_18937,N_12962,N_12971);
or U18938 (N_18938,N_11229,N_14550);
nor U18939 (N_18939,N_10985,N_11629);
nor U18940 (N_18940,N_12411,N_13206);
nor U18941 (N_18941,N_12811,N_12305);
nor U18942 (N_18942,N_11729,N_12509);
nand U18943 (N_18943,N_13188,N_12473);
nor U18944 (N_18944,N_13666,N_12209);
nor U18945 (N_18945,N_13797,N_14872);
and U18946 (N_18946,N_13466,N_10691);
nand U18947 (N_18947,N_10119,N_13094);
nor U18948 (N_18948,N_13666,N_14196);
and U18949 (N_18949,N_12534,N_11356);
and U18950 (N_18950,N_11089,N_12574);
and U18951 (N_18951,N_11101,N_14411);
and U18952 (N_18952,N_10506,N_10309);
and U18953 (N_18953,N_13490,N_12895);
or U18954 (N_18954,N_14727,N_11193);
or U18955 (N_18955,N_10519,N_14011);
nor U18956 (N_18956,N_13196,N_12554);
nor U18957 (N_18957,N_12734,N_13184);
nor U18958 (N_18958,N_12087,N_13265);
or U18959 (N_18959,N_14532,N_12237);
nand U18960 (N_18960,N_10341,N_10727);
and U18961 (N_18961,N_13633,N_11458);
or U18962 (N_18962,N_11254,N_14066);
or U18963 (N_18963,N_13600,N_13947);
and U18964 (N_18964,N_11654,N_14696);
and U18965 (N_18965,N_13129,N_12722);
or U18966 (N_18966,N_14364,N_14464);
and U18967 (N_18967,N_12653,N_11065);
and U18968 (N_18968,N_12615,N_10524);
nand U18969 (N_18969,N_14645,N_12268);
nor U18970 (N_18970,N_14242,N_10600);
and U18971 (N_18971,N_11455,N_10319);
and U18972 (N_18972,N_12586,N_12212);
nor U18973 (N_18973,N_12325,N_13398);
nand U18974 (N_18974,N_14978,N_12300);
nor U18975 (N_18975,N_11090,N_13931);
nor U18976 (N_18976,N_10868,N_12724);
and U18977 (N_18977,N_14061,N_13931);
and U18978 (N_18978,N_12502,N_10142);
nor U18979 (N_18979,N_14809,N_11613);
nand U18980 (N_18980,N_13631,N_11133);
nor U18981 (N_18981,N_10810,N_11755);
or U18982 (N_18982,N_13834,N_14666);
nand U18983 (N_18983,N_12481,N_14837);
or U18984 (N_18984,N_10258,N_12961);
and U18985 (N_18985,N_14832,N_14857);
nor U18986 (N_18986,N_12520,N_10083);
and U18987 (N_18987,N_11844,N_11817);
and U18988 (N_18988,N_11359,N_12910);
nor U18989 (N_18989,N_13069,N_13703);
and U18990 (N_18990,N_12473,N_12511);
nor U18991 (N_18991,N_12231,N_14597);
nor U18992 (N_18992,N_13239,N_10073);
nor U18993 (N_18993,N_10845,N_11491);
nor U18994 (N_18994,N_11984,N_11873);
and U18995 (N_18995,N_13815,N_12092);
nand U18996 (N_18996,N_12493,N_12886);
and U18997 (N_18997,N_11440,N_11573);
nand U18998 (N_18998,N_12840,N_11141);
nor U18999 (N_18999,N_11444,N_11805);
nor U19000 (N_19000,N_14918,N_10703);
nand U19001 (N_19001,N_13738,N_11296);
nor U19002 (N_19002,N_14069,N_12503);
nand U19003 (N_19003,N_10600,N_14131);
nand U19004 (N_19004,N_11625,N_12093);
nor U19005 (N_19005,N_12038,N_12970);
and U19006 (N_19006,N_12822,N_14747);
nand U19007 (N_19007,N_11858,N_13367);
nand U19008 (N_19008,N_14998,N_12296);
and U19009 (N_19009,N_11761,N_14131);
nand U19010 (N_19010,N_13230,N_11735);
nor U19011 (N_19011,N_10097,N_12639);
and U19012 (N_19012,N_11782,N_14024);
nor U19013 (N_19013,N_13668,N_11222);
and U19014 (N_19014,N_14465,N_11459);
nor U19015 (N_19015,N_10880,N_11268);
or U19016 (N_19016,N_13278,N_14531);
nand U19017 (N_19017,N_10258,N_13431);
or U19018 (N_19018,N_10435,N_14129);
or U19019 (N_19019,N_13543,N_12025);
or U19020 (N_19020,N_12714,N_14819);
nor U19021 (N_19021,N_13063,N_14735);
and U19022 (N_19022,N_10566,N_10367);
nand U19023 (N_19023,N_11009,N_11136);
nand U19024 (N_19024,N_12111,N_11090);
or U19025 (N_19025,N_13066,N_13336);
or U19026 (N_19026,N_14523,N_13001);
or U19027 (N_19027,N_13177,N_11301);
and U19028 (N_19028,N_14389,N_11203);
nor U19029 (N_19029,N_14542,N_14903);
and U19030 (N_19030,N_10969,N_14977);
and U19031 (N_19031,N_11514,N_14985);
and U19032 (N_19032,N_11351,N_12524);
and U19033 (N_19033,N_14168,N_13956);
nand U19034 (N_19034,N_13141,N_10341);
or U19035 (N_19035,N_11811,N_13095);
and U19036 (N_19036,N_14407,N_11304);
and U19037 (N_19037,N_10689,N_14107);
nand U19038 (N_19038,N_12278,N_12427);
nand U19039 (N_19039,N_10399,N_11272);
nand U19040 (N_19040,N_10902,N_14485);
nor U19041 (N_19041,N_13213,N_12439);
or U19042 (N_19042,N_11884,N_14534);
or U19043 (N_19043,N_13520,N_12119);
nor U19044 (N_19044,N_14483,N_10765);
or U19045 (N_19045,N_12120,N_12583);
nor U19046 (N_19046,N_10964,N_13527);
nand U19047 (N_19047,N_12987,N_12792);
nor U19048 (N_19048,N_14238,N_13960);
nand U19049 (N_19049,N_14626,N_10790);
or U19050 (N_19050,N_14954,N_14207);
and U19051 (N_19051,N_12575,N_11721);
nand U19052 (N_19052,N_10090,N_12965);
nor U19053 (N_19053,N_13879,N_10809);
and U19054 (N_19054,N_11256,N_12339);
nor U19055 (N_19055,N_14753,N_13488);
nor U19056 (N_19056,N_11431,N_11395);
nand U19057 (N_19057,N_11872,N_11617);
nand U19058 (N_19058,N_11646,N_10514);
nor U19059 (N_19059,N_10805,N_13181);
and U19060 (N_19060,N_11936,N_14001);
or U19061 (N_19061,N_14352,N_11983);
or U19062 (N_19062,N_13275,N_14624);
nor U19063 (N_19063,N_13071,N_13035);
nor U19064 (N_19064,N_12282,N_14078);
xor U19065 (N_19065,N_14029,N_13815);
or U19066 (N_19066,N_11602,N_13751);
nor U19067 (N_19067,N_12526,N_13835);
and U19068 (N_19068,N_12973,N_10306);
or U19069 (N_19069,N_11193,N_11871);
xnor U19070 (N_19070,N_10518,N_12046);
nor U19071 (N_19071,N_13798,N_13750);
or U19072 (N_19072,N_14510,N_11537);
and U19073 (N_19073,N_12126,N_14870);
nand U19074 (N_19074,N_14039,N_11778);
nor U19075 (N_19075,N_14497,N_13346);
and U19076 (N_19076,N_10753,N_11902);
nand U19077 (N_19077,N_13271,N_10902);
xnor U19078 (N_19078,N_11476,N_10455);
nor U19079 (N_19079,N_14059,N_11737);
nand U19080 (N_19080,N_10557,N_10839);
nand U19081 (N_19081,N_13669,N_10017);
and U19082 (N_19082,N_14741,N_10811);
or U19083 (N_19083,N_14715,N_12584);
and U19084 (N_19084,N_11306,N_13364);
or U19085 (N_19085,N_10797,N_12783);
nor U19086 (N_19086,N_10928,N_10142);
nand U19087 (N_19087,N_11916,N_11450);
nand U19088 (N_19088,N_13873,N_14872);
nor U19089 (N_19089,N_14964,N_14919);
and U19090 (N_19090,N_12499,N_13071);
nand U19091 (N_19091,N_10759,N_12963);
or U19092 (N_19092,N_12272,N_10643);
and U19093 (N_19093,N_13944,N_11023);
or U19094 (N_19094,N_13031,N_12149);
nand U19095 (N_19095,N_12285,N_11271);
and U19096 (N_19096,N_11994,N_14463);
or U19097 (N_19097,N_13908,N_13793);
and U19098 (N_19098,N_13308,N_14477);
nor U19099 (N_19099,N_10493,N_12702);
nand U19100 (N_19100,N_13625,N_10403);
or U19101 (N_19101,N_14154,N_11187);
nand U19102 (N_19102,N_13465,N_11760);
nand U19103 (N_19103,N_10143,N_13029);
nor U19104 (N_19104,N_10764,N_14192);
and U19105 (N_19105,N_11526,N_13901);
nand U19106 (N_19106,N_13789,N_11748);
and U19107 (N_19107,N_14483,N_12213);
nor U19108 (N_19108,N_10840,N_13530);
nand U19109 (N_19109,N_10803,N_11661);
nor U19110 (N_19110,N_10898,N_10538);
nand U19111 (N_19111,N_14103,N_13008);
nand U19112 (N_19112,N_14291,N_14693);
nor U19113 (N_19113,N_12189,N_13208);
nand U19114 (N_19114,N_12227,N_13175);
nor U19115 (N_19115,N_10414,N_13932);
or U19116 (N_19116,N_14563,N_13620);
or U19117 (N_19117,N_14147,N_14488);
nor U19118 (N_19118,N_14142,N_14862);
nor U19119 (N_19119,N_12225,N_13149);
nor U19120 (N_19120,N_14864,N_12919);
and U19121 (N_19121,N_13996,N_10398);
nor U19122 (N_19122,N_11184,N_12382);
nor U19123 (N_19123,N_11443,N_13125);
and U19124 (N_19124,N_12473,N_12071);
and U19125 (N_19125,N_10939,N_14834);
nand U19126 (N_19126,N_13042,N_14102);
nor U19127 (N_19127,N_14141,N_13063);
nand U19128 (N_19128,N_13620,N_10106);
and U19129 (N_19129,N_12175,N_12159);
nor U19130 (N_19130,N_12985,N_13312);
nor U19131 (N_19131,N_11560,N_11864);
nor U19132 (N_19132,N_12453,N_12142);
and U19133 (N_19133,N_13731,N_14690);
nand U19134 (N_19134,N_12218,N_10643);
nand U19135 (N_19135,N_13033,N_12914);
and U19136 (N_19136,N_11220,N_13286);
nand U19137 (N_19137,N_10151,N_13948);
nor U19138 (N_19138,N_11344,N_10135);
or U19139 (N_19139,N_14832,N_12882);
or U19140 (N_19140,N_12907,N_10261);
and U19141 (N_19141,N_13253,N_11052);
or U19142 (N_19142,N_13155,N_13446);
nor U19143 (N_19143,N_12434,N_10978);
nor U19144 (N_19144,N_11831,N_10465);
nor U19145 (N_19145,N_11189,N_13832);
or U19146 (N_19146,N_13522,N_14095);
nor U19147 (N_19147,N_13931,N_10194);
nor U19148 (N_19148,N_13164,N_10924);
or U19149 (N_19149,N_13439,N_10865);
and U19150 (N_19150,N_10689,N_13476);
or U19151 (N_19151,N_11431,N_11853);
or U19152 (N_19152,N_13244,N_10575);
nand U19153 (N_19153,N_10803,N_13729);
or U19154 (N_19154,N_14840,N_13986);
or U19155 (N_19155,N_11071,N_14866);
and U19156 (N_19156,N_11130,N_13319);
nand U19157 (N_19157,N_12679,N_12200);
and U19158 (N_19158,N_12453,N_11108);
or U19159 (N_19159,N_14202,N_13314);
or U19160 (N_19160,N_13202,N_12500);
and U19161 (N_19161,N_10284,N_11828);
or U19162 (N_19162,N_12371,N_14610);
or U19163 (N_19163,N_13687,N_13686);
and U19164 (N_19164,N_10713,N_14954);
nor U19165 (N_19165,N_14781,N_14621);
and U19166 (N_19166,N_10779,N_13606);
nor U19167 (N_19167,N_12601,N_14380);
nand U19168 (N_19168,N_11377,N_11232);
and U19169 (N_19169,N_10525,N_13269);
and U19170 (N_19170,N_14018,N_11789);
nand U19171 (N_19171,N_12820,N_11331);
or U19172 (N_19172,N_11149,N_11114);
and U19173 (N_19173,N_11333,N_10831);
and U19174 (N_19174,N_10056,N_11259);
nand U19175 (N_19175,N_11785,N_13154);
or U19176 (N_19176,N_11553,N_11928);
or U19177 (N_19177,N_10639,N_11242);
and U19178 (N_19178,N_11548,N_13078);
nand U19179 (N_19179,N_13594,N_10748);
or U19180 (N_19180,N_14871,N_12459);
nand U19181 (N_19181,N_12327,N_12497);
and U19182 (N_19182,N_11613,N_12010);
nor U19183 (N_19183,N_10856,N_14055);
nand U19184 (N_19184,N_14126,N_13428);
or U19185 (N_19185,N_13388,N_11694);
nand U19186 (N_19186,N_11930,N_10759);
nor U19187 (N_19187,N_14220,N_10700);
and U19188 (N_19188,N_10888,N_12316);
nand U19189 (N_19189,N_10164,N_13674);
nor U19190 (N_19190,N_14998,N_13495);
nand U19191 (N_19191,N_12001,N_10517);
or U19192 (N_19192,N_10465,N_12009);
or U19193 (N_19193,N_14678,N_11460);
nor U19194 (N_19194,N_12534,N_11763);
and U19195 (N_19195,N_10992,N_13440);
nor U19196 (N_19196,N_12136,N_11231);
and U19197 (N_19197,N_12955,N_12303);
nor U19198 (N_19198,N_10887,N_14862);
and U19199 (N_19199,N_11527,N_13968);
or U19200 (N_19200,N_14647,N_14662);
nand U19201 (N_19201,N_12957,N_10154);
or U19202 (N_19202,N_14928,N_11041);
nand U19203 (N_19203,N_12057,N_14726);
xnor U19204 (N_19204,N_11696,N_11274);
nor U19205 (N_19205,N_13453,N_13729);
nor U19206 (N_19206,N_14818,N_13838);
xnor U19207 (N_19207,N_10149,N_13747);
nor U19208 (N_19208,N_14733,N_13387);
nor U19209 (N_19209,N_11418,N_11593);
and U19210 (N_19210,N_13204,N_11625);
nand U19211 (N_19211,N_12739,N_12453);
nand U19212 (N_19212,N_12042,N_14482);
or U19213 (N_19213,N_10276,N_14171);
nand U19214 (N_19214,N_14507,N_11070);
nor U19215 (N_19215,N_13743,N_12086);
nand U19216 (N_19216,N_11416,N_12477);
nor U19217 (N_19217,N_13011,N_11013);
nor U19218 (N_19218,N_12818,N_11474);
nor U19219 (N_19219,N_10276,N_10749);
nor U19220 (N_19220,N_11846,N_14514);
or U19221 (N_19221,N_13267,N_12831);
nor U19222 (N_19222,N_11247,N_14350);
and U19223 (N_19223,N_12977,N_11164);
or U19224 (N_19224,N_11083,N_13927);
nor U19225 (N_19225,N_13874,N_14231);
and U19226 (N_19226,N_12488,N_14722);
and U19227 (N_19227,N_10001,N_13345);
and U19228 (N_19228,N_13089,N_14801);
nand U19229 (N_19229,N_11120,N_14063);
or U19230 (N_19230,N_12719,N_14792);
nor U19231 (N_19231,N_10725,N_14763);
or U19232 (N_19232,N_14803,N_11719);
nand U19233 (N_19233,N_10066,N_12556);
nor U19234 (N_19234,N_10258,N_14088);
nor U19235 (N_19235,N_13007,N_12724);
nand U19236 (N_19236,N_11257,N_13373);
xnor U19237 (N_19237,N_10929,N_14331);
or U19238 (N_19238,N_14301,N_10879);
nand U19239 (N_19239,N_14916,N_13767);
or U19240 (N_19240,N_10873,N_10956);
and U19241 (N_19241,N_14125,N_14758);
or U19242 (N_19242,N_14790,N_14119);
nor U19243 (N_19243,N_10807,N_11634);
nand U19244 (N_19244,N_13092,N_10183);
or U19245 (N_19245,N_14183,N_13733);
and U19246 (N_19246,N_10699,N_12312);
nand U19247 (N_19247,N_10247,N_13511);
nor U19248 (N_19248,N_11175,N_13748);
xor U19249 (N_19249,N_13881,N_10789);
nand U19250 (N_19250,N_10626,N_11535);
and U19251 (N_19251,N_11935,N_14065);
or U19252 (N_19252,N_10248,N_14970);
and U19253 (N_19253,N_13015,N_11522);
and U19254 (N_19254,N_12387,N_14965);
or U19255 (N_19255,N_14546,N_14085);
and U19256 (N_19256,N_10723,N_12834);
or U19257 (N_19257,N_13132,N_12667);
nand U19258 (N_19258,N_11220,N_14942);
nand U19259 (N_19259,N_13216,N_14070);
or U19260 (N_19260,N_14936,N_11566);
and U19261 (N_19261,N_13520,N_14890);
and U19262 (N_19262,N_13555,N_14289);
and U19263 (N_19263,N_12551,N_14513);
nor U19264 (N_19264,N_12447,N_14052);
nand U19265 (N_19265,N_10973,N_10892);
and U19266 (N_19266,N_13244,N_13643);
nand U19267 (N_19267,N_12874,N_13953);
and U19268 (N_19268,N_12263,N_11223);
and U19269 (N_19269,N_14357,N_12391);
and U19270 (N_19270,N_11879,N_14321);
and U19271 (N_19271,N_10148,N_11118);
nor U19272 (N_19272,N_10173,N_14521);
and U19273 (N_19273,N_11747,N_12939);
nor U19274 (N_19274,N_12940,N_12872);
or U19275 (N_19275,N_10358,N_13364);
or U19276 (N_19276,N_10425,N_13770);
or U19277 (N_19277,N_14832,N_14977);
nor U19278 (N_19278,N_13370,N_10088);
and U19279 (N_19279,N_11302,N_11867);
nand U19280 (N_19280,N_11913,N_11093);
or U19281 (N_19281,N_14593,N_12295);
and U19282 (N_19282,N_10522,N_11649);
nand U19283 (N_19283,N_14741,N_11056);
or U19284 (N_19284,N_13844,N_14578);
nand U19285 (N_19285,N_14516,N_10911);
nand U19286 (N_19286,N_10308,N_12643);
and U19287 (N_19287,N_14217,N_10113);
and U19288 (N_19288,N_13221,N_11612);
nor U19289 (N_19289,N_14862,N_11998);
or U19290 (N_19290,N_14196,N_14168);
nand U19291 (N_19291,N_11448,N_11997);
nor U19292 (N_19292,N_12301,N_11672);
or U19293 (N_19293,N_13877,N_12983);
nand U19294 (N_19294,N_14766,N_10818);
nor U19295 (N_19295,N_13664,N_13110);
or U19296 (N_19296,N_12605,N_11746);
and U19297 (N_19297,N_14020,N_13511);
and U19298 (N_19298,N_10946,N_11161);
xor U19299 (N_19299,N_10804,N_13129);
nor U19300 (N_19300,N_14410,N_13506);
and U19301 (N_19301,N_12575,N_13613);
nand U19302 (N_19302,N_13286,N_14184);
nand U19303 (N_19303,N_13254,N_10402);
nor U19304 (N_19304,N_10279,N_14204);
nand U19305 (N_19305,N_12841,N_13426);
or U19306 (N_19306,N_10282,N_14566);
and U19307 (N_19307,N_14230,N_11800);
or U19308 (N_19308,N_12374,N_12130);
nand U19309 (N_19309,N_13307,N_10428);
nand U19310 (N_19310,N_13273,N_11244);
nand U19311 (N_19311,N_11787,N_10316);
and U19312 (N_19312,N_11386,N_11679);
nand U19313 (N_19313,N_10829,N_10799);
or U19314 (N_19314,N_10942,N_12040);
or U19315 (N_19315,N_10807,N_12213);
nor U19316 (N_19316,N_11346,N_12427);
and U19317 (N_19317,N_10852,N_10801);
or U19318 (N_19318,N_12550,N_12344);
and U19319 (N_19319,N_13232,N_11567);
nand U19320 (N_19320,N_13720,N_12546);
and U19321 (N_19321,N_14907,N_11586);
nor U19322 (N_19322,N_12170,N_11003);
or U19323 (N_19323,N_11276,N_14891);
and U19324 (N_19324,N_13345,N_10027);
or U19325 (N_19325,N_13701,N_10593);
or U19326 (N_19326,N_14529,N_12121);
or U19327 (N_19327,N_12197,N_12023);
or U19328 (N_19328,N_10260,N_10097);
xor U19329 (N_19329,N_13499,N_13724);
and U19330 (N_19330,N_14943,N_10399);
and U19331 (N_19331,N_11893,N_10001);
nand U19332 (N_19332,N_10061,N_11264);
nor U19333 (N_19333,N_14180,N_14396);
or U19334 (N_19334,N_11474,N_12744);
nor U19335 (N_19335,N_14039,N_10761);
or U19336 (N_19336,N_12101,N_11355);
and U19337 (N_19337,N_13819,N_12775);
xor U19338 (N_19338,N_14538,N_11511);
nand U19339 (N_19339,N_10458,N_13802);
or U19340 (N_19340,N_14038,N_13353);
nand U19341 (N_19341,N_13775,N_12500);
or U19342 (N_19342,N_14214,N_12298);
or U19343 (N_19343,N_14258,N_14448);
and U19344 (N_19344,N_10689,N_11682);
or U19345 (N_19345,N_12973,N_12102);
or U19346 (N_19346,N_11830,N_12743);
nand U19347 (N_19347,N_13174,N_14570);
nor U19348 (N_19348,N_10109,N_10697);
or U19349 (N_19349,N_12853,N_12759);
nor U19350 (N_19350,N_13214,N_14985);
nand U19351 (N_19351,N_13296,N_12316);
nand U19352 (N_19352,N_12325,N_10322);
nand U19353 (N_19353,N_10633,N_12958);
or U19354 (N_19354,N_12663,N_10912);
nand U19355 (N_19355,N_12258,N_10540);
xor U19356 (N_19356,N_13913,N_11564);
nor U19357 (N_19357,N_11346,N_12286);
and U19358 (N_19358,N_10708,N_11694);
nor U19359 (N_19359,N_12655,N_10698);
nor U19360 (N_19360,N_13162,N_10068);
or U19361 (N_19361,N_13461,N_10588);
and U19362 (N_19362,N_11751,N_14053);
nand U19363 (N_19363,N_12299,N_10705);
nand U19364 (N_19364,N_11915,N_10488);
nor U19365 (N_19365,N_11782,N_14254);
or U19366 (N_19366,N_14314,N_10346);
xor U19367 (N_19367,N_10334,N_13748);
nand U19368 (N_19368,N_11783,N_13857);
and U19369 (N_19369,N_14283,N_13041);
and U19370 (N_19370,N_13286,N_11758);
nor U19371 (N_19371,N_10604,N_12567);
nor U19372 (N_19372,N_14029,N_11879);
nor U19373 (N_19373,N_13682,N_11624);
and U19374 (N_19374,N_12927,N_11869);
and U19375 (N_19375,N_14206,N_12841);
nor U19376 (N_19376,N_12500,N_14945);
nor U19377 (N_19377,N_14725,N_10604);
nand U19378 (N_19378,N_12222,N_14876);
and U19379 (N_19379,N_11877,N_11081);
xnor U19380 (N_19380,N_14693,N_12587);
and U19381 (N_19381,N_11309,N_14256);
xnor U19382 (N_19382,N_13659,N_10967);
nand U19383 (N_19383,N_10601,N_12416);
or U19384 (N_19384,N_14125,N_11439);
or U19385 (N_19385,N_11982,N_13283);
nand U19386 (N_19386,N_11433,N_14475);
nor U19387 (N_19387,N_11338,N_10266);
nand U19388 (N_19388,N_12777,N_10928);
or U19389 (N_19389,N_13499,N_11036);
and U19390 (N_19390,N_14786,N_14674);
and U19391 (N_19391,N_12226,N_12724);
and U19392 (N_19392,N_12466,N_14931);
or U19393 (N_19393,N_10712,N_10767);
nand U19394 (N_19394,N_10718,N_10152);
nor U19395 (N_19395,N_10595,N_12975);
xnor U19396 (N_19396,N_13034,N_12161);
nand U19397 (N_19397,N_11445,N_12662);
and U19398 (N_19398,N_11428,N_13259);
nor U19399 (N_19399,N_14681,N_14609);
nand U19400 (N_19400,N_13250,N_14558);
nor U19401 (N_19401,N_12159,N_10521);
and U19402 (N_19402,N_10135,N_12606);
or U19403 (N_19403,N_13813,N_13891);
or U19404 (N_19404,N_13735,N_11666);
nand U19405 (N_19405,N_14011,N_11555);
and U19406 (N_19406,N_14525,N_10481);
nor U19407 (N_19407,N_10530,N_11809);
and U19408 (N_19408,N_11432,N_14580);
or U19409 (N_19409,N_10950,N_10138);
nand U19410 (N_19410,N_12522,N_13277);
nor U19411 (N_19411,N_14439,N_14751);
nor U19412 (N_19412,N_14774,N_12158);
or U19413 (N_19413,N_14915,N_11042);
xnor U19414 (N_19414,N_14255,N_14597);
xnor U19415 (N_19415,N_12798,N_14195);
nor U19416 (N_19416,N_10562,N_12300);
and U19417 (N_19417,N_14172,N_11015);
and U19418 (N_19418,N_13940,N_11585);
or U19419 (N_19419,N_14042,N_11816);
and U19420 (N_19420,N_12719,N_10018);
nand U19421 (N_19421,N_11739,N_11880);
nand U19422 (N_19422,N_14366,N_11273);
nand U19423 (N_19423,N_13919,N_11857);
or U19424 (N_19424,N_14656,N_10022);
and U19425 (N_19425,N_11557,N_13632);
and U19426 (N_19426,N_14513,N_14420);
and U19427 (N_19427,N_12920,N_12965);
nor U19428 (N_19428,N_12667,N_10684);
or U19429 (N_19429,N_12139,N_10396);
and U19430 (N_19430,N_10459,N_13167);
nor U19431 (N_19431,N_10856,N_13868);
nor U19432 (N_19432,N_12178,N_12710);
nand U19433 (N_19433,N_13806,N_14994);
nand U19434 (N_19434,N_10183,N_13542);
and U19435 (N_19435,N_11591,N_14993);
nand U19436 (N_19436,N_12973,N_11234);
nand U19437 (N_19437,N_14712,N_13694);
or U19438 (N_19438,N_11563,N_13667);
nor U19439 (N_19439,N_11995,N_12027);
or U19440 (N_19440,N_14495,N_14511);
or U19441 (N_19441,N_11348,N_11591);
or U19442 (N_19442,N_10693,N_14486);
and U19443 (N_19443,N_13276,N_12744);
nand U19444 (N_19444,N_11782,N_12506);
nor U19445 (N_19445,N_13399,N_13244);
nand U19446 (N_19446,N_13887,N_13714);
nand U19447 (N_19447,N_14442,N_14804);
and U19448 (N_19448,N_10762,N_10420);
nor U19449 (N_19449,N_13813,N_10352);
or U19450 (N_19450,N_12499,N_10684);
or U19451 (N_19451,N_11668,N_13363);
xnor U19452 (N_19452,N_14391,N_14052);
nand U19453 (N_19453,N_12208,N_10705);
xor U19454 (N_19454,N_14754,N_10404);
or U19455 (N_19455,N_14673,N_12832);
nor U19456 (N_19456,N_13617,N_11835);
and U19457 (N_19457,N_14896,N_13206);
or U19458 (N_19458,N_10459,N_11188);
nand U19459 (N_19459,N_10303,N_10780);
nor U19460 (N_19460,N_11824,N_14791);
nand U19461 (N_19461,N_11575,N_14749);
nor U19462 (N_19462,N_10061,N_10923);
nand U19463 (N_19463,N_13835,N_11272);
nand U19464 (N_19464,N_13799,N_10640);
or U19465 (N_19465,N_13690,N_14838);
and U19466 (N_19466,N_10341,N_13557);
nor U19467 (N_19467,N_13405,N_13793);
and U19468 (N_19468,N_14941,N_12302);
and U19469 (N_19469,N_13049,N_13778);
nor U19470 (N_19470,N_13612,N_11225);
nor U19471 (N_19471,N_10149,N_11877);
and U19472 (N_19472,N_11589,N_10921);
nor U19473 (N_19473,N_14705,N_13342);
and U19474 (N_19474,N_14231,N_12790);
nand U19475 (N_19475,N_14436,N_12627);
or U19476 (N_19476,N_12226,N_13736);
nand U19477 (N_19477,N_11425,N_14581);
and U19478 (N_19478,N_14790,N_14144);
nor U19479 (N_19479,N_14459,N_10220);
nand U19480 (N_19480,N_13516,N_10920);
and U19481 (N_19481,N_14837,N_14190);
nand U19482 (N_19482,N_14971,N_11674);
nand U19483 (N_19483,N_11988,N_14987);
and U19484 (N_19484,N_13668,N_14452);
xor U19485 (N_19485,N_11392,N_10355);
and U19486 (N_19486,N_10104,N_12730);
nand U19487 (N_19487,N_13586,N_10625);
or U19488 (N_19488,N_11482,N_10592);
or U19489 (N_19489,N_11242,N_12728);
or U19490 (N_19490,N_12794,N_11742);
nand U19491 (N_19491,N_10856,N_12570);
nand U19492 (N_19492,N_11884,N_10268);
nor U19493 (N_19493,N_11031,N_11834);
nand U19494 (N_19494,N_14223,N_13989);
or U19495 (N_19495,N_13656,N_13122);
xnor U19496 (N_19496,N_13033,N_14083);
nand U19497 (N_19497,N_10102,N_12355);
and U19498 (N_19498,N_10070,N_13289);
xnor U19499 (N_19499,N_14166,N_13668);
nor U19500 (N_19500,N_14216,N_10369);
and U19501 (N_19501,N_10197,N_12819);
nor U19502 (N_19502,N_12726,N_10013);
or U19503 (N_19503,N_12499,N_13267);
nand U19504 (N_19504,N_12969,N_14232);
nor U19505 (N_19505,N_11158,N_14083);
nor U19506 (N_19506,N_10885,N_10453);
nor U19507 (N_19507,N_11634,N_13139);
or U19508 (N_19508,N_11221,N_13603);
or U19509 (N_19509,N_14713,N_13190);
or U19510 (N_19510,N_11845,N_10104);
or U19511 (N_19511,N_12789,N_13993);
nand U19512 (N_19512,N_11531,N_12783);
and U19513 (N_19513,N_11000,N_14905);
nor U19514 (N_19514,N_10229,N_11976);
nor U19515 (N_19515,N_14856,N_14640);
nand U19516 (N_19516,N_12831,N_11299);
nor U19517 (N_19517,N_12614,N_12542);
or U19518 (N_19518,N_13234,N_14108);
or U19519 (N_19519,N_10846,N_13656);
and U19520 (N_19520,N_10958,N_11044);
nor U19521 (N_19521,N_11099,N_11693);
or U19522 (N_19522,N_10773,N_14899);
nor U19523 (N_19523,N_12487,N_12387);
or U19524 (N_19524,N_12063,N_13875);
or U19525 (N_19525,N_13750,N_10646);
or U19526 (N_19526,N_10282,N_11913);
or U19527 (N_19527,N_14758,N_13503);
nor U19528 (N_19528,N_13415,N_14787);
nor U19529 (N_19529,N_11407,N_12986);
nand U19530 (N_19530,N_13245,N_12819);
nor U19531 (N_19531,N_10533,N_12032);
or U19532 (N_19532,N_14379,N_12727);
and U19533 (N_19533,N_12424,N_11148);
or U19534 (N_19534,N_10966,N_11865);
or U19535 (N_19535,N_11511,N_11223);
or U19536 (N_19536,N_10114,N_11738);
xnor U19537 (N_19537,N_10394,N_13680);
or U19538 (N_19538,N_14169,N_11825);
nor U19539 (N_19539,N_12961,N_11063);
xnor U19540 (N_19540,N_10417,N_13473);
nor U19541 (N_19541,N_13032,N_11376);
or U19542 (N_19542,N_12105,N_12229);
nor U19543 (N_19543,N_11592,N_10486);
nand U19544 (N_19544,N_14018,N_11042);
or U19545 (N_19545,N_11874,N_14634);
nor U19546 (N_19546,N_12473,N_10642);
or U19547 (N_19547,N_14669,N_10087);
or U19548 (N_19548,N_14313,N_12841);
nand U19549 (N_19549,N_11831,N_14729);
or U19550 (N_19550,N_13766,N_11691);
and U19551 (N_19551,N_14019,N_12759);
nand U19552 (N_19552,N_14928,N_10275);
and U19553 (N_19553,N_11249,N_10305);
and U19554 (N_19554,N_12322,N_10483);
nand U19555 (N_19555,N_13930,N_12758);
or U19556 (N_19556,N_12919,N_13466);
and U19557 (N_19557,N_12748,N_12262);
or U19558 (N_19558,N_10660,N_11908);
or U19559 (N_19559,N_14075,N_14481);
nand U19560 (N_19560,N_12063,N_13898);
and U19561 (N_19561,N_13450,N_11969);
or U19562 (N_19562,N_11272,N_13951);
nor U19563 (N_19563,N_10349,N_10632);
nor U19564 (N_19564,N_11475,N_12598);
nor U19565 (N_19565,N_10172,N_11685);
nor U19566 (N_19566,N_14167,N_12620);
nand U19567 (N_19567,N_10501,N_13266);
or U19568 (N_19568,N_11416,N_11503);
nor U19569 (N_19569,N_12052,N_14732);
or U19570 (N_19570,N_10455,N_12136);
or U19571 (N_19571,N_12797,N_13997);
nor U19572 (N_19572,N_10345,N_11747);
or U19573 (N_19573,N_14824,N_11394);
or U19574 (N_19574,N_14486,N_13671);
and U19575 (N_19575,N_14764,N_13258);
nor U19576 (N_19576,N_14275,N_10793);
nand U19577 (N_19577,N_10395,N_11843);
and U19578 (N_19578,N_12673,N_10124);
and U19579 (N_19579,N_12031,N_10667);
and U19580 (N_19580,N_11844,N_13106);
or U19581 (N_19581,N_12305,N_11380);
or U19582 (N_19582,N_10199,N_13055);
nand U19583 (N_19583,N_14452,N_14628);
nor U19584 (N_19584,N_11149,N_12812);
nand U19585 (N_19585,N_13054,N_14649);
nand U19586 (N_19586,N_10888,N_13009);
or U19587 (N_19587,N_13205,N_13263);
or U19588 (N_19588,N_10808,N_11069);
nand U19589 (N_19589,N_11695,N_13822);
or U19590 (N_19590,N_14030,N_10277);
nand U19591 (N_19591,N_14512,N_10586);
nor U19592 (N_19592,N_11956,N_12591);
or U19593 (N_19593,N_12640,N_11336);
nor U19594 (N_19594,N_13354,N_12773);
or U19595 (N_19595,N_10199,N_12972);
xor U19596 (N_19596,N_12684,N_11676);
xor U19597 (N_19597,N_12727,N_13348);
nor U19598 (N_19598,N_14617,N_14242);
and U19599 (N_19599,N_11664,N_13445);
nand U19600 (N_19600,N_10685,N_10342);
or U19601 (N_19601,N_13170,N_14156);
nand U19602 (N_19602,N_13177,N_10182);
nor U19603 (N_19603,N_14624,N_10147);
and U19604 (N_19604,N_11279,N_14406);
or U19605 (N_19605,N_14983,N_10099);
nand U19606 (N_19606,N_12735,N_11754);
nand U19607 (N_19607,N_11041,N_12600);
nand U19608 (N_19608,N_11128,N_10836);
and U19609 (N_19609,N_10638,N_13431);
nor U19610 (N_19610,N_11766,N_14634);
and U19611 (N_19611,N_14546,N_13295);
nor U19612 (N_19612,N_14753,N_13761);
nor U19613 (N_19613,N_14393,N_14854);
nand U19614 (N_19614,N_11417,N_13305);
and U19615 (N_19615,N_14888,N_11960);
nand U19616 (N_19616,N_12152,N_14175);
nor U19617 (N_19617,N_11340,N_12097);
or U19618 (N_19618,N_11440,N_12975);
nand U19619 (N_19619,N_10838,N_12333);
nor U19620 (N_19620,N_12098,N_12108);
nand U19621 (N_19621,N_14137,N_10430);
nand U19622 (N_19622,N_13601,N_12218);
and U19623 (N_19623,N_12373,N_13102);
and U19624 (N_19624,N_12616,N_11514);
nand U19625 (N_19625,N_10112,N_14863);
and U19626 (N_19626,N_12113,N_11399);
and U19627 (N_19627,N_10267,N_12234);
nor U19628 (N_19628,N_11623,N_12794);
nand U19629 (N_19629,N_12696,N_12235);
nor U19630 (N_19630,N_11293,N_12414);
nand U19631 (N_19631,N_11362,N_13792);
nand U19632 (N_19632,N_11349,N_13713);
and U19633 (N_19633,N_12649,N_11955);
nor U19634 (N_19634,N_12524,N_10065);
xnor U19635 (N_19635,N_12550,N_14978);
and U19636 (N_19636,N_14768,N_14956);
nand U19637 (N_19637,N_14321,N_13127);
nor U19638 (N_19638,N_12420,N_14167);
nand U19639 (N_19639,N_10807,N_13514);
and U19640 (N_19640,N_12226,N_13374);
or U19641 (N_19641,N_10264,N_11315);
nor U19642 (N_19642,N_12213,N_14327);
and U19643 (N_19643,N_13758,N_11188);
and U19644 (N_19644,N_13693,N_14293);
or U19645 (N_19645,N_14373,N_14186);
nor U19646 (N_19646,N_12611,N_10651);
or U19647 (N_19647,N_10558,N_11549);
nand U19648 (N_19648,N_10011,N_12247);
and U19649 (N_19649,N_14510,N_13165);
nand U19650 (N_19650,N_14912,N_14606);
or U19651 (N_19651,N_14717,N_14590);
nor U19652 (N_19652,N_10445,N_12936);
and U19653 (N_19653,N_12904,N_14312);
and U19654 (N_19654,N_10921,N_14270);
and U19655 (N_19655,N_12517,N_14000);
and U19656 (N_19656,N_11353,N_14667);
nor U19657 (N_19657,N_12162,N_13215);
nor U19658 (N_19658,N_13814,N_12148);
nor U19659 (N_19659,N_12244,N_11548);
and U19660 (N_19660,N_12267,N_12692);
xnor U19661 (N_19661,N_11393,N_10385);
nor U19662 (N_19662,N_13100,N_13499);
or U19663 (N_19663,N_12156,N_13160);
and U19664 (N_19664,N_13925,N_12828);
nor U19665 (N_19665,N_12516,N_13174);
and U19666 (N_19666,N_12909,N_12602);
nor U19667 (N_19667,N_10201,N_13877);
and U19668 (N_19668,N_12469,N_12256);
xnor U19669 (N_19669,N_14730,N_13782);
or U19670 (N_19670,N_12189,N_14909);
or U19671 (N_19671,N_13605,N_10193);
nand U19672 (N_19672,N_10953,N_11881);
nand U19673 (N_19673,N_10606,N_13382);
nand U19674 (N_19674,N_10045,N_11608);
nand U19675 (N_19675,N_10979,N_11029);
and U19676 (N_19676,N_14140,N_12217);
nand U19677 (N_19677,N_14008,N_11074);
or U19678 (N_19678,N_12332,N_10538);
and U19679 (N_19679,N_14896,N_14578);
and U19680 (N_19680,N_14335,N_10111);
and U19681 (N_19681,N_10558,N_12970);
nand U19682 (N_19682,N_10070,N_13513);
or U19683 (N_19683,N_13633,N_13318);
nor U19684 (N_19684,N_11784,N_10782);
nand U19685 (N_19685,N_14039,N_14642);
nand U19686 (N_19686,N_10556,N_14277);
and U19687 (N_19687,N_12844,N_14991);
and U19688 (N_19688,N_10314,N_11868);
xnor U19689 (N_19689,N_14750,N_14692);
nor U19690 (N_19690,N_10754,N_11200);
nor U19691 (N_19691,N_14597,N_13780);
or U19692 (N_19692,N_10987,N_12439);
nor U19693 (N_19693,N_13545,N_11871);
xor U19694 (N_19694,N_12476,N_14345);
and U19695 (N_19695,N_12596,N_11415);
nor U19696 (N_19696,N_11495,N_12117);
nand U19697 (N_19697,N_12359,N_14456);
and U19698 (N_19698,N_12379,N_14920);
nor U19699 (N_19699,N_10293,N_12390);
xor U19700 (N_19700,N_12707,N_14602);
and U19701 (N_19701,N_13801,N_14262);
xnor U19702 (N_19702,N_10275,N_10172);
nand U19703 (N_19703,N_10754,N_11211);
or U19704 (N_19704,N_13728,N_10264);
nor U19705 (N_19705,N_13782,N_14248);
nor U19706 (N_19706,N_14111,N_13855);
nor U19707 (N_19707,N_14148,N_13744);
nand U19708 (N_19708,N_14540,N_12820);
nor U19709 (N_19709,N_13268,N_13505);
nand U19710 (N_19710,N_11237,N_14220);
nor U19711 (N_19711,N_11606,N_13547);
nor U19712 (N_19712,N_14728,N_13337);
and U19713 (N_19713,N_14847,N_14515);
or U19714 (N_19714,N_10728,N_12768);
nor U19715 (N_19715,N_12860,N_11950);
nand U19716 (N_19716,N_10595,N_12589);
nand U19717 (N_19717,N_14651,N_13709);
nor U19718 (N_19718,N_14926,N_10163);
and U19719 (N_19719,N_13667,N_12965);
and U19720 (N_19720,N_11003,N_10772);
or U19721 (N_19721,N_10362,N_11128);
and U19722 (N_19722,N_10858,N_14047);
nor U19723 (N_19723,N_10511,N_13644);
nand U19724 (N_19724,N_12420,N_13843);
or U19725 (N_19725,N_14546,N_11639);
nand U19726 (N_19726,N_12079,N_11044);
nand U19727 (N_19727,N_11051,N_14659);
nand U19728 (N_19728,N_14032,N_14314);
nor U19729 (N_19729,N_14290,N_13123);
nand U19730 (N_19730,N_14078,N_14947);
nor U19731 (N_19731,N_10150,N_11924);
nand U19732 (N_19732,N_12525,N_13423);
and U19733 (N_19733,N_11721,N_12874);
and U19734 (N_19734,N_13868,N_12267);
nand U19735 (N_19735,N_11355,N_11885);
nor U19736 (N_19736,N_14644,N_10655);
or U19737 (N_19737,N_14956,N_13543);
nor U19738 (N_19738,N_11672,N_11999);
or U19739 (N_19739,N_11220,N_13031);
or U19740 (N_19740,N_13623,N_11947);
and U19741 (N_19741,N_10473,N_11597);
nor U19742 (N_19742,N_14844,N_10364);
and U19743 (N_19743,N_10075,N_14803);
and U19744 (N_19744,N_13279,N_10000);
nor U19745 (N_19745,N_14953,N_14769);
and U19746 (N_19746,N_12672,N_13095);
and U19747 (N_19747,N_12416,N_11412);
and U19748 (N_19748,N_14099,N_12830);
nor U19749 (N_19749,N_12681,N_10049);
and U19750 (N_19750,N_10984,N_11379);
nor U19751 (N_19751,N_14525,N_10971);
nand U19752 (N_19752,N_11725,N_10305);
nor U19753 (N_19753,N_13255,N_13993);
and U19754 (N_19754,N_12382,N_13333);
or U19755 (N_19755,N_13057,N_12008);
and U19756 (N_19756,N_12231,N_10280);
nor U19757 (N_19757,N_10741,N_10619);
nand U19758 (N_19758,N_11135,N_10209);
or U19759 (N_19759,N_12120,N_13000);
or U19760 (N_19760,N_14031,N_10440);
nor U19761 (N_19761,N_11401,N_12961);
or U19762 (N_19762,N_14177,N_12693);
and U19763 (N_19763,N_13757,N_12610);
nor U19764 (N_19764,N_14760,N_11103);
nand U19765 (N_19765,N_10093,N_13595);
nor U19766 (N_19766,N_14154,N_13321);
and U19767 (N_19767,N_13129,N_13810);
or U19768 (N_19768,N_12262,N_14085);
and U19769 (N_19769,N_10978,N_13670);
or U19770 (N_19770,N_11191,N_14438);
nor U19771 (N_19771,N_12521,N_11859);
nand U19772 (N_19772,N_13388,N_14731);
nand U19773 (N_19773,N_11714,N_10135);
and U19774 (N_19774,N_14847,N_12124);
or U19775 (N_19775,N_13110,N_11114);
nand U19776 (N_19776,N_14457,N_14919);
nor U19777 (N_19777,N_11383,N_14314);
and U19778 (N_19778,N_11782,N_11609);
and U19779 (N_19779,N_13060,N_10142);
or U19780 (N_19780,N_11884,N_14127);
nand U19781 (N_19781,N_11772,N_12088);
or U19782 (N_19782,N_12422,N_11691);
nand U19783 (N_19783,N_11102,N_10956);
or U19784 (N_19784,N_12163,N_10252);
or U19785 (N_19785,N_10339,N_11560);
nor U19786 (N_19786,N_12148,N_14894);
nor U19787 (N_19787,N_14595,N_12478);
xnor U19788 (N_19788,N_12029,N_14645);
nand U19789 (N_19789,N_10742,N_14327);
and U19790 (N_19790,N_10129,N_13648);
or U19791 (N_19791,N_14735,N_11207);
nor U19792 (N_19792,N_11121,N_14933);
nand U19793 (N_19793,N_12259,N_13615);
and U19794 (N_19794,N_11671,N_14250);
nand U19795 (N_19795,N_14931,N_11387);
nand U19796 (N_19796,N_13786,N_12584);
or U19797 (N_19797,N_10188,N_11522);
and U19798 (N_19798,N_10131,N_11967);
nor U19799 (N_19799,N_10542,N_14283);
nand U19800 (N_19800,N_10556,N_12363);
or U19801 (N_19801,N_13975,N_13118);
and U19802 (N_19802,N_12374,N_12202);
nand U19803 (N_19803,N_12157,N_13262);
nand U19804 (N_19804,N_14405,N_10322);
and U19805 (N_19805,N_14716,N_13321);
nor U19806 (N_19806,N_14544,N_14343);
or U19807 (N_19807,N_13930,N_12803);
and U19808 (N_19808,N_12957,N_10963);
nand U19809 (N_19809,N_13008,N_11791);
nand U19810 (N_19810,N_11876,N_14634);
nand U19811 (N_19811,N_14922,N_12550);
nand U19812 (N_19812,N_11583,N_14474);
and U19813 (N_19813,N_12358,N_13256);
or U19814 (N_19814,N_14709,N_14942);
and U19815 (N_19815,N_12543,N_14603);
nor U19816 (N_19816,N_12954,N_13002);
nor U19817 (N_19817,N_12151,N_10541);
nand U19818 (N_19818,N_14844,N_13562);
and U19819 (N_19819,N_14832,N_12528);
nor U19820 (N_19820,N_11296,N_10813);
or U19821 (N_19821,N_11405,N_13637);
and U19822 (N_19822,N_14223,N_10526);
nand U19823 (N_19823,N_13079,N_10316);
nand U19824 (N_19824,N_11313,N_12913);
or U19825 (N_19825,N_10124,N_13728);
nor U19826 (N_19826,N_11247,N_14358);
nor U19827 (N_19827,N_13925,N_13447);
nor U19828 (N_19828,N_10620,N_10956);
or U19829 (N_19829,N_10037,N_12981);
or U19830 (N_19830,N_12931,N_10250);
nand U19831 (N_19831,N_12805,N_14699);
nor U19832 (N_19832,N_14962,N_14423);
nor U19833 (N_19833,N_11680,N_14108);
xnor U19834 (N_19834,N_10446,N_11109);
nor U19835 (N_19835,N_11793,N_13191);
and U19836 (N_19836,N_14957,N_13012);
nand U19837 (N_19837,N_13370,N_12207);
nand U19838 (N_19838,N_14437,N_10843);
or U19839 (N_19839,N_14570,N_14289);
nor U19840 (N_19840,N_11379,N_10050);
and U19841 (N_19841,N_13908,N_13020);
or U19842 (N_19842,N_11865,N_13680);
and U19843 (N_19843,N_10302,N_12298);
or U19844 (N_19844,N_10152,N_10294);
nand U19845 (N_19845,N_13202,N_13916);
nand U19846 (N_19846,N_10316,N_11702);
nor U19847 (N_19847,N_11251,N_10727);
or U19848 (N_19848,N_13482,N_11230);
or U19849 (N_19849,N_11746,N_12292);
nor U19850 (N_19850,N_14270,N_11925);
and U19851 (N_19851,N_14341,N_14635);
or U19852 (N_19852,N_10969,N_11670);
xnor U19853 (N_19853,N_11574,N_13605);
and U19854 (N_19854,N_11255,N_13111);
nand U19855 (N_19855,N_12932,N_14548);
and U19856 (N_19856,N_11263,N_13594);
nor U19857 (N_19857,N_14966,N_10903);
or U19858 (N_19858,N_10837,N_14012);
and U19859 (N_19859,N_13822,N_10805);
or U19860 (N_19860,N_11759,N_10850);
nand U19861 (N_19861,N_10157,N_10214);
and U19862 (N_19862,N_14573,N_12449);
and U19863 (N_19863,N_12357,N_11545);
and U19864 (N_19864,N_12692,N_10318);
and U19865 (N_19865,N_14483,N_12570);
nand U19866 (N_19866,N_11098,N_10340);
and U19867 (N_19867,N_12059,N_13555);
nand U19868 (N_19868,N_13914,N_11676);
and U19869 (N_19869,N_13547,N_12017);
nand U19870 (N_19870,N_12702,N_11303);
nor U19871 (N_19871,N_12555,N_13404);
nand U19872 (N_19872,N_11328,N_14976);
nand U19873 (N_19873,N_10129,N_12609);
and U19874 (N_19874,N_12976,N_14410);
nor U19875 (N_19875,N_11103,N_12571);
and U19876 (N_19876,N_11521,N_12844);
nor U19877 (N_19877,N_14554,N_13630);
nand U19878 (N_19878,N_10914,N_13918);
and U19879 (N_19879,N_12124,N_14541);
xnor U19880 (N_19880,N_13942,N_14394);
or U19881 (N_19881,N_10993,N_10235);
nand U19882 (N_19882,N_14815,N_12636);
nand U19883 (N_19883,N_10187,N_10208);
or U19884 (N_19884,N_10590,N_12723);
nand U19885 (N_19885,N_14808,N_13943);
and U19886 (N_19886,N_14238,N_11605);
nor U19887 (N_19887,N_13600,N_14465);
or U19888 (N_19888,N_10872,N_10891);
nand U19889 (N_19889,N_12433,N_12058);
nand U19890 (N_19890,N_10313,N_13786);
or U19891 (N_19891,N_12804,N_10200);
nor U19892 (N_19892,N_14077,N_11320);
nor U19893 (N_19893,N_10096,N_14020);
nand U19894 (N_19894,N_12098,N_12863);
and U19895 (N_19895,N_13967,N_12174);
nor U19896 (N_19896,N_12386,N_10572);
nor U19897 (N_19897,N_13442,N_12635);
and U19898 (N_19898,N_13563,N_14435);
xor U19899 (N_19899,N_13714,N_14196);
nand U19900 (N_19900,N_10816,N_14300);
nand U19901 (N_19901,N_10494,N_12002);
and U19902 (N_19902,N_12302,N_14816);
nand U19903 (N_19903,N_11524,N_12158);
nand U19904 (N_19904,N_12645,N_12083);
nand U19905 (N_19905,N_12161,N_13750);
nand U19906 (N_19906,N_13319,N_12865);
nor U19907 (N_19907,N_13246,N_13106);
nand U19908 (N_19908,N_12865,N_14703);
nor U19909 (N_19909,N_12882,N_13479);
nand U19910 (N_19910,N_13209,N_12213);
nor U19911 (N_19911,N_14271,N_12510);
and U19912 (N_19912,N_14156,N_11257);
nand U19913 (N_19913,N_12229,N_11816);
and U19914 (N_19914,N_14253,N_10019);
or U19915 (N_19915,N_13079,N_10787);
or U19916 (N_19916,N_10011,N_10462);
and U19917 (N_19917,N_12962,N_14163);
nor U19918 (N_19918,N_11841,N_10993);
nor U19919 (N_19919,N_10777,N_11219);
and U19920 (N_19920,N_14643,N_12151);
nor U19921 (N_19921,N_10399,N_12325);
and U19922 (N_19922,N_12010,N_13466);
or U19923 (N_19923,N_14648,N_14296);
and U19924 (N_19924,N_11539,N_13707);
nand U19925 (N_19925,N_11985,N_13037);
and U19926 (N_19926,N_14652,N_14212);
and U19927 (N_19927,N_14703,N_14133);
and U19928 (N_19928,N_12323,N_10783);
and U19929 (N_19929,N_14866,N_13897);
nor U19930 (N_19930,N_11672,N_12873);
and U19931 (N_19931,N_12831,N_13634);
and U19932 (N_19932,N_11729,N_11847);
and U19933 (N_19933,N_11780,N_13850);
and U19934 (N_19934,N_10865,N_13752);
or U19935 (N_19935,N_10505,N_13411);
nand U19936 (N_19936,N_14033,N_12427);
and U19937 (N_19937,N_10023,N_11618);
nor U19938 (N_19938,N_10730,N_14041);
nand U19939 (N_19939,N_12468,N_12448);
nand U19940 (N_19940,N_10458,N_14357);
nand U19941 (N_19941,N_14711,N_11013);
nor U19942 (N_19942,N_12529,N_10095);
and U19943 (N_19943,N_12263,N_14767);
and U19944 (N_19944,N_14566,N_13152);
or U19945 (N_19945,N_14412,N_14803);
or U19946 (N_19946,N_12179,N_14579);
and U19947 (N_19947,N_11248,N_14090);
or U19948 (N_19948,N_11417,N_14770);
nor U19949 (N_19949,N_14265,N_13332);
nand U19950 (N_19950,N_14642,N_10002);
nand U19951 (N_19951,N_13551,N_14657);
or U19952 (N_19952,N_10739,N_10427);
or U19953 (N_19953,N_13905,N_12845);
and U19954 (N_19954,N_10324,N_13295);
nor U19955 (N_19955,N_10827,N_13148);
or U19956 (N_19956,N_13037,N_12362);
nand U19957 (N_19957,N_14878,N_12843);
or U19958 (N_19958,N_11778,N_12277);
nor U19959 (N_19959,N_13667,N_12126);
or U19960 (N_19960,N_10601,N_10721);
or U19961 (N_19961,N_13554,N_13971);
nor U19962 (N_19962,N_14361,N_12748);
nor U19963 (N_19963,N_11279,N_13763);
or U19964 (N_19964,N_12397,N_11231);
nor U19965 (N_19965,N_11355,N_10852);
nand U19966 (N_19966,N_11004,N_10253);
or U19967 (N_19967,N_11378,N_12689);
nand U19968 (N_19968,N_11334,N_13926);
nand U19969 (N_19969,N_14192,N_13728);
and U19970 (N_19970,N_14267,N_13930);
nor U19971 (N_19971,N_11445,N_14350);
and U19972 (N_19972,N_13289,N_11066);
nand U19973 (N_19973,N_12229,N_13710);
nor U19974 (N_19974,N_13219,N_10706);
nor U19975 (N_19975,N_13812,N_11802);
or U19976 (N_19976,N_13372,N_11788);
or U19977 (N_19977,N_11205,N_13370);
and U19978 (N_19978,N_10915,N_13922);
nand U19979 (N_19979,N_10267,N_14086);
or U19980 (N_19980,N_13183,N_12873);
xor U19981 (N_19981,N_14354,N_14654);
nand U19982 (N_19982,N_13712,N_10222);
or U19983 (N_19983,N_10752,N_14850);
nand U19984 (N_19984,N_10005,N_13025);
or U19985 (N_19985,N_13016,N_13166);
or U19986 (N_19986,N_10879,N_10502);
nand U19987 (N_19987,N_13521,N_14519);
or U19988 (N_19988,N_13834,N_11571);
nand U19989 (N_19989,N_14548,N_14202);
and U19990 (N_19990,N_10438,N_12371);
nand U19991 (N_19991,N_12019,N_14772);
nor U19992 (N_19992,N_13615,N_10612);
or U19993 (N_19993,N_11411,N_13922);
nand U19994 (N_19994,N_13364,N_11696);
nor U19995 (N_19995,N_14972,N_10007);
nand U19996 (N_19996,N_11958,N_11728);
and U19997 (N_19997,N_11217,N_12339);
and U19998 (N_19998,N_13636,N_10081);
xnor U19999 (N_19999,N_11722,N_13352);
nor UO_0 (O_0,N_15207,N_15247);
or UO_1 (O_1,N_17038,N_18148);
nor UO_2 (O_2,N_15546,N_18631);
nand UO_3 (O_3,N_15887,N_15954);
or UO_4 (O_4,N_17736,N_17768);
xor UO_5 (O_5,N_18888,N_15896);
nor UO_6 (O_6,N_18845,N_19828);
or UO_7 (O_7,N_17695,N_19440);
nand UO_8 (O_8,N_18803,N_16276);
or UO_9 (O_9,N_17881,N_17385);
or UO_10 (O_10,N_17898,N_18167);
or UO_11 (O_11,N_19352,N_17505);
and UO_12 (O_12,N_18059,N_17131);
and UO_13 (O_13,N_19726,N_18010);
nand UO_14 (O_14,N_15504,N_18553);
nor UO_15 (O_15,N_18207,N_15112);
or UO_16 (O_16,N_18800,N_17412);
nand UO_17 (O_17,N_17691,N_16447);
nor UO_18 (O_18,N_18231,N_16397);
nor UO_19 (O_19,N_18530,N_16284);
nand UO_20 (O_20,N_18972,N_15241);
or UO_21 (O_21,N_18725,N_19649);
or UO_22 (O_22,N_18532,N_18844);
xor UO_23 (O_23,N_18158,N_16123);
nor UO_24 (O_24,N_17745,N_17375);
or UO_25 (O_25,N_18661,N_17462);
and UO_26 (O_26,N_19261,N_19326);
or UO_27 (O_27,N_15117,N_17861);
nor UO_28 (O_28,N_18163,N_17342);
and UO_29 (O_29,N_19190,N_17628);
and UO_30 (O_30,N_19107,N_17598);
xor UO_31 (O_31,N_18622,N_19579);
or UO_32 (O_32,N_16705,N_19318);
nand UO_33 (O_33,N_15271,N_17864);
or UO_34 (O_34,N_18193,N_16528);
and UO_35 (O_35,N_16780,N_19841);
nand UO_36 (O_36,N_15399,N_17978);
nor UO_37 (O_37,N_15046,N_17698);
or UO_38 (O_38,N_18420,N_16790);
nor UO_39 (O_39,N_18921,N_17594);
xnor UO_40 (O_40,N_18048,N_17617);
nand UO_41 (O_41,N_15044,N_17220);
nand UO_42 (O_42,N_15171,N_15964);
nand UO_43 (O_43,N_16329,N_16717);
nand UO_44 (O_44,N_19877,N_18541);
nand UO_45 (O_45,N_16738,N_18700);
or UO_46 (O_46,N_16268,N_15377);
nor UO_47 (O_47,N_19565,N_18597);
and UO_48 (O_48,N_19388,N_15909);
nor UO_49 (O_49,N_17688,N_15113);
and UO_50 (O_50,N_18664,N_18166);
nor UO_51 (O_51,N_15227,N_17339);
nand UO_52 (O_52,N_18766,N_16275);
nor UO_53 (O_53,N_18240,N_19934);
and UO_54 (O_54,N_15703,N_18102);
nor UO_55 (O_55,N_18300,N_18284);
or UO_56 (O_56,N_19913,N_16849);
nand UO_57 (O_57,N_16024,N_18660);
nand UO_58 (O_58,N_19720,N_17297);
nor UO_59 (O_59,N_18069,N_19397);
or UO_60 (O_60,N_18692,N_19781);
and UO_61 (O_61,N_17447,N_17895);
or UO_62 (O_62,N_18577,N_18246);
nand UO_63 (O_63,N_15657,N_17459);
nand UO_64 (O_64,N_16159,N_17254);
and UO_65 (O_65,N_15806,N_15834);
nor UO_66 (O_66,N_19818,N_18364);
and UO_67 (O_67,N_16627,N_15622);
nand UO_68 (O_68,N_18268,N_17017);
and UO_69 (O_69,N_17818,N_15977);
xnor UO_70 (O_70,N_15124,N_15865);
nor UO_71 (O_71,N_15267,N_15899);
nor UO_72 (O_72,N_17524,N_17085);
nor UO_73 (O_73,N_19942,N_18647);
and UO_74 (O_74,N_18445,N_18105);
nor UO_75 (O_75,N_19060,N_15201);
and UO_76 (O_76,N_19810,N_19552);
and UO_77 (O_77,N_15232,N_17785);
or UO_78 (O_78,N_15572,N_18269);
nor UO_79 (O_79,N_19027,N_19082);
nand UO_80 (O_80,N_17371,N_15364);
and UO_81 (O_81,N_19186,N_18855);
and UO_82 (O_82,N_18644,N_17416);
nor UO_83 (O_83,N_17904,N_18579);
nor UO_84 (O_84,N_17007,N_15734);
nand UO_85 (O_85,N_19219,N_15177);
and UO_86 (O_86,N_15198,N_18956);
and UO_87 (O_87,N_18161,N_15035);
or UO_88 (O_88,N_19614,N_16917);
or UO_89 (O_89,N_19271,N_17843);
nand UO_90 (O_90,N_16131,N_15666);
or UO_91 (O_91,N_15995,N_15273);
nor UO_92 (O_92,N_16238,N_18683);
or UO_93 (O_93,N_18098,N_15683);
nor UO_94 (O_94,N_16523,N_19036);
nand UO_95 (O_95,N_16454,N_15619);
nand UO_96 (O_96,N_18607,N_18441);
or UO_97 (O_97,N_17384,N_16052);
and UO_98 (O_98,N_15808,N_19247);
xnor UO_99 (O_99,N_17253,N_15006);
and UO_100 (O_100,N_15159,N_19324);
or UO_101 (O_101,N_17854,N_18990);
nor UO_102 (O_102,N_18582,N_15292);
nand UO_103 (O_103,N_18772,N_19092);
and UO_104 (O_104,N_18017,N_15386);
nor UO_105 (O_105,N_19322,N_18241);
or UO_106 (O_106,N_17621,N_19829);
nand UO_107 (O_107,N_17146,N_19385);
and UO_108 (O_108,N_15243,N_15797);
nand UO_109 (O_109,N_17012,N_17465);
and UO_110 (O_110,N_19795,N_19497);
or UO_111 (O_111,N_19545,N_17392);
or UO_112 (O_112,N_19081,N_17859);
and UO_113 (O_113,N_16128,N_18278);
and UO_114 (O_114,N_19445,N_19379);
nand UO_115 (O_115,N_17779,N_18083);
nand UO_116 (O_116,N_18789,N_17696);
or UO_117 (O_117,N_19991,N_16300);
nand UO_118 (O_118,N_17756,N_19333);
nand UO_119 (O_119,N_18400,N_17863);
and UO_120 (O_120,N_15099,N_18708);
and UO_121 (O_121,N_16007,N_15553);
nor UO_122 (O_122,N_19155,N_19124);
or UO_123 (O_123,N_16824,N_18760);
nor UO_124 (O_124,N_15017,N_18162);
nand UO_125 (O_125,N_17379,N_19629);
and UO_126 (O_126,N_15296,N_16870);
and UO_127 (O_127,N_18698,N_15036);
nor UO_128 (O_128,N_15134,N_17064);
nor UO_129 (O_129,N_15939,N_16187);
nor UO_130 (O_130,N_18677,N_17522);
nand UO_131 (O_131,N_18715,N_17489);
nand UO_132 (O_132,N_17453,N_18810);
nand UO_133 (O_133,N_17047,N_18629);
and UO_134 (O_134,N_15290,N_18601);
nor UO_135 (O_135,N_15209,N_17817);
nand UO_136 (O_136,N_19235,N_16237);
xnor UO_137 (O_137,N_17508,N_15969);
and UO_138 (O_138,N_15277,N_17430);
or UO_139 (O_139,N_15219,N_16614);
nand UO_140 (O_140,N_19238,N_16195);
or UO_141 (O_141,N_15993,N_15252);
nand UO_142 (O_142,N_17813,N_17989);
nand UO_143 (O_143,N_16292,N_18520);
nor UO_144 (O_144,N_15809,N_15753);
and UO_145 (O_145,N_17263,N_15677);
nor UO_146 (O_146,N_15642,N_16994);
nand UO_147 (O_147,N_16440,N_16953);
and UO_148 (O_148,N_16189,N_15968);
nand UO_149 (O_149,N_19211,N_19712);
or UO_150 (O_150,N_16465,N_15525);
or UO_151 (O_151,N_15437,N_18122);
nand UO_152 (O_152,N_16346,N_18765);
nor UO_153 (O_153,N_18668,N_15568);
nand UO_154 (O_154,N_17751,N_15772);
nand UO_155 (O_155,N_17543,N_17221);
nand UO_156 (O_156,N_15557,N_16344);
and UO_157 (O_157,N_16038,N_17580);
nand UO_158 (O_158,N_19150,N_18230);
nand UO_159 (O_159,N_15987,N_17003);
and UO_160 (O_160,N_16243,N_17265);
and UO_161 (O_161,N_15533,N_15002);
nand UO_162 (O_162,N_15349,N_19536);
nor UO_163 (O_163,N_18223,N_17656);
nand UO_164 (O_164,N_15980,N_17260);
nand UO_165 (O_165,N_18709,N_15878);
nor UO_166 (O_166,N_19910,N_15024);
and UO_167 (O_167,N_15732,N_18662);
nor UO_168 (O_168,N_15283,N_15374);
nand UO_169 (O_169,N_15752,N_16646);
xnor UO_170 (O_170,N_19508,N_16574);
nor UO_171 (O_171,N_15693,N_16772);
nand UO_172 (O_172,N_17850,N_15297);
and UO_173 (O_173,N_19197,N_18878);
nor UO_174 (O_174,N_18266,N_16339);
nand UO_175 (O_175,N_19967,N_19122);
nor UO_176 (O_176,N_18831,N_15358);
or UO_177 (O_177,N_15549,N_18562);
nand UO_178 (O_178,N_16039,N_16242);
nand UO_179 (O_179,N_19601,N_15327);
or UO_180 (O_180,N_19513,N_16168);
or UO_181 (O_181,N_17532,N_18355);
or UO_182 (O_182,N_15242,N_18947);
nand UO_183 (O_183,N_17041,N_18707);
nand UO_184 (O_184,N_19452,N_16282);
or UO_185 (O_185,N_18596,N_19477);
nor UO_186 (O_186,N_17944,N_19022);
nor UO_187 (O_187,N_19628,N_18904);
and UO_188 (O_188,N_17644,N_19807);
and UO_189 (O_189,N_17960,N_19944);
or UO_190 (O_190,N_19104,N_17721);
nand UO_191 (O_191,N_17481,N_18464);
nand UO_192 (O_192,N_18636,N_18090);
or UO_193 (O_193,N_16821,N_16632);
xnor UO_194 (O_194,N_18834,N_17726);
or UO_195 (O_195,N_18711,N_18503);
or UO_196 (O_196,N_15883,N_16756);
or UO_197 (O_197,N_17952,N_18914);
nor UO_198 (O_198,N_17896,N_17588);
or UO_199 (O_199,N_16909,N_19459);
and UO_200 (O_200,N_16768,N_15420);
and UO_201 (O_201,N_17790,N_16732);
and UO_202 (O_202,N_19222,N_16345);
nand UO_203 (O_203,N_15301,N_16901);
or UO_204 (O_204,N_17305,N_19947);
or UO_205 (O_205,N_19835,N_18665);
or UO_206 (O_206,N_19564,N_19689);
nand UO_207 (O_207,N_16303,N_16659);
nor UO_208 (O_208,N_15765,N_17499);
and UO_209 (O_209,N_19031,N_15331);
nor UO_210 (O_210,N_15418,N_16351);
and UO_211 (O_211,N_17821,N_17974);
nand UO_212 (O_212,N_18000,N_16661);
nand UO_213 (O_213,N_15895,N_18043);
nand UO_214 (O_214,N_16137,N_19411);
nor UO_215 (O_215,N_19655,N_17706);
and UO_216 (O_216,N_18965,N_19193);
nor UO_217 (O_217,N_15239,N_17879);
nor UO_218 (O_218,N_19303,N_15914);
nor UO_219 (O_219,N_17124,N_17727);
or UO_220 (O_220,N_19347,N_15066);
and UO_221 (O_221,N_19986,N_17390);
or UO_222 (O_222,N_19773,N_16514);
nor UO_223 (O_223,N_19364,N_17202);
and UO_224 (O_224,N_15270,N_16557);
and UO_225 (O_225,N_18523,N_18469);
nor UO_226 (O_226,N_17699,N_15789);
or UO_227 (O_227,N_19831,N_17538);
nor UO_228 (O_228,N_17548,N_18933);
nand UO_229 (O_229,N_15366,N_17278);
or UO_230 (O_230,N_17283,N_19381);
nand UO_231 (O_231,N_15545,N_16998);
nor UO_232 (O_232,N_18885,N_18141);
xnor UO_233 (O_233,N_19691,N_17559);
nor UO_234 (O_234,N_18455,N_16012);
and UO_235 (O_235,N_18643,N_19623);
or UO_236 (O_236,N_18669,N_15527);
nor UO_237 (O_237,N_18026,N_19468);
and UO_238 (O_238,N_17271,N_15396);
nor UO_239 (O_239,N_18500,N_18257);
and UO_240 (O_240,N_17894,N_19024);
and UO_241 (O_241,N_17592,N_19741);
and UO_242 (O_242,N_16660,N_19774);
nand UO_243 (O_243,N_19064,N_17631);
nor UO_244 (O_244,N_17217,N_18843);
and UO_245 (O_245,N_16882,N_17516);
and UO_246 (O_246,N_16822,N_15829);
xor UO_247 (O_247,N_17053,N_17069);
nor UO_248 (O_248,N_16420,N_19849);
nor UO_249 (O_249,N_19112,N_16079);
and UO_250 (O_250,N_17030,N_17378);
and UO_251 (O_251,N_17052,N_15014);
and UO_252 (O_252,N_19899,N_19383);
nand UO_253 (O_253,N_15000,N_18035);
nand UO_254 (O_254,N_17608,N_18496);
or UO_255 (O_255,N_18454,N_17860);
or UO_256 (O_256,N_17201,N_19685);
or UO_257 (O_257,N_17345,N_19591);
xor UO_258 (O_258,N_18493,N_15330);
or UO_259 (O_259,N_17561,N_19615);
nand UO_260 (O_260,N_16393,N_16879);
nor UO_261 (O_261,N_19253,N_17147);
and UO_262 (O_262,N_18738,N_17060);
nor UO_263 (O_263,N_17585,N_18199);
and UO_264 (O_264,N_15173,N_19259);
nand UO_265 (O_265,N_19350,N_16899);
or UO_266 (O_266,N_17761,N_18699);
or UO_267 (O_267,N_15139,N_19932);
nor UO_268 (O_268,N_17391,N_17661);
and UO_269 (O_269,N_16766,N_16025);
nor UO_270 (O_270,N_19474,N_19195);
nand UO_271 (O_271,N_16507,N_18435);
and UO_272 (O_272,N_18805,N_16640);
nand UO_273 (O_273,N_17852,N_16874);
or UO_274 (O_274,N_17777,N_18391);
nand UO_275 (O_275,N_16515,N_15257);
and UO_276 (O_276,N_16372,N_15653);
and UO_277 (O_277,N_17191,N_15083);
nand UO_278 (O_278,N_15302,N_18077);
or UO_279 (O_279,N_16531,N_19862);
or UO_280 (O_280,N_19787,N_19786);
nand UO_281 (O_281,N_15620,N_19729);
nor UO_282 (O_282,N_15361,N_16207);
and UO_283 (O_283,N_15060,N_17510);
and UO_284 (O_284,N_15352,N_15750);
and UO_285 (O_285,N_19679,N_17868);
nor UO_286 (O_286,N_19061,N_18369);
or UO_287 (O_287,N_18070,N_18906);
and UO_288 (O_288,N_15833,N_18081);
nand UO_289 (O_289,N_15792,N_16852);
nor UO_290 (O_290,N_19782,N_17326);
nor UO_291 (O_291,N_16075,N_19077);
and UO_292 (O_292,N_18979,N_18955);
nand UO_293 (O_293,N_15151,N_15554);
nand UO_294 (O_294,N_15652,N_17786);
nand UO_295 (O_295,N_18650,N_19788);
nand UO_296 (O_296,N_18305,N_16014);
and UO_297 (O_297,N_18630,N_19426);
and UO_298 (O_298,N_18440,N_15400);
and UO_299 (O_299,N_16382,N_16844);
nand UO_300 (O_300,N_19283,N_16807);
nand UO_301 (O_301,N_18412,N_17106);
and UO_302 (O_302,N_15764,N_16349);
nand UO_303 (O_303,N_16020,N_16133);
or UO_304 (O_304,N_18014,N_15921);
nor UO_305 (O_305,N_16516,N_18483);
nor UO_306 (O_306,N_16982,N_17975);
nand UO_307 (O_307,N_18600,N_16094);
nand UO_308 (O_308,N_19724,N_16833);
nand UO_309 (O_309,N_15212,N_15773);
nand UO_310 (O_310,N_15673,N_18809);
xor UO_311 (O_311,N_17571,N_16903);
or UO_312 (O_312,N_19804,N_17110);
nand UO_313 (O_313,N_18802,N_15254);
or UO_314 (O_314,N_19309,N_19470);
nor UO_315 (O_315,N_15015,N_17888);
nand UO_316 (O_316,N_17545,N_15595);
or UO_317 (O_317,N_19727,N_17834);
nand UO_318 (O_318,N_16234,N_17259);
nand UO_319 (O_319,N_19548,N_15021);
and UO_320 (O_320,N_17244,N_15233);
or UO_321 (O_321,N_18624,N_15803);
or UO_322 (O_322,N_19073,N_15991);
nor UO_323 (O_323,N_19071,N_16777);
or UO_324 (O_324,N_18652,N_19609);
nand UO_325 (O_325,N_16047,N_17484);
xor UO_326 (O_326,N_16127,N_19864);
or UO_327 (O_327,N_18253,N_16138);
or UO_328 (O_328,N_16375,N_16022);
or UO_329 (O_329,N_15088,N_15532);
or UO_330 (O_330,N_15517,N_16965);
nor UO_331 (O_331,N_16011,N_19941);
or UO_332 (O_332,N_15452,N_19659);
nor UO_333 (O_333,N_19936,N_15263);
and UO_334 (O_334,N_17930,N_19055);
or UO_335 (O_335,N_18084,N_17724);
or UO_336 (O_336,N_16323,N_16190);
and UO_337 (O_337,N_15704,N_17317);
nand UO_338 (O_338,N_15119,N_19054);
nand UO_339 (O_339,N_15222,N_19097);
nor UO_340 (O_340,N_18310,N_17066);
or UO_341 (O_341,N_18609,N_18040);
nor UO_342 (O_342,N_15316,N_17166);
nor UO_343 (O_343,N_18675,N_15160);
nand UO_344 (O_344,N_17501,N_18555);
xor UO_345 (O_345,N_17008,N_19549);
and UO_346 (O_346,N_18276,N_18539);
and UO_347 (O_347,N_15027,N_17179);
nor UO_348 (O_348,N_18327,N_18901);
and UO_349 (O_349,N_17054,N_15537);
or UO_350 (O_350,N_15538,N_17076);
and UO_351 (O_351,N_16122,N_17373);
or UO_352 (O_352,N_18036,N_17021);
or UO_353 (O_353,N_18864,N_18206);
nand UO_354 (O_354,N_17674,N_19242);
nand UO_355 (O_355,N_15678,N_19417);
or UO_356 (O_356,N_16692,N_15794);
nand UO_357 (O_357,N_16930,N_18477);
nand UO_358 (O_358,N_18150,N_17029);
nor UO_359 (O_359,N_17540,N_17527);
nor UO_360 (O_360,N_16169,N_19286);
or UO_361 (O_361,N_15972,N_15246);
nand UO_362 (O_362,N_18958,N_18212);
nor UO_363 (O_363,N_19768,N_15512);
nand UO_364 (O_364,N_19769,N_18663);
and UO_365 (O_365,N_16222,N_16206);
and UO_366 (O_366,N_17748,N_19879);
nor UO_367 (O_367,N_15491,N_15672);
and UO_368 (O_368,N_15612,N_18112);
and UO_369 (O_369,N_17258,N_16224);
nand UO_370 (O_370,N_18130,N_17370);
nor UO_371 (O_371,N_18786,N_16348);
xnor UO_372 (O_372,N_19147,N_17331);
and UO_373 (O_373,N_16320,N_17184);
nand UO_374 (O_374,N_19269,N_16194);
or UO_375 (O_375,N_16708,N_15583);
and UO_376 (O_376,N_19707,N_17822);
xor UO_377 (O_377,N_18872,N_15466);
nand UO_378 (O_378,N_17095,N_17840);
nor UO_379 (O_379,N_19393,N_19546);
nand UO_380 (O_380,N_16477,N_15949);
and UO_381 (O_381,N_18585,N_15266);
and UO_382 (O_382,N_16799,N_15928);
nor UO_383 (O_383,N_15394,N_17100);
or UO_384 (O_384,N_18263,N_19871);
nor UO_385 (O_385,N_16117,N_17846);
nor UO_386 (O_386,N_18450,N_16464);
nand UO_387 (O_387,N_15069,N_18976);
nand UO_388 (O_388,N_19044,N_15278);
or UO_389 (O_389,N_16435,N_16662);
and UO_390 (O_390,N_17294,N_19585);
nor UO_391 (O_391,N_18678,N_15070);
nor UO_392 (O_392,N_15234,N_18874);
and UO_393 (O_393,N_19931,N_16309);
nor UO_394 (O_394,N_16394,N_16157);
or UO_395 (O_395,N_17377,N_17870);
nor UO_396 (O_396,N_19358,N_17193);
and UO_397 (O_397,N_16954,N_19923);
nor UO_398 (O_398,N_17452,N_16257);
and UO_399 (O_399,N_15244,N_19858);
and UO_400 (O_400,N_17145,N_19686);
nand UO_401 (O_401,N_18104,N_15231);
or UO_402 (O_402,N_15728,N_18818);
and UO_403 (O_403,N_16726,N_17943);
and UO_404 (O_404,N_18823,N_15197);
nor UO_405 (O_405,N_16318,N_18016);
nor UO_406 (O_406,N_16993,N_19502);
nand UO_407 (O_407,N_15691,N_17094);
nor UO_408 (O_408,N_17606,N_18794);
nand UO_409 (O_409,N_15716,N_15579);
and UO_410 (O_410,N_19050,N_19144);
nand UO_411 (O_411,N_16484,N_19684);
nor UO_412 (O_412,N_19711,N_16296);
or UO_413 (O_413,N_17243,N_17582);
nand UO_414 (O_414,N_18606,N_15598);
and UO_415 (O_415,N_17919,N_17133);
nand UO_416 (O_416,N_18255,N_19698);
nor UO_417 (O_417,N_16827,N_18881);
and UO_418 (O_418,N_17990,N_19291);
or UO_419 (O_419,N_19052,N_16980);
or UO_420 (O_420,N_19883,N_15956);
nand UO_421 (O_421,N_15880,N_18549);
nor UO_422 (O_422,N_16907,N_18209);
nand UO_423 (O_423,N_17684,N_17921);
nor UO_424 (O_424,N_18728,N_16403);
nor UO_425 (O_425,N_17274,N_15255);
nand UO_426 (O_426,N_15810,N_15503);
and UO_427 (O_427,N_15093,N_19802);
nand UO_428 (O_428,N_17097,N_19436);
nor UO_429 (O_429,N_18264,N_17167);
nand UO_430 (O_430,N_18646,N_15974);
nor UO_431 (O_431,N_15966,N_16856);
nor UO_432 (O_432,N_17065,N_18515);
nand UO_433 (O_433,N_16266,N_17494);
nor UO_434 (O_434,N_15260,N_16703);
and UO_435 (O_435,N_18381,N_15611);
nor UO_436 (O_436,N_15047,N_17206);
nor UO_437 (O_437,N_17048,N_19688);
xnor UO_438 (O_438,N_16648,N_15042);
nor UO_439 (O_439,N_15940,N_19439);
and UO_440 (O_440,N_15641,N_19701);
and UO_441 (O_441,N_17196,N_18024);
nor UO_442 (O_442,N_15830,N_17507);
or UO_443 (O_443,N_17568,N_17366);
and UO_444 (O_444,N_17519,N_17675);
nand UO_445 (O_445,N_15767,N_16164);
or UO_446 (O_446,N_19007,N_19984);
nor UO_447 (O_447,N_15821,N_16791);
and UO_448 (O_448,N_15250,N_16212);
or UO_449 (O_449,N_16830,N_16728);
nand UO_450 (O_450,N_19570,N_17645);
nor UO_451 (O_451,N_16143,N_15646);
nand UO_452 (O_452,N_17577,N_16286);
nor UO_453 (O_453,N_18682,N_18586);
and UO_454 (O_454,N_17405,N_15488);
or UO_455 (O_455,N_19392,N_18931);
xnor UO_456 (O_456,N_18639,N_18769);
or UO_457 (O_457,N_18525,N_18071);
xor UO_458 (O_458,N_19517,N_15220);
and UO_459 (O_459,N_19086,N_15314);
or UO_460 (O_460,N_15056,N_16505);
or UO_461 (O_461,N_16379,N_18067);
nor UO_462 (O_462,N_19997,N_18186);
nor UO_463 (O_463,N_17738,N_17472);
nor UO_464 (O_464,N_17406,N_18128);
nand UO_465 (O_465,N_15344,N_17766);
nand UO_466 (O_466,N_18753,N_18838);
nor UO_467 (O_467,N_16126,N_18929);
nand UO_468 (O_468,N_15147,N_17403);
and UO_469 (O_469,N_15105,N_18820);
nand UO_470 (O_470,N_16831,N_17630);
nor UO_471 (O_471,N_15674,N_17410);
nor UO_472 (O_472,N_15226,N_19413);
nor UO_473 (O_473,N_16369,N_15032);
and UO_474 (O_474,N_15188,N_17648);
xor UO_475 (O_475,N_17009,N_18336);
and UO_476 (O_476,N_19485,N_16955);
xor UO_477 (O_477,N_18127,N_18868);
or UO_478 (O_478,N_15900,N_19895);
nand UO_479 (O_479,N_15749,N_18814);
nand UO_480 (O_480,N_18171,N_18808);
or UO_481 (O_481,N_16293,N_19406);
nor UO_482 (O_482,N_19654,N_15441);
nor UO_483 (O_483,N_16325,N_17000);
nand UO_484 (O_484,N_18157,N_15607);
and UO_485 (O_485,N_16975,N_18877);
nor UO_486 (O_486,N_19911,N_17351);
and UO_487 (O_487,N_15229,N_17463);
nand UO_488 (O_488,N_16838,N_18841);
and UO_489 (O_489,N_18739,N_17735);
and UO_490 (O_490,N_18853,N_16801);
and UO_491 (O_491,N_15681,N_18468);
or UO_492 (O_492,N_15339,N_15106);
nand UO_493 (O_493,N_16620,N_18120);
nand UO_494 (O_494,N_19187,N_15846);
nand UO_495 (O_495,N_18100,N_19836);
or UO_496 (O_496,N_16102,N_18544);
and UO_497 (O_497,N_19161,N_16600);
xnor UO_498 (O_498,N_16905,N_16272);
nor UO_499 (O_499,N_16295,N_16943);
or UO_500 (O_500,N_18082,N_15748);
and UO_501 (O_501,N_19343,N_15994);
or UO_502 (O_502,N_18351,N_15096);
nand UO_503 (O_503,N_19047,N_16865);
or UO_504 (O_504,N_15990,N_15843);
nand UO_505 (O_505,N_17947,N_16937);
nor UO_506 (O_506,N_17533,N_18466);
or UO_507 (O_507,N_17525,N_16742);
nand UO_508 (O_508,N_16654,N_15550);
or UO_509 (O_509,N_19710,N_19850);
nor UO_510 (O_510,N_15054,N_17937);
or UO_511 (O_511,N_19059,N_19140);
nand UO_512 (O_512,N_19066,N_17487);
nor UO_513 (O_513,N_18177,N_17117);
and UO_514 (O_514,N_15321,N_19014);
nand UO_515 (O_515,N_18258,N_19550);
and UO_516 (O_516,N_18227,N_16679);
nor UO_517 (O_517,N_17694,N_15285);
nor UO_518 (O_518,N_19535,N_19493);
nand UO_519 (O_519,N_17640,N_17480);
nor UO_520 (O_520,N_17603,N_16361);
and UO_521 (O_521,N_16846,N_16065);
or UO_522 (O_522,N_17150,N_18564);
nand UO_523 (O_523,N_15543,N_15867);
nor UO_524 (O_524,N_16405,N_16563);
and UO_525 (O_525,N_16932,N_18706);
nand UO_526 (O_526,N_16804,N_18220);
nand UO_527 (O_527,N_16125,N_19926);
or UO_528 (O_528,N_17273,N_16962);
nor UO_529 (O_529,N_15697,N_19945);
nand UO_530 (O_530,N_19040,N_19376);
or UO_531 (O_531,N_18970,N_18546);
nor UO_532 (O_532,N_16926,N_18299);
nand UO_533 (O_533,N_19216,N_17589);
nor UO_534 (O_534,N_18376,N_15205);
or UO_535 (O_535,N_19205,N_19897);
or UO_536 (O_536,N_18107,N_15562);
and UO_537 (O_537,N_18414,N_19290);
and UO_538 (O_538,N_15798,N_17677);
and UO_539 (O_539,N_17241,N_17639);
nor UO_540 (O_540,N_19265,N_17611);
and UO_541 (O_541,N_18094,N_16028);
and UO_542 (O_542,N_15086,N_16594);
or UO_543 (O_543,N_15081,N_16248);
nand UO_544 (O_544,N_17848,N_17584);
nand UO_545 (O_545,N_19884,N_16040);
nor UO_546 (O_546,N_16305,N_15665);
nand UO_547 (O_547,N_17972,N_19526);
or UO_548 (O_548,N_17513,N_18494);
and UO_549 (O_549,N_18882,N_16816);
nand UO_550 (O_550,N_19761,N_15917);
and UO_551 (O_551,N_19043,N_19045);
nand UO_552 (O_552,N_19421,N_19232);
nand UO_553 (O_553,N_19427,N_18502);
nand UO_554 (O_554,N_19657,N_19301);
nand UO_555 (O_555,N_15332,N_15819);
nand UO_556 (O_556,N_15982,N_15778);
or UO_557 (O_557,N_17077,N_18136);
or UO_558 (O_558,N_19577,N_16721);
nor UO_559 (O_559,N_18179,N_15034);
and UO_560 (O_560,N_19718,N_16097);
nor UO_561 (O_561,N_16843,N_16267);
and UO_562 (O_562,N_18621,N_19605);
and UO_563 (O_563,N_18557,N_16274);
nand UO_564 (O_564,N_15952,N_19213);
nand UO_565 (O_565,N_17825,N_18243);
nand UO_566 (O_566,N_18417,N_19034);
nor UO_567 (O_567,N_18865,N_19037);
nor UO_568 (O_568,N_19298,N_17194);
nand UO_569 (O_569,N_17662,N_18149);
xnor UO_570 (O_570,N_19904,N_18824);
or UO_571 (O_571,N_18971,N_17215);
or UO_572 (O_572,N_19201,N_16067);
or UO_573 (O_573,N_16245,N_16753);
or UO_574 (O_574,N_19455,N_16327);
nand UO_575 (O_575,N_16139,N_15788);
or UO_576 (O_576,N_19438,N_17121);
nand UO_577 (O_577,N_17090,N_16045);
and UO_578 (O_578,N_15790,N_15502);
nand UO_579 (O_579,N_19606,N_16335);
nand UO_580 (O_580,N_17423,N_16685);
nor UO_581 (O_581,N_19403,N_17720);
nand UO_582 (O_582,N_18487,N_15937);
nand UO_583 (O_583,N_18776,N_19412);
and UO_584 (O_584,N_18531,N_18019);
xnor UO_585 (O_585,N_16407,N_17212);
or UO_586 (O_586,N_19764,N_19987);
xor UO_587 (O_587,N_18078,N_19728);
or UO_588 (O_588,N_19390,N_16495);
and UO_589 (O_589,N_18062,N_17329);
and UO_590 (O_590,N_19958,N_16432);
and UO_591 (O_591,N_17732,N_15606);
and UO_592 (O_592,N_16630,N_16588);
xnor UO_593 (O_593,N_19217,N_18146);
and UO_594 (O_594,N_17743,N_18667);
nand UO_595 (O_595,N_15999,N_18115);
or UO_596 (O_596,N_18687,N_17087);
or UO_597 (O_597,N_19273,N_19320);
or UO_598 (O_598,N_19172,N_19437);
or UO_599 (O_599,N_16021,N_18889);
nand UO_600 (O_600,N_19976,N_18001);
or UO_601 (O_601,N_16938,N_15800);
nand UO_602 (O_602,N_15265,N_16444);
nand UO_603 (O_603,N_18403,N_15961);
nand UO_604 (O_604,N_19083,N_17016);
nor UO_605 (O_605,N_18797,N_19896);
nand UO_606 (O_606,N_15238,N_18324);
and UO_607 (O_607,N_15464,N_15153);
nand UO_608 (O_608,N_15820,N_19483);
or UO_609 (O_609,N_16355,N_18799);
nand UO_610 (O_610,N_16216,N_16214);
nor UO_611 (O_611,N_16536,N_15943);
or UO_612 (O_612,N_15370,N_15904);
nor UO_613 (O_613,N_17300,N_19506);
or UO_614 (O_614,N_16891,N_15508);
and UO_615 (O_615,N_18983,N_18842);
nand UO_616 (O_616,N_16560,N_17986);
and UO_617 (O_617,N_17929,N_18695);
and UO_618 (O_618,N_18119,N_17409);
nand UO_619 (O_619,N_17174,N_15299);
and UO_620 (O_620,N_15080,N_19363);
nand UO_621 (O_621,N_19880,N_15392);
and UO_622 (O_622,N_18840,N_15354);
and UO_623 (O_623,N_16701,N_19975);
and UO_624 (O_624,N_15120,N_16285);
nand UO_625 (O_625,N_19510,N_18205);
and UO_626 (O_626,N_18697,N_19642);
or UO_627 (O_627,N_16152,N_19907);
and UO_628 (O_628,N_15165,N_18461);
or UO_629 (O_629,N_18294,N_17778);
nor UO_630 (O_630,N_16106,N_15476);
and UO_631 (O_631,N_19739,N_17013);
nand UO_632 (O_632,N_17977,N_15998);
and UO_633 (O_633,N_18771,N_18499);
or UO_634 (O_634,N_15718,N_17264);
nand UO_635 (O_635,N_19117,N_17512);
and UO_636 (O_636,N_19794,N_17902);
or UO_637 (O_637,N_16252,N_17230);
xor UO_638 (O_638,N_19593,N_19640);
and UO_639 (O_639,N_15648,N_19543);
nand UO_640 (O_640,N_18517,N_17700);
nor UO_641 (O_641,N_18833,N_18430);
nor UO_642 (O_642,N_17040,N_15138);
and UO_643 (O_643,N_19011,N_18283);
and UO_644 (O_644,N_15643,N_18160);
nor UO_645 (O_645,N_19738,N_16493);
and UO_646 (O_646,N_15610,N_16991);
nand UO_647 (O_647,N_19604,N_16716);
nor UO_648 (O_648,N_19021,N_16621);
nand UO_649 (O_649,N_16553,N_18628);
nor UO_650 (O_650,N_19928,N_18387);
nand UO_651 (O_651,N_18007,N_19557);
and UO_652 (O_652,N_15720,N_18518);
nand UO_653 (O_653,N_15126,N_15811);
nand UO_654 (O_654,N_16881,N_17926);
and UO_655 (O_655,N_19270,N_15919);
or UO_656 (O_656,N_19520,N_16510);
or UO_657 (O_657,N_16615,N_19530);
nand UO_658 (O_658,N_15225,N_19713);
or UO_659 (O_659,N_15567,N_19859);
nor UO_660 (O_660,N_16076,N_19157);
xor UO_661 (O_661,N_17467,N_18325);
nand UO_662 (O_662,N_15814,N_18792);
and UO_663 (O_663,N_18784,N_19395);
and UO_664 (O_664,N_15578,N_15986);
nor UO_665 (O_665,N_15319,N_16458);
or UO_666 (O_666,N_18627,N_19812);
nand UO_667 (O_667,N_18702,N_19359);
or UO_668 (O_668,N_15451,N_18615);
and UO_669 (O_669,N_16841,N_19842);
and UO_670 (O_670,N_15818,N_16974);
and UO_671 (O_671,N_15127,N_17324);
or UO_672 (O_672,N_19429,N_17419);
nor UO_673 (O_673,N_15028,N_17627);
and UO_674 (O_674,N_19002,N_19948);
nor UO_675 (O_675,N_16262,N_15492);
nand UO_676 (O_676,N_16568,N_17886);
and UO_677 (O_677,N_15582,N_15615);
nand UO_678 (O_678,N_19743,N_15116);
nor UO_679 (O_679,N_16561,N_19620);
or UO_680 (O_680,N_19519,N_18770);
nand UO_681 (O_681,N_15671,N_16914);
and UO_682 (O_682,N_15875,N_15362);
nand UO_683 (O_683,N_16526,N_16334);
nor UO_684 (O_684,N_19625,N_19498);
nor UO_685 (O_685,N_17875,N_15409);
nand UO_686 (O_686,N_18056,N_19631);
or UO_687 (O_687,N_15667,N_15712);
or UO_688 (O_688,N_16987,N_19357);
and UO_689 (O_689,N_15346,N_15858);
or UO_690 (O_690,N_17749,N_16219);
and UO_691 (O_691,N_15132,N_17438);
nand UO_692 (O_692,N_19108,N_16787);
nor UO_693 (O_693,N_18642,N_18038);
or UO_694 (O_694,N_17932,N_18755);
nand UO_695 (O_695,N_18658,N_17031);
and UO_696 (O_696,N_18567,N_16091);
nor UO_697 (O_697,N_15011,N_19454);
nor UO_698 (O_698,N_15484,N_18724);
nor UO_699 (O_699,N_16573,N_15886);
nor UO_700 (O_700,N_16482,N_17006);
and UO_701 (O_701,N_17394,N_19571);
or UO_702 (O_702,N_18032,N_18195);
and UO_703 (O_703,N_19142,N_18835);
and UO_704 (O_704,N_15016,N_18522);
nand UO_705 (O_705,N_18169,N_15180);
nand UO_706 (O_706,N_15783,N_15862);
nand UO_707 (O_707,N_18409,N_18986);
nor UO_708 (O_708,N_15058,N_18302);
nand UO_709 (O_709,N_18311,N_17246);
and UO_710 (O_710,N_16919,N_16304);
and UO_711 (O_711,N_18846,N_17374);
and UO_712 (O_712,N_15143,N_16871);
or UO_713 (O_713,N_18740,N_19775);
and UO_714 (O_714,N_15812,N_17893);
nor UO_715 (O_715,N_19171,N_16474);
and UO_716 (O_716,N_15528,N_17441);
or UO_717 (O_717,N_15908,N_15347);
or UO_718 (O_718,N_17554,N_17600);
nand UO_719 (O_719,N_18618,N_19678);
and UO_720 (O_720,N_17924,N_18994);
and UO_721 (O_721,N_15920,N_17961);
nand UO_722 (O_722,N_18061,N_16636);
nand UO_723 (O_723,N_18337,N_19048);
nand UO_724 (O_724,N_18096,N_16806);
and UO_725 (O_725,N_16984,N_18576);
nor UO_726 (O_726,N_16723,N_18170);
and UO_727 (O_727,N_16313,N_19183);
or UO_728 (O_728,N_17858,N_15530);
nand UO_729 (O_729,N_18584,N_15318);
or UO_730 (O_730,N_19174,N_18222);
and UO_731 (O_731,N_16888,N_15852);
nand UO_732 (O_732,N_17633,N_18908);
nand UO_733 (O_733,N_15689,N_15523);
or UO_734 (O_734,N_18962,N_19237);
xor UO_735 (O_735,N_15022,N_18861);
nor UO_736 (O_736,N_19130,N_16572);
or UO_737 (O_737,N_16567,N_15325);
nand UO_738 (O_738,N_15701,N_15387);
and UO_739 (O_739,N_15779,N_18423);
and UO_740 (O_740,N_18811,N_15618);
xnor UO_741 (O_741,N_16604,N_17182);
nor UO_742 (O_742,N_18952,N_15632);
nand UO_743 (O_743,N_18261,N_19168);
and UO_744 (O_744,N_16951,N_17357);
or UO_745 (O_745,N_16539,N_19813);
nand UO_746 (O_746,N_19467,N_15844);
and UO_747 (O_747,N_15658,N_19749);
and UO_748 (O_748,N_15861,N_19093);
nor UO_749 (O_749,N_17425,N_18912);
nand UO_750 (O_750,N_17676,N_18866);
and UO_751 (O_751,N_16118,N_19258);
or UO_752 (O_752,N_17470,N_18457);
and UO_753 (O_753,N_19537,N_15787);
and UO_754 (O_754,N_15341,N_18306);
nor UO_755 (O_755,N_19404,N_15406);
or UO_756 (O_756,N_19337,N_19875);
and UO_757 (O_757,N_17478,N_15916);
nand UO_758 (O_758,N_17951,N_16631);
or UO_759 (O_759,N_18887,N_15340);
and UO_760 (O_760,N_19461,N_16239);
and UO_761 (O_761,N_19328,N_16743);
or UO_762 (O_762,N_19784,N_17413);
nand UO_763 (O_763,N_15312,N_19463);
or UO_764 (O_764,N_19793,N_18727);
nand UO_765 (O_765,N_17309,N_16100);
and UO_766 (O_766,N_16972,N_17776);
nor UO_767 (O_767,N_19198,N_16936);
nor UO_768 (O_768,N_19178,N_15019);
and UO_769 (O_769,N_15731,N_17605);
nor UO_770 (O_770,N_18396,N_18935);
nor UO_771 (O_771,N_17760,N_18599);
nand UO_772 (O_772,N_18072,N_18453);
nor UO_773 (O_773,N_15249,N_16298);
or UO_774 (O_774,N_17015,N_16933);
and UO_775 (O_775,N_18259,N_17033);
or UO_776 (O_776,N_17074,N_16570);
and UO_777 (O_777,N_18182,N_17753);
and UO_778 (O_778,N_17344,N_17401);
nand UO_779 (O_779,N_15211,N_15414);
nand UO_780 (O_780,N_16036,N_16099);
or UO_781 (O_781,N_17810,N_18705);
or UO_782 (O_782,N_15288,N_16198);
nand UO_783 (O_783,N_15506,N_17387);
nand UO_784 (O_784,N_16098,N_17332);
xor UO_785 (O_785,N_15603,N_16306);
and UO_786 (O_786,N_15813,N_18593);
nand UO_787 (O_787,N_18757,N_17650);
nor UO_788 (O_788,N_17995,N_18188);
nand UO_789 (O_789,N_19572,N_16461);
or UO_790 (O_790,N_18431,N_17551);
nand UO_791 (O_791,N_19837,N_19974);
or UO_792 (O_792,N_16322,N_19597);
nor UO_793 (O_793,N_19203,N_17399);
or UO_794 (O_794,N_18091,N_16616);
xnor UO_795 (O_795,N_16380,N_17722);
nand UO_796 (O_796,N_18481,N_16008);
or UO_797 (O_797,N_15453,N_19566);
nand UO_798 (O_798,N_18894,N_19342);
xnor UO_799 (O_799,N_18554,N_19339);
or UO_800 (O_800,N_15942,N_17874);
and UO_801 (O_801,N_16452,N_16488);
or UO_802 (O_802,N_15140,N_17856);
nor UO_803 (O_803,N_18201,N_15470);
and UO_804 (O_804,N_19100,N_17839);
and UO_805 (O_805,N_15446,N_19330);
nand UO_806 (O_806,N_15805,N_17654);
nand UO_807 (O_807,N_18475,N_19087);
nand UO_808 (O_808,N_19733,N_17075);
or UO_809 (O_809,N_16324,N_16217);
nand UO_810 (O_810,N_19826,N_19632);
and UO_811 (O_811,N_15569,N_16053);
or UO_812 (O_812,N_18967,N_19422);
nor UO_813 (O_813,N_16326,N_15494);
xnor UO_814 (O_814,N_15510,N_16332);
nor UO_815 (O_815,N_19569,N_18068);
nor UO_816 (O_816,N_18298,N_16030);
or UO_817 (O_817,N_16460,N_16694);
and UO_818 (O_818,N_15755,N_19058);
or UO_819 (O_819,N_15328,N_18598);
and UO_820 (O_820,N_18485,N_16386);
nor UO_821 (O_821,N_19218,N_15481);
nand UO_822 (O_822,N_17437,N_15992);
or UO_823 (O_823,N_18117,N_17758);
and UO_824 (O_824,N_18680,N_18611);
and UO_825 (O_825,N_15450,N_15541);
nand UO_826 (O_826,N_15675,N_16815);
nand UO_827 (O_827,N_16210,N_16399);
nor UO_828 (O_828,N_19499,N_18527);
xor UO_829 (O_829,N_15873,N_17448);
nand UO_830 (O_830,N_16836,N_16864);
or UO_831 (O_831,N_17687,N_16658);
or UO_832 (O_832,N_19963,N_15548);
or UO_833 (O_833,N_17652,N_16535);
nor UO_834 (O_834,N_17155,N_15026);
nand UO_835 (O_835,N_19874,N_16209);
nor UO_836 (O_836,N_18884,N_18625);
nor UO_837 (O_837,N_19255,N_17411);
xor UO_838 (O_838,N_16370,N_15981);
nor UO_839 (O_839,N_16160,N_16530);
nand UO_840 (O_840,N_18462,N_18859);
and UO_841 (O_841,N_16941,N_16789);
nor UO_842 (O_842,N_16851,N_18854);
nand UO_843 (O_843,N_16913,N_19448);
xor UO_844 (O_844,N_15148,N_18583);
nand UO_845 (O_845,N_15662,N_16782);
or UO_846 (O_846,N_19725,N_17987);
and UO_847 (O_847,N_19873,N_17549);
nor UO_848 (O_848,N_18641,N_16592);
nand UO_849 (O_849,N_16130,N_18913);
and UO_850 (O_850,N_19619,N_18353);
nand UO_851 (O_851,N_15841,N_15625);
and UO_852 (O_852,N_19834,N_17641);
or UO_853 (O_853,N_19370,N_16192);
nand UO_854 (O_854,N_16605,N_15593);
or UO_855 (O_855,N_16223,N_19616);
or UO_856 (O_856,N_15967,N_15082);
or UO_857 (O_857,N_18374,N_16450);
and UO_858 (O_858,N_19751,N_15587);
nand UO_859 (O_859,N_15879,N_19418);
xor UO_860 (O_860,N_16765,N_17836);
and UO_861 (O_861,N_18415,N_15713);
and UO_862 (O_862,N_15150,N_17198);
nand UO_863 (O_863,N_17130,N_16672);
and UO_864 (O_864,N_18528,N_18350);
nand UO_865 (O_865,N_15957,N_16376);
and UO_866 (O_866,N_19224,N_18418);
or UO_867 (O_867,N_19999,N_19966);
nor UO_868 (O_868,N_16371,N_17020);
or UO_869 (O_869,N_16725,N_18719);
nand UO_870 (O_870,N_16087,N_19182);
or UO_871 (O_871,N_19994,N_19523);
and UO_872 (O_872,N_19644,N_15334);
nand UO_873 (O_873,N_16569,N_17144);
nor UO_874 (O_874,N_18612,N_15149);
xnor UO_875 (O_875,N_19177,N_17770);
or UO_876 (O_876,N_19906,N_19257);
and UO_877 (O_877,N_15194,N_15473);
or UO_878 (O_878,N_15710,N_17976);
and UO_879 (O_879,N_19409,N_15078);
nor UO_880 (O_880,N_15141,N_16719);
and UO_881 (O_881,N_18393,N_16341);
xnor UO_882 (O_882,N_16156,N_18953);
nand UO_883 (O_883,N_18510,N_16311);
nor UO_884 (O_884,N_15432,N_19141);
nand UO_885 (O_885,N_16340,N_16082);
and UO_886 (O_886,N_15426,N_17067);
nand UO_887 (O_887,N_18342,N_16607);
xnor UO_888 (O_888,N_18752,N_19241);
nor UO_889 (O_889,N_19015,N_16817);
or UO_890 (O_890,N_18559,N_16653);
nand UO_891 (O_891,N_15656,N_19068);
or UO_892 (O_892,N_15596,N_16596);
nor UO_893 (O_893,N_19446,N_17787);
nand UO_894 (O_894,N_18368,N_16035);
nor UO_895 (O_895,N_19785,N_19617);
and UO_896 (O_896,N_15585,N_19449);
or UO_897 (O_897,N_15699,N_17686);
or UO_898 (O_898,N_15375,N_19332);
nand UO_899 (O_899,N_15597,N_18588);
or UO_900 (O_900,N_19340,N_17638);
nor UO_901 (O_901,N_15955,N_18943);
or UO_902 (O_902,N_15098,N_17578);
and UO_903 (O_903,N_16281,N_15262);
and UO_904 (O_904,N_17811,N_16489);
nor UO_905 (O_905,N_18742,N_18547);
nor UO_906 (O_906,N_16033,N_15191);
nand UO_907 (O_907,N_18203,N_16855);
nor UO_908 (O_908,N_15053,N_17955);
nor UO_909 (O_909,N_15947,N_16112);
nor UO_910 (O_910,N_19652,N_15114);
or UO_911 (O_911,N_15115,N_18910);
or UO_912 (O_912,N_16670,N_15682);
xor UO_913 (O_913,N_15281,N_16041);
nor UO_914 (O_914,N_16299,N_15730);
nand UO_915 (O_915,N_16288,N_17049);
nor UO_916 (O_916,N_16820,N_19028);
or UO_917 (O_917,N_15317,N_19008);
or UO_918 (O_918,N_15664,N_18095);
or UO_919 (O_919,N_15007,N_16709);
nand UO_920 (O_920,N_16086,N_15690);
nor UO_921 (O_921,N_15398,N_18399);
or UO_922 (O_922,N_16459,N_17238);
nor UO_923 (O_923,N_17180,N_15012);
nor UO_924 (O_924,N_18563,N_16696);
nor UO_925 (O_925,N_16231,N_15757);
xnor UO_926 (O_926,N_19734,N_17468);
and UO_927 (O_927,N_19647,N_18159);
and UO_928 (O_928,N_15931,N_18548);
xnor UO_929 (O_929,N_17704,N_19220);
and UO_930 (O_930,N_15739,N_16733);
nand UO_931 (O_931,N_18224,N_18319);
or UO_932 (O_932,N_17725,N_15357);
nand UO_933 (O_933,N_18285,N_17705);
and UO_934 (O_934,N_18291,N_16666);
or UO_935 (O_935,N_15294,N_18932);
and UO_936 (O_936,N_19316,N_18829);
or UO_937 (O_937,N_19900,N_16263);
and UO_938 (O_938,N_19432,N_19414);
nor UO_939 (O_939,N_17941,N_16957);
nand UO_940 (O_940,N_19854,N_19956);
or UO_941 (O_941,N_16188,N_17051);
or UO_942 (O_942,N_17546,N_18168);
or UO_943 (O_943,N_16896,N_16287);
or UO_944 (O_944,N_18408,N_19962);
or UO_945 (O_945,N_17939,N_15558);
xor UO_946 (O_946,N_16802,N_16534);
nor UO_947 (O_947,N_19544,N_18949);
nand UO_948 (O_948,N_15828,N_17226);
nand UO_949 (O_949,N_15350,N_17702);
nor UO_950 (O_950,N_19915,N_17969);
nand UO_951 (O_951,N_17092,N_16096);
nor UO_952 (O_952,N_16863,N_16509);
and UO_953 (O_953,N_19072,N_18495);
nand UO_954 (O_954,N_17765,N_18514);
xor UO_955 (O_955,N_16254,N_16582);
nor UO_956 (O_956,N_17312,N_17328);
nor UO_957 (O_957,N_15381,N_16665);
nor UO_958 (O_958,N_19188,N_16835);
or UO_959 (O_959,N_19581,N_16294);
and UO_960 (O_960,N_17426,N_16163);
and UO_961 (O_961,N_17731,N_17539);
or UO_962 (O_962,N_16316,N_19914);
nand UO_963 (O_963,N_19277,N_16555);
or UO_964 (O_964,N_18655,N_18915);
nor UO_965 (O_965,N_15065,N_18950);
and UO_966 (O_966,N_15351,N_16009);
nand UO_967 (O_967,N_17093,N_19965);
and UO_968 (O_968,N_18080,N_16103);
nor UO_969 (O_969,N_16060,N_19630);
and UO_970 (O_970,N_17830,N_18063);
and UO_971 (O_971,N_15214,N_16637);
xnor UO_972 (O_972,N_17797,N_15343);
nand UO_973 (O_973,N_17010,N_15649);
nor UO_974 (O_974,N_15574,N_19925);
nor UO_975 (O_975,N_19872,N_17653);
nor UO_976 (O_976,N_16754,N_15694);
or UO_977 (O_977,N_16898,N_18459);
nor UO_978 (O_978,N_18075,N_17908);
nor UO_979 (O_979,N_19151,N_18613);
or UO_980 (O_980,N_17190,N_15824);
nand UO_981 (O_981,N_19700,N_17270);
nor UO_982 (O_982,N_15456,N_15705);
or UO_983 (O_983,N_15025,N_19191);
nand UO_984 (O_984,N_15985,N_15605);
nand UO_985 (O_985,N_17299,N_19353);
or UO_986 (O_986,N_19709,N_15628);
or UO_987 (O_987,N_16436,N_15010);
nand UO_988 (O_988,N_19026,N_16512);
xor UO_989 (O_989,N_19663,N_19504);
nor UO_990 (O_990,N_17376,N_18999);
nor UO_991 (O_991,N_17431,N_15471);
nand UO_992 (O_992,N_18064,N_15877);
and UO_993 (O_993,N_16221,N_16414);
nor UO_994 (O_994,N_16713,N_17980);
nand UO_995 (O_995,N_18113,N_15145);
nand UO_996 (O_996,N_16017,N_16774);
nor UO_997 (O_997,N_17088,N_18046);
xnor UO_998 (O_998,N_17869,N_17716);
nor UO_999 (O_999,N_16861,N_16072);
nand UO_1000 (O_1000,N_15684,N_15483);
xnor UO_1001 (O_1001,N_15337,N_18726);
and UO_1002 (O_1002,N_16729,N_19264);
nor UO_1003 (O_1003,N_15845,N_17767);
nand UO_1004 (O_1004,N_16876,N_18126);
nand UO_1005 (O_1005,N_17427,N_19918);
nor UO_1006 (O_1006,N_15723,N_19525);
or UO_1007 (O_1007,N_15190,N_15478);
and UO_1008 (O_1008,N_17136,N_17055);
or UO_1009 (O_1009,N_19909,N_15575);
nand UO_1010 (O_1010,N_16587,N_17799);
nor UO_1011 (O_1011,N_19622,N_16781);
or UO_1012 (O_1012,N_16966,N_16291);
nand UO_1013 (O_1013,N_15206,N_15303);
and UO_1014 (O_1014,N_16811,N_16032);
or UO_1015 (O_1015,N_15457,N_19254);
nor UO_1016 (O_1016,N_17157,N_16062);
nor UO_1017 (O_1017,N_16508,N_17139);
nor UO_1018 (O_1018,N_15411,N_19384);
nand UO_1019 (O_1019,N_19063,N_18280);
nor UO_1020 (O_1020,N_18565,N_15542);
and UO_1021 (O_1021,N_16230,N_17954);
and UO_1022 (O_1022,N_17984,N_16911);
or UO_1023 (O_1023,N_17752,N_15474);
nand UO_1024 (O_1024,N_18262,N_15560);
or UO_1025 (O_1025,N_19078,N_19401);
nand UO_1026 (O_1026,N_19766,N_16973);
or UO_1027 (O_1027,N_15072,N_17319);
or UO_1028 (O_1028,N_17701,N_16900);
and UO_1029 (O_1029,N_17775,N_17068);
nand UO_1030 (O_1030,N_16449,N_15235);
and UO_1031 (O_1031,N_19716,N_15280);
or UO_1032 (O_1032,N_17880,N_17432);
nand UO_1033 (O_1033,N_17535,N_19067);
and UO_1034 (O_1034,N_19759,N_18954);
nor UO_1035 (O_1035,N_16378,N_16317);
or UO_1036 (O_1036,N_18345,N_16853);
or UO_1037 (O_1037,N_16959,N_17809);
and UO_1038 (O_1038,N_18674,N_16289);
or UO_1039 (O_1039,N_17341,N_16442);
nor UO_1040 (O_1040,N_17398,N_16069);
and UO_1041 (O_1041,N_18603,N_15536);
or UO_1042 (O_1042,N_18346,N_16923);
nor UO_1043 (O_1043,N_17587,N_16960);
and UO_1044 (O_1044,N_15592,N_19199);
or UO_1045 (O_1045,N_18537,N_17579);
or UO_1046 (O_1046,N_15905,N_19304);
nor UO_1047 (O_1047,N_15518,N_15851);
or UO_1048 (O_1048,N_18501,N_17816);
or UO_1049 (O_1049,N_19553,N_17322);
and UO_1050 (O_1050,N_16823,N_16247);
or UO_1051 (O_1051,N_18178,N_17759);
or UO_1052 (O_1052,N_18340,N_19294);
or UO_1053 (O_1053,N_17884,N_19580);
nor UO_1054 (O_1054,N_19170,N_17454);
nor UO_1055 (O_1055,N_17872,N_16271);
or UO_1056 (O_1056,N_17707,N_19542);
nor UO_1057 (O_1057,N_17433,N_15780);
or UO_1058 (O_1058,N_18509,N_15376);
and UO_1059 (O_1059,N_18511,N_19533);
or UO_1060 (O_1060,N_19215,N_15185);
and UO_1061 (O_1061,N_17835,N_15839);
nor UO_1062 (O_1062,N_17566,N_18879);
and UO_1063 (O_1063,N_15529,N_15962);
nand UO_1064 (O_1064,N_18762,N_16121);
nor UO_1065 (O_1065,N_18002,N_15064);
or UO_1066 (O_1066,N_17383,N_15609);
nor UO_1067 (O_1067,N_19166,N_19808);
and UO_1068 (O_1068,N_16059,N_19758);
nand UO_1069 (O_1069,N_17247,N_19408);
nand UO_1070 (O_1070,N_19641,N_18192);
and UO_1071 (O_1071,N_18645,N_17086);
nand UO_1072 (O_1072,N_18569,N_18787);
nand UO_1073 (O_1073,N_16409,N_18286);
and UO_1074 (O_1074,N_18634,N_17105);
nand UO_1075 (O_1075,N_17320,N_17801);
or UO_1076 (O_1076,N_18385,N_16635);
or UO_1077 (O_1077,N_18432,N_16918);
nor UO_1078 (O_1078,N_18356,N_19501);
nand UO_1079 (O_1079,N_17708,N_16678);
xnor UO_1080 (O_1080,N_18785,N_18890);
or UO_1081 (O_1081,N_15192,N_17812);
or UO_1082 (O_1082,N_19338,N_15761);
and UO_1083 (O_1083,N_17288,N_16803);
nor UO_1084 (O_1084,N_17602,N_17028);
or UO_1085 (O_1085,N_15033,N_17509);
nand UO_1086 (O_1086,N_16466,N_16887);
nand UO_1087 (O_1087,N_17449,N_19146);
or UO_1088 (O_1088,N_17192,N_16749);
and UO_1089 (O_1089,N_18470,N_18279);
and UO_1090 (O_1090,N_18703,N_17338);
nand UO_1091 (O_1091,N_15372,N_16176);
and UO_1092 (O_1092,N_16996,N_16434);
and UO_1093 (O_1093,N_19056,N_15599);
and UO_1094 (O_1094,N_19843,N_17330);
and UO_1095 (O_1095,N_17291,N_18328);
and UO_1096 (O_1096,N_15910,N_16149);
and UO_1097 (O_1097,N_16417,N_17327);
or UO_1098 (O_1098,N_19833,N_15722);
xnor UO_1099 (O_1099,N_16958,N_16227);
and UO_1100 (O_1100,N_16691,N_15953);
nor UO_1101 (O_1101,N_18977,N_15817);
or UO_1102 (O_1102,N_18898,N_16667);
nand UO_1103 (O_1103,N_16350,N_18540);
nand UO_1104 (O_1104,N_15763,N_15715);
and UO_1105 (O_1105,N_18446,N_15333);
nand UO_1106 (O_1106,N_16935,N_18815);
or UO_1107 (O_1107,N_17388,N_18106);
nor UO_1108 (O_1108,N_18957,N_16867);
or UO_1109 (O_1109,N_17343,N_19669);
or UO_1110 (O_1110,N_15970,N_15449);
or UO_1111 (O_1111,N_15001,N_19653);
nand UO_1112 (O_1112,N_18076,N_19148);
nand UO_1113 (O_1113,N_17945,N_17763);
xnor UO_1114 (O_1114,N_15356,N_19820);
and UO_1115 (O_1115,N_19491,N_15199);
or UO_1116 (O_1116,N_17208,N_19486);
nand UO_1117 (O_1117,N_15482,N_15412);
nand UO_1118 (O_1118,N_18551,N_15874);
nand UO_1119 (O_1119,N_17239,N_17232);
or UO_1120 (O_1120,N_16693,N_19348);
nor UO_1121 (O_1121,N_15218,N_15434);
or UO_1122 (O_1122,N_16034,N_15062);
and UO_1123 (O_1123,N_16908,N_19120);
and UO_1124 (O_1124,N_16328,N_15371);
or UO_1125 (O_1125,N_17889,N_18216);
nor UO_1126 (O_1126,N_17151,N_19888);
nand UO_1127 (O_1127,N_19416,N_19603);
nor UO_1128 (O_1128,N_15079,N_18145);
and UO_1129 (O_1129,N_17214,N_16109);
nor UO_1130 (O_1130,N_16544,N_15898);
nand UO_1131 (O_1131,N_18219,N_18295);
or UO_1132 (O_1132,N_15415,N_18413);
or UO_1133 (O_1133,N_17350,N_19838);
nand UO_1134 (O_1134,N_19110,N_15676);
and UO_1135 (O_1135,N_19460,N_16124);
or UO_1136 (O_1136,N_17804,N_16504);
and UO_1137 (O_1137,N_19208,N_18111);
and UO_1138 (O_1138,N_17081,N_15121);
or UO_1139 (O_1139,N_16412,N_19336);
nor UO_1140 (O_1140,N_16562,N_17176);
nor UO_1141 (O_1141,N_18301,N_16457);
and UO_1142 (O_1142,N_19041,N_16365);
nand UO_1143 (O_1143,N_18850,N_19827);
and UO_1144 (O_1144,N_16391,N_16389);
or UO_1145 (O_1145,N_19830,N_18989);
or UO_1146 (O_1146,N_15863,N_19682);
or UO_1147 (O_1147,N_18039,N_18434);
nand UO_1148 (O_1148,N_18610,N_19916);
xnor UO_1149 (O_1149,N_17604,N_18744);
or UO_1150 (O_1150,N_19748,N_16114);
nand UO_1151 (O_1151,N_16520,N_15915);
and UO_1152 (O_1152,N_16686,N_18247);
or UO_1153 (O_1153,N_17730,N_16794);
or UO_1154 (O_1154,N_18507,N_16080);
or UO_1155 (O_1155,N_17746,N_17882);
nand UO_1156 (O_1156,N_16746,N_16398);
nand UO_1157 (O_1157,N_15631,N_19816);
and UO_1158 (O_1158,N_19551,N_19250);
nand UO_1159 (O_1159,N_15023,N_16663);
and UO_1160 (O_1160,N_17070,N_16218);
nor UO_1161 (O_1161,N_16255,N_18436);
nor UO_1162 (O_1162,N_18235,N_16545);
or UO_1163 (O_1163,N_17657,N_18296);
and UO_1164 (O_1164,N_18047,N_18595);
nor UO_1165 (O_1165,N_15685,N_17404);
or UO_1166 (O_1166,N_18147,N_15050);
nand UO_1167 (O_1167,N_16599,N_17072);
nor UO_1168 (O_1168,N_16770,N_16448);
and UO_1169 (O_1169,N_18992,N_19143);
or UO_1170 (O_1170,N_19458,N_19740);
nor UO_1171 (O_1171,N_15519,N_17335);
and UO_1172 (O_1172,N_16463,N_19018);
and UO_1173 (O_1173,N_19231,N_15832);
and UO_1174 (O_1174,N_19524,N_17583);
and UO_1175 (O_1175,N_18573,N_19249);
or UO_1176 (O_1176,N_19703,N_18384);
nand UO_1177 (O_1177,N_16704,N_16722);
or UO_1178 (O_1178,N_15687,N_17789);
or UO_1179 (O_1179,N_18213,N_18478);
nand UO_1180 (O_1180,N_18545,N_18343);
nand UO_1181 (O_1181,N_17386,N_18066);
nor UO_1182 (O_1182,N_15390,N_17424);
xnor UO_1183 (O_1183,N_15166,N_19760);
and UO_1184 (O_1184,N_16147,N_15454);
nand UO_1185 (O_1185,N_15091,N_19163);
and UO_1186 (O_1186,N_19476,N_15882);
nor UO_1187 (O_1187,N_19755,N_19005);
nor UO_1188 (O_1188,N_19280,N_17792);
xnor UO_1189 (O_1189,N_15436,N_19049);
nor UO_1190 (O_1190,N_15289,N_19670);
and UO_1191 (O_1191,N_18099,N_15490);
nor UO_1192 (O_1192,N_19274,N_17360);
or UO_1193 (O_1193,N_17878,N_17349);
nand UO_1194 (O_1194,N_18194,N_15004);
or UO_1195 (O_1195,N_15184,N_16525);
and UO_1196 (O_1196,N_18681,N_17515);
nand UO_1197 (O_1197,N_17296,N_18995);
nor UO_1198 (O_1198,N_16166,N_19797);
nand UO_1199 (O_1199,N_15369,N_19745);
nor UO_1200 (O_1200,N_17714,N_17354);
or UO_1201 (O_1201,N_18471,N_17256);
nor UO_1202 (O_1202,N_18320,N_19789);
nor UO_1203 (O_1203,N_15776,N_18991);
or UO_1204 (O_1204,N_15902,N_18397);
and UO_1205 (O_1205,N_19441,N_17272);
nand UO_1206 (O_1206,N_18758,N_18734);
or UO_1207 (O_1207,N_16990,N_18277);
and UO_1208 (O_1208,N_15565,N_15825);
nand UO_1209 (O_1209,N_17293,N_19567);
or UO_1210 (O_1210,N_16948,N_18427);
nor UO_1211 (O_1211,N_17717,N_15695);
and UO_1212 (O_1212,N_16758,N_17340);
nor UO_1213 (O_1213,N_17805,N_16135);
or UO_1214 (O_1214,N_19792,N_15407);
nor UO_1215 (O_1215,N_15439,N_16814);
or UO_1216 (O_1216,N_15762,N_19996);
nand UO_1217 (O_1217,N_18512,N_15923);
or UO_1218 (O_1218,N_18918,N_17358);
or UO_1219 (O_1219,N_18021,N_15300);
nor UO_1220 (O_1220,N_18869,N_16331);
and UO_1221 (O_1221,N_15584,N_15965);
or UO_1222 (O_1222,N_15707,N_16942);
nor UO_1223 (O_1223,N_16651,N_17796);
and UO_1224 (O_1224,N_18380,N_16543);
and UO_1225 (O_1225,N_19902,N_17689);
nand UO_1226 (O_1226,N_18109,N_18849);
nand UO_1227 (O_1227,N_18927,N_17575);
nand UO_1228 (O_1228,N_18333,N_17521);
and UO_1229 (O_1229,N_16540,N_18452);
and UO_1230 (O_1230,N_15089,N_17853);
or UO_1231 (O_1231,N_18964,N_19982);
and UO_1232 (O_1232,N_16120,N_16576);
or UO_1233 (O_1233,N_15782,N_18847);
nor UO_1234 (O_1234,N_18492,N_17948);
or UO_1235 (O_1235,N_18352,N_19398);
or UO_1236 (O_1236,N_15826,N_17011);
nor UO_1237 (O_1237,N_16727,N_15950);
nor UO_1238 (O_1238,N_18271,N_18451);
nand UO_1239 (O_1239,N_17940,N_15799);
and UO_1240 (O_1240,N_17928,N_19331);
and UO_1241 (O_1241,N_16205,N_15202);
nor UO_1242 (O_1242,N_15911,N_19189);
or UO_1243 (O_1243,N_17269,N_16381);
nor UO_1244 (O_1244,N_15854,N_15419);
and UO_1245 (O_1245,N_18749,N_17958);
and UO_1246 (O_1246,N_17871,N_15272);
nand UO_1247 (O_1247,N_19981,N_17402);
nor UO_1248 (O_1248,N_15781,N_16202);
nor UO_1249 (O_1249,N_17181,N_16362);
and UO_1250 (O_1250,N_19244,N_17022);
nand UO_1251 (O_1251,N_18591,N_15514);
and UO_1252 (O_1252,N_16426,N_19435);
nor UO_1253 (O_1253,N_17555,N_15282);
or UO_1254 (O_1254,N_18489,N_15324);
nand UO_1255 (O_1255,N_16353,N_17658);
or UO_1256 (O_1256,N_16601,N_15061);
or UO_1257 (O_1257,N_16424,N_17161);
nor UO_1258 (O_1258,N_18313,N_17564);
nand UO_1259 (O_1259,N_19695,N_16013);
nand UO_1260 (O_1260,N_16480,N_16439);
nor UO_1261 (O_1261,N_15410,N_17071);
nor UO_1262 (O_1262,N_15576,N_18331);
nand UO_1263 (O_1263,N_18873,N_16095);
nor UO_1264 (O_1264,N_16001,N_19662);
and UO_1265 (O_1265,N_18181,N_18125);
nor UO_1266 (O_1266,N_19919,N_19176);
and UO_1267 (O_1267,N_19638,N_19892);
nand UO_1268 (O_1268,N_19263,N_18410);
or UO_1269 (O_1269,N_15320,N_18281);
nor UO_1270 (O_1270,N_19223,N_19136);
or UO_1271 (O_1271,N_16513,N_15258);
nor UO_1272 (O_1272,N_17153,N_15284);
and UO_1273 (O_1273,N_16810,N_18173);
and UO_1274 (O_1274,N_15714,N_15751);
nor UO_1275 (O_1275,N_16677,N_16314);
and UO_1276 (O_1276,N_17043,N_17415);
or UO_1277 (O_1277,N_18969,N_15958);
and UO_1278 (O_1278,N_17574,N_18790);
and UO_1279 (O_1279,N_18272,N_18444);
nand UO_1280 (O_1280,N_16931,N_15373);
or UO_1281 (O_1281,N_15084,N_16699);
or UO_1282 (O_1282,N_18759,N_18052);
or UO_1283 (O_1283,N_15329,N_17934);
nor UO_1284 (O_1284,N_19380,N_15049);
and UO_1285 (O_1285,N_16015,N_15563);
and UO_1286 (O_1286,N_19717,N_15111);
or UO_1287 (O_1287,N_17670,N_16105);
nand UO_1288 (O_1288,N_19431,N_18367);
nor UO_1289 (O_1289,N_18260,N_15721);
nor UO_1290 (O_1290,N_19473,N_19935);
nand UO_1291 (O_1291,N_17024,N_16884);
and UO_1292 (O_1292,N_18783,N_16613);
and UO_1293 (O_1293,N_16795,N_19194);
and UO_1294 (O_1294,N_17610,N_16225);
nand UO_1295 (O_1295,N_15571,N_17119);
nand UO_1296 (O_1296,N_19479,N_16952);
or UO_1297 (O_1297,N_17709,N_19180);
nand UO_1298 (O_1298,N_15368,N_18750);
nand UO_1299 (O_1299,N_15101,N_16321);
or UO_1300 (O_1300,N_16939,N_17044);
nand UO_1301 (O_1301,N_17996,N_18233);
or UO_1302 (O_1302,N_19878,N_17276);
and UO_1303 (O_1303,N_17227,N_15217);
or UO_1304 (O_1304,N_16585,N_18428);
and UO_1305 (O_1305,N_16392,N_16433);
and UO_1306 (O_1306,N_15534,N_15383);
nand UO_1307 (O_1307,N_19387,N_17103);
nand UO_1308 (O_1308,N_15759,N_16740);
or UO_1309 (O_1309,N_16136,N_19998);
nor UO_1310 (O_1310,N_19621,N_17037);
and UO_1311 (O_1311,N_18604,N_15551);
and UO_1312 (O_1312,N_18960,N_19600);
or UO_1313 (O_1313,N_16104,N_18922);
nor UO_1314 (O_1314,N_18044,N_15564);
nor UO_1315 (O_1315,N_17737,N_18968);
nand UO_1316 (O_1316,N_15555,N_19080);
xnor UO_1317 (O_1317,N_18791,N_16750);
and UO_1318 (O_1318,N_19715,N_17899);
nor UO_1319 (O_1319,N_17059,N_18226);
nor UO_1320 (O_1320,N_16475,N_18360);
nand UO_1321 (O_1321,N_15405,N_18087);
nor UO_1322 (O_1322,N_18379,N_15941);
or UO_1323 (O_1323,N_15796,N_16915);
nor UO_1324 (O_1324,N_15866,N_16116);
nor UO_1325 (O_1325,N_18536,N_18903);
and UO_1326 (O_1326,N_17165,N_18312);
nor UO_1327 (O_1327,N_15013,N_18354);
and UO_1328 (O_1328,N_16556,N_15313);
or UO_1329 (O_1329,N_19464,N_16968);
nand UO_1330 (O_1330,N_16419,N_19799);
and UO_1331 (O_1331,N_19109,N_16148);
and UO_1332 (O_1332,N_18497,N_15771);
and UO_1333 (O_1333,N_15604,N_15477);
and UO_1334 (O_1334,N_19832,N_19953);
nand UO_1335 (O_1335,N_16797,N_17831);
and UO_1336 (O_1336,N_16809,N_18988);
or UO_1337 (O_1337,N_17523,N_16140);
xor UO_1338 (O_1338,N_19179,N_15462);
nor UO_1339 (O_1339,N_19995,N_19137);
and UO_1340 (O_1340,N_15181,N_18438);
nand UO_1341 (O_1341,N_15433,N_15860);
nor UO_1342 (O_1342,N_17369,N_15700);
and UO_1343 (O_1343,N_19285,N_17089);
and UO_1344 (O_1344,N_18781,N_16928);
or UO_1345 (O_1345,N_17096,N_18375);
nor UO_1346 (O_1346,N_16813,N_17397);
or UO_1347 (O_1347,N_15073,N_16904);
or UO_1348 (O_1348,N_19084,N_15651);
and UO_1349 (O_1349,N_15385,N_19824);
and UO_1350 (O_1350,N_16269,N_19677);
and UO_1351 (O_1351,N_16064,N_19103);
or UO_1352 (O_1352,N_17586,N_15588);
and UO_1353 (O_1353,N_17672,N_16402);
nor UO_1354 (O_1354,N_15380,N_15570);
and UO_1355 (O_1355,N_18297,N_18897);
nand UO_1356 (O_1356,N_19844,N_18717);
nor UO_1357 (O_1357,N_17483,N_18778);
and UO_1358 (O_1358,N_18491,N_17563);
and UO_1359 (O_1359,N_16575,N_18458);
and UO_1360 (O_1360,N_18137,N_16664);
or UO_1361 (O_1361,N_17833,N_19365);
and UO_1362 (O_1362,N_18270,N_15063);
nor UO_1363 (O_1363,N_16347,N_19360);
nand UO_1364 (O_1364,N_18543,N_19227);
and UO_1365 (O_1365,N_16260,N_17261);
nand UO_1366 (O_1366,N_16387,N_19989);
and UO_1367 (O_1367,N_15158,N_19484);
and UO_1368 (O_1368,N_19425,N_19369);
and UO_1369 (O_1369,N_17502,N_15655);
or UO_1370 (O_1370,N_19671,N_15161);
nand UO_1371 (O_1371,N_17445,N_19924);
or UO_1372 (O_1372,N_17697,N_15591);
or UO_1373 (O_1373,N_17873,N_16115);
nand UO_1374 (O_1374,N_16043,N_16042);
nand UO_1375 (O_1375,N_16697,N_15594);
nor UO_1376 (O_1376,N_17135,N_19650);
nor UO_1377 (O_1377,N_15745,N_19375);
nand UO_1378 (O_1378,N_18238,N_17393);
nand UO_1379 (O_1379,N_15311,N_18867);
and UO_1380 (O_1380,N_16453,N_16541);
and UO_1381 (O_1381,N_15425,N_16633);
or UO_1382 (O_1382,N_18649,N_18851);
nand UO_1383 (O_1383,N_19088,N_19541);
nor UO_1384 (O_1384,N_17325,N_18349);
nand UO_1385 (O_1385,N_17642,N_16680);
and UO_1386 (O_1386,N_16499,N_17625);
nor UO_1387 (O_1387,N_15876,N_15640);
or UO_1388 (O_1388,N_19125,N_18366);
nor UO_1389 (O_1389,N_16671,N_17595);
and UO_1390 (O_1390,N_19038,N_19532);
and UO_1391 (O_1391,N_19396,N_16204);
or UO_1392 (O_1392,N_17101,N_19722);
nand UO_1393 (O_1393,N_16845,N_15367);
and UO_1394 (O_1394,N_19870,N_16249);
nor UO_1395 (O_1395,N_15005,N_16173);
xor UO_1396 (O_1396,N_16134,N_18447);
and UO_1397 (O_1397,N_16144,N_17851);
and UO_1398 (O_1398,N_18429,N_17983);
and UO_1399 (O_1399,N_15509,N_18876);
nor UO_1400 (O_1400,N_16866,N_16850);
or UO_1401 (O_1401,N_15960,N_18321);
or UO_1402 (O_1402,N_16706,N_18633);
or UO_1403 (O_1403,N_16649,N_15382);
nand UO_1404 (O_1404,N_18748,N_19389);
nand UO_1405 (O_1405,N_18925,N_18395);
nor UO_1406 (O_1406,N_15659,N_15306);
and UO_1407 (O_1407,N_18924,N_17718);
nor UO_1408 (O_1408,N_19196,N_19323);
or UO_1409 (O_1409,N_15237,N_19296);
or UO_1410 (O_1410,N_17793,N_15744);
nand UO_1411 (O_1411,N_18716,N_16366);
or UO_1412 (O_1412,N_19017,N_15868);
nor UO_1413 (O_1413,N_16979,N_16519);
or UO_1414 (O_1414,N_15444,N_16315);
nand UO_1415 (O_1415,N_15497,N_16425);
or UO_1416 (O_1416,N_19306,N_17883);
xnor UO_1417 (O_1417,N_16174,N_16868);
or UO_1418 (O_1418,N_19972,N_16609);
or UO_1419 (O_1419,N_15770,N_18426);
nor UO_1420 (O_1420,N_18318,N_19295);
and UO_1421 (O_1421,N_15336,N_18656);
and UO_1422 (O_1422,N_17526,N_16564);
nor UO_1423 (O_1423,N_19315,N_19825);
nand UO_1424 (O_1424,N_16878,N_18987);
or UO_1425 (O_1425,N_19200,N_15480);
nor UO_1426 (O_1426,N_18023,N_19377);
nor UO_1427 (O_1427,N_16739,N_15636);
and UO_1428 (O_1428,N_15213,N_16003);
nor UO_1429 (O_1429,N_16847,N_18614);
or UO_1430 (O_1430,N_19287,N_16798);
nand UO_1431 (O_1431,N_15100,N_17576);
or UO_1432 (O_1432,N_19023,N_15189);
nor UO_1433 (O_1433,N_15295,N_15353);
nand UO_1434 (O_1434,N_19618,N_15174);
or UO_1435 (O_1435,N_17237,N_17845);
nor UO_1436 (O_1436,N_16547,N_19308);
and UO_1437 (O_1437,N_16360,N_16734);
and UO_1438 (O_1438,N_16618,N_16551);
nor UO_1439 (O_1439,N_15630,N_16927);
nand UO_1440 (O_1440,N_18388,N_16675);
and UO_1441 (O_1441,N_17991,N_16612);
and UO_1442 (O_1442,N_18140,N_15635);
nor UO_1443 (O_1443,N_15686,N_19559);
nand UO_1444 (O_1444,N_16092,N_19115);
nand UO_1445 (O_1445,N_17626,N_19889);
nand UO_1446 (O_1446,N_17446,N_15801);
or UO_1447 (O_1447,N_18289,N_15256);
nand UO_1448 (O_1448,N_16441,N_15430);
and UO_1449 (O_1449,N_16338,N_16081);
nor UO_1450 (O_1450,N_18196,N_16542);
nand UO_1451 (O_1451,N_17303,N_17788);
xnor UO_1452 (O_1452,N_19076,N_19651);
xor UO_1453 (O_1453,N_19478,N_17762);
or UO_1454 (O_1454,N_18074,N_19317);
nand UO_1455 (O_1455,N_18041,N_16297);
and UO_1456 (O_1456,N_18839,N_17569);
or UO_1457 (O_1457,N_16051,N_17451);
nor UO_1458 (O_1458,N_19469,N_15835);
or UO_1459 (O_1459,N_16145,N_19062);
nor UO_1460 (O_1460,N_16590,N_17183);
and UO_1461 (O_1461,N_15807,N_19305);
or UO_1462 (O_1462,N_16244,N_19434);
nor UO_1463 (O_1463,N_15175,N_18701);
and UO_1464 (O_1464,N_18334,N_16786);
nor UO_1465 (O_1465,N_17137,N_19020);
or UO_1466 (O_1466,N_19921,N_18498);
nand UO_1467 (O_1467,N_18273,N_17210);
or UO_1468 (O_1468,N_17655,N_16997);
nor UO_1469 (O_1469,N_15608,N_17632);
and UO_1470 (O_1470,N_16241,N_16358);
and UO_1471 (O_1471,N_16110,N_19779);
xor UO_1472 (O_1472,N_17906,N_19514);
or UO_1473 (O_1473,N_16496,N_16193);
nor UO_1474 (O_1474,N_16132,N_18732);
and UO_1475 (O_1475,N_18975,N_16529);
nand UO_1476 (O_1476,N_18773,N_18694);
nor UO_1477 (O_1477,N_17876,N_19664);
and UO_1478 (O_1478,N_17613,N_17903);
nand UO_1479 (O_1479,N_15176,N_16479);
or UO_1480 (O_1480,N_19547,N_18886);
and UO_1481 (O_1481,N_18290,N_18042);
nor UO_1482 (O_1482,N_15539,N_18088);
nor UO_1483 (O_1483,N_18348,N_19492);
nor UO_1484 (O_1484,N_19256,N_16628);
and UO_1485 (O_1485,N_15463,N_19527);
and UO_1486 (O_1486,N_17849,N_19578);
or UO_1487 (O_1487,N_18793,N_18568);
nor UO_1488 (O_1488,N_17993,N_17485);
or UO_1489 (O_1489,N_19490,N_15733);
and UO_1490 (O_1490,N_18693,N_19105);
nand UO_1491 (O_1491,N_15775,N_18747);
or UO_1492 (O_1492,N_15738,N_19181);
or UO_1493 (O_1493,N_15179,N_18508);
nor UO_1494 (O_1494,N_15216,N_19750);
and UO_1495 (O_1495,N_15059,N_17039);
nand UO_1496 (O_1496,N_16437,N_18250);
or UO_1497 (O_1497,N_18155,N_15156);
nor UO_1498 (O_1498,N_19658,N_17420);
and UO_1499 (O_1499,N_18229,N_16785);
or UO_1500 (O_1500,N_16063,N_19248);
and UO_1501 (O_1501,N_19228,N_17250);
nand UO_1502 (O_1502,N_18132,N_16259);
nor UO_1503 (O_1503,N_18028,N_15627);
and UO_1504 (O_1504,N_19423,N_16676);
or UO_1505 (O_1505,N_18164,N_19428);
nor UO_1506 (O_1506,N_16232,N_15784);
or UO_1507 (O_1507,N_17680,N_16491);
nand UO_1508 (O_1508,N_17414,N_19588);
nand UO_1509 (O_1509,N_19973,N_18449);
and UO_1510 (O_1510,N_17281,N_17514);
or UO_1511 (O_1511,N_18101,N_17795);
nand UO_1512 (O_1512,N_16084,N_17159);
nand UO_1513 (O_1513,N_16333,N_18154);
nand UO_1514 (O_1514,N_16343,N_19496);
and UO_1515 (O_1515,N_15559,N_18358);
nand UO_1516 (O_1516,N_15342,N_18626);
and UO_1517 (O_1517,N_15493,N_16645);
and UO_1518 (O_1518,N_16857,N_19447);
nor UO_1519 (O_1519,N_17063,N_16698);
or UO_1520 (O_1520,N_16010,N_15236);
and UO_1521 (O_1521,N_18402,N_18187);
and UO_1522 (O_1522,N_16848,N_18058);
or UO_1523 (O_1523,N_15601,N_15850);
or UO_1524 (O_1524,N_17890,N_17289);
and UO_1525 (O_1525,N_19978,N_19293);
and UO_1526 (O_1526,N_17922,N_19809);
nor UO_1527 (O_1527,N_18718,N_16642);
nand UO_1528 (O_1528,N_18242,N_17892);
nand UO_1529 (O_1529,N_16988,N_18529);
and UO_1530 (O_1530,N_15109,N_18060);
and UO_1531 (O_1531,N_16196,N_17782);
nand UO_1532 (O_1532,N_16184,N_17900);
or UO_1533 (O_1533,N_19354,N_19127);
nand UO_1534 (O_1534,N_16054,N_19051);
nor UO_1535 (O_1535,N_17755,N_18779);
nor UO_1536 (O_1536,N_19866,N_19851);
nand UO_1537 (O_1537,N_16714,N_19310);
nor UO_1538 (O_1538,N_17615,N_17663);
nor UO_1539 (O_1539,N_18917,N_18774);
or UO_1540 (O_1540,N_16178,N_17491);
or UO_1541 (O_1541,N_19311,N_17591);
or UO_1542 (O_1542,N_16956,N_18390);
nand UO_1543 (O_1543,N_15881,N_17034);
nand UO_1544 (O_1544,N_19776,N_16363);
nor UO_1545 (O_1545,N_18896,N_18165);
and UO_1546 (O_1546,N_16862,N_18359);
nor UO_1547 (O_1547,N_15144,N_16170);
nand UO_1548 (O_1548,N_16228,N_15424);
nor UO_1549 (O_1549,N_19560,N_17368);
nor UO_1550 (O_1550,N_19032,N_18198);
nor UO_1551 (O_1551,N_18433,N_15725);
and UO_1552 (O_1552,N_19245,N_17597);
nand UO_1553 (O_1553,N_19920,N_16374);
nor UO_1554 (O_1554,N_17643,N_17311);
nand UO_1555 (O_1555,N_16151,N_18516);
nand UO_1556 (O_1556,N_16565,N_18210);
or UO_1557 (O_1557,N_18899,N_15253);
nand UO_1558 (O_1558,N_15856,N_17407);
nand UO_1559 (O_1559,N_15894,N_17609);
and UO_1560 (O_1560,N_19927,N_19746);
or UO_1561 (O_1561,N_16818,N_18329);
nand UO_1562 (O_1562,N_18558,N_17728);
and UO_1563 (O_1563,N_19633,N_15095);
or UO_1564 (O_1564,N_18437,N_16413);
nand UO_1565 (O_1565,N_17476,N_17946);
and UO_1566 (O_1566,N_16430,N_18330);
nor UO_1567 (O_1567,N_15248,N_17252);
nand UO_1568 (O_1568,N_18696,N_17170);
nor UO_1569 (O_1569,N_18197,N_16687);
nand UO_1570 (O_1570,N_17098,N_18862);
nor UO_1571 (O_1571,N_19152,N_19030);
or UO_1572 (O_1572,N_19512,N_19754);
nor UO_1573 (O_1573,N_15945,N_18589);
nor UO_1574 (O_1574,N_17019,N_19576);
nor UO_1575 (O_1575,N_18594,N_17607);
and UO_1576 (O_1576,N_15455,N_18659);
nor UO_1577 (O_1577,N_17363,N_16837);
nand UO_1578 (O_1578,N_17757,N_17337);
or UO_1579 (O_1579,N_18926,N_19001);
or UO_1580 (O_1580,N_17517,N_18745);
nand UO_1581 (O_1581,N_16235,N_18895);
and UO_1582 (O_1582,N_19957,N_19912);
or UO_1583 (O_1583,N_18684,N_18637);
nor UO_1584 (O_1584,N_19374,N_19135);
or UO_1585 (O_1585,N_19643,N_18282);
or UO_1586 (O_1586,N_16668,N_15760);
and UO_1587 (O_1587,N_16253,N_15193);
nand UO_1588 (O_1588,N_16462,N_15076);
and UO_1589 (O_1589,N_18691,N_15891);
nand UO_1590 (O_1590,N_18288,N_19602);
or UO_1591 (O_1591,N_18978,N_18025);
or UO_1592 (O_1592,N_18821,N_16532);
nor UO_1593 (O_1593,N_19737,N_19821);
nand UO_1594 (O_1594,N_18425,N_19099);
and UO_1595 (O_1595,N_19167,N_16623);
or UO_1596 (O_1596,N_17865,N_15634);
nand UO_1597 (O_1597,N_16583,N_19865);
nor UO_1598 (O_1598,N_18670,N_16005);
or UO_1599 (O_1599,N_17651,N_16342);
or UO_1600 (O_1600,N_18767,N_17719);
nor UO_1601 (O_1601,N_19173,N_18804);
nor UO_1602 (O_1602,N_18114,N_19840);
and UO_1603 (O_1603,N_17531,N_15848);
nand UO_1604 (O_1604,N_19887,N_18049);
nor UO_1605 (O_1605,N_18221,N_19674);
nand UO_1606 (O_1606,N_17417,N_17683);
or UO_1607 (O_1607,N_18422,N_17599);
nor UO_1608 (O_1608,N_19102,N_19648);
nor UO_1609 (O_1609,N_15322,N_19687);
and UO_1610 (O_1610,N_16312,N_15864);
xnor UO_1611 (O_1611,N_16066,N_18825);
or UO_1612 (O_1612,N_19681,N_18254);
nand UO_1613 (O_1613,N_17216,N_19443);
and UO_1614 (O_1614,N_17593,N_17629);
nor UO_1615 (O_1615,N_15907,N_15305);
and UO_1616 (O_1616,N_19268,N_18826);
nand UO_1617 (O_1617,N_15071,N_18249);
nand UO_1618 (O_1618,N_16478,N_19806);
or UO_1619 (O_1619,N_17267,N_19415);
and UO_1620 (O_1620,N_17808,N_18712);
or UO_1621 (O_1621,N_16521,N_18361);
nand UO_1622 (O_1622,N_17971,N_19626);
and UO_1623 (O_1623,N_17581,N_17560);
nor UO_1624 (O_1624,N_16023,N_18945);
or UO_1625 (O_1625,N_17482,N_16019);
and UO_1626 (O_1626,N_18309,N_16872);
nor UO_1627 (O_1627,N_18248,N_15680);
nand UO_1628 (O_1628,N_17245,N_16029);
nor UO_1629 (O_1629,N_16201,N_16924);
and UO_1630 (O_1630,N_19101,N_15008);
nor UO_1631 (O_1631,N_16606,N_17205);
and UO_1632 (O_1632,N_17292,N_15849);
nand UO_1633 (O_1633,N_17918,N_18401);
nor UO_1634 (O_1634,N_15912,N_15129);
and UO_1635 (O_1635,N_17062,N_16336);
and UO_1636 (O_1636,N_18373,N_19704);
nand UO_1637 (O_1637,N_17565,N_17457);
or UO_1638 (O_1638,N_18110,N_19857);
nor UO_1639 (O_1639,N_17005,N_17080);
nor UO_1640 (O_1640,N_16940,N_19980);
nor UO_1641 (O_1641,N_18480,N_18966);
nor UO_1642 (O_1642,N_15223,N_16213);
nor UO_1643 (O_1643,N_19009,N_15566);
nand UO_1644 (O_1644,N_17916,N_16829);
or UO_1645 (O_1645,N_15200,N_16431);
and UO_1646 (O_1646,N_18029,N_16626);
and UO_1647 (O_1647,N_17160,N_17122);
nor UO_1648 (O_1648,N_19518,N_19531);
or UO_1649 (O_1649,N_19845,N_15645);
nand UO_1650 (O_1650,N_17803,N_19752);
or UO_1651 (O_1651,N_17622,N_15485);
or UO_1652 (O_1652,N_15938,N_17998);
or UO_1653 (O_1653,N_17112,N_18946);
nand UO_1654 (O_1654,N_15644,N_16910);
nand UO_1655 (O_1655,N_17466,N_18775);
xor UO_1656 (O_1656,N_17784,N_18371);
nor UO_1657 (O_1657,N_19706,N_19977);
nor UO_1658 (O_1658,N_15183,N_19344);
or UO_1659 (O_1659,N_19822,N_19680);
or UO_1660 (O_1660,N_17914,N_17620);
or UO_1661 (O_1661,N_16763,N_19790);
nor UO_1662 (O_1662,N_16162,N_17506);
nor UO_1663 (O_1663,N_16111,N_15447);
or UO_1664 (O_1664,N_15360,N_16580);
nand UO_1665 (O_1665,N_17619,N_17042);
nand UO_1666 (O_1666,N_16702,N_17129);
and UO_1667 (O_1667,N_16527,N_15075);
and UO_1668 (O_1668,N_19465,N_17679);
xor UO_1669 (O_1669,N_16368,N_19214);
nand UO_1670 (O_1670,N_15639,N_18764);
nand UO_1671 (O_1671,N_17113,N_15378);
nand UO_1672 (O_1672,N_16183,N_19430);
and UO_1673 (O_1673,N_16476,N_19505);
and UO_1674 (O_1674,N_19302,N_17534);
nor UO_1675 (O_1675,N_16652,N_15836);
and UO_1676 (O_1676,N_19882,N_19239);
nor UO_1677 (O_1677,N_15903,N_19070);
nor UO_1678 (O_1678,N_16016,N_15475);
or UO_1679 (O_1679,N_18185,N_18761);
nand UO_1680 (O_1680,N_18421,N_17942);
and UO_1681 (O_1681,N_16456,N_16383);
nand UO_1682 (O_1682,N_15944,N_19094);
nand UO_1683 (O_1683,N_17035,N_16566);
and UO_1684 (O_1684,N_17058,N_18763);
nand UO_1685 (O_1685,N_15793,N_17025);
and UO_1686 (O_1686,N_18721,N_19736);
or UO_1687 (O_1687,N_17713,N_18798);
and UO_1688 (O_1688,N_18782,N_17999);
and UO_1689 (O_1689,N_16741,N_17970);
nor UO_1690 (O_1690,N_16674,N_17115);
nand UO_1691 (O_1691,N_16945,N_15511);
nor UO_1692 (O_1692,N_15355,N_18228);
and UO_1693 (O_1693,N_15440,N_17703);
or UO_1694 (O_1694,N_17026,N_16552);
or UO_1695 (O_1695,N_16048,N_18768);
and UO_1696 (O_1696,N_18832,N_19368);
nand UO_1697 (O_1697,N_16641,N_16710);
nand UO_1698 (O_1698,N_15688,N_19702);
nand UO_1699 (O_1699,N_17590,N_17134);
and UO_1700 (O_1700,N_19325,N_17422);
or UO_1701 (O_1701,N_17963,N_19362);
nand UO_1702 (O_1702,N_17346,N_15465);
nor UO_1703 (O_1703,N_16443,N_19762);
or UO_1704 (O_1704,N_15445,N_16922);
nand UO_1705 (O_1705,N_16792,N_16058);
nor UO_1706 (O_1706,N_18473,N_16226);
nor UO_1707 (O_1707,N_15827,N_16418);
and UO_1708 (O_1708,N_17460,N_19511);
nor UO_1709 (O_1709,N_18341,N_19798);
and UO_1710 (O_1710,N_19646,N_18439);
and UO_1711 (O_1711,N_16071,N_18570);
nor UO_1712 (O_1712,N_15274,N_16390);
nand UO_1713 (O_1713,N_18416,N_19329);
nand UO_1714 (O_1714,N_18307,N_18817);
nor UO_1715 (O_1715,N_19791,N_18383);
and UO_1716 (O_1716,N_16584,N_15215);
or UO_1717 (O_1717,N_17536,N_17550);
nor UO_1718 (O_1718,N_16995,N_19690);
or UO_1719 (O_1719,N_15182,N_15496);
nand UO_1720 (O_1720,N_19154,N_16764);
or UO_1721 (O_1721,N_18003,N_16644);
nand UO_1722 (O_1722,N_16759,N_18004);
and UO_1723 (O_1723,N_15154,N_17956);
or UO_1724 (O_1724,N_18807,N_16842);
or UO_1725 (O_1725,N_18827,N_15038);
xor UO_1726 (O_1726,N_18981,N_17236);
and UO_1727 (O_1727,N_16401,N_18323);
nand UO_1728 (O_1728,N_19817,N_18339);
or UO_1729 (O_1729,N_17968,N_15108);
nor UO_1730 (O_1730,N_18556,N_19554);
nor UO_1731 (O_1731,N_15577,N_19634);
and UO_1732 (O_1732,N_18476,N_17032);
nand UO_1733 (O_1733,N_15428,N_15988);
nor UO_1734 (O_1734,N_18474,N_15102);
or UO_1735 (O_1735,N_18729,N_17240);
or UO_1736 (O_1736,N_18731,N_18256);
or UO_1737 (O_1737,N_18189,N_15009);
or UO_1738 (O_1738,N_17207,N_16395);
nor UO_1739 (O_1739,N_16683,N_16934);
nor UO_1740 (O_1740,N_17158,N_18676);
nand UO_1741 (O_1741,N_17083,N_19908);
or UO_1742 (O_1742,N_17635,N_17280);
nor UO_1743 (O_1743,N_19012,N_15758);
and UO_1744 (O_1744,N_18398,N_16155);
and UO_1745 (O_1745,N_15769,N_19852);
nor UO_1746 (O_1746,N_18139,N_15427);
nand UO_1747 (O_1747,N_17154,N_15740);
nor UO_1748 (O_1748,N_15934,N_17197);
nor UO_1749 (O_1749,N_18382,N_18151);
nor UO_1750 (O_1750,N_17492,N_19419);
and UO_1751 (O_1751,N_16989,N_17474);
and UO_1752 (O_1752,N_19288,N_19714);
nor UO_1753 (O_1753,N_17056,N_19847);
nand UO_1754 (O_1754,N_16404,N_16421);
nand UO_1755 (O_1755,N_19481,N_19132);
and UO_1756 (O_1756,N_19692,N_19985);
nor UO_1757 (O_1757,N_16985,N_19391);
or UO_1758 (O_1758,N_19823,N_15756);
nor UO_1759 (O_1759,N_16748,N_17242);
and UO_1760 (O_1760,N_18816,N_18460);
nor UO_1761 (O_1761,N_17301,N_15269);
or UO_1762 (O_1762,N_15498,N_16720);
or UO_1763 (O_1763,N_19399,N_19184);
nand UO_1764 (O_1764,N_19016,N_15094);
nor UO_1765 (O_1765,N_19371,N_17057);
or UO_1766 (O_1766,N_18338,N_16964);
or UO_1767 (O_1767,N_16902,N_19165);
nor UO_1768 (O_1768,N_17623,N_18651);
or UO_1769 (O_1769,N_18581,N_19952);
or UO_1770 (O_1770,N_15741,N_17082);
nand UO_1771 (O_1771,N_15804,N_18572);
or UO_1772 (O_1772,N_15822,N_15837);
nand UO_1773 (O_1773,N_16078,N_17897);
and UO_1774 (O_1774,N_18215,N_15442);
nor UO_1775 (O_1775,N_16611,N_16586);
or UO_1776 (O_1776,N_17912,N_17552);
nor UO_1777 (O_1777,N_17367,N_17464);
and UO_1778 (O_1778,N_19938,N_18679);
nor UO_1779 (O_1779,N_15884,N_17200);
and UO_1780 (O_1780,N_16925,N_15581);
nand UO_1781 (O_1781,N_17891,N_17547);
or UO_1782 (O_1782,N_15890,N_18251);
or UO_1783 (O_1783,N_17823,N_19672);
nand UO_1784 (O_1784,N_16446,N_18129);
or UO_1785 (O_1785,N_18542,N_17225);
or UO_1786 (O_1786,N_19456,N_18722);
nor UO_1787 (O_1787,N_18236,N_17428);
xnor UO_1788 (O_1788,N_16650,N_19162);
nor UO_1789 (O_1789,N_17901,N_19159);
nand UO_1790 (O_1790,N_19471,N_16150);
nor UO_1791 (O_1791,N_19803,N_19855);
nand UO_1792 (O_1792,N_15178,N_16538);
nor UO_1793 (O_1793,N_19753,N_17213);
nand UO_1794 (O_1794,N_16638,N_15128);
nor UO_1795 (O_1795,N_15240,N_15983);
and UO_1796 (O_1796,N_16971,N_17733);
or UO_1797 (O_1797,N_18860,N_15472);
or UO_1798 (O_1798,N_17923,N_17073);
nand UO_1799 (O_1799,N_15040,N_19003);
nor UO_1800 (O_1800,N_17141,N_18941);
or UO_1801 (O_1801,N_18287,N_16229);
or UO_1802 (O_1802,N_16471,N_19444);
nor UO_1803 (O_1803,N_19156,N_16061);
nand UO_1804 (O_1804,N_18304,N_16854);
and UO_1805 (O_1805,N_18389,N_19608);
nand UO_1806 (O_1806,N_15556,N_17711);
or UO_1807 (O_1807,N_16438,N_18009);
or UO_1808 (O_1808,N_18980,N_15489);
and UO_1809 (O_1809,N_16373,N_15230);
nor UO_1810 (O_1810,N_19314,N_17262);
and UO_1811 (O_1811,N_16367,N_17185);
or UO_1812 (O_1812,N_16796,N_19033);
nor UO_1813 (O_1813,N_16455,N_19489);
and UO_1814 (O_1814,N_15906,N_19665);
nor UO_1815 (O_1815,N_17364,N_17195);
or UO_1816 (O_1816,N_19243,N_17665);
nor UO_1817 (O_1817,N_18275,N_19035);
or UO_1818 (O_1818,N_19085,N_15633);
and UO_1819 (O_1819,N_19558,N_16897);
or UO_1820 (O_1820,N_16625,N_18316);
and UO_1821 (O_1821,N_17774,N_19951);
nor UO_1822 (O_1822,N_16470,N_17734);
and UO_1823 (O_1823,N_19503,N_19267);
nor UO_1824 (O_1824,N_19128,N_19420);
and UO_1825 (O_1825,N_19673,N_19771);
nand UO_1826 (O_1826,N_19509,N_16186);
nor UO_1827 (O_1827,N_15561,N_15507);
or UO_1828 (O_1828,N_15169,N_18909);
and UO_1829 (O_1829,N_19529,N_18690);
or UO_1830 (O_1830,N_15323,N_16191);
and UO_1831 (O_1831,N_15196,N_15614);
nor UO_1832 (O_1832,N_16236,N_19929);
and UO_1833 (O_1833,N_15573,N_18602);
nor UO_1834 (O_1834,N_19801,N_17931);
or UO_1835 (O_1835,N_18822,N_15501);
nand UO_1836 (O_1836,N_17837,N_19262);
and UO_1837 (O_1837,N_16037,N_16411);
or UO_1838 (O_1838,N_19000,N_16757);
or UO_1839 (O_1839,N_16707,N_18754);
nand UO_1840 (O_1840,N_18363,N_16858);
and UO_1841 (O_1841,N_17333,N_18020);
and UO_1842 (O_1842,N_16180,N_19767);
nor UO_1843 (O_1843,N_15531,N_18751);
or UO_1844 (O_1844,N_16673,N_16885);
and UO_1845 (O_1845,N_15893,N_15859);
and UO_1846 (O_1846,N_15932,N_15515);
and UO_1847 (O_1847,N_18561,N_19230);
and UO_1848 (O_1848,N_16624,N_19400);
and UO_1849 (O_1849,N_16745,N_18796);
or UO_1850 (O_1850,N_19210,N_16006);
or UO_1851 (O_1851,N_16046,N_16415);
or UO_1852 (O_1852,N_15816,N_19079);
or UO_1853 (O_1853,N_19057,N_16161);
nand UO_1854 (O_1854,N_17442,N_16055);
and UO_1855 (O_1855,N_19300,N_16181);
nand UO_1856 (O_1856,N_15979,N_17498);
and UO_1857 (O_1857,N_19442,N_17529);
nor UO_1858 (O_1858,N_18928,N_18005);
nand UO_1859 (O_1859,N_18143,N_16406);
xnor UO_1860 (O_1860,N_15831,N_16537);
or UO_1861 (O_1861,N_19867,N_17486);
nor UO_1862 (O_1862,N_19666,N_16983);
nand UO_1863 (O_1863,N_17671,N_19282);
nand UO_1864 (O_1864,N_19361,N_17233);
or UO_1865 (O_1865,N_17542,N_19402);
and UO_1866 (O_1866,N_19853,N_19394);
and UO_1867 (O_1867,N_16427,N_17381);
nand UO_1868 (O_1868,N_17018,N_18996);
or UO_1869 (O_1869,N_19860,N_19940);
nor UO_1870 (O_1870,N_17495,N_16859);
and UO_1871 (O_1871,N_16976,N_15706);
or UO_1872 (O_1872,N_15186,N_16487);
or UO_1873 (O_1873,N_16946,N_16778);
nor UO_1874 (O_1874,N_15709,N_19133);
nand UO_1875 (O_1875,N_19694,N_18012);
nand UO_1876 (O_1876,N_17750,N_18093);
nor UO_1877 (O_1877,N_16873,N_16608);
nand UO_1878 (O_1878,N_16265,N_15168);
or UO_1879 (O_1879,N_16981,N_18086);
nor UO_1880 (O_1880,N_15310,N_19661);
or UO_1881 (O_1881,N_18985,N_17209);
nand UO_1882 (O_1882,N_15068,N_17829);
and UO_1883 (O_1883,N_15629,N_19656);
or UO_1884 (O_1884,N_18245,N_17637);
nand UO_1885 (O_1885,N_18819,N_17188);
and UO_1886 (O_1886,N_17178,N_17389);
and UO_1887 (O_1887,N_16639,N_15162);
nand UO_1888 (O_1888,N_16912,N_16800);
nor UO_1889 (O_1889,N_17395,N_15897);
and UO_1890 (O_1890,N_15245,N_19983);
xnor UO_1891 (O_1891,N_17321,N_17910);
nand UO_1892 (O_1892,N_19583,N_15930);
nand UO_1893 (O_1893,N_18934,N_15338);
nand UO_1894 (O_1894,N_15823,N_15221);
xnor UO_1895 (O_1895,N_17994,N_19905);
nand UO_1896 (O_1896,N_16090,N_16068);
and UO_1897 (O_1897,N_18124,N_17562);
or UO_1898 (O_1898,N_16049,N_17479);
nand UO_1899 (O_1899,N_16788,N_17444);
or UO_1900 (O_1900,N_19074,N_15187);
or UO_1901 (O_1901,N_18880,N_15291);
nor UO_1902 (O_1902,N_17171,N_18961);
and UO_1903 (O_1903,N_17953,N_16077);
and UO_1904 (O_1904,N_18617,N_18448);
or UO_1905 (O_1905,N_16949,N_19696);
nor UO_1906 (O_1906,N_15133,N_18657);
and UO_1907 (O_1907,N_15110,N_17111);
nor UO_1908 (O_1908,N_16158,N_17646);
or UO_1909 (O_1909,N_15975,N_18714);
or UO_1910 (O_1910,N_18202,N_19341);
or UO_1911 (O_1911,N_18015,N_19251);
and UO_1912 (O_1912,N_17163,N_19069);
nor UO_1913 (O_1913,N_15616,N_19327);
nor UO_1914 (O_1914,N_18566,N_18911);
nand UO_1915 (O_1915,N_16577,N_15654);
nand UO_1916 (O_1916,N_15443,N_18959);
or UO_1917 (O_1917,N_15045,N_19937);
or UO_1918 (O_1918,N_18138,N_16469);
nor UO_1919 (O_1919,N_19472,N_18590);
and UO_1920 (O_1920,N_15870,N_16718);
and UO_1921 (O_1921,N_19450,N_16167);
or UO_1922 (O_1922,N_19278,N_19584);
nand UO_1923 (O_1923,N_15623,N_18534);
and UO_1924 (O_1924,N_16622,N_18689);
and UO_1925 (O_1925,N_15729,N_16088);
nand UO_1926 (O_1926,N_18116,N_16422);
nor UO_1927 (O_1927,N_18073,N_16688);
or UO_1928 (O_1928,N_17490,N_19378);
and UO_1929 (O_1929,N_17780,N_15363);
nand UO_1930 (O_1930,N_15384,N_18806);
and UO_1931 (O_1931,N_19226,N_17102);
nand UO_1932 (O_1932,N_18524,N_17298);
nor UO_1933 (O_1933,N_17156,N_18654);
and UO_1934 (O_1934,N_19636,N_19345);
nand UO_1935 (O_1935,N_15535,N_16775);
and UO_1936 (O_1936,N_17690,N_19993);
or UO_1937 (O_1937,N_15698,N_16429);
nor UO_1938 (O_1938,N_19134,N_15090);
and UO_1939 (O_1939,N_17429,N_16762);
and UO_1940 (O_1940,N_19592,N_15670);
nor UO_1941 (O_1941,N_17138,N_16805);
nand UO_1942 (O_1942,N_19770,N_16860);
or UO_1943 (O_1943,N_16279,N_17541);
nand UO_1944 (O_1944,N_16558,N_16481);
or UO_1945 (O_1945,N_19356,N_19410);
nand UO_1946 (O_1946,N_19868,N_15795);
nor UO_1947 (O_1947,N_18405,N_15746);
and UO_1948 (O_1948,N_18688,N_15304);
and UO_1949 (O_1949,N_18424,N_15268);
nand UO_1950 (O_1950,N_18937,N_18144);
and UO_1951 (O_1951,N_19312,N_16165);
and UO_1952 (O_1952,N_15711,N_19131);
nand UO_1953 (O_1953,N_17747,N_17078);
nand UO_1954 (O_1954,N_16602,N_16277);
and UO_1955 (O_1955,N_19252,N_18852);
or UO_1956 (O_1956,N_18963,N_18211);
nor UO_1957 (O_1957,N_15516,N_15404);
nand UO_1958 (O_1958,N_15487,N_16492);
xor UO_1959 (O_1959,N_19970,N_19881);
and UO_1960 (O_1960,N_15393,N_19599);
or UO_1961 (O_1961,N_19355,N_16093);
and UO_1962 (O_1962,N_15157,N_19113);
or UO_1963 (O_1963,N_19979,N_17791);
nand UO_1964 (O_1964,N_17302,N_19861);
nand UO_1965 (O_1965,N_19366,N_16893);
nand UO_1966 (O_1966,N_19676,N_19275);
and UO_1967 (O_1967,N_15933,N_17744);
and UO_1968 (O_1968,N_16731,N_16408);
nor UO_1969 (O_1969,N_18482,N_18057);
nand UO_1970 (O_1970,N_17769,N_17439);
and UO_1971 (O_1971,N_17421,N_18134);
nand UO_1972 (O_1972,N_18180,N_16018);
nand UO_1973 (O_1973,N_19839,N_15997);
or UO_1974 (O_1974,N_16119,N_16337);
and UO_1975 (O_1975,N_18905,N_17235);
and UO_1976 (O_1976,N_15724,N_16869);
xor UO_1977 (O_1977,N_19969,N_15164);
nor UO_1978 (O_1978,N_15203,N_19886);
nand UO_1979 (O_1979,N_19627,N_17436);
nand UO_1980 (O_1980,N_19949,N_15948);
nand UO_1981 (O_1981,N_15074,N_17177);
or UO_1982 (O_1982,N_19765,N_15018);
nor UO_1983 (O_1983,N_15505,N_16747);
or UO_1984 (O_1984,N_15717,N_17798);
nand UO_1985 (O_1985,N_17518,N_16485);
and UO_1986 (O_1986,N_17249,N_19111);
and UO_1987 (O_1987,N_18174,N_18743);
nand UO_1988 (O_1988,N_17362,N_18357);
nand UO_1989 (O_1989,N_18232,N_19946);
nand UO_1990 (O_1990,N_17982,N_18237);
and UO_1991 (O_1991,N_16776,N_17318);
and UO_1992 (O_1992,N_15869,N_18560);
nand UO_1993 (O_1993,N_18801,N_19699);
or UO_1994 (O_1994,N_15030,N_17290);
nand UO_1995 (O_1995,N_18055,N_17528);
nor UO_1996 (O_1996,N_19856,N_17815);
and UO_1997 (O_1997,N_19522,N_15261);
nor UO_1998 (O_1998,N_15458,N_15971);
nor UO_1999 (O_1999,N_16357,N_15624);
and UO_2000 (O_2000,N_18467,N_19284);
and UO_2001 (O_2001,N_19645,N_16593);
or UO_2002 (O_2002,N_15468,N_15092);
nor UO_2003 (O_2003,N_18404,N_16735);
or UO_2004 (O_2004,N_15448,N_15135);
nor UO_2005 (O_2005,N_16233,N_17992);
and UO_2006 (O_2006,N_15417,N_17967);
nor UO_2007 (O_2007,N_18919,N_17911);
nand UO_2008 (O_2008,N_18973,N_18635);
nand UO_2009 (O_2009,N_19129,N_19961);
nor UO_2010 (O_2010,N_17219,N_15152);
nor UO_2011 (O_2011,N_17669,N_19386);
nand UO_2012 (O_2012,N_16490,N_18443);
nand UO_2013 (O_2013,N_15668,N_19240);
nand UO_2014 (O_2014,N_16773,N_19697);
nand UO_2015 (O_2015,N_17493,N_16992);
nand UO_2016 (O_2016,N_16503,N_18550);
and UO_2017 (O_2017,N_17802,N_18133);
or UO_2018 (O_2018,N_15524,N_19164);
and UO_2019 (O_2019,N_17927,N_16967);
nor UO_2020 (O_2020,N_16689,N_16629);
or UO_2021 (O_2021,N_19988,N_18172);
and UO_2022 (O_2022,N_18795,N_15210);
nor UO_2023 (O_2023,N_18456,N_17530);
and UO_2024 (O_2024,N_16712,N_19515);
xnor UO_2025 (O_2025,N_16416,N_15984);
or UO_2026 (O_2026,N_15737,N_16203);
or UO_2027 (O_2027,N_17223,N_18370);
nand UO_2028 (O_2028,N_16085,N_18045);
nor UO_2029 (O_2029,N_17618,N_18616);
nor UO_2030 (O_2030,N_17148,N_18930);
or UO_2031 (O_2031,N_15719,N_16056);
or UO_2032 (O_2032,N_17229,N_19457);
or UO_2033 (O_2033,N_18152,N_18118);
and UO_2034 (O_2034,N_19757,N_17544);
or UO_2035 (O_2035,N_19540,N_19307);
nand UO_2036 (O_2036,N_19139,N_17488);
nand UO_2037 (O_2037,N_17681,N_15637);
and UO_2038 (O_2038,N_16177,N_19990);
or UO_2039 (O_2039,N_15925,N_16681);
nor UO_2040 (O_2040,N_17286,N_15647);
nor UO_2041 (O_2041,N_17570,N_19229);
or UO_2042 (O_2042,N_16736,N_17036);
nor UO_2043 (O_2043,N_18234,N_19894);
and UO_2044 (O_2044,N_17173,N_17771);
or UO_2045 (O_2045,N_17537,N_16589);
nor UO_2046 (O_2046,N_16200,N_16264);
nor UO_2047 (O_2047,N_16559,N_18394);
nor UO_2048 (O_2048,N_16330,N_19624);
or UO_2049 (O_2049,N_19233,N_17985);
nand UO_2050 (O_2050,N_19613,N_18018);
nor UO_2051 (O_2051,N_18673,N_17316);
and UO_2052 (O_2052,N_17162,N_18274);
and UO_2053 (O_2053,N_19805,N_16524);
nor UO_2054 (O_2054,N_16385,N_19236);
nand UO_2055 (O_2055,N_19153,N_15052);
or UO_2056 (O_2056,N_16273,N_17118);
nor UO_2057 (O_2057,N_18939,N_18710);
nor UO_2058 (O_2058,N_17125,N_19721);
nand UO_2059 (O_2059,N_19006,N_15051);
nand UO_2060 (O_2060,N_17211,N_15122);
nor UO_2061 (O_2061,N_19319,N_15276);
nand UO_2062 (O_2062,N_19575,N_15467);
nand UO_2063 (O_2063,N_19594,N_15590);
nor UO_2064 (O_2064,N_19943,N_18623);
and UO_2065 (O_2065,N_16220,N_19939);
and UO_2066 (O_2066,N_17500,N_16423);
nand UO_2067 (O_2067,N_18065,N_19610);
xor UO_2068 (O_2068,N_15626,N_15118);
nand UO_2069 (O_2069,N_15123,N_15293);
nand UO_2070 (O_2070,N_19289,N_17450);
or UO_2071 (O_2071,N_16044,N_19260);
or UO_2072 (O_2072,N_18620,N_18580);
and UO_2073 (O_2073,N_16506,N_18856);
or UO_2074 (O_2074,N_18592,N_17511);
or UO_2075 (O_2075,N_17295,N_19175);
nand UO_2076 (O_2076,N_18936,N_16026);
and UO_2077 (O_2077,N_19276,N_16283);
nor UO_2078 (O_2078,N_19819,N_16571);
or UO_2079 (O_2079,N_18587,N_17120);
nand UO_2080 (O_2080,N_16533,N_15855);
and UO_2081 (O_2081,N_19138,N_18378);
nor UO_2082 (O_2082,N_19708,N_18033);
nor UO_2083 (O_2083,N_17740,N_19780);
and UO_2084 (O_2084,N_17668,N_15929);
or UO_2085 (O_2085,N_15163,N_17023);
nor UO_2086 (O_2086,N_19272,N_19095);
nor UO_2087 (O_2087,N_17877,N_15479);
nor UO_2088 (O_2088,N_16468,N_16617);
nor UO_2089 (O_2089,N_15402,N_19098);
nand UO_2090 (O_2090,N_15669,N_15586);
nand UO_2091 (O_2091,N_18533,N_16250);
nand UO_2092 (O_2092,N_15500,N_15989);
nand UO_2093 (O_2093,N_18828,N_19590);
and UO_2094 (O_2094,N_18317,N_17826);
nor UO_2095 (O_2095,N_18858,N_17660);
nand UO_2096 (O_2096,N_18175,N_19772);
or UO_2097 (O_2097,N_19019,N_18730);
nor UO_2098 (O_2098,N_17123,N_19574);
and UO_2099 (O_2099,N_19010,N_16522);
and UO_2100 (O_2100,N_18153,N_15125);
nand UO_2101 (O_2101,N_16963,N_17231);
nand UO_2102 (O_2102,N_15660,N_15621);
nand UO_2103 (O_2103,N_19116,N_15298);
or UO_2104 (O_2104,N_18672,N_19595);
nand UO_2105 (O_2105,N_15613,N_15422);
nand UO_2106 (O_2106,N_15838,N_19538);
or UO_2107 (O_2107,N_18735,N_18848);
and UO_2108 (O_2108,N_16002,N_18504);
nand UO_2109 (O_2109,N_18575,N_15857);
nor UO_2110 (O_2110,N_17027,N_18079);
nor UO_2111 (O_2111,N_17866,N_17002);
and UO_2112 (O_2112,N_17172,N_19335);
nand UO_2113 (O_2113,N_15842,N_19573);
or UO_2114 (O_2114,N_18535,N_18780);
nand UO_2115 (O_2115,N_16784,N_16146);
nor UO_2116 (O_2116,N_16793,N_19611);
and UO_2117 (O_2117,N_19901,N_16356);
and UO_2118 (O_2118,N_19876,N_17045);
and UO_2119 (O_2119,N_18521,N_18484);
nand UO_2120 (O_2120,N_17764,N_15552);
nor UO_2121 (O_2121,N_17255,N_18666);
and UO_2122 (O_2122,N_18875,N_18519);
nand UO_2123 (O_2123,N_15901,N_15996);
or UO_2124 (O_2124,N_17396,N_16724);
nor UO_2125 (O_2125,N_17855,N_17365);
and UO_2126 (O_2126,N_19922,N_19683);
nand UO_2127 (O_2127,N_17348,N_15170);
xor UO_2128 (O_2128,N_15107,N_19119);
and UO_2129 (O_2129,N_18265,N_17666);
or UO_2130 (O_2130,N_19954,N_16101);
and UO_2131 (O_2131,N_18736,N_18156);
nor UO_2132 (O_2132,N_15379,N_17475);
nand UO_2133 (O_2133,N_17315,N_19126);
nand UO_2134 (O_2134,N_16906,N_17862);
and UO_2135 (O_2135,N_17773,N_16171);
or UO_2136 (O_2136,N_17933,N_15388);
xnor UO_2137 (O_2137,N_18648,N_15918);
and UO_2138 (O_2138,N_16027,N_19451);
xor UO_2139 (O_2139,N_16400,N_16761);
nand UO_2140 (O_2140,N_17612,N_16472);
and UO_2141 (O_2141,N_19693,N_17806);
and UO_2142 (O_2142,N_17443,N_19321);
xor UO_2143 (O_2143,N_18619,N_18746);
nor UO_2144 (O_2144,N_15251,N_17455);
and UO_2145 (O_2145,N_17116,N_16388);
nor UO_2146 (O_2146,N_17832,N_19587);
and UO_2147 (O_2147,N_15600,N_19675);
nor UO_2148 (O_2148,N_16500,N_16595);
and UO_2149 (O_2149,N_16969,N_16700);
nor UO_2150 (O_2150,N_19930,N_17222);
nor UO_2151 (O_2151,N_15973,N_19169);
nor UO_2152 (O_2152,N_18308,N_18027);
and UO_2153 (O_2153,N_17962,N_19500);
nand UO_2154 (O_2154,N_17557,N_17224);
or UO_2155 (O_2155,N_19637,N_16270);
or UO_2156 (O_2156,N_18632,N_16771);
or UO_2157 (O_2157,N_15020,N_16977);
and UO_2158 (O_2158,N_17844,N_16108);
and UO_2159 (O_2159,N_15103,N_18997);
xnor UO_2160 (O_2160,N_19121,N_17282);
and UO_2161 (O_2161,N_15228,N_15935);
and UO_2162 (O_2162,N_17572,N_16308);
or UO_2163 (O_2163,N_17400,N_17667);
and UO_2164 (O_2164,N_17739,N_16246);
nand UO_2165 (O_2165,N_19158,N_18900);
nor UO_2166 (O_2166,N_16834,N_16690);
or UO_2167 (O_2167,N_16554,N_17614);
or UO_2168 (O_2168,N_18685,N_17692);
nand UO_2169 (O_2169,N_15167,N_17957);
or UO_2170 (O_2170,N_17277,N_17820);
nor UO_2171 (O_2171,N_18733,N_15840);
nor UO_2172 (O_2172,N_15097,N_17885);
nand UO_2173 (O_2173,N_15264,N_16498);
nand UO_2174 (O_2174,N_19433,N_16812);
nand UO_2175 (O_2175,N_19487,N_17132);
nor UO_2176 (O_2176,N_18085,N_16310);
nand UO_2177 (O_2177,N_19719,N_17997);
and UO_2178 (O_2178,N_18314,N_19266);
nand UO_2179 (O_2179,N_19090,N_16760);
or UO_2180 (O_2180,N_17800,N_19815);
and UO_2181 (O_2181,N_16779,N_18974);
nor UO_2182 (O_2182,N_16384,N_15389);
nand UO_2183 (O_2183,N_18053,N_18552);
or UO_2184 (O_2184,N_19582,N_17471);
and UO_2185 (O_2185,N_19480,N_17794);
nand UO_2186 (O_2186,N_17936,N_16669);
nand UO_2187 (O_2187,N_18998,N_18239);
nor UO_2188 (O_2188,N_18135,N_16597);
xor UO_2189 (O_2189,N_16073,N_15039);
nand UO_2190 (O_2190,N_17336,N_18013);
or UO_2191 (O_2191,N_17114,N_17988);
nor UO_2192 (O_2192,N_17458,N_18486);
or UO_2193 (O_2193,N_17634,N_18993);
and UO_2194 (O_2194,N_19346,N_16894);
or UO_2195 (O_2195,N_16467,N_17814);
nor UO_2196 (O_2196,N_19893,N_19903);
or UO_2197 (O_2197,N_16877,N_15029);
nor UO_2198 (O_2198,N_17520,N_15224);
nand UO_2199 (O_2199,N_16890,N_17496);
or UO_2200 (O_2200,N_19145,N_16886);
nand UO_2201 (O_2201,N_18505,N_17084);
or UO_2202 (O_2202,N_17079,N_19933);
nor UO_2203 (O_2203,N_18176,N_15815);
nand UO_2204 (O_2204,N_18392,N_19192);
or UO_2205 (O_2205,N_17218,N_19039);
nor UO_2206 (O_2206,N_19488,N_19635);
nor UO_2207 (O_2207,N_19898,N_16089);
or UO_2208 (O_2208,N_15747,N_16261);
and UO_2209 (O_2209,N_19742,N_16598);
or UO_2210 (O_2210,N_18411,N_17710);
nand UO_2211 (O_2211,N_18050,N_16755);
or UO_2212 (O_2212,N_19763,N_19660);
nand UO_2213 (O_2213,N_17104,N_17248);
nand UO_2214 (O_2214,N_16307,N_16518);
or UO_2215 (O_2215,N_15936,N_18813);
nand UO_2216 (O_2216,N_15922,N_18571);
and UO_2217 (O_2217,N_17356,N_16783);
nand UO_2218 (O_2218,N_15589,N_16657);
nand UO_2219 (O_2219,N_18490,N_18837);
and UO_2220 (O_2220,N_17109,N_17307);
or UO_2221 (O_2221,N_17469,N_16154);
and UO_2222 (O_2222,N_15889,N_15461);
nor UO_2223 (O_2223,N_15650,N_16280);
and UO_2224 (O_2224,N_18183,N_16258);
or UO_2225 (O_2225,N_17473,N_19279);
or UO_2226 (O_2226,N_15307,N_16769);
nand UO_2227 (O_2227,N_19589,N_15309);
nand UO_2228 (O_2228,N_17558,N_19106);
nand UO_2229 (O_2229,N_16070,N_18419);
xor UO_2230 (O_2230,N_15365,N_16619);
or UO_2231 (O_2231,N_19281,N_19013);
and UO_2232 (O_2232,N_19053,N_18857);
xor UO_2233 (O_2233,N_15802,N_15888);
nor UO_2234 (O_2234,N_16947,N_17624);
nor UO_2235 (O_2235,N_15766,N_16832);
or UO_2236 (O_2236,N_19292,N_16511);
or UO_2237 (O_2237,N_17285,N_19334);
or UO_2238 (O_2238,N_15708,N_19607);
nor UO_2239 (O_2239,N_18538,N_19118);
nand UO_2240 (O_2240,N_18372,N_18982);
or UO_2241 (O_2241,N_18951,N_15104);
or UO_2242 (O_2242,N_18940,N_16410);
or UO_2243 (O_2243,N_16744,N_17168);
or UO_2244 (O_2244,N_17440,N_19025);
and UO_2245 (O_2245,N_19004,N_18315);
nor UO_2246 (O_2246,N_18322,N_17418);
nor UO_2247 (O_2247,N_19992,N_15871);
nor UO_2248 (O_2248,N_17434,N_19475);
xnor UO_2249 (O_2249,N_16578,N_15768);
and UO_2250 (O_2250,N_19596,N_15335);
or UO_2251 (O_2251,N_15345,N_15395);
nand UO_2252 (O_2252,N_17187,N_16711);
or UO_2253 (O_2253,N_18488,N_18513);
or UO_2254 (O_2254,N_17313,N_17920);
nor UO_2255 (O_2255,N_16634,N_15777);
nand UO_2256 (O_2256,N_16751,N_19732);
nor UO_2257 (O_2257,N_18217,N_15172);
or UO_2258 (O_2258,N_17359,N_15638);
nor UO_2259 (O_2259,N_17091,N_19123);
nor UO_2260 (O_2260,N_19800,N_19796);
nor UO_2261 (O_2261,N_15401,N_19955);
nand UO_2262 (O_2262,N_17857,N_19114);
and UO_2263 (O_2263,N_16695,N_15580);
nor UO_2264 (O_2264,N_18332,N_17867);
xor UO_2265 (O_2265,N_16129,N_16682);
and UO_2266 (O_2266,N_19091,N_19234);
and UO_2267 (O_2267,N_19065,N_18200);
nor UO_2268 (O_2268,N_17310,N_17573);
and UO_2269 (O_2269,N_16986,N_16251);
nor UO_2270 (O_2270,N_16473,N_18407);
nand UO_2271 (O_2271,N_15087,N_18777);
or UO_2272 (O_2272,N_16921,N_15959);
nand UO_2273 (O_2273,N_19730,N_19668);
or UO_2274 (O_2274,N_16354,N_19206);
or UO_2275 (O_2275,N_15279,N_16944);
or UO_2276 (O_2276,N_19561,N_17204);
nor UO_2277 (O_2277,N_18741,N_19846);
or UO_2278 (O_2278,N_16999,N_18142);
nor UO_2279 (O_2279,N_15726,N_16548);
nor UO_2280 (O_2280,N_16643,N_16892);
or UO_2281 (O_2281,N_19096,N_16185);
nand UO_2282 (O_2282,N_18605,N_16684);
nand UO_2283 (O_2283,N_18463,N_19705);
xor UO_2284 (O_2284,N_16929,N_17907);
nor UO_2285 (O_2285,N_17938,N_15041);
nor UO_2286 (O_2286,N_15540,N_15892);
nand UO_2287 (O_2287,N_17596,N_16074);
or UO_2288 (O_2288,N_18031,N_16517);
or UO_2289 (O_2289,N_19556,N_17199);
nor UO_2290 (O_2290,N_16179,N_18103);
xor UO_2291 (O_2291,N_18123,N_16883);
nand UO_2292 (O_2292,N_16377,N_18479);
nor UO_2293 (O_2293,N_19382,N_15520);
and UO_2294 (O_2294,N_18812,N_15048);
nor UO_2295 (O_2295,N_17461,N_18006);
or UO_2296 (O_2296,N_15924,N_15469);
and UO_2297 (O_2297,N_16767,N_15696);
and UO_2298 (O_2298,N_15976,N_19960);
nand UO_2299 (O_2299,N_18893,N_19297);
or UO_2300 (O_2300,N_17234,N_16950);
and UO_2301 (O_2301,N_18406,N_15348);
nand UO_2302 (O_2302,N_18344,N_16730);
or UO_2303 (O_2303,N_17323,N_15926);
or UO_2304 (O_2304,N_17408,N_17142);
nor UO_2305 (O_2305,N_17126,N_17275);
nor UO_2306 (O_2306,N_17712,N_17601);
and UO_2307 (O_2307,N_15459,N_15142);
and UO_2308 (O_2308,N_18984,N_17772);
nand UO_2309 (O_2309,N_18756,N_16141);
nor UO_2310 (O_2310,N_18362,N_15259);
and UO_2311 (O_2311,N_17915,N_17905);
nor UO_2312 (O_2312,N_15547,N_15391);
or UO_2313 (O_2313,N_15486,N_15397);
or UO_2314 (O_2314,N_17279,N_17847);
and UO_2315 (O_2315,N_18938,N_15286);
and UO_2316 (O_2316,N_15774,N_17636);
or UO_2317 (O_2317,N_18671,N_15522);
nand UO_2318 (O_2318,N_19612,N_16752);
or UO_2319 (O_2319,N_19756,N_16839);
and UO_2320 (O_2320,N_17567,N_16319);
and UO_2321 (O_2321,N_15431,N_15438);
xnor UO_2322 (O_2322,N_17959,N_19521);
or UO_2323 (O_2323,N_17251,N_19494);
nand UO_2324 (O_2324,N_18871,N_16826);
and UO_2325 (O_2325,N_16175,N_19246);
xor UO_2326 (O_2326,N_17169,N_17308);
xnor UO_2327 (O_2327,N_17828,N_16199);
nand UO_2328 (O_2328,N_19209,N_18653);
or UO_2329 (O_2329,N_16142,N_16502);
and UO_2330 (O_2330,N_18022,N_19453);
nand UO_2331 (O_2331,N_15513,N_15526);
or UO_2332 (O_2332,N_19950,N_18863);
or UO_2333 (O_2333,N_18335,N_17715);
or UO_2334 (O_2334,N_19372,N_18225);
or UO_2335 (O_2335,N_15785,N_17781);
xnor UO_2336 (O_2336,N_16364,N_19212);
nand UO_2337 (O_2337,N_15885,N_18713);
nand UO_2338 (O_2338,N_15735,N_17050);
and UO_2339 (O_2339,N_15057,N_19299);
or UO_2340 (O_2340,N_15204,N_19185);
nor UO_2341 (O_2341,N_15003,N_18011);
and UO_2342 (O_2342,N_17266,N_16920);
nand UO_2343 (O_2343,N_18252,N_16197);
or UO_2344 (O_2344,N_17553,N_19598);
or UO_2345 (O_2345,N_15031,N_17965);
and UO_2346 (O_2346,N_17143,N_16172);
nor UO_2347 (O_2347,N_17616,N_19917);
nor UO_2348 (O_2348,N_18214,N_17729);
nor UO_2349 (O_2349,N_18292,N_19971);
or UO_2350 (O_2350,N_15067,N_16961);
nand UO_2351 (O_2351,N_18737,N_17966);
nand UO_2352 (O_2352,N_17284,N_18720);
and UO_2353 (O_2353,N_19885,N_19639);
and UO_2354 (O_2354,N_18326,N_19869);
nor UO_2355 (O_2355,N_16916,N_17127);
nand UO_2356 (O_2356,N_15495,N_19149);
or UO_2357 (O_2357,N_15416,N_19968);
and UO_2358 (O_2358,N_17203,N_15872);
nor UO_2359 (O_2359,N_18034,N_16352);
nor UO_2360 (O_2360,N_19089,N_17838);
nor UO_2361 (O_2361,N_15847,N_18830);
and UO_2362 (O_2362,N_15077,N_18916);
and UO_2363 (O_2363,N_18303,N_19891);
or UO_2364 (O_2364,N_18942,N_15544);
nand UO_2365 (O_2365,N_17108,N_16610);
nor UO_2366 (O_2366,N_15131,N_15951);
or UO_2367 (O_2367,N_17456,N_15679);
or UO_2368 (O_2368,N_19516,N_18377);
xnor UO_2369 (O_2369,N_16451,N_17925);
and UO_2370 (O_2370,N_15287,N_19563);
nor UO_2371 (O_2371,N_17827,N_17186);
nor UO_2372 (O_2372,N_16970,N_16737);
xor UO_2373 (O_2373,N_18030,N_17001);
nand UO_2374 (O_2374,N_15326,N_19204);
or UO_2375 (O_2375,N_15692,N_19202);
and UO_2376 (O_2376,N_17742,N_18892);
nand UO_2377 (O_2377,N_17314,N_15736);
nand UO_2378 (O_2378,N_16655,N_18208);
or UO_2379 (O_2379,N_19667,N_18907);
or UO_2380 (O_2380,N_17004,N_15743);
nor UO_2381 (O_2381,N_17935,N_19482);
and UO_2382 (O_2382,N_16880,N_15946);
or UO_2383 (O_2383,N_18526,N_16182);
or UO_2384 (O_2384,N_15155,N_18365);
and UO_2385 (O_2385,N_16240,N_16825);
or UO_2386 (O_2386,N_17435,N_17352);
nor UO_2387 (O_2387,N_17741,N_17228);
nand UO_2388 (O_2388,N_17128,N_17723);
nor UO_2389 (O_2389,N_17964,N_18051);
or UO_2390 (O_2390,N_18723,N_17807);
nor UO_2391 (O_2391,N_18506,N_19424);
nor UO_2392 (O_2392,N_17361,N_19373);
and UO_2393 (O_2393,N_18574,N_16549);
nand UO_2394 (O_2394,N_15742,N_19959);
and UO_2395 (O_2395,N_15617,N_18204);
nor UO_2396 (O_2396,N_16808,N_17382);
or UO_2397 (O_2397,N_18442,N_15195);
and UO_2398 (O_2398,N_17842,N_17917);
nor UO_2399 (O_2399,N_16428,N_16497);
nor UO_2400 (O_2400,N_16278,N_15403);
or UO_2401 (O_2401,N_17647,N_18267);
and UO_2402 (O_2402,N_18293,N_18008);
nand UO_2403 (O_2403,N_15853,N_15130);
and UO_2404 (O_2404,N_15429,N_19811);
and UO_2405 (O_2405,N_18923,N_15727);
or UO_2406 (O_2406,N_17909,N_18054);
nor UO_2407 (O_2407,N_17673,N_16359);
nor UO_2408 (O_2408,N_18244,N_17046);
and UO_2409 (O_2409,N_19313,N_18948);
and UO_2410 (O_2410,N_16486,N_19528);
nor UO_2411 (O_2411,N_15791,N_16050);
nand UO_2412 (O_2412,N_15308,N_16301);
or UO_2413 (O_2413,N_17353,N_18836);
or UO_2414 (O_2414,N_19848,N_17973);
and UO_2415 (O_2415,N_18883,N_15275);
and UO_2416 (O_2416,N_18472,N_19351);
or UO_2417 (O_2417,N_17304,N_17380);
nand UO_2418 (O_2418,N_19462,N_15602);
and UO_2419 (O_2419,N_15315,N_18190);
or UO_2420 (O_2420,N_19349,N_18920);
and UO_2421 (O_2421,N_17175,N_16396);
and UO_2422 (O_2422,N_15043,N_19747);
nor UO_2423 (O_2423,N_17685,N_18788);
or UO_2424 (O_2424,N_17477,N_17979);
nor UO_2425 (O_2425,N_15663,N_17347);
or UO_2426 (O_2426,N_15421,N_16483);
nand UO_2427 (O_2427,N_19042,N_16000);
and UO_2428 (O_2428,N_16290,N_16302);
nand UO_2429 (O_2429,N_17556,N_17504);
or UO_2430 (O_2430,N_16215,N_18184);
nor UO_2431 (O_2431,N_15754,N_19555);
nand UO_2432 (O_2432,N_16031,N_17824);
or UO_2433 (O_2433,N_18704,N_15913);
nor UO_2434 (O_2434,N_19777,N_19783);
or UO_2435 (O_2435,N_18686,N_16647);
and UO_2436 (O_2436,N_17497,N_15359);
xor UO_2437 (O_2437,N_17140,N_19160);
nand UO_2438 (O_2438,N_17950,N_16083);
nand UO_2439 (O_2439,N_17152,N_17355);
and UO_2440 (O_2440,N_16057,N_16579);
nor UO_2441 (O_2441,N_15055,N_19407);
nand UO_2442 (O_2442,N_17306,N_17659);
nor UO_2443 (O_2443,N_17887,N_19466);
and UO_2444 (O_2444,N_15136,N_18108);
and UO_2445 (O_2445,N_17783,N_19075);
nor UO_2446 (O_2446,N_16978,N_17189);
and UO_2447 (O_2447,N_17099,N_16546);
nor UO_2448 (O_2448,N_17372,N_16113);
or UO_2449 (O_2449,N_16875,N_17014);
or UO_2450 (O_2450,N_17819,N_19562);
nor UO_2451 (O_2451,N_17257,N_19367);
or UO_2452 (O_2452,N_18891,N_17107);
and UO_2453 (O_2453,N_18465,N_18191);
and UO_2454 (O_2454,N_17841,N_16715);
nor UO_2455 (O_2455,N_19221,N_18089);
nand UO_2456 (O_2456,N_16494,N_15408);
or UO_2457 (O_2457,N_19495,N_16208);
nor UO_2458 (O_2458,N_15499,N_19405);
nor UO_2459 (O_2459,N_17949,N_16581);
or UO_2460 (O_2460,N_18608,N_17503);
nor UO_2461 (O_2461,N_17682,N_18578);
or UO_2462 (O_2462,N_18944,N_16107);
nor UO_2463 (O_2463,N_17334,N_19890);
and UO_2464 (O_2464,N_16153,N_18386);
nor UO_2465 (O_2465,N_17693,N_17268);
nor UO_2466 (O_2466,N_15085,N_16256);
or UO_2467 (O_2467,N_17678,N_19539);
nor UO_2468 (O_2468,N_18870,N_18092);
or UO_2469 (O_2469,N_17649,N_15146);
and UO_2470 (O_2470,N_15786,N_15978);
nand UO_2471 (O_2471,N_15927,N_15037);
or UO_2472 (O_2472,N_16445,N_15702);
nand UO_2473 (O_2473,N_19723,N_17149);
or UO_2474 (O_2474,N_17754,N_19744);
nor UO_2475 (O_2475,N_18638,N_19534);
and UO_2476 (O_2476,N_18347,N_15460);
and UO_2477 (O_2477,N_18037,N_19863);
or UO_2478 (O_2478,N_18218,N_16895);
and UO_2479 (O_2479,N_16211,N_15413);
nand UO_2480 (O_2480,N_16591,N_15435);
nor UO_2481 (O_2481,N_18097,N_18121);
and UO_2482 (O_2482,N_19029,N_19735);
nor UO_2483 (O_2483,N_18640,N_15963);
or UO_2484 (O_2484,N_17981,N_17664);
and UO_2485 (O_2485,N_15661,N_17061);
or UO_2486 (O_2486,N_15208,N_17287);
nand UO_2487 (O_2487,N_16550,N_15423);
or UO_2488 (O_2488,N_16004,N_16501);
nand UO_2489 (O_2489,N_18131,N_19207);
or UO_2490 (O_2490,N_19964,N_19225);
nor UO_2491 (O_2491,N_18902,N_16840);
nand UO_2492 (O_2492,N_16889,N_15521);
nand UO_2493 (O_2493,N_16603,N_15137);
or UO_2494 (O_2494,N_16656,N_17913);
nor UO_2495 (O_2495,N_17164,N_19046);
nand UO_2496 (O_2496,N_19731,N_19586);
and UO_2497 (O_2497,N_19778,N_19507);
and UO_2498 (O_2498,N_16819,N_19568);
or UO_2499 (O_2499,N_19814,N_16828);
endmodule