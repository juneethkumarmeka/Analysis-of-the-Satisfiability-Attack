module basic_1000_10000_1500_4_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_634,In_856);
nand U1 (N_1,In_246,In_91);
nand U2 (N_2,In_290,In_54);
nand U3 (N_3,In_212,In_975);
nand U4 (N_4,In_579,In_673);
and U5 (N_5,In_82,In_0);
and U6 (N_6,In_731,In_776);
and U7 (N_7,In_779,In_648);
and U8 (N_8,In_245,In_156);
and U9 (N_9,In_869,In_842);
nand U10 (N_10,In_332,In_665);
or U11 (N_11,In_461,In_352);
xnor U12 (N_12,In_734,In_284);
and U13 (N_13,In_220,In_31);
or U14 (N_14,In_580,In_900);
or U15 (N_15,In_918,In_688);
nor U16 (N_16,In_68,In_594);
or U17 (N_17,In_355,In_961);
nand U18 (N_18,In_824,In_478);
nand U19 (N_19,In_985,In_769);
nor U20 (N_20,In_440,In_368);
and U21 (N_21,In_158,In_655);
nand U22 (N_22,In_135,In_996);
nor U23 (N_23,In_690,In_520);
and U24 (N_24,In_118,In_744);
or U25 (N_25,In_818,In_637);
xor U26 (N_26,In_765,In_871);
nor U27 (N_27,In_854,In_739);
nand U28 (N_28,In_396,In_259);
xor U29 (N_29,In_325,In_280);
xor U30 (N_30,In_9,In_979);
and U31 (N_31,In_834,In_173);
nand U32 (N_32,In_953,In_906);
xnor U33 (N_33,In_131,In_586);
and U34 (N_34,In_968,In_606);
nor U35 (N_35,In_73,In_514);
xor U36 (N_36,In_194,In_11);
xnor U37 (N_37,In_427,In_149);
nand U38 (N_38,In_452,In_876);
or U39 (N_39,In_242,In_923);
xor U40 (N_40,In_881,In_130);
nand U41 (N_41,In_970,In_879);
nor U42 (N_42,In_201,In_140);
nand U43 (N_43,In_784,In_311);
xnor U44 (N_44,In_342,In_340);
xor U45 (N_45,In_182,In_184);
xnor U46 (N_46,In_473,In_510);
nor U47 (N_47,In_525,In_597);
nand U48 (N_48,In_30,In_12);
nand U49 (N_49,In_963,In_123);
xnor U50 (N_50,In_70,In_945);
xnor U51 (N_51,In_449,In_202);
nand U52 (N_52,In_708,In_71);
and U53 (N_53,In_113,In_470);
nand U54 (N_54,In_800,In_518);
or U55 (N_55,In_115,In_134);
and U56 (N_56,In_385,In_763);
nor U57 (N_57,In_468,In_837);
and U58 (N_58,In_602,In_767);
nor U59 (N_59,In_86,In_614);
and U60 (N_60,In_629,In_335);
xor U61 (N_61,In_926,In_236);
nand U62 (N_62,In_79,In_787);
or U63 (N_63,In_962,In_974);
or U64 (N_64,In_406,In_596);
nand U65 (N_65,In_475,In_491);
nand U66 (N_66,In_551,In_388);
nor U67 (N_67,In_600,In_395);
and U68 (N_68,In_568,In_747);
nor U69 (N_69,In_746,In_870);
or U70 (N_70,In_270,In_691);
or U71 (N_71,In_289,In_847);
nand U72 (N_72,In_277,In_208);
or U73 (N_73,In_896,In_296);
nor U74 (N_74,In_171,In_556);
or U75 (N_75,In_503,In_840);
xnor U76 (N_76,In_183,In_790);
or U77 (N_77,In_102,In_852);
xor U78 (N_78,In_728,In_861);
nand U79 (N_79,In_207,In_855);
and U80 (N_80,In_213,In_61);
or U81 (N_81,In_720,In_210);
nor U82 (N_82,In_110,In_932);
xnor U83 (N_83,In_345,In_257);
nand U84 (N_84,In_867,In_766);
xnor U85 (N_85,In_38,In_741);
nor U86 (N_86,In_114,In_391);
and U87 (N_87,In_294,In_628);
and U88 (N_88,In_901,In_850);
xor U89 (N_89,In_999,In_365);
nand U90 (N_90,In_862,In_612);
xnor U91 (N_91,In_951,In_694);
or U92 (N_92,In_451,In_549);
nor U93 (N_93,In_160,In_826);
and U94 (N_94,In_682,In_1);
xnor U95 (N_95,In_922,In_442);
and U96 (N_96,In_557,In_838);
nand U97 (N_97,In_804,In_84);
or U98 (N_98,In_785,In_490);
nor U99 (N_99,In_439,In_796);
xor U100 (N_100,In_816,In_947);
xnor U101 (N_101,In_959,In_987);
nor U102 (N_102,In_904,In_578);
xnor U103 (N_103,In_89,In_316);
nand U104 (N_104,In_954,In_434);
and U105 (N_105,In_209,In_788);
xor U106 (N_106,In_991,In_735);
or U107 (N_107,In_370,In_76);
or U108 (N_108,In_77,In_255);
or U109 (N_109,In_295,In_320);
or U110 (N_110,In_562,In_402);
nor U111 (N_111,In_833,In_431);
or U112 (N_112,In_423,In_969);
or U113 (N_113,In_39,In_567);
or U114 (N_114,In_550,In_367);
or U115 (N_115,In_692,In_531);
xor U116 (N_116,In_249,In_821);
and U117 (N_117,In_832,In_40);
or U118 (N_118,In_541,In_193);
nor U119 (N_119,In_438,In_920);
nor U120 (N_120,In_492,In_302);
nand U121 (N_121,In_87,In_122);
nand U122 (N_122,In_573,In_234);
and U123 (N_123,In_774,In_286);
nand U124 (N_124,In_253,In_155);
or U125 (N_125,In_712,In_248);
xnor U126 (N_126,In_482,In_943);
and U127 (N_127,In_15,In_757);
or U128 (N_128,In_453,In_725);
nor U129 (N_129,In_143,In_397);
or U130 (N_130,In_559,In_481);
or U131 (N_131,In_946,In_955);
nand U132 (N_132,In_458,In_374);
nor U133 (N_133,In_530,In_146);
and U134 (N_134,In_351,In_697);
or U135 (N_135,In_237,In_254);
or U136 (N_136,In_915,In_74);
nor U137 (N_137,In_732,In_886);
or U138 (N_138,In_174,In_601);
or U139 (N_139,In_807,In_719);
nor U140 (N_140,In_334,In_211);
nand U141 (N_141,In_125,In_252);
or U142 (N_142,In_69,In_882);
nor U143 (N_143,In_674,In_401);
nor U144 (N_144,In_398,In_136);
nor U145 (N_145,In_474,In_772);
xor U146 (N_146,In_263,In_362);
nand U147 (N_147,In_233,In_812);
and U148 (N_148,In_321,In_545);
nor U149 (N_149,In_190,In_306);
nor U150 (N_150,In_144,In_327);
or U151 (N_151,In_792,In_166);
or U152 (N_152,In_815,In_686);
xor U153 (N_153,In_843,In_866);
nor U154 (N_154,In_786,In_319);
xor U155 (N_155,In_226,In_200);
and U156 (N_156,In_808,In_643);
nand U157 (N_157,In_456,In_488);
nor U158 (N_158,In_783,In_262);
and U159 (N_159,In_811,In_21);
and U160 (N_160,In_749,In_161);
nand U161 (N_161,In_275,In_25);
and U162 (N_162,In_960,In_828);
nand U163 (N_163,In_639,In_126);
nand U164 (N_164,In_417,In_799);
or U165 (N_165,In_803,In_446);
and U166 (N_166,In_758,In_436);
or U167 (N_167,In_225,In_934);
nor U168 (N_168,In_264,In_657);
nand U169 (N_169,In_661,In_891);
xor U170 (N_170,In_421,In_420);
and U171 (N_171,In_930,In_20);
xor U172 (N_172,In_291,In_328);
nand U173 (N_173,In_221,In_384);
xnor U174 (N_174,In_56,In_888);
nor U175 (N_175,In_464,In_768);
xnor U176 (N_176,In_369,In_971);
nor U177 (N_177,In_713,In_825);
nor U178 (N_178,In_952,In_874);
and U179 (N_179,In_309,In_724);
xor U180 (N_180,In_98,In_572);
nor U181 (N_181,In_455,In_375);
nor U182 (N_182,In_459,In_469);
and U183 (N_183,In_10,In_159);
nand U184 (N_184,In_889,In_487);
xor U185 (N_185,In_917,In_517);
and U186 (N_186,In_244,In_903);
nand U187 (N_187,In_293,In_693);
xnor U188 (N_188,In_631,In_312);
nor U189 (N_189,In_479,In_218);
and U190 (N_190,In_329,In_885);
xor U191 (N_191,In_83,In_680);
xnor U192 (N_192,In_145,In_878);
or U193 (N_193,In_829,In_499);
nor U194 (N_194,In_192,In_152);
or U195 (N_195,In_288,In_34);
and U196 (N_196,In_48,In_256);
and U197 (N_197,In_495,In_528);
and U198 (N_198,In_989,In_887);
nand U199 (N_199,In_120,In_186);
or U200 (N_200,In_644,In_623);
nand U201 (N_201,In_515,In_860);
or U202 (N_202,In_88,In_6);
and U203 (N_203,In_791,In_409);
and U204 (N_204,In_872,In_611);
and U205 (N_205,In_511,In_343);
or U206 (N_206,In_205,In_260);
or U207 (N_207,In_875,In_621);
nor U208 (N_208,In_645,In_63);
or U209 (N_209,In_323,In_378);
nand U210 (N_210,In_18,In_179);
or U211 (N_211,In_718,In_809);
or U212 (N_212,In_435,In_32);
xor U213 (N_213,In_506,In_806);
nand U214 (N_214,In_933,In_51);
nand U215 (N_215,In_589,In_373);
nand U216 (N_216,In_138,In_188);
or U217 (N_217,In_273,In_675);
and U218 (N_218,In_627,In_711);
and U219 (N_219,In_232,In_777);
nor U220 (N_220,In_700,In_668);
nand U221 (N_221,In_169,In_267);
and U222 (N_222,In_865,In_705);
or U223 (N_223,In_995,In_723);
nor U224 (N_224,In_948,In_677);
or U225 (N_225,In_868,In_425);
nor U226 (N_226,In_571,In_949);
nand U227 (N_227,In_941,In_973);
nand U228 (N_228,In_419,In_782);
and U229 (N_229,In_507,In_727);
nor U230 (N_230,In_215,In_574);
xor U231 (N_231,In_582,In_607);
xnor U232 (N_232,In_914,In_992);
nand U233 (N_233,In_921,In_957);
nor U234 (N_234,In_199,In_781);
and U235 (N_235,In_685,In_14);
nand U236 (N_236,In_383,In_181);
xor U237 (N_237,In_990,In_465);
and U238 (N_238,In_229,In_944);
xor U239 (N_239,In_128,In_658);
nand U240 (N_240,In_737,In_372);
nor U241 (N_241,In_736,In_641);
nand U242 (N_242,In_981,In_392);
and U243 (N_243,In_471,In_33);
and U244 (N_244,In_44,In_195);
nor U245 (N_245,In_618,In_537);
nor U246 (N_246,In_448,In_617);
and U247 (N_247,In_432,In_381);
nor U248 (N_248,In_976,In_356);
nand U249 (N_249,In_78,In_544);
nor U250 (N_250,In_911,In_738);
nor U251 (N_251,In_346,In_137);
nor U252 (N_252,In_997,In_780);
nor U253 (N_253,In_897,In_980);
nor U254 (N_254,In_415,In_937);
nor U255 (N_255,In_908,In_984);
xnor U256 (N_256,In_927,In_462);
or U257 (N_257,In_170,In_65);
nand U258 (N_258,In_521,In_216);
or U259 (N_259,In_116,In_928);
or U260 (N_260,In_303,In_42);
nor U261 (N_261,In_710,In_50);
xor U262 (N_262,In_743,In_197);
or U263 (N_263,In_247,In_52);
or U264 (N_264,In_43,In_827);
and U265 (N_265,In_111,In_543);
or U266 (N_266,In_2,In_287);
xor U267 (N_267,In_411,In_377);
or U268 (N_268,In_104,In_272);
nor U269 (N_269,In_412,In_85);
nand U270 (N_270,In_533,In_271);
xnor U271 (N_271,In_986,In_929);
xnor U272 (N_272,In_912,In_22);
or U273 (N_273,In_656,In_844);
and U274 (N_274,In_576,In_106);
and U275 (N_275,In_467,In_466);
nand U276 (N_276,In_925,In_715);
nor U277 (N_277,In_733,In_307);
or U278 (N_278,In_638,In_347);
or U279 (N_279,In_240,In_297);
and U280 (N_280,In_709,In_49);
nor U281 (N_281,In_336,In_622);
nand U282 (N_282,In_413,In_555);
and U283 (N_283,In_414,In_36);
nand U284 (N_284,In_707,In_176);
nand U285 (N_285,In_938,In_841);
or U286 (N_286,In_222,In_793);
and U287 (N_287,In_721,In_157);
and U288 (N_288,In_848,In_717);
xnor U289 (N_289,In_164,In_552);
nor U290 (N_290,In_105,In_112);
nor U291 (N_291,In_62,In_390);
xnor U292 (N_292,In_433,In_554);
and U293 (N_293,In_745,In_539);
nor U294 (N_294,In_967,In_814);
nand U295 (N_295,In_298,In_29);
or U296 (N_296,In_310,In_588);
or U297 (N_297,In_142,In_317);
and U298 (N_298,In_133,In_858);
nor U299 (N_299,In_836,In_810);
xor U300 (N_300,In_513,In_585);
xor U301 (N_301,In_99,In_817);
or U302 (N_302,In_163,In_258);
and U303 (N_303,In_24,In_857);
nor U304 (N_304,In_41,In_823);
xnor U305 (N_305,In_523,In_109);
or U306 (N_306,In_662,In_407);
and U307 (N_307,In_95,In_742);
nand U308 (N_308,In_416,In_714);
nor U309 (N_309,In_379,In_204);
or U310 (N_310,In_338,In_57);
xnor U311 (N_311,In_331,In_304);
nor U312 (N_312,In_94,In_172);
nor U313 (N_313,In_505,In_129);
or U314 (N_314,In_910,In_266);
and U315 (N_315,In_498,In_651);
or U316 (N_316,In_426,In_380);
and U317 (N_317,In_935,In_972);
or U318 (N_318,In_687,In_563);
and U319 (N_319,In_250,In_584);
nor U320 (N_320,In_701,In_667);
xnor U321 (N_321,In_97,In_382);
nor U322 (N_322,In_178,In_67);
and U323 (N_323,In_292,In_931);
nor U324 (N_324,In_909,In_353);
nand U325 (N_325,In_450,In_616);
nand U326 (N_326,In_845,In_529);
nand U327 (N_327,In_532,In_13);
nor U328 (N_328,In_595,In_276);
and U329 (N_329,In_484,In_239);
and U330 (N_330,In_626,In_536);
nand U331 (N_331,In_496,In_28);
nor U332 (N_332,In_96,In_154);
nand U333 (N_333,In_350,In_704);
nand U334 (N_334,In_604,In_168);
nand U335 (N_335,In_268,In_630);
and U336 (N_336,In_359,In_647);
nor U337 (N_337,In_569,In_472);
nand U338 (N_338,In_940,In_447);
or U339 (N_339,In_764,In_441);
and U340 (N_340,In_592,In_75);
nor U341 (N_341,In_366,In_561);
and U342 (N_342,In_820,In_399);
nor U343 (N_343,In_8,In_101);
nand U344 (N_344,In_750,In_805);
nand U345 (N_345,In_180,In_902);
nand U346 (N_346,In_357,In_919);
nor U347 (N_347,In_802,In_924);
nand U348 (N_348,In_666,In_830);
or U349 (N_349,In_534,In_486);
and U350 (N_350,In_587,In_660);
nand U351 (N_351,In_650,In_877);
xnor U352 (N_352,In_620,In_740);
xor U353 (N_353,In_653,In_35);
and U354 (N_354,In_679,In_635);
nor U355 (N_355,In_333,In_227);
nand U356 (N_356,In_408,In_497);
or U357 (N_357,In_983,In_393);
nand U358 (N_358,In_801,In_880);
nor U359 (N_359,In_219,In_754);
or U360 (N_360,In_978,In_760);
xor U361 (N_361,In_894,In_548);
nand U362 (N_362,In_994,In_299);
and U363 (N_363,In_939,In_913);
nor U364 (N_364,In_354,In_613);
nor U365 (N_365,In_835,In_813);
nor U366 (N_366,In_19,In_16);
xor U367 (N_367,In_422,In_851);
nor U368 (N_368,In_203,In_640);
and U369 (N_369,In_608,In_722);
xor U370 (N_370,In_993,In_17);
nand U371 (N_371,In_535,In_863);
nand U372 (N_372,In_956,In_771);
nand U373 (N_373,In_936,In_527);
nand U374 (N_374,In_753,In_755);
nor U375 (N_375,In_706,In_214);
nor U376 (N_376,In_494,In_798);
or U377 (N_377,In_916,In_235);
nand U378 (N_378,In_403,In_404);
xnor U379 (N_379,In_698,In_437);
nor U380 (N_380,In_93,In_890);
and U381 (N_381,In_577,In_907);
nand U382 (N_382,In_389,In_965);
and U383 (N_383,In_699,In_90);
nand U384 (N_384,In_560,In_405);
or U385 (N_385,In_565,In_37);
xor U386 (N_386,In_703,In_859);
xnor U387 (N_387,In_301,In_274);
xnor U388 (N_388,In_483,In_324);
xnor U389 (N_389,In_726,In_341);
nor U390 (N_390,In_278,In_669);
or U391 (N_391,In_66,In_477);
and U392 (N_392,In_175,In_831);
xnor U393 (N_393,In_187,In_230);
nor U394 (N_394,In_598,In_326);
nor U395 (N_395,In_678,In_748);
and U396 (N_396,In_189,In_26);
or U397 (N_397,In_558,In_376);
and U398 (N_398,In_261,In_313);
and U399 (N_399,In_898,In_609);
or U400 (N_400,In_371,In_581);
nand U401 (N_401,In_53,In_676);
nor U402 (N_402,In_58,In_873);
nand U403 (N_403,In_55,In_633);
nand U404 (N_404,In_251,In_538);
nor U405 (N_405,In_729,In_684);
and U406 (N_406,In_443,In_241);
nor U407 (N_407,In_636,In_778);
xor U408 (N_408,In_162,In_958);
xor U409 (N_409,In_476,In_337);
or U410 (N_410,In_315,In_540);
nand U411 (N_411,In_547,In_72);
and U412 (N_412,In_762,In_400);
nand U413 (N_413,In_387,In_198);
nand U414 (N_414,In_615,In_654);
xor U415 (N_415,In_839,In_348);
and U416 (N_416,In_853,In_480);
nand U417 (N_417,In_206,In_689);
or U418 (N_418,In_4,In_45);
or U419 (N_419,In_493,In_27);
xor U420 (N_420,In_759,In_141);
nor U421 (N_421,In_695,In_509);
and U422 (N_422,In_716,In_117);
nand U423 (N_423,In_454,In_121);
nand U424 (N_424,In_512,In_167);
xnor U425 (N_425,In_982,In_864);
or U426 (N_426,In_964,In_457);
nand U427 (N_427,In_108,In_883);
nand U428 (N_428,In_730,In_150);
nor U429 (N_429,In_279,In_500);
nor U430 (N_430,In_761,In_794);
xnor U431 (N_431,In_81,In_504);
nor U432 (N_432,In_895,In_671);
nand U433 (N_433,In_147,In_23);
nand U434 (N_434,In_905,In_224);
nor U435 (N_435,In_223,In_575);
or U436 (N_436,In_508,In_463);
or U437 (N_437,In_683,In_652);
and U438 (N_438,In_7,In_893);
nand U439 (N_439,In_265,In_314);
xor U440 (N_440,In_564,In_430);
and U441 (N_441,In_132,In_217);
xor U442 (N_442,In_501,In_702);
nor U443 (N_443,In_770,In_489);
nor U444 (N_444,In_165,In_542);
and U445 (N_445,In_177,In_360);
xnor U446 (N_446,In_46,In_269);
nand U447 (N_447,In_119,In_460);
nor U448 (N_448,In_153,In_899);
or U449 (N_449,In_445,In_308);
xnor U450 (N_450,In_566,In_591);
nand U451 (N_451,In_364,In_522);
and U452 (N_452,In_191,In_977);
nor U453 (N_453,In_139,In_305);
nand U454 (N_454,In_752,In_649);
xnor U455 (N_455,In_349,In_5);
or U456 (N_456,In_625,In_599);
xor U457 (N_457,In_59,In_570);
nor U458 (N_458,In_428,In_526);
and U459 (N_459,In_322,In_281);
and U460 (N_460,In_282,In_361);
xnor U461 (N_461,In_358,In_664);
xnor U462 (N_462,In_546,In_231);
nor U463 (N_463,In_60,In_797);
xnor U464 (N_464,In_751,In_795);
nor U465 (N_465,In_363,In_127);
xor U466 (N_466,In_988,In_502);
nor U467 (N_467,In_386,In_646);
xnor U468 (N_468,In_819,In_80);
nor U469 (N_469,In_775,In_485);
nand U470 (N_470,In_424,In_756);
or U471 (N_471,In_283,In_410);
or U472 (N_472,In_300,In_663);
nand U473 (N_473,In_672,In_892);
nand U474 (N_474,In_444,In_124);
and U475 (N_475,In_344,In_519);
nor U476 (N_476,In_47,In_998);
and U477 (N_477,In_681,In_64);
nand U478 (N_478,In_670,In_942);
xnor U479 (N_479,In_966,In_822);
nor U480 (N_480,In_330,In_632);
nand U481 (N_481,In_151,In_950);
xnor U482 (N_482,In_285,In_243);
or U483 (N_483,In_553,In_846);
or U484 (N_484,In_318,In_605);
xor U485 (N_485,In_659,In_418);
or U486 (N_486,In_593,In_196);
nor U487 (N_487,In_228,In_429);
xnor U488 (N_488,In_583,In_516);
nand U489 (N_489,In_3,In_773);
nand U490 (N_490,In_849,In_590);
and U491 (N_491,In_789,In_394);
or U492 (N_492,In_696,In_92);
and U493 (N_493,In_148,In_603);
xnor U494 (N_494,In_100,In_238);
nor U495 (N_495,In_524,In_619);
nand U496 (N_496,In_185,In_610);
and U497 (N_497,In_103,In_624);
or U498 (N_498,In_642,In_107);
and U499 (N_499,In_339,In_884);
and U500 (N_500,In_948,In_465);
or U501 (N_501,In_281,In_121);
and U502 (N_502,In_27,In_116);
nor U503 (N_503,In_550,In_997);
xor U504 (N_504,In_789,In_452);
or U505 (N_505,In_352,In_66);
and U506 (N_506,In_198,In_361);
or U507 (N_507,In_485,In_218);
nor U508 (N_508,In_272,In_240);
or U509 (N_509,In_926,In_132);
nor U510 (N_510,In_412,In_335);
nor U511 (N_511,In_566,In_381);
or U512 (N_512,In_922,In_654);
and U513 (N_513,In_531,In_280);
nor U514 (N_514,In_290,In_879);
nand U515 (N_515,In_553,In_467);
or U516 (N_516,In_767,In_423);
nor U517 (N_517,In_261,In_342);
and U518 (N_518,In_812,In_677);
or U519 (N_519,In_958,In_244);
xnor U520 (N_520,In_437,In_155);
xnor U521 (N_521,In_433,In_237);
xor U522 (N_522,In_121,In_671);
nand U523 (N_523,In_48,In_283);
nor U524 (N_524,In_432,In_672);
nand U525 (N_525,In_628,In_879);
xor U526 (N_526,In_854,In_401);
and U527 (N_527,In_822,In_608);
nand U528 (N_528,In_520,In_88);
or U529 (N_529,In_162,In_269);
nor U530 (N_530,In_998,In_266);
and U531 (N_531,In_468,In_191);
xor U532 (N_532,In_471,In_468);
and U533 (N_533,In_877,In_293);
xnor U534 (N_534,In_326,In_908);
nor U535 (N_535,In_491,In_457);
nor U536 (N_536,In_805,In_143);
or U537 (N_537,In_973,In_706);
xor U538 (N_538,In_821,In_776);
nor U539 (N_539,In_482,In_130);
nor U540 (N_540,In_162,In_135);
nand U541 (N_541,In_434,In_697);
xnor U542 (N_542,In_773,In_942);
nand U543 (N_543,In_987,In_598);
xnor U544 (N_544,In_126,In_496);
or U545 (N_545,In_239,In_974);
or U546 (N_546,In_70,In_804);
nor U547 (N_547,In_783,In_412);
nor U548 (N_548,In_320,In_497);
xor U549 (N_549,In_211,In_562);
nor U550 (N_550,In_494,In_529);
and U551 (N_551,In_600,In_278);
xnor U552 (N_552,In_15,In_734);
nor U553 (N_553,In_185,In_601);
and U554 (N_554,In_973,In_720);
nand U555 (N_555,In_927,In_890);
or U556 (N_556,In_71,In_840);
or U557 (N_557,In_277,In_92);
and U558 (N_558,In_610,In_846);
nor U559 (N_559,In_430,In_172);
nor U560 (N_560,In_957,In_820);
xnor U561 (N_561,In_640,In_142);
nor U562 (N_562,In_411,In_491);
and U563 (N_563,In_270,In_342);
or U564 (N_564,In_497,In_968);
or U565 (N_565,In_609,In_382);
and U566 (N_566,In_695,In_909);
and U567 (N_567,In_889,In_105);
nor U568 (N_568,In_675,In_783);
xor U569 (N_569,In_836,In_976);
and U570 (N_570,In_762,In_208);
and U571 (N_571,In_428,In_503);
or U572 (N_572,In_535,In_453);
or U573 (N_573,In_45,In_553);
nand U574 (N_574,In_850,In_347);
nor U575 (N_575,In_57,In_960);
nand U576 (N_576,In_892,In_687);
nand U577 (N_577,In_166,In_716);
xnor U578 (N_578,In_297,In_666);
xnor U579 (N_579,In_532,In_980);
and U580 (N_580,In_970,In_590);
xor U581 (N_581,In_124,In_451);
nand U582 (N_582,In_643,In_238);
nand U583 (N_583,In_139,In_218);
nor U584 (N_584,In_39,In_705);
and U585 (N_585,In_498,In_808);
nor U586 (N_586,In_316,In_368);
or U587 (N_587,In_756,In_771);
or U588 (N_588,In_669,In_763);
or U589 (N_589,In_23,In_114);
or U590 (N_590,In_746,In_132);
and U591 (N_591,In_34,In_468);
nand U592 (N_592,In_986,In_686);
nand U593 (N_593,In_669,In_524);
xnor U594 (N_594,In_504,In_892);
nor U595 (N_595,In_441,In_567);
xor U596 (N_596,In_679,In_765);
xor U597 (N_597,In_450,In_225);
and U598 (N_598,In_118,In_87);
or U599 (N_599,In_835,In_643);
nor U600 (N_600,In_825,In_528);
or U601 (N_601,In_326,In_391);
xnor U602 (N_602,In_28,In_521);
nor U603 (N_603,In_805,In_435);
xor U604 (N_604,In_884,In_618);
xor U605 (N_605,In_627,In_43);
xnor U606 (N_606,In_883,In_416);
nor U607 (N_607,In_910,In_16);
and U608 (N_608,In_46,In_177);
nand U609 (N_609,In_776,In_792);
nand U610 (N_610,In_223,In_749);
xor U611 (N_611,In_446,In_499);
nor U612 (N_612,In_58,In_126);
and U613 (N_613,In_347,In_58);
xnor U614 (N_614,In_16,In_322);
or U615 (N_615,In_741,In_434);
nor U616 (N_616,In_80,In_340);
xnor U617 (N_617,In_610,In_914);
or U618 (N_618,In_604,In_781);
or U619 (N_619,In_859,In_669);
xnor U620 (N_620,In_786,In_693);
nand U621 (N_621,In_345,In_249);
and U622 (N_622,In_300,In_673);
nand U623 (N_623,In_69,In_1);
nor U624 (N_624,In_171,In_581);
nor U625 (N_625,In_84,In_571);
nand U626 (N_626,In_254,In_526);
nor U627 (N_627,In_878,In_914);
nand U628 (N_628,In_115,In_361);
xor U629 (N_629,In_581,In_524);
or U630 (N_630,In_299,In_248);
xor U631 (N_631,In_615,In_976);
xor U632 (N_632,In_359,In_76);
and U633 (N_633,In_500,In_282);
or U634 (N_634,In_661,In_118);
nand U635 (N_635,In_63,In_922);
and U636 (N_636,In_459,In_68);
and U637 (N_637,In_441,In_306);
nor U638 (N_638,In_807,In_305);
nand U639 (N_639,In_154,In_564);
nor U640 (N_640,In_120,In_475);
nand U641 (N_641,In_722,In_935);
and U642 (N_642,In_102,In_963);
nand U643 (N_643,In_153,In_529);
nand U644 (N_644,In_998,In_121);
nor U645 (N_645,In_347,In_637);
nand U646 (N_646,In_335,In_959);
and U647 (N_647,In_537,In_436);
nor U648 (N_648,In_193,In_415);
nand U649 (N_649,In_511,In_333);
or U650 (N_650,In_459,In_528);
nand U651 (N_651,In_446,In_480);
and U652 (N_652,In_154,In_948);
and U653 (N_653,In_709,In_649);
nor U654 (N_654,In_978,In_678);
xnor U655 (N_655,In_710,In_695);
or U656 (N_656,In_603,In_382);
or U657 (N_657,In_152,In_623);
xor U658 (N_658,In_170,In_74);
xnor U659 (N_659,In_952,In_797);
xnor U660 (N_660,In_176,In_547);
or U661 (N_661,In_438,In_917);
or U662 (N_662,In_823,In_531);
nand U663 (N_663,In_844,In_910);
and U664 (N_664,In_904,In_395);
nor U665 (N_665,In_533,In_664);
nand U666 (N_666,In_107,In_212);
or U667 (N_667,In_984,In_580);
or U668 (N_668,In_141,In_289);
xnor U669 (N_669,In_776,In_298);
or U670 (N_670,In_725,In_52);
or U671 (N_671,In_705,In_195);
and U672 (N_672,In_983,In_40);
xor U673 (N_673,In_825,In_988);
and U674 (N_674,In_884,In_460);
or U675 (N_675,In_407,In_813);
nand U676 (N_676,In_960,In_988);
and U677 (N_677,In_660,In_519);
and U678 (N_678,In_519,In_839);
nand U679 (N_679,In_840,In_334);
xnor U680 (N_680,In_933,In_791);
and U681 (N_681,In_882,In_933);
nand U682 (N_682,In_896,In_198);
and U683 (N_683,In_610,In_519);
and U684 (N_684,In_612,In_931);
xnor U685 (N_685,In_158,In_182);
nor U686 (N_686,In_940,In_226);
or U687 (N_687,In_599,In_181);
nand U688 (N_688,In_542,In_740);
and U689 (N_689,In_306,In_34);
nand U690 (N_690,In_468,In_666);
xnor U691 (N_691,In_778,In_103);
nor U692 (N_692,In_876,In_911);
or U693 (N_693,In_665,In_36);
xnor U694 (N_694,In_467,In_713);
xnor U695 (N_695,In_801,In_417);
nand U696 (N_696,In_894,In_638);
or U697 (N_697,In_977,In_644);
nand U698 (N_698,In_269,In_881);
or U699 (N_699,In_182,In_570);
or U700 (N_700,In_460,In_937);
xnor U701 (N_701,In_764,In_352);
or U702 (N_702,In_407,In_229);
xor U703 (N_703,In_538,In_674);
nand U704 (N_704,In_294,In_234);
or U705 (N_705,In_626,In_75);
or U706 (N_706,In_998,In_174);
xnor U707 (N_707,In_206,In_326);
xnor U708 (N_708,In_224,In_363);
nor U709 (N_709,In_440,In_907);
xnor U710 (N_710,In_845,In_481);
or U711 (N_711,In_349,In_679);
or U712 (N_712,In_302,In_902);
or U713 (N_713,In_639,In_642);
xor U714 (N_714,In_952,In_193);
or U715 (N_715,In_194,In_825);
xnor U716 (N_716,In_521,In_534);
nand U717 (N_717,In_618,In_302);
or U718 (N_718,In_450,In_325);
nor U719 (N_719,In_191,In_562);
nand U720 (N_720,In_332,In_413);
or U721 (N_721,In_909,In_599);
nand U722 (N_722,In_791,In_0);
nand U723 (N_723,In_514,In_302);
and U724 (N_724,In_937,In_786);
or U725 (N_725,In_638,In_883);
and U726 (N_726,In_881,In_779);
or U727 (N_727,In_80,In_700);
xor U728 (N_728,In_339,In_142);
or U729 (N_729,In_418,In_923);
or U730 (N_730,In_625,In_411);
and U731 (N_731,In_840,In_195);
nand U732 (N_732,In_757,In_530);
nand U733 (N_733,In_109,In_965);
or U734 (N_734,In_990,In_669);
nand U735 (N_735,In_877,In_484);
nand U736 (N_736,In_251,In_102);
nand U737 (N_737,In_871,In_625);
and U738 (N_738,In_599,In_141);
nand U739 (N_739,In_288,In_835);
and U740 (N_740,In_101,In_904);
or U741 (N_741,In_923,In_534);
or U742 (N_742,In_405,In_626);
or U743 (N_743,In_244,In_489);
or U744 (N_744,In_72,In_597);
and U745 (N_745,In_615,In_734);
xnor U746 (N_746,In_388,In_387);
or U747 (N_747,In_7,In_841);
xor U748 (N_748,In_357,In_367);
nand U749 (N_749,In_237,In_513);
and U750 (N_750,In_452,In_214);
nor U751 (N_751,In_865,In_535);
or U752 (N_752,In_657,In_196);
nand U753 (N_753,In_955,In_927);
xor U754 (N_754,In_676,In_739);
xor U755 (N_755,In_620,In_640);
and U756 (N_756,In_228,In_242);
nor U757 (N_757,In_69,In_156);
or U758 (N_758,In_174,In_50);
or U759 (N_759,In_776,In_847);
nand U760 (N_760,In_64,In_373);
nor U761 (N_761,In_208,In_438);
nand U762 (N_762,In_435,In_254);
xor U763 (N_763,In_337,In_767);
and U764 (N_764,In_581,In_123);
nand U765 (N_765,In_3,In_319);
nor U766 (N_766,In_387,In_726);
or U767 (N_767,In_946,In_8);
nor U768 (N_768,In_437,In_482);
and U769 (N_769,In_801,In_50);
and U770 (N_770,In_934,In_996);
nand U771 (N_771,In_287,In_657);
nor U772 (N_772,In_462,In_576);
and U773 (N_773,In_244,In_250);
xnor U774 (N_774,In_647,In_802);
and U775 (N_775,In_884,In_833);
nor U776 (N_776,In_218,In_982);
nor U777 (N_777,In_283,In_359);
nand U778 (N_778,In_114,In_279);
and U779 (N_779,In_179,In_636);
nand U780 (N_780,In_351,In_910);
nand U781 (N_781,In_61,In_636);
and U782 (N_782,In_577,In_515);
xor U783 (N_783,In_389,In_729);
xor U784 (N_784,In_912,In_64);
nand U785 (N_785,In_771,In_246);
nand U786 (N_786,In_144,In_233);
xnor U787 (N_787,In_695,In_543);
nand U788 (N_788,In_26,In_210);
xor U789 (N_789,In_491,In_950);
nor U790 (N_790,In_522,In_555);
xor U791 (N_791,In_610,In_585);
or U792 (N_792,In_395,In_286);
and U793 (N_793,In_371,In_608);
or U794 (N_794,In_696,In_958);
or U795 (N_795,In_750,In_876);
xor U796 (N_796,In_268,In_400);
xor U797 (N_797,In_367,In_493);
xnor U798 (N_798,In_216,In_479);
nor U799 (N_799,In_118,In_72);
xnor U800 (N_800,In_941,In_281);
nand U801 (N_801,In_856,In_9);
nand U802 (N_802,In_754,In_971);
and U803 (N_803,In_662,In_840);
nand U804 (N_804,In_639,In_631);
nor U805 (N_805,In_212,In_472);
nand U806 (N_806,In_765,In_970);
nand U807 (N_807,In_286,In_701);
nand U808 (N_808,In_47,In_719);
or U809 (N_809,In_802,In_48);
xnor U810 (N_810,In_971,In_742);
xnor U811 (N_811,In_253,In_932);
nor U812 (N_812,In_305,In_632);
and U813 (N_813,In_596,In_761);
nand U814 (N_814,In_238,In_302);
nand U815 (N_815,In_531,In_402);
xor U816 (N_816,In_340,In_85);
nor U817 (N_817,In_290,In_91);
nor U818 (N_818,In_855,In_378);
xor U819 (N_819,In_457,In_817);
nand U820 (N_820,In_25,In_340);
and U821 (N_821,In_175,In_252);
or U822 (N_822,In_797,In_977);
or U823 (N_823,In_429,In_880);
nor U824 (N_824,In_394,In_437);
xor U825 (N_825,In_522,In_854);
and U826 (N_826,In_707,In_988);
xor U827 (N_827,In_73,In_372);
nand U828 (N_828,In_641,In_335);
nor U829 (N_829,In_381,In_169);
xnor U830 (N_830,In_450,In_706);
xor U831 (N_831,In_704,In_987);
and U832 (N_832,In_713,In_476);
nand U833 (N_833,In_21,In_427);
nor U834 (N_834,In_281,In_940);
xnor U835 (N_835,In_389,In_296);
xnor U836 (N_836,In_975,In_115);
xor U837 (N_837,In_285,In_728);
nand U838 (N_838,In_525,In_520);
nor U839 (N_839,In_938,In_505);
nor U840 (N_840,In_581,In_324);
and U841 (N_841,In_989,In_636);
and U842 (N_842,In_165,In_410);
and U843 (N_843,In_953,In_726);
xor U844 (N_844,In_98,In_138);
nor U845 (N_845,In_696,In_457);
xor U846 (N_846,In_595,In_806);
nor U847 (N_847,In_375,In_800);
xor U848 (N_848,In_166,In_884);
or U849 (N_849,In_361,In_878);
nand U850 (N_850,In_776,In_278);
xor U851 (N_851,In_259,In_645);
nor U852 (N_852,In_907,In_516);
and U853 (N_853,In_692,In_798);
nor U854 (N_854,In_548,In_993);
or U855 (N_855,In_954,In_222);
nor U856 (N_856,In_16,In_231);
and U857 (N_857,In_102,In_432);
or U858 (N_858,In_276,In_236);
and U859 (N_859,In_555,In_146);
and U860 (N_860,In_661,In_113);
xor U861 (N_861,In_375,In_871);
nor U862 (N_862,In_751,In_376);
xor U863 (N_863,In_83,In_1);
nor U864 (N_864,In_3,In_936);
and U865 (N_865,In_48,In_692);
and U866 (N_866,In_313,In_516);
or U867 (N_867,In_98,In_748);
nor U868 (N_868,In_312,In_481);
nand U869 (N_869,In_835,In_190);
nand U870 (N_870,In_3,In_638);
and U871 (N_871,In_148,In_200);
nand U872 (N_872,In_376,In_25);
nand U873 (N_873,In_957,In_352);
xor U874 (N_874,In_112,In_973);
nor U875 (N_875,In_803,In_828);
nor U876 (N_876,In_875,In_627);
nand U877 (N_877,In_244,In_61);
and U878 (N_878,In_295,In_102);
nand U879 (N_879,In_68,In_465);
xor U880 (N_880,In_98,In_996);
or U881 (N_881,In_408,In_368);
and U882 (N_882,In_118,In_286);
nor U883 (N_883,In_39,In_803);
nand U884 (N_884,In_496,In_597);
nand U885 (N_885,In_701,In_597);
or U886 (N_886,In_37,In_247);
xnor U887 (N_887,In_784,In_870);
or U888 (N_888,In_346,In_923);
nand U889 (N_889,In_916,In_984);
xnor U890 (N_890,In_652,In_40);
xnor U891 (N_891,In_812,In_517);
nor U892 (N_892,In_190,In_700);
and U893 (N_893,In_722,In_104);
nand U894 (N_894,In_927,In_275);
or U895 (N_895,In_954,In_815);
or U896 (N_896,In_66,In_272);
nor U897 (N_897,In_909,In_137);
nand U898 (N_898,In_731,In_610);
nand U899 (N_899,In_778,In_868);
and U900 (N_900,In_304,In_980);
nor U901 (N_901,In_171,In_723);
nor U902 (N_902,In_212,In_556);
and U903 (N_903,In_49,In_241);
and U904 (N_904,In_48,In_739);
nor U905 (N_905,In_280,In_650);
nor U906 (N_906,In_186,In_915);
nor U907 (N_907,In_69,In_367);
xor U908 (N_908,In_700,In_94);
nor U909 (N_909,In_593,In_826);
nand U910 (N_910,In_935,In_639);
nand U911 (N_911,In_502,In_571);
and U912 (N_912,In_523,In_385);
and U913 (N_913,In_166,In_639);
nand U914 (N_914,In_888,In_972);
xor U915 (N_915,In_794,In_375);
nor U916 (N_916,In_589,In_419);
nor U917 (N_917,In_31,In_971);
and U918 (N_918,In_62,In_980);
nor U919 (N_919,In_197,In_40);
and U920 (N_920,In_324,In_13);
and U921 (N_921,In_125,In_896);
or U922 (N_922,In_106,In_425);
nand U923 (N_923,In_436,In_437);
or U924 (N_924,In_67,In_121);
or U925 (N_925,In_168,In_670);
or U926 (N_926,In_340,In_317);
xnor U927 (N_927,In_364,In_181);
and U928 (N_928,In_30,In_242);
and U929 (N_929,In_337,In_338);
xnor U930 (N_930,In_105,In_761);
or U931 (N_931,In_677,In_427);
nand U932 (N_932,In_997,In_846);
nand U933 (N_933,In_599,In_555);
nor U934 (N_934,In_97,In_940);
nor U935 (N_935,In_893,In_534);
xor U936 (N_936,In_963,In_905);
nand U937 (N_937,In_894,In_916);
nor U938 (N_938,In_896,In_218);
xnor U939 (N_939,In_465,In_975);
nor U940 (N_940,In_606,In_663);
or U941 (N_941,In_126,In_130);
nor U942 (N_942,In_15,In_768);
nor U943 (N_943,In_627,In_106);
xnor U944 (N_944,In_661,In_935);
xor U945 (N_945,In_400,In_955);
nand U946 (N_946,In_208,In_962);
and U947 (N_947,In_354,In_257);
nor U948 (N_948,In_885,In_658);
or U949 (N_949,In_525,In_622);
nor U950 (N_950,In_228,In_921);
nor U951 (N_951,In_738,In_327);
or U952 (N_952,In_133,In_958);
xor U953 (N_953,In_293,In_792);
nor U954 (N_954,In_527,In_715);
nor U955 (N_955,In_48,In_369);
nand U956 (N_956,In_47,In_640);
and U957 (N_957,In_603,In_637);
nor U958 (N_958,In_850,In_707);
and U959 (N_959,In_866,In_78);
nand U960 (N_960,In_663,In_382);
or U961 (N_961,In_529,In_874);
xor U962 (N_962,In_178,In_132);
nor U963 (N_963,In_435,In_935);
nand U964 (N_964,In_841,In_288);
nor U965 (N_965,In_931,In_316);
nand U966 (N_966,In_389,In_52);
xnor U967 (N_967,In_458,In_431);
or U968 (N_968,In_298,In_903);
xor U969 (N_969,In_229,In_429);
xor U970 (N_970,In_584,In_578);
and U971 (N_971,In_152,In_131);
nor U972 (N_972,In_394,In_379);
and U973 (N_973,In_751,In_864);
nor U974 (N_974,In_737,In_191);
nand U975 (N_975,In_167,In_817);
nor U976 (N_976,In_638,In_785);
xor U977 (N_977,In_172,In_436);
nor U978 (N_978,In_736,In_24);
xor U979 (N_979,In_217,In_352);
xor U980 (N_980,In_717,In_194);
nor U981 (N_981,In_531,In_966);
nor U982 (N_982,In_335,In_534);
nor U983 (N_983,In_447,In_91);
or U984 (N_984,In_205,In_402);
nand U985 (N_985,In_786,In_105);
and U986 (N_986,In_282,In_45);
nor U987 (N_987,In_335,In_179);
or U988 (N_988,In_892,In_953);
xor U989 (N_989,In_792,In_107);
and U990 (N_990,In_770,In_227);
and U991 (N_991,In_203,In_778);
or U992 (N_992,In_839,In_978);
nor U993 (N_993,In_105,In_593);
nor U994 (N_994,In_627,In_85);
and U995 (N_995,In_89,In_280);
and U996 (N_996,In_298,In_593);
nor U997 (N_997,In_410,In_985);
and U998 (N_998,In_266,In_10);
nor U999 (N_999,In_721,In_399);
nor U1000 (N_1000,In_871,In_809);
or U1001 (N_1001,In_281,In_310);
and U1002 (N_1002,In_336,In_833);
nand U1003 (N_1003,In_140,In_313);
or U1004 (N_1004,In_377,In_326);
and U1005 (N_1005,In_587,In_851);
nand U1006 (N_1006,In_894,In_35);
nand U1007 (N_1007,In_22,In_662);
nand U1008 (N_1008,In_153,In_473);
nor U1009 (N_1009,In_959,In_697);
xor U1010 (N_1010,In_62,In_12);
nand U1011 (N_1011,In_744,In_260);
or U1012 (N_1012,In_796,In_495);
xor U1013 (N_1013,In_103,In_994);
nor U1014 (N_1014,In_935,In_524);
xnor U1015 (N_1015,In_129,In_337);
nand U1016 (N_1016,In_578,In_529);
or U1017 (N_1017,In_357,In_710);
nand U1018 (N_1018,In_524,In_756);
xor U1019 (N_1019,In_90,In_1);
and U1020 (N_1020,In_797,In_305);
xnor U1021 (N_1021,In_649,In_555);
or U1022 (N_1022,In_283,In_794);
and U1023 (N_1023,In_565,In_668);
nor U1024 (N_1024,In_367,In_447);
or U1025 (N_1025,In_100,In_170);
nand U1026 (N_1026,In_105,In_205);
nor U1027 (N_1027,In_56,In_634);
nor U1028 (N_1028,In_66,In_473);
or U1029 (N_1029,In_383,In_188);
or U1030 (N_1030,In_689,In_631);
xor U1031 (N_1031,In_517,In_318);
xnor U1032 (N_1032,In_884,In_235);
nor U1033 (N_1033,In_440,In_479);
nand U1034 (N_1034,In_395,In_696);
nand U1035 (N_1035,In_888,In_644);
or U1036 (N_1036,In_710,In_953);
and U1037 (N_1037,In_284,In_346);
nor U1038 (N_1038,In_627,In_920);
xor U1039 (N_1039,In_994,In_381);
and U1040 (N_1040,In_123,In_829);
and U1041 (N_1041,In_582,In_698);
or U1042 (N_1042,In_291,In_222);
and U1043 (N_1043,In_925,In_473);
xnor U1044 (N_1044,In_799,In_615);
or U1045 (N_1045,In_285,In_468);
or U1046 (N_1046,In_85,In_407);
nand U1047 (N_1047,In_612,In_722);
nand U1048 (N_1048,In_58,In_893);
nand U1049 (N_1049,In_134,In_318);
nor U1050 (N_1050,In_846,In_54);
nand U1051 (N_1051,In_464,In_263);
xor U1052 (N_1052,In_787,In_950);
and U1053 (N_1053,In_977,In_570);
nand U1054 (N_1054,In_464,In_748);
nor U1055 (N_1055,In_243,In_177);
nand U1056 (N_1056,In_300,In_454);
nor U1057 (N_1057,In_919,In_580);
or U1058 (N_1058,In_279,In_272);
nor U1059 (N_1059,In_745,In_415);
and U1060 (N_1060,In_397,In_925);
nor U1061 (N_1061,In_15,In_345);
nand U1062 (N_1062,In_335,In_514);
xnor U1063 (N_1063,In_74,In_884);
xnor U1064 (N_1064,In_959,In_29);
nand U1065 (N_1065,In_995,In_955);
or U1066 (N_1066,In_263,In_468);
xnor U1067 (N_1067,In_299,In_530);
nand U1068 (N_1068,In_352,In_554);
or U1069 (N_1069,In_484,In_79);
nand U1070 (N_1070,In_107,In_647);
or U1071 (N_1071,In_319,In_196);
nand U1072 (N_1072,In_68,In_394);
xor U1073 (N_1073,In_388,In_477);
or U1074 (N_1074,In_758,In_85);
or U1075 (N_1075,In_798,In_586);
nand U1076 (N_1076,In_514,In_220);
or U1077 (N_1077,In_777,In_338);
xnor U1078 (N_1078,In_581,In_907);
nand U1079 (N_1079,In_624,In_512);
nand U1080 (N_1080,In_84,In_432);
nand U1081 (N_1081,In_733,In_446);
xor U1082 (N_1082,In_751,In_35);
nor U1083 (N_1083,In_133,In_971);
xor U1084 (N_1084,In_60,In_698);
xnor U1085 (N_1085,In_372,In_747);
and U1086 (N_1086,In_420,In_464);
xnor U1087 (N_1087,In_928,In_917);
and U1088 (N_1088,In_8,In_894);
xor U1089 (N_1089,In_985,In_729);
and U1090 (N_1090,In_756,In_227);
and U1091 (N_1091,In_108,In_231);
and U1092 (N_1092,In_170,In_388);
xor U1093 (N_1093,In_329,In_655);
nand U1094 (N_1094,In_519,In_597);
xnor U1095 (N_1095,In_312,In_633);
nand U1096 (N_1096,In_317,In_48);
or U1097 (N_1097,In_792,In_458);
nor U1098 (N_1098,In_840,In_564);
xor U1099 (N_1099,In_25,In_162);
xor U1100 (N_1100,In_631,In_585);
nand U1101 (N_1101,In_273,In_665);
nand U1102 (N_1102,In_111,In_724);
nor U1103 (N_1103,In_688,In_146);
or U1104 (N_1104,In_722,In_526);
or U1105 (N_1105,In_307,In_892);
nand U1106 (N_1106,In_475,In_347);
nand U1107 (N_1107,In_579,In_190);
or U1108 (N_1108,In_344,In_656);
nand U1109 (N_1109,In_522,In_749);
nand U1110 (N_1110,In_597,In_554);
nand U1111 (N_1111,In_264,In_817);
nand U1112 (N_1112,In_845,In_867);
nand U1113 (N_1113,In_881,In_196);
and U1114 (N_1114,In_356,In_402);
and U1115 (N_1115,In_144,In_898);
nand U1116 (N_1116,In_66,In_549);
and U1117 (N_1117,In_637,In_420);
nand U1118 (N_1118,In_405,In_934);
or U1119 (N_1119,In_473,In_671);
nand U1120 (N_1120,In_65,In_955);
or U1121 (N_1121,In_270,In_19);
and U1122 (N_1122,In_743,In_672);
nand U1123 (N_1123,In_105,In_878);
and U1124 (N_1124,In_770,In_776);
or U1125 (N_1125,In_410,In_532);
nand U1126 (N_1126,In_790,In_850);
and U1127 (N_1127,In_180,In_564);
xor U1128 (N_1128,In_909,In_862);
or U1129 (N_1129,In_756,In_715);
or U1130 (N_1130,In_520,In_138);
or U1131 (N_1131,In_375,In_487);
nand U1132 (N_1132,In_112,In_484);
nor U1133 (N_1133,In_893,In_611);
nor U1134 (N_1134,In_153,In_34);
xnor U1135 (N_1135,In_743,In_903);
nand U1136 (N_1136,In_960,In_118);
and U1137 (N_1137,In_654,In_255);
and U1138 (N_1138,In_820,In_101);
nand U1139 (N_1139,In_358,In_826);
or U1140 (N_1140,In_947,In_638);
or U1141 (N_1141,In_143,In_885);
nor U1142 (N_1142,In_944,In_470);
nor U1143 (N_1143,In_678,In_487);
or U1144 (N_1144,In_880,In_839);
nand U1145 (N_1145,In_645,In_400);
nor U1146 (N_1146,In_409,In_735);
nand U1147 (N_1147,In_302,In_337);
nand U1148 (N_1148,In_721,In_365);
nor U1149 (N_1149,In_53,In_400);
or U1150 (N_1150,In_290,In_550);
and U1151 (N_1151,In_396,In_869);
nor U1152 (N_1152,In_335,In_852);
nand U1153 (N_1153,In_775,In_955);
xnor U1154 (N_1154,In_124,In_890);
xor U1155 (N_1155,In_971,In_678);
nor U1156 (N_1156,In_459,In_877);
or U1157 (N_1157,In_163,In_631);
nor U1158 (N_1158,In_527,In_953);
or U1159 (N_1159,In_225,In_2);
nor U1160 (N_1160,In_794,In_588);
or U1161 (N_1161,In_608,In_228);
or U1162 (N_1162,In_151,In_829);
nor U1163 (N_1163,In_621,In_287);
or U1164 (N_1164,In_108,In_545);
xnor U1165 (N_1165,In_298,In_564);
nand U1166 (N_1166,In_159,In_948);
and U1167 (N_1167,In_213,In_553);
or U1168 (N_1168,In_148,In_747);
and U1169 (N_1169,In_235,In_610);
nand U1170 (N_1170,In_506,In_851);
nor U1171 (N_1171,In_526,In_249);
or U1172 (N_1172,In_33,In_953);
and U1173 (N_1173,In_416,In_228);
nand U1174 (N_1174,In_960,In_880);
nand U1175 (N_1175,In_52,In_938);
nor U1176 (N_1176,In_16,In_353);
and U1177 (N_1177,In_894,In_980);
and U1178 (N_1178,In_356,In_81);
or U1179 (N_1179,In_548,In_834);
and U1180 (N_1180,In_465,In_664);
and U1181 (N_1181,In_465,In_871);
or U1182 (N_1182,In_938,In_971);
nor U1183 (N_1183,In_294,In_59);
or U1184 (N_1184,In_604,In_189);
nor U1185 (N_1185,In_423,In_960);
nor U1186 (N_1186,In_387,In_589);
and U1187 (N_1187,In_576,In_77);
and U1188 (N_1188,In_513,In_366);
and U1189 (N_1189,In_512,In_433);
and U1190 (N_1190,In_938,In_984);
nand U1191 (N_1191,In_993,In_78);
or U1192 (N_1192,In_425,In_281);
nand U1193 (N_1193,In_807,In_662);
or U1194 (N_1194,In_245,In_67);
and U1195 (N_1195,In_603,In_445);
or U1196 (N_1196,In_166,In_323);
and U1197 (N_1197,In_49,In_14);
nand U1198 (N_1198,In_245,In_138);
and U1199 (N_1199,In_744,In_964);
and U1200 (N_1200,In_969,In_873);
nand U1201 (N_1201,In_828,In_471);
nand U1202 (N_1202,In_849,In_536);
xor U1203 (N_1203,In_122,In_805);
nand U1204 (N_1204,In_616,In_334);
xnor U1205 (N_1205,In_67,In_140);
nor U1206 (N_1206,In_462,In_84);
or U1207 (N_1207,In_73,In_283);
nand U1208 (N_1208,In_770,In_643);
nor U1209 (N_1209,In_155,In_369);
xor U1210 (N_1210,In_241,In_472);
nand U1211 (N_1211,In_261,In_358);
nor U1212 (N_1212,In_427,In_844);
xnor U1213 (N_1213,In_962,In_885);
nand U1214 (N_1214,In_58,In_438);
xor U1215 (N_1215,In_899,In_983);
and U1216 (N_1216,In_250,In_491);
nand U1217 (N_1217,In_889,In_30);
or U1218 (N_1218,In_891,In_359);
nand U1219 (N_1219,In_559,In_540);
nand U1220 (N_1220,In_456,In_354);
or U1221 (N_1221,In_503,In_736);
or U1222 (N_1222,In_490,In_397);
xnor U1223 (N_1223,In_809,In_684);
nor U1224 (N_1224,In_385,In_312);
or U1225 (N_1225,In_831,In_479);
nor U1226 (N_1226,In_375,In_973);
or U1227 (N_1227,In_384,In_580);
xnor U1228 (N_1228,In_644,In_251);
nor U1229 (N_1229,In_199,In_476);
xor U1230 (N_1230,In_978,In_282);
nor U1231 (N_1231,In_731,In_751);
nor U1232 (N_1232,In_174,In_361);
nor U1233 (N_1233,In_59,In_900);
xor U1234 (N_1234,In_453,In_968);
nand U1235 (N_1235,In_484,In_646);
nor U1236 (N_1236,In_569,In_360);
nand U1237 (N_1237,In_156,In_267);
and U1238 (N_1238,In_151,In_226);
xor U1239 (N_1239,In_840,In_328);
or U1240 (N_1240,In_905,In_367);
nor U1241 (N_1241,In_989,In_621);
xor U1242 (N_1242,In_302,In_994);
nand U1243 (N_1243,In_268,In_961);
and U1244 (N_1244,In_358,In_809);
or U1245 (N_1245,In_516,In_185);
and U1246 (N_1246,In_362,In_74);
nand U1247 (N_1247,In_514,In_773);
nand U1248 (N_1248,In_626,In_98);
nand U1249 (N_1249,In_426,In_207);
xor U1250 (N_1250,In_398,In_821);
or U1251 (N_1251,In_598,In_756);
nor U1252 (N_1252,In_279,In_328);
xnor U1253 (N_1253,In_964,In_222);
xor U1254 (N_1254,In_845,In_814);
or U1255 (N_1255,In_684,In_284);
and U1256 (N_1256,In_793,In_458);
nor U1257 (N_1257,In_277,In_84);
nor U1258 (N_1258,In_609,In_736);
nor U1259 (N_1259,In_762,In_678);
nand U1260 (N_1260,In_358,In_394);
xnor U1261 (N_1261,In_449,In_679);
or U1262 (N_1262,In_224,In_335);
or U1263 (N_1263,In_803,In_600);
xnor U1264 (N_1264,In_910,In_740);
nor U1265 (N_1265,In_96,In_678);
nor U1266 (N_1266,In_127,In_254);
nor U1267 (N_1267,In_10,In_509);
or U1268 (N_1268,In_63,In_750);
nand U1269 (N_1269,In_631,In_819);
xor U1270 (N_1270,In_562,In_434);
nor U1271 (N_1271,In_665,In_431);
nand U1272 (N_1272,In_93,In_490);
nor U1273 (N_1273,In_336,In_498);
and U1274 (N_1274,In_600,In_775);
and U1275 (N_1275,In_753,In_230);
or U1276 (N_1276,In_497,In_404);
and U1277 (N_1277,In_632,In_967);
and U1278 (N_1278,In_721,In_111);
xor U1279 (N_1279,In_420,In_121);
xnor U1280 (N_1280,In_654,In_992);
and U1281 (N_1281,In_907,In_108);
nor U1282 (N_1282,In_263,In_283);
nand U1283 (N_1283,In_909,In_882);
nor U1284 (N_1284,In_240,In_503);
or U1285 (N_1285,In_182,In_232);
xnor U1286 (N_1286,In_829,In_477);
or U1287 (N_1287,In_632,In_846);
or U1288 (N_1288,In_29,In_104);
nand U1289 (N_1289,In_555,In_420);
or U1290 (N_1290,In_605,In_114);
nor U1291 (N_1291,In_724,In_304);
nor U1292 (N_1292,In_941,In_411);
nand U1293 (N_1293,In_496,In_282);
or U1294 (N_1294,In_232,In_673);
nand U1295 (N_1295,In_618,In_565);
and U1296 (N_1296,In_801,In_414);
nand U1297 (N_1297,In_905,In_547);
nand U1298 (N_1298,In_337,In_996);
nor U1299 (N_1299,In_568,In_41);
nand U1300 (N_1300,In_594,In_732);
and U1301 (N_1301,In_190,In_472);
nand U1302 (N_1302,In_878,In_646);
xor U1303 (N_1303,In_779,In_367);
nor U1304 (N_1304,In_373,In_950);
nand U1305 (N_1305,In_916,In_849);
nor U1306 (N_1306,In_616,In_967);
or U1307 (N_1307,In_23,In_722);
nand U1308 (N_1308,In_306,In_72);
nand U1309 (N_1309,In_793,In_935);
or U1310 (N_1310,In_152,In_474);
nor U1311 (N_1311,In_204,In_911);
and U1312 (N_1312,In_98,In_152);
nor U1313 (N_1313,In_962,In_914);
or U1314 (N_1314,In_773,In_483);
or U1315 (N_1315,In_246,In_195);
xor U1316 (N_1316,In_245,In_762);
nand U1317 (N_1317,In_996,In_715);
and U1318 (N_1318,In_393,In_535);
nor U1319 (N_1319,In_824,In_700);
and U1320 (N_1320,In_435,In_249);
nor U1321 (N_1321,In_595,In_724);
nand U1322 (N_1322,In_307,In_656);
nor U1323 (N_1323,In_737,In_232);
nand U1324 (N_1324,In_748,In_266);
or U1325 (N_1325,In_35,In_771);
or U1326 (N_1326,In_784,In_623);
nand U1327 (N_1327,In_74,In_444);
or U1328 (N_1328,In_146,In_27);
or U1329 (N_1329,In_296,In_460);
and U1330 (N_1330,In_625,In_174);
or U1331 (N_1331,In_185,In_704);
xnor U1332 (N_1332,In_797,In_264);
xor U1333 (N_1333,In_970,In_773);
nand U1334 (N_1334,In_980,In_963);
nand U1335 (N_1335,In_681,In_527);
nor U1336 (N_1336,In_552,In_987);
xor U1337 (N_1337,In_69,In_901);
and U1338 (N_1338,In_930,In_744);
and U1339 (N_1339,In_843,In_725);
nand U1340 (N_1340,In_437,In_140);
or U1341 (N_1341,In_6,In_794);
and U1342 (N_1342,In_141,In_222);
nor U1343 (N_1343,In_78,In_535);
nand U1344 (N_1344,In_329,In_105);
or U1345 (N_1345,In_756,In_881);
nand U1346 (N_1346,In_664,In_998);
xnor U1347 (N_1347,In_626,In_779);
and U1348 (N_1348,In_707,In_948);
and U1349 (N_1349,In_958,In_28);
and U1350 (N_1350,In_51,In_440);
nor U1351 (N_1351,In_585,In_656);
nand U1352 (N_1352,In_926,In_96);
nor U1353 (N_1353,In_109,In_542);
nand U1354 (N_1354,In_419,In_204);
xnor U1355 (N_1355,In_108,In_490);
and U1356 (N_1356,In_601,In_21);
xor U1357 (N_1357,In_850,In_145);
nor U1358 (N_1358,In_923,In_809);
xnor U1359 (N_1359,In_719,In_908);
nor U1360 (N_1360,In_563,In_595);
or U1361 (N_1361,In_159,In_695);
xnor U1362 (N_1362,In_136,In_73);
xor U1363 (N_1363,In_296,In_986);
nand U1364 (N_1364,In_56,In_115);
and U1365 (N_1365,In_306,In_802);
xnor U1366 (N_1366,In_906,In_602);
and U1367 (N_1367,In_950,In_908);
xor U1368 (N_1368,In_621,In_346);
or U1369 (N_1369,In_485,In_536);
nand U1370 (N_1370,In_428,In_692);
and U1371 (N_1371,In_344,In_936);
nor U1372 (N_1372,In_769,In_8);
or U1373 (N_1373,In_333,In_889);
nand U1374 (N_1374,In_118,In_389);
and U1375 (N_1375,In_873,In_960);
xnor U1376 (N_1376,In_597,In_720);
nor U1377 (N_1377,In_768,In_691);
and U1378 (N_1378,In_68,In_411);
nor U1379 (N_1379,In_299,In_561);
nand U1380 (N_1380,In_995,In_11);
nand U1381 (N_1381,In_597,In_286);
xor U1382 (N_1382,In_342,In_900);
nand U1383 (N_1383,In_760,In_67);
xnor U1384 (N_1384,In_340,In_717);
and U1385 (N_1385,In_999,In_555);
or U1386 (N_1386,In_202,In_860);
nor U1387 (N_1387,In_676,In_407);
or U1388 (N_1388,In_61,In_956);
nand U1389 (N_1389,In_858,In_492);
xnor U1390 (N_1390,In_381,In_231);
nor U1391 (N_1391,In_559,In_772);
nand U1392 (N_1392,In_374,In_452);
and U1393 (N_1393,In_419,In_2);
or U1394 (N_1394,In_527,In_307);
xnor U1395 (N_1395,In_257,In_921);
xnor U1396 (N_1396,In_707,In_296);
and U1397 (N_1397,In_621,In_549);
and U1398 (N_1398,In_228,In_32);
nor U1399 (N_1399,In_419,In_216);
nor U1400 (N_1400,In_219,In_878);
and U1401 (N_1401,In_48,In_543);
or U1402 (N_1402,In_167,In_36);
nor U1403 (N_1403,In_9,In_224);
xnor U1404 (N_1404,In_407,In_809);
nand U1405 (N_1405,In_985,In_774);
xor U1406 (N_1406,In_441,In_193);
and U1407 (N_1407,In_709,In_625);
nor U1408 (N_1408,In_77,In_934);
nor U1409 (N_1409,In_459,In_876);
nand U1410 (N_1410,In_44,In_820);
nand U1411 (N_1411,In_348,In_435);
nor U1412 (N_1412,In_696,In_382);
or U1413 (N_1413,In_413,In_495);
and U1414 (N_1414,In_799,In_777);
nand U1415 (N_1415,In_108,In_719);
xor U1416 (N_1416,In_439,In_873);
nand U1417 (N_1417,In_398,In_859);
and U1418 (N_1418,In_821,In_580);
xor U1419 (N_1419,In_523,In_791);
nor U1420 (N_1420,In_700,In_860);
and U1421 (N_1421,In_988,In_853);
xnor U1422 (N_1422,In_209,In_473);
or U1423 (N_1423,In_545,In_930);
and U1424 (N_1424,In_706,In_312);
nor U1425 (N_1425,In_847,In_881);
xnor U1426 (N_1426,In_74,In_718);
nand U1427 (N_1427,In_609,In_386);
nor U1428 (N_1428,In_865,In_544);
and U1429 (N_1429,In_649,In_827);
nor U1430 (N_1430,In_451,In_505);
nand U1431 (N_1431,In_59,In_550);
nor U1432 (N_1432,In_311,In_453);
or U1433 (N_1433,In_375,In_98);
nor U1434 (N_1434,In_435,In_452);
nand U1435 (N_1435,In_870,In_766);
and U1436 (N_1436,In_348,In_68);
and U1437 (N_1437,In_870,In_445);
or U1438 (N_1438,In_808,In_13);
or U1439 (N_1439,In_129,In_522);
xor U1440 (N_1440,In_286,In_379);
or U1441 (N_1441,In_45,In_734);
nor U1442 (N_1442,In_140,In_887);
nand U1443 (N_1443,In_161,In_492);
nor U1444 (N_1444,In_719,In_364);
nand U1445 (N_1445,In_546,In_528);
and U1446 (N_1446,In_796,In_251);
or U1447 (N_1447,In_349,In_637);
nand U1448 (N_1448,In_939,In_729);
or U1449 (N_1449,In_788,In_594);
or U1450 (N_1450,In_604,In_830);
and U1451 (N_1451,In_3,In_78);
and U1452 (N_1452,In_967,In_307);
nor U1453 (N_1453,In_717,In_302);
xor U1454 (N_1454,In_431,In_255);
nor U1455 (N_1455,In_725,In_25);
nor U1456 (N_1456,In_17,In_927);
xor U1457 (N_1457,In_954,In_532);
nor U1458 (N_1458,In_269,In_70);
xnor U1459 (N_1459,In_867,In_274);
and U1460 (N_1460,In_685,In_282);
nor U1461 (N_1461,In_767,In_412);
and U1462 (N_1462,In_808,In_797);
xnor U1463 (N_1463,In_862,In_543);
nor U1464 (N_1464,In_195,In_677);
and U1465 (N_1465,In_96,In_960);
nor U1466 (N_1466,In_77,In_134);
xnor U1467 (N_1467,In_906,In_804);
xor U1468 (N_1468,In_216,In_741);
nand U1469 (N_1469,In_676,In_370);
and U1470 (N_1470,In_254,In_181);
nor U1471 (N_1471,In_115,In_870);
or U1472 (N_1472,In_481,In_275);
nor U1473 (N_1473,In_209,In_93);
xnor U1474 (N_1474,In_738,In_387);
or U1475 (N_1475,In_979,In_184);
and U1476 (N_1476,In_82,In_819);
or U1477 (N_1477,In_954,In_799);
and U1478 (N_1478,In_614,In_833);
nand U1479 (N_1479,In_554,In_515);
nor U1480 (N_1480,In_129,In_475);
and U1481 (N_1481,In_815,In_715);
nor U1482 (N_1482,In_834,In_496);
or U1483 (N_1483,In_120,In_809);
xor U1484 (N_1484,In_569,In_295);
nand U1485 (N_1485,In_920,In_967);
or U1486 (N_1486,In_39,In_176);
nor U1487 (N_1487,In_349,In_588);
nor U1488 (N_1488,In_186,In_773);
nor U1489 (N_1489,In_327,In_259);
and U1490 (N_1490,In_925,In_144);
nand U1491 (N_1491,In_795,In_513);
nand U1492 (N_1492,In_437,In_148);
xor U1493 (N_1493,In_699,In_325);
and U1494 (N_1494,In_25,In_749);
nor U1495 (N_1495,In_57,In_730);
or U1496 (N_1496,In_537,In_751);
nor U1497 (N_1497,In_807,In_704);
nand U1498 (N_1498,In_973,In_656);
nand U1499 (N_1499,In_203,In_498);
nand U1500 (N_1500,In_705,In_884);
and U1501 (N_1501,In_17,In_187);
nor U1502 (N_1502,In_141,In_735);
and U1503 (N_1503,In_322,In_258);
nor U1504 (N_1504,In_352,In_628);
and U1505 (N_1505,In_194,In_862);
xnor U1506 (N_1506,In_375,In_111);
and U1507 (N_1507,In_528,In_238);
or U1508 (N_1508,In_949,In_620);
or U1509 (N_1509,In_48,In_881);
or U1510 (N_1510,In_440,In_850);
xor U1511 (N_1511,In_502,In_607);
or U1512 (N_1512,In_668,In_523);
or U1513 (N_1513,In_582,In_263);
nand U1514 (N_1514,In_771,In_305);
xor U1515 (N_1515,In_10,In_254);
xnor U1516 (N_1516,In_944,In_549);
nor U1517 (N_1517,In_653,In_44);
and U1518 (N_1518,In_193,In_976);
nor U1519 (N_1519,In_833,In_852);
or U1520 (N_1520,In_62,In_994);
or U1521 (N_1521,In_992,In_60);
nand U1522 (N_1522,In_670,In_680);
xor U1523 (N_1523,In_475,In_232);
xnor U1524 (N_1524,In_409,In_266);
nor U1525 (N_1525,In_798,In_874);
nor U1526 (N_1526,In_636,In_135);
xor U1527 (N_1527,In_261,In_678);
nor U1528 (N_1528,In_182,In_824);
or U1529 (N_1529,In_999,In_459);
xor U1530 (N_1530,In_589,In_422);
xor U1531 (N_1531,In_640,In_323);
nor U1532 (N_1532,In_491,In_472);
nand U1533 (N_1533,In_506,In_16);
xor U1534 (N_1534,In_462,In_774);
or U1535 (N_1535,In_349,In_327);
xnor U1536 (N_1536,In_956,In_631);
or U1537 (N_1537,In_512,In_859);
xor U1538 (N_1538,In_938,In_899);
xnor U1539 (N_1539,In_191,In_621);
nor U1540 (N_1540,In_977,In_694);
nand U1541 (N_1541,In_301,In_800);
or U1542 (N_1542,In_127,In_152);
nand U1543 (N_1543,In_314,In_247);
xor U1544 (N_1544,In_164,In_724);
and U1545 (N_1545,In_190,In_635);
xnor U1546 (N_1546,In_263,In_246);
or U1547 (N_1547,In_633,In_301);
or U1548 (N_1548,In_621,In_335);
nand U1549 (N_1549,In_511,In_414);
nor U1550 (N_1550,In_88,In_480);
nor U1551 (N_1551,In_382,In_135);
nor U1552 (N_1552,In_581,In_255);
and U1553 (N_1553,In_535,In_722);
xor U1554 (N_1554,In_304,In_67);
or U1555 (N_1555,In_578,In_362);
nor U1556 (N_1556,In_459,In_307);
nor U1557 (N_1557,In_13,In_292);
or U1558 (N_1558,In_420,In_191);
nand U1559 (N_1559,In_70,In_17);
nor U1560 (N_1560,In_359,In_219);
nor U1561 (N_1561,In_842,In_279);
and U1562 (N_1562,In_490,In_710);
nand U1563 (N_1563,In_327,In_392);
xnor U1564 (N_1564,In_221,In_94);
nand U1565 (N_1565,In_112,In_705);
and U1566 (N_1566,In_537,In_273);
nand U1567 (N_1567,In_646,In_711);
nand U1568 (N_1568,In_481,In_107);
nor U1569 (N_1569,In_667,In_590);
xnor U1570 (N_1570,In_596,In_937);
and U1571 (N_1571,In_65,In_152);
nand U1572 (N_1572,In_951,In_226);
or U1573 (N_1573,In_448,In_377);
nor U1574 (N_1574,In_810,In_543);
and U1575 (N_1575,In_986,In_309);
xor U1576 (N_1576,In_698,In_330);
nor U1577 (N_1577,In_56,In_357);
xor U1578 (N_1578,In_994,In_377);
xor U1579 (N_1579,In_492,In_390);
xnor U1580 (N_1580,In_497,In_66);
nor U1581 (N_1581,In_575,In_887);
nor U1582 (N_1582,In_260,In_629);
nand U1583 (N_1583,In_138,In_19);
xor U1584 (N_1584,In_416,In_256);
and U1585 (N_1585,In_266,In_834);
or U1586 (N_1586,In_761,In_734);
nor U1587 (N_1587,In_671,In_639);
or U1588 (N_1588,In_8,In_902);
and U1589 (N_1589,In_818,In_219);
nor U1590 (N_1590,In_664,In_669);
or U1591 (N_1591,In_366,In_40);
xor U1592 (N_1592,In_513,In_857);
and U1593 (N_1593,In_383,In_215);
nor U1594 (N_1594,In_863,In_782);
xor U1595 (N_1595,In_253,In_721);
and U1596 (N_1596,In_681,In_25);
nand U1597 (N_1597,In_28,In_45);
nor U1598 (N_1598,In_112,In_811);
nand U1599 (N_1599,In_184,In_400);
xnor U1600 (N_1600,In_658,In_482);
nand U1601 (N_1601,In_490,In_653);
nand U1602 (N_1602,In_170,In_437);
nand U1603 (N_1603,In_807,In_872);
and U1604 (N_1604,In_759,In_322);
or U1605 (N_1605,In_398,In_491);
xnor U1606 (N_1606,In_510,In_827);
nor U1607 (N_1607,In_524,In_376);
and U1608 (N_1608,In_895,In_980);
nor U1609 (N_1609,In_996,In_534);
nand U1610 (N_1610,In_113,In_29);
or U1611 (N_1611,In_749,In_635);
nand U1612 (N_1612,In_261,In_15);
or U1613 (N_1613,In_869,In_84);
and U1614 (N_1614,In_319,In_501);
nor U1615 (N_1615,In_178,In_264);
nand U1616 (N_1616,In_268,In_38);
xnor U1617 (N_1617,In_891,In_830);
and U1618 (N_1618,In_583,In_327);
or U1619 (N_1619,In_834,In_970);
nor U1620 (N_1620,In_499,In_716);
xnor U1621 (N_1621,In_964,In_196);
nor U1622 (N_1622,In_309,In_481);
nor U1623 (N_1623,In_581,In_191);
or U1624 (N_1624,In_516,In_631);
and U1625 (N_1625,In_678,In_93);
or U1626 (N_1626,In_307,In_709);
or U1627 (N_1627,In_479,In_435);
xor U1628 (N_1628,In_637,In_865);
or U1629 (N_1629,In_568,In_320);
and U1630 (N_1630,In_903,In_670);
xor U1631 (N_1631,In_651,In_18);
xnor U1632 (N_1632,In_411,In_25);
nand U1633 (N_1633,In_723,In_606);
nor U1634 (N_1634,In_104,In_788);
or U1635 (N_1635,In_456,In_128);
or U1636 (N_1636,In_594,In_815);
or U1637 (N_1637,In_43,In_788);
nor U1638 (N_1638,In_487,In_626);
or U1639 (N_1639,In_845,In_246);
xnor U1640 (N_1640,In_33,In_694);
nand U1641 (N_1641,In_52,In_754);
and U1642 (N_1642,In_586,In_422);
or U1643 (N_1643,In_619,In_748);
nor U1644 (N_1644,In_588,In_188);
nand U1645 (N_1645,In_362,In_37);
xor U1646 (N_1646,In_742,In_679);
or U1647 (N_1647,In_721,In_933);
nor U1648 (N_1648,In_304,In_489);
and U1649 (N_1649,In_645,In_459);
or U1650 (N_1650,In_17,In_212);
and U1651 (N_1651,In_172,In_924);
and U1652 (N_1652,In_166,In_814);
nor U1653 (N_1653,In_967,In_473);
xor U1654 (N_1654,In_413,In_684);
and U1655 (N_1655,In_581,In_19);
nor U1656 (N_1656,In_415,In_741);
or U1657 (N_1657,In_334,In_359);
nand U1658 (N_1658,In_66,In_452);
nand U1659 (N_1659,In_268,In_788);
xor U1660 (N_1660,In_281,In_957);
nand U1661 (N_1661,In_373,In_46);
nand U1662 (N_1662,In_291,In_665);
nor U1663 (N_1663,In_665,In_225);
nand U1664 (N_1664,In_202,In_32);
and U1665 (N_1665,In_817,In_7);
nor U1666 (N_1666,In_205,In_206);
nand U1667 (N_1667,In_237,In_267);
and U1668 (N_1668,In_631,In_739);
nor U1669 (N_1669,In_906,In_51);
xor U1670 (N_1670,In_951,In_605);
nor U1671 (N_1671,In_551,In_661);
xor U1672 (N_1672,In_908,In_364);
xor U1673 (N_1673,In_60,In_784);
or U1674 (N_1674,In_386,In_314);
and U1675 (N_1675,In_490,In_957);
nand U1676 (N_1676,In_318,In_617);
nor U1677 (N_1677,In_539,In_603);
and U1678 (N_1678,In_408,In_986);
xor U1679 (N_1679,In_730,In_809);
nor U1680 (N_1680,In_592,In_993);
and U1681 (N_1681,In_762,In_536);
nand U1682 (N_1682,In_198,In_120);
and U1683 (N_1683,In_681,In_991);
nor U1684 (N_1684,In_29,In_757);
xor U1685 (N_1685,In_819,In_507);
and U1686 (N_1686,In_49,In_486);
and U1687 (N_1687,In_260,In_540);
nor U1688 (N_1688,In_677,In_54);
and U1689 (N_1689,In_759,In_92);
or U1690 (N_1690,In_188,In_721);
and U1691 (N_1691,In_656,In_665);
nor U1692 (N_1692,In_339,In_960);
xnor U1693 (N_1693,In_920,In_70);
nor U1694 (N_1694,In_291,In_387);
and U1695 (N_1695,In_417,In_395);
xor U1696 (N_1696,In_373,In_746);
nor U1697 (N_1697,In_863,In_279);
and U1698 (N_1698,In_693,In_45);
nand U1699 (N_1699,In_229,In_576);
and U1700 (N_1700,In_370,In_488);
nand U1701 (N_1701,In_165,In_656);
and U1702 (N_1702,In_991,In_810);
xor U1703 (N_1703,In_250,In_296);
nand U1704 (N_1704,In_177,In_956);
xor U1705 (N_1705,In_150,In_18);
or U1706 (N_1706,In_159,In_698);
and U1707 (N_1707,In_573,In_342);
or U1708 (N_1708,In_527,In_136);
or U1709 (N_1709,In_100,In_42);
and U1710 (N_1710,In_88,In_762);
nand U1711 (N_1711,In_868,In_680);
nand U1712 (N_1712,In_697,In_347);
or U1713 (N_1713,In_377,In_988);
nor U1714 (N_1714,In_929,In_980);
xnor U1715 (N_1715,In_550,In_689);
or U1716 (N_1716,In_932,In_646);
nand U1717 (N_1717,In_280,In_769);
and U1718 (N_1718,In_567,In_474);
nor U1719 (N_1719,In_110,In_250);
nand U1720 (N_1720,In_43,In_179);
and U1721 (N_1721,In_850,In_826);
nor U1722 (N_1722,In_37,In_583);
and U1723 (N_1723,In_120,In_770);
and U1724 (N_1724,In_42,In_210);
nand U1725 (N_1725,In_775,In_480);
xor U1726 (N_1726,In_37,In_605);
nor U1727 (N_1727,In_301,In_530);
or U1728 (N_1728,In_783,In_623);
nor U1729 (N_1729,In_599,In_960);
or U1730 (N_1730,In_432,In_447);
nor U1731 (N_1731,In_678,In_645);
nor U1732 (N_1732,In_650,In_746);
xor U1733 (N_1733,In_649,In_477);
xnor U1734 (N_1734,In_221,In_722);
and U1735 (N_1735,In_583,In_862);
nand U1736 (N_1736,In_614,In_3);
nand U1737 (N_1737,In_599,In_488);
nor U1738 (N_1738,In_175,In_790);
nor U1739 (N_1739,In_205,In_269);
nor U1740 (N_1740,In_874,In_344);
xnor U1741 (N_1741,In_374,In_858);
or U1742 (N_1742,In_747,In_952);
nand U1743 (N_1743,In_222,In_307);
nand U1744 (N_1744,In_141,In_443);
or U1745 (N_1745,In_437,In_619);
or U1746 (N_1746,In_321,In_123);
and U1747 (N_1747,In_589,In_686);
xor U1748 (N_1748,In_819,In_100);
nand U1749 (N_1749,In_619,In_372);
nor U1750 (N_1750,In_77,In_758);
nand U1751 (N_1751,In_35,In_327);
nand U1752 (N_1752,In_388,In_62);
nor U1753 (N_1753,In_648,In_50);
nand U1754 (N_1754,In_31,In_816);
nor U1755 (N_1755,In_650,In_231);
nor U1756 (N_1756,In_446,In_488);
nor U1757 (N_1757,In_308,In_107);
nand U1758 (N_1758,In_34,In_622);
and U1759 (N_1759,In_402,In_997);
and U1760 (N_1760,In_439,In_830);
or U1761 (N_1761,In_915,In_928);
or U1762 (N_1762,In_404,In_286);
nor U1763 (N_1763,In_110,In_688);
xor U1764 (N_1764,In_617,In_533);
xnor U1765 (N_1765,In_795,In_718);
nand U1766 (N_1766,In_265,In_14);
nor U1767 (N_1767,In_469,In_614);
nor U1768 (N_1768,In_540,In_234);
or U1769 (N_1769,In_281,In_235);
or U1770 (N_1770,In_735,In_385);
nand U1771 (N_1771,In_269,In_38);
and U1772 (N_1772,In_974,In_423);
xnor U1773 (N_1773,In_778,In_374);
or U1774 (N_1774,In_892,In_736);
xnor U1775 (N_1775,In_800,In_43);
and U1776 (N_1776,In_940,In_846);
nand U1777 (N_1777,In_469,In_51);
or U1778 (N_1778,In_562,In_19);
nor U1779 (N_1779,In_122,In_450);
and U1780 (N_1780,In_704,In_920);
xor U1781 (N_1781,In_46,In_699);
nor U1782 (N_1782,In_70,In_340);
or U1783 (N_1783,In_33,In_90);
xnor U1784 (N_1784,In_950,In_121);
nor U1785 (N_1785,In_951,In_994);
nor U1786 (N_1786,In_424,In_402);
xor U1787 (N_1787,In_686,In_674);
nor U1788 (N_1788,In_841,In_486);
nor U1789 (N_1789,In_473,In_389);
xor U1790 (N_1790,In_890,In_816);
and U1791 (N_1791,In_411,In_94);
nor U1792 (N_1792,In_364,In_516);
and U1793 (N_1793,In_153,In_671);
or U1794 (N_1794,In_665,In_412);
nand U1795 (N_1795,In_229,In_892);
and U1796 (N_1796,In_847,In_711);
xor U1797 (N_1797,In_836,In_884);
and U1798 (N_1798,In_397,In_79);
or U1799 (N_1799,In_173,In_411);
or U1800 (N_1800,In_588,In_462);
nor U1801 (N_1801,In_496,In_311);
or U1802 (N_1802,In_812,In_440);
xor U1803 (N_1803,In_709,In_383);
nand U1804 (N_1804,In_907,In_481);
or U1805 (N_1805,In_599,In_292);
or U1806 (N_1806,In_636,In_874);
xor U1807 (N_1807,In_776,In_164);
and U1808 (N_1808,In_532,In_216);
or U1809 (N_1809,In_73,In_130);
nor U1810 (N_1810,In_221,In_150);
xor U1811 (N_1811,In_423,In_124);
and U1812 (N_1812,In_600,In_708);
or U1813 (N_1813,In_233,In_724);
nor U1814 (N_1814,In_730,In_226);
and U1815 (N_1815,In_760,In_549);
xnor U1816 (N_1816,In_994,In_403);
xor U1817 (N_1817,In_607,In_331);
xor U1818 (N_1818,In_421,In_687);
and U1819 (N_1819,In_25,In_857);
nor U1820 (N_1820,In_86,In_940);
or U1821 (N_1821,In_317,In_792);
xnor U1822 (N_1822,In_327,In_582);
nor U1823 (N_1823,In_953,In_545);
and U1824 (N_1824,In_710,In_158);
xnor U1825 (N_1825,In_510,In_115);
nor U1826 (N_1826,In_346,In_152);
or U1827 (N_1827,In_288,In_491);
and U1828 (N_1828,In_500,In_879);
or U1829 (N_1829,In_802,In_176);
and U1830 (N_1830,In_816,In_333);
or U1831 (N_1831,In_951,In_133);
nand U1832 (N_1832,In_192,In_127);
xnor U1833 (N_1833,In_886,In_512);
and U1834 (N_1834,In_358,In_994);
xor U1835 (N_1835,In_403,In_516);
xnor U1836 (N_1836,In_161,In_523);
xnor U1837 (N_1837,In_467,In_365);
nand U1838 (N_1838,In_125,In_43);
or U1839 (N_1839,In_635,In_382);
or U1840 (N_1840,In_367,In_916);
xor U1841 (N_1841,In_511,In_421);
xor U1842 (N_1842,In_886,In_42);
or U1843 (N_1843,In_577,In_680);
nor U1844 (N_1844,In_308,In_443);
and U1845 (N_1845,In_384,In_377);
or U1846 (N_1846,In_434,In_991);
and U1847 (N_1847,In_130,In_700);
or U1848 (N_1848,In_428,In_482);
nor U1849 (N_1849,In_211,In_647);
xor U1850 (N_1850,In_997,In_835);
xor U1851 (N_1851,In_893,In_801);
nand U1852 (N_1852,In_743,In_640);
xnor U1853 (N_1853,In_588,In_697);
or U1854 (N_1854,In_146,In_835);
nand U1855 (N_1855,In_135,In_760);
nand U1856 (N_1856,In_725,In_163);
and U1857 (N_1857,In_766,In_177);
or U1858 (N_1858,In_931,In_135);
and U1859 (N_1859,In_452,In_263);
or U1860 (N_1860,In_974,In_455);
xor U1861 (N_1861,In_320,In_569);
nand U1862 (N_1862,In_597,In_969);
xnor U1863 (N_1863,In_289,In_938);
and U1864 (N_1864,In_978,In_809);
xor U1865 (N_1865,In_954,In_496);
xor U1866 (N_1866,In_789,In_602);
nand U1867 (N_1867,In_152,In_388);
nor U1868 (N_1868,In_980,In_682);
and U1869 (N_1869,In_307,In_321);
and U1870 (N_1870,In_999,In_302);
nor U1871 (N_1871,In_413,In_880);
and U1872 (N_1872,In_219,In_907);
and U1873 (N_1873,In_93,In_298);
xor U1874 (N_1874,In_525,In_646);
xnor U1875 (N_1875,In_466,In_677);
or U1876 (N_1876,In_209,In_960);
xor U1877 (N_1877,In_648,In_118);
nor U1878 (N_1878,In_311,In_495);
nor U1879 (N_1879,In_410,In_110);
xnor U1880 (N_1880,In_147,In_792);
xnor U1881 (N_1881,In_826,In_691);
and U1882 (N_1882,In_531,In_165);
nand U1883 (N_1883,In_606,In_131);
xnor U1884 (N_1884,In_941,In_320);
and U1885 (N_1885,In_904,In_903);
xor U1886 (N_1886,In_928,In_388);
or U1887 (N_1887,In_820,In_881);
nor U1888 (N_1888,In_147,In_997);
or U1889 (N_1889,In_211,In_756);
xor U1890 (N_1890,In_961,In_527);
or U1891 (N_1891,In_346,In_297);
nand U1892 (N_1892,In_364,In_586);
nor U1893 (N_1893,In_626,In_193);
nand U1894 (N_1894,In_451,In_678);
and U1895 (N_1895,In_396,In_394);
and U1896 (N_1896,In_245,In_622);
and U1897 (N_1897,In_442,In_471);
xnor U1898 (N_1898,In_109,In_9);
or U1899 (N_1899,In_655,In_979);
xnor U1900 (N_1900,In_976,In_391);
nor U1901 (N_1901,In_248,In_372);
or U1902 (N_1902,In_850,In_816);
and U1903 (N_1903,In_939,In_377);
nor U1904 (N_1904,In_601,In_233);
xnor U1905 (N_1905,In_958,In_319);
or U1906 (N_1906,In_910,In_852);
nand U1907 (N_1907,In_121,In_898);
nand U1908 (N_1908,In_844,In_53);
and U1909 (N_1909,In_183,In_909);
xnor U1910 (N_1910,In_863,In_719);
or U1911 (N_1911,In_176,In_118);
nor U1912 (N_1912,In_676,In_769);
xnor U1913 (N_1913,In_402,In_775);
nand U1914 (N_1914,In_491,In_970);
nor U1915 (N_1915,In_594,In_98);
or U1916 (N_1916,In_919,In_391);
xor U1917 (N_1917,In_189,In_888);
or U1918 (N_1918,In_469,In_718);
xor U1919 (N_1919,In_409,In_308);
nand U1920 (N_1920,In_289,In_159);
or U1921 (N_1921,In_11,In_907);
nor U1922 (N_1922,In_523,In_675);
xor U1923 (N_1923,In_306,In_442);
and U1924 (N_1924,In_529,In_205);
and U1925 (N_1925,In_168,In_559);
or U1926 (N_1926,In_524,In_35);
nand U1927 (N_1927,In_469,In_642);
or U1928 (N_1928,In_237,In_622);
and U1929 (N_1929,In_673,In_192);
nor U1930 (N_1930,In_408,In_693);
or U1931 (N_1931,In_50,In_78);
xnor U1932 (N_1932,In_389,In_713);
nor U1933 (N_1933,In_725,In_191);
nand U1934 (N_1934,In_228,In_791);
or U1935 (N_1935,In_317,In_149);
or U1936 (N_1936,In_721,In_468);
or U1937 (N_1937,In_966,In_714);
nand U1938 (N_1938,In_193,In_211);
xnor U1939 (N_1939,In_102,In_744);
xnor U1940 (N_1940,In_738,In_909);
xnor U1941 (N_1941,In_148,In_265);
xor U1942 (N_1942,In_679,In_839);
nor U1943 (N_1943,In_737,In_921);
or U1944 (N_1944,In_407,In_437);
nand U1945 (N_1945,In_820,In_852);
xor U1946 (N_1946,In_607,In_395);
nand U1947 (N_1947,In_299,In_548);
and U1948 (N_1948,In_220,In_688);
xnor U1949 (N_1949,In_80,In_184);
xnor U1950 (N_1950,In_72,In_269);
or U1951 (N_1951,In_371,In_230);
nand U1952 (N_1952,In_740,In_276);
and U1953 (N_1953,In_697,In_473);
nand U1954 (N_1954,In_33,In_911);
xnor U1955 (N_1955,In_808,In_942);
or U1956 (N_1956,In_528,In_988);
nand U1957 (N_1957,In_61,In_191);
and U1958 (N_1958,In_435,In_446);
or U1959 (N_1959,In_443,In_507);
xor U1960 (N_1960,In_776,In_882);
or U1961 (N_1961,In_114,In_245);
or U1962 (N_1962,In_201,In_562);
nand U1963 (N_1963,In_825,In_386);
nor U1964 (N_1964,In_579,In_635);
and U1965 (N_1965,In_144,In_827);
or U1966 (N_1966,In_282,In_558);
nand U1967 (N_1967,In_891,In_42);
nand U1968 (N_1968,In_886,In_32);
or U1969 (N_1969,In_980,In_634);
xnor U1970 (N_1970,In_42,In_923);
xor U1971 (N_1971,In_144,In_497);
and U1972 (N_1972,In_700,In_119);
or U1973 (N_1973,In_247,In_567);
xor U1974 (N_1974,In_723,In_41);
and U1975 (N_1975,In_694,In_194);
or U1976 (N_1976,In_103,In_589);
nor U1977 (N_1977,In_510,In_818);
nand U1978 (N_1978,In_533,In_561);
and U1979 (N_1979,In_289,In_492);
nor U1980 (N_1980,In_392,In_562);
or U1981 (N_1981,In_844,In_828);
xnor U1982 (N_1982,In_910,In_142);
xnor U1983 (N_1983,In_162,In_806);
nand U1984 (N_1984,In_870,In_649);
nor U1985 (N_1985,In_878,In_661);
xnor U1986 (N_1986,In_796,In_879);
nand U1987 (N_1987,In_793,In_540);
xnor U1988 (N_1988,In_590,In_747);
or U1989 (N_1989,In_186,In_664);
xnor U1990 (N_1990,In_788,In_135);
or U1991 (N_1991,In_564,In_527);
and U1992 (N_1992,In_975,In_133);
nor U1993 (N_1993,In_967,In_567);
nand U1994 (N_1994,In_460,In_5);
nor U1995 (N_1995,In_275,In_522);
nor U1996 (N_1996,In_549,In_222);
and U1997 (N_1997,In_803,In_786);
and U1998 (N_1998,In_275,In_110);
nand U1999 (N_1999,In_166,In_176);
xnor U2000 (N_2000,In_219,In_784);
xnor U2001 (N_2001,In_361,In_720);
and U2002 (N_2002,In_416,In_260);
xor U2003 (N_2003,In_852,In_931);
and U2004 (N_2004,In_951,In_484);
and U2005 (N_2005,In_165,In_941);
nor U2006 (N_2006,In_381,In_980);
xnor U2007 (N_2007,In_997,In_966);
or U2008 (N_2008,In_34,In_370);
xnor U2009 (N_2009,In_224,In_635);
or U2010 (N_2010,In_71,In_398);
nor U2011 (N_2011,In_754,In_816);
or U2012 (N_2012,In_697,In_142);
or U2013 (N_2013,In_352,In_114);
nand U2014 (N_2014,In_562,In_759);
xnor U2015 (N_2015,In_31,In_984);
nor U2016 (N_2016,In_150,In_8);
nor U2017 (N_2017,In_136,In_675);
nor U2018 (N_2018,In_307,In_212);
and U2019 (N_2019,In_27,In_352);
xnor U2020 (N_2020,In_151,In_828);
or U2021 (N_2021,In_529,In_77);
nor U2022 (N_2022,In_681,In_526);
xor U2023 (N_2023,In_372,In_352);
nor U2024 (N_2024,In_700,In_754);
nor U2025 (N_2025,In_528,In_886);
nand U2026 (N_2026,In_163,In_152);
nand U2027 (N_2027,In_556,In_271);
or U2028 (N_2028,In_580,In_319);
or U2029 (N_2029,In_330,In_961);
nor U2030 (N_2030,In_611,In_832);
and U2031 (N_2031,In_842,In_24);
nor U2032 (N_2032,In_847,In_992);
nand U2033 (N_2033,In_159,In_893);
and U2034 (N_2034,In_155,In_57);
nor U2035 (N_2035,In_848,In_188);
xnor U2036 (N_2036,In_696,In_965);
xor U2037 (N_2037,In_98,In_465);
xnor U2038 (N_2038,In_885,In_156);
nor U2039 (N_2039,In_57,In_259);
xor U2040 (N_2040,In_413,In_674);
xnor U2041 (N_2041,In_368,In_80);
nor U2042 (N_2042,In_314,In_764);
nor U2043 (N_2043,In_233,In_951);
xor U2044 (N_2044,In_212,In_931);
and U2045 (N_2045,In_898,In_884);
or U2046 (N_2046,In_540,In_879);
nand U2047 (N_2047,In_503,In_831);
and U2048 (N_2048,In_677,In_142);
nand U2049 (N_2049,In_751,In_721);
nor U2050 (N_2050,In_972,In_186);
nor U2051 (N_2051,In_379,In_840);
nand U2052 (N_2052,In_827,In_893);
xor U2053 (N_2053,In_602,In_305);
nand U2054 (N_2054,In_674,In_439);
or U2055 (N_2055,In_22,In_371);
and U2056 (N_2056,In_271,In_292);
xnor U2057 (N_2057,In_822,In_236);
nor U2058 (N_2058,In_140,In_314);
nand U2059 (N_2059,In_131,In_864);
and U2060 (N_2060,In_978,In_880);
nor U2061 (N_2061,In_887,In_359);
nand U2062 (N_2062,In_62,In_749);
nand U2063 (N_2063,In_770,In_37);
or U2064 (N_2064,In_248,In_24);
nand U2065 (N_2065,In_88,In_563);
or U2066 (N_2066,In_437,In_97);
nand U2067 (N_2067,In_614,In_104);
nor U2068 (N_2068,In_422,In_394);
nand U2069 (N_2069,In_299,In_765);
and U2070 (N_2070,In_528,In_120);
and U2071 (N_2071,In_181,In_915);
and U2072 (N_2072,In_142,In_779);
or U2073 (N_2073,In_863,In_846);
nand U2074 (N_2074,In_932,In_447);
and U2075 (N_2075,In_304,In_879);
nand U2076 (N_2076,In_42,In_697);
and U2077 (N_2077,In_198,In_326);
nand U2078 (N_2078,In_199,In_418);
nand U2079 (N_2079,In_832,In_545);
nand U2080 (N_2080,In_749,In_67);
or U2081 (N_2081,In_47,In_264);
nand U2082 (N_2082,In_740,In_670);
nand U2083 (N_2083,In_223,In_847);
nor U2084 (N_2084,In_802,In_316);
xnor U2085 (N_2085,In_358,In_549);
and U2086 (N_2086,In_48,In_915);
or U2087 (N_2087,In_157,In_934);
nor U2088 (N_2088,In_56,In_54);
nor U2089 (N_2089,In_38,In_493);
nand U2090 (N_2090,In_709,In_832);
nand U2091 (N_2091,In_803,In_179);
nor U2092 (N_2092,In_562,In_49);
and U2093 (N_2093,In_531,In_432);
nor U2094 (N_2094,In_165,In_839);
nand U2095 (N_2095,In_245,In_682);
nand U2096 (N_2096,In_856,In_784);
nor U2097 (N_2097,In_885,In_43);
or U2098 (N_2098,In_60,In_806);
xnor U2099 (N_2099,In_60,In_310);
or U2100 (N_2100,In_182,In_866);
nand U2101 (N_2101,In_661,In_801);
and U2102 (N_2102,In_234,In_845);
xor U2103 (N_2103,In_431,In_760);
nand U2104 (N_2104,In_934,In_359);
nand U2105 (N_2105,In_552,In_183);
and U2106 (N_2106,In_377,In_879);
nor U2107 (N_2107,In_22,In_651);
nor U2108 (N_2108,In_165,In_99);
and U2109 (N_2109,In_7,In_775);
and U2110 (N_2110,In_684,In_208);
or U2111 (N_2111,In_898,In_37);
or U2112 (N_2112,In_214,In_54);
nor U2113 (N_2113,In_573,In_340);
nor U2114 (N_2114,In_996,In_926);
nor U2115 (N_2115,In_317,In_888);
nand U2116 (N_2116,In_435,In_750);
xor U2117 (N_2117,In_988,In_234);
xnor U2118 (N_2118,In_297,In_328);
nor U2119 (N_2119,In_706,In_177);
nor U2120 (N_2120,In_832,In_115);
nor U2121 (N_2121,In_187,In_195);
nor U2122 (N_2122,In_914,In_946);
nand U2123 (N_2123,In_0,In_372);
xnor U2124 (N_2124,In_711,In_514);
xnor U2125 (N_2125,In_873,In_940);
and U2126 (N_2126,In_886,In_643);
and U2127 (N_2127,In_357,In_444);
xor U2128 (N_2128,In_365,In_479);
and U2129 (N_2129,In_466,In_442);
xor U2130 (N_2130,In_432,In_903);
nand U2131 (N_2131,In_98,In_878);
nor U2132 (N_2132,In_67,In_904);
nand U2133 (N_2133,In_100,In_903);
nor U2134 (N_2134,In_470,In_704);
or U2135 (N_2135,In_619,In_521);
nand U2136 (N_2136,In_120,In_357);
nor U2137 (N_2137,In_293,In_726);
or U2138 (N_2138,In_877,In_859);
and U2139 (N_2139,In_86,In_539);
or U2140 (N_2140,In_661,In_530);
and U2141 (N_2141,In_386,In_182);
nor U2142 (N_2142,In_110,In_287);
and U2143 (N_2143,In_858,In_874);
nand U2144 (N_2144,In_771,In_128);
xnor U2145 (N_2145,In_871,In_516);
nand U2146 (N_2146,In_957,In_754);
and U2147 (N_2147,In_6,In_565);
and U2148 (N_2148,In_303,In_533);
nor U2149 (N_2149,In_881,In_972);
nor U2150 (N_2150,In_316,In_120);
nand U2151 (N_2151,In_112,In_664);
nor U2152 (N_2152,In_902,In_49);
or U2153 (N_2153,In_277,In_679);
and U2154 (N_2154,In_352,In_884);
nor U2155 (N_2155,In_721,In_637);
or U2156 (N_2156,In_165,In_834);
nor U2157 (N_2157,In_158,In_127);
and U2158 (N_2158,In_284,In_542);
xnor U2159 (N_2159,In_450,In_712);
nor U2160 (N_2160,In_369,In_775);
nor U2161 (N_2161,In_15,In_67);
and U2162 (N_2162,In_760,In_5);
xor U2163 (N_2163,In_21,In_286);
xor U2164 (N_2164,In_185,In_812);
xnor U2165 (N_2165,In_772,In_238);
xor U2166 (N_2166,In_182,In_293);
nor U2167 (N_2167,In_124,In_734);
nand U2168 (N_2168,In_925,In_438);
xor U2169 (N_2169,In_959,In_137);
nor U2170 (N_2170,In_758,In_90);
and U2171 (N_2171,In_332,In_947);
nor U2172 (N_2172,In_903,In_86);
nor U2173 (N_2173,In_771,In_553);
nor U2174 (N_2174,In_749,In_315);
or U2175 (N_2175,In_216,In_512);
xor U2176 (N_2176,In_543,In_789);
xnor U2177 (N_2177,In_408,In_5);
xnor U2178 (N_2178,In_454,In_836);
nand U2179 (N_2179,In_956,In_738);
nor U2180 (N_2180,In_361,In_895);
nand U2181 (N_2181,In_849,In_488);
xnor U2182 (N_2182,In_28,In_994);
nand U2183 (N_2183,In_97,In_57);
and U2184 (N_2184,In_232,In_179);
or U2185 (N_2185,In_202,In_808);
and U2186 (N_2186,In_765,In_121);
xnor U2187 (N_2187,In_78,In_158);
or U2188 (N_2188,In_911,In_119);
nand U2189 (N_2189,In_926,In_67);
nor U2190 (N_2190,In_285,In_769);
xnor U2191 (N_2191,In_730,In_667);
nor U2192 (N_2192,In_604,In_406);
nand U2193 (N_2193,In_937,In_269);
nor U2194 (N_2194,In_779,In_4);
xnor U2195 (N_2195,In_390,In_583);
or U2196 (N_2196,In_732,In_875);
or U2197 (N_2197,In_502,In_962);
and U2198 (N_2198,In_602,In_312);
nor U2199 (N_2199,In_674,In_682);
nor U2200 (N_2200,In_823,In_83);
or U2201 (N_2201,In_970,In_234);
and U2202 (N_2202,In_864,In_211);
xnor U2203 (N_2203,In_196,In_726);
nand U2204 (N_2204,In_30,In_642);
xnor U2205 (N_2205,In_368,In_812);
or U2206 (N_2206,In_226,In_652);
nor U2207 (N_2207,In_88,In_461);
or U2208 (N_2208,In_474,In_801);
or U2209 (N_2209,In_363,In_370);
nand U2210 (N_2210,In_998,In_59);
nor U2211 (N_2211,In_278,In_747);
and U2212 (N_2212,In_742,In_668);
or U2213 (N_2213,In_445,In_695);
nand U2214 (N_2214,In_906,In_308);
nand U2215 (N_2215,In_819,In_34);
xor U2216 (N_2216,In_330,In_864);
xnor U2217 (N_2217,In_247,In_150);
and U2218 (N_2218,In_829,In_841);
xor U2219 (N_2219,In_243,In_795);
and U2220 (N_2220,In_492,In_165);
or U2221 (N_2221,In_884,In_675);
nand U2222 (N_2222,In_477,In_524);
nor U2223 (N_2223,In_251,In_873);
xnor U2224 (N_2224,In_72,In_601);
nor U2225 (N_2225,In_280,In_736);
and U2226 (N_2226,In_502,In_828);
and U2227 (N_2227,In_327,In_494);
nor U2228 (N_2228,In_80,In_151);
or U2229 (N_2229,In_0,In_646);
and U2230 (N_2230,In_922,In_492);
or U2231 (N_2231,In_260,In_216);
or U2232 (N_2232,In_248,In_904);
nor U2233 (N_2233,In_580,In_564);
nor U2234 (N_2234,In_791,In_986);
xnor U2235 (N_2235,In_478,In_114);
xnor U2236 (N_2236,In_9,In_192);
and U2237 (N_2237,In_15,In_930);
nor U2238 (N_2238,In_828,In_201);
and U2239 (N_2239,In_296,In_457);
and U2240 (N_2240,In_437,In_865);
nor U2241 (N_2241,In_233,In_935);
nor U2242 (N_2242,In_590,In_532);
nor U2243 (N_2243,In_685,In_943);
or U2244 (N_2244,In_810,In_364);
nor U2245 (N_2245,In_582,In_536);
or U2246 (N_2246,In_723,In_210);
xnor U2247 (N_2247,In_990,In_829);
or U2248 (N_2248,In_686,In_410);
nand U2249 (N_2249,In_150,In_428);
and U2250 (N_2250,In_953,In_260);
nand U2251 (N_2251,In_39,In_951);
and U2252 (N_2252,In_863,In_133);
nand U2253 (N_2253,In_9,In_310);
and U2254 (N_2254,In_566,In_272);
xor U2255 (N_2255,In_135,In_850);
and U2256 (N_2256,In_860,In_877);
and U2257 (N_2257,In_178,In_868);
nor U2258 (N_2258,In_446,In_240);
nor U2259 (N_2259,In_856,In_925);
and U2260 (N_2260,In_816,In_603);
nor U2261 (N_2261,In_474,In_253);
nand U2262 (N_2262,In_108,In_121);
nor U2263 (N_2263,In_923,In_746);
and U2264 (N_2264,In_149,In_93);
and U2265 (N_2265,In_750,In_616);
xnor U2266 (N_2266,In_959,In_71);
or U2267 (N_2267,In_202,In_764);
xor U2268 (N_2268,In_729,In_105);
nor U2269 (N_2269,In_762,In_908);
or U2270 (N_2270,In_70,In_626);
and U2271 (N_2271,In_695,In_601);
nor U2272 (N_2272,In_285,In_246);
and U2273 (N_2273,In_7,In_744);
nor U2274 (N_2274,In_991,In_103);
nand U2275 (N_2275,In_958,In_849);
and U2276 (N_2276,In_115,In_546);
or U2277 (N_2277,In_656,In_454);
or U2278 (N_2278,In_75,In_931);
nand U2279 (N_2279,In_309,In_852);
nand U2280 (N_2280,In_373,In_785);
or U2281 (N_2281,In_139,In_155);
and U2282 (N_2282,In_344,In_526);
and U2283 (N_2283,In_222,In_639);
and U2284 (N_2284,In_423,In_230);
nor U2285 (N_2285,In_109,In_179);
xor U2286 (N_2286,In_260,In_34);
nand U2287 (N_2287,In_5,In_119);
nand U2288 (N_2288,In_788,In_326);
nor U2289 (N_2289,In_845,In_730);
or U2290 (N_2290,In_152,In_432);
xnor U2291 (N_2291,In_643,In_895);
nor U2292 (N_2292,In_228,In_480);
xor U2293 (N_2293,In_843,In_616);
nor U2294 (N_2294,In_136,In_559);
or U2295 (N_2295,In_482,In_846);
xor U2296 (N_2296,In_732,In_322);
xor U2297 (N_2297,In_715,In_112);
or U2298 (N_2298,In_830,In_533);
nor U2299 (N_2299,In_987,In_885);
or U2300 (N_2300,In_475,In_765);
nor U2301 (N_2301,In_308,In_819);
xor U2302 (N_2302,In_306,In_267);
xnor U2303 (N_2303,In_974,In_566);
nor U2304 (N_2304,In_742,In_801);
and U2305 (N_2305,In_478,In_741);
or U2306 (N_2306,In_69,In_982);
nor U2307 (N_2307,In_197,In_217);
xnor U2308 (N_2308,In_650,In_327);
xor U2309 (N_2309,In_894,In_354);
xor U2310 (N_2310,In_338,In_779);
nor U2311 (N_2311,In_189,In_695);
or U2312 (N_2312,In_673,In_450);
nor U2313 (N_2313,In_113,In_79);
and U2314 (N_2314,In_899,In_274);
nand U2315 (N_2315,In_324,In_944);
or U2316 (N_2316,In_282,In_903);
and U2317 (N_2317,In_975,In_369);
xor U2318 (N_2318,In_7,In_319);
nand U2319 (N_2319,In_970,In_14);
and U2320 (N_2320,In_960,In_816);
xor U2321 (N_2321,In_858,In_538);
and U2322 (N_2322,In_435,In_875);
nor U2323 (N_2323,In_234,In_542);
or U2324 (N_2324,In_303,In_548);
or U2325 (N_2325,In_469,In_400);
or U2326 (N_2326,In_995,In_438);
nand U2327 (N_2327,In_385,In_79);
xor U2328 (N_2328,In_992,In_397);
and U2329 (N_2329,In_885,In_615);
xnor U2330 (N_2330,In_586,In_108);
or U2331 (N_2331,In_805,In_884);
and U2332 (N_2332,In_466,In_88);
xor U2333 (N_2333,In_822,In_226);
xnor U2334 (N_2334,In_164,In_857);
or U2335 (N_2335,In_62,In_403);
xnor U2336 (N_2336,In_679,In_283);
xor U2337 (N_2337,In_487,In_825);
and U2338 (N_2338,In_539,In_451);
and U2339 (N_2339,In_42,In_990);
nand U2340 (N_2340,In_675,In_937);
nor U2341 (N_2341,In_560,In_480);
and U2342 (N_2342,In_24,In_448);
nor U2343 (N_2343,In_581,In_518);
nand U2344 (N_2344,In_789,In_778);
and U2345 (N_2345,In_270,In_636);
xnor U2346 (N_2346,In_196,In_707);
nor U2347 (N_2347,In_265,In_767);
nor U2348 (N_2348,In_429,In_552);
and U2349 (N_2349,In_916,In_6);
xor U2350 (N_2350,In_345,In_220);
nand U2351 (N_2351,In_99,In_196);
and U2352 (N_2352,In_654,In_623);
xnor U2353 (N_2353,In_652,In_121);
or U2354 (N_2354,In_511,In_76);
nor U2355 (N_2355,In_983,In_134);
nor U2356 (N_2356,In_505,In_121);
nand U2357 (N_2357,In_442,In_972);
or U2358 (N_2358,In_253,In_906);
and U2359 (N_2359,In_832,In_12);
nand U2360 (N_2360,In_373,In_258);
or U2361 (N_2361,In_698,In_447);
and U2362 (N_2362,In_741,In_552);
xnor U2363 (N_2363,In_88,In_982);
or U2364 (N_2364,In_277,In_116);
nor U2365 (N_2365,In_967,In_880);
nand U2366 (N_2366,In_99,In_56);
nand U2367 (N_2367,In_274,In_430);
nor U2368 (N_2368,In_315,In_408);
nor U2369 (N_2369,In_576,In_393);
nor U2370 (N_2370,In_222,In_301);
or U2371 (N_2371,In_859,In_819);
or U2372 (N_2372,In_440,In_509);
or U2373 (N_2373,In_771,In_725);
or U2374 (N_2374,In_306,In_522);
or U2375 (N_2375,In_944,In_185);
or U2376 (N_2376,In_843,In_356);
and U2377 (N_2377,In_128,In_719);
nor U2378 (N_2378,In_696,In_137);
nand U2379 (N_2379,In_397,In_474);
and U2380 (N_2380,In_370,In_524);
xor U2381 (N_2381,In_968,In_278);
xnor U2382 (N_2382,In_701,In_282);
and U2383 (N_2383,In_391,In_230);
and U2384 (N_2384,In_551,In_74);
or U2385 (N_2385,In_286,In_175);
nand U2386 (N_2386,In_568,In_834);
or U2387 (N_2387,In_69,In_137);
nor U2388 (N_2388,In_377,In_998);
nor U2389 (N_2389,In_609,In_215);
xor U2390 (N_2390,In_258,In_191);
xor U2391 (N_2391,In_305,In_372);
xor U2392 (N_2392,In_340,In_927);
xnor U2393 (N_2393,In_505,In_232);
xnor U2394 (N_2394,In_869,In_261);
nand U2395 (N_2395,In_85,In_915);
or U2396 (N_2396,In_914,In_667);
nand U2397 (N_2397,In_205,In_991);
nor U2398 (N_2398,In_976,In_916);
or U2399 (N_2399,In_880,In_996);
xor U2400 (N_2400,In_328,In_399);
xor U2401 (N_2401,In_160,In_156);
or U2402 (N_2402,In_567,In_770);
nor U2403 (N_2403,In_392,In_565);
nor U2404 (N_2404,In_136,In_112);
and U2405 (N_2405,In_311,In_818);
xor U2406 (N_2406,In_250,In_194);
xnor U2407 (N_2407,In_790,In_614);
nor U2408 (N_2408,In_84,In_251);
and U2409 (N_2409,In_437,In_221);
xnor U2410 (N_2410,In_569,In_310);
and U2411 (N_2411,In_374,In_796);
and U2412 (N_2412,In_350,In_565);
or U2413 (N_2413,In_166,In_552);
nand U2414 (N_2414,In_639,In_678);
nand U2415 (N_2415,In_215,In_37);
nor U2416 (N_2416,In_578,In_582);
or U2417 (N_2417,In_794,In_783);
nor U2418 (N_2418,In_196,In_813);
xor U2419 (N_2419,In_332,In_113);
nor U2420 (N_2420,In_531,In_7);
and U2421 (N_2421,In_511,In_793);
and U2422 (N_2422,In_723,In_702);
xor U2423 (N_2423,In_737,In_399);
or U2424 (N_2424,In_342,In_195);
xor U2425 (N_2425,In_356,In_468);
nand U2426 (N_2426,In_250,In_314);
nand U2427 (N_2427,In_402,In_310);
and U2428 (N_2428,In_143,In_546);
or U2429 (N_2429,In_525,In_891);
xnor U2430 (N_2430,In_333,In_499);
nand U2431 (N_2431,In_325,In_383);
nor U2432 (N_2432,In_611,In_946);
or U2433 (N_2433,In_51,In_630);
nor U2434 (N_2434,In_417,In_42);
or U2435 (N_2435,In_45,In_797);
and U2436 (N_2436,In_913,In_568);
nor U2437 (N_2437,In_589,In_956);
xnor U2438 (N_2438,In_102,In_696);
or U2439 (N_2439,In_544,In_600);
nand U2440 (N_2440,In_795,In_611);
nor U2441 (N_2441,In_579,In_423);
nand U2442 (N_2442,In_759,In_486);
or U2443 (N_2443,In_145,In_950);
or U2444 (N_2444,In_781,In_374);
xor U2445 (N_2445,In_390,In_396);
nand U2446 (N_2446,In_38,In_161);
nor U2447 (N_2447,In_758,In_651);
nor U2448 (N_2448,In_53,In_160);
nor U2449 (N_2449,In_240,In_980);
and U2450 (N_2450,In_80,In_753);
nand U2451 (N_2451,In_183,In_351);
nor U2452 (N_2452,In_860,In_73);
xnor U2453 (N_2453,In_990,In_394);
xor U2454 (N_2454,In_832,In_37);
nand U2455 (N_2455,In_255,In_945);
or U2456 (N_2456,In_173,In_623);
nor U2457 (N_2457,In_425,In_483);
xnor U2458 (N_2458,In_157,In_256);
nor U2459 (N_2459,In_603,In_949);
or U2460 (N_2460,In_962,In_921);
nand U2461 (N_2461,In_784,In_300);
or U2462 (N_2462,In_65,In_743);
nand U2463 (N_2463,In_151,In_948);
nand U2464 (N_2464,In_208,In_271);
nand U2465 (N_2465,In_734,In_683);
nand U2466 (N_2466,In_508,In_544);
or U2467 (N_2467,In_242,In_861);
or U2468 (N_2468,In_696,In_602);
xnor U2469 (N_2469,In_4,In_69);
nor U2470 (N_2470,In_854,In_468);
and U2471 (N_2471,In_709,In_111);
nor U2472 (N_2472,In_171,In_305);
xnor U2473 (N_2473,In_708,In_612);
and U2474 (N_2474,In_532,In_905);
nor U2475 (N_2475,In_408,In_924);
and U2476 (N_2476,In_480,In_441);
nor U2477 (N_2477,In_342,In_604);
or U2478 (N_2478,In_95,In_609);
or U2479 (N_2479,In_459,In_585);
and U2480 (N_2480,In_360,In_768);
xor U2481 (N_2481,In_289,In_926);
nand U2482 (N_2482,In_229,In_640);
nor U2483 (N_2483,In_576,In_404);
nor U2484 (N_2484,In_655,In_602);
and U2485 (N_2485,In_676,In_583);
nor U2486 (N_2486,In_147,In_559);
and U2487 (N_2487,In_152,In_752);
and U2488 (N_2488,In_762,In_573);
xnor U2489 (N_2489,In_78,In_399);
nand U2490 (N_2490,In_829,In_334);
nor U2491 (N_2491,In_488,In_366);
nand U2492 (N_2492,In_942,In_156);
nor U2493 (N_2493,In_935,In_191);
and U2494 (N_2494,In_990,In_57);
nand U2495 (N_2495,In_498,In_694);
or U2496 (N_2496,In_695,In_369);
xor U2497 (N_2497,In_623,In_98);
and U2498 (N_2498,In_252,In_374);
and U2499 (N_2499,In_719,In_771);
nand U2500 (N_2500,N_60,N_1988);
and U2501 (N_2501,N_2492,N_896);
and U2502 (N_2502,N_1672,N_919);
nor U2503 (N_2503,N_2217,N_1558);
nor U2504 (N_2504,N_2037,N_161);
nor U2505 (N_2505,N_115,N_376);
nor U2506 (N_2506,N_686,N_236);
and U2507 (N_2507,N_2189,N_1641);
or U2508 (N_2508,N_2075,N_1744);
and U2509 (N_2509,N_229,N_1208);
xnor U2510 (N_2510,N_2303,N_1766);
nor U2511 (N_2511,N_136,N_1459);
and U2512 (N_2512,N_1767,N_2074);
or U2513 (N_2513,N_423,N_2481);
xnor U2514 (N_2514,N_324,N_1762);
or U2515 (N_2515,N_1981,N_1263);
xnor U2516 (N_2516,N_853,N_1800);
nand U2517 (N_2517,N_1940,N_166);
xnor U2518 (N_2518,N_884,N_542);
and U2519 (N_2519,N_204,N_1354);
and U2520 (N_2520,N_2200,N_7);
and U2521 (N_2521,N_304,N_1086);
nor U2522 (N_2522,N_2426,N_429);
or U2523 (N_2523,N_1039,N_1649);
xor U2524 (N_2524,N_794,N_1728);
xor U2525 (N_2525,N_1786,N_1544);
or U2526 (N_2526,N_1187,N_2375);
or U2527 (N_2527,N_840,N_186);
xnor U2528 (N_2528,N_1640,N_1332);
nor U2529 (N_2529,N_1624,N_994);
or U2530 (N_2530,N_2272,N_1137);
nand U2531 (N_2531,N_1328,N_347);
and U2532 (N_2532,N_874,N_1983);
xnor U2533 (N_2533,N_1235,N_798);
nor U2534 (N_2534,N_1169,N_2252);
nor U2535 (N_2535,N_1694,N_691);
and U2536 (N_2536,N_974,N_2030);
nor U2537 (N_2537,N_962,N_774);
or U2538 (N_2538,N_87,N_14);
and U2539 (N_2539,N_883,N_1524);
and U2540 (N_2540,N_1740,N_1618);
nand U2541 (N_2541,N_1548,N_992);
xor U2542 (N_2542,N_1690,N_768);
xor U2543 (N_2543,N_850,N_394);
nand U2544 (N_2544,N_632,N_1069);
nor U2545 (N_2545,N_1247,N_173);
or U2546 (N_2546,N_1484,N_854);
nand U2547 (N_2547,N_1696,N_1635);
nor U2548 (N_2548,N_598,N_1099);
and U2549 (N_2549,N_286,N_1140);
and U2550 (N_2550,N_135,N_2162);
nand U2551 (N_2551,N_799,N_1188);
xnor U2552 (N_2552,N_1523,N_495);
xnor U2553 (N_2553,N_1571,N_1449);
nor U2554 (N_2554,N_25,N_248);
xor U2555 (N_2555,N_206,N_2296);
nand U2556 (N_2556,N_1103,N_1772);
or U2557 (N_2557,N_1645,N_1859);
nor U2558 (N_2558,N_1415,N_2236);
nand U2559 (N_2559,N_1985,N_801);
xor U2560 (N_2560,N_2137,N_191);
nand U2561 (N_2561,N_594,N_1477);
or U2562 (N_2562,N_2202,N_510);
xor U2563 (N_2563,N_952,N_552);
nor U2564 (N_2564,N_2154,N_616);
and U2565 (N_2565,N_508,N_771);
nand U2566 (N_2566,N_537,N_543);
nor U2567 (N_2567,N_966,N_809);
or U2568 (N_2568,N_739,N_2175);
and U2569 (N_2569,N_1301,N_1688);
xor U2570 (N_2570,N_1977,N_231);
or U2571 (N_2571,N_1002,N_255);
and U2572 (N_2572,N_1280,N_1578);
nand U2573 (N_2573,N_1525,N_2003);
xor U2574 (N_2574,N_1220,N_1828);
and U2575 (N_2575,N_497,N_1982);
or U2576 (N_2576,N_1053,N_219);
and U2577 (N_2577,N_1612,N_1092);
nor U2578 (N_2578,N_348,N_708);
nor U2579 (N_2579,N_326,N_144);
and U2580 (N_2580,N_1036,N_649);
xnor U2581 (N_2581,N_1918,N_1898);
nand U2582 (N_2582,N_2483,N_1979);
and U2583 (N_2583,N_417,N_398);
and U2584 (N_2584,N_886,N_2312);
nor U2585 (N_2585,N_312,N_343);
nand U2586 (N_2586,N_1711,N_1619);
nand U2587 (N_2587,N_1458,N_1359);
and U2588 (N_2588,N_448,N_1933);
or U2589 (N_2589,N_1031,N_1734);
or U2590 (N_2590,N_609,N_2011);
xnor U2591 (N_2591,N_1972,N_357);
nor U2592 (N_2592,N_1242,N_728);
or U2593 (N_2593,N_1952,N_1543);
nor U2594 (N_2594,N_1147,N_1264);
xnor U2595 (N_2595,N_1156,N_785);
or U2596 (N_2596,N_1133,N_2216);
or U2597 (N_2597,N_2027,N_1349);
nor U2598 (N_2598,N_496,N_2320);
or U2599 (N_2599,N_477,N_869);
and U2600 (N_2600,N_789,N_2371);
and U2601 (N_2601,N_1335,N_778);
nor U2602 (N_2602,N_1120,N_1849);
or U2603 (N_2603,N_290,N_1228);
and U2604 (N_2604,N_205,N_877);
xor U2605 (N_2605,N_1342,N_2329);
or U2606 (N_2606,N_2226,N_182);
or U2607 (N_2607,N_2335,N_381);
and U2608 (N_2608,N_48,N_2254);
nor U2609 (N_2609,N_737,N_574);
or U2610 (N_2610,N_1588,N_2260);
nand U2611 (N_2611,N_1437,N_2013);
and U2612 (N_2612,N_984,N_1617);
and U2613 (N_2613,N_1807,N_1087);
nor U2614 (N_2614,N_989,N_1648);
nor U2615 (N_2615,N_1100,N_199);
or U2616 (N_2616,N_1655,N_1260);
and U2617 (N_2617,N_2125,N_656);
xor U2618 (N_2618,N_386,N_67);
nand U2619 (N_2619,N_1470,N_1546);
and U2620 (N_2620,N_1240,N_1621);
xor U2621 (N_2621,N_400,N_1320);
nand U2622 (N_2622,N_2392,N_291);
xnor U2623 (N_2623,N_791,N_2359);
or U2624 (N_2624,N_1602,N_1950);
or U2625 (N_2625,N_1316,N_1013);
and U2626 (N_2626,N_137,N_842);
nand U2627 (N_2627,N_2211,N_479);
or U2628 (N_2628,N_2423,N_1501);
or U2629 (N_2629,N_648,N_1582);
nand U2630 (N_2630,N_498,N_1575);
or U2631 (N_2631,N_350,N_162);
nand U2632 (N_2632,N_2106,N_300);
nand U2633 (N_2633,N_2077,N_1680);
or U2634 (N_2634,N_2184,N_936);
nand U2635 (N_2635,N_727,N_1045);
or U2636 (N_2636,N_1441,N_1285);
or U2637 (N_2637,N_262,N_333);
nor U2638 (N_2638,N_2326,N_2008);
nor U2639 (N_2639,N_2454,N_1936);
nor U2640 (N_2640,N_2070,N_1178);
nand U2641 (N_2641,N_401,N_1564);
xor U2642 (N_2642,N_1846,N_1268);
and U2643 (N_2643,N_242,N_714);
or U2644 (N_2644,N_1255,N_113);
xor U2645 (N_2645,N_1684,N_1817);
xor U2646 (N_2646,N_1337,N_1889);
nor U2647 (N_2647,N_2484,N_421);
nand U2648 (N_2648,N_1079,N_57);
or U2649 (N_2649,N_514,N_1853);
nand U2650 (N_2650,N_518,N_482);
or U2651 (N_2651,N_1196,N_271);
or U2652 (N_2652,N_276,N_155);
nor U2653 (N_2653,N_1445,N_1225);
nand U2654 (N_2654,N_1256,N_577);
nor U2655 (N_2655,N_701,N_564);
nor U2656 (N_2656,N_1463,N_2357);
and U2657 (N_2657,N_561,N_504);
nor U2658 (N_2658,N_1905,N_1651);
and U2659 (N_2659,N_2036,N_2177);
xor U2660 (N_2660,N_122,N_1585);
xnor U2661 (N_2661,N_897,N_1888);
nand U2662 (N_2662,N_1408,N_1175);
xor U2663 (N_2663,N_724,N_351);
nand U2664 (N_2664,N_211,N_671);
and U2665 (N_2665,N_991,N_377);
nand U2666 (N_2666,N_1610,N_744);
or U2667 (N_2667,N_761,N_1897);
or U2668 (N_2668,N_71,N_2048);
nor U2669 (N_2669,N_1996,N_1643);
nand U2670 (N_2670,N_230,N_194);
nor U2671 (N_2671,N_473,N_439);
nor U2672 (N_2672,N_2132,N_1644);
nor U2673 (N_2673,N_1822,N_2085);
nand U2674 (N_2674,N_321,N_1490);
nor U2675 (N_2675,N_501,N_1662);
xor U2676 (N_2676,N_318,N_767);
xor U2677 (N_2677,N_409,N_1334);
or U2678 (N_2678,N_1001,N_2327);
or U2679 (N_2679,N_328,N_2174);
nor U2680 (N_2680,N_1191,N_1413);
nand U2681 (N_2681,N_1839,N_576);
or U2682 (N_2682,N_1452,N_237);
and U2683 (N_2683,N_2348,N_1901);
nand U2684 (N_2684,N_2034,N_2355);
nor U2685 (N_2685,N_391,N_867);
or U2686 (N_2686,N_2005,N_85);
nand U2687 (N_2687,N_1903,N_2373);
nand U2688 (N_2688,N_306,N_1414);
and U2689 (N_2689,N_615,N_340);
nor U2690 (N_2690,N_1357,N_2430);
and U2691 (N_2691,N_1238,N_2025);
nor U2692 (N_2692,N_2315,N_726);
or U2693 (N_2693,N_1955,N_132);
and U2694 (N_2694,N_965,N_2449);
xnor U2695 (N_2695,N_1628,N_1946);
nor U2696 (N_2696,N_844,N_1161);
nand U2697 (N_2697,N_388,N_650);
nor U2698 (N_2698,N_1974,N_1537);
xnor U2699 (N_2699,N_646,N_1833);
nand U2700 (N_2700,N_1658,N_2240);
and U2701 (N_2701,N_2369,N_1234);
and U2702 (N_2702,N_1632,N_160);
or U2703 (N_2703,N_2097,N_1394);
nor U2704 (N_2704,N_639,N_13);
and U2705 (N_2705,N_1884,N_1384);
or U2706 (N_2706,N_847,N_720);
nor U2707 (N_2707,N_1150,N_525);
or U2708 (N_2708,N_1410,N_2149);
nand U2709 (N_2709,N_1713,N_1131);
and U2710 (N_2710,N_256,N_346);
and U2711 (N_2711,N_1925,N_2229);
nand U2712 (N_2712,N_1197,N_1868);
nand U2713 (N_2713,N_1138,N_116);
or U2714 (N_2714,N_1840,N_178);
xor U2715 (N_2715,N_133,N_112);
nand U2716 (N_2716,N_1479,N_1948);
xnor U2717 (N_2717,N_2495,N_1451);
and U2718 (N_2718,N_2385,N_1347);
nor U2719 (N_2719,N_123,N_218);
nand U2720 (N_2720,N_749,N_1552);
nor U2721 (N_2721,N_630,N_1751);
and U2722 (N_2722,N_418,N_1080);
nor U2723 (N_2723,N_2246,N_2311);
or U2724 (N_2724,N_772,N_1035);
nor U2725 (N_2725,N_1870,N_1792);
nand U2726 (N_2726,N_2403,N_179);
nor U2727 (N_2727,N_1560,N_1497);
xor U2728 (N_2728,N_1218,N_1094);
nand U2729 (N_2729,N_1217,N_924);
nand U2730 (N_2730,N_1465,N_2398);
or U2731 (N_2731,N_750,N_1143);
nor U2732 (N_2732,N_2394,N_1485);
nand U2733 (N_2733,N_2119,N_2076);
nor U2734 (N_2734,N_1442,N_895);
nor U2735 (N_2735,N_371,N_2056);
or U2736 (N_2736,N_1124,N_1504);
and U2737 (N_2737,N_294,N_2069);
or U2738 (N_2738,N_364,N_2039);
xor U2739 (N_2739,N_2087,N_1883);
nand U2740 (N_2740,N_169,N_1266);
and U2741 (N_2741,N_1388,N_1064);
xnor U2742 (N_2742,N_1542,N_466);
or U2743 (N_2743,N_1233,N_121);
xor U2744 (N_2744,N_2278,N_2455);
nand U2745 (N_2745,N_314,N_1496);
nand U2746 (N_2746,N_550,N_1062);
nand U2747 (N_2747,N_2288,N_1741);
or U2748 (N_2748,N_431,N_814);
nor U2749 (N_2749,N_913,N_1024);
nand U2750 (N_2750,N_1689,N_387);
nor U2751 (N_2751,N_437,N_950);
nor U2752 (N_2752,N_1406,N_1421);
nor U2753 (N_2753,N_669,N_2224);
nor U2754 (N_2754,N_1427,N_1787);
xor U2755 (N_2755,N_297,N_683);
nand U2756 (N_2756,N_385,N_1167);
nor U2757 (N_2757,N_2147,N_2109);
nor U2758 (N_2758,N_1142,N_915);
nand U2759 (N_2759,N_1698,N_1554);
and U2760 (N_2760,N_1721,N_2409);
nor U2761 (N_2761,N_390,N_2294);
or U2762 (N_2762,N_1104,N_1960);
or U2763 (N_2763,N_354,N_1916);
nor U2764 (N_2764,N_1180,N_828);
and U2765 (N_2765,N_1522,N_2464);
xor U2766 (N_2766,N_891,N_157);
xor U2767 (N_2767,N_1719,N_2165);
xor U2768 (N_2768,N_1227,N_6);
or U2769 (N_2769,N_1540,N_661);
nor U2770 (N_2770,N_130,N_2204);
and U2771 (N_2771,N_754,N_511);
xnor U2772 (N_2772,N_1710,N_1935);
xnor U2773 (N_2773,N_494,N_105);
or U2774 (N_2774,N_1170,N_806);
and U2775 (N_2775,N_1153,N_1892);
xnor U2776 (N_2776,N_49,N_2400);
nor U2777 (N_2777,N_545,N_1848);
xnor U2778 (N_2778,N_2286,N_1381);
xor U2779 (N_2779,N_1195,N_2052);
nand U2780 (N_2780,N_463,N_579);
xor U2781 (N_2781,N_1789,N_2350);
xor U2782 (N_2782,N_2159,N_777);
or U2783 (N_2783,N_1385,N_921);
xor U2784 (N_2784,N_1732,N_269);
xnor U2785 (N_2785,N_1364,N_344);
and U2786 (N_2786,N_2295,N_1887);
and U2787 (N_2787,N_19,N_2466);
nor U2788 (N_2788,N_900,N_841);
and U2789 (N_2789,N_1203,N_1857);
nor U2790 (N_2790,N_308,N_585);
xnor U2791 (N_2791,N_2459,N_699);
nand U2792 (N_2792,N_1404,N_277);
nor U2793 (N_2793,N_1919,N_1596);
or U2794 (N_2794,N_2401,N_1182);
and U2795 (N_2795,N_303,N_109);
and U2796 (N_2796,N_360,N_1184);
and U2797 (N_2797,N_1049,N_1924);
nand U2798 (N_2798,N_515,N_534);
nor U2799 (N_2799,N_1693,N_11);
nor U2800 (N_2800,N_356,N_1148);
or U2801 (N_2801,N_1980,N_1174);
nand U2802 (N_2802,N_503,N_667);
or U2803 (N_2803,N_1825,N_982);
or U2804 (N_2804,N_1516,N_912);
nor U2805 (N_2805,N_196,N_2480);
and U2806 (N_2806,N_2412,N_2437);
nand U2807 (N_2807,N_2482,N_2133);
xnor U2808 (N_2808,N_2485,N_436);
and U2809 (N_2809,N_643,N_1251);
or U2810 (N_2810,N_2117,N_1854);
nand U2811 (N_2811,N_792,N_1638);
or U2812 (N_2812,N_8,N_1829);
and U2813 (N_2813,N_863,N_1683);
or U2814 (N_2814,N_1056,N_2156);
and U2815 (N_2815,N_745,N_78);
and U2816 (N_2816,N_627,N_2230);
xnor U2817 (N_2817,N_1101,N_2095);
and U2818 (N_2818,N_2193,N_2298);
nor U2819 (N_2819,N_2170,N_2469);
or U2820 (N_2820,N_2264,N_2237);
nor U2821 (N_2821,N_1378,N_1566);
and U2822 (N_2822,N_2407,N_1011);
nand U2823 (N_2823,N_301,N_1937);
nor U2824 (N_2824,N_128,N_1577);
xnor U2825 (N_2825,N_30,N_601);
nor U2826 (N_2826,N_1893,N_143);
or U2827 (N_2827,N_1304,N_1539);
nor U2828 (N_2828,N_365,N_35);
xnor U2829 (N_2829,N_1014,N_488);
or U2830 (N_2830,N_688,N_198);
and U2831 (N_2831,N_311,N_389);
and U2832 (N_2832,N_2247,N_1000);
or U2833 (N_2833,N_568,N_2098);
xor U2834 (N_2834,N_1436,N_110);
or U2835 (N_2835,N_730,N_1863);
xor U2836 (N_2836,N_1674,N_2225);
or U2837 (N_2837,N_97,N_1754);
or U2838 (N_2838,N_1418,N_1878);
xor U2839 (N_2839,N_1922,N_1760);
xor U2840 (N_2840,N_2166,N_948);
nand U2841 (N_2841,N_1112,N_1951);
nand U2842 (N_2842,N_673,N_209);
or U2843 (N_2843,N_2171,N_119);
xor U2844 (N_2844,N_118,N_415);
or U2845 (N_2845,N_1269,N_784);
and U2846 (N_2846,N_1764,N_1277);
xnor U2847 (N_2847,N_1181,N_1252);
nand U2848 (N_2848,N_70,N_2141);
nand U2849 (N_2849,N_2404,N_1811);
nand U2850 (N_2850,N_695,N_378);
or U2851 (N_2851,N_1928,N_796);
or U2852 (N_2852,N_241,N_1111);
or U2853 (N_2853,N_961,N_848);
xnor U2854 (N_2854,N_1369,N_1550);
nor U2855 (N_2855,N_760,N_2364);
nand U2856 (N_2856,N_77,N_933);
nor U2857 (N_2857,N_1325,N_1289);
or U2858 (N_2858,N_2362,N_943);
nor U2859 (N_2859,N_1007,N_2094);
and U2860 (N_2860,N_743,N_575);
and U2861 (N_2861,N_625,N_213);
xnor U2862 (N_2862,N_1670,N_1093);
nor U2863 (N_2863,N_190,N_142);
and U2864 (N_2864,N_2091,N_2049);
nor U2865 (N_2865,N_2339,N_1726);
or U2866 (N_2866,N_894,N_837);
xnor U2867 (N_2867,N_5,N_2122);
nor U2868 (N_2868,N_292,N_1396);
nor U2869 (N_2869,N_947,N_1611);
and U2870 (N_2870,N_2448,N_679);
nand U2871 (N_2871,N_597,N_1561);
xnor U2872 (N_2872,N_539,N_1494);
nor U2873 (N_2873,N_316,N_412);
and U2874 (N_2874,N_697,N_124);
or U2875 (N_2875,N_138,N_1753);
nand U2876 (N_2876,N_535,N_2196);
or U2877 (N_2877,N_998,N_711);
xor U2878 (N_2878,N_247,N_670);
nand U2879 (N_2879,N_1842,N_2231);
xnor U2880 (N_2880,N_233,N_425);
xnor U2881 (N_2881,N_2410,N_634);
nor U2882 (N_2882,N_461,N_981);
and U2883 (N_2883,N_1030,N_1439);
and U2884 (N_2884,N_2358,N_92);
nor U2885 (N_2885,N_2243,N_1229);
and U2886 (N_2886,N_1351,N_2256);
or U2887 (N_2887,N_403,N_90);
or U2888 (N_2888,N_1959,N_2197);
and U2889 (N_2889,N_621,N_325);
or U2890 (N_2890,N_1834,N_21);
nor U2891 (N_2891,N_1348,N_1293);
nor U2892 (N_2892,N_2057,N_1376);
or U2893 (N_2893,N_846,N_820);
and U2894 (N_2894,N_1215,N_918);
xor U2895 (N_2895,N_1082,N_1222);
nor U2896 (N_2896,N_1701,N_657);
and U2897 (N_2897,N_1579,N_2372);
nand U2898 (N_2898,N_323,N_2379);
and U2899 (N_2899,N_1749,N_460);
nand U2900 (N_2900,N_1659,N_2351);
nor U2901 (N_2901,N_2429,N_275);
nor U2902 (N_2902,N_935,N_2274);
nor U2903 (N_2903,N_1686,N_1282);
and U2904 (N_2904,N_9,N_631);
or U2905 (N_2905,N_706,N_2282);
nor U2906 (N_2906,N_1291,N_956);
nor U2907 (N_2907,N_548,N_1652);
xor U2908 (N_2908,N_1483,N_249);
and U2909 (N_2909,N_452,N_239);
nor U2910 (N_2910,N_1295,N_873);
and U2911 (N_2911,N_1570,N_2107);
nand U2912 (N_2912,N_2150,N_2082);
or U2913 (N_2913,N_1627,N_1791);
nand U2914 (N_2914,N_2059,N_959);
xnor U2915 (N_2915,N_1294,N_938);
xnor U2916 (N_2916,N_259,N_2472);
nand U2917 (N_2917,N_1292,N_129);
xor U2918 (N_2918,N_1914,N_762);
or U2919 (N_2919,N_2065,N_64);
nor U2920 (N_2920,N_441,N_1041);
xor U2921 (N_2921,N_1341,N_516);
xor U2922 (N_2922,N_1654,N_941);
xnor U2923 (N_2923,N_1130,N_313);
or U2924 (N_2924,N_2227,N_1243);
xnor U2925 (N_2925,N_2354,N_2363);
nor U2926 (N_2926,N_512,N_2461);
nor U2927 (N_2927,N_972,N_1032);
and U2928 (N_2928,N_1038,N_544);
nand U2929 (N_2929,N_1874,N_293);
nor U2930 (N_2930,N_1164,N_214);
or U2931 (N_2931,N_1606,N_928);
nor U2932 (N_2932,N_1867,N_1144);
or U2933 (N_2933,N_2103,N_1391);
and U2934 (N_2934,N_2179,N_2038);
nand U2935 (N_2935,N_805,N_2279);
or U2936 (N_2936,N_2284,N_1474);
nor U2937 (N_2937,N_2062,N_1812);
xor U2938 (N_2938,N_1317,N_2276);
or U2939 (N_2939,N_2185,N_2478);
xor U2940 (N_2940,N_2233,N_2058);
xor U2941 (N_2941,N_1373,N_1089);
nor U2942 (N_2942,N_945,N_628);
nand U2943 (N_2943,N_1581,N_2218);
xor U2944 (N_2944,N_2389,N_1300);
or U2945 (N_2945,N_2341,N_1827);
xor U2946 (N_2946,N_1746,N_1116);
xnor U2947 (N_2947,N_1343,N_363);
nor U2948 (N_2948,N_1118,N_1372);
xor U2949 (N_2949,N_2411,N_99);
nor U2950 (N_2950,N_1583,N_1679);
or U2951 (N_2951,N_1530,N_2121);
nor U2952 (N_2952,N_2489,N_140);
xor U2953 (N_2953,N_1476,N_1318);
xnor U2954 (N_2954,N_335,N_1303);
xor U2955 (N_2955,N_1070,N_2089);
xnor U2956 (N_2956,N_1920,N_84);
or U2957 (N_2957,N_95,N_2436);
nand U2958 (N_2958,N_1042,N_2110);
xnor U2959 (N_2959,N_803,N_4);
nand U2960 (N_2960,N_651,N_822);
nand U2961 (N_2961,N_602,N_1250);
xnor U2962 (N_2962,N_624,N_1986);
xor U2963 (N_2963,N_1315,N_1083);
xnor U2964 (N_2964,N_148,N_1499);
nor U2965 (N_2965,N_2157,N_2380);
xnor U2966 (N_2966,N_1739,N_1425);
nand U2967 (N_2967,N_91,N_833);
nor U2968 (N_2968,N_1605,N_1122);
xor U2969 (N_2969,N_2381,N_2050);
or U2970 (N_2970,N_302,N_1879);
or U2971 (N_2971,N_2353,N_680);
or U2972 (N_2972,N_1068,N_1017);
and U2973 (N_2973,N_456,N_1660);
or U2974 (N_2974,N_1508,N_310);
nor U2975 (N_2975,N_339,N_849);
nor U2976 (N_2976,N_396,N_907);
and U2977 (N_2977,N_2467,N_1995);
nand U2978 (N_2978,N_619,N_816);
xor U2979 (N_2979,N_1616,N_888);
xnor U2980 (N_2980,N_1160,N_234);
nor U2981 (N_2981,N_979,N_766);
xnor U2982 (N_2982,N_2245,N_1194);
nor U2983 (N_2983,N_184,N_1488);
nor U2984 (N_2984,N_1352,N_1681);
and U2985 (N_2985,N_414,N_1482);
nor U2986 (N_2986,N_1119,N_1448);
xor U2987 (N_2987,N_2004,N_295);
or U2988 (N_2988,N_200,N_1498);
and U2989 (N_2989,N_1712,N_838);
nor U2990 (N_2990,N_776,N_1793);
or U2991 (N_2991,N_2374,N_15);
nand U2992 (N_2992,N_1063,N_382);
nand U2993 (N_2993,N_759,N_723);
nand U2994 (N_2994,N_315,N_875);
xor U2995 (N_2995,N_920,N_487);
nor U2996 (N_2996,N_2328,N_1779);
and U2997 (N_2997,N_2192,N_2061);
and U2998 (N_2998,N_940,N_2305);
xor U2999 (N_2999,N_977,N_2266);
nor U3000 (N_3000,N_1214,N_1966);
nor U3001 (N_3001,N_1908,N_1275);
or U3002 (N_3002,N_464,N_2064);
nor U3003 (N_3003,N_53,N_2386);
xor U3004 (N_3004,N_523,N_1139);
and U3005 (N_3005,N_1756,N_2222);
and U3006 (N_3006,N_1327,N_1661);
nor U3007 (N_3007,N_1043,N_1492);
and U3008 (N_3008,N_76,N_2477);
and U3009 (N_3009,N_2118,N_108);
or U3010 (N_3010,N_384,N_42);
nor U3011 (N_3011,N_1346,N_1154);
nand U3012 (N_3012,N_1345,N_1900);
xor U3013 (N_3013,N_1747,N_43);
nand U3014 (N_3014,N_2248,N_2301);
nor U3015 (N_3015,N_880,N_1306);
or U3016 (N_3016,N_158,N_2391);
xor U3017 (N_3017,N_61,N_1896);
and U3018 (N_3018,N_509,N_1424);
nand U3019 (N_3019,N_826,N_735);
and U3020 (N_3020,N_1665,N_1431);
nor U3021 (N_3021,N_1253,N_284);
or U3022 (N_3022,N_923,N_1675);
and U3023 (N_3023,N_600,N_36);
nand U3024 (N_3024,N_1858,N_153);
or U3025 (N_3025,N_2012,N_1037);
xnor U3026 (N_3026,N_2308,N_193);
or U3027 (N_3027,N_1095,N_380);
xor U3028 (N_3028,N_978,N_1515);
or U3029 (N_3029,N_282,N_2205);
or U3030 (N_3030,N_34,N_1190);
nand U3031 (N_3031,N_1307,N_645);
or U3032 (N_3032,N_2144,N_821);
nor U3033 (N_3033,N_582,N_1088);
nand U3034 (N_3034,N_1374,N_467);
nor U3035 (N_3035,N_2126,N_563);
nand U3036 (N_3036,N_1844,N_1664);
nand U3037 (N_3037,N_1949,N_1964);
or U3038 (N_3038,N_445,N_1395);
xor U3039 (N_3039,N_2383,N_1417);
or U3040 (N_3040,N_2242,N_1048);
nor U3041 (N_3041,N_995,N_555);
or U3042 (N_3042,N_1869,N_2138);
or U3043 (N_3043,N_2131,N_2015);
and U3044 (N_3044,N_1860,N_2425);
and U3045 (N_3045,N_1909,N_606);
or U3046 (N_3046,N_1899,N_1666);
nor U3047 (N_3047,N_1797,N_1895);
and U3048 (N_3048,N_1034,N_725);
or U3049 (N_3049,N_2151,N_892);
xor U3050 (N_3050,N_775,N_1267);
nor U3051 (N_3051,N_1028,N_580);
nand U3052 (N_3052,N_964,N_462);
nand U3053 (N_3053,N_1363,N_1305);
nand U3054 (N_3054,N_1818,N_2124);
nand U3055 (N_3055,N_672,N_1177);
nor U3056 (N_3056,N_652,N_2323);
xor U3057 (N_3057,N_1832,N_1473);
nor U3058 (N_3058,N_851,N_1531);
nand U3059 (N_3059,N_1375,N_1393);
and U3060 (N_3060,N_2388,N_868);
nor U3061 (N_3061,N_1387,N_2029);
or U3062 (N_3062,N_361,N_1769);
nand U3063 (N_3063,N_557,N_1904);
xor U3064 (N_3064,N_1379,N_2263);
nor U3065 (N_3065,N_272,N_207);
nor U3066 (N_3066,N_1962,N_1796);
and U3067 (N_3067,N_51,N_827);
and U3068 (N_3068,N_2152,N_188);
or U3069 (N_3069,N_1447,N_1625);
xor U3070 (N_3070,N_245,N_46);
xnor U3071 (N_3071,N_562,N_2261);
nand U3072 (N_3072,N_2120,N_1890);
or U3073 (N_3073,N_855,N_1804);
and U3074 (N_3074,N_1894,N_1005);
or U3075 (N_3075,N_1202,N_526);
or U3076 (N_3076,N_1505,N_1457);
xnor U3077 (N_3077,N_2271,N_2199);
nor U3078 (N_3078,N_134,N_1510);
or U3079 (N_3079,N_154,N_274);
xnor U3080 (N_3080,N_2215,N_1957);
xnor U3081 (N_3081,N_859,N_2476);
xnor U3082 (N_3082,N_689,N_2127);
or U3083 (N_3083,N_2285,N_1313);
and U3084 (N_3084,N_1529,N_329);
nor U3085 (N_3085,N_871,N_559);
nor U3086 (N_3086,N_107,N_428);
nor U3087 (N_3087,N_101,N_156);
or U3088 (N_3088,N_2447,N_1580);
and U3089 (N_3089,N_1368,N_1692);
xnor U3090 (N_3090,N_1830,N_1132);
and U3091 (N_3091,N_1423,N_1434);
xnor U3092 (N_3092,N_1273,N_963);
nand U3093 (N_3093,N_2283,N_352);
and U3094 (N_3094,N_716,N_1020);
nand U3095 (N_3095,N_1881,N_96);
xnor U3096 (N_3096,N_2273,N_1623);
nand U3097 (N_3097,N_1416,N_1731);
or U3098 (N_3098,N_1274,N_296);
and U3099 (N_3099,N_1814,N_696);
nor U3100 (N_3100,N_1547,N_934);
nand U3101 (N_3101,N_404,N_1135);
or U3102 (N_3102,N_560,N_32);
nor U3103 (N_3103,N_2128,N_2330);
nor U3104 (N_3104,N_1033,N_317);
nand U3105 (N_3105,N_2427,N_17);
and U3106 (N_3106,N_223,N_410);
nor U3107 (N_3107,N_2033,N_2035);
and U3108 (N_3108,N_1430,N_710);
or U3109 (N_3109,N_2130,N_1517);
xnor U3110 (N_3110,N_808,N_80);
nand U3111 (N_3111,N_2347,N_1403);
nand U3112 (N_3112,N_1961,N_131);
nand U3113 (N_3113,N_10,N_2458);
nand U3114 (N_3114,N_653,N_929);
nand U3115 (N_3115,N_203,N_746);
and U3116 (N_3116,N_738,N_1377);
nor U3117 (N_3117,N_287,N_599);
and U3118 (N_3118,N_1486,N_852);
xor U3119 (N_3119,N_1,N_864);
nor U3120 (N_3120,N_901,N_330);
xnor U3121 (N_3121,N_126,N_2182);
or U3122 (N_3122,N_861,N_1362);
nand U3123 (N_3123,N_117,N_2249);
xnor U3124 (N_3124,N_1535,N_1631);
xor U3125 (N_3125,N_970,N_1906);
and U3126 (N_3126,N_2014,N_1353);
nand U3127 (N_3127,N_44,N_866);
xor U3128 (N_3128,N_729,N_183);
nand U3129 (N_3129,N_1758,N_2220);
nand U3130 (N_3130,N_971,N_2203);
nor U3131 (N_3131,N_320,N_1489);
nand U3132 (N_3132,N_807,N_626);
xor U3133 (N_3133,N_406,N_1009);
nor U3134 (N_3134,N_208,N_1261);
xor U3135 (N_3135,N_1944,N_2470);
or U3136 (N_3136,N_1090,N_1568);
and U3137 (N_3137,N_2186,N_2016);
and U3138 (N_3138,N_2304,N_899);
or U3139 (N_3139,N_1735,N_986);
and U3140 (N_3140,N_63,N_270);
xor U3141 (N_3141,N_149,N_2306);
nor U3142 (N_3142,N_1736,N_1450);
nor U3143 (N_3143,N_783,N_106);
nor U3144 (N_3144,N_1390,N_997);
and U3145 (N_3145,N_2451,N_1994);
nand U3146 (N_3146,N_65,N_422);
nor U3147 (N_3147,N_2376,N_1750);
and U3148 (N_3148,N_362,N_2418);
and U3149 (N_3149,N_450,N_1271);
or U3150 (N_3150,N_593,N_2232);
or U3151 (N_3151,N_932,N_1555);
and U3152 (N_3152,N_719,N_1246);
xnor U3153 (N_3153,N_590,N_327);
nand U3154 (N_3154,N_1278,N_1836);
xor U3155 (N_3155,N_712,N_2079);
nand U3156 (N_3156,N_1549,N_780);
or U3157 (N_3157,N_2167,N_1682);
nand U3158 (N_3158,N_973,N_195);
nand U3159 (N_3159,N_416,N_1358);
xor U3160 (N_3160,N_1412,N_1471);
nor U3161 (N_3161,N_1943,N_2251);
and U3162 (N_3162,N_1397,N_2112);
nor U3163 (N_3163,N_1464,N_856);
nor U3164 (N_3164,N_1748,N_499);
nand U3165 (N_3165,N_147,N_2063);
and U3166 (N_3166,N_1134,N_1805);
nor U3167 (N_3167,N_2390,N_1074);
xnor U3168 (N_3168,N_1149,N_1730);
nand U3169 (N_3169,N_839,N_623);
nand U3170 (N_3170,N_120,N_1557);
and U3171 (N_3171,N_1113,N_707);
and U3172 (N_3172,N_1685,N_567);
and U3173 (N_3173,N_1040,N_1073);
xnor U3174 (N_3174,N_368,N_522);
or U3175 (N_3175,N_2377,N_1129);
nand U3176 (N_3176,N_309,N_469);
nand U3177 (N_3177,N_531,N_2491);
and U3178 (N_3178,N_94,N_2343);
and U3179 (N_3179,N_1121,N_261);
or U3180 (N_3180,N_1598,N_1865);
xnor U3181 (N_3181,N_553,N_1468);
or U3182 (N_3182,N_1367,N_1503);
nand U3183 (N_3183,N_433,N_1407);
and U3184 (N_3184,N_2433,N_226);
nand U3185 (N_3185,N_817,N_1563);
or U3186 (N_3186,N_1921,N_1286);
xor U3187 (N_3187,N_860,N_786);
nand U3188 (N_3188,N_800,N_1193);
nand U3189 (N_3189,N_2114,N_1487);
or U3190 (N_3190,N_1422,N_675);
xnor U3191 (N_3191,N_2268,N_1221);
nor U3192 (N_3192,N_740,N_1173);
or U3193 (N_3193,N_2161,N_870);
nand U3194 (N_3194,N_2223,N_1259);
and U3195 (N_3195,N_1287,N_399);
and U3196 (N_3196,N_2017,N_1224);
nor U3197 (N_3197,N_1567,N_2319);
nand U3198 (N_3198,N_1738,N_2023);
xnor U3199 (N_3199,N_2191,N_111);
nor U3200 (N_3200,N_1945,N_2235);
nor U3201 (N_3201,N_1990,N_1847);
and U3202 (N_3202,N_170,N_1553);
or U3203 (N_3203,N_769,N_1022);
nor U3204 (N_3204,N_2053,N_1475);
nor U3205 (N_3205,N_592,N_1622);
and U3206 (N_3206,N_765,N_1845);
or U3207 (N_3207,N_2275,N_2244);
nand U3208 (N_3208,N_2072,N_1199);
or U3209 (N_3209,N_1528,N_506);
xor U3210 (N_3210,N_969,N_1254);
and U3211 (N_3211,N_2486,N_1219);
and U3212 (N_3212,N_189,N_393);
xor U3213 (N_3213,N_1671,N_185);
xor U3214 (N_3214,N_2209,N_215);
nor U3215 (N_3215,N_1158,N_457);
or U3216 (N_3216,N_659,N_2420);
and U3217 (N_3217,N_812,N_283);
nor U3218 (N_3218,N_1072,N_1803);
xor U3219 (N_3219,N_1722,N_1010);
or U3220 (N_3220,N_2292,N_2145);
xnor U3221 (N_3221,N_1603,N_641);
nand U3222 (N_3222,N_2443,N_1650);
or U3223 (N_3223,N_1613,N_674);
nand U3224 (N_3224,N_2083,N_72);
nor U3225 (N_3225,N_1536,N_1975);
and U3226 (N_3226,N_2020,N_288);
nor U3227 (N_3227,N_82,N_647);
and U3228 (N_3228,N_2101,N_407);
xor U3229 (N_3229,N_1495,N_1521);
and U3230 (N_3230,N_558,N_2417);
nand U3231 (N_3231,N_319,N_210);
nand U3232 (N_3232,N_1782,N_2396);
or U3233 (N_3233,N_1281,N_908);
xnor U3234 (N_3234,N_644,N_3);
nor U3235 (N_3235,N_451,N_1023);
xnor U3236 (N_3236,N_1755,N_1724);
nand U3237 (N_3237,N_618,N_1071);
or U3238 (N_3238,N_1123,N_1856);
and U3239 (N_3239,N_2291,N_1128);
nand U3240 (N_3240,N_1084,N_1340);
or U3241 (N_3241,N_1044,N_1929);
nand U3242 (N_3242,N_2100,N_1861);
or U3243 (N_3243,N_1212,N_2287);
xnor U3244 (N_3244,N_2368,N_476);
and U3245 (N_3245,N_1389,N_2456);
nor U3246 (N_3246,N_1207,N_698);
nand U3247 (N_3247,N_2361,N_444);
and U3248 (N_3248,N_824,N_1003);
and U3249 (N_3249,N_718,N_1774);
nand U3250 (N_3250,N_1519,N_139);
nand U3251 (N_3251,N_960,N_637);
nand U3252 (N_3252,N_1871,N_1912);
xor U3253 (N_3253,N_458,N_1667);
nand U3254 (N_3254,N_1117,N_478);
and U3255 (N_3255,N_175,N_1270);
nor U3256 (N_3256,N_1469,N_45);
xor U3257 (N_3257,N_1541,N_2258);
or U3258 (N_3258,N_252,N_341);
and U3259 (N_3259,N_243,N_926);
and U3260 (N_3260,N_40,N_305);
or U3261 (N_3261,N_1607,N_2498);
nor U3262 (N_3262,N_1788,N_541);
or U3263 (N_3263,N_1015,N_1841);
nand U3264 (N_3264,N_1308,N_1366);
nor U3265 (N_3265,N_1299,N_773);
nor U3266 (N_3266,N_1444,N_589);
nor U3267 (N_3267,N_2297,N_165);
nand U3268 (N_3268,N_1969,N_2321);
nand U3269 (N_3269,N_2419,N_1077);
and U3270 (N_3270,N_2160,N_1402);
xor U3271 (N_3271,N_937,N_2086);
xor U3272 (N_3272,N_432,N_125);
nand U3273 (N_3273,N_1050,N_1910);
nand U3274 (N_3274,N_2473,N_353);
or U3275 (N_3275,N_52,N_2210);
nor U3276 (N_3276,N_622,N_755);
xor U3277 (N_3277,N_267,N_1877);
nor U3278 (N_3278,N_944,N_736);
nor U3279 (N_3279,N_1593,N_1875);
and U3280 (N_3280,N_2257,N_2302);
nand U3281 (N_3281,N_58,N_700);
xor U3282 (N_3282,N_74,N_1743);
xor U3283 (N_3283,N_2032,N_1330);
nand U3284 (N_3284,N_2183,N_538);
nand U3285 (N_3285,N_1763,N_885);
xor U3286 (N_3286,N_2493,N_2463);
nor U3287 (N_3287,N_2228,N_1771);
and U3288 (N_3288,N_980,N_1329);
and U3289 (N_3289,N_150,N_1723);
and U3290 (N_3290,N_1699,N_1838);
and U3291 (N_3291,N_612,N_2241);
and U3292 (N_3292,N_411,N_583);
or U3293 (N_3293,N_1614,N_658);
and U3294 (N_3294,N_1545,N_280);
nand U3295 (N_3295,N_1098,N_1586);
or U3296 (N_3296,N_232,N_264);
and U3297 (N_3297,N_2349,N_665);
nand U3298 (N_3298,N_2009,N_1176);
nor U3299 (N_3299,N_2113,N_1386);
xnor U3300 (N_3300,N_1344,N_1850);
nand U3301 (N_3301,N_611,N_468);
xnor U3302 (N_3302,N_2136,N_660);
nand U3303 (N_3303,N_1886,N_1562);
and U3304 (N_3304,N_1400,N_1106);
nor U3305 (N_3305,N_1314,N_829);
nand U3306 (N_3306,N_832,N_2336);
nor U3307 (N_3307,N_1051,N_1873);
and U3308 (N_3308,N_62,N_902);
and U3309 (N_3309,N_951,N_1941);
and U3310 (N_3310,N_1795,N_1157);
nand U3311 (N_3311,N_2024,N_2045);
xor U3312 (N_3312,N_88,N_1331);
nand U3313 (N_3313,N_434,N_50);
nand U3314 (N_3314,N_1599,N_2422);
nand U3315 (N_3315,N_235,N_2382);
and U3316 (N_3316,N_1882,N_797);
nor U3317 (N_3317,N_2115,N_2428);
and U3318 (N_3318,N_273,N_1572);
nor U3319 (N_3319,N_1851,N_990);
or U3320 (N_3320,N_2201,N_413);
xor U3321 (N_3321,N_1998,N_815);
nor U3322 (N_3322,N_1230,N_1239);
or U3323 (N_3323,N_2445,N_608);
xnor U3324 (N_3324,N_664,N_571);
nand U3325 (N_3325,N_151,N_666);
xor U3326 (N_3326,N_747,N_2395);
and U3327 (N_3327,N_910,N_565);
or U3328 (N_3328,N_757,N_1810);
nand U3329 (N_3329,N_2105,N_1806);
xor U3330 (N_3330,N_471,N_1707);
and U3331 (N_3331,N_1725,N_1970);
or U3332 (N_3332,N_1820,N_939);
nor U3333 (N_3333,N_603,N_1991);
and U3334 (N_3334,N_440,N_1232);
or U3335 (N_3335,N_27,N_2081);
and U3336 (N_3336,N_244,N_905);
nand U3337 (N_3337,N_332,N_1630);
nor U3338 (N_3338,N_2322,N_2468);
or U3339 (N_3339,N_1405,N_480);
or U3340 (N_3340,N_629,N_663);
or U3341 (N_3341,N_690,N_1205);
nand U3342 (N_3342,N_1008,N_1025);
nand U3343 (N_3343,N_2440,N_713);
nand U3344 (N_3344,N_1060,N_795);
nand U3345 (N_3345,N_446,N_694);
and U3346 (N_3346,N_722,N_197);
xnor U3347 (N_3347,N_876,N_781);
nor U3348 (N_3348,N_68,N_830);
nand U3349 (N_3349,N_2239,N_748);
or U3350 (N_3350,N_1636,N_168);
or U3351 (N_3351,N_1026,N_1165);
nor U3352 (N_3352,N_455,N_227);
nand U3353 (N_3353,N_1262,N_1697);
nand U3354 (N_3354,N_1608,N_1152);
and U3355 (N_3355,N_1716,N_2356);
nand U3356 (N_3356,N_2168,N_289);
or U3357 (N_3357,N_872,N_1752);
nor U3358 (N_3358,N_946,N_1783);
or U3359 (N_3359,N_1365,N_2494);
and U3360 (N_3360,N_383,N_2408);
nor U3361 (N_3361,N_1934,N_668);
nand U3362 (N_3362,N_1057,N_2188);
xor U3363 (N_3363,N_2046,N_1637);
and U3364 (N_3364,N_278,N_682);
xnor U3365 (N_3365,N_2099,N_1727);
nand U3366 (N_3366,N_999,N_31);
nor U3367 (N_3367,N_220,N_345);
xnor U3368 (N_3368,N_1126,N_453);
and U3369 (N_3369,N_2255,N_904);
nor U3370 (N_3370,N_2090,N_2352);
xnor U3371 (N_3371,N_1185,N_2402);
nand U3372 (N_3372,N_2010,N_1162);
or U3373 (N_3373,N_2318,N_2307);
nand U3374 (N_3374,N_16,N_1866);
or U3375 (N_3375,N_2206,N_1075);
or U3376 (N_3376,N_500,N_2123);
and U3377 (N_3377,N_1370,N_392);
xnor U3378 (N_3378,N_1102,N_367);
or U3379 (N_3379,N_1597,N_370);
xor U3380 (N_3380,N_1663,N_474);
xor U3381 (N_3381,N_1018,N_470);
xor U3382 (N_3382,N_1745,N_159);
nand U3383 (N_3383,N_349,N_224);
xnor U3384 (N_3384,N_887,N_492);
and U3385 (N_3385,N_532,N_1513);
or U3386 (N_3386,N_1507,N_1907);
nand U3387 (N_3387,N_942,N_1551);
and U3388 (N_3388,N_201,N_253);
nand U3389 (N_3389,N_790,N_465);
xnor U3390 (N_3390,N_2290,N_1478);
nor U3391 (N_3391,N_1046,N_931);
nand U3392 (N_3392,N_1004,N_2153);
nor U3393 (N_3393,N_379,N_2158);
nor U3394 (N_3394,N_1759,N_1454);
and U3395 (N_3395,N_2367,N_1321);
or U3396 (N_3396,N_1272,N_2414);
nand U3397 (N_3397,N_2142,N_167);
and U3398 (N_3398,N_281,N_566);
and U3399 (N_3399,N_472,N_1702);
nor U3400 (N_3400,N_2176,N_909);
xnor U3401 (N_3401,N_2019,N_779);
and U3402 (N_3402,N_604,N_192);
xnor U3403 (N_3403,N_1226,N_1956);
xnor U3404 (N_3404,N_75,N_1592);
nor U3405 (N_3405,N_1785,N_12);
xnor U3406 (N_3406,N_2277,N_1231);
xor U3407 (N_3407,N_322,N_570);
and U3408 (N_3408,N_1211,N_1695);
and U3409 (N_3409,N_1107,N_102);
and U3410 (N_3410,N_520,N_1978);
nor U3411 (N_3411,N_1704,N_2434);
and U3412 (N_3412,N_733,N_770);
and U3413 (N_3413,N_533,N_187);
and U3414 (N_3414,N_23,N_1356);
nand U3415 (N_3415,N_1669,N_893);
nor U3416 (N_3416,N_1216,N_2194);
nor U3417 (N_3417,N_1506,N_1283);
nor U3418 (N_3418,N_334,N_547);
and U3419 (N_3419,N_1257,N_2006);
and U3420 (N_3420,N_1574,N_2340);
and U3421 (N_3421,N_1114,N_751);
nand U3422 (N_3422,N_146,N_1775);
nor U3423 (N_3423,N_1078,N_426);
nor U3424 (N_3424,N_1065,N_1371);
and U3425 (N_3425,N_2021,N_1279);
nor U3426 (N_3426,N_1676,N_2325);
xnor U3427 (N_3427,N_1967,N_1718);
xnor U3428 (N_3428,N_358,N_2253);
nor U3429 (N_3429,N_2093,N_2462);
nand U3430 (N_3430,N_1824,N_2299);
or U3431 (N_3431,N_1958,N_1518);
nor U3432 (N_3432,N_1615,N_402);
nor U3433 (N_3433,N_1297,N_2441);
nor U3434 (N_3434,N_2397,N_2324);
nand U3435 (N_3435,N_1059,N_33);
nor U3436 (N_3436,N_1757,N_1245);
xnor U3437 (N_3437,N_1333,N_857);
xnor U3438 (N_3438,N_372,N_93);
and U3439 (N_3439,N_342,N_1171);
nand U3440 (N_3440,N_1136,N_1213);
xnor U3441 (N_3441,N_22,N_2406);
or U3442 (N_3442,N_975,N_958);
nor U3443 (N_3443,N_1819,N_1815);
nor U3444 (N_3444,N_862,N_1891);
xnor U3445 (N_3445,N_1428,N_1326);
xnor U3446 (N_3446,N_1913,N_2146);
and U3447 (N_3447,N_1831,N_588);
and U3448 (N_3448,N_831,N_1993);
or U3449 (N_3449,N_83,N_702);
xor U3450 (N_3450,N_238,N_1186);
and U3451 (N_3451,N_29,N_916);
or U3452 (N_3452,N_1105,N_1462);
or U3453 (N_3453,N_1989,N_100);
xor U3454 (N_3454,N_1923,N_610);
xor U3455 (N_3455,N_1236,N_2337);
or U3456 (N_3456,N_1872,N_1097);
nor U3457 (N_3457,N_481,N_2002);
nand U3458 (N_3458,N_836,N_1802);
and U3459 (N_3459,N_692,N_435);
nor U3460 (N_3460,N_1705,N_2092);
or U3461 (N_3461,N_89,N_181);
nor U3462 (N_3462,N_1715,N_2405);
xor U3463 (N_3463,N_573,N_843);
nor U3464 (N_3464,N_1355,N_1204);
nor U3465 (N_3465,N_1626,N_2169);
nor U3466 (N_3466,N_2439,N_596);
and U3467 (N_3467,N_2333,N_529);
nor U3468 (N_3468,N_1502,N_2479);
nor U3469 (N_3469,N_26,N_1125);
nand U3470 (N_3470,N_890,N_2424);
and U3471 (N_3471,N_1446,N_405);
nand U3472 (N_3472,N_2365,N_176);
nor U3473 (N_3473,N_1311,N_721);
or U3474 (N_3474,N_1241,N_1911);
and U3475 (N_3475,N_519,N_1527);
or U3476 (N_3476,N_1633,N_408);
and U3477 (N_3477,N_1141,N_1455);
or U3478 (N_3478,N_715,N_957);
nor U3479 (N_3479,N_86,N_2180);
xor U3480 (N_3480,N_2071,N_587);
xor U3481 (N_3481,N_447,N_540);
nor U3482 (N_3482,N_1360,N_299);
xor U3483 (N_3483,N_1794,N_172);
nand U3484 (N_3484,N_2338,N_1420);
xnor U3485 (N_3485,N_2499,N_804);
nor U3486 (N_3486,N_676,N_2096);
and U3487 (N_3487,N_2366,N_988);
nor U3488 (N_3488,N_260,N_1383);
xor U3489 (N_3489,N_1930,N_1336);
xor U3490 (N_3490,N_1350,N_424);
and U3491 (N_3491,N_1514,N_2000);
xnor U3492 (N_3492,N_1917,N_1151);
and U3493 (N_3493,N_2178,N_1999);
nand U3494 (N_3494,N_2055,N_2043);
xor U3495 (N_3495,N_756,N_1826);
and U3496 (N_3496,N_1159,N_1380);
xor U3497 (N_3497,N_2139,N_1511);
nor U3498 (N_3498,N_1480,N_914);
or U3499 (N_3499,N_1798,N_2148);
or U3500 (N_3500,N_1382,N_2488);
nand U3501 (N_3501,N_279,N_1189);
nor U3502 (N_3502,N_81,N_967);
nor U3503 (N_3503,N_1864,N_2164);
xnor U3504 (N_3504,N_265,N_2250);
nor U3505 (N_3505,N_1703,N_2346);
nor U3506 (N_3506,N_2415,N_569);
xor U3507 (N_3507,N_640,N_486);
and U3508 (N_3508,N_2344,N_1183);
nand U3509 (N_3509,N_1248,N_47);
or U3510 (N_3510,N_2028,N_258);
xnor U3511 (N_3511,N_1109,N_2134);
and U3512 (N_3512,N_1493,N_1729);
nand U3513 (N_3513,N_2,N_103);
and U3514 (N_3514,N_307,N_246);
nor U3515 (N_3515,N_2475,N_1284);
or U3516 (N_3516,N_802,N_2084);
and U3517 (N_3517,N_1801,N_1127);
and U3518 (N_3518,N_1398,N_2444);
and U3519 (N_3519,N_1594,N_1223);
xor U3520 (N_3520,N_752,N_1052);
xor U3521 (N_3521,N_2207,N_163);
xor U3522 (N_3522,N_1837,N_337);
xor U3523 (N_3523,N_2088,N_180);
or U3524 (N_3524,N_2073,N_1201);
nor U3525 (N_3525,N_442,N_793);
xnor U3526 (N_3526,N_216,N_810);
nor U3527 (N_3527,N_2384,N_1085);
or U3528 (N_3528,N_427,N_1773);
xnor U3529 (N_3529,N_1312,N_911);
or U3530 (N_3530,N_1461,N_1790);
nor U3531 (N_3531,N_24,N_2413);
or U3532 (N_3532,N_1456,N_38);
nor U3533 (N_3533,N_607,N_263);
and U3534 (N_3534,N_1601,N_1433);
nand U3535 (N_3535,N_987,N_202);
or U3536 (N_3536,N_268,N_1885);
nor U3537 (N_3537,N_2465,N_922);
nand U3538 (N_3538,N_1296,N_642);
xnor U3539 (N_3539,N_419,N_1932);
and U3540 (N_3540,N_1717,N_1629);
xor U3541 (N_3541,N_1249,N_1163);
xnor U3542 (N_3542,N_1021,N_152);
xnor U3543 (N_3543,N_1784,N_489);
nor U3544 (N_3544,N_1809,N_2078);
nand U3545 (N_3545,N_1687,N_1855);
or U3546 (N_3546,N_2234,N_2416);
nor U3547 (N_3547,N_1573,N_1813);
or U3548 (N_3548,N_2496,N_586);
or U3549 (N_3549,N_1512,N_127);
and U3550 (N_3550,N_459,N_1590);
nand U3551 (N_3551,N_1055,N_79);
nand U3552 (N_3552,N_177,N_2190);
and U3553 (N_3553,N_1902,N_1467);
xnor U3554 (N_3554,N_2435,N_1559);
nand U3555 (N_3555,N_1409,N_925);
nor U3556 (N_3556,N_1061,N_1620);
and U3557 (N_3557,N_2399,N_1984);
nor U3558 (N_3558,N_1288,N_2267);
xor U3559 (N_3559,N_171,N_638);
xnor U3560 (N_3560,N_2051,N_2446);
nand U3561 (N_3561,N_2259,N_1781);
nand U3562 (N_3562,N_1209,N_2474);
xnor U3563 (N_3563,N_430,N_1265);
xor U3564 (N_3564,N_2393,N_1976);
xnor U3565 (N_3565,N_1938,N_536);
and U3566 (N_3566,N_1108,N_1526);
xnor U3567 (N_3567,N_811,N_2457);
and U3568 (N_3568,N_834,N_212);
and U3569 (N_3569,N_2438,N_521);
xor U3570 (N_3570,N_98,N_1862);
xor U3571 (N_3571,N_517,N_2104);
nand U3572 (N_3572,N_2102,N_1799);
or U3573 (N_3573,N_818,N_1992);
and U3574 (N_3574,N_1210,N_373);
nor U3575 (N_3575,N_395,N_898);
nand U3576 (N_3576,N_2281,N_1997);
nand U3577 (N_3577,N_878,N_1429);
nand U3578 (N_3578,N_1192,N_1006);
nor U3579 (N_3579,N_1823,N_620);
and U3580 (N_3580,N_369,N_1646);
nor U3581 (N_3581,N_613,N_141);
nand U3582 (N_3582,N_1319,N_2007);
and U3583 (N_3583,N_1714,N_1500);
nand U3584 (N_3584,N_1096,N_2173);
nand U3585 (N_3585,N_927,N_581);
nor U3586 (N_3586,N_1963,N_1411);
or U3587 (N_3587,N_1534,N_2042);
and U3588 (N_3588,N_222,N_2213);
nor U3589 (N_3589,N_1954,N_551);
nand U3590 (N_3590,N_2080,N_1647);
and U3591 (N_3591,N_949,N_1533);
and U3592 (N_3592,N_2453,N_903);
xor U3593 (N_3593,N_1324,N_1339);
nor U3594 (N_3594,N_2041,N_1584);
nor U3595 (N_3595,N_2040,N_475);
and U3596 (N_3596,N_764,N_225);
and U3597 (N_3597,N_2313,N_2310);
or U3598 (N_3598,N_763,N_1742);
and U3599 (N_3599,N_703,N_930);
xnor U3600 (N_3600,N_823,N_2143);
and U3601 (N_3601,N_2293,N_338);
nand U3602 (N_3602,N_881,N_1466);
nor U3603 (N_3603,N_882,N_528);
nand U3604 (N_3604,N_554,N_375);
and U3605 (N_3605,N_1673,N_955);
or U3606 (N_3606,N_983,N_1438);
xnor U3607 (N_3607,N_145,N_1737);
xor U3608 (N_3608,N_705,N_2135);
or U3609 (N_3609,N_1440,N_2421);
and U3610 (N_3610,N_819,N_578);
or U3611 (N_3611,N_2172,N_1401);
nand U3612 (N_3612,N_1609,N_1765);
nor U3613 (N_3613,N_1852,N_906);
nor U3614 (N_3614,N_1426,N_753);
nand U3615 (N_3615,N_953,N_617);
nand U3616 (N_3616,N_2060,N_454);
nor U3617 (N_3617,N_2018,N_217);
or U3618 (N_3618,N_493,N_732);
and U3619 (N_3619,N_1926,N_1677);
nand U3620 (N_3620,N_2378,N_1915);
nand U3621 (N_3621,N_858,N_2067);
xnor U3622 (N_3622,N_1947,N_2309);
or U3623 (N_3623,N_240,N_483);
and U3624 (N_3624,N_2026,N_2129);
xnor U3625 (N_3625,N_1166,N_2116);
nor U3626 (N_3626,N_2195,N_693);
and U3627 (N_3627,N_1155,N_1843);
nor U3628 (N_3628,N_1392,N_1678);
or U3629 (N_3629,N_1538,N_73);
or U3630 (N_3630,N_1973,N_2269);
or U3631 (N_3631,N_835,N_374);
or U3632 (N_3632,N_2265,N_41);
xor U3633 (N_3633,N_1604,N_2431);
or U3634 (N_3634,N_2066,N_677);
nor U3635 (N_3635,N_251,N_572);
xnor U3636 (N_3636,N_1091,N_1939);
nand U3637 (N_3637,N_507,N_2212);
and U3638 (N_3638,N_1776,N_1460);
nor U3639 (N_3639,N_484,N_2219);
xnor U3640 (N_3640,N_1691,N_1302);
nand U3641 (N_3641,N_635,N_37);
nor U3642 (N_3642,N_1338,N_1653);
nand U3643 (N_3643,N_1777,N_2068);
and U3644 (N_3644,N_39,N_2460);
xnor U3645 (N_3645,N_2370,N_685);
and U3646 (N_3646,N_1029,N_1298);
and U3647 (N_3647,N_2262,N_1968);
xnor U3648 (N_3648,N_254,N_654);
nor U3649 (N_3649,N_1816,N_443);
or U3650 (N_3650,N_1058,N_1322);
or U3651 (N_3651,N_2345,N_556);
or U3652 (N_3652,N_1435,N_2471);
nor U3653 (N_3653,N_845,N_717);
and U3654 (N_3654,N_1168,N_1509);
nor U3655 (N_3655,N_687,N_1146);
or U3656 (N_3656,N_614,N_1432);
and U3657 (N_3657,N_917,N_741);
nor U3658 (N_3658,N_505,N_985);
xor U3659 (N_3659,N_174,N_1323);
and U3660 (N_3660,N_636,N_2022);
and U3661 (N_3661,N_1258,N_56);
or U3662 (N_3662,N_114,N_221);
and U3663 (N_3663,N_104,N_734);
nor U3664 (N_3664,N_1110,N_1067);
nor U3665 (N_3665,N_1115,N_59);
xnor U3666 (N_3666,N_2208,N_2221);
and U3667 (N_3667,N_1634,N_1309);
xor U3668 (N_3668,N_549,N_1076);
and U3669 (N_3669,N_66,N_595);
and U3670 (N_3670,N_1145,N_2270);
and U3671 (N_3671,N_1821,N_788);
and U3672 (N_3672,N_1310,N_2163);
nor U3673 (N_3673,N_678,N_584);
nand U3674 (N_3674,N_1709,N_2044);
nor U3675 (N_3675,N_1971,N_2317);
nand U3676 (N_3676,N_1657,N_2452);
or U3677 (N_3677,N_2054,N_2314);
and U3678 (N_3678,N_524,N_2187);
xor U3679 (N_3679,N_2111,N_1778);
or U3680 (N_3680,N_996,N_1244);
nor U3681 (N_3681,N_266,N_1443);
xor U3682 (N_3682,N_1668,N_366);
or U3683 (N_3683,N_2238,N_490);
xnor U3684 (N_3684,N_1708,N_2490);
xnor U3685 (N_3685,N_2001,N_787);
and U3686 (N_3686,N_1876,N_731);
nand U3687 (N_3687,N_2487,N_1880);
nor U3688 (N_3688,N_1808,N_546);
or U3689 (N_3689,N_1587,N_1081);
or U3690 (N_3690,N_228,N_2155);
or U3691 (N_3691,N_1556,N_1453);
nand U3692 (N_3692,N_1472,N_2387);
and U3693 (N_3693,N_485,N_1066);
xor U3694 (N_3694,N_2450,N_1012);
xnor U3695 (N_3695,N_20,N_1700);
nand U3696 (N_3696,N_250,N_2047);
and U3697 (N_3697,N_605,N_420);
or U3698 (N_3698,N_54,N_591);
or U3699 (N_3699,N_285,N_527);
nor U3700 (N_3700,N_1576,N_502);
xor U3701 (N_3701,N_742,N_18);
and U3702 (N_3702,N_1290,N_1835);
nand U3703 (N_3703,N_359,N_1931);
xnor U3704 (N_3704,N_1953,N_2214);
nand U3705 (N_3705,N_1768,N_1532);
nand U3706 (N_3706,N_709,N_2334);
nand U3707 (N_3707,N_1770,N_879);
xnor U3708 (N_3708,N_1047,N_1965);
xor U3709 (N_3709,N_1491,N_1019);
xor U3710 (N_3710,N_2316,N_1591);
nor U3711 (N_3711,N_1200,N_2198);
and U3712 (N_3712,N_2342,N_28);
nor U3713 (N_3713,N_1027,N_2181);
nor U3714 (N_3714,N_1569,N_1589);
nor U3715 (N_3715,N_684,N_1399);
xnor U3716 (N_3716,N_1642,N_1595);
nand U3717 (N_3717,N_0,N_1276);
xor U3718 (N_3718,N_633,N_2360);
xnor U3719 (N_3719,N_1172,N_1987);
and U3720 (N_3720,N_257,N_813);
nand U3721 (N_3721,N_1600,N_758);
or U3722 (N_3722,N_993,N_1179);
nor U3723 (N_3723,N_1780,N_782);
or U3724 (N_3724,N_2432,N_2140);
and U3725 (N_3725,N_889,N_2332);
and U3726 (N_3726,N_1927,N_1706);
nand U3727 (N_3727,N_1733,N_2031);
and U3728 (N_3728,N_1656,N_1361);
xor U3729 (N_3729,N_1419,N_1198);
and U3730 (N_3730,N_1565,N_298);
nand U3731 (N_3731,N_1016,N_55);
or U3732 (N_3732,N_1761,N_1481);
or U3733 (N_3733,N_530,N_655);
or U3734 (N_3734,N_1237,N_825);
and U3735 (N_3735,N_2289,N_1720);
nor U3736 (N_3736,N_2280,N_69);
xnor U3737 (N_3737,N_976,N_449);
and U3738 (N_3738,N_1206,N_968);
xnor U3739 (N_3739,N_865,N_681);
nor U3740 (N_3740,N_438,N_1942);
nor U3741 (N_3741,N_2108,N_2331);
or U3742 (N_3742,N_1054,N_164);
xnor U3743 (N_3743,N_2300,N_331);
nor U3744 (N_3744,N_704,N_662);
nor U3745 (N_3745,N_1639,N_491);
nand U3746 (N_3746,N_2497,N_2442);
or U3747 (N_3747,N_355,N_336);
xor U3748 (N_3748,N_954,N_397);
and U3749 (N_3749,N_1520,N_513);
nor U3750 (N_3750,N_610,N_1960);
and U3751 (N_3751,N_2204,N_565);
nor U3752 (N_3752,N_1242,N_2370);
and U3753 (N_3753,N_1259,N_1083);
or U3754 (N_3754,N_2245,N_657);
nand U3755 (N_3755,N_657,N_1602);
or U3756 (N_3756,N_1787,N_1084);
or U3757 (N_3757,N_1942,N_1822);
and U3758 (N_3758,N_236,N_255);
nand U3759 (N_3759,N_2436,N_1705);
nand U3760 (N_3760,N_2337,N_1506);
xor U3761 (N_3761,N_1289,N_332);
nand U3762 (N_3762,N_2258,N_893);
or U3763 (N_3763,N_1593,N_1569);
nand U3764 (N_3764,N_620,N_1702);
nor U3765 (N_3765,N_99,N_876);
and U3766 (N_3766,N_2127,N_2445);
nor U3767 (N_3767,N_947,N_908);
or U3768 (N_3768,N_96,N_631);
and U3769 (N_3769,N_1648,N_141);
and U3770 (N_3770,N_92,N_1564);
xor U3771 (N_3771,N_1865,N_658);
nand U3772 (N_3772,N_360,N_749);
or U3773 (N_3773,N_577,N_2362);
nand U3774 (N_3774,N_2357,N_2358);
xor U3775 (N_3775,N_126,N_600);
and U3776 (N_3776,N_1055,N_119);
nor U3777 (N_3777,N_413,N_2066);
or U3778 (N_3778,N_989,N_2012);
nor U3779 (N_3779,N_2100,N_500);
or U3780 (N_3780,N_1026,N_2029);
nor U3781 (N_3781,N_2326,N_1637);
and U3782 (N_3782,N_2081,N_1016);
and U3783 (N_3783,N_485,N_207);
and U3784 (N_3784,N_33,N_2415);
nor U3785 (N_3785,N_1216,N_2191);
and U3786 (N_3786,N_996,N_2367);
nor U3787 (N_3787,N_1172,N_1211);
and U3788 (N_3788,N_392,N_755);
nand U3789 (N_3789,N_324,N_1834);
or U3790 (N_3790,N_1597,N_226);
or U3791 (N_3791,N_525,N_178);
nand U3792 (N_3792,N_1118,N_308);
nand U3793 (N_3793,N_577,N_757);
and U3794 (N_3794,N_2383,N_1156);
nand U3795 (N_3795,N_1648,N_2027);
nand U3796 (N_3796,N_1942,N_1170);
or U3797 (N_3797,N_1363,N_1990);
nor U3798 (N_3798,N_138,N_978);
or U3799 (N_3799,N_1226,N_2244);
nor U3800 (N_3800,N_2353,N_2094);
xnor U3801 (N_3801,N_2019,N_690);
xnor U3802 (N_3802,N_6,N_76);
xnor U3803 (N_3803,N_1689,N_1038);
nor U3804 (N_3804,N_1418,N_1161);
nand U3805 (N_3805,N_1000,N_944);
and U3806 (N_3806,N_113,N_783);
and U3807 (N_3807,N_1622,N_1365);
and U3808 (N_3808,N_2302,N_1657);
xor U3809 (N_3809,N_354,N_1765);
xor U3810 (N_3810,N_2045,N_457);
and U3811 (N_3811,N_431,N_1905);
xnor U3812 (N_3812,N_449,N_1199);
and U3813 (N_3813,N_1397,N_2188);
nand U3814 (N_3814,N_1636,N_2136);
nor U3815 (N_3815,N_2113,N_733);
or U3816 (N_3816,N_2242,N_853);
or U3817 (N_3817,N_2356,N_599);
and U3818 (N_3818,N_2343,N_993);
or U3819 (N_3819,N_451,N_2441);
or U3820 (N_3820,N_748,N_1610);
xor U3821 (N_3821,N_763,N_1188);
and U3822 (N_3822,N_1490,N_954);
and U3823 (N_3823,N_603,N_152);
xor U3824 (N_3824,N_413,N_1322);
nor U3825 (N_3825,N_2056,N_2115);
or U3826 (N_3826,N_1393,N_477);
nand U3827 (N_3827,N_1881,N_1321);
and U3828 (N_3828,N_678,N_1692);
and U3829 (N_3829,N_197,N_2267);
nor U3830 (N_3830,N_263,N_1324);
and U3831 (N_3831,N_31,N_814);
or U3832 (N_3832,N_1631,N_46);
and U3833 (N_3833,N_521,N_1580);
and U3834 (N_3834,N_2347,N_152);
xor U3835 (N_3835,N_191,N_547);
and U3836 (N_3836,N_502,N_588);
and U3837 (N_3837,N_2286,N_1559);
and U3838 (N_3838,N_1705,N_1850);
nand U3839 (N_3839,N_116,N_2228);
or U3840 (N_3840,N_213,N_1172);
and U3841 (N_3841,N_2139,N_1186);
nand U3842 (N_3842,N_1610,N_1428);
nand U3843 (N_3843,N_337,N_2077);
nor U3844 (N_3844,N_515,N_1323);
xnor U3845 (N_3845,N_1844,N_326);
xor U3846 (N_3846,N_1650,N_789);
nor U3847 (N_3847,N_458,N_186);
nand U3848 (N_3848,N_339,N_1787);
and U3849 (N_3849,N_528,N_729);
xor U3850 (N_3850,N_985,N_1041);
nand U3851 (N_3851,N_1632,N_165);
and U3852 (N_3852,N_2110,N_1621);
nor U3853 (N_3853,N_1752,N_1797);
nor U3854 (N_3854,N_1674,N_1962);
and U3855 (N_3855,N_442,N_2000);
nand U3856 (N_3856,N_1075,N_856);
nand U3857 (N_3857,N_1739,N_235);
and U3858 (N_3858,N_284,N_1815);
nand U3859 (N_3859,N_640,N_451);
or U3860 (N_3860,N_1801,N_2131);
or U3861 (N_3861,N_2042,N_958);
nand U3862 (N_3862,N_1466,N_187);
nand U3863 (N_3863,N_1045,N_2210);
xnor U3864 (N_3864,N_930,N_1917);
xor U3865 (N_3865,N_1053,N_1846);
and U3866 (N_3866,N_110,N_840);
or U3867 (N_3867,N_1508,N_1211);
nor U3868 (N_3868,N_1239,N_452);
xor U3869 (N_3869,N_1455,N_397);
and U3870 (N_3870,N_307,N_413);
nor U3871 (N_3871,N_2009,N_2265);
or U3872 (N_3872,N_1424,N_1838);
xor U3873 (N_3873,N_187,N_664);
and U3874 (N_3874,N_1622,N_319);
xor U3875 (N_3875,N_393,N_742);
xnor U3876 (N_3876,N_685,N_6);
nand U3877 (N_3877,N_66,N_929);
nand U3878 (N_3878,N_476,N_1543);
nor U3879 (N_3879,N_1043,N_934);
and U3880 (N_3880,N_872,N_2056);
or U3881 (N_3881,N_140,N_2419);
and U3882 (N_3882,N_1425,N_2211);
and U3883 (N_3883,N_862,N_16);
nor U3884 (N_3884,N_2379,N_2385);
nor U3885 (N_3885,N_349,N_183);
and U3886 (N_3886,N_453,N_2295);
nand U3887 (N_3887,N_2252,N_2057);
or U3888 (N_3888,N_2358,N_1420);
xnor U3889 (N_3889,N_1602,N_1691);
xor U3890 (N_3890,N_99,N_892);
and U3891 (N_3891,N_1943,N_294);
and U3892 (N_3892,N_2033,N_64);
or U3893 (N_3893,N_336,N_1087);
nor U3894 (N_3894,N_20,N_200);
nand U3895 (N_3895,N_2125,N_983);
nand U3896 (N_3896,N_671,N_1952);
and U3897 (N_3897,N_1016,N_2303);
xnor U3898 (N_3898,N_2271,N_588);
and U3899 (N_3899,N_247,N_232);
or U3900 (N_3900,N_550,N_2094);
and U3901 (N_3901,N_1972,N_700);
nor U3902 (N_3902,N_1194,N_1849);
or U3903 (N_3903,N_1030,N_1582);
nand U3904 (N_3904,N_2079,N_804);
nor U3905 (N_3905,N_1791,N_1959);
xnor U3906 (N_3906,N_1884,N_1516);
nor U3907 (N_3907,N_1711,N_243);
or U3908 (N_3908,N_887,N_2070);
nor U3909 (N_3909,N_2452,N_2294);
or U3910 (N_3910,N_1477,N_2486);
and U3911 (N_3911,N_1473,N_2467);
or U3912 (N_3912,N_1848,N_595);
nor U3913 (N_3913,N_248,N_370);
xnor U3914 (N_3914,N_1823,N_1944);
or U3915 (N_3915,N_1693,N_560);
nor U3916 (N_3916,N_437,N_673);
nor U3917 (N_3917,N_1724,N_994);
and U3918 (N_3918,N_927,N_1727);
nand U3919 (N_3919,N_102,N_286);
and U3920 (N_3920,N_257,N_913);
nor U3921 (N_3921,N_794,N_1084);
or U3922 (N_3922,N_706,N_832);
and U3923 (N_3923,N_370,N_187);
nor U3924 (N_3924,N_2209,N_65);
or U3925 (N_3925,N_1831,N_1852);
or U3926 (N_3926,N_304,N_924);
nor U3927 (N_3927,N_1109,N_1127);
and U3928 (N_3928,N_1184,N_1646);
nor U3929 (N_3929,N_597,N_221);
xnor U3930 (N_3930,N_1198,N_484);
nand U3931 (N_3931,N_638,N_903);
xor U3932 (N_3932,N_2404,N_2060);
nor U3933 (N_3933,N_475,N_2184);
xnor U3934 (N_3934,N_790,N_1845);
xor U3935 (N_3935,N_1468,N_1615);
and U3936 (N_3936,N_354,N_1501);
xnor U3937 (N_3937,N_793,N_1722);
and U3938 (N_3938,N_1076,N_1867);
nor U3939 (N_3939,N_2274,N_1743);
nor U3940 (N_3940,N_835,N_2495);
nand U3941 (N_3941,N_682,N_624);
nor U3942 (N_3942,N_1938,N_69);
or U3943 (N_3943,N_2338,N_2250);
and U3944 (N_3944,N_967,N_833);
nor U3945 (N_3945,N_49,N_2177);
and U3946 (N_3946,N_229,N_787);
xor U3947 (N_3947,N_2139,N_699);
xnor U3948 (N_3948,N_713,N_1060);
or U3949 (N_3949,N_1168,N_985);
xnor U3950 (N_3950,N_191,N_1703);
or U3951 (N_3951,N_669,N_345);
nand U3952 (N_3952,N_932,N_607);
or U3953 (N_3953,N_2309,N_446);
xor U3954 (N_3954,N_1450,N_1243);
or U3955 (N_3955,N_382,N_635);
or U3956 (N_3956,N_452,N_699);
or U3957 (N_3957,N_2456,N_1711);
nand U3958 (N_3958,N_1409,N_80);
nand U3959 (N_3959,N_2314,N_1699);
and U3960 (N_3960,N_1647,N_2437);
or U3961 (N_3961,N_1611,N_225);
nor U3962 (N_3962,N_752,N_1548);
or U3963 (N_3963,N_315,N_1792);
xor U3964 (N_3964,N_2014,N_434);
or U3965 (N_3965,N_431,N_1157);
nand U3966 (N_3966,N_1838,N_2468);
and U3967 (N_3967,N_861,N_1940);
xnor U3968 (N_3968,N_2011,N_1168);
nand U3969 (N_3969,N_682,N_1424);
nand U3970 (N_3970,N_220,N_883);
and U3971 (N_3971,N_1521,N_1745);
xor U3972 (N_3972,N_1032,N_2198);
and U3973 (N_3973,N_357,N_463);
nor U3974 (N_3974,N_123,N_2489);
or U3975 (N_3975,N_1449,N_1886);
or U3976 (N_3976,N_1161,N_1250);
or U3977 (N_3977,N_1974,N_551);
and U3978 (N_3978,N_1183,N_159);
or U3979 (N_3979,N_2061,N_637);
nor U3980 (N_3980,N_1925,N_666);
xor U3981 (N_3981,N_783,N_1878);
xor U3982 (N_3982,N_2340,N_857);
nor U3983 (N_3983,N_774,N_194);
nand U3984 (N_3984,N_1392,N_1802);
xor U3985 (N_3985,N_2482,N_288);
or U3986 (N_3986,N_1984,N_965);
nand U3987 (N_3987,N_2003,N_1628);
or U3988 (N_3988,N_1487,N_2184);
and U3989 (N_3989,N_1659,N_1113);
nor U3990 (N_3990,N_1147,N_23);
nand U3991 (N_3991,N_399,N_1750);
or U3992 (N_3992,N_1022,N_2238);
and U3993 (N_3993,N_2440,N_60);
xnor U3994 (N_3994,N_1367,N_2293);
nor U3995 (N_3995,N_1988,N_1158);
nand U3996 (N_3996,N_498,N_703);
or U3997 (N_3997,N_176,N_178);
xor U3998 (N_3998,N_1461,N_278);
xnor U3999 (N_3999,N_1172,N_2238);
nor U4000 (N_4000,N_1157,N_1903);
and U4001 (N_4001,N_1232,N_1464);
xor U4002 (N_4002,N_2222,N_2267);
and U4003 (N_4003,N_1262,N_2006);
nor U4004 (N_4004,N_426,N_2373);
nor U4005 (N_4005,N_2413,N_1798);
and U4006 (N_4006,N_2340,N_1596);
nand U4007 (N_4007,N_405,N_1619);
nand U4008 (N_4008,N_180,N_2197);
and U4009 (N_4009,N_2109,N_2473);
xor U4010 (N_4010,N_676,N_446);
xnor U4011 (N_4011,N_2067,N_1616);
xor U4012 (N_4012,N_10,N_2011);
and U4013 (N_4013,N_1914,N_1168);
or U4014 (N_4014,N_1791,N_582);
xor U4015 (N_4015,N_2438,N_2225);
or U4016 (N_4016,N_757,N_11);
nor U4017 (N_4017,N_288,N_381);
and U4018 (N_4018,N_2285,N_1195);
nand U4019 (N_4019,N_2349,N_348);
nand U4020 (N_4020,N_1579,N_211);
and U4021 (N_4021,N_960,N_311);
nor U4022 (N_4022,N_301,N_394);
and U4023 (N_4023,N_415,N_2372);
xnor U4024 (N_4024,N_2301,N_842);
xnor U4025 (N_4025,N_520,N_1042);
xnor U4026 (N_4026,N_1868,N_1727);
or U4027 (N_4027,N_1828,N_1318);
and U4028 (N_4028,N_39,N_731);
nand U4029 (N_4029,N_385,N_171);
and U4030 (N_4030,N_417,N_1249);
and U4031 (N_4031,N_498,N_1436);
nand U4032 (N_4032,N_2381,N_2247);
nor U4033 (N_4033,N_710,N_73);
and U4034 (N_4034,N_1313,N_494);
xor U4035 (N_4035,N_2019,N_588);
and U4036 (N_4036,N_1534,N_1317);
nor U4037 (N_4037,N_89,N_264);
nand U4038 (N_4038,N_144,N_1686);
or U4039 (N_4039,N_2096,N_1383);
and U4040 (N_4040,N_2227,N_1462);
nor U4041 (N_4041,N_611,N_813);
nor U4042 (N_4042,N_1174,N_1028);
and U4043 (N_4043,N_578,N_1301);
nor U4044 (N_4044,N_1822,N_2431);
and U4045 (N_4045,N_599,N_1867);
xnor U4046 (N_4046,N_1478,N_1808);
nor U4047 (N_4047,N_1636,N_1074);
or U4048 (N_4048,N_2242,N_707);
xnor U4049 (N_4049,N_1705,N_368);
and U4050 (N_4050,N_1646,N_1787);
nand U4051 (N_4051,N_1753,N_1896);
nand U4052 (N_4052,N_340,N_1466);
nor U4053 (N_4053,N_993,N_2142);
and U4054 (N_4054,N_802,N_1186);
xor U4055 (N_4055,N_1984,N_2342);
and U4056 (N_4056,N_488,N_2412);
nand U4057 (N_4057,N_2067,N_938);
xnor U4058 (N_4058,N_2173,N_241);
nor U4059 (N_4059,N_895,N_17);
nor U4060 (N_4060,N_742,N_881);
or U4061 (N_4061,N_1091,N_177);
xnor U4062 (N_4062,N_1090,N_2210);
and U4063 (N_4063,N_532,N_816);
nor U4064 (N_4064,N_624,N_1409);
xor U4065 (N_4065,N_2146,N_142);
or U4066 (N_4066,N_836,N_881);
or U4067 (N_4067,N_2206,N_1868);
and U4068 (N_4068,N_2027,N_44);
or U4069 (N_4069,N_2407,N_2318);
and U4070 (N_4070,N_1702,N_577);
and U4071 (N_4071,N_1053,N_1240);
xor U4072 (N_4072,N_1807,N_123);
and U4073 (N_4073,N_1416,N_114);
and U4074 (N_4074,N_1050,N_2353);
or U4075 (N_4075,N_1403,N_1061);
or U4076 (N_4076,N_1003,N_1955);
or U4077 (N_4077,N_861,N_735);
or U4078 (N_4078,N_681,N_514);
nand U4079 (N_4079,N_1040,N_1407);
nor U4080 (N_4080,N_2234,N_2238);
and U4081 (N_4081,N_770,N_449);
and U4082 (N_4082,N_778,N_125);
nor U4083 (N_4083,N_1218,N_1252);
nor U4084 (N_4084,N_1118,N_2183);
nor U4085 (N_4085,N_529,N_1461);
nor U4086 (N_4086,N_2232,N_1431);
and U4087 (N_4087,N_1101,N_257);
and U4088 (N_4088,N_1851,N_1097);
xnor U4089 (N_4089,N_168,N_997);
nand U4090 (N_4090,N_1836,N_822);
nand U4091 (N_4091,N_2045,N_2252);
and U4092 (N_4092,N_484,N_1601);
xor U4093 (N_4093,N_1877,N_150);
or U4094 (N_4094,N_695,N_536);
xnor U4095 (N_4095,N_167,N_1050);
and U4096 (N_4096,N_1643,N_2370);
and U4097 (N_4097,N_1285,N_1933);
and U4098 (N_4098,N_1032,N_2378);
and U4099 (N_4099,N_2044,N_213);
nor U4100 (N_4100,N_556,N_2453);
xnor U4101 (N_4101,N_282,N_2040);
nand U4102 (N_4102,N_893,N_1993);
and U4103 (N_4103,N_1766,N_1167);
xnor U4104 (N_4104,N_233,N_1294);
nor U4105 (N_4105,N_2090,N_1511);
xnor U4106 (N_4106,N_829,N_1714);
xor U4107 (N_4107,N_1266,N_279);
and U4108 (N_4108,N_632,N_94);
and U4109 (N_4109,N_197,N_449);
and U4110 (N_4110,N_840,N_130);
xor U4111 (N_4111,N_1623,N_183);
nand U4112 (N_4112,N_1130,N_907);
xor U4113 (N_4113,N_2074,N_2155);
nor U4114 (N_4114,N_2466,N_2429);
xnor U4115 (N_4115,N_509,N_2371);
or U4116 (N_4116,N_2242,N_1995);
and U4117 (N_4117,N_1984,N_2020);
and U4118 (N_4118,N_346,N_928);
and U4119 (N_4119,N_1297,N_2106);
and U4120 (N_4120,N_2112,N_56);
and U4121 (N_4121,N_798,N_1839);
or U4122 (N_4122,N_1888,N_200);
nand U4123 (N_4123,N_2142,N_2476);
nor U4124 (N_4124,N_2484,N_2374);
and U4125 (N_4125,N_1295,N_1343);
and U4126 (N_4126,N_2010,N_1191);
xor U4127 (N_4127,N_1130,N_681);
or U4128 (N_4128,N_2443,N_1229);
nand U4129 (N_4129,N_1896,N_1021);
nand U4130 (N_4130,N_1045,N_231);
nor U4131 (N_4131,N_2226,N_2127);
nand U4132 (N_4132,N_1438,N_1708);
or U4133 (N_4133,N_1201,N_672);
xor U4134 (N_4134,N_2112,N_2132);
nand U4135 (N_4135,N_1499,N_318);
xnor U4136 (N_4136,N_1048,N_1374);
or U4137 (N_4137,N_1913,N_1454);
nor U4138 (N_4138,N_1403,N_2404);
nand U4139 (N_4139,N_2076,N_1076);
or U4140 (N_4140,N_553,N_253);
nand U4141 (N_4141,N_994,N_999);
and U4142 (N_4142,N_1042,N_986);
xnor U4143 (N_4143,N_836,N_1912);
nand U4144 (N_4144,N_1251,N_1916);
xor U4145 (N_4145,N_452,N_1561);
or U4146 (N_4146,N_1162,N_764);
xnor U4147 (N_4147,N_352,N_579);
or U4148 (N_4148,N_1326,N_1762);
nor U4149 (N_4149,N_1713,N_1838);
nand U4150 (N_4150,N_1000,N_1313);
xnor U4151 (N_4151,N_1654,N_2403);
nor U4152 (N_4152,N_1225,N_1796);
nor U4153 (N_4153,N_381,N_2241);
xor U4154 (N_4154,N_755,N_142);
or U4155 (N_4155,N_1370,N_1983);
xnor U4156 (N_4156,N_373,N_1240);
xor U4157 (N_4157,N_2134,N_418);
xor U4158 (N_4158,N_122,N_1332);
nor U4159 (N_4159,N_2305,N_1428);
nor U4160 (N_4160,N_2007,N_1314);
nand U4161 (N_4161,N_350,N_508);
and U4162 (N_4162,N_1672,N_386);
nand U4163 (N_4163,N_925,N_1570);
and U4164 (N_4164,N_1229,N_129);
nor U4165 (N_4165,N_137,N_2368);
or U4166 (N_4166,N_606,N_580);
xor U4167 (N_4167,N_809,N_1173);
and U4168 (N_4168,N_2487,N_1708);
nor U4169 (N_4169,N_2468,N_2035);
or U4170 (N_4170,N_698,N_994);
xnor U4171 (N_4171,N_1019,N_428);
and U4172 (N_4172,N_1417,N_1603);
nor U4173 (N_4173,N_1242,N_89);
xnor U4174 (N_4174,N_608,N_1194);
xnor U4175 (N_4175,N_1794,N_706);
and U4176 (N_4176,N_132,N_2100);
nand U4177 (N_4177,N_2257,N_2015);
xnor U4178 (N_4178,N_35,N_77);
nand U4179 (N_4179,N_254,N_2172);
nand U4180 (N_4180,N_33,N_474);
nand U4181 (N_4181,N_1007,N_2461);
and U4182 (N_4182,N_2278,N_397);
nor U4183 (N_4183,N_700,N_1461);
and U4184 (N_4184,N_892,N_330);
nand U4185 (N_4185,N_861,N_2142);
xnor U4186 (N_4186,N_1564,N_990);
nor U4187 (N_4187,N_988,N_321);
nand U4188 (N_4188,N_1925,N_146);
or U4189 (N_4189,N_849,N_1458);
xnor U4190 (N_4190,N_234,N_286);
and U4191 (N_4191,N_100,N_1618);
nor U4192 (N_4192,N_1025,N_1997);
nor U4193 (N_4193,N_1056,N_1453);
and U4194 (N_4194,N_1310,N_749);
or U4195 (N_4195,N_1178,N_898);
and U4196 (N_4196,N_747,N_2408);
and U4197 (N_4197,N_1312,N_628);
or U4198 (N_4198,N_2274,N_550);
nand U4199 (N_4199,N_2362,N_556);
nand U4200 (N_4200,N_1014,N_199);
nand U4201 (N_4201,N_494,N_2361);
xnor U4202 (N_4202,N_1757,N_1593);
nand U4203 (N_4203,N_718,N_248);
xnor U4204 (N_4204,N_734,N_883);
and U4205 (N_4205,N_2273,N_815);
nor U4206 (N_4206,N_335,N_1109);
nor U4207 (N_4207,N_89,N_184);
or U4208 (N_4208,N_23,N_2436);
nor U4209 (N_4209,N_150,N_111);
xnor U4210 (N_4210,N_1857,N_2498);
nand U4211 (N_4211,N_1505,N_210);
or U4212 (N_4212,N_286,N_1336);
and U4213 (N_4213,N_2227,N_517);
and U4214 (N_4214,N_1757,N_69);
and U4215 (N_4215,N_1866,N_79);
nand U4216 (N_4216,N_614,N_1471);
and U4217 (N_4217,N_2346,N_499);
and U4218 (N_4218,N_1729,N_746);
nand U4219 (N_4219,N_1449,N_286);
xor U4220 (N_4220,N_1835,N_1183);
xnor U4221 (N_4221,N_697,N_2201);
nor U4222 (N_4222,N_1524,N_965);
or U4223 (N_4223,N_1216,N_1534);
xor U4224 (N_4224,N_2165,N_1948);
or U4225 (N_4225,N_467,N_582);
and U4226 (N_4226,N_2470,N_1596);
xnor U4227 (N_4227,N_1100,N_1023);
and U4228 (N_4228,N_1080,N_2019);
xor U4229 (N_4229,N_989,N_690);
nand U4230 (N_4230,N_745,N_281);
or U4231 (N_4231,N_1042,N_1035);
nand U4232 (N_4232,N_1696,N_475);
nand U4233 (N_4233,N_2145,N_381);
nand U4234 (N_4234,N_269,N_839);
nor U4235 (N_4235,N_1408,N_242);
and U4236 (N_4236,N_1454,N_54);
and U4237 (N_4237,N_2081,N_1559);
and U4238 (N_4238,N_1873,N_1954);
and U4239 (N_4239,N_166,N_1150);
nor U4240 (N_4240,N_696,N_444);
nand U4241 (N_4241,N_2112,N_1587);
nand U4242 (N_4242,N_2400,N_1250);
and U4243 (N_4243,N_1902,N_1322);
xor U4244 (N_4244,N_1317,N_2205);
nor U4245 (N_4245,N_1986,N_642);
nor U4246 (N_4246,N_248,N_1734);
and U4247 (N_4247,N_886,N_876);
nand U4248 (N_4248,N_595,N_1539);
and U4249 (N_4249,N_1913,N_1839);
xnor U4250 (N_4250,N_1838,N_2146);
xnor U4251 (N_4251,N_1038,N_117);
xor U4252 (N_4252,N_605,N_538);
or U4253 (N_4253,N_2176,N_565);
nor U4254 (N_4254,N_1862,N_701);
nor U4255 (N_4255,N_1315,N_1988);
nor U4256 (N_4256,N_2371,N_799);
and U4257 (N_4257,N_2395,N_60);
nor U4258 (N_4258,N_850,N_1772);
and U4259 (N_4259,N_1234,N_2162);
and U4260 (N_4260,N_1642,N_2111);
nand U4261 (N_4261,N_303,N_2287);
nand U4262 (N_4262,N_1610,N_2132);
and U4263 (N_4263,N_1342,N_828);
nand U4264 (N_4264,N_1815,N_199);
nor U4265 (N_4265,N_345,N_1252);
and U4266 (N_4266,N_3,N_676);
nor U4267 (N_4267,N_1789,N_1521);
nor U4268 (N_4268,N_1577,N_1266);
or U4269 (N_4269,N_2035,N_1988);
xor U4270 (N_4270,N_137,N_1490);
or U4271 (N_4271,N_2455,N_285);
and U4272 (N_4272,N_2326,N_583);
or U4273 (N_4273,N_1733,N_1171);
nand U4274 (N_4274,N_2398,N_1209);
or U4275 (N_4275,N_2172,N_519);
or U4276 (N_4276,N_1910,N_1149);
nand U4277 (N_4277,N_2047,N_2072);
nor U4278 (N_4278,N_1180,N_1717);
nor U4279 (N_4279,N_582,N_1106);
and U4280 (N_4280,N_1586,N_1450);
nand U4281 (N_4281,N_2027,N_2054);
xor U4282 (N_4282,N_616,N_657);
or U4283 (N_4283,N_445,N_1651);
or U4284 (N_4284,N_1258,N_1143);
xor U4285 (N_4285,N_1667,N_381);
xnor U4286 (N_4286,N_2193,N_1034);
xor U4287 (N_4287,N_617,N_205);
and U4288 (N_4288,N_1491,N_1805);
nand U4289 (N_4289,N_2300,N_997);
nand U4290 (N_4290,N_1742,N_710);
or U4291 (N_4291,N_1395,N_1046);
and U4292 (N_4292,N_2135,N_567);
and U4293 (N_4293,N_1231,N_171);
and U4294 (N_4294,N_2324,N_1823);
and U4295 (N_4295,N_876,N_1374);
xor U4296 (N_4296,N_392,N_813);
nor U4297 (N_4297,N_2273,N_174);
xor U4298 (N_4298,N_416,N_2291);
nand U4299 (N_4299,N_332,N_602);
nor U4300 (N_4300,N_2075,N_550);
nand U4301 (N_4301,N_2390,N_1639);
nor U4302 (N_4302,N_277,N_1103);
xor U4303 (N_4303,N_142,N_263);
nand U4304 (N_4304,N_1178,N_845);
or U4305 (N_4305,N_344,N_97);
nor U4306 (N_4306,N_1064,N_1);
nand U4307 (N_4307,N_448,N_250);
xnor U4308 (N_4308,N_683,N_1194);
nand U4309 (N_4309,N_569,N_715);
xnor U4310 (N_4310,N_2336,N_472);
xor U4311 (N_4311,N_1065,N_873);
xor U4312 (N_4312,N_298,N_639);
xor U4313 (N_4313,N_2087,N_2158);
or U4314 (N_4314,N_2498,N_2270);
nor U4315 (N_4315,N_2249,N_1713);
xnor U4316 (N_4316,N_1852,N_1654);
or U4317 (N_4317,N_2019,N_1630);
nor U4318 (N_4318,N_2340,N_941);
and U4319 (N_4319,N_1256,N_1658);
or U4320 (N_4320,N_810,N_874);
or U4321 (N_4321,N_2123,N_2057);
nand U4322 (N_4322,N_151,N_585);
xor U4323 (N_4323,N_772,N_117);
nand U4324 (N_4324,N_1508,N_1283);
and U4325 (N_4325,N_2495,N_1606);
and U4326 (N_4326,N_1352,N_628);
nand U4327 (N_4327,N_774,N_2352);
and U4328 (N_4328,N_1051,N_2191);
xor U4329 (N_4329,N_1285,N_524);
or U4330 (N_4330,N_1414,N_1282);
nor U4331 (N_4331,N_178,N_310);
and U4332 (N_4332,N_346,N_39);
xor U4333 (N_4333,N_785,N_601);
nand U4334 (N_4334,N_137,N_1002);
nor U4335 (N_4335,N_1478,N_2217);
and U4336 (N_4336,N_2084,N_2214);
and U4337 (N_4337,N_1277,N_2343);
and U4338 (N_4338,N_1292,N_1741);
and U4339 (N_4339,N_423,N_767);
nor U4340 (N_4340,N_1428,N_2447);
and U4341 (N_4341,N_842,N_2457);
or U4342 (N_4342,N_363,N_1512);
or U4343 (N_4343,N_599,N_278);
nor U4344 (N_4344,N_1977,N_1601);
nand U4345 (N_4345,N_286,N_1111);
or U4346 (N_4346,N_319,N_1722);
nand U4347 (N_4347,N_1435,N_1164);
xnor U4348 (N_4348,N_811,N_145);
or U4349 (N_4349,N_346,N_1288);
and U4350 (N_4350,N_1886,N_299);
nor U4351 (N_4351,N_1322,N_1408);
and U4352 (N_4352,N_362,N_2281);
nand U4353 (N_4353,N_1733,N_2213);
nor U4354 (N_4354,N_2346,N_1908);
xnor U4355 (N_4355,N_1744,N_2048);
or U4356 (N_4356,N_944,N_946);
nor U4357 (N_4357,N_1179,N_458);
nor U4358 (N_4358,N_1746,N_2009);
and U4359 (N_4359,N_2348,N_1179);
and U4360 (N_4360,N_252,N_247);
nand U4361 (N_4361,N_2450,N_296);
xnor U4362 (N_4362,N_1111,N_1061);
nand U4363 (N_4363,N_244,N_1539);
nand U4364 (N_4364,N_2339,N_1330);
nor U4365 (N_4365,N_1070,N_383);
nand U4366 (N_4366,N_167,N_1150);
xor U4367 (N_4367,N_2216,N_59);
nand U4368 (N_4368,N_1627,N_2027);
and U4369 (N_4369,N_1893,N_1353);
nor U4370 (N_4370,N_471,N_2174);
nand U4371 (N_4371,N_1919,N_1923);
nand U4372 (N_4372,N_1943,N_315);
and U4373 (N_4373,N_1059,N_172);
nand U4374 (N_4374,N_1774,N_1447);
nand U4375 (N_4375,N_541,N_1400);
or U4376 (N_4376,N_407,N_195);
nand U4377 (N_4377,N_598,N_1778);
or U4378 (N_4378,N_861,N_1107);
xnor U4379 (N_4379,N_1647,N_2301);
xnor U4380 (N_4380,N_930,N_959);
or U4381 (N_4381,N_2305,N_426);
nor U4382 (N_4382,N_1484,N_870);
or U4383 (N_4383,N_1268,N_1319);
nand U4384 (N_4384,N_420,N_857);
nor U4385 (N_4385,N_36,N_1034);
nor U4386 (N_4386,N_2044,N_2381);
and U4387 (N_4387,N_557,N_1689);
nand U4388 (N_4388,N_1040,N_1251);
or U4389 (N_4389,N_1205,N_1173);
xor U4390 (N_4390,N_330,N_947);
xor U4391 (N_4391,N_695,N_574);
and U4392 (N_4392,N_1145,N_1849);
or U4393 (N_4393,N_576,N_1313);
xor U4394 (N_4394,N_1142,N_2309);
nor U4395 (N_4395,N_979,N_2438);
nor U4396 (N_4396,N_1696,N_2089);
nand U4397 (N_4397,N_1520,N_93);
nand U4398 (N_4398,N_425,N_1711);
nand U4399 (N_4399,N_630,N_1471);
or U4400 (N_4400,N_1917,N_1363);
nand U4401 (N_4401,N_617,N_1292);
xor U4402 (N_4402,N_1791,N_202);
nor U4403 (N_4403,N_1399,N_2475);
nand U4404 (N_4404,N_228,N_411);
and U4405 (N_4405,N_1102,N_2013);
nand U4406 (N_4406,N_2096,N_2063);
xnor U4407 (N_4407,N_1269,N_458);
or U4408 (N_4408,N_748,N_1933);
or U4409 (N_4409,N_1468,N_466);
nand U4410 (N_4410,N_343,N_451);
or U4411 (N_4411,N_1797,N_1182);
nand U4412 (N_4412,N_1311,N_545);
nor U4413 (N_4413,N_586,N_1580);
or U4414 (N_4414,N_1853,N_707);
xnor U4415 (N_4415,N_1986,N_2480);
nor U4416 (N_4416,N_2183,N_1751);
nor U4417 (N_4417,N_1821,N_475);
nand U4418 (N_4418,N_1646,N_1570);
xnor U4419 (N_4419,N_133,N_1662);
nand U4420 (N_4420,N_1549,N_1101);
nor U4421 (N_4421,N_1511,N_1814);
nand U4422 (N_4422,N_134,N_1005);
nand U4423 (N_4423,N_1748,N_2024);
nand U4424 (N_4424,N_758,N_717);
xor U4425 (N_4425,N_66,N_586);
nor U4426 (N_4426,N_55,N_1754);
nand U4427 (N_4427,N_2313,N_200);
nor U4428 (N_4428,N_308,N_2483);
nor U4429 (N_4429,N_1059,N_1148);
xor U4430 (N_4430,N_359,N_2061);
or U4431 (N_4431,N_2160,N_2050);
nand U4432 (N_4432,N_756,N_2159);
nor U4433 (N_4433,N_2004,N_365);
or U4434 (N_4434,N_1813,N_2343);
nor U4435 (N_4435,N_1657,N_364);
and U4436 (N_4436,N_46,N_1432);
nor U4437 (N_4437,N_1763,N_2139);
and U4438 (N_4438,N_39,N_1608);
xnor U4439 (N_4439,N_1586,N_1163);
xnor U4440 (N_4440,N_1532,N_1181);
and U4441 (N_4441,N_350,N_2351);
xor U4442 (N_4442,N_40,N_150);
xnor U4443 (N_4443,N_2290,N_1392);
xor U4444 (N_4444,N_937,N_877);
nor U4445 (N_4445,N_689,N_922);
or U4446 (N_4446,N_1494,N_1511);
and U4447 (N_4447,N_133,N_1503);
nand U4448 (N_4448,N_324,N_26);
or U4449 (N_4449,N_1008,N_791);
xor U4450 (N_4450,N_1682,N_519);
and U4451 (N_4451,N_1726,N_316);
xnor U4452 (N_4452,N_1214,N_1394);
nand U4453 (N_4453,N_78,N_2025);
xnor U4454 (N_4454,N_1342,N_2471);
nor U4455 (N_4455,N_47,N_945);
xor U4456 (N_4456,N_45,N_2115);
and U4457 (N_4457,N_1761,N_1737);
nor U4458 (N_4458,N_678,N_1104);
nor U4459 (N_4459,N_1065,N_1330);
nor U4460 (N_4460,N_1482,N_478);
nand U4461 (N_4461,N_175,N_167);
nor U4462 (N_4462,N_421,N_1086);
nor U4463 (N_4463,N_1628,N_1034);
and U4464 (N_4464,N_2401,N_487);
nand U4465 (N_4465,N_932,N_1801);
and U4466 (N_4466,N_2230,N_2337);
and U4467 (N_4467,N_605,N_666);
or U4468 (N_4468,N_711,N_176);
nor U4469 (N_4469,N_1691,N_697);
and U4470 (N_4470,N_2466,N_104);
or U4471 (N_4471,N_179,N_497);
nor U4472 (N_4472,N_763,N_1291);
nand U4473 (N_4473,N_2492,N_1679);
nor U4474 (N_4474,N_891,N_941);
xnor U4475 (N_4475,N_1118,N_2214);
nand U4476 (N_4476,N_2278,N_1802);
nand U4477 (N_4477,N_617,N_1675);
nand U4478 (N_4478,N_856,N_933);
or U4479 (N_4479,N_1643,N_97);
or U4480 (N_4480,N_1991,N_2319);
nor U4481 (N_4481,N_605,N_1598);
nor U4482 (N_4482,N_626,N_1963);
nor U4483 (N_4483,N_1234,N_733);
xor U4484 (N_4484,N_2483,N_97);
nor U4485 (N_4485,N_1986,N_2308);
and U4486 (N_4486,N_2254,N_2089);
nor U4487 (N_4487,N_1983,N_392);
or U4488 (N_4488,N_1271,N_504);
and U4489 (N_4489,N_1879,N_2222);
and U4490 (N_4490,N_1315,N_2266);
or U4491 (N_4491,N_2215,N_428);
or U4492 (N_4492,N_1588,N_1019);
xor U4493 (N_4493,N_1929,N_1023);
nand U4494 (N_4494,N_1430,N_1654);
xor U4495 (N_4495,N_1828,N_1608);
and U4496 (N_4496,N_360,N_584);
xor U4497 (N_4497,N_1051,N_491);
or U4498 (N_4498,N_1711,N_231);
and U4499 (N_4499,N_693,N_308);
and U4500 (N_4500,N_42,N_2398);
or U4501 (N_4501,N_458,N_363);
and U4502 (N_4502,N_1342,N_1532);
nand U4503 (N_4503,N_2077,N_859);
nor U4504 (N_4504,N_1915,N_1158);
and U4505 (N_4505,N_475,N_233);
and U4506 (N_4506,N_2283,N_1257);
xor U4507 (N_4507,N_1388,N_1231);
nand U4508 (N_4508,N_783,N_1674);
nor U4509 (N_4509,N_1639,N_134);
nand U4510 (N_4510,N_1365,N_1969);
and U4511 (N_4511,N_272,N_2217);
xor U4512 (N_4512,N_1161,N_1168);
xor U4513 (N_4513,N_751,N_1601);
and U4514 (N_4514,N_1119,N_957);
or U4515 (N_4515,N_1838,N_650);
nand U4516 (N_4516,N_1662,N_656);
or U4517 (N_4517,N_1505,N_2251);
nor U4518 (N_4518,N_338,N_1966);
xnor U4519 (N_4519,N_923,N_1346);
xor U4520 (N_4520,N_1090,N_399);
and U4521 (N_4521,N_1186,N_1457);
xor U4522 (N_4522,N_280,N_924);
nor U4523 (N_4523,N_364,N_1283);
nand U4524 (N_4524,N_52,N_984);
nand U4525 (N_4525,N_838,N_145);
or U4526 (N_4526,N_991,N_2117);
nor U4527 (N_4527,N_384,N_1349);
xor U4528 (N_4528,N_2432,N_930);
nor U4529 (N_4529,N_1331,N_1364);
xnor U4530 (N_4530,N_2313,N_1390);
nand U4531 (N_4531,N_359,N_574);
or U4532 (N_4532,N_105,N_956);
and U4533 (N_4533,N_892,N_718);
xor U4534 (N_4534,N_258,N_929);
nor U4535 (N_4535,N_242,N_1039);
xor U4536 (N_4536,N_1694,N_643);
or U4537 (N_4537,N_1932,N_1309);
xor U4538 (N_4538,N_559,N_1558);
and U4539 (N_4539,N_908,N_1300);
nor U4540 (N_4540,N_622,N_698);
nor U4541 (N_4541,N_1325,N_416);
nand U4542 (N_4542,N_2,N_1115);
nand U4543 (N_4543,N_1195,N_969);
xnor U4544 (N_4544,N_1405,N_2206);
and U4545 (N_4545,N_2240,N_232);
and U4546 (N_4546,N_1485,N_538);
or U4547 (N_4547,N_713,N_1810);
nand U4548 (N_4548,N_1819,N_1259);
and U4549 (N_4549,N_1745,N_490);
nand U4550 (N_4550,N_1822,N_2248);
or U4551 (N_4551,N_113,N_1487);
xor U4552 (N_4552,N_648,N_1813);
nor U4553 (N_4553,N_1308,N_2302);
nand U4554 (N_4554,N_1236,N_850);
nor U4555 (N_4555,N_1549,N_1912);
or U4556 (N_4556,N_2421,N_1164);
and U4557 (N_4557,N_206,N_1317);
nor U4558 (N_4558,N_354,N_359);
or U4559 (N_4559,N_1491,N_2159);
and U4560 (N_4560,N_1862,N_1440);
or U4561 (N_4561,N_116,N_70);
nand U4562 (N_4562,N_1114,N_1022);
nand U4563 (N_4563,N_200,N_1382);
and U4564 (N_4564,N_1896,N_2178);
or U4565 (N_4565,N_1108,N_1022);
nor U4566 (N_4566,N_2123,N_2408);
or U4567 (N_4567,N_2017,N_1739);
or U4568 (N_4568,N_1425,N_974);
and U4569 (N_4569,N_2111,N_1205);
or U4570 (N_4570,N_803,N_2075);
and U4571 (N_4571,N_359,N_364);
nand U4572 (N_4572,N_869,N_2459);
and U4573 (N_4573,N_2167,N_606);
and U4574 (N_4574,N_1656,N_788);
nand U4575 (N_4575,N_1991,N_2343);
or U4576 (N_4576,N_636,N_2415);
and U4577 (N_4577,N_335,N_2433);
or U4578 (N_4578,N_2191,N_198);
nand U4579 (N_4579,N_1404,N_1801);
nand U4580 (N_4580,N_900,N_2012);
nand U4581 (N_4581,N_1289,N_247);
xor U4582 (N_4582,N_1485,N_402);
xor U4583 (N_4583,N_1143,N_613);
or U4584 (N_4584,N_2262,N_1881);
nand U4585 (N_4585,N_869,N_2453);
and U4586 (N_4586,N_1309,N_1706);
nor U4587 (N_4587,N_455,N_684);
xor U4588 (N_4588,N_450,N_2359);
and U4589 (N_4589,N_330,N_862);
xor U4590 (N_4590,N_1323,N_1972);
nor U4591 (N_4591,N_2473,N_1879);
or U4592 (N_4592,N_2251,N_823);
or U4593 (N_4593,N_1750,N_2264);
xnor U4594 (N_4594,N_2254,N_635);
nor U4595 (N_4595,N_1499,N_862);
or U4596 (N_4596,N_11,N_745);
nor U4597 (N_4597,N_2413,N_79);
nor U4598 (N_4598,N_610,N_1225);
nor U4599 (N_4599,N_2114,N_423);
and U4600 (N_4600,N_127,N_1185);
nor U4601 (N_4601,N_2369,N_598);
nor U4602 (N_4602,N_1751,N_2052);
and U4603 (N_4603,N_2028,N_644);
and U4604 (N_4604,N_224,N_1097);
and U4605 (N_4605,N_1192,N_1643);
nand U4606 (N_4606,N_1857,N_2266);
nand U4607 (N_4607,N_1897,N_739);
nand U4608 (N_4608,N_1591,N_2377);
xnor U4609 (N_4609,N_995,N_2439);
and U4610 (N_4610,N_457,N_1440);
and U4611 (N_4611,N_2300,N_356);
nand U4612 (N_4612,N_929,N_2213);
or U4613 (N_4613,N_2060,N_2116);
or U4614 (N_4614,N_2052,N_1211);
xnor U4615 (N_4615,N_1013,N_1762);
nor U4616 (N_4616,N_2307,N_1629);
nand U4617 (N_4617,N_587,N_2054);
nand U4618 (N_4618,N_1624,N_855);
nor U4619 (N_4619,N_1167,N_573);
or U4620 (N_4620,N_1517,N_2398);
nor U4621 (N_4621,N_2122,N_1699);
or U4622 (N_4622,N_1990,N_591);
nand U4623 (N_4623,N_2232,N_481);
xor U4624 (N_4624,N_1195,N_42);
xor U4625 (N_4625,N_2193,N_711);
and U4626 (N_4626,N_2462,N_1009);
xor U4627 (N_4627,N_2316,N_976);
nand U4628 (N_4628,N_619,N_2379);
or U4629 (N_4629,N_1978,N_1902);
or U4630 (N_4630,N_1139,N_701);
or U4631 (N_4631,N_1796,N_2084);
nor U4632 (N_4632,N_1087,N_56);
xnor U4633 (N_4633,N_1276,N_552);
nor U4634 (N_4634,N_769,N_19);
or U4635 (N_4635,N_2320,N_1320);
or U4636 (N_4636,N_2336,N_1103);
nor U4637 (N_4637,N_1010,N_2097);
or U4638 (N_4638,N_368,N_1090);
nor U4639 (N_4639,N_219,N_1458);
or U4640 (N_4640,N_532,N_486);
nor U4641 (N_4641,N_2417,N_714);
or U4642 (N_4642,N_1427,N_1227);
nand U4643 (N_4643,N_651,N_2321);
nand U4644 (N_4644,N_156,N_408);
or U4645 (N_4645,N_2017,N_2421);
xor U4646 (N_4646,N_1829,N_123);
and U4647 (N_4647,N_1874,N_1022);
and U4648 (N_4648,N_1851,N_503);
nor U4649 (N_4649,N_345,N_1916);
or U4650 (N_4650,N_2203,N_1699);
nor U4651 (N_4651,N_2319,N_2436);
nor U4652 (N_4652,N_2220,N_487);
and U4653 (N_4653,N_391,N_2080);
nor U4654 (N_4654,N_2498,N_172);
nor U4655 (N_4655,N_1027,N_2043);
nor U4656 (N_4656,N_2096,N_1327);
xor U4657 (N_4657,N_1216,N_256);
nor U4658 (N_4658,N_1210,N_1389);
or U4659 (N_4659,N_1473,N_587);
xnor U4660 (N_4660,N_2441,N_2279);
and U4661 (N_4661,N_250,N_602);
and U4662 (N_4662,N_132,N_1025);
and U4663 (N_4663,N_1696,N_932);
nand U4664 (N_4664,N_1073,N_201);
and U4665 (N_4665,N_2001,N_2035);
or U4666 (N_4666,N_308,N_1781);
and U4667 (N_4667,N_144,N_888);
and U4668 (N_4668,N_2322,N_350);
nand U4669 (N_4669,N_878,N_2062);
or U4670 (N_4670,N_1050,N_1829);
nor U4671 (N_4671,N_2126,N_2339);
xnor U4672 (N_4672,N_1254,N_1895);
and U4673 (N_4673,N_2454,N_55);
or U4674 (N_4674,N_119,N_1622);
nand U4675 (N_4675,N_1981,N_1236);
and U4676 (N_4676,N_1876,N_1202);
xnor U4677 (N_4677,N_376,N_1865);
xnor U4678 (N_4678,N_2206,N_1154);
xor U4679 (N_4679,N_1033,N_1352);
nor U4680 (N_4680,N_1973,N_128);
or U4681 (N_4681,N_872,N_74);
or U4682 (N_4682,N_2183,N_1713);
and U4683 (N_4683,N_1372,N_1963);
xor U4684 (N_4684,N_578,N_1823);
and U4685 (N_4685,N_79,N_1280);
and U4686 (N_4686,N_841,N_2336);
xor U4687 (N_4687,N_1656,N_853);
or U4688 (N_4688,N_2148,N_2023);
xnor U4689 (N_4689,N_242,N_421);
nor U4690 (N_4690,N_2254,N_219);
nor U4691 (N_4691,N_2416,N_766);
and U4692 (N_4692,N_404,N_371);
nand U4693 (N_4693,N_30,N_1036);
nor U4694 (N_4694,N_133,N_2396);
nor U4695 (N_4695,N_1018,N_2351);
xnor U4696 (N_4696,N_679,N_62);
nand U4697 (N_4697,N_715,N_1430);
nand U4698 (N_4698,N_259,N_2180);
nor U4699 (N_4699,N_351,N_384);
nor U4700 (N_4700,N_1691,N_196);
or U4701 (N_4701,N_128,N_2181);
nand U4702 (N_4702,N_661,N_1601);
nand U4703 (N_4703,N_13,N_202);
or U4704 (N_4704,N_1114,N_680);
xor U4705 (N_4705,N_2037,N_1102);
or U4706 (N_4706,N_1887,N_420);
nor U4707 (N_4707,N_1546,N_174);
or U4708 (N_4708,N_711,N_1411);
or U4709 (N_4709,N_378,N_1446);
xor U4710 (N_4710,N_711,N_2122);
xor U4711 (N_4711,N_628,N_2301);
nand U4712 (N_4712,N_1795,N_876);
and U4713 (N_4713,N_1017,N_1622);
or U4714 (N_4714,N_1825,N_214);
nand U4715 (N_4715,N_599,N_2226);
xor U4716 (N_4716,N_2420,N_606);
and U4717 (N_4717,N_1128,N_1818);
nand U4718 (N_4718,N_1620,N_216);
or U4719 (N_4719,N_1182,N_1391);
xnor U4720 (N_4720,N_283,N_376);
nor U4721 (N_4721,N_1302,N_370);
and U4722 (N_4722,N_2115,N_1078);
or U4723 (N_4723,N_220,N_2144);
nor U4724 (N_4724,N_429,N_305);
nor U4725 (N_4725,N_1857,N_2445);
xor U4726 (N_4726,N_1659,N_981);
nor U4727 (N_4727,N_2325,N_602);
or U4728 (N_4728,N_1853,N_1238);
nand U4729 (N_4729,N_156,N_2047);
xor U4730 (N_4730,N_343,N_1167);
nand U4731 (N_4731,N_104,N_1473);
and U4732 (N_4732,N_2032,N_2392);
or U4733 (N_4733,N_1192,N_1936);
xor U4734 (N_4734,N_2379,N_1122);
nor U4735 (N_4735,N_158,N_1275);
nor U4736 (N_4736,N_1729,N_1025);
or U4737 (N_4737,N_577,N_1857);
xor U4738 (N_4738,N_225,N_2489);
and U4739 (N_4739,N_2102,N_890);
and U4740 (N_4740,N_954,N_1662);
nand U4741 (N_4741,N_2440,N_1185);
or U4742 (N_4742,N_61,N_1558);
xnor U4743 (N_4743,N_2442,N_1);
xor U4744 (N_4744,N_204,N_1776);
or U4745 (N_4745,N_2327,N_2379);
nand U4746 (N_4746,N_1720,N_496);
or U4747 (N_4747,N_144,N_67);
or U4748 (N_4748,N_117,N_809);
nor U4749 (N_4749,N_1472,N_1129);
or U4750 (N_4750,N_1880,N_1743);
xnor U4751 (N_4751,N_156,N_1678);
or U4752 (N_4752,N_198,N_1643);
and U4753 (N_4753,N_567,N_573);
xnor U4754 (N_4754,N_1427,N_813);
xor U4755 (N_4755,N_75,N_559);
and U4756 (N_4756,N_2167,N_832);
and U4757 (N_4757,N_1617,N_2326);
nor U4758 (N_4758,N_259,N_1959);
xnor U4759 (N_4759,N_164,N_281);
xor U4760 (N_4760,N_489,N_2265);
and U4761 (N_4761,N_842,N_273);
xor U4762 (N_4762,N_721,N_2165);
or U4763 (N_4763,N_2240,N_1490);
and U4764 (N_4764,N_218,N_1904);
nor U4765 (N_4765,N_161,N_285);
or U4766 (N_4766,N_1453,N_470);
and U4767 (N_4767,N_467,N_967);
and U4768 (N_4768,N_1613,N_2293);
or U4769 (N_4769,N_309,N_197);
nand U4770 (N_4770,N_44,N_187);
and U4771 (N_4771,N_2352,N_2361);
nor U4772 (N_4772,N_2044,N_1133);
nand U4773 (N_4773,N_1385,N_954);
or U4774 (N_4774,N_1346,N_2466);
xor U4775 (N_4775,N_1572,N_789);
nor U4776 (N_4776,N_1822,N_33);
or U4777 (N_4777,N_2460,N_1222);
and U4778 (N_4778,N_102,N_640);
or U4779 (N_4779,N_187,N_37);
nand U4780 (N_4780,N_1535,N_441);
xnor U4781 (N_4781,N_2438,N_1224);
nor U4782 (N_4782,N_587,N_1308);
and U4783 (N_4783,N_67,N_507);
and U4784 (N_4784,N_551,N_1832);
nand U4785 (N_4785,N_2328,N_1722);
or U4786 (N_4786,N_1017,N_2158);
or U4787 (N_4787,N_415,N_741);
and U4788 (N_4788,N_378,N_458);
nor U4789 (N_4789,N_1524,N_2488);
xnor U4790 (N_4790,N_1400,N_2440);
or U4791 (N_4791,N_1738,N_1065);
xor U4792 (N_4792,N_2489,N_321);
nand U4793 (N_4793,N_1820,N_71);
nand U4794 (N_4794,N_1117,N_512);
xnor U4795 (N_4795,N_1696,N_2296);
nor U4796 (N_4796,N_580,N_2061);
and U4797 (N_4797,N_866,N_1567);
and U4798 (N_4798,N_1896,N_2016);
nor U4799 (N_4799,N_595,N_179);
nand U4800 (N_4800,N_140,N_186);
or U4801 (N_4801,N_672,N_702);
nand U4802 (N_4802,N_391,N_1592);
nor U4803 (N_4803,N_1761,N_1025);
xor U4804 (N_4804,N_1357,N_877);
xor U4805 (N_4805,N_2479,N_1185);
and U4806 (N_4806,N_137,N_1813);
nand U4807 (N_4807,N_2191,N_2391);
nand U4808 (N_4808,N_1316,N_1269);
xor U4809 (N_4809,N_938,N_2406);
nor U4810 (N_4810,N_895,N_1972);
nor U4811 (N_4811,N_586,N_1350);
and U4812 (N_4812,N_90,N_779);
nor U4813 (N_4813,N_569,N_230);
or U4814 (N_4814,N_2362,N_854);
xnor U4815 (N_4815,N_1419,N_2137);
nand U4816 (N_4816,N_1153,N_1928);
nand U4817 (N_4817,N_1669,N_1372);
xnor U4818 (N_4818,N_1629,N_667);
nand U4819 (N_4819,N_2266,N_55);
or U4820 (N_4820,N_730,N_605);
xor U4821 (N_4821,N_1182,N_1299);
and U4822 (N_4822,N_1283,N_2222);
nand U4823 (N_4823,N_2244,N_1188);
nand U4824 (N_4824,N_1344,N_2030);
nor U4825 (N_4825,N_661,N_847);
or U4826 (N_4826,N_1316,N_1344);
xor U4827 (N_4827,N_774,N_2415);
and U4828 (N_4828,N_1253,N_1328);
or U4829 (N_4829,N_661,N_76);
nand U4830 (N_4830,N_1220,N_1785);
nor U4831 (N_4831,N_2375,N_665);
nor U4832 (N_4832,N_1040,N_1125);
or U4833 (N_4833,N_1673,N_409);
and U4834 (N_4834,N_2110,N_671);
nand U4835 (N_4835,N_1728,N_2393);
nor U4836 (N_4836,N_1672,N_1363);
xnor U4837 (N_4837,N_1723,N_1135);
or U4838 (N_4838,N_7,N_448);
nand U4839 (N_4839,N_366,N_72);
or U4840 (N_4840,N_804,N_216);
and U4841 (N_4841,N_1581,N_1140);
nand U4842 (N_4842,N_731,N_2334);
xnor U4843 (N_4843,N_315,N_434);
or U4844 (N_4844,N_1809,N_912);
or U4845 (N_4845,N_846,N_244);
and U4846 (N_4846,N_1660,N_1743);
nand U4847 (N_4847,N_265,N_2231);
nor U4848 (N_4848,N_2239,N_1734);
nor U4849 (N_4849,N_810,N_1308);
nor U4850 (N_4850,N_1863,N_1406);
nand U4851 (N_4851,N_1337,N_2025);
and U4852 (N_4852,N_948,N_1090);
or U4853 (N_4853,N_259,N_2453);
nor U4854 (N_4854,N_1093,N_773);
or U4855 (N_4855,N_1481,N_2324);
xor U4856 (N_4856,N_1256,N_1869);
or U4857 (N_4857,N_1396,N_1152);
nor U4858 (N_4858,N_2417,N_2155);
xnor U4859 (N_4859,N_858,N_2473);
and U4860 (N_4860,N_1903,N_167);
xnor U4861 (N_4861,N_145,N_1614);
nor U4862 (N_4862,N_1133,N_699);
xnor U4863 (N_4863,N_331,N_570);
xnor U4864 (N_4864,N_1310,N_1002);
nor U4865 (N_4865,N_569,N_421);
and U4866 (N_4866,N_970,N_162);
nand U4867 (N_4867,N_1877,N_2324);
nor U4868 (N_4868,N_1289,N_2466);
nand U4869 (N_4869,N_1616,N_1533);
nor U4870 (N_4870,N_1582,N_1933);
or U4871 (N_4871,N_95,N_1787);
and U4872 (N_4872,N_880,N_2336);
nand U4873 (N_4873,N_285,N_2343);
or U4874 (N_4874,N_355,N_1591);
and U4875 (N_4875,N_2392,N_1859);
nor U4876 (N_4876,N_151,N_1138);
nand U4877 (N_4877,N_610,N_1714);
nand U4878 (N_4878,N_2339,N_1498);
xor U4879 (N_4879,N_395,N_1531);
xor U4880 (N_4880,N_116,N_817);
nand U4881 (N_4881,N_483,N_1058);
nor U4882 (N_4882,N_2320,N_1473);
or U4883 (N_4883,N_2440,N_858);
nand U4884 (N_4884,N_1459,N_2224);
or U4885 (N_4885,N_416,N_1828);
and U4886 (N_4886,N_2202,N_1576);
nor U4887 (N_4887,N_94,N_1520);
or U4888 (N_4888,N_374,N_2057);
nand U4889 (N_4889,N_192,N_2195);
or U4890 (N_4890,N_2048,N_2031);
or U4891 (N_4891,N_1317,N_139);
or U4892 (N_4892,N_2095,N_1791);
nor U4893 (N_4893,N_669,N_531);
and U4894 (N_4894,N_1435,N_1315);
or U4895 (N_4895,N_2150,N_354);
nand U4896 (N_4896,N_563,N_2331);
nor U4897 (N_4897,N_1409,N_1299);
nand U4898 (N_4898,N_282,N_1484);
and U4899 (N_4899,N_2141,N_1867);
xor U4900 (N_4900,N_1341,N_132);
nand U4901 (N_4901,N_1728,N_1980);
or U4902 (N_4902,N_797,N_444);
and U4903 (N_4903,N_2284,N_769);
nand U4904 (N_4904,N_2420,N_1298);
nand U4905 (N_4905,N_1186,N_1616);
or U4906 (N_4906,N_1157,N_1758);
nand U4907 (N_4907,N_1868,N_1729);
and U4908 (N_4908,N_578,N_167);
and U4909 (N_4909,N_309,N_2470);
and U4910 (N_4910,N_2361,N_2029);
or U4911 (N_4911,N_1131,N_65);
xnor U4912 (N_4912,N_324,N_1901);
and U4913 (N_4913,N_1333,N_1979);
nand U4914 (N_4914,N_769,N_2038);
or U4915 (N_4915,N_1061,N_684);
nor U4916 (N_4916,N_490,N_42);
xnor U4917 (N_4917,N_1989,N_2463);
xor U4918 (N_4918,N_318,N_1924);
and U4919 (N_4919,N_1289,N_702);
and U4920 (N_4920,N_1312,N_1532);
nor U4921 (N_4921,N_1855,N_1818);
nand U4922 (N_4922,N_1772,N_2250);
and U4923 (N_4923,N_463,N_1101);
nor U4924 (N_4924,N_1095,N_585);
nand U4925 (N_4925,N_700,N_636);
nor U4926 (N_4926,N_1806,N_2278);
or U4927 (N_4927,N_1869,N_929);
and U4928 (N_4928,N_1174,N_2023);
xnor U4929 (N_4929,N_2097,N_770);
or U4930 (N_4930,N_2444,N_781);
and U4931 (N_4931,N_2263,N_475);
nand U4932 (N_4932,N_602,N_320);
xor U4933 (N_4933,N_38,N_1367);
nand U4934 (N_4934,N_206,N_2432);
or U4935 (N_4935,N_1460,N_2255);
xnor U4936 (N_4936,N_2425,N_1781);
and U4937 (N_4937,N_1933,N_541);
nor U4938 (N_4938,N_206,N_2204);
nand U4939 (N_4939,N_73,N_1733);
nand U4940 (N_4940,N_265,N_589);
or U4941 (N_4941,N_2435,N_216);
nor U4942 (N_4942,N_2119,N_1588);
xnor U4943 (N_4943,N_2365,N_1674);
xnor U4944 (N_4944,N_87,N_545);
nand U4945 (N_4945,N_1232,N_1751);
nor U4946 (N_4946,N_2108,N_1736);
xor U4947 (N_4947,N_1517,N_298);
and U4948 (N_4948,N_2363,N_254);
and U4949 (N_4949,N_293,N_1494);
nand U4950 (N_4950,N_220,N_2249);
nor U4951 (N_4951,N_2107,N_631);
nand U4952 (N_4952,N_1663,N_2084);
or U4953 (N_4953,N_2310,N_2156);
and U4954 (N_4954,N_1991,N_1510);
or U4955 (N_4955,N_1906,N_1383);
and U4956 (N_4956,N_849,N_2104);
nand U4957 (N_4957,N_1763,N_2447);
nand U4958 (N_4958,N_1642,N_1081);
xnor U4959 (N_4959,N_206,N_2119);
and U4960 (N_4960,N_1551,N_2146);
and U4961 (N_4961,N_1980,N_2232);
xor U4962 (N_4962,N_2187,N_711);
or U4963 (N_4963,N_244,N_2086);
and U4964 (N_4964,N_1847,N_143);
or U4965 (N_4965,N_1212,N_1867);
and U4966 (N_4966,N_1147,N_2184);
xnor U4967 (N_4967,N_507,N_536);
nor U4968 (N_4968,N_347,N_1125);
and U4969 (N_4969,N_1754,N_1600);
or U4970 (N_4970,N_2173,N_1847);
and U4971 (N_4971,N_1795,N_1182);
xor U4972 (N_4972,N_635,N_362);
or U4973 (N_4973,N_765,N_1107);
or U4974 (N_4974,N_2172,N_1167);
nor U4975 (N_4975,N_2333,N_1665);
or U4976 (N_4976,N_802,N_2223);
nand U4977 (N_4977,N_1712,N_827);
or U4978 (N_4978,N_271,N_2160);
or U4979 (N_4979,N_1547,N_972);
nor U4980 (N_4980,N_2354,N_519);
nor U4981 (N_4981,N_1465,N_174);
and U4982 (N_4982,N_1687,N_1519);
nor U4983 (N_4983,N_754,N_289);
and U4984 (N_4984,N_82,N_1697);
xor U4985 (N_4985,N_983,N_1754);
nand U4986 (N_4986,N_1770,N_1351);
or U4987 (N_4987,N_2137,N_217);
or U4988 (N_4988,N_1729,N_756);
nor U4989 (N_4989,N_2159,N_142);
and U4990 (N_4990,N_1362,N_306);
nand U4991 (N_4991,N_526,N_2268);
nand U4992 (N_4992,N_581,N_2260);
nand U4993 (N_4993,N_1415,N_346);
nor U4994 (N_4994,N_1176,N_1341);
nor U4995 (N_4995,N_1455,N_2271);
nand U4996 (N_4996,N_314,N_1978);
or U4997 (N_4997,N_340,N_627);
nand U4998 (N_4998,N_2180,N_2495);
xnor U4999 (N_4999,N_2203,N_1012);
nand U5000 (N_5000,N_4633,N_3078);
xnor U5001 (N_5001,N_4483,N_3382);
or U5002 (N_5002,N_4681,N_4552);
nand U5003 (N_5003,N_3011,N_3587);
nor U5004 (N_5004,N_3397,N_4987);
or U5005 (N_5005,N_4243,N_3888);
xnor U5006 (N_5006,N_4600,N_2709);
nor U5007 (N_5007,N_3164,N_2855);
nand U5008 (N_5008,N_4773,N_2752);
nor U5009 (N_5009,N_4171,N_4732);
or U5010 (N_5010,N_3714,N_4988);
nor U5011 (N_5011,N_3291,N_3904);
nor U5012 (N_5012,N_3407,N_4686);
xnor U5013 (N_5013,N_4366,N_4185);
and U5014 (N_5014,N_3566,N_4093);
nand U5015 (N_5015,N_3393,N_4113);
and U5016 (N_5016,N_3831,N_3353);
xor U5017 (N_5017,N_3372,N_3383);
nand U5018 (N_5018,N_3176,N_4809);
and U5019 (N_5019,N_4606,N_4588);
xor U5020 (N_5020,N_3613,N_2947);
nor U5021 (N_5021,N_2745,N_3442);
nand U5022 (N_5022,N_2776,N_4638);
nor U5023 (N_5023,N_3694,N_4038);
nor U5024 (N_5024,N_4969,N_3650);
and U5025 (N_5025,N_3314,N_3321);
nand U5026 (N_5026,N_4830,N_3192);
nor U5027 (N_5027,N_3903,N_3057);
xnor U5028 (N_5028,N_3367,N_4709);
nand U5029 (N_5029,N_3546,N_4948);
and U5030 (N_5030,N_4438,N_2889);
and U5031 (N_5031,N_4540,N_4872);
xnor U5032 (N_5032,N_3932,N_2800);
and U5033 (N_5033,N_3626,N_4693);
nor U5034 (N_5034,N_2618,N_3070);
or U5035 (N_5035,N_3081,N_4747);
or U5036 (N_5036,N_3523,N_2827);
nand U5037 (N_5037,N_4912,N_2857);
nor U5038 (N_5038,N_4324,N_4610);
xnor U5039 (N_5039,N_2711,N_4542);
or U5040 (N_5040,N_2999,N_4248);
nand U5041 (N_5041,N_3247,N_4719);
xnor U5042 (N_5042,N_2706,N_4420);
and U5043 (N_5043,N_3118,N_4331);
nor U5044 (N_5044,N_3340,N_3162);
nor U5045 (N_5045,N_3708,N_4429);
xnor U5046 (N_5046,N_4503,N_3717);
nor U5047 (N_5047,N_4471,N_4280);
or U5048 (N_5048,N_4323,N_4843);
and U5049 (N_5049,N_4805,N_2829);
nand U5050 (N_5050,N_4617,N_4364);
and U5051 (N_5051,N_3837,N_3283);
nand U5052 (N_5052,N_4590,N_3661);
and U5053 (N_5053,N_2750,N_2818);
or U5054 (N_5054,N_4487,N_2665);
nor U5055 (N_5055,N_3489,N_4906);
and U5056 (N_5056,N_3352,N_3312);
xor U5057 (N_5057,N_3834,N_4742);
and U5058 (N_5058,N_4309,N_2995);
nor U5059 (N_5059,N_4739,N_2982);
and U5060 (N_5060,N_3278,N_3400);
and U5061 (N_5061,N_4463,N_3119);
nor U5062 (N_5062,N_4522,N_4581);
nor U5063 (N_5063,N_3189,N_3555);
nor U5064 (N_5064,N_2799,N_2977);
or U5065 (N_5065,N_3728,N_3270);
or U5066 (N_5066,N_2795,N_2727);
and U5067 (N_5067,N_3971,N_3540);
or U5068 (N_5068,N_2737,N_2527);
nor U5069 (N_5069,N_4683,N_2761);
nor U5070 (N_5070,N_2983,N_3193);
and U5071 (N_5071,N_4338,N_3521);
xor U5072 (N_5072,N_2622,N_4138);
nand U5073 (N_5073,N_3204,N_3020);
nand U5074 (N_5074,N_4075,N_4343);
nor U5075 (N_5075,N_4791,N_3260);
nor U5076 (N_5076,N_4180,N_4135);
and U5077 (N_5077,N_4209,N_2524);
or U5078 (N_5078,N_3537,N_4382);
xor U5079 (N_5079,N_3207,N_3706);
nor U5080 (N_5080,N_4435,N_4431);
and U5081 (N_5081,N_2601,N_4557);
nor U5082 (N_5082,N_3474,N_4777);
nand U5083 (N_5083,N_3990,N_4716);
nor U5084 (N_5084,N_4611,N_4721);
nand U5085 (N_5085,N_3104,N_3210);
or U5086 (N_5086,N_2949,N_4114);
xnor U5087 (N_5087,N_3785,N_4145);
or U5088 (N_5088,N_2671,N_3544);
nor U5089 (N_5089,N_2648,N_4266);
xor U5090 (N_5090,N_4751,N_3362);
or U5091 (N_5091,N_4104,N_2748);
or U5092 (N_5092,N_4211,N_4886);
xor U5093 (N_5093,N_2842,N_2511);
nand U5094 (N_5094,N_2550,N_4986);
nand U5095 (N_5095,N_4879,N_3775);
nand U5096 (N_5096,N_2990,N_4735);
and U5097 (N_5097,N_3951,N_4692);
or U5098 (N_5098,N_4359,N_3236);
nand U5099 (N_5099,N_4291,N_3478);
nor U5100 (N_5100,N_4713,N_2871);
and U5101 (N_5101,N_4937,N_4608);
and U5102 (N_5102,N_4785,N_4949);
nand U5103 (N_5103,N_4636,N_4406);
xor U5104 (N_5104,N_4015,N_3360);
nor U5105 (N_5105,N_3701,N_3106);
nand U5106 (N_5106,N_3859,N_4007);
xnor U5107 (N_5107,N_4149,N_4860);
or U5108 (N_5108,N_4458,N_3581);
xnor U5109 (N_5109,N_4449,N_3058);
nor U5110 (N_5110,N_2803,N_4575);
or U5111 (N_5111,N_2839,N_4302);
or U5112 (N_5112,N_4694,N_4155);
nor U5113 (N_5113,N_2720,N_3033);
or U5114 (N_5114,N_3909,N_4946);
and U5115 (N_5115,N_3941,N_4231);
nand U5116 (N_5116,N_4861,N_3818);
and U5117 (N_5117,N_3102,N_4369);
nand U5118 (N_5118,N_2812,N_3813);
nand U5119 (N_5119,N_4717,N_2814);
and U5120 (N_5120,N_3525,N_3497);
xnor U5121 (N_5121,N_2951,N_4904);
or U5122 (N_5122,N_4288,N_3042);
nor U5123 (N_5123,N_2735,N_4237);
and U5124 (N_5124,N_4762,N_3456);
and U5125 (N_5125,N_3799,N_3730);
and U5126 (N_5126,N_3562,N_2661);
nor U5127 (N_5127,N_2876,N_4898);
nor U5128 (N_5128,N_3361,N_2603);
and U5129 (N_5129,N_2915,N_2656);
or U5130 (N_5130,N_2673,N_2683);
or U5131 (N_5131,N_3606,N_3590);
xnor U5132 (N_5132,N_4178,N_3366);
nand U5133 (N_5133,N_3745,N_4482);
nand U5134 (N_5134,N_4193,N_2798);
or U5135 (N_5135,N_2877,N_2846);
xnor U5136 (N_5136,N_3296,N_3095);
nor U5137 (N_5137,N_4790,N_4476);
and U5138 (N_5138,N_4472,N_3844);
nand U5139 (N_5139,N_4400,N_4335);
xnor U5140 (N_5140,N_4797,N_4485);
nor U5141 (N_5141,N_2591,N_3695);
and U5142 (N_5142,N_2721,N_4412);
and U5143 (N_5143,N_4853,N_3823);
and U5144 (N_5144,N_2614,N_4350);
nand U5145 (N_5145,N_3824,N_3451);
nor U5146 (N_5146,N_2731,N_4268);
nor U5147 (N_5147,N_3527,N_3486);
nor U5148 (N_5148,N_3053,N_3879);
and U5149 (N_5149,N_2697,N_4940);
or U5150 (N_5150,N_4258,N_4652);
or U5151 (N_5151,N_3698,N_2584);
or U5152 (N_5152,N_3069,N_3174);
and U5153 (N_5153,N_3392,N_4955);
and U5154 (N_5154,N_3638,N_3809);
xor U5155 (N_5155,N_2617,N_2912);
or U5156 (N_5156,N_4976,N_4062);
and U5157 (N_5157,N_4405,N_2736);
xor U5158 (N_5158,N_4441,N_4033);
nand U5159 (N_5159,N_4819,N_3461);
and U5160 (N_5160,N_4547,N_4784);
nand U5161 (N_5161,N_4439,N_3940);
xnor U5162 (N_5162,N_4461,N_4598);
nand U5163 (N_5163,N_4232,N_3465);
and U5164 (N_5164,N_4004,N_2627);
and U5165 (N_5165,N_2950,N_2961);
xnor U5166 (N_5166,N_4068,N_4097);
nand U5167 (N_5167,N_4817,N_4945);
and U5168 (N_5168,N_2934,N_3394);
and U5169 (N_5169,N_2922,N_2694);
nand U5170 (N_5170,N_3226,N_3403);
xnor U5171 (N_5171,N_3284,N_3761);
or U5172 (N_5172,N_3666,N_2675);
or U5173 (N_5173,N_3711,N_2941);
xor U5174 (N_5174,N_3607,N_3950);
xnor U5175 (N_5175,N_3750,N_4105);
nand U5176 (N_5176,N_3239,N_3111);
and U5177 (N_5177,N_4665,N_4251);
xor U5178 (N_5178,N_4909,N_4753);
and U5179 (N_5179,N_2868,N_2732);
nand U5180 (N_5180,N_4000,N_4714);
and U5181 (N_5181,N_2900,N_3578);
and U5182 (N_5182,N_3025,N_2521);
or U5183 (N_5183,N_3303,N_3026);
nand U5184 (N_5184,N_4034,N_4357);
and U5185 (N_5185,N_4964,N_4725);
nor U5186 (N_5186,N_3219,N_4842);
nand U5187 (N_5187,N_3059,N_3691);
or U5188 (N_5188,N_2780,N_4261);
nand U5189 (N_5189,N_4179,N_4867);
nand U5190 (N_5190,N_2640,N_4219);
xnor U5191 (N_5191,N_2851,N_4066);
and U5192 (N_5192,N_3787,N_4915);
xnor U5193 (N_5193,N_4025,N_4152);
xnor U5194 (N_5194,N_4883,N_2817);
or U5195 (N_5195,N_3519,N_3633);
or U5196 (N_5196,N_3333,N_2597);
nand U5197 (N_5197,N_4101,N_2699);
xnor U5198 (N_5198,N_4602,N_3071);
or U5199 (N_5199,N_4531,N_4414);
nand U5200 (N_5200,N_2880,N_3052);
nor U5201 (N_5201,N_3722,N_3100);
or U5202 (N_5202,N_3565,N_4440);
xor U5203 (N_5203,N_2526,N_2952);
and U5204 (N_5204,N_4174,N_3122);
or U5205 (N_5205,N_3402,N_3178);
xor U5206 (N_5206,N_3826,N_2739);
and U5207 (N_5207,N_4279,N_4409);
nor U5208 (N_5208,N_3543,N_3846);
or U5209 (N_5209,N_2960,N_2548);
xnor U5210 (N_5210,N_2894,N_2634);
xor U5211 (N_5211,N_2978,N_3601);
xor U5212 (N_5212,N_4035,N_4908);
xnor U5213 (N_5213,N_4927,N_4119);
xor U5214 (N_5214,N_2596,N_3384);
and U5215 (N_5215,N_2593,N_3757);
nand U5216 (N_5216,N_4727,N_4653);
nor U5217 (N_5217,N_3028,N_3965);
nor U5218 (N_5218,N_3452,N_4162);
or U5219 (N_5219,N_3037,N_2542);
nor U5220 (N_5220,N_2652,N_2967);
and U5221 (N_5221,N_4183,N_2859);
nor U5222 (N_5222,N_3449,N_4120);
or U5223 (N_5223,N_2805,N_3356);
or U5224 (N_5224,N_3657,N_3986);
xor U5225 (N_5225,N_3013,N_3096);
nor U5226 (N_5226,N_3789,N_4844);
or U5227 (N_5227,N_3079,N_3018);
xor U5228 (N_5228,N_3238,N_2605);
and U5229 (N_5229,N_4783,N_2775);
and U5230 (N_5230,N_4954,N_2802);
xor U5231 (N_5231,N_4074,N_3862);
or U5232 (N_5232,N_2623,N_2756);
nor U5233 (N_5233,N_3195,N_4477);
or U5234 (N_5234,N_4534,N_2559);
or U5235 (N_5235,N_4130,N_3265);
nand U5236 (N_5236,N_3840,N_4859);
or U5237 (N_5237,N_3737,N_4204);
and U5238 (N_5238,N_3589,N_3499);
nand U5239 (N_5239,N_4579,N_4161);
nand U5240 (N_5240,N_3330,N_2964);
xor U5241 (N_5241,N_4466,N_3476);
xnor U5242 (N_5242,N_2535,N_3365);
nor U5243 (N_5243,N_4082,N_4868);
xnor U5244 (N_5244,N_2534,N_3970);
nor U5245 (N_5245,N_3632,N_3983);
or U5246 (N_5246,N_3213,N_2808);
nand U5247 (N_5247,N_4985,N_3343);
nor U5248 (N_5248,N_4148,N_4698);
xnor U5249 (N_5249,N_4275,N_3148);
xnor U5250 (N_5250,N_2822,N_3389);
nor U5251 (N_5251,N_3437,N_4071);
nand U5252 (N_5252,N_2718,N_2836);
or U5253 (N_5253,N_4666,N_4895);
or U5254 (N_5254,N_4601,N_4604);
xor U5255 (N_5255,N_4787,N_2589);
or U5256 (N_5256,N_4222,N_3894);
and U5257 (N_5257,N_4271,N_4580);
nor U5258 (N_5258,N_2670,N_4123);
or U5259 (N_5259,N_4761,N_2549);
nor U5260 (N_5260,N_3067,N_3976);
and U5261 (N_5261,N_4277,N_3997);
nand U5262 (N_5262,N_4930,N_4630);
nor U5263 (N_5263,N_2519,N_3268);
or U5264 (N_5264,N_4939,N_4848);
nor U5265 (N_5265,N_4432,N_4234);
nand U5266 (N_5266,N_4917,N_4831);
xor U5267 (N_5267,N_4298,N_3252);
xor U5268 (N_5268,N_3446,N_2804);
nand U5269 (N_5269,N_3072,N_4107);
nand U5270 (N_5270,N_3036,N_3861);
xor U5271 (N_5271,N_3736,N_3504);
and U5272 (N_5272,N_2588,N_3954);
nor U5273 (N_5273,N_3723,N_3006);
and U5274 (N_5274,N_3082,N_4584);
and U5275 (N_5275,N_3492,N_2541);
nand U5276 (N_5276,N_3700,N_3586);
xnor U5277 (N_5277,N_4555,N_4168);
xor U5278 (N_5278,N_4620,N_4320);
nand U5279 (N_5279,N_4850,N_2753);
nand U5280 (N_5280,N_4064,N_4896);
nand U5281 (N_5281,N_3858,N_2561);
and U5282 (N_5282,N_3772,N_3426);
xnor U5283 (N_5283,N_3713,N_3864);
or U5284 (N_5284,N_3167,N_4589);
and U5285 (N_5285,N_4933,N_2663);
and U5286 (N_5286,N_4746,N_3132);
or U5287 (N_5287,N_3784,N_3803);
and U5288 (N_5288,N_3323,N_4292);
xor U5289 (N_5289,N_4743,N_2908);
or U5290 (N_5290,N_4392,N_3960);
or U5291 (N_5291,N_2708,N_4203);
nor U5292 (N_5292,N_3438,N_2907);
nand U5293 (N_5293,N_4259,N_4257);
nand U5294 (N_5294,N_4173,N_2807);
xor U5295 (N_5295,N_4659,N_4926);
nand U5296 (N_5296,N_3625,N_4253);
nor U5297 (N_5297,N_2998,N_4923);
nor U5298 (N_5298,N_4778,N_2508);
nand U5299 (N_5299,N_3806,N_2937);
or U5300 (N_5300,N_4265,N_3375);
nand U5301 (N_5301,N_4703,N_3275);
and U5302 (N_5302,N_4866,N_3161);
nand U5303 (N_5303,N_3910,N_3863);
and U5304 (N_5304,N_4142,N_2556);
xor U5305 (N_5305,N_3931,N_2646);
nand U5306 (N_5306,N_3399,N_4958);
xor U5307 (N_5307,N_2782,N_4078);
and U5308 (N_5308,N_3202,N_2959);
and U5309 (N_5309,N_4565,N_3667);
nor U5310 (N_5310,N_3038,N_3410);
xor U5311 (N_5311,N_4942,N_2560);
nor U5312 (N_5312,N_3988,N_4088);
or U5313 (N_5313,N_4479,N_4526);
and U5314 (N_5314,N_4413,N_4996);
and U5315 (N_5315,N_3927,N_3001);
and U5316 (N_5316,N_3536,N_4497);
nand U5317 (N_5317,N_3506,N_4799);
nor U5318 (N_5318,N_4974,N_4404);
xnor U5319 (N_5319,N_3501,N_4658);
or U5320 (N_5320,N_3724,N_3891);
and U5321 (N_5321,N_3748,N_3311);
or U5322 (N_5322,N_2783,N_3792);
xor U5323 (N_5323,N_3947,N_4934);
nor U5324 (N_5324,N_3849,N_2791);
or U5325 (N_5325,N_4318,N_4544);
xor U5326 (N_5326,N_4260,N_4558);
or U5327 (N_5327,N_3630,N_3307);
nand U5328 (N_5328,N_4944,N_3703);
and U5329 (N_5329,N_4533,N_3777);
and U5330 (N_5330,N_4635,N_2766);
xor U5331 (N_5331,N_4614,N_3182);
or U5332 (N_5332,N_3429,N_3767);
nand U5333 (N_5333,N_3884,N_3290);
xnor U5334 (N_5334,N_4530,N_3170);
xnor U5335 (N_5335,N_3257,N_3117);
or U5336 (N_5336,N_3583,N_2760);
nand U5337 (N_5337,N_4273,N_4982);
or U5338 (N_5338,N_3845,N_4637);
xnor U5339 (N_5339,N_2975,N_2628);
xor U5340 (N_5340,N_3160,N_4643);
or U5341 (N_5341,N_4046,N_3682);
and U5342 (N_5342,N_3422,N_4158);
nor U5343 (N_5343,N_4084,N_4192);
and U5344 (N_5344,N_2893,N_3793);
nand U5345 (N_5345,N_3526,N_3301);
nor U5346 (N_5346,N_4206,N_3743);
nand U5347 (N_5347,N_4083,N_3600);
nor U5348 (N_5348,N_3250,N_3670);
nor U5349 (N_5349,N_3575,N_3808);
and U5350 (N_5350,N_4668,N_3658);
xnor U5351 (N_5351,N_3224,N_4052);
nor U5352 (N_5352,N_2738,N_4786);
nand U5353 (N_5353,N_3348,N_4815);
xor U5354 (N_5354,N_2897,N_4577);
nor U5355 (N_5355,N_4514,N_4621);
xnor U5356 (N_5356,N_3008,N_3842);
and U5357 (N_5357,N_3277,N_2693);
and U5358 (N_5358,N_3327,N_4215);
nand U5359 (N_5359,N_3075,N_3967);
xor U5360 (N_5360,N_3535,N_3851);
or U5361 (N_5361,N_3163,N_3496);
xnor U5362 (N_5362,N_2759,N_4972);
nand U5363 (N_5363,N_3386,N_3066);
or U5364 (N_5364,N_4319,N_3105);
and U5365 (N_5365,N_3573,N_2910);
and U5366 (N_5366,N_2828,N_3593);
and U5367 (N_5367,N_3783,N_3493);
nand U5368 (N_5368,N_3597,N_4294);
nor U5369 (N_5369,N_3147,N_3232);
nand U5370 (N_5370,N_3261,N_4663);
and U5371 (N_5371,N_4792,N_4656);
or U5372 (N_5372,N_2644,N_2532);
or U5373 (N_5373,N_3009,N_3716);
and U5374 (N_5374,N_4607,N_3896);
nor U5375 (N_5375,N_2779,N_2996);
or U5376 (N_5376,N_4593,N_4447);
or U5377 (N_5377,N_3672,N_3430);
xnor U5378 (N_5378,N_2764,N_3871);
nor U5379 (N_5379,N_4498,N_2568);
xor U5380 (N_5380,N_4150,N_4037);
and U5381 (N_5381,N_4838,N_3952);
or U5382 (N_5382,N_3991,N_3557);
nand U5383 (N_5383,N_3503,N_3801);
xor U5384 (N_5384,N_2672,N_3612);
xor U5385 (N_5385,N_2987,N_3217);
or U5386 (N_5386,N_4303,N_3432);
and U5387 (N_5387,N_4704,N_3076);
xor U5388 (N_5388,N_3387,N_3516);
and U5389 (N_5389,N_3322,N_2856);
or U5390 (N_5390,N_4510,N_4421);
nand U5391 (N_5391,N_4640,N_3300);
and U5392 (N_5392,N_2754,N_2666);
and U5393 (N_5393,N_2520,N_2724);
nor U5394 (N_5394,N_4067,N_4774);
or U5395 (N_5395,N_4375,N_3917);
xnor U5396 (N_5396,N_4176,N_4385);
nand U5397 (N_5397,N_3194,N_4801);
xnor U5398 (N_5398,N_3796,N_4172);
nand U5399 (N_5399,N_4613,N_3928);
and U5400 (N_5400,N_2680,N_4213);
nor U5401 (N_5401,N_4631,N_4040);
xor U5402 (N_5402,N_3628,N_3732);
xnor U5403 (N_5403,N_4766,N_3098);
xnor U5404 (N_5404,N_3689,N_3596);
or U5405 (N_5405,N_3398,N_3532);
and U5406 (N_5406,N_2890,N_3620);
nor U5407 (N_5407,N_3335,N_3766);
and U5408 (N_5408,N_4833,N_3520);
and U5409 (N_5409,N_4221,N_3240);
and U5410 (N_5410,N_2801,N_4768);
and U5411 (N_5411,N_4239,N_2792);
and U5412 (N_5412,N_3010,N_4316);
nor U5413 (N_5413,N_4835,N_3996);
nand U5414 (N_5414,N_3051,N_4326);
xnor U5415 (N_5415,N_4009,N_2566);
nor U5416 (N_5416,N_3355,N_2531);
nor U5417 (N_5417,N_4169,N_4134);
or U5418 (N_5418,N_4803,N_4595);
nand U5419 (N_5419,N_4187,N_3481);
nor U5420 (N_5420,N_3688,N_3999);
xor U5421 (N_5421,N_3417,N_2957);
xor U5422 (N_5422,N_3376,N_2899);
and U5423 (N_5423,N_3614,N_3897);
and U5424 (N_5424,N_3924,N_4468);
xor U5425 (N_5425,N_2544,N_4442);
nand U5426 (N_5426,N_3550,N_3734);
nand U5427 (N_5427,N_3822,N_4451);
or U5428 (N_5428,N_2674,N_2863);
or U5429 (N_5429,N_4810,N_3077);
and U5430 (N_5430,N_4676,N_2744);
nand U5431 (N_5431,N_3594,N_3244);
xor U5432 (N_5432,N_2611,N_3948);
or U5433 (N_5433,N_3308,N_2948);
nand U5434 (N_5434,N_4016,N_4157);
nand U5435 (N_5435,N_3973,N_4373);
xor U5436 (N_5436,N_4549,N_3378);
or U5437 (N_5437,N_3279,N_4019);
and U5438 (N_5438,N_4994,N_2682);
nand U5439 (N_5439,N_3720,N_4314);
xor U5440 (N_5440,N_4328,N_4042);
nand U5441 (N_5441,N_3293,N_4377);
and U5442 (N_5442,N_4165,N_3144);
nand U5443 (N_5443,N_4769,N_2954);
or U5444 (N_5444,N_2633,N_4023);
or U5445 (N_5445,N_4979,N_4099);
and U5446 (N_5446,N_4226,N_4532);
or U5447 (N_5447,N_2579,N_2621);
or U5448 (N_5448,N_3755,N_3440);
or U5449 (N_5449,N_3545,N_4117);
xnor U5450 (N_5450,N_3774,N_4395);
and U5451 (N_5451,N_4333,N_4196);
and U5452 (N_5452,N_4388,N_4465);
xnor U5453 (N_5453,N_4153,N_3073);
or U5454 (N_5454,N_3740,N_4551);
nor U5455 (N_5455,N_4837,N_4781);
or U5456 (N_5456,N_4699,N_3227);
and U5457 (N_5457,N_4685,N_4748);
or U5458 (N_5458,N_3462,N_2658);
nor U5459 (N_5459,N_2785,N_4163);
and U5460 (N_5460,N_4851,N_4864);
nor U5461 (N_5461,N_4151,N_4055);
and U5462 (N_5462,N_2522,N_2729);
xnor U5463 (N_5463,N_2710,N_3479);
nor U5464 (N_5464,N_3805,N_2831);
nor U5465 (N_5465,N_3396,N_4327);
or U5466 (N_5466,N_2562,N_2882);
xnor U5467 (N_5467,N_2892,N_2590);
or U5468 (N_5468,N_2516,N_3153);
or U5469 (N_5469,N_4332,N_4654);
or U5470 (N_5470,N_4847,N_3175);
xnor U5471 (N_5471,N_2825,N_4334);
nor U5472 (N_5472,N_4336,N_4384);
nand U5473 (N_5473,N_4745,N_3778);
xnor U5474 (N_5474,N_2505,N_4235);
nor U5475 (N_5475,N_2686,N_4885);
nand U5476 (N_5476,N_4182,N_3794);
xnor U5477 (N_5477,N_2972,N_3867);
and U5478 (N_5478,N_4020,N_4529);
nor U5479 (N_5479,N_4518,N_2848);
xnor U5480 (N_5480,N_3739,N_4081);
nor U5481 (N_5481,N_4367,N_3123);
or U5482 (N_5482,N_2958,N_4936);
nor U5483 (N_5483,N_3031,N_4457);
xor U5484 (N_5484,N_2813,N_4228);
nand U5485 (N_5485,N_2850,N_4242);
and U5486 (N_5486,N_4548,N_4619);
and U5487 (N_5487,N_3487,N_3919);
or U5488 (N_5488,N_3332,N_3780);
nor U5489 (N_5489,N_3401,N_4370);
nor U5490 (N_5490,N_3149,N_2837);
xor U5491 (N_5491,N_3431,N_3024);
xor U5492 (N_5492,N_2629,N_4975);
nor U5493 (N_5493,N_3807,N_3627);
or U5494 (N_5494,N_3531,N_3878);
nand U5495 (N_5495,N_4649,N_3134);
or U5496 (N_5496,N_2870,N_4486);
and U5497 (N_5497,N_3855,N_4587);
nor U5498 (N_5498,N_4629,N_2655);
nor U5499 (N_5499,N_3032,N_3317);
nand U5500 (N_5500,N_4789,N_4845);
nor U5501 (N_5501,N_4205,N_2707);
or U5502 (N_5502,N_4752,N_4089);
xor U5503 (N_5503,N_4349,N_2503);
nand U5504 (N_5504,N_4300,N_4018);
and U5505 (N_5505,N_4870,N_3469);
xor U5506 (N_5506,N_3364,N_2914);
nor U5507 (N_5507,N_4511,N_3381);
nand U5508 (N_5508,N_4919,N_4711);
nor U5509 (N_5509,N_3453,N_3668);
xor U5510 (N_5510,N_3513,N_2530);
nand U5511 (N_5511,N_2700,N_4024);
nor U5512 (N_5512,N_4596,N_3580);
or U5513 (N_5513,N_4921,N_3223);
nand U5514 (N_5514,N_3443,N_4473);
nand U5515 (N_5515,N_4858,N_4823);
or U5516 (N_5516,N_4398,N_2860);
or U5517 (N_5517,N_4684,N_3591);
or U5518 (N_5518,N_4943,N_3690);
xor U5519 (N_5519,N_2545,N_3758);
xor U5520 (N_5520,N_2965,N_2678);
xnor U5521 (N_5521,N_3572,N_3121);
or U5522 (N_5522,N_3379,N_4424);
and U5523 (N_5523,N_4462,N_2845);
and U5524 (N_5524,N_3242,N_2630);
nand U5525 (N_5525,N_2659,N_3336);
nor U5526 (N_5526,N_4755,N_3005);
xnor U5527 (N_5527,N_2970,N_4583);
or U5528 (N_5528,N_3064,N_3712);
nand U5529 (N_5529,N_3084,N_4798);
nand U5530 (N_5530,N_3480,N_4563);
nor U5531 (N_5531,N_4116,N_3873);
xnor U5532 (N_5532,N_3357,N_3272);
nand U5533 (N_5533,N_3889,N_4307);
xnor U5534 (N_5534,N_4278,N_4678);
nand U5535 (N_5535,N_3434,N_4470);
nor U5536 (N_5536,N_3972,N_2704);
nand U5537 (N_5537,N_3659,N_2650);
nand U5538 (N_5538,N_4133,N_3533);
nand U5539 (N_5539,N_4723,N_4981);
nor U5540 (N_5540,N_4128,N_3377);
nand U5541 (N_5541,N_3518,N_2849);
or U5542 (N_5542,N_2938,N_3812);
nand U5543 (N_5543,N_3380,N_3299);
and U5544 (N_5544,N_3187,N_4478);
and U5545 (N_5545,N_2616,N_4290);
and U5546 (N_5546,N_4679,N_4539);
or U5547 (N_5547,N_2502,N_4141);
or U5548 (N_5548,N_4521,N_3918);
nand U5549 (N_5549,N_3751,N_3528);
and U5550 (N_5550,N_4423,N_4632);
or U5551 (N_5551,N_2687,N_3856);
or U5552 (N_5552,N_4993,N_2558);
and U5553 (N_5553,N_4496,N_3145);
and U5554 (N_5554,N_2540,N_3615);
nand U5555 (N_5555,N_3942,N_4804);
nor U5556 (N_5556,N_2925,N_4793);
and U5557 (N_5557,N_4664,N_4063);
nand U5558 (N_5558,N_3517,N_2895);
and U5559 (N_5559,N_3498,N_3112);
xor U5560 (N_5560,N_2636,N_3548);
xor U5561 (N_5561,N_4582,N_3570);
nor U5562 (N_5562,N_3158,N_4190);
nor U5563 (N_5563,N_3872,N_4507);
xor U5564 (N_5564,N_3251,N_2547);
xnor U5565 (N_5565,N_4296,N_4094);
xnor U5566 (N_5566,N_3687,N_4876);
and U5567 (N_5567,N_4903,N_2835);
nand U5568 (N_5568,N_2574,N_2769);
and U5569 (N_5569,N_3155,N_4682);
xor U5570 (N_5570,N_4928,N_3779);
and U5571 (N_5571,N_3412,N_4156);
and U5572 (N_5572,N_2858,N_4573);
or U5573 (N_5573,N_2942,N_2865);
xor U5574 (N_5574,N_3460,N_4269);
nand U5575 (N_5575,N_3363,N_4091);
and U5576 (N_5576,N_4059,N_2507);
xnor U5577 (N_5577,N_3610,N_4962);
xor U5578 (N_5578,N_4856,N_4184);
xor U5579 (N_5579,N_3524,N_4216);
or U5580 (N_5580,N_2928,N_3819);
nand U5581 (N_5581,N_4997,N_2577);
nand U5582 (N_5582,N_4378,N_3491);
nand U5583 (N_5583,N_3140,N_4389);
and U5584 (N_5584,N_3103,N_4543);
nand U5585 (N_5585,N_4829,N_3993);
and U5586 (N_5586,N_4990,N_4970);
nand U5587 (N_5587,N_2660,N_4281);
nor U5588 (N_5588,N_4391,N_2525);
xnor U5589 (N_5589,N_4706,N_4475);
xor U5590 (N_5590,N_4794,N_3289);
nor U5591 (N_5591,N_4841,N_2677);
or U5592 (N_5592,N_4136,N_4760);
and U5593 (N_5593,N_3448,N_4077);
and U5594 (N_5594,N_4836,N_3003);
and U5595 (N_5595,N_3048,N_4553);
nand U5596 (N_5596,N_2509,N_3944);
nand U5597 (N_5597,N_2793,N_2554);
and U5598 (N_5598,N_3416,N_4325);
nor U5599 (N_5599,N_2598,N_4562);
or U5600 (N_5600,N_3848,N_3825);
nor U5601 (N_5601,N_3342,N_3920);
nand U5602 (N_5602,N_2684,N_2788);
or U5603 (N_5603,N_4779,N_4489);
and U5604 (N_5604,N_3652,N_4578);
or U5605 (N_5605,N_3354,N_4566);
nand U5606 (N_5606,N_4984,N_4929);
xor U5607 (N_5607,N_4967,N_3127);
nand U5608 (N_5608,N_2790,N_3159);
nor U5609 (N_5609,N_3880,N_3040);
nand U5610 (N_5610,N_2615,N_4857);
or U5611 (N_5611,N_4115,N_2513);
or U5612 (N_5612,N_4217,N_4159);
or U5613 (N_5613,N_4198,N_2833);
nand U5614 (N_5614,N_2797,N_3709);
nor U5615 (N_5615,N_4999,N_4775);
xor U5616 (N_5616,N_4110,N_4240);
nor U5617 (N_5617,N_4626,N_2852);
xor U5618 (N_5618,N_3014,N_3868);
nand U5619 (N_5619,N_2689,N_3141);
or U5620 (N_5620,N_2703,N_4076);
or U5621 (N_5621,N_4493,N_3514);
nand U5622 (N_5622,N_4834,N_3371);
and U5623 (N_5623,N_4344,N_3838);
nand U5624 (N_5624,N_2774,N_4622);
nand U5625 (N_5625,N_4983,N_4623);
or U5626 (N_5626,N_2555,N_3344);
nand U5627 (N_5627,N_4846,N_4031);
nor U5628 (N_5628,N_3964,N_3345);
or U5629 (N_5629,N_4050,N_4670);
or U5630 (N_5630,N_3542,N_3325);
or U5631 (N_5631,N_3902,N_4935);
or U5632 (N_5632,N_4087,N_3113);
nor U5633 (N_5633,N_4065,N_4036);
nand U5634 (N_5634,N_4989,N_4425);
and U5635 (N_5635,N_2538,N_3205);
nor U5636 (N_5636,N_4492,N_2571);
and U5637 (N_5637,N_2887,N_2923);
nor U5638 (N_5638,N_3093,N_4674);
nand U5639 (N_5639,N_3899,N_4402);
nor U5640 (N_5640,N_2913,N_3907);
and U5641 (N_5641,N_3669,N_4645);
nand U5642 (N_5642,N_4605,N_3171);
nand U5643 (N_5643,N_4559,N_4545);
nor U5644 (N_5644,N_3618,N_2875);
and U5645 (N_5645,N_3457,N_3165);
and U5646 (N_5646,N_2667,N_2796);
nand U5647 (N_5647,N_3349,N_3231);
nand U5648 (N_5648,N_3468,N_3905);
nand U5649 (N_5649,N_3248,N_2819);
nor U5650 (N_5650,N_3866,N_3428);
nand U5651 (N_5651,N_3571,N_2546);
or U5652 (N_5652,N_2712,N_3259);
nor U5653 (N_5653,N_2984,N_2992);
xnor U5654 (N_5654,N_4893,N_4306);
nand U5655 (N_5655,N_4255,N_4188);
or U5656 (N_5656,N_2625,N_2705);
nand U5657 (N_5657,N_4875,N_2758);
and U5658 (N_5658,N_2717,N_4224);
or U5659 (N_5659,N_3992,N_4740);
or U5660 (N_5660,N_3211,N_4862);
nand U5661 (N_5661,N_4570,N_4047);
nand U5662 (N_5662,N_2637,N_3634);
xor U5663 (N_5663,N_3875,N_4871);
xnor U5664 (N_5664,N_3177,N_4017);
nor U5665 (N_5665,N_4586,N_2955);
or U5666 (N_5666,N_2722,N_3235);
nand U5667 (N_5667,N_3190,N_4770);
nor U5668 (N_5668,N_3146,N_3749);
and U5669 (N_5669,N_4132,N_4832);
nand U5670 (N_5670,N_3326,N_3933);
xnor U5671 (N_5671,N_3644,N_4363);
xnor U5672 (N_5672,N_3925,N_4852);
xnor U5673 (N_5673,N_4448,N_3198);
nor U5674 (N_5674,N_3243,N_2504);
xnor U5675 (N_5675,N_4428,N_4572);
nor U5676 (N_5676,N_4311,N_2878);
xor U5677 (N_5677,N_3966,N_4609);
nand U5678 (N_5678,N_4167,N_3923);
nor U5679 (N_5679,N_3080,N_4634);
xor U5680 (N_5680,N_4109,N_4963);
nand U5681 (N_5681,N_3839,N_3643);
nand U5682 (N_5682,N_4121,N_3172);
or U5683 (N_5683,N_4728,N_4505);
or U5684 (N_5684,N_3636,N_4356);
nor U5685 (N_5685,N_2647,N_4700);
and U5686 (N_5686,N_2901,N_4720);
nor U5687 (N_5687,N_4754,N_4651);
nand U5688 (N_5688,N_4100,N_3642);
xor U5689 (N_5689,N_3621,N_3350);
nand U5690 (N_5690,N_4427,N_3890);
nand U5691 (N_5691,N_4828,N_2943);
nor U5692 (N_5692,N_3262,N_3568);
nor U5693 (N_5693,N_4208,N_4701);
nand U5694 (N_5694,N_2945,N_3814);
nand U5695 (N_5695,N_4264,N_4647);
nand U5696 (N_5696,N_3370,N_4108);
nand U5697 (N_5697,N_4445,N_2864);
xnor U5698 (N_5698,N_4661,N_2733);
or U5699 (N_5699,N_3833,N_4197);
nand U5700 (N_5700,N_3212,N_2966);
or U5701 (N_5701,N_4460,N_4374);
xor U5702 (N_5702,N_2695,N_4881);
nand U5703 (N_5703,N_4561,N_4189);
nand U5704 (N_5704,N_4199,N_3843);
xnor U5705 (N_5705,N_3552,N_4905);
nor U5706 (N_5706,N_3769,N_4029);
nor U5707 (N_5707,N_3811,N_4252);
nor U5708 (N_5708,N_2726,N_3921);
or U5709 (N_5709,N_4995,N_3264);
nand U5710 (N_5710,N_4001,N_3423);
and U5711 (N_5711,N_3221,N_3419);
or U5712 (N_5712,N_2778,N_3047);
nand U5713 (N_5713,N_3912,N_4782);
nand U5714 (N_5714,N_4376,N_2939);
nand U5715 (N_5715,N_2931,N_3684);
nor U5716 (N_5716,N_3483,N_4569);
nor U5717 (N_5717,N_4304,N_3310);
xor U5718 (N_5718,N_2715,N_3413);
and U5719 (N_5719,N_2968,N_4574);
nor U5720 (N_5720,N_3725,N_3062);
nor U5721 (N_5721,N_4057,N_4528);
nand U5722 (N_5722,N_3044,N_3138);
and U5723 (N_5723,N_4080,N_3598);
xnor U5724 (N_5724,N_4434,N_3771);
nor U5725 (N_5725,N_3249,N_4550);
nor U5726 (N_5726,N_3439,N_2669);
and U5727 (N_5727,N_4315,N_3865);
and U5728 (N_5728,N_4200,N_3271);
nor U5729 (N_5729,N_2768,N_3609);
or U5730 (N_5730,N_2638,N_4814);
nor U5731 (N_5731,N_4899,N_3624);
xnor U5732 (N_5732,N_4276,N_2714);
xor U5733 (N_5733,N_4005,N_2573);
or U5734 (N_5734,N_3276,N_4355);
nor U5735 (N_5735,N_3294,N_4491);
xor U5736 (N_5736,N_4286,N_3782);
xor U5737 (N_5737,N_3979,N_4454);
nor U5738 (N_5738,N_3466,N_4102);
nand U5739 (N_5739,N_4696,N_2929);
and U5740 (N_5740,N_4950,N_3768);
and U5741 (N_5741,N_3561,N_2654);
or U5742 (N_5742,N_2909,N_2518);
nor U5743 (N_5743,N_3295,N_2570);
or U5744 (N_5744,N_2500,N_2787);
xor U5745 (N_5745,N_3369,N_2932);
or U5746 (N_5746,N_4118,N_4337);
or U5747 (N_5747,N_2989,N_3874);
nor U5748 (N_5748,N_4513,N_4646);
nand U5749 (N_5749,N_3599,N_3893);
nor U5750 (N_5750,N_4131,N_3334);
and U5751 (N_5751,N_4112,N_4655);
xor U5752 (N_5752,N_3631,N_2956);
nor U5753 (N_5753,N_4293,N_2888);
xor U5754 (N_5754,N_3984,N_4880);
xnor U5755 (N_5755,N_3567,N_3685);
and U5756 (N_5756,N_3273,N_3841);
nor U5757 (N_5757,N_4236,N_4339);
nor U5758 (N_5758,N_4399,N_2991);
nor U5759 (N_5759,N_4688,N_2773);
nor U5760 (N_5760,N_4744,N_2921);
nor U5761 (N_5761,N_3280,N_4960);
or U5762 (N_5762,N_3441,N_3206);
xor U5763 (N_5763,N_3680,N_3196);
nand U5764 (N_5764,N_3662,N_4267);
nand U5765 (N_5765,N_4807,N_3676);
and U5766 (N_5766,N_4455,N_3229);
nand U5767 (N_5767,N_2924,N_3829);
or U5768 (N_5768,N_4418,N_3619);
and U5769 (N_5769,N_4957,N_4910);
and U5770 (N_5770,N_3553,N_2730);
or U5771 (N_5771,N_4992,N_2765);
nor U5772 (N_5772,N_4780,N_4597);
xor U5773 (N_5773,N_2781,N_4365);
nor U5774 (N_5774,N_3225,N_3564);
or U5775 (N_5775,N_4865,N_2815);
nor U5776 (N_5776,N_4524,N_4289);
xnor U5777 (N_5777,N_3915,N_4695);
nor U5778 (N_5778,N_4387,N_3929);
xor U5779 (N_5779,N_3029,N_3126);
nand U5780 (N_5780,N_2832,N_2624);
nand U5781 (N_5781,N_3458,N_3045);
xor U5782 (N_5782,N_4317,N_4379);
nor U5783 (N_5783,N_3554,N_4446);
or U5784 (N_5784,N_4044,N_3847);
and U5785 (N_5785,N_2944,N_3090);
nand U5786 (N_5786,N_4043,N_2904);
and U5787 (N_5787,N_2632,N_4771);
nor U5788 (N_5788,N_4900,N_2824);
nand U5789 (N_5789,N_3368,N_4026);
nor U5790 (N_5790,N_3510,N_4628);
nor U5791 (N_5791,N_4008,N_4873);
nor U5792 (N_5792,N_3351,N_3373);
nand U5793 (N_5793,N_4538,N_3604);
nor U5794 (N_5794,N_4687,N_4767);
and U5795 (N_5795,N_3331,N_2581);
or U5796 (N_5796,N_3208,N_4506);
xor U5797 (N_5797,N_3420,N_4523);
xnor U5798 (N_5798,N_3405,N_4764);
and U5799 (N_5799,N_2529,N_3962);
and U5800 (N_5800,N_3945,N_3056);
nand U5801 (N_5801,N_4362,N_3943);
or U5802 (N_5802,N_4884,N_3753);
nor U5803 (N_5803,N_4372,N_4122);
or U5804 (N_5804,N_2552,N_2840);
xnor U5805 (N_5805,N_3852,N_3298);
and U5806 (N_5806,N_4947,N_4069);
nor U5807 (N_5807,N_3637,N_4508);
and U5808 (N_5808,N_4127,N_3956);
and U5809 (N_5809,N_3004,N_3718);
nor U5810 (N_5810,N_3339,N_2688);
nor U5811 (N_5811,N_2997,N_3608);
nand U5812 (N_5812,N_3715,N_2595);
or U5813 (N_5813,N_3816,N_3157);
and U5814 (N_5814,N_3109,N_3649);
nand U5815 (N_5815,N_4126,N_2728);
xor U5816 (N_5816,N_2620,N_3922);
nor U5817 (N_5817,N_3623,N_4096);
nand U5818 (N_5818,N_3085,N_2935);
or U5819 (N_5819,N_3256,N_3595);
nand U5820 (N_5820,N_4371,N_4351);
or U5821 (N_5821,N_3395,N_4381);
and U5822 (N_5822,N_4991,N_4697);
xnor U5823 (N_5823,N_4436,N_3538);
and U5824 (N_5824,N_2512,N_2643);
nand U5825 (N_5825,N_4233,N_2946);
and U5826 (N_5826,N_4014,N_3651);
nor U5827 (N_5827,N_3409,N_3602);
nand U5828 (N_5828,N_3083,N_2916);
and U5829 (N_5829,N_4305,N_3287);
nand U5830 (N_5830,N_3585,N_3756);
and U5831 (N_5831,N_4616,N_3021);
nor U5832 (N_5832,N_2533,N_4129);
xor U5833 (N_5833,N_3641,N_2971);
nand U5834 (N_5834,N_4913,N_4612);
or U5835 (N_5835,N_2553,N_3472);
or U5836 (N_5836,N_3681,N_2767);
xnor U5837 (N_5837,N_3228,N_3981);
nor U5838 (N_5838,N_3108,N_4603);
nor U5839 (N_5839,N_2772,N_3188);
or U5840 (N_5840,N_2981,N_3746);
and U5841 (N_5841,N_3302,N_4849);
or U5842 (N_5842,N_3828,N_4011);
and U5843 (N_5843,N_4641,N_3114);
nor U5844 (N_5844,N_2582,N_2879);
and U5845 (N_5845,N_2830,N_3470);
nor U5846 (N_5846,N_4877,N_4826);
xnor U5847 (N_5847,N_3857,N_3218);
and U5848 (N_5848,N_3515,N_4124);
nand U5849 (N_5849,N_4459,N_4535);
xnor U5850 (N_5850,N_3655,N_3197);
and U5851 (N_5851,N_3560,N_4058);
nand U5852 (N_5852,N_2649,N_3220);
or U5853 (N_5853,N_4085,N_3490);
xor U5854 (N_5854,N_3731,N_3473);
nand U5855 (N_5855,N_3686,N_4140);
and U5856 (N_5856,N_2881,N_4730);
nand U5857 (N_5857,N_2575,N_3129);
nand U5858 (N_5858,N_4354,N_3485);
nand U5859 (N_5859,N_3241,N_3222);
nand U5860 (N_5860,N_3166,N_3445);
nand U5861 (N_5861,N_4887,N_4287);
nor U5862 (N_5862,N_3374,N_2569);
xor U5863 (N_5863,N_2930,N_4854);
and U5864 (N_5864,N_4393,N_4882);
and U5865 (N_5865,N_4564,N_4401);
nor U5866 (N_5866,N_3696,N_4966);
nor U5867 (N_5867,N_3579,N_4715);
xnor U5868 (N_5868,N_3763,N_4662);
or U5869 (N_5869,N_3267,N_4953);
nand U5870 (N_5870,N_4708,N_4827);
nor U5871 (N_5871,N_3292,N_3887);
nand U5872 (N_5872,N_3946,N_4920);
nor U5873 (N_5873,N_3463,N_3017);
or U5874 (N_5874,N_2635,N_3169);
nand U5875 (N_5875,N_4022,N_4690);
or U5876 (N_5876,N_3742,N_3060);
nand U5877 (N_5877,N_3424,N_3977);
and U5878 (N_5878,N_3124,N_3926);
and U5879 (N_5879,N_3237,N_4924);
and U5880 (N_5880,N_2528,N_4737);
and U5881 (N_5881,N_2631,N_3895);
nand U5882 (N_5882,N_4749,N_3156);
or U5883 (N_5883,N_3201,N_2962);
nor U5884 (N_5884,N_3994,N_4519);
nor U5885 (N_5885,N_4464,N_3754);
or U5886 (N_5886,N_4396,N_4490);
or U5887 (N_5887,N_4504,N_4433);
or U5888 (N_5888,N_4045,N_3663);
nand U5889 (N_5889,N_2810,N_4223);
nand U5890 (N_5890,N_4925,N_2514);
or U5891 (N_5891,N_4869,N_3135);
and U5892 (N_5892,N_3209,N_4229);
or U5893 (N_5893,N_2543,N_3041);
and U5894 (N_5894,N_4890,N_3529);
and U5895 (N_5895,N_3930,N_2823);
nor U5896 (N_5896,N_4672,N_3002);
and U5897 (N_5897,N_3741,N_3136);
xnor U5898 (N_5898,N_3411,N_2746);
xnor U5899 (N_5899,N_2844,N_4299);
and U5900 (N_5900,N_3735,N_4191);
nand U5901 (N_5901,N_3914,N_3693);
xor U5902 (N_5902,N_4250,N_4952);
nand U5903 (N_5903,N_4244,N_3131);
nor U5904 (N_5904,N_4207,N_4262);
xor U5905 (N_5905,N_2551,N_3549);
and U5906 (N_5906,N_4002,N_2883);
nand U5907 (N_5907,N_4757,N_3050);
and U5908 (N_5908,N_4139,N_3150);
nor U5909 (N_5909,N_3815,N_3710);
nor U5910 (N_5910,N_4657,N_4353);
or U5911 (N_5911,N_4731,N_3563);
nor U5912 (N_5912,N_3835,N_4763);
xor U5913 (N_5913,N_4541,N_2940);
nor U5914 (N_5914,N_4027,N_4348);
xor U5915 (N_5915,N_3115,N_2662);
xor U5916 (N_5916,N_3234,N_3603);
xnor U5917 (N_5917,N_3512,N_3646);
nor U5918 (N_5918,N_2685,N_2862);
or U5919 (N_5919,N_4125,N_3306);
xor U5920 (N_5920,N_4509,N_4284);
and U5921 (N_5921,N_3987,N_3982);
and U5922 (N_5922,N_3937,N_4285);
xor U5923 (N_5923,N_4456,N_3494);
and U5924 (N_5924,N_3319,N_3883);
nor U5925 (N_5925,N_3584,N_4301);
or U5926 (N_5926,N_3315,N_4567);
nor U5927 (N_5927,N_2980,N_3274);
and U5928 (N_5928,N_4386,N_3892);
or U5929 (N_5929,N_3035,N_4802);
and U5930 (N_5930,N_3675,N_3522);
xor U5931 (N_5931,N_4677,N_2701);
or U5932 (N_5932,N_3556,N_3255);
nand U5933 (N_5933,N_4426,N_4313);
nor U5934 (N_5934,N_3617,N_3582);
nor U5935 (N_5935,N_2743,N_3969);
nor U5936 (N_5936,N_3061,N_4175);
xor U5937 (N_5937,N_4095,N_3199);
or U5938 (N_5938,N_3246,N_3645);
xnor U5939 (N_5939,N_3938,N_3039);
xnor U5940 (N_5940,N_4051,N_2645);
and U5941 (N_5941,N_3949,N_2580);
nand U5942 (N_5942,N_4397,N_4086);
and U5943 (N_5943,N_4980,N_3484);
nand U5944 (N_5944,N_3541,N_3898);
nor U5945 (N_5945,N_4878,N_3421);
and U5946 (N_5946,N_4006,N_3810);
and U5947 (N_5947,N_4147,N_3324);
xnor U5948 (N_5948,N_3989,N_3577);
nor U5949 (N_5949,N_4352,N_2517);
nor U5950 (N_5950,N_3027,N_4556);
or U5951 (N_5951,N_3776,N_2641);
and U5952 (N_5952,N_3804,N_4090);
and U5953 (N_5953,N_2885,N_4705);
nand U5954 (N_5954,N_3616,N_3648);
xnor U5955 (N_5955,N_2873,N_4707);
xor U5956 (N_5956,N_4669,N_2676);
or U5957 (N_5957,N_3055,N_4246);
nand U5958 (N_5958,N_4410,N_4515);
nand U5959 (N_5959,N_2578,N_2539);
nor U5960 (N_5960,N_4776,N_2642);
xnor U5961 (N_5961,N_4484,N_3391);
nand U5962 (N_5962,N_4170,N_3677);
nor U5963 (N_5963,N_4437,N_4932);
xor U5964 (N_5964,N_3022,N_2537);
xor U5965 (N_5965,N_3882,N_2612);
and U5966 (N_5966,N_3850,N_4795);
nor U5967 (N_5967,N_3673,N_4897);
nor U5968 (N_5968,N_4054,N_2841);
nand U5969 (N_5969,N_4956,N_3764);
and U5970 (N_5970,N_3854,N_3049);
xnor U5971 (N_5971,N_4111,N_4941);
xnor U5972 (N_5972,N_4624,N_3015);
xnor U5973 (N_5973,N_2523,N_4227);
and U5974 (N_5974,N_3019,N_3653);
or U5975 (N_5975,N_2891,N_2600);
xor U5976 (N_5976,N_3500,N_4469);
or U5977 (N_5977,N_4691,N_3759);
and U5978 (N_5978,N_2613,N_3415);
or U5979 (N_5979,N_3414,N_3635);
or U5980 (N_5980,N_4914,N_4297);
xor U5981 (N_5981,N_4618,N_4765);
nand U5982 (N_5982,N_2651,N_2639);
xor U5983 (N_5983,N_2691,N_3046);
nor U5984 (N_5984,N_2747,N_3418);
and U5985 (N_5985,N_4594,N_3404);
xnor U5986 (N_5986,N_3574,N_2657);
nor U5987 (N_5987,N_3953,N_4736);
nor U5988 (N_5988,N_4030,N_4321);
or U5989 (N_5989,N_3877,N_4734);
or U5990 (N_5990,N_2755,N_2866);
or U5991 (N_5991,N_4053,N_3347);
nor U5992 (N_5992,N_3832,N_3269);
nor U5993 (N_5993,N_2607,N_3089);
nor U5994 (N_5994,N_3853,N_3692);
nand U5995 (N_5995,N_4591,N_4911);
nand U5996 (N_5996,N_3961,N_2861);
nand U5997 (N_5997,N_3125,N_4825);
nand U5998 (N_5998,N_3281,N_4874);
nand U5999 (N_5999,N_4164,N_3341);
xnor U6000 (N_6000,N_2834,N_2963);
xor U6001 (N_6001,N_4345,N_3916);
and U6002 (N_6002,N_4520,N_2626);
and U6003 (N_6003,N_4390,N_3328);
xor U6004 (N_6004,N_2936,N_3800);
nor U6005 (N_6005,N_3101,N_4272);
and U6006 (N_6006,N_4702,N_3034);
xor U6007 (N_6007,N_3911,N_4481);
or U6008 (N_6008,N_3467,N_3744);
nand U6009 (N_6009,N_4592,N_3959);
nor U6010 (N_6010,N_3647,N_4186);
nand U6011 (N_6011,N_2751,N_3068);
or U6012 (N_6012,N_3978,N_2608);
nand U6013 (N_6013,N_3475,N_3786);
and U6014 (N_6014,N_3975,N_4738);
xor U6015 (N_6015,N_4416,N_4998);
or U6016 (N_6016,N_4274,N_2816);
nand U6017 (N_6017,N_2994,N_3304);
and U6018 (N_6018,N_2719,N_4812);
or U6019 (N_6019,N_3534,N_3704);
xnor U6020 (N_6020,N_4500,N_3705);
or U6021 (N_6021,N_4394,N_2789);
and U6022 (N_6022,N_2749,N_3427);
and U6023 (N_6023,N_3886,N_3087);
xnor U6024 (N_6024,N_3530,N_4571);
xor U6025 (N_6025,N_2668,N_2809);
xnor U6026 (N_6026,N_4201,N_3507);
and U6027 (N_6027,N_2602,N_3191);
or U6028 (N_6028,N_2771,N_4049);
xnor U6029 (N_6029,N_2806,N_4689);
and U6030 (N_6030,N_3980,N_4901);
nor U6031 (N_6031,N_3110,N_4012);
nand U6032 (N_6032,N_2606,N_2933);
nand U6033 (N_6033,N_3288,N_4072);
nand U6034 (N_6034,N_3509,N_4021);
or U6035 (N_6035,N_3908,N_4813);
and U6036 (N_6036,N_2698,N_4889);
xor U6037 (N_6037,N_4888,N_4092);
and U6038 (N_6038,N_3913,N_2953);
nand U6039 (N_6039,N_3881,N_3985);
or U6040 (N_6040,N_4729,N_3065);
nor U6041 (N_6041,N_3817,N_4247);
or U6042 (N_6042,N_4383,N_2564);
xnor U6043 (N_6043,N_4806,N_3656);
or U6044 (N_6044,N_3203,N_3120);
nor U6045 (N_6045,N_4443,N_2898);
xor U6046 (N_6046,N_4417,N_3974);
nor U6047 (N_6047,N_3097,N_4070);
or U6048 (N_6048,N_4143,N_4361);
nand U6049 (N_6049,N_4056,N_3781);
or U6050 (N_6050,N_3007,N_3702);
nor U6051 (N_6051,N_3385,N_4079);
nand U6052 (N_6052,N_4772,N_3558);
and U6053 (N_6053,N_3752,N_4977);
or U6054 (N_6054,N_4973,N_3086);
nand U6055 (N_6055,N_3282,N_4907);
and U6056 (N_6056,N_2696,N_4450);
nand U6057 (N_6057,N_3447,N_3939);
xnor U6058 (N_6058,N_3253,N_2501);
nand U6059 (N_6059,N_4340,N_3254);
or U6060 (N_6060,N_2506,N_3186);
nand U6061 (N_6061,N_2576,N_3665);
and U6062 (N_6062,N_4218,N_4650);
xor U6063 (N_6063,N_4312,N_4822);
and U6064 (N_6064,N_4675,N_4965);
and U6065 (N_6065,N_2567,N_2838);
nand U6066 (N_6066,N_4902,N_4922);
and U6067 (N_6067,N_3337,N_3173);
nand U6068 (N_6068,N_4820,N_4282);
and U6069 (N_6069,N_4839,N_3495);
xor U6070 (N_6070,N_2969,N_4615);
nor U6071 (N_6071,N_4028,N_3678);
and U6072 (N_6072,N_3152,N_4671);
nand U6073 (N_6073,N_3729,N_3074);
and U6074 (N_6074,N_2820,N_4821);
nand U6075 (N_6075,N_3063,N_4951);
xor U6076 (N_6076,N_3030,N_4741);
xor U6077 (N_6077,N_4722,N_3230);
or U6078 (N_6078,N_2886,N_3320);
nor U6079 (N_6079,N_2853,N_3406);
nor U6080 (N_6080,N_3459,N_3869);
xnor U6081 (N_6081,N_3727,N_2777);
nor U6082 (N_6082,N_4106,N_3329);
nor U6083 (N_6083,N_4788,N_4978);
nand U6084 (N_6084,N_3901,N_4824);
xor U6085 (N_6085,N_3471,N_4512);
nor U6086 (N_6086,N_4796,N_4494);
xor U6087 (N_6087,N_3697,N_4329);
nand U6088 (N_6088,N_3200,N_2723);
xnor U6089 (N_6089,N_3245,N_3936);
nand U6090 (N_6090,N_3233,N_2610);
nand U6091 (N_6091,N_2905,N_3143);
and U6092 (N_6092,N_4249,N_3699);
and U6093 (N_6093,N_3455,N_2974);
xor U6094 (N_6094,N_3318,N_3346);
nor U6095 (N_6095,N_4452,N_3180);
and U6096 (N_6096,N_3539,N_3605);
xnor U6097 (N_6097,N_4931,N_4800);
nor U6098 (N_6098,N_3821,N_3133);
xnor U6099 (N_6099,N_2763,N_3827);
nand U6100 (N_6100,N_3860,N_2563);
or U6101 (N_6101,N_2918,N_3436);
and U6102 (N_6102,N_3995,N_4599);
or U6103 (N_6103,N_4144,N_3957);
xor U6104 (N_6104,N_4639,N_2762);
and U6105 (N_6105,N_4467,N_2911);
nand U6106 (N_6106,N_4308,N_3639);
nand U6107 (N_6107,N_3802,N_3963);
and U6108 (N_6108,N_4039,N_4576);
xor U6109 (N_6109,N_4238,N_4444);
or U6110 (N_6110,N_2679,N_3023);
nor U6111 (N_6111,N_4718,N_4160);
xor U6112 (N_6112,N_3683,N_3464);
nand U6113 (N_6113,N_2565,N_4855);
nor U6114 (N_6114,N_4961,N_3266);
and U6115 (N_6115,N_4342,N_4256);
nand U6116 (N_6116,N_2713,N_4517);
nand U6117 (N_6117,N_4214,N_3660);
or U6118 (N_6118,N_3128,N_2917);
and U6119 (N_6119,N_3765,N_2826);
nand U6120 (N_6120,N_3390,N_4488);
xor U6121 (N_6121,N_4710,N_4560);
and U6122 (N_6122,N_4032,N_4212);
xor U6123 (N_6123,N_3885,N_3508);
nor U6124 (N_6124,N_3679,N_3482);
or U6125 (N_6125,N_3099,N_4195);
nor U6126 (N_6126,N_4137,N_2757);
and U6127 (N_6127,N_4667,N_3285);
xnor U6128 (N_6128,N_2734,N_2854);
nor U6129 (N_6129,N_3263,N_3091);
nand U6130 (N_6130,N_2869,N_3359);
and U6131 (N_6131,N_2690,N_2692);
nand U6132 (N_6132,N_3216,N_3998);
nand U6133 (N_6133,N_4726,N_3900);
xnor U6134 (N_6134,N_2583,N_4568);
and U6135 (N_6135,N_4181,N_4330);
nor U6136 (N_6136,N_4750,N_4368);
or U6137 (N_6137,N_2742,N_2515);
xor U6138 (N_6138,N_4003,N_4680);
and U6139 (N_6139,N_3094,N_3733);
nand U6140 (N_6140,N_4103,N_3316);
nor U6141 (N_6141,N_2784,N_4811);
nor U6142 (N_6142,N_4010,N_4048);
nand U6143 (N_6143,N_2821,N_3425);
and U6144 (N_6144,N_2725,N_2585);
or U6145 (N_6145,N_4527,N_2619);
nor U6146 (N_6146,N_3790,N_4408);
and U6147 (N_6147,N_4938,N_4380);
nand U6148 (N_6148,N_3214,N_4422);
nor U6149 (N_6149,N_3588,N_3958);
or U6150 (N_6150,N_3000,N_4724);
xnor U6151 (N_6151,N_4295,N_2740);
and U6152 (N_6152,N_4407,N_3762);
nand U6153 (N_6153,N_4346,N_3408);
nor U6154 (N_6154,N_3488,N_3154);
and U6155 (N_6155,N_3569,N_4347);
xnor U6156 (N_6156,N_3454,N_3433);
xnor U6157 (N_6157,N_4892,N_3435);
or U6158 (N_6158,N_2786,N_2985);
xor U6159 (N_6159,N_3450,N_4894);
nor U6160 (N_6160,N_3388,N_2867);
xnor U6161 (N_6161,N_4495,N_3016);
nand U6162 (N_6162,N_2919,N_3559);
nor U6163 (N_6163,N_2770,N_4210);
nor U6164 (N_6164,N_4756,N_3622);
and U6165 (N_6165,N_3760,N_4585);
and U6166 (N_6166,N_3092,N_3139);
nor U6167 (N_6167,N_3151,N_4013);
xnor U6168 (N_6168,N_2993,N_3870);
xor U6169 (N_6169,N_2884,N_4245);
nand U6170 (N_6170,N_4918,N_3054);
nor U6171 (N_6171,N_4310,N_3934);
or U6172 (N_6172,N_2926,N_2976);
nor U6173 (N_6173,N_3088,N_3185);
nor U6174 (N_6174,N_3576,N_4673);
nor U6175 (N_6175,N_3012,N_2903);
nor U6176 (N_6176,N_3738,N_3215);
and U6177 (N_6177,N_3830,N_4241);
xor U6178 (N_6178,N_3747,N_4816);
xor U6179 (N_6179,N_4840,N_2986);
and U6180 (N_6180,N_4322,N_3444);
nand U6181 (N_6181,N_3654,N_3797);
and U6182 (N_6182,N_3968,N_4411);
xor U6183 (N_6183,N_3547,N_2741);
xor U6184 (N_6184,N_3297,N_2920);
nor U6185 (N_6185,N_4660,N_4502);
and U6186 (N_6186,N_2592,N_4453);
and U6187 (N_6187,N_4154,N_4959);
or U6188 (N_6188,N_3726,N_4270);
nand U6189 (N_6189,N_3286,N_4546);
or U6190 (N_6190,N_2664,N_3640);
and U6191 (N_6191,N_4263,N_3795);
and U6192 (N_6192,N_3629,N_3935);
nor U6193 (N_6193,N_3671,N_3338);
nor U6194 (N_6194,N_4225,N_2847);
and U6195 (N_6195,N_3179,N_2572);
nand U6196 (N_6196,N_3477,N_4254);
or U6197 (N_6197,N_3820,N_3664);
nor U6198 (N_6198,N_3181,N_4098);
nand U6199 (N_6199,N_2927,N_4525);
or U6200 (N_6200,N_4537,N_3505);
nor U6201 (N_6201,N_3183,N_2609);
xor U6202 (N_6202,N_4642,N_2794);
nand U6203 (N_6203,N_2653,N_4863);
nor U6204 (N_6204,N_4733,N_4430);
and U6205 (N_6205,N_4283,N_2843);
or U6206 (N_6206,N_3168,N_4061);
nand U6207 (N_6207,N_2599,N_3719);
nor U6208 (N_6208,N_3798,N_2510);
nand U6209 (N_6209,N_3258,N_4166);
nand U6210 (N_6210,N_3511,N_2557);
nand U6211 (N_6211,N_2811,N_2874);
or U6212 (N_6212,N_4146,N_4480);
and U6213 (N_6213,N_4808,N_4968);
and U6214 (N_6214,N_2988,N_4358);
xnor U6215 (N_6215,N_4536,N_2902);
xnor U6216 (N_6216,N_4419,N_2979);
or U6217 (N_6217,N_2896,N_2594);
nor U6218 (N_6218,N_3721,N_3107);
or U6219 (N_6219,N_3906,N_4516);
and U6220 (N_6220,N_3791,N_2586);
xnor U6221 (N_6221,N_3305,N_4230);
nand U6222 (N_6222,N_3358,N_4360);
nor U6223 (N_6223,N_4202,N_2906);
nand U6224 (N_6224,N_4554,N_3551);
xor U6225 (N_6225,N_4916,N_3313);
xnor U6226 (N_6226,N_3309,N_3116);
xnor U6227 (N_6227,N_2587,N_4041);
and U6228 (N_6228,N_2536,N_4474);
nor U6229 (N_6229,N_4060,N_4415);
nand U6230 (N_6230,N_3773,N_4403);
and U6231 (N_6231,N_4501,N_4220);
nor U6232 (N_6232,N_4644,N_4194);
and U6233 (N_6233,N_3955,N_4758);
or U6234 (N_6234,N_3770,N_3674);
or U6235 (N_6235,N_4712,N_2702);
and U6236 (N_6236,N_4499,N_3611);
and U6237 (N_6237,N_4648,N_3137);
nor U6238 (N_6238,N_3836,N_3502);
or U6239 (N_6239,N_4971,N_4818);
xnor U6240 (N_6240,N_3184,N_4177);
nand U6241 (N_6241,N_4625,N_2872);
and U6242 (N_6242,N_3043,N_2973);
and U6243 (N_6243,N_3142,N_3130);
and U6244 (N_6244,N_4073,N_3876);
or U6245 (N_6245,N_4341,N_3788);
nor U6246 (N_6246,N_4891,N_3592);
or U6247 (N_6247,N_3707,N_2716);
or U6248 (N_6248,N_2681,N_4759);
and U6249 (N_6249,N_4627,N_2604);
xnor U6250 (N_6250,N_3080,N_3516);
and U6251 (N_6251,N_3633,N_4001);
nor U6252 (N_6252,N_4051,N_2812);
xnor U6253 (N_6253,N_4244,N_3902);
nor U6254 (N_6254,N_3017,N_3006);
and U6255 (N_6255,N_4997,N_3894);
nand U6256 (N_6256,N_3174,N_3877);
xor U6257 (N_6257,N_3602,N_2610);
or U6258 (N_6258,N_4366,N_4412);
nor U6259 (N_6259,N_4709,N_3069);
nand U6260 (N_6260,N_2565,N_3612);
nor U6261 (N_6261,N_4527,N_3110);
or U6262 (N_6262,N_3150,N_2920);
xnor U6263 (N_6263,N_4712,N_4247);
nand U6264 (N_6264,N_4105,N_3941);
nand U6265 (N_6265,N_3932,N_4385);
nand U6266 (N_6266,N_3339,N_2641);
and U6267 (N_6267,N_4653,N_3701);
nand U6268 (N_6268,N_3810,N_4252);
nand U6269 (N_6269,N_3400,N_3829);
nand U6270 (N_6270,N_3541,N_4657);
xor U6271 (N_6271,N_3774,N_3455);
nand U6272 (N_6272,N_4762,N_4476);
and U6273 (N_6273,N_4150,N_3909);
nand U6274 (N_6274,N_3323,N_4918);
nor U6275 (N_6275,N_4806,N_3779);
xor U6276 (N_6276,N_3983,N_2854);
and U6277 (N_6277,N_3139,N_2808);
nor U6278 (N_6278,N_2871,N_3946);
nor U6279 (N_6279,N_3701,N_4664);
xnor U6280 (N_6280,N_4644,N_3940);
nor U6281 (N_6281,N_4731,N_3633);
nand U6282 (N_6282,N_3170,N_3954);
nor U6283 (N_6283,N_3207,N_4574);
and U6284 (N_6284,N_4045,N_3571);
xor U6285 (N_6285,N_4335,N_4275);
or U6286 (N_6286,N_3002,N_3596);
nor U6287 (N_6287,N_3231,N_4593);
or U6288 (N_6288,N_4176,N_3319);
and U6289 (N_6289,N_4464,N_3482);
or U6290 (N_6290,N_4846,N_4977);
nor U6291 (N_6291,N_4403,N_4163);
nor U6292 (N_6292,N_2928,N_3982);
nand U6293 (N_6293,N_2563,N_4055);
or U6294 (N_6294,N_4318,N_2626);
and U6295 (N_6295,N_2843,N_4873);
and U6296 (N_6296,N_2811,N_4075);
or U6297 (N_6297,N_4651,N_4960);
nand U6298 (N_6298,N_2546,N_4342);
xnor U6299 (N_6299,N_4318,N_3454);
nand U6300 (N_6300,N_4655,N_4882);
xnor U6301 (N_6301,N_3443,N_3729);
or U6302 (N_6302,N_3922,N_2920);
or U6303 (N_6303,N_4759,N_4016);
and U6304 (N_6304,N_3606,N_2838);
or U6305 (N_6305,N_3941,N_4285);
or U6306 (N_6306,N_3716,N_3340);
xor U6307 (N_6307,N_4353,N_3630);
xnor U6308 (N_6308,N_3519,N_3110);
xnor U6309 (N_6309,N_4389,N_4147);
nor U6310 (N_6310,N_4095,N_4093);
and U6311 (N_6311,N_3530,N_4214);
and U6312 (N_6312,N_4934,N_4037);
nor U6313 (N_6313,N_2517,N_4999);
nor U6314 (N_6314,N_3689,N_3867);
nor U6315 (N_6315,N_4037,N_2702);
nor U6316 (N_6316,N_4470,N_2547);
nor U6317 (N_6317,N_4626,N_4995);
nand U6318 (N_6318,N_3788,N_3700);
xnor U6319 (N_6319,N_2794,N_2886);
nand U6320 (N_6320,N_3834,N_3231);
and U6321 (N_6321,N_4987,N_4503);
and U6322 (N_6322,N_3621,N_3277);
nor U6323 (N_6323,N_3274,N_2996);
nor U6324 (N_6324,N_4715,N_3979);
nor U6325 (N_6325,N_3770,N_2988);
nor U6326 (N_6326,N_4361,N_3318);
xnor U6327 (N_6327,N_4388,N_3216);
nor U6328 (N_6328,N_4004,N_4247);
nand U6329 (N_6329,N_4181,N_3581);
nor U6330 (N_6330,N_3383,N_3258);
nor U6331 (N_6331,N_3866,N_2627);
or U6332 (N_6332,N_2598,N_3942);
or U6333 (N_6333,N_3934,N_3388);
or U6334 (N_6334,N_4050,N_3379);
or U6335 (N_6335,N_4334,N_3559);
or U6336 (N_6336,N_3144,N_3251);
nand U6337 (N_6337,N_2813,N_3197);
nor U6338 (N_6338,N_4115,N_3076);
nor U6339 (N_6339,N_3514,N_4655);
or U6340 (N_6340,N_2694,N_4696);
xnor U6341 (N_6341,N_3464,N_4984);
or U6342 (N_6342,N_3225,N_4067);
nand U6343 (N_6343,N_3461,N_4397);
or U6344 (N_6344,N_3540,N_4473);
xnor U6345 (N_6345,N_4097,N_2888);
and U6346 (N_6346,N_3719,N_3515);
and U6347 (N_6347,N_3488,N_2584);
and U6348 (N_6348,N_3372,N_4248);
xnor U6349 (N_6349,N_3355,N_4695);
or U6350 (N_6350,N_3367,N_3189);
nand U6351 (N_6351,N_4656,N_2881);
and U6352 (N_6352,N_2606,N_2819);
xor U6353 (N_6353,N_4599,N_3541);
and U6354 (N_6354,N_3628,N_3500);
xor U6355 (N_6355,N_3477,N_2770);
and U6356 (N_6356,N_2596,N_3169);
xnor U6357 (N_6357,N_3493,N_4844);
xnor U6358 (N_6358,N_4057,N_3935);
and U6359 (N_6359,N_3727,N_3028);
nand U6360 (N_6360,N_4341,N_3448);
and U6361 (N_6361,N_4226,N_3952);
and U6362 (N_6362,N_3876,N_2987);
nor U6363 (N_6363,N_2726,N_4380);
xnor U6364 (N_6364,N_4137,N_4648);
and U6365 (N_6365,N_2601,N_4053);
xor U6366 (N_6366,N_2564,N_2983);
and U6367 (N_6367,N_3481,N_3532);
and U6368 (N_6368,N_4748,N_4717);
nand U6369 (N_6369,N_3856,N_3701);
nand U6370 (N_6370,N_4825,N_4201);
nand U6371 (N_6371,N_4750,N_3014);
or U6372 (N_6372,N_4009,N_2695);
xor U6373 (N_6373,N_3673,N_4976);
or U6374 (N_6374,N_3863,N_3876);
or U6375 (N_6375,N_4387,N_3453);
and U6376 (N_6376,N_3237,N_2716);
and U6377 (N_6377,N_4995,N_3036);
nor U6378 (N_6378,N_4478,N_3754);
and U6379 (N_6379,N_3419,N_4817);
nand U6380 (N_6380,N_4578,N_2694);
or U6381 (N_6381,N_4839,N_2966);
nand U6382 (N_6382,N_3399,N_3600);
nor U6383 (N_6383,N_4009,N_2561);
and U6384 (N_6384,N_3118,N_3679);
nor U6385 (N_6385,N_4043,N_3783);
nor U6386 (N_6386,N_2783,N_4006);
nor U6387 (N_6387,N_3749,N_3592);
xnor U6388 (N_6388,N_4538,N_3506);
nor U6389 (N_6389,N_4917,N_4071);
or U6390 (N_6390,N_3912,N_3646);
or U6391 (N_6391,N_3783,N_2862);
and U6392 (N_6392,N_2882,N_3665);
and U6393 (N_6393,N_3725,N_4092);
nand U6394 (N_6394,N_3733,N_4550);
nor U6395 (N_6395,N_4683,N_3371);
nand U6396 (N_6396,N_4877,N_3802);
nor U6397 (N_6397,N_4321,N_4873);
xnor U6398 (N_6398,N_4106,N_4436);
xor U6399 (N_6399,N_4730,N_3194);
xor U6400 (N_6400,N_3659,N_4549);
nor U6401 (N_6401,N_4958,N_4938);
nor U6402 (N_6402,N_3767,N_4410);
nand U6403 (N_6403,N_4407,N_3980);
nor U6404 (N_6404,N_3061,N_2984);
or U6405 (N_6405,N_4930,N_3328);
xnor U6406 (N_6406,N_3784,N_4689);
nand U6407 (N_6407,N_3490,N_4104);
xor U6408 (N_6408,N_4033,N_2561);
xor U6409 (N_6409,N_4202,N_2889);
nor U6410 (N_6410,N_4387,N_4824);
nand U6411 (N_6411,N_4435,N_4573);
or U6412 (N_6412,N_2867,N_4836);
nor U6413 (N_6413,N_3181,N_3543);
xnor U6414 (N_6414,N_4188,N_2778);
and U6415 (N_6415,N_3257,N_3267);
xor U6416 (N_6416,N_2582,N_2532);
nor U6417 (N_6417,N_4684,N_4653);
and U6418 (N_6418,N_4529,N_4705);
or U6419 (N_6419,N_3114,N_3086);
nor U6420 (N_6420,N_4940,N_3608);
nor U6421 (N_6421,N_4420,N_3001);
nand U6422 (N_6422,N_4804,N_4438);
or U6423 (N_6423,N_4652,N_3011);
nor U6424 (N_6424,N_4050,N_3200);
nor U6425 (N_6425,N_4331,N_4092);
nand U6426 (N_6426,N_4459,N_3147);
xnor U6427 (N_6427,N_2600,N_2561);
and U6428 (N_6428,N_3423,N_3680);
nand U6429 (N_6429,N_4552,N_3799);
nand U6430 (N_6430,N_3207,N_4455);
nand U6431 (N_6431,N_4171,N_3842);
or U6432 (N_6432,N_4048,N_3044);
xnor U6433 (N_6433,N_4522,N_3368);
nand U6434 (N_6434,N_4780,N_2649);
or U6435 (N_6435,N_4701,N_3068);
nand U6436 (N_6436,N_3887,N_2658);
nor U6437 (N_6437,N_4707,N_3255);
xnor U6438 (N_6438,N_4454,N_2546);
or U6439 (N_6439,N_2696,N_4236);
nand U6440 (N_6440,N_4993,N_3342);
nor U6441 (N_6441,N_3052,N_4212);
and U6442 (N_6442,N_3296,N_3607);
and U6443 (N_6443,N_4533,N_2894);
nor U6444 (N_6444,N_3980,N_3752);
or U6445 (N_6445,N_3880,N_3277);
or U6446 (N_6446,N_2532,N_4177);
and U6447 (N_6447,N_3963,N_4261);
xor U6448 (N_6448,N_2631,N_4788);
nor U6449 (N_6449,N_3417,N_4234);
nand U6450 (N_6450,N_2720,N_4484);
and U6451 (N_6451,N_2615,N_3402);
and U6452 (N_6452,N_3786,N_4640);
xor U6453 (N_6453,N_2998,N_3038);
xor U6454 (N_6454,N_3213,N_4751);
nor U6455 (N_6455,N_4123,N_4729);
xnor U6456 (N_6456,N_4146,N_4885);
or U6457 (N_6457,N_4563,N_4562);
nand U6458 (N_6458,N_3782,N_4224);
xnor U6459 (N_6459,N_3800,N_3524);
and U6460 (N_6460,N_3549,N_2577);
xor U6461 (N_6461,N_2674,N_3054);
xor U6462 (N_6462,N_4196,N_3363);
and U6463 (N_6463,N_3145,N_3243);
xnor U6464 (N_6464,N_4106,N_3587);
and U6465 (N_6465,N_3538,N_4752);
xnor U6466 (N_6466,N_3608,N_3411);
and U6467 (N_6467,N_3690,N_3875);
nor U6468 (N_6468,N_2787,N_3381);
xnor U6469 (N_6469,N_3530,N_3337);
xnor U6470 (N_6470,N_3633,N_3612);
or U6471 (N_6471,N_4639,N_2840);
and U6472 (N_6472,N_4952,N_2909);
or U6473 (N_6473,N_3870,N_2655);
xor U6474 (N_6474,N_4701,N_4283);
xor U6475 (N_6475,N_4964,N_4910);
or U6476 (N_6476,N_3852,N_3747);
nor U6477 (N_6477,N_4419,N_3072);
or U6478 (N_6478,N_4500,N_2934);
xnor U6479 (N_6479,N_3095,N_3818);
nand U6480 (N_6480,N_4236,N_3012);
nor U6481 (N_6481,N_4777,N_4004);
nor U6482 (N_6482,N_3374,N_3326);
nand U6483 (N_6483,N_3881,N_3701);
nor U6484 (N_6484,N_3213,N_3458);
and U6485 (N_6485,N_3053,N_2963);
and U6486 (N_6486,N_4329,N_4420);
and U6487 (N_6487,N_4655,N_4413);
or U6488 (N_6488,N_3798,N_2775);
xnor U6489 (N_6489,N_3685,N_3184);
xnor U6490 (N_6490,N_4260,N_3358);
or U6491 (N_6491,N_3704,N_2737);
nand U6492 (N_6492,N_4019,N_2549);
xor U6493 (N_6493,N_4620,N_4023);
nand U6494 (N_6494,N_3792,N_3804);
nor U6495 (N_6495,N_2947,N_2518);
xor U6496 (N_6496,N_3636,N_4485);
and U6497 (N_6497,N_4260,N_2774);
xnor U6498 (N_6498,N_4087,N_4629);
or U6499 (N_6499,N_3840,N_4053);
nand U6500 (N_6500,N_4895,N_4812);
and U6501 (N_6501,N_4805,N_2545);
nor U6502 (N_6502,N_3580,N_4154);
nor U6503 (N_6503,N_3560,N_2891);
or U6504 (N_6504,N_4451,N_4472);
nand U6505 (N_6505,N_3949,N_4304);
nor U6506 (N_6506,N_2976,N_4316);
or U6507 (N_6507,N_4447,N_2673);
nand U6508 (N_6508,N_2900,N_4804);
xor U6509 (N_6509,N_3439,N_2587);
or U6510 (N_6510,N_3874,N_3702);
nand U6511 (N_6511,N_4674,N_4712);
xnor U6512 (N_6512,N_2716,N_3471);
nor U6513 (N_6513,N_4503,N_4096);
nor U6514 (N_6514,N_3447,N_3857);
nor U6515 (N_6515,N_2960,N_4057);
xor U6516 (N_6516,N_4106,N_3816);
xnor U6517 (N_6517,N_4522,N_3656);
and U6518 (N_6518,N_2953,N_3160);
xnor U6519 (N_6519,N_2551,N_3372);
xnor U6520 (N_6520,N_4204,N_3237);
nor U6521 (N_6521,N_4823,N_3491);
and U6522 (N_6522,N_3745,N_4394);
and U6523 (N_6523,N_3453,N_3986);
and U6524 (N_6524,N_4559,N_2672);
or U6525 (N_6525,N_3065,N_2741);
nand U6526 (N_6526,N_3024,N_3550);
and U6527 (N_6527,N_4948,N_3267);
or U6528 (N_6528,N_2653,N_3670);
nor U6529 (N_6529,N_2525,N_2715);
and U6530 (N_6530,N_3227,N_4835);
xnor U6531 (N_6531,N_2591,N_2997);
nand U6532 (N_6532,N_4129,N_3554);
or U6533 (N_6533,N_3791,N_3752);
xor U6534 (N_6534,N_4730,N_4166);
xnor U6535 (N_6535,N_3423,N_2766);
xnor U6536 (N_6536,N_2742,N_2654);
nor U6537 (N_6537,N_4219,N_3216);
nand U6538 (N_6538,N_3697,N_2771);
nor U6539 (N_6539,N_2764,N_3768);
nor U6540 (N_6540,N_3344,N_3123);
nor U6541 (N_6541,N_3233,N_4154);
or U6542 (N_6542,N_3181,N_4201);
nor U6543 (N_6543,N_2506,N_4979);
or U6544 (N_6544,N_4032,N_2531);
and U6545 (N_6545,N_4216,N_4943);
nand U6546 (N_6546,N_3295,N_3385);
and U6547 (N_6547,N_3756,N_3698);
nand U6548 (N_6548,N_2975,N_4456);
or U6549 (N_6549,N_3809,N_4357);
nor U6550 (N_6550,N_3654,N_3496);
and U6551 (N_6551,N_4042,N_3301);
xor U6552 (N_6552,N_3891,N_3667);
or U6553 (N_6553,N_3726,N_4066);
nand U6554 (N_6554,N_4998,N_3711);
and U6555 (N_6555,N_3619,N_2568);
nor U6556 (N_6556,N_3386,N_3052);
and U6557 (N_6557,N_2559,N_4690);
nor U6558 (N_6558,N_3876,N_4308);
nor U6559 (N_6559,N_3974,N_4131);
nand U6560 (N_6560,N_4500,N_2778);
and U6561 (N_6561,N_2735,N_4325);
nor U6562 (N_6562,N_4925,N_3294);
nand U6563 (N_6563,N_4346,N_4261);
xnor U6564 (N_6564,N_3753,N_3046);
xor U6565 (N_6565,N_3920,N_2746);
nor U6566 (N_6566,N_2566,N_4708);
nand U6567 (N_6567,N_2595,N_4794);
nor U6568 (N_6568,N_3329,N_4716);
and U6569 (N_6569,N_4795,N_3996);
xnor U6570 (N_6570,N_3185,N_3074);
nand U6571 (N_6571,N_3619,N_2588);
or U6572 (N_6572,N_3666,N_3271);
nor U6573 (N_6573,N_3892,N_3599);
nand U6574 (N_6574,N_3663,N_3881);
or U6575 (N_6575,N_4558,N_3941);
and U6576 (N_6576,N_2975,N_3513);
or U6577 (N_6577,N_2834,N_4011);
or U6578 (N_6578,N_4191,N_3982);
xor U6579 (N_6579,N_3753,N_3491);
or U6580 (N_6580,N_3302,N_3628);
or U6581 (N_6581,N_4015,N_3428);
nand U6582 (N_6582,N_3793,N_2753);
or U6583 (N_6583,N_3816,N_4374);
xnor U6584 (N_6584,N_4677,N_2983);
xor U6585 (N_6585,N_3934,N_4317);
xnor U6586 (N_6586,N_2878,N_2705);
nand U6587 (N_6587,N_2684,N_4033);
nand U6588 (N_6588,N_2810,N_4874);
and U6589 (N_6589,N_4462,N_2675);
and U6590 (N_6590,N_3743,N_4901);
nor U6591 (N_6591,N_3378,N_4406);
nor U6592 (N_6592,N_3781,N_2931);
or U6593 (N_6593,N_2558,N_4665);
nor U6594 (N_6594,N_3006,N_4301);
nand U6595 (N_6595,N_4076,N_3184);
and U6596 (N_6596,N_3109,N_2723);
nor U6597 (N_6597,N_4222,N_3474);
and U6598 (N_6598,N_3472,N_4829);
nand U6599 (N_6599,N_4401,N_2923);
or U6600 (N_6600,N_4367,N_4599);
nor U6601 (N_6601,N_2811,N_4555);
and U6602 (N_6602,N_4492,N_2577);
or U6603 (N_6603,N_3201,N_4492);
nand U6604 (N_6604,N_4754,N_4938);
and U6605 (N_6605,N_4868,N_3632);
xor U6606 (N_6606,N_3163,N_2914);
nor U6607 (N_6607,N_4837,N_3095);
nand U6608 (N_6608,N_4455,N_3622);
or U6609 (N_6609,N_2914,N_2717);
and U6610 (N_6610,N_2522,N_2859);
nor U6611 (N_6611,N_4988,N_4663);
xnor U6612 (N_6612,N_3318,N_4508);
xnor U6613 (N_6613,N_3752,N_4866);
and U6614 (N_6614,N_3009,N_3779);
nor U6615 (N_6615,N_3832,N_3723);
nor U6616 (N_6616,N_2787,N_3665);
nor U6617 (N_6617,N_3154,N_4088);
or U6618 (N_6618,N_4869,N_3495);
xor U6619 (N_6619,N_3386,N_4371);
and U6620 (N_6620,N_4806,N_3932);
and U6621 (N_6621,N_4299,N_2814);
nand U6622 (N_6622,N_3413,N_4536);
xor U6623 (N_6623,N_4003,N_4425);
nand U6624 (N_6624,N_2708,N_3382);
or U6625 (N_6625,N_3715,N_4578);
nand U6626 (N_6626,N_4372,N_4812);
nand U6627 (N_6627,N_3548,N_2711);
or U6628 (N_6628,N_4648,N_3398);
nor U6629 (N_6629,N_4445,N_3272);
nand U6630 (N_6630,N_2703,N_3835);
nand U6631 (N_6631,N_4835,N_2910);
nor U6632 (N_6632,N_3664,N_4332);
nor U6633 (N_6633,N_4182,N_4485);
xor U6634 (N_6634,N_3541,N_4778);
and U6635 (N_6635,N_3358,N_3857);
nor U6636 (N_6636,N_3578,N_2673);
and U6637 (N_6637,N_4114,N_3164);
xnor U6638 (N_6638,N_3159,N_2690);
and U6639 (N_6639,N_3095,N_4434);
or U6640 (N_6640,N_4371,N_4435);
and U6641 (N_6641,N_3459,N_3412);
nor U6642 (N_6642,N_4807,N_3009);
xor U6643 (N_6643,N_4600,N_4760);
nand U6644 (N_6644,N_3691,N_2823);
nand U6645 (N_6645,N_4219,N_2527);
nand U6646 (N_6646,N_2943,N_4656);
xnor U6647 (N_6647,N_3339,N_2574);
or U6648 (N_6648,N_3340,N_3803);
xor U6649 (N_6649,N_4994,N_3196);
and U6650 (N_6650,N_2697,N_3227);
and U6651 (N_6651,N_4445,N_4011);
nand U6652 (N_6652,N_2767,N_2718);
nor U6653 (N_6653,N_3647,N_2656);
nand U6654 (N_6654,N_4297,N_4412);
xnor U6655 (N_6655,N_3601,N_2590);
nand U6656 (N_6656,N_4124,N_3599);
nor U6657 (N_6657,N_3502,N_4536);
nand U6658 (N_6658,N_3343,N_3649);
and U6659 (N_6659,N_4387,N_3901);
nand U6660 (N_6660,N_4862,N_4306);
nand U6661 (N_6661,N_2686,N_3426);
nor U6662 (N_6662,N_3376,N_3110);
xor U6663 (N_6663,N_2988,N_4220);
or U6664 (N_6664,N_3587,N_4486);
xnor U6665 (N_6665,N_2905,N_3410);
nand U6666 (N_6666,N_3089,N_4610);
xnor U6667 (N_6667,N_3595,N_4669);
and U6668 (N_6668,N_3006,N_4844);
nand U6669 (N_6669,N_3176,N_3650);
and U6670 (N_6670,N_4744,N_3273);
xor U6671 (N_6671,N_3154,N_4338);
or U6672 (N_6672,N_3746,N_2735);
nor U6673 (N_6673,N_3018,N_3005);
nor U6674 (N_6674,N_3081,N_3777);
nor U6675 (N_6675,N_4160,N_4476);
and U6676 (N_6676,N_3139,N_3789);
or U6677 (N_6677,N_3970,N_4249);
and U6678 (N_6678,N_3651,N_2992);
or U6679 (N_6679,N_4659,N_4205);
nand U6680 (N_6680,N_4104,N_2877);
xnor U6681 (N_6681,N_3441,N_3499);
or U6682 (N_6682,N_3747,N_4093);
and U6683 (N_6683,N_4382,N_4712);
nor U6684 (N_6684,N_4569,N_2670);
and U6685 (N_6685,N_4325,N_2836);
nor U6686 (N_6686,N_3773,N_2861);
nand U6687 (N_6687,N_4661,N_3809);
or U6688 (N_6688,N_4290,N_3402);
and U6689 (N_6689,N_3255,N_4214);
or U6690 (N_6690,N_3097,N_2994);
nand U6691 (N_6691,N_2989,N_4746);
or U6692 (N_6692,N_2585,N_3731);
nand U6693 (N_6693,N_3599,N_3718);
and U6694 (N_6694,N_4844,N_3504);
nor U6695 (N_6695,N_3422,N_4892);
nand U6696 (N_6696,N_3714,N_2755);
xnor U6697 (N_6697,N_3219,N_3725);
and U6698 (N_6698,N_3593,N_3834);
or U6699 (N_6699,N_4594,N_3011);
nor U6700 (N_6700,N_3025,N_3355);
and U6701 (N_6701,N_4450,N_4266);
nand U6702 (N_6702,N_4513,N_3153);
xnor U6703 (N_6703,N_3290,N_3930);
nor U6704 (N_6704,N_4073,N_4776);
and U6705 (N_6705,N_3554,N_3400);
and U6706 (N_6706,N_2952,N_3402);
and U6707 (N_6707,N_4166,N_3228);
and U6708 (N_6708,N_3093,N_4155);
nor U6709 (N_6709,N_3287,N_3193);
nor U6710 (N_6710,N_3572,N_4498);
xnor U6711 (N_6711,N_3246,N_3623);
nand U6712 (N_6712,N_4739,N_3807);
xor U6713 (N_6713,N_4397,N_2583);
xor U6714 (N_6714,N_3725,N_4958);
and U6715 (N_6715,N_4193,N_3295);
and U6716 (N_6716,N_4014,N_4377);
and U6717 (N_6717,N_4590,N_2854);
or U6718 (N_6718,N_3226,N_3653);
or U6719 (N_6719,N_2772,N_3902);
xor U6720 (N_6720,N_4575,N_2983);
or U6721 (N_6721,N_4760,N_2997);
or U6722 (N_6722,N_3816,N_4237);
and U6723 (N_6723,N_2708,N_3944);
xor U6724 (N_6724,N_4505,N_3397);
and U6725 (N_6725,N_4022,N_2816);
xor U6726 (N_6726,N_4409,N_2742);
nand U6727 (N_6727,N_4892,N_3525);
nand U6728 (N_6728,N_2599,N_4124);
xnor U6729 (N_6729,N_2559,N_2797);
nand U6730 (N_6730,N_4710,N_4664);
and U6731 (N_6731,N_2710,N_4646);
xnor U6732 (N_6732,N_4706,N_2739);
nor U6733 (N_6733,N_4400,N_3462);
xnor U6734 (N_6734,N_4292,N_3493);
or U6735 (N_6735,N_4232,N_3227);
nor U6736 (N_6736,N_2556,N_3015);
xnor U6737 (N_6737,N_4141,N_4687);
or U6738 (N_6738,N_3147,N_4817);
xnor U6739 (N_6739,N_3073,N_2615);
nor U6740 (N_6740,N_3727,N_3947);
or U6741 (N_6741,N_3396,N_3169);
or U6742 (N_6742,N_4764,N_4536);
xor U6743 (N_6743,N_4802,N_4698);
or U6744 (N_6744,N_3140,N_4759);
and U6745 (N_6745,N_4050,N_3234);
nor U6746 (N_6746,N_4803,N_2635);
nand U6747 (N_6747,N_3239,N_2686);
or U6748 (N_6748,N_4335,N_2548);
nor U6749 (N_6749,N_4616,N_3798);
or U6750 (N_6750,N_4267,N_3825);
and U6751 (N_6751,N_4336,N_4904);
xnor U6752 (N_6752,N_3221,N_2664);
nand U6753 (N_6753,N_4919,N_4921);
nor U6754 (N_6754,N_4459,N_2743);
and U6755 (N_6755,N_3027,N_3204);
nand U6756 (N_6756,N_3646,N_2777);
xor U6757 (N_6757,N_4119,N_4681);
nor U6758 (N_6758,N_4304,N_4303);
nand U6759 (N_6759,N_2593,N_4073);
or U6760 (N_6760,N_4010,N_3040);
nor U6761 (N_6761,N_4561,N_4355);
and U6762 (N_6762,N_3431,N_4588);
and U6763 (N_6763,N_4647,N_4941);
nand U6764 (N_6764,N_4788,N_3320);
nand U6765 (N_6765,N_4886,N_2632);
or U6766 (N_6766,N_3048,N_4782);
or U6767 (N_6767,N_2978,N_3889);
or U6768 (N_6768,N_3056,N_4673);
nand U6769 (N_6769,N_3265,N_2525);
or U6770 (N_6770,N_4876,N_3182);
xnor U6771 (N_6771,N_2500,N_3166);
nor U6772 (N_6772,N_3023,N_3336);
nor U6773 (N_6773,N_2585,N_4932);
and U6774 (N_6774,N_4279,N_4064);
nand U6775 (N_6775,N_3805,N_4293);
or U6776 (N_6776,N_4893,N_3589);
xor U6777 (N_6777,N_4164,N_4634);
or U6778 (N_6778,N_4068,N_2695);
nand U6779 (N_6779,N_4642,N_3279);
xor U6780 (N_6780,N_4915,N_4965);
or U6781 (N_6781,N_4870,N_3046);
nor U6782 (N_6782,N_4164,N_3441);
nor U6783 (N_6783,N_2675,N_4498);
nor U6784 (N_6784,N_2966,N_4972);
or U6785 (N_6785,N_2849,N_3875);
nand U6786 (N_6786,N_2876,N_3989);
nand U6787 (N_6787,N_4386,N_4760);
nand U6788 (N_6788,N_4841,N_2737);
nand U6789 (N_6789,N_4918,N_2807);
nor U6790 (N_6790,N_4132,N_4443);
xnor U6791 (N_6791,N_4531,N_4513);
xor U6792 (N_6792,N_3013,N_3248);
xor U6793 (N_6793,N_4981,N_2807);
nor U6794 (N_6794,N_4357,N_2640);
xor U6795 (N_6795,N_3119,N_3700);
or U6796 (N_6796,N_2581,N_3934);
nor U6797 (N_6797,N_4291,N_2631);
xor U6798 (N_6798,N_3340,N_4681);
and U6799 (N_6799,N_3610,N_3651);
or U6800 (N_6800,N_3133,N_4592);
nand U6801 (N_6801,N_4977,N_4562);
or U6802 (N_6802,N_4979,N_4494);
xor U6803 (N_6803,N_2636,N_3137);
nor U6804 (N_6804,N_2520,N_4887);
nand U6805 (N_6805,N_4547,N_4205);
xor U6806 (N_6806,N_3662,N_4412);
xnor U6807 (N_6807,N_2794,N_4695);
or U6808 (N_6808,N_3874,N_4828);
or U6809 (N_6809,N_2872,N_3523);
nor U6810 (N_6810,N_3938,N_3960);
xnor U6811 (N_6811,N_2989,N_4712);
nand U6812 (N_6812,N_4544,N_4716);
nand U6813 (N_6813,N_4062,N_2742);
and U6814 (N_6814,N_4308,N_4882);
and U6815 (N_6815,N_3017,N_4527);
nor U6816 (N_6816,N_4100,N_4249);
xnor U6817 (N_6817,N_3328,N_3342);
xor U6818 (N_6818,N_3903,N_2680);
xnor U6819 (N_6819,N_3502,N_3046);
nor U6820 (N_6820,N_4562,N_3693);
or U6821 (N_6821,N_4573,N_3353);
or U6822 (N_6822,N_3055,N_4660);
and U6823 (N_6823,N_4138,N_3274);
and U6824 (N_6824,N_3406,N_4172);
nand U6825 (N_6825,N_3116,N_2885);
and U6826 (N_6826,N_4350,N_4256);
nand U6827 (N_6827,N_3385,N_3428);
xnor U6828 (N_6828,N_3953,N_3577);
and U6829 (N_6829,N_2717,N_3066);
and U6830 (N_6830,N_2748,N_3090);
xor U6831 (N_6831,N_2687,N_4364);
or U6832 (N_6832,N_3357,N_4210);
or U6833 (N_6833,N_3147,N_3274);
nor U6834 (N_6834,N_3798,N_3012);
and U6835 (N_6835,N_4117,N_3120);
and U6836 (N_6836,N_3055,N_3227);
and U6837 (N_6837,N_3709,N_4439);
or U6838 (N_6838,N_2911,N_4201);
nand U6839 (N_6839,N_3091,N_2655);
and U6840 (N_6840,N_4327,N_3779);
nand U6841 (N_6841,N_4455,N_4292);
or U6842 (N_6842,N_2607,N_3316);
nor U6843 (N_6843,N_2988,N_3181);
nor U6844 (N_6844,N_4693,N_3666);
and U6845 (N_6845,N_3144,N_2986);
nand U6846 (N_6846,N_2935,N_4640);
nand U6847 (N_6847,N_3677,N_3648);
nor U6848 (N_6848,N_3665,N_4490);
nand U6849 (N_6849,N_3763,N_2555);
or U6850 (N_6850,N_2658,N_2539);
nor U6851 (N_6851,N_3114,N_3566);
nand U6852 (N_6852,N_3056,N_3465);
or U6853 (N_6853,N_3717,N_4113);
xor U6854 (N_6854,N_2591,N_4447);
or U6855 (N_6855,N_4454,N_3266);
nor U6856 (N_6856,N_2519,N_4539);
or U6857 (N_6857,N_2981,N_3513);
or U6858 (N_6858,N_3427,N_3880);
or U6859 (N_6859,N_4015,N_4621);
and U6860 (N_6860,N_2962,N_4394);
or U6861 (N_6861,N_3932,N_4943);
and U6862 (N_6862,N_4487,N_4027);
nor U6863 (N_6863,N_4234,N_3960);
and U6864 (N_6864,N_4369,N_4755);
nor U6865 (N_6865,N_4953,N_4291);
xnor U6866 (N_6866,N_3369,N_3249);
and U6867 (N_6867,N_3265,N_3146);
or U6868 (N_6868,N_3667,N_4026);
nor U6869 (N_6869,N_4761,N_3892);
or U6870 (N_6870,N_3892,N_2776);
xnor U6871 (N_6871,N_4271,N_3020);
nand U6872 (N_6872,N_3612,N_4746);
xor U6873 (N_6873,N_2998,N_4338);
and U6874 (N_6874,N_4498,N_2708);
nor U6875 (N_6875,N_4350,N_4778);
xnor U6876 (N_6876,N_4770,N_4328);
nand U6877 (N_6877,N_3144,N_3097);
nand U6878 (N_6878,N_3528,N_4612);
or U6879 (N_6879,N_3897,N_3239);
and U6880 (N_6880,N_3500,N_4623);
and U6881 (N_6881,N_3619,N_4199);
and U6882 (N_6882,N_2649,N_4670);
xnor U6883 (N_6883,N_3122,N_3877);
and U6884 (N_6884,N_4850,N_3811);
xnor U6885 (N_6885,N_4429,N_2854);
nand U6886 (N_6886,N_4625,N_3714);
xor U6887 (N_6887,N_3545,N_2999);
and U6888 (N_6888,N_4122,N_2751);
xnor U6889 (N_6889,N_3905,N_4407);
xor U6890 (N_6890,N_3648,N_2611);
nand U6891 (N_6891,N_2521,N_2784);
and U6892 (N_6892,N_4610,N_4605);
and U6893 (N_6893,N_3094,N_3156);
and U6894 (N_6894,N_4969,N_4381);
or U6895 (N_6895,N_3019,N_3376);
nand U6896 (N_6896,N_2952,N_3206);
xnor U6897 (N_6897,N_4828,N_4139);
or U6898 (N_6898,N_4165,N_4588);
xor U6899 (N_6899,N_3247,N_4911);
xor U6900 (N_6900,N_3840,N_3371);
xnor U6901 (N_6901,N_3171,N_4550);
or U6902 (N_6902,N_3747,N_4237);
xnor U6903 (N_6903,N_3082,N_3938);
xnor U6904 (N_6904,N_3980,N_4530);
and U6905 (N_6905,N_3351,N_3068);
nor U6906 (N_6906,N_2655,N_4823);
nor U6907 (N_6907,N_3064,N_4703);
or U6908 (N_6908,N_2643,N_4375);
xnor U6909 (N_6909,N_3078,N_4521);
or U6910 (N_6910,N_4564,N_4663);
or U6911 (N_6911,N_3523,N_3472);
and U6912 (N_6912,N_3505,N_3796);
nor U6913 (N_6913,N_4809,N_2723);
nand U6914 (N_6914,N_2997,N_2517);
nand U6915 (N_6915,N_3829,N_3448);
xnor U6916 (N_6916,N_4861,N_4926);
xor U6917 (N_6917,N_3218,N_3842);
and U6918 (N_6918,N_3768,N_4137);
or U6919 (N_6919,N_2844,N_3664);
and U6920 (N_6920,N_2894,N_3924);
xor U6921 (N_6921,N_3917,N_4161);
or U6922 (N_6922,N_3049,N_2886);
and U6923 (N_6923,N_4982,N_4769);
and U6924 (N_6924,N_2767,N_3835);
xnor U6925 (N_6925,N_3473,N_2635);
nor U6926 (N_6926,N_4719,N_4516);
xnor U6927 (N_6927,N_4371,N_3134);
xnor U6928 (N_6928,N_4129,N_3898);
nand U6929 (N_6929,N_3753,N_4771);
or U6930 (N_6930,N_4905,N_4111);
nor U6931 (N_6931,N_4007,N_2666);
xnor U6932 (N_6932,N_4188,N_4541);
and U6933 (N_6933,N_3603,N_4449);
xnor U6934 (N_6934,N_4999,N_4663);
and U6935 (N_6935,N_3288,N_3032);
nor U6936 (N_6936,N_3553,N_2670);
nor U6937 (N_6937,N_4548,N_3056);
nor U6938 (N_6938,N_3279,N_3569);
nand U6939 (N_6939,N_4604,N_2856);
and U6940 (N_6940,N_3707,N_4033);
or U6941 (N_6941,N_2990,N_3879);
and U6942 (N_6942,N_2574,N_3367);
or U6943 (N_6943,N_3349,N_4775);
or U6944 (N_6944,N_3769,N_4347);
or U6945 (N_6945,N_3936,N_2947);
nand U6946 (N_6946,N_3846,N_3278);
nor U6947 (N_6947,N_2867,N_3737);
nor U6948 (N_6948,N_3378,N_2669);
or U6949 (N_6949,N_4127,N_3799);
nand U6950 (N_6950,N_3594,N_3325);
nand U6951 (N_6951,N_4853,N_3779);
nand U6952 (N_6952,N_3832,N_2858);
or U6953 (N_6953,N_2593,N_3706);
xnor U6954 (N_6954,N_2994,N_4812);
xor U6955 (N_6955,N_3503,N_4591);
nand U6956 (N_6956,N_4975,N_2604);
nor U6957 (N_6957,N_4848,N_3940);
nor U6958 (N_6958,N_3164,N_4383);
and U6959 (N_6959,N_4905,N_4913);
xor U6960 (N_6960,N_3038,N_4820);
nor U6961 (N_6961,N_3032,N_2730);
or U6962 (N_6962,N_4025,N_2673);
nand U6963 (N_6963,N_3395,N_3186);
or U6964 (N_6964,N_4404,N_2731);
and U6965 (N_6965,N_3113,N_2919);
nor U6966 (N_6966,N_4602,N_2728);
nand U6967 (N_6967,N_4100,N_3822);
nor U6968 (N_6968,N_4744,N_4684);
xnor U6969 (N_6969,N_3451,N_4170);
xnor U6970 (N_6970,N_4551,N_3132);
nor U6971 (N_6971,N_3767,N_3858);
and U6972 (N_6972,N_2654,N_3350);
and U6973 (N_6973,N_3193,N_3192);
nand U6974 (N_6974,N_4753,N_2919);
and U6975 (N_6975,N_4741,N_4695);
nand U6976 (N_6976,N_3459,N_4141);
xor U6977 (N_6977,N_4848,N_4553);
nand U6978 (N_6978,N_4581,N_3250);
or U6979 (N_6979,N_4185,N_4670);
or U6980 (N_6980,N_3435,N_4976);
xnor U6981 (N_6981,N_4580,N_3953);
and U6982 (N_6982,N_4329,N_2904);
nand U6983 (N_6983,N_4177,N_4767);
nand U6984 (N_6984,N_4521,N_3952);
nor U6985 (N_6985,N_3838,N_4779);
nor U6986 (N_6986,N_4404,N_3116);
xnor U6987 (N_6987,N_4559,N_3381);
nor U6988 (N_6988,N_4823,N_2547);
xor U6989 (N_6989,N_4309,N_3135);
and U6990 (N_6990,N_3026,N_2582);
nor U6991 (N_6991,N_4792,N_4051);
nor U6992 (N_6992,N_2927,N_4437);
xor U6993 (N_6993,N_3245,N_3684);
nand U6994 (N_6994,N_3193,N_4996);
and U6995 (N_6995,N_2924,N_4883);
nand U6996 (N_6996,N_4275,N_4289);
nand U6997 (N_6997,N_4851,N_2778);
xnor U6998 (N_6998,N_4109,N_4177);
nor U6999 (N_6999,N_4817,N_3155);
xor U7000 (N_7000,N_2773,N_3361);
and U7001 (N_7001,N_2985,N_3044);
or U7002 (N_7002,N_4996,N_4181);
xor U7003 (N_7003,N_3058,N_3734);
or U7004 (N_7004,N_4678,N_2830);
nand U7005 (N_7005,N_4654,N_4990);
nor U7006 (N_7006,N_2772,N_3449);
and U7007 (N_7007,N_3274,N_4774);
and U7008 (N_7008,N_3207,N_4377);
xnor U7009 (N_7009,N_2613,N_3452);
nand U7010 (N_7010,N_3805,N_2631);
or U7011 (N_7011,N_2989,N_4735);
xor U7012 (N_7012,N_3407,N_2861);
nand U7013 (N_7013,N_3360,N_4792);
or U7014 (N_7014,N_2817,N_2972);
xor U7015 (N_7015,N_3608,N_4066);
nand U7016 (N_7016,N_3469,N_4973);
nor U7017 (N_7017,N_4296,N_2688);
nor U7018 (N_7018,N_3341,N_4829);
xor U7019 (N_7019,N_3578,N_2873);
and U7020 (N_7020,N_3872,N_3448);
or U7021 (N_7021,N_4611,N_3061);
nor U7022 (N_7022,N_4947,N_4642);
and U7023 (N_7023,N_4997,N_4400);
and U7024 (N_7024,N_2768,N_4170);
xor U7025 (N_7025,N_2779,N_4712);
xnor U7026 (N_7026,N_4904,N_4993);
and U7027 (N_7027,N_3181,N_3606);
nand U7028 (N_7028,N_2906,N_4821);
and U7029 (N_7029,N_2972,N_3755);
nand U7030 (N_7030,N_3553,N_2935);
nand U7031 (N_7031,N_4856,N_3900);
nand U7032 (N_7032,N_2715,N_4887);
and U7033 (N_7033,N_2859,N_4928);
nand U7034 (N_7034,N_3073,N_4903);
xnor U7035 (N_7035,N_3852,N_3451);
nor U7036 (N_7036,N_4722,N_4158);
xor U7037 (N_7037,N_2557,N_2641);
xnor U7038 (N_7038,N_2645,N_4871);
xor U7039 (N_7039,N_4128,N_4657);
or U7040 (N_7040,N_2894,N_3351);
and U7041 (N_7041,N_3454,N_4357);
and U7042 (N_7042,N_3671,N_4813);
or U7043 (N_7043,N_4419,N_2767);
and U7044 (N_7044,N_4774,N_3892);
or U7045 (N_7045,N_3655,N_3315);
or U7046 (N_7046,N_3091,N_4887);
nor U7047 (N_7047,N_3863,N_3196);
and U7048 (N_7048,N_2558,N_3062);
nand U7049 (N_7049,N_4497,N_4279);
nand U7050 (N_7050,N_3522,N_4026);
nand U7051 (N_7051,N_2545,N_4047);
nor U7052 (N_7052,N_4110,N_4485);
or U7053 (N_7053,N_2936,N_2552);
and U7054 (N_7054,N_3989,N_3088);
or U7055 (N_7055,N_4214,N_3299);
xor U7056 (N_7056,N_2689,N_4064);
nand U7057 (N_7057,N_3753,N_4673);
and U7058 (N_7058,N_4478,N_4098);
or U7059 (N_7059,N_2724,N_4977);
xor U7060 (N_7060,N_4133,N_3357);
xnor U7061 (N_7061,N_3961,N_3932);
nand U7062 (N_7062,N_3555,N_4772);
or U7063 (N_7063,N_2936,N_3321);
nor U7064 (N_7064,N_3354,N_2971);
nor U7065 (N_7065,N_4255,N_4894);
and U7066 (N_7066,N_4202,N_4478);
nor U7067 (N_7067,N_4528,N_4517);
xnor U7068 (N_7068,N_2803,N_4434);
or U7069 (N_7069,N_3067,N_4052);
nand U7070 (N_7070,N_4163,N_4096);
and U7071 (N_7071,N_4394,N_3656);
nor U7072 (N_7072,N_3562,N_3026);
and U7073 (N_7073,N_3954,N_3194);
nand U7074 (N_7074,N_2860,N_3078);
xnor U7075 (N_7075,N_4917,N_2694);
nor U7076 (N_7076,N_4631,N_4826);
xnor U7077 (N_7077,N_4138,N_3041);
and U7078 (N_7078,N_2514,N_3622);
and U7079 (N_7079,N_2957,N_3848);
nor U7080 (N_7080,N_3003,N_4505);
and U7081 (N_7081,N_4554,N_4220);
and U7082 (N_7082,N_2730,N_2589);
and U7083 (N_7083,N_2512,N_2712);
or U7084 (N_7084,N_3103,N_4840);
nand U7085 (N_7085,N_4016,N_4220);
nor U7086 (N_7086,N_3542,N_4236);
or U7087 (N_7087,N_3702,N_3179);
nand U7088 (N_7088,N_4730,N_4980);
xor U7089 (N_7089,N_3930,N_4997);
nor U7090 (N_7090,N_3862,N_4562);
and U7091 (N_7091,N_3278,N_4131);
xnor U7092 (N_7092,N_3342,N_3432);
and U7093 (N_7093,N_4225,N_3585);
or U7094 (N_7094,N_2658,N_3244);
and U7095 (N_7095,N_3483,N_2806);
nor U7096 (N_7096,N_4888,N_2630);
nand U7097 (N_7097,N_3819,N_3094);
xnor U7098 (N_7098,N_4853,N_4783);
or U7099 (N_7099,N_3320,N_3105);
xor U7100 (N_7100,N_2649,N_4321);
nor U7101 (N_7101,N_3943,N_4712);
or U7102 (N_7102,N_4647,N_3592);
nor U7103 (N_7103,N_4286,N_3908);
or U7104 (N_7104,N_3325,N_3562);
xor U7105 (N_7105,N_4110,N_4243);
xnor U7106 (N_7106,N_4492,N_4871);
or U7107 (N_7107,N_3834,N_3729);
xor U7108 (N_7108,N_4872,N_4747);
and U7109 (N_7109,N_2895,N_4594);
nor U7110 (N_7110,N_4894,N_3858);
and U7111 (N_7111,N_2665,N_3597);
xor U7112 (N_7112,N_3443,N_4718);
xor U7113 (N_7113,N_4380,N_3591);
nand U7114 (N_7114,N_3338,N_4595);
xnor U7115 (N_7115,N_3044,N_4449);
nor U7116 (N_7116,N_4208,N_3376);
and U7117 (N_7117,N_4569,N_4711);
nor U7118 (N_7118,N_4681,N_4478);
xnor U7119 (N_7119,N_2994,N_4749);
or U7120 (N_7120,N_2714,N_2832);
nor U7121 (N_7121,N_4622,N_4844);
or U7122 (N_7122,N_4861,N_2921);
or U7123 (N_7123,N_3401,N_3996);
or U7124 (N_7124,N_4834,N_4707);
nor U7125 (N_7125,N_2865,N_4880);
xor U7126 (N_7126,N_4283,N_2645);
nor U7127 (N_7127,N_3522,N_3261);
or U7128 (N_7128,N_4696,N_3469);
nor U7129 (N_7129,N_4581,N_4696);
nor U7130 (N_7130,N_2813,N_3483);
nor U7131 (N_7131,N_2684,N_3414);
xnor U7132 (N_7132,N_2529,N_3817);
nand U7133 (N_7133,N_4939,N_4970);
and U7134 (N_7134,N_3279,N_4584);
xnor U7135 (N_7135,N_3863,N_2684);
or U7136 (N_7136,N_2684,N_4135);
and U7137 (N_7137,N_2699,N_3085);
xnor U7138 (N_7138,N_4927,N_2579);
or U7139 (N_7139,N_3041,N_3690);
and U7140 (N_7140,N_3425,N_3552);
nor U7141 (N_7141,N_4418,N_4507);
xor U7142 (N_7142,N_4583,N_2953);
or U7143 (N_7143,N_4596,N_4631);
and U7144 (N_7144,N_4405,N_4507);
and U7145 (N_7145,N_4797,N_4339);
and U7146 (N_7146,N_2876,N_2790);
xnor U7147 (N_7147,N_3906,N_3602);
nor U7148 (N_7148,N_4851,N_3619);
xnor U7149 (N_7149,N_2652,N_3996);
or U7150 (N_7150,N_2861,N_2843);
or U7151 (N_7151,N_2545,N_4667);
and U7152 (N_7152,N_4979,N_3089);
xnor U7153 (N_7153,N_3132,N_2873);
nand U7154 (N_7154,N_2623,N_4178);
or U7155 (N_7155,N_2965,N_3814);
and U7156 (N_7156,N_3933,N_4093);
or U7157 (N_7157,N_4729,N_4404);
xor U7158 (N_7158,N_4112,N_3399);
nor U7159 (N_7159,N_2704,N_3093);
and U7160 (N_7160,N_3639,N_3339);
nor U7161 (N_7161,N_3452,N_4536);
or U7162 (N_7162,N_3631,N_2651);
and U7163 (N_7163,N_4239,N_4734);
xor U7164 (N_7164,N_4271,N_4259);
or U7165 (N_7165,N_4340,N_2990);
xnor U7166 (N_7166,N_2676,N_4288);
nor U7167 (N_7167,N_3255,N_2933);
nor U7168 (N_7168,N_3401,N_3416);
xnor U7169 (N_7169,N_3363,N_4534);
nor U7170 (N_7170,N_4197,N_4299);
or U7171 (N_7171,N_3897,N_4023);
and U7172 (N_7172,N_2585,N_3103);
nor U7173 (N_7173,N_4663,N_3651);
nor U7174 (N_7174,N_4893,N_3718);
nor U7175 (N_7175,N_2519,N_2734);
nand U7176 (N_7176,N_4432,N_3780);
nor U7177 (N_7177,N_2920,N_3180);
xor U7178 (N_7178,N_4247,N_4515);
xnor U7179 (N_7179,N_3662,N_4262);
xor U7180 (N_7180,N_3543,N_2888);
xor U7181 (N_7181,N_3151,N_2596);
nand U7182 (N_7182,N_4646,N_2750);
and U7183 (N_7183,N_3927,N_4445);
and U7184 (N_7184,N_3680,N_4634);
nor U7185 (N_7185,N_4425,N_2832);
or U7186 (N_7186,N_2935,N_3858);
xnor U7187 (N_7187,N_3722,N_4126);
and U7188 (N_7188,N_4408,N_3531);
nand U7189 (N_7189,N_3604,N_4171);
or U7190 (N_7190,N_2542,N_3134);
nand U7191 (N_7191,N_4527,N_4217);
or U7192 (N_7192,N_2772,N_3189);
or U7193 (N_7193,N_4062,N_4848);
or U7194 (N_7194,N_4539,N_4477);
and U7195 (N_7195,N_4238,N_4677);
nand U7196 (N_7196,N_3428,N_4309);
and U7197 (N_7197,N_3284,N_3813);
xnor U7198 (N_7198,N_2621,N_3736);
and U7199 (N_7199,N_4779,N_4673);
xor U7200 (N_7200,N_4406,N_3079);
nor U7201 (N_7201,N_2934,N_3070);
nand U7202 (N_7202,N_4065,N_3083);
nor U7203 (N_7203,N_4613,N_2872);
xor U7204 (N_7204,N_4803,N_4454);
xor U7205 (N_7205,N_3612,N_3117);
and U7206 (N_7206,N_4983,N_3099);
or U7207 (N_7207,N_3923,N_3597);
and U7208 (N_7208,N_3250,N_3525);
nor U7209 (N_7209,N_4275,N_3313);
nand U7210 (N_7210,N_2603,N_2605);
or U7211 (N_7211,N_4739,N_3268);
nand U7212 (N_7212,N_4695,N_4943);
xnor U7213 (N_7213,N_4641,N_4216);
xor U7214 (N_7214,N_4801,N_4944);
nor U7215 (N_7215,N_3184,N_2657);
nor U7216 (N_7216,N_3033,N_4058);
xor U7217 (N_7217,N_3739,N_2640);
xor U7218 (N_7218,N_4955,N_3848);
nand U7219 (N_7219,N_3459,N_4717);
nor U7220 (N_7220,N_4611,N_3087);
and U7221 (N_7221,N_4485,N_4256);
xnor U7222 (N_7222,N_4058,N_4584);
nand U7223 (N_7223,N_4844,N_4280);
nand U7224 (N_7224,N_2556,N_3027);
nor U7225 (N_7225,N_3651,N_2903);
nor U7226 (N_7226,N_3539,N_2675);
or U7227 (N_7227,N_4189,N_3813);
nand U7228 (N_7228,N_2834,N_3809);
and U7229 (N_7229,N_4398,N_3023);
nand U7230 (N_7230,N_3976,N_3682);
xor U7231 (N_7231,N_3963,N_3885);
xor U7232 (N_7232,N_4083,N_4489);
nand U7233 (N_7233,N_3973,N_3989);
or U7234 (N_7234,N_4497,N_2645);
nor U7235 (N_7235,N_4728,N_4082);
and U7236 (N_7236,N_3772,N_4423);
xor U7237 (N_7237,N_2885,N_3369);
nand U7238 (N_7238,N_3244,N_3047);
nor U7239 (N_7239,N_2775,N_3456);
or U7240 (N_7240,N_4626,N_2835);
xnor U7241 (N_7241,N_4814,N_4150);
nand U7242 (N_7242,N_3287,N_4399);
nand U7243 (N_7243,N_3008,N_4141);
nor U7244 (N_7244,N_3718,N_4162);
nor U7245 (N_7245,N_4447,N_3413);
and U7246 (N_7246,N_2620,N_4512);
and U7247 (N_7247,N_4631,N_3642);
xnor U7248 (N_7248,N_3297,N_3284);
xor U7249 (N_7249,N_4039,N_3915);
xor U7250 (N_7250,N_4839,N_4194);
nor U7251 (N_7251,N_3639,N_4234);
xnor U7252 (N_7252,N_3202,N_3421);
xor U7253 (N_7253,N_2881,N_4779);
xnor U7254 (N_7254,N_3310,N_3073);
or U7255 (N_7255,N_2659,N_4379);
nand U7256 (N_7256,N_3314,N_4056);
nor U7257 (N_7257,N_3869,N_4310);
nor U7258 (N_7258,N_4141,N_4981);
and U7259 (N_7259,N_4751,N_3832);
or U7260 (N_7260,N_4287,N_3152);
and U7261 (N_7261,N_3331,N_3545);
nor U7262 (N_7262,N_3838,N_2843);
nand U7263 (N_7263,N_3550,N_4544);
nand U7264 (N_7264,N_3960,N_3868);
nand U7265 (N_7265,N_3518,N_4457);
nand U7266 (N_7266,N_4012,N_2673);
nor U7267 (N_7267,N_4703,N_3435);
or U7268 (N_7268,N_2507,N_4873);
xor U7269 (N_7269,N_4776,N_2610);
and U7270 (N_7270,N_4922,N_4973);
and U7271 (N_7271,N_3086,N_3969);
or U7272 (N_7272,N_3648,N_2693);
nand U7273 (N_7273,N_3879,N_3494);
or U7274 (N_7274,N_2637,N_4994);
and U7275 (N_7275,N_2945,N_3468);
nor U7276 (N_7276,N_4187,N_4877);
and U7277 (N_7277,N_4340,N_4003);
nand U7278 (N_7278,N_3087,N_3105);
nor U7279 (N_7279,N_2875,N_4227);
xor U7280 (N_7280,N_3780,N_3053);
nor U7281 (N_7281,N_3738,N_3843);
nand U7282 (N_7282,N_3076,N_3481);
nand U7283 (N_7283,N_4481,N_4999);
or U7284 (N_7284,N_4884,N_3155);
nor U7285 (N_7285,N_4763,N_4205);
nor U7286 (N_7286,N_4495,N_3649);
or U7287 (N_7287,N_2664,N_2647);
nor U7288 (N_7288,N_3963,N_4326);
or U7289 (N_7289,N_3993,N_4349);
xor U7290 (N_7290,N_3212,N_4605);
nand U7291 (N_7291,N_3076,N_3443);
and U7292 (N_7292,N_3437,N_4593);
and U7293 (N_7293,N_4313,N_2530);
xnor U7294 (N_7294,N_3666,N_3012);
or U7295 (N_7295,N_4310,N_2961);
or U7296 (N_7296,N_3994,N_4033);
and U7297 (N_7297,N_4465,N_2916);
nor U7298 (N_7298,N_4741,N_4465);
and U7299 (N_7299,N_3791,N_2911);
nor U7300 (N_7300,N_3147,N_4842);
and U7301 (N_7301,N_4113,N_3200);
xor U7302 (N_7302,N_4692,N_3134);
xor U7303 (N_7303,N_4332,N_2849);
xor U7304 (N_7304,N_4919,N_4856);
nand U7305 (N_7305,N_4741,N_4992);
or U7306 (N_7306,N_3226,N_4920);
or U7307 (N_7307,N_4712,N_4219);
xnor U7308 (N_7308,N_4743,N_2991);
nand U7309 (N_7309,N_3795,N_3277);
or U7310 (N_7310,N_2767,N_3409);
nand U7311 (N_7311,N_3701,N_2506);
or U7312 (N_7312,N_3280,N_3860);
and U7313 (N_7313,N_4018,N_3442);
or U7314 (N_7314,N_3942,N_4014);
nand U7315 (N_7315,N_3761,N_4469);
nand U7316 (N_7316,N_4550,N_4356);
and U7317 (N_7317,N_2781,N_3963);
or U7318 (N_7318,N_4815,N_3485);
xnor U7319 (N_7319,N_3331,N_2861);
nand U7320 (N_7320,N_3696,N_3389);
nand U7321 (N_7321,N_2670,N_4225);
nor U7322 (N_7322,N_4967,N_4070);
or U7323 (N_7323,N_3087,N_4614);
nand U7324 (N_7324,N_4386,N_4548);
and U7325 (N_7325,N_3798,N_3518);
nor U7326 (N_7326,N_3495,N_4883);
xor U7327 (N_7327,N_4423,N_4242);
nand U7328 (N_7328,N_4057,N_3476);
nor U7329 (N_7329,N_2511,N_4171);
or U7330 (N_7330,N_3793,N_4941);
and U7331 (N_7331,N_3285,N_2861);
or U7332 (N_7332,N_3216,N_3264);
and U7333 (N_7333,N_3685,N_4753);
nor U7334 (N_7334,N_3224,N_3560);
xor U7335 (N_7335,N_4703,N_3639);
or U7336 (N_7336,N_4679,N_4202);
and U7337 (N_7337,N_3119,N_3486);
nor U7338 (N_7338,N_4044,N_2910);
nor U7339 (N_7339,N_4712,N_4550);
or U7340 (N_7340,N_2803,N_4304);
and U7341 (N_7341,N_4827,N_3302);
xor U7342 (N_7342,N_2706,N_4923);
nor U7343 (N_7343,N_3279,N_4383);
xnor U7344 (N_7344,N_3344,N_3890);
xor U7345 (N_7345,N_3624,N_4485);
and U7346 (N_7346,N_2806,N_3033);
nand U7347 (N_7347,N_3186,N_4974);
nand U7348 (N_7348,N_4048,N_2791);
xor U7349 (N_7349,N_4548,N_4667);
nor U7350 (N_7350,N_2586,N_2734);
xnor U7351 (N_7351,N_2948,N_3941);
nor U7352 (N_7352,N_3046,N_4543);
nand U7353 (N_7353,N_3527,N_4672);
or U7354 (N_7354,N_3168,N_3628);
xnor U7355 (N_7355,N_3248,N_3141);
nand U7356 (N_7356,N_3166,N_4493);
nand U7357 (N_7357,N_4996,N_3379);
xor U7358 (N_7358,N_2652,N_2972);
and U7359 (N_7359,N_4347,N_3495);
nand U7360 (N_7360,N_4601,N_2645);
xnor U7361 (N_7361,N_4509,N_2853);
and U7362 (N_7362,N_4871,N_3984);
and U7363 (N_7363,N_4096,N_3606);
and U7364 (N_7364,N_4739,N_4277);
or U7365 (N_7365,N_3426,N_4875);
xnor U7366 (N_7366,N_2819,N_3107);
nand U7367 (N_7367,N_4274,N_4277);
and U7368 (N_7368,N_3957,N_3663);
xor U7369 (N_7369,N_4035,N_4474);
nor U7370 (N_7370,N_4999,N_3013);
xor U7371 (N_7371,N_4136,N_4265);
nand U7372 (N_7372,N_4740,N_3878);
or U7373 (N_7373,N_3950,N_4606);
xor U7374 (N_7374,N_4987,N_4185);
nand U7375 (N_7375,N_4866,N_2597);
nor U7376 (N_7376,N_2771,N_4881);
nand U7377 (N_7377,N_4692,N_3463);
or U7378 (N_7378,N_4469,N_4993);
and U7379 (N_7379,N_2918,N_3222);
nand U7380 (N_7380,N_3271,N_3601);
xor U7381 (N_7381,N_2623,N_4811);
nand U7382 (N_7382,N_2727,N_3119);
nand U7383 (N_7383,N_4230,N_4348);
nor U7384 (N_7384,N_2978,N_3990);
or U7385 (N_7385,N_4109,N_2587);
and U7386 (N_7386,N_3500,N_3566);
nor U7387 (N_7387,N_4347,N_2732);
nor U7388 (N_7388,N_4946,N_4865);
and U7389 (N_7389,N_4862,N_2849);
nor U7390 (N_7390,N_4525,N_3587);
and U7391 (N_7391,N_2591,N_4411);
nor U7392 (N_7392,N_2916,N_3020);
or U7393 (N_7393,N_4580,N_4285);
nor U7394 (N_7394,N_2854,N_4474);
nand U7395 (N_7395,N_4182,N_4949);
xnor U7396 (N_7396,N_4726,N_4188);
or U7397 (N_7397,N_3809,N_3759);
nand U7398 (N_7398,N_2919,N_3242);
xor U7399 (N_7399,N_3144,N_3745);
and U7400 (N_7400,N_4302,N_4692);
nand U7401 (N_7401,N_4911,N_4073);
and U7402 (N_7402,N_4762,N_2989);
nand U7403 (N_7403,N_3609,N_2808);
or U7404 (N_7404,N_3362,N_2564);
nor U7405 (N_7405,N_4385,N_4712);
nor U7406 (N_7406,N_3394,N_2507);
and U7407 (N_7407,N_2581,N_3654);
xor U7408 (N_7408,N_3120,N_2543);
nor U7409 (N_7409,N_4396,N_4281);
or U7410 (N_7410,N_2674,N_4206);
or U7411 (N_7411,N_4754,N_4592);
xor U7412 (N_7412,N_3911,N_3217);
or U7413 (N_7413,N_4334,N_2678);
and U7414 (N_7414,N_3893,N_4241);
and U7415 (N_7415,N_4086,N_3067);
or U7416 (N_7416,N_3193,N_3332);
nand U7417 (N_7417,N_2720,N_3358);
nand U7418 (N_7418,N_4277,N_3053);
nand U7419 (N_7419,N_4523,N_3702);
nor U7420 (N_7420,N_4550,N_2784);
nor U7421 (N_7421,N_2844,N_3402);
nand U7422 (N_7422,N_2619,N_4254);
xnor U7423 (N_7423,N_2581,N_2851);
or U7424 (N_7424,N_4505,N_3496);
or U7425 (N_7425,N_4094,N_2824);
and U7426 (N_7426,N_2889,N_4651);
or U7427 (N_7427,N_2595,N_4940);
nor U7428 (N_7428,N_2843,N_2797);
nand U7429 (N_7429,N_3172,N_3958);
or U7430 (N_7430,N_4610,N_3992);
nor U7431 (N_7431,N_4861,N_4460);
and U7432 (N_7432,N_4910,N_3848);
nand U7433 (N_7433,N_3548,N_3506);
xnor U7434 (N_7434,N_3976,N_3352);
or U7435 (N_7435,N_3718,N_3967);
xnor U7436 (N_7436,N_3818,N_4573);
xnor U7437 (N_7437,N_3738,N_3829);
nor U7438 (N_7438,N_4607,N_3944);
and U7439 (N_7439,N_3952,N_4335);
nand U7440 (N_7440,N_4073,N_4538);
xor U7441 (N_7441,N_2961,N_4891);
xor U7442 (N_7442,N_3648,N_3176);
nand U7443 (N_7443,N_3245,N_4762);
xnor U7444 (N_7444,N_4202,N_3469);
and U7445 (N_7445,N_4569,N_4894);
and U7446 (N_7446,N_4954,N_2959);
nor U7447 (N_7447,N_2752,N_4886);
and U7448 (N_7448,N_3527,N_3362);
xor U7449 (N_7449,N_4846,N_4922);
nand U7450 (N_7450,N_3628,N_4659);
nor U7451 (N_7451,N_4843,N_4950);
nand U7452 (N_7452,N_4077,N_3772);
xor U7453 (N_7453,N_2577,N_3668);
xor U7454 (N_7454,N_3582,N_4537);
or U7455 (N_7455,N_4807,N_2760);
or U7456 (N_7456,N_2806,N_4711);
or U7457 (N_7457,N_3321,N_3218);
or U7458 (N_7458,N_2571,N_2626);
nand U7459 (N_7459,N_3057,N_4587);
xnor U7460 (N_7460,N_2790,N_3940);
xor U7461 (N_7461,N_3728,N_4722);
nor U7462 (N_7462,N_2688,N_3625);
nor U7463 (N_7463,N_3026,N_4935);
or U7464 (N_7464,N_2510,N_4748);
and U7465 (N_7465,N_2710,N_2691);
nor U7466 (N_7466,N_4403,N_3887);
xor U7467 (N_7467,N_2647,N_4991);
and U7468 (N_7468,N_4209,N_3315);
nand U7469 (N_7469,N_3608,N_4511);
nor U7470 (N_7470,N_4211,N_3396);
nor U7471 (N_7471,N_3261,N_3909);
nor U7472 (N_7472,N_3348,N_2711);
xor U7473 (N_7473,N_3204,N_3215);
and U7474 (N_7474,N_3071,N_4330);
nor U7475 (N_7475,N_4016,N_4272);
nor U7476 (N_7476,N_2741,N_4508);
nand U7477 (N_7477,N_4367,N_3298);
and U7478 (N_7478,N_3164,N_4926);
nor U7479 (N_7479,N_3373,N_3113);
xnor U7480 (N_7480,N_4236,N_3420);
and U7481 (N_7481,N_2752,N_2965);
or U7482 (N_7482,N_4786,N_4824);
xnor U7483 (N_7483,N_4481,N_4985);
nor U7484 (N_7484,N_2598,N_2905);
nand U7485 (N_7485,N_4453,N_2769);
and U7486 (N_7486,N_4229,N_2555);
or U7487 (N_7487,N_4944,N_2691);
nand U7488 (N_7488,N_3693,N_3417);
and U7489 (N_7489,N_2937,N_3999);
and U7490 (N_7490,N_2704,N_3678);
and U7491 (N_7491,N_4422,N_3713);
xor U7492 (N_7492,N_3231,N_4691);
or U7493 (N_7493,N_4948,N_3114);
nor U7494 (N_7494,N_4580,N_4527);
nor U7495 (N_7495,N_2513,N_3508);
nor U7496 (N_7496,N_3165,N_4297);
nor U7497 (N_7497,N_2897,N_4725);
nor U7498 (N_7498,N_2987,N_4989);
xor U7499 (N_7499,N_3693,N_2693);
nor U7500 (N_7500,N_7327,N_5732);
xor U7501 (N_7501,N_6017,N_6091);
nor U7502 (N_7502,N_6198,N_7194);
and U7503 (N_7503,N_6263,N_5590);
nor U7504 (N_7504,N_5088,N_5481);
nor U7505 (N_7505,N_5875,N_5010);
nor U7506 (N_7506,N_7385,N_6480);
nor U7507 (N_7507,N_5025,N_5707);
nor U7508 (N_7508,N_5258,N_6462);
nand U7509 (N_7509,N_5505,N_6486);
nand U7510 (N_7510,N_5754,N_6718);
nand U7511 (N_7511,N_5457,N_7190);
xnor U7512 (N_7512,N_5578,N_6339);
xnor U7513 (N_7513,N_6770,N_5842);
nor U7514 (N_7514,N_7313,N_6870);
nand U7515 (N_7515,N_5735,N_6428);
nand U7516 (N_7516,N_6891,N_5397);
nand U7517 (N_7517,N_5325,N_7472);
or U7518 (N_7518,N_6020,N_6210);
nor U7519 (N_7519,N_5169,N_7391);
nand U7520 (N_7520,N_5129,N_6081);
nand U7521 (N_7521,N_6888,N_6244);
and U7522 (N_7522,N_7417,N_5133);
or U7523 (N_7523,N_7119,N_5761);
xnor U7524 (N_7524,N_7229,N_7309);
xnor U7525 (N_7525,N_6335,N_7478);
nor U7526 (N_7526,N_6687,N_7438);
and U7527 (N_7527,N_6556,N_5062);
nor U7528 (N_7528,N_7228,N_5790);
nor U7529 (N_7529,N_6952,N_5065);
or U7530 (N_7530,N_5806,N_5529);
and U7531 (N_7531,N_6893,N_5681);
nor U7532 (N_7532,N_6748,N_6076);
nor U7533 (N_7533,N_6588,N_6746);
xnor U7534 (N_7534,N_7328,N_5771);
nor U7535 (N_7535,N_5094,N_6761);
nor U7536 (N_7536,N_6875,N_6729);
xor U7537 (N_7537,N_5278,N_6752);
or U7538 (N_7538,N_6955,N_6125);
nor U7539 (N_7539,N_7428,N_5988);
or U7540 (N_7540,N_5112,N_7020);
nor U7541 (N_7541,N_7348,N_6540);
and U7542 (N_7542,N_5615,N_5952);
nor U7543 (N_7543,N_7463,N_6913);
xnor U7544 (N_7544,N_6485,N_6171);
nor U7545 (N_7545,N_5138,N_5955);
or U7546 (N_7546,N_7330,N_7186);
nand U7547 (N_7547,N_7234,N_5423);
or U7548 (N_7548,N_6211,N_6987);
xor U7549 (N_7549,N_6663,N_7097);
or U7550 (N_7550,N_7439,N_5912);
nand U7551 (N_7551,N_7296,N_6995);
nand U7552 (N_7552,N_6622,N_7344);
and U7553 (N_7553,N_5610,N_6242);
or U7554 (N_7554,N_6157,N_6307);
nand U7555 (N_7555,N_7487,N_6253);
or U7556 (N_7556,N_6403,N_5555);
or U7557 (N_7557,N_5731,N_5626);
xor U7558 (N_7558,N_5388,N_5204);
nand U7559 (N_7559,N_5897,N_5880);
nor U7560 (N_7560,N_5121,N_6438);
nor U7561 (N_7561,N_5437,N_6484);
nand U7562 (N_7562,N_6859,N_5178);
nor U7563 (N_7563,N_6224,N_5327);
nor U7564 (N_7564,N_5131,N_5623);
nor U7565 (N_7565,N_7100,N_5276);
nand U7566 (N_7566,N_7095,N_6424);
or U7567 (N_7567,N_6539,N_6175);
nor U7568 (N_7568,N_5510,N_6133);
nor U7569 (N_7569,N_6231,N_5639);
and U7570 (N_7570,N_5476,N_7267);
xnor U7571 (N_7571,N_6492,N_6047);
nor U7572 (N_7572,N_5796,N_6319);
nand U7573 (N_7573,N_7282,N_5666);
nand U7574 (N_7574,N_6958,N_5192);
xnor U7575 (N_7575,N_6002,N_5648);
or U7576 (N_7576,N_5398,N_7078);
and U7577 (N_7577,N_6034,N_6083);
nand U7578 (N_7578,N_6431,N_6361);
nand U7579 (N_7579,N_6032,N_6408);
nor U7580 (N_7580,N_5745,N_6837);
or U7581 (N_7581,N_6576,N_6367);
or U7582 (N_7582,N_6964,N_6828);
nand U7583 (N_7583,N_5242,N_6804);
xor U7584 (N_7584,N_5292,N_6168);
nand U7585 (N_7585,N_6145,N_5873);
nand U7586 (N_7586,N_5917,N_5033);
nor U7587 (N_7587,N_5037,N_6510);
xnor U7588 (N_7588,N_6344,N_5698);
xnor U7589 (N_7589,N_5838,N_7044);
nor U7590 (N_7590,N_7007,N_5050);
nor U7591 (N_7591,N_6978,N_7323);
or U7592 (N_7592,N_6291,N_6625);
nand U7593 (N_7593,N_5531,N_6940);
and U7594 (N_7594,N_5056,N_6983);
nor U7595 (N_7595,N_5057,N_6765);
nor U7596 (N_7596,N_6222,N_6392);
nand U7597 (N_7597,N_6632,N_7202);
xor U7598 (N_7598,N_7305,N_5090);
nand U7599 (N_7599,N_5554,N_5458);
nand U7600 (N_7600,N_6406,N_7294);
and U7601 (N_7601,N_7429,N_5528);
nor U7602 (N_7602,N_6283,N_6690);
or U7603 (N_7603,N_5272,N_6483);
nand U7604 (N_7604,N_6743,N_5283);
and U7605 (N_7605,N_5871,N_6548);
nand U7606 (N_7606,N_6694,N_6144);
and U7607 (N_7607,N_6310,N_5940);
or U7608 (N_7608,N_5798,N_7466);
and U7609 (N_7609,N_7031,N_5307);
or U7610 (N_7610,N_5225,N_5218);
nand U7611 (N_7611,N_7217,N_6608);
and U7612 (N_7612,N_6898,N_7378);
nor U7613 (N_7613,N_6093,N_6401);
nand U7614 (N_7614,N_5817,N_6973);
and U7615 (N_7615,N_6085,N_5456);
or U7616 (N_7616,N_5768,N_5730);
nor U7617 (N_7617,N_6751,N_6302);
or U7618 (N_7618,N_6531,N_5947);
and U7619 (N_7619,N_7374,N_6365);
nand U7620 (N_7620,N_5215,N_6584);
nor U7621 (N_7621,N_6174,N_7103);
xnor U7622 (N_7622,N_7373,N_5644);
nor U7623 (N_7623,N_7084,N_6792);
or U7624 (N_7624,N_5643,N_6985);
and U7625 (N_7625,N_6557,N_7060);
xor U7626 (N_7626,N_6703,N_6391);
or U7627 (N_7627,N_6228,N_6195);
xor U7628 (N_7628,N_5994,N_5862);
xnor U7629 (N_7629,N_5937,N_7467);
and U7630 (N_7630,N_7037,N_5699);
nand U7631 (N_7631,N_5713,N_6778);
xnor U7632 (N_7632,N_6030,N_6794);
or U7633 (N_7633,N_6960,N_5500);
or U7634 (N_7634,N_6239,N_5690);
nand U7635 (N_7635,N_7134,N_6721);
nor U7636 (N_7636,N_7405,N_5332);
and U7637 (N_7637,N_6838,N_6653);
nor U7638 (N_7638,N_5434,N_7314);
and U7639 (N_7639,N_5585,N_5575);
xor U7640 (N_7640,N_6087,N_5155);
xor U7641 (N_7641,N_7003,N_6027);
xor U7642 (N_7642,N_5650,N_7226);
nand U7643 (N_7643,N_6165,N_6123);
nand U7644 (N_7644,N_6044,N_6241);
xnor U7645 (N_7645,N_5011,N_5723);
xor U7646 (N_7646,N_5816,N_5141);
nor U7647 (N_7647,N_5603,N_6250);
xnor U7648 (N_7648,N_6710,N_6142);
xnor U7649 (N_7649,N_5651,N_7244);
nand U7650 (N_7650,N_6790,N_5609);
nand U7651 (N_7651,N_5162,N_6885);
or U7652 (N_7652,N_7086,N_6803);
or U7653 (N_7653,N_5377,N_6399);
xnor U7654 (N_7654,N_6153,N_5508);
or U7655 (N_7655,N_7360,N_5087);
or U7656 (N_7656,N_5200,N_7163);
nand U7657 (N_7657,N_5928,N_6349);
or U7658 (N_7658,N_5509,N_5341);
nor U7659 (N_7659,N_5156,N_6180);
and U7660 (N_7660,N_7106,N_6275);
nor U7661 (N_7661,N_7193,N_5966);
and U7662 (N_7662,N_5188,N_5413);
nor U7663 (N_7663,N_6207,N_6443);
or U7664 (N_7664,N_5302,N_5645);
xnor U7665 (N_7665,N_5891,N_7208);
or U7666 (N_7666,N_6733,N_6696);
xnor U7667 (N_7667,N_5887,N_7087);
and U7668 (N_7668,N_6327,N_5911);
nor U7669 (N_7669,N_6836,N_6639);
nand U7670 (N_7670,N_5657,N_5562);
nor U7671 (N_7671,N_6376,N_5636);
nor U7672 (N_7672,N_5054,N_6582);
nand U7673 (N_7673,N_6693,N_5211);
or U7674 (N_7674,N_6173,N_5962);
or U7675 (N_7675,N_6422,N_5985);
nor U7676 (N_7676,N_6533,N_5685);
xnor U7677 (N_7677,N_7138,N_5736);
or U7678 (N_7678,N_6905,N_5426);
nand U7679 (N_7679,N_5261,N_5244);
xnor U7680 (N_7680,N_5535,N_6309);
and U7681 (N_7681,N_6661,N_5007);
nor U7682 (N_7682,N_6966,N_7338);
xnor U7683 (N_7683,N_7337,N_5052);
nor U7684 (N_7684,N_6234,N_6516);
nor U7685 (N_7685,N_5755,N_5637);
and U7686 (N_7686,N_6706,N_7312);
nand U7687 (N_7687,N_7158,N_7231);
or U7688 (N_7688,N_5320,N_6990);
xor U7689 (N_7689,N_6256,N_6644);
and U7690 (N_7690,N_5829,N_7030);
xnor U7691 (N_7691,N_7235,N_6835);
nor U7692 (N_7692,N_6954,N_5284);
and U7693 (N_7693,N_6596,N_5684);
xor U7694 (N_7694,N_6612,N_5104);
nor U7695 (N_7695,N_5346,N_5385);
nand U7696 (N_7696,N_6411,N_6342);
and U7697 (N_7697,N_7280,N_5611);
nor U7698 (N_7698,N_7383,N_5652);
nor U7699 (N_7699,N_6611,N_5918);
nand U7700 (N_7700,N_7301,N_5709);
xnor U7701 (N_7701,N_6839,N_7347);
nor U7702 (N_7702,N_6301,N_5879);
xnor U7703 (N_7703,N_6050,N_6763);
and U7704 (N_7704,N_7413,N_5980);
or U7705 (N_7705,N_6923,N_5117);
xor U7706 (N_7706,N_6979,N_5975);
and U7707 (N_7707,N_6633,N_6200);
xnor U7708 (N_7708,N_6605,N_7041);
xnor U7709 (N_7709,N_7443,N_5961);
nor U7710 (N_7710,N_5759,N_5976);
and U7711 (N_7711,N_6638,N_5447);
nor U7712 (N_7712,N_5391,N_5137);
nor U7713 (N_7713,N_7033,N_7082);
or U7714 (N_7714,N_5970,N_7247);
or U7715 (N_7715,N_6230,N_5522);
or U7716 (N_7716,N_5749,N_5223);
nand U7717 (N_7717,N_7341,N_7075);
and U7718 (N_7718,N_7461,N_5371);
nor U7719 (N_7719,N_5614,N_7488);
xnor U7720 (N_7720,N_6992,N_5146);
or U7721 (N_7721,N_6380,N_6537);
nor U7722 (N_7722,N_6164,N_6854);
nand U7723 (N_7723,N_6345,N_6936);
nand U7724 (N_7724,N_6248,N_6779);
xnor U7725 (N_7725,N_6521,N_6813);
nor U7726 (N_7726,N_5436,N_7257);
nor U7727 (N_7727,N_6042,N_5496);
and U7728 (N_7728,N_5794,N_6645);
or U7729 (N_7729,N_6387,N_5805);
xor U7730 (N_7730,N_6613,N_5473);
and U7731 (N_7731,N_7076,N_6282);
xnor U7732 (N_7732,N_6969,N_7046);
nand U7733 (N_7733,N_7480,N_6128);
or U7734 (N_7734,N_5919,N_7427);
nor U7735 (N_7735,N_5486,N_5837);
xnor U7736 (N_7736,N_6143,N_5519);
nor U7737 (N_7737,N_7079,N_6353);
xnor U7738 (N_7738,N_7148,N_6815);
nand U7739 (N_7739,N_7418,N_5586);
nor U7740 (N_7740,N_6102,N_5285);
or U7741 (N_7741,N_5064,N_6225);
xor U7742 (N_7742,N_5275,N_5809);
and U7743 (N_7743,N_5116,N_6331);
nor U7744 (N_7744,N_6997,N_6993);
or U7745 (N_7745,N_6865,N_5420);
nand U7746 (N_7746,N_5334,N_5905);
and U7747 (N_7747,N_5471,N_5118);
or U7748 (N_7748,N_6481,N_5299);
xor U7749 (N_7749,N_6129,N_7315);
nand U7750 (N_7750,N_6500,N_6773);
or U7751 (N_7751,N_6324,N_6927);
and U7752 (N_7752,N_5414,N_6218);
nor U7753 (N_7753,N_5596,N_5232);
and U7754 (N_7754,N_5366,N_5881);
nor U7755 (N_7755,N_6212,N_6853);
nor U7756 (N_7756,N_5392,N_7483);
or U7757 (N_7757,N_5948,N_6495);
xor U7758 (N_7758,N_6595,N_6354);
or U7759 (N_7759,N_5716,N_6829);
nor U7760 (N_7760,N_5950,N_7400);
and U7761 (N_7761,N_6160,N_6886);
or U7762 (N_7762,N_5857,N_6429);
or U7763 (N_7763,N_6744,N_7140);
nand U7764 (N_7764,N_5265,N_5804);
nand U7765 (N_7765,N_5892,N_5597);
and U7766 (N_7766,N_7069,N_5222);
and U7767 (N_7767,N_6251,N_6460);
or U7768 (N_7768,N_5679,N_6541);
or U7769 (N_7769,N_7090,N_6038);
nor U7770 (N_7770,N_5963,N_5167);
nand U7771 (N_7771,N_7214,N_7384);
and U7772 (N_7772,N_7269,N_5973);
or U7773 (N_7773,N_7062,N_7394);
and U7774 (N_7774,N_6255,N_5799);
nor U7775 (N_7775,N_5144,N_5579);
nand U7776 (N_7776,N_7320,N_7449);
xnor U7777 (N_7777,N_7210,N_5939);
or U7778 (N_7778,N_5309,N_5972);
xor U7779 (N_7779,N_6514,N_5708);
or U7780 (N_7780,N_6294,N_5402);
nand U7781 (N_7781,N_7113,N_7489);
and U7782 (N_7782,N_6172,N_6238);
and U7783 (N_7783,N_5328,N_7331);
and U7784 (N_7784,N_6926,N_6941);
or U7785 (N_7785,N_7232,N_7408);
nand U7786 (N_7786,N_6780,N_6151);
and U7787 (N_7787,N_6432,N_6845);
or U7788 (N_7788,N_6665,N_6092);
nor U7789 (N_7789,N_7256,N_6303);
nor U7790 (N_7790,N_5608,N_6683);
and U7791 (N_7791,N_5105,N_5686);
nor U7792 (N_7792,N_6702,N_5164);
and U7793 (N_7793,N_6243,N_6107);
or U7794 (N_7794,N_7189,N_6720);
nand U7795 (N_7795,N_5274,N_6385);
or U7796 (N_7796,N_6842,N_6415);
or U7797 (N_7797,N_5989,N_5375);
and U7798 (N_7798,N_7107,N_5381);
nor U7799 (N_7799,N_6866,N_6598);
xor U7800 (N_7800,N_5789,N_6674);
and U7801 (N_7801,N_6318,N_6560);
nor U7802 (N_7802,N_6215,N_6784);
and U7803 (N_7803,N_5002,N_6581);
and U7804 (N_7804,N_6202,N_6860);
or U7805 (N_7805,N_6336,N_5019);
nor U7806 (N_7806,N_5938,N_7261);
xnor U7807 (N_7807,N_7419,N_5495);
and U7808 (N_7808,N_6101,N_6205);
or U7809 (N_7809,N_6197,N_5537);
nand U7810 (N_7810,N_6651,N_6642);
xnor U7811 (N_7811,N_6728,N_6932);
xor U7812 (N_7812,N_6777,N_6452);
or U7813 (N_7813,N_7333,N_6634);
xor U7814 (N_7814,N_5560,N_5259);
nand U7815 (N_7815,N_5633,N_5815);
and U7816 (N_7816,N_5358,N_7343);
and U7817 (N_7817,N_5360,N_6360);
nand U7818 (N_7818,N_5159,N_5901);
and U7819 (N_7819,N_7000,N_7105);
xnor U7820 (N_7820,N_5077,N_7137);
and U7821 (N_7821,N_6589,N_5240);
and U7822 (N_7822,N_5210,N_6209);
nor U7823 (N_7823,N_7368,N_6446);
and U7824 (N_7824,N_6191,N_5689);
xor U7825 (N_7825,N_7045,N_7054);
nor U7826 (N_7826,N_5110,N_6061);
xnor U7827 (N_7827,N_5766,N_6781);
and U7828 (N_7828,N_6158,N_6447);
or U7829 (N_7829,N_5093,N_5914);
xnor U7830 (N_7830,N_7034,N_5108);
or U7831 (N_7831,N_6602,N_7155);
or U7832 (N_7832,N_5329,N_5147);
xnor U7833 (N_7833,N_5321,N_5123);
and U7834 (N_7834,N_5557,N_5737);
and U7835 (N_7835,N_5477,N_6848);
or U7836 (N_7836,N_6322,N_6497);
and U7837 (N_7837,N_5827,N_7211);
or U7838 (N_7838,N_7319,N_7445);
nand U7839 (N_7839,N_6583,N_5593);
xor U7840 (N_7840,N_7104,N_7136);
nand U7841 (N_7841,N_7259,N_7083);
or U7842 (N_7842,N_6742,N_5181);
and U7843 (N_7843,N_6536,N_5929);
or U7844 (N_7844,N_6668,N_6019);
nor U7845 (N_7845,N_5605,N_7205);
nor U7846 (N_7846,N_5287,N_5154);
nand U7847 (N_7847,N_5694,N_7285);
nand U7848 (N_7848,N_7156,N_5017);
or U7849 (N_7849,N_5527,N_5864);
nand U7850 (N_7850,N_5570,N_6922);
and U7851 (N_7851,N_7474,N_5517);
xor U7852 (N_7852,N_6071,N_6149);
nor U7853 (N_7853,N_7273,N_7064);
and U7854 (N_7854,N_5965,N_5670);
xor U7855 (N_7855,N_7289,N_5170);
nand U7856 (N_7856,N_5843,N_5903);
or U7857 (N_7857,N_5834,N_6490);
nand U7858 (N_7858,N_6098,N_5642);
nand U7859 (N_7859,N_6688,N_6998);
nor U7860 (N_7860,N_5251,N_6599);
nand U7861 (N_7861,N_6919,N_5801);
nor U7862 (N_7862,N_7127,N_6442);
and U7863 (N_7863,N_7017,N_5602);
nand U7864 (N_7864,N_7410,N_6700);
or U7865 (N_7865,N_5673,N_5493);
nand U7866 (N_7866,N_6635,N_5290);
xnor U7867 (N_7867,N_7067,N_5581);
nand U7868 (N_7868,N_5422,N_6570);
or U7869 (N_7869,N_6561,N_5721);
nand U7870 (N_7870,N_5565,N_5536);
xor U7871 (N_7871,N_7420,N_6914);
nand U7872 (N_7872,N_6802,N_5907);
nor U7873 (N_7873,N_5368,N_6585);
nor U7874 (N_7874,N_6730,N_5807);
or U7875 (N_7875,N_5479,N_7481);
and U7876 (N_7876,N_5559,N_6329);
and U7877 (N_7877,N_5810,N_6279);
or U7878 (N_7878,N_6678,N_6321);
xor U7879 (N_7879,N_6325,N_5780);
nand U7880 (N_7880,N_7122,N_7126);
or U7881 (N_7881,N_6025,N_6265);
nor U7882 (N_7882,N_5782,N_5151);
and U7883 (N_7883,N_7304,N_5692);
nand U7884 (N_7884,N_6768,N_7180);
nand U7885 (N_7885,N_6226,N_6136);
and U7886 (N_7886,N_6811,N_5130);
nor U7887 (N_7887,N_6031,N_5595);
nor U7888 (N_7888,N_5055,N_7018);
and U7889 (N_7889,N_6343,N_6405);
or U7890 (N_7890,N_6935,N_7306);
xnor U7891 (N_7891,N_6827,N_6734);
nand U7892 (N_7892,N_7133,N_6461);
nand U7893 (N_7893,N_6760,N_7184);
or U7894 (N_7894,N_5483,N_7065);
or U7895 (N_7895,N_6788,N_5427);
or U7896 (N_7896,N_7262,N_6006);
nor U7897 (N_7897,N_6762,N_5859);
and U7898 (N_7898,N_6412,N_5040);
nor U7899 (N_7899,N_7224,N_6769);
and U7900 (N_7900,N_5069,N_6397);
and U7901 (N_7901,N_6362,N_7376);
nand U7902 (N_7902,N_5467,N_6194);
nand U7903 (N_7903,N_5468,N_6227);
or U7904 (N_7904,N_7219,N_7006);
xnor U7905 (N_7905,N_6039,N_5606);
or U7906 (N_7906,N_6333,N_5540);
and U7907 (N_7907,N_7218,N_6989);
nand U7908 (N_7908,N_5221,N_7380);
and U7909 (N_7909,N_5811,N_5812);
nand U7910 (N_7910,N_7302,N_6188);
and U7911 (N_7911,N_5601,N_5649);
nand U7912 (N_7912,N_7249,N_7188);
xor U7913 (N_7913,N_7171,N_5693);
nor U7914 (N_7914,N_6317,N_6474);
nor U7915 (N_7915,N_6482,N_5830);
nand U7916 (N_7916,N_7390,N_7022);
nand U7917 (N_7917,N_5561,N_5813);
nor U7918 (N_7918,N_7477,N_7317);
nand U7919 (N_7919,N_5418,N_5035);
xnor U7920 (N_7920,N_7275,N_6108);
nor U7921 (N_7921,N_5742,N_5788);
and U7922 (N_7922,N_5526,N_5910);
xnor U7923 (N_7923,N_7270,N_5335);
nand U7924 (N_7924,N_5410,N_5852);
or U7925 (N_7925,N_5543,N_5899);
and U7926 (N_7926,N_6963,N_6867);
nor U7927 (N_7927,N_7416,N_5044);
and U7928 (N_7928,N_7293,N_6819);
nor U7929 (N_7929,N_5260,N_6909);
and U7930 (N_7930,N_5992,N_7063);
and U7931 (N_7931,N_5342,N_6915);
and U7932 (N_7932,N_6808,N_5501);
xnor U7933 (N_7933,N_5298,N_7375);
or U7934 (N_7934,N_6106,N_7146);
nand U7935 (N_7935,N_6924,N_6357);
or U7936 (N_7936,N_5854,N_5209);
or U7937 (N_7937,N_5148,N_6089);
nand U7938 (N_7938,N_5710,N_5201);
or U7939 (N_7939,N_5149,N_6503);
xnor U7940 (N_7940,N_7425,N_7009);
and U7941 (N_7941,N_6273,N_5853);
nand U7942 (N_7942,N_7142,N_7411);
xnor U7943 (N_7943,N_5550,N_5969);
nand U7944 (N_7944,N_5856,N_5818);
xor U7945 (N_7945,N_6300,N_6064);
xor U7946 (N_7946,N_5765,N_6375);
nand U7947 (N_7947,N_6126,N_6040);
nor U7948 (N_7948,N_5851,N_5814);
and U7949 (N_7949,N_7476,N_5520);
and U7950 (N_7950,N_6359,N_6847);
nor U7951 (N_7951,N_7011,N_5008);
nand U7952 (N_7952,N_6080,N_6286);
xor U7953 (N_7953,N_5861,N_5741);
or U7954 (N_7954,N_5701,N_5573);
or U7955 (N_7955,N_5173,N_5998);
xor U7956 (N_7956,N_5424,N_7237);
nand U7957 (N_7957,N_6766,N_6564);
nor U7958 (N_7958,N_6003,N_5262);
or U7959 (N_7959,N_6593,N_6701);
and U7960 (N_7960,N_5835,N_7465);
or U7961 (N_7961,N_6756,N_6176);
and U7962 (N_7962,N_6912,N_5653);
xor U7963 (N_7963,N_5444,N_7080);
xor U7964 (N_7964,N_6208,N_5179);
or U7965 (N_7965,N_6364,N_7109);
nor U7966 (N_7966,N_7396,N_5791);
nand U7967 (N_7967,N_5785,N_6559);
xnor U7968 (N_7968,N_5844,N_5115);
xor U7969 (N_7969,N_5311,N_6505);
nand U7970 (N_7970,N_6348,N_5340);
xnor U7971 (N_7971,N_6394,N_6161);
or U7972 (N_7972,N_6135,N_7329);
nand U7973 (N_7973,N_7177,N_5401);
nand U7974 (N_7974,N_7287,N_5691);
and U7975 (N_7975,N_7367,N_5568);
and U7976 (N_7976,N_7216,N_7191);
and U7977 (N_7977,N_7207,N_7495);
nor U7978 (N_7978,N_5722,N_7014);
or U7979 (N_7979,N_7403,N_6834);
or U7980 (N_7980,N_6988,N_6072);
nand U7981 (N_7981,N_5412,N_6757);
xor U7982 (N_7982,N_6782,N_5359);
xnor U7983 (N_7983,N_5647,N_5408);
nand U7984 (N_7984,N_7241,N_5616);
nand U7985 (N_7985,N_6229,N_7036);
nand U7986 (N_7986,N_5126,N_6373);
and U7987 (N_7987,N_5982,N_5564);
nand U7988 (N_7988,N_6871,N_5697);
and U7989 (N_7989,N_5630,N_6942);
nor U7990 (N_7990,N_5226,N_7209);
or U7991 (N_7991,N_6352,N_6159);
and U7992 (N_7992,N_7243,N_5865);
xnor U7993 (N_7993,N_5631,N_7268);
or U7994 (N_7994,N_6920,N_7169);
xnor U7995 (N_7995,N_6214,N_6455);
or U7996 (N_7996,N_5959,N_5042);
nand U7997 (N_7997,N_7451,N_6896);
nand U7998 (N_7998,N_7272,N_6627);
xor U7999 (N_7999,N_5866,N_7094);
and U8000 (N_8000,N_6725,N_6413);
nor U8001 (N_8001,N_7143,N_6874);
nor U8002 (N_8002,N_6190,N_5999);
nor U8003 (N_8003,N_6587,N_6809);
and U8004 (N_8004,N_6213,N_5993);
nand U8005 (N_8005,N_6697,N_5665);
or U8006 (N_8006,N_5549,N_5877);
and U8007 (N_8007,N_6463,N_6272);
nor U8008 (N_8008,N_6120,N_5066);
or U8009 (N_8009,N_7166,N_6798);
and U8010 (N_8010,N_5431,N_5619);
and U8011 (N_8011,N_6410,N_6947);
or U8012 (N_8012,N_6116,N_5256);
xor U8013 (N_8013,N_6805,N_6551);
nor U8014 (N_8014,N_5049,N_7164);
nand U8015 (N_8015,N_6555,N_5795);
xnor U8016 (N_8016,N_6767,N_5802);
nor U8017 (N_8017,N_6501,N_7212);
or U8018 (N_8018,N_7406,N_5208);
nand U8019 (N_8019,N_7342,N_5589);
and U8020 (N_8020,N_6689,N_5416);
or U8021 (N_8021,N_7318,N_6685);
nor U8022 (N_8022,N_7175,N_6615);
or U8023 (N_8023,N_6755,N_6939);
nand U8024 (N_8024,N_6671,N_7182);
or U8025 (N_8025,N_7026,N_6386);
nand U8026 (N_8026,N_5361,N_6110);
xnor U8027 (N_8027,N_6673,N_6013);
nand U8028 (N_8028,N_7021,N_5705);
xor U8029 (N_8029,N_7493,N_5655);
nand U8030 (N_8030,N_6946,N_6904);
nor U8031 (N_8031,N_7458,N_6592);
nand U8032 (N_8032,N_5230,N_7423);
nand U8033 (N_8033,N_6529,N_6712);
nand U8034 (N_8034,N_7025,N_6822);
nand U8035 (N_8035,N_6196,N_7371);
nor U8036 (N_8036,N_7002,N_6618);
nand U8037 (N_8037,N_6840,N_5793);
nor U8038 (N_8038,N_5640,N_6028);
xnor U8039 (N_8039,N_5687,N_7324);
nor U8040 (N_8040,N_5482,N_7172);
xnor U8041 (N_8041,N_5846,N_7242);
or U8042 (N_8042,N_6513,N_6393);
and U8043 (N_8043,N_5625,N_6049);
and U8044 (N_8044,N_6054,N_6470);
nand U8045 (N_8045,N_5072,N_6862);
or U8046 (N_8046,N_7444,N_6005);
xnor U8047 (N_8047,N_6137,N_5484);
nor U8048 (N_8048,N_7311,N_5499);
and U8049 (N_8049,N_5452,N_6723);
or U8050 (N_8050,N_6046,N_6313);
nand U8051 (N_8051,N_6818,N_6737);
xor U8052 (N_8052,N_5711,N_5632);
and U8053 (N_8053,N_6311,N_6715);
nand U8054 (N_8054,N_5028,N_5516);
and U8055 (N_8055,N_6314,N_5525);
or U8056 (N_8056,N_6400,N_6538);
xor U8057 (N_8057,N_6532,N_7154);
xnor U8058 (N_8058,N_6917,N_7468);
nor U8059 (N_8059,N_6472,N_6414);
xor U8060 (N_8060,N_6929,N_7081);
and U8061 (N_8061,N_6672,N_7027);
nor U8062 (N_8062,N_6789,N_7366);
xnor U8063 (N_8063,N_6270,N_5488);
nor U8064 (N_8064,N_6041,N_5034);
nand U8065 (N_8065,N_5213,N_5883);
nand U8066 (N_8066,N_6379,N_5680);
and U8067 (N_8067,N_5943,N_5250);
or U8068 (N_8068,N_6907,N_7409);
xor U8069 (N_8069,N_5503,N_6109);
xor U8070 (N_8070,N_6018,N_5125);
xor U8071 (N_8071,N_7130,N_5855);
xnor U8072 (N_8072,N_7199,N_5061);
and U8073 (N_8073,N_5354,N_7139);
or U8074 (N_8074,N_7434,N_6236);
or U8075 (N_8075,N_7252,N_7424);
and U8076 (N_8076,N_5005,N_6390);
and U8077 (N_8077,N_6974,N_5556);
or U8078 (N_8078,N_7415,N_7038);
or U8079 (N_8079,N_5800,N_6658);
or U8080 (N_8080,N_6011,N_5386);
nand U8081 (N_8081,N_5305,N_7471);
nand U8082 (N_8082,N_6670,N_5622);
or U8083 (N_8083,N_5091,N_6350);
and U8084 (N_8084,N_6857,N_6258);
xnor U8085 (N_8085,N_6628,N_5454);
and U8086 (N_8086,N_6449,N_5682);
xor U8087 (N_8087,N_5466,N_5336);
or U8088 (N_8088,N_7388,N_6036);
nor U8089 (N_8089,N_5239,N_7077);
nand U8090 (N_8090,N_6271,N_5548);
or U8091 (N_8091,N_7150,N_6965);
and U8092 (N_8092,N_7290,N_5498);
nand U8093 (N_8093,N_5338,N_5583);
or U8094 (N_8094,N_5207,N_6140);
nand U8095 (N_8095,N_6910,N_5460);
xnor U8096 (N_8096,N_6433,N_5070);
nor U8097 (N_8097,N_6707,N_5238);
nand U8098 (N_8098,N_5355,N_6363);
nand U8099 (N_8099,N_6878,N_5363);
nand U8100 (N_8100,N_5580,N_5081);
xor U8101 (N_8101,N_6630,N_6285);
and U8102 (N_8102,N_5744,N_5808);
nor U8103 (N_8103,N_5820,N_6894);
xor U8104 (N_8104,N_5926,N_6187);
xor U8105 (N_8105,N_6192,N_5497);
and U8106 (N_8106,N_6118,N_5518);
and U8107 (N_8107,N_5433,N_6681);
xor U8108 (N_8108,N_6527,N_5584);
nor U8109 (N_8109,N_5964,N_6469);
nor U8110 (N_8110,N_5190,N_5333);
nand U8111 (N_8111,N_6841,N_5435);
and U8112 (N_8112,N_6150,N_6477);
nor U8113 (N_8113,N_6856,N_7131);
nand U8114 (N_8114,N_6558,N_5990);
xnor U8115 (N_8115,N_6468,N_7070);
or U8116 (N_8116,N_6814,N_6021);
or U8117 (N_8117,N_6572,N_6975);
and U8118 (N_8118,N_5107,N_5674);
nor U8119 (N_8119,N_5205,N_7236);
and U8120 (N_8120,N_7454,N_6423);
xor U8121 (N_8121,N_6852,N_7457);
nand U8122 (N_8122,N_6962,N_6580);
and U8123 (N_8123,N_7364,N_6439);
or U8124 (N_8124,N_6793,N_6015);
or U8125 (N_8125,N_7200,N_5119);
or U8126 (N_8126,N_5776,N_5174);
xor U8127 (N_8127,N_5252,N_6082);
or U8128 (N_8128,N_7308,N_6851);
xor U8129 (N_8129,N_6563,N_5445);
xnor U8130 (N_8130,N_6996,N_6577);
nor U8131 (N_8131,N_5863,N_6825);
xor U8132 (N_8132,N_5930,N_5539);
nor U8133 (N_8133,N_7432,N_5894);
and U8134 (N_8134,N_5758,N_5143);
or U8135 (N_8135,N_6786,N_5474);
nand U8136 (N_8136,N_5442,N_5661);
nand U8137 (N_8137,N_5430,N_5604);
and U8138 (N_8138,N_6420,N_6680);
and U8139 (N_8139,N_5120,N_6055);
nand U8140 (N_8140,N_7223,N_7450);
nor U8141 (N_8141,N_6573,N_7151);
and U8142 (N_8142,N_6499,N_6546);
nor U8143 (N_8143,N_5783,N_6620);
nor U8144 (N_8144,N_7145,N_6245);
nand U8145 (N_8145,N_7121,N_5797);
nand U8146 (N_8146,N_5158,N_7401);
nor U8147 (N_8147,N_5612,N_5746);
and U8148 (N_8148,N_5944,N_5004);
nand U8149 (N_8149,N_7332,N_7430);
and U8150 (N_8150,N_6293,N_6649);
nand U8151 (N_8151,N_6378,N_5449);
or U8152 (N_8152,N_7222,N_6384);
xnor U8153 (N_8153,N_5715,N_7431);
nor U8154 (N_8154,N_5667,N_5280);
nor U8155 (N_8155,N_7015,N_5153);
nand U8156 (N_8156,N_6304,N_6824);
and U8157 (N_8157,N_6407,N_6496);
nand U8158 (N_8158,N_6185,N_6986);
and U8159 (N_8159,N_7162,N_7295);
nor U8160 (N_8160,N_7052,N_5097);
nand U8161 (N_8161,N_7051,N_7359);
nor U8162 (N_8162,N_5825,N_5316);
or U8163 (N_8163,N_6016,N_6177);
nand U8164 (N_8164,N_6418,N_6552);
and U8165 (N_8165,N_6456,N_5113);
or U8166 (N_8166,N_6249,N_5051);
or U8167 (N_8167,N_6037,N_7353);
nor U8168 (N_8168,N_6654,N_5076);
and U8169 (N_8169,N_6043,N_7433);
and U8170 (N_8170,N_6750,N_5323);
nor U8171 (N_8171,N_6869,N_5638);
nand U8172 (N_8172,N_7115,N_5127);
nand U8173 (N_8173,N_5921,N_7019);
nand U8174 (N_8174,N_6121,N_6235);
xnor U8175 (N_8175,N_5695,N_7455);
nor U8176 (N_8176,N_6717,N_5182);
and U8177 (N_8177,N_5831,N_7464);
and U8178 (N_8178,N_6607,N_5628);
or U8179 (N_8179,N_5451,N_6545);
nand U8180 (N_8180,N_5176,N_7407);
nand U8181 (N_8181,N_5157,N_5821);
nand U8182 (N_8182,N_5229,N_5348);
nor U8183 (N_8183,N_7393,N_5515);
xnor U8184 (N_8184,N_7178,N_5165);
nand U8185 (N_8185,N_6059,N_7230);
nand U8186 (N_8186,N_7250,N_5312);
nand U8187 (N_8187,N_6502,N_5869);
nor U8188 (N_8188,N_7096,N_5646);
nor U8189 (N_8189,N_5395,N_6772);
and U8190 (N_8190,N_6254,N_7074);
nand U8191 (N_8191,N_6489,N_6094);
or U8192 (N_8192,N_5246,N_5850);
and U8193 (N_8193,N_6276,N_5032);
xor U8194 (N_8194,N_5078,N_6058);
or U8195 (N_8195,N_5634,N_6604);
and U8196 (N_8196,N_6525,N_6014);
and U8197 (N_8197,N_7058,N_7462);
nand U8198 (N_8198,N_5577,N_6719);
nand U8199 (N_8199,N_7001,N_6534);
nor U8200 (N_8200,N_5524,N_5839);
xor U8201 (N_8201,N_6902,N_5664);
and U8202 (N_8202,N_6493,N_6982);
nand U8203 (N_8203,N_6830,N_7355);
or U8204 (N_8204,N_5198,N_6981);
and U8205 (N_8205,N_5196,N_6783);
or U8206 (N_8206,N_6921,N_5885);
or U8207 (N_8207,N_7402,N_6872);
and U8208 (N_8208,N_6068,N_6295);
and U8209 (N_8209,N_7201,N_5824);
xnor U8210 (N_8210,N_5075,N_7125);
xnor U8211 (N_8211,N_6938,N_7258);
or U8212 (N_8212,N_6156,N_6381);
nor U8213 (N_8213,N_6826,N_5884);
nand U8214 (N_8214,N_6682,N_5487);
nor U8215 (N_8215,N_6522,N_6201);
nor U8216 (N_8216,N_5347,N_5502);
xnor U8217 (N_8217,N_5641,N_5833);
or U8218 (N_8218,N_7215,N_6843);
nor U8219 (N_8219,N_6667,N_5013);
and U8220 (N_8220,N_5739,N_6863);
nor U8221 (N_8221,N_5356,N_6617);
xor U8222 (N_8222,N_6745,N_6203);
or U8223 (N_8223,N_7093,N_5547);
and U8224 (N_8224,N_6347,N_5995);
nor U8225 (N_8225,N_5703,N_6930);
nor U8226 (N_8226,N_7028,N_5016);
xnor U8227 (N_8227,N_5688,N_5840);
xor U8228 (N_8228,N_5784,N_6252);
nor U8229 (N_8229,N_6264,N_5934);
nor U8230 (N_8230,N_6119,N_6591);
nand U8231 (N_8231,N_5874,N_5023);
nor U8232 (N_8232,N_5282,N_6507);
and U8233 (N_8233,N_6609,N_6193);
nor U8234 (N_8234,N_5935,N_6574);
nand U8235 (N_8235,N_6112,N_7157);
nand U8236 (N_8236,N_5512,N_6024);
nor U8237 (N_8237,N_6099,N_7437);
nor U8238 (N_8238,N_6566,N_5494);
nor U8239 (N_8239,N_7152,N_5286);
nor U8240 (N_8240,N_5111,N_5507);
xnor U8241 (N_8241,N_7057,N_6754);
nand U8242 (N_8242,N_6186,N_5345);
nand U8243 (N_8243,N_6261,N_7300);
or U8244 (N_8244,N_6267,N_7283);
and U8245 (N_8245,N_6154,N_6646);
nor U8246 (N_8246,N_5216,N_6749);
nor U8247 (N_8247,N_6679,N_7448);
nand U8248 (N_8248,N_6660,N_5770);
or U8249 (N_8249,N_6799,N_7240);
nor U8250 (N_8250,N_5163,N_5683);
xor U8251 (N_8251,N_5576,N_7363);
or U8252 (N_8252,N_5199,N_6686);
nor U8253 (N_8253,N_7196,N_6033);
and U8254 (N_8254,N_5747,N_6440);
and U8255 (N_8255,N_6465,N_5942);
nor U8256 (N_8256,N_6800,N_6844);
nand U8257 (N_8257,N_5318,N_6931);
and U8258 (N_8258,N_6308,N_6961);
nor U8259 (N_8259,N_5082,N_5981);
xnor U8260 (N_8260,N_6138,N_7108);
nor U8261 (N_8261,N_5906,N_5367);
nand U8262 (N_8262,N_5085,N_5823);
and U8263 (N_8263,N_7292,N_7135);
xnor U8264 (N_8264,N_5195,N_5668);
nand U8265 (N_8265,N_6656,N_5924);
nand U8266 (N_8266,N_6579,N_6736);
and U8267 (N_8267,N_6925,N_5591);
xor U8268 (N_8268,N_6009,N_7349);
xor U8269 (N_8269,N_5220,N_5478);
and U8270 (N_8270,N_5872,N_6070);
and U8271 (N_8271,N_6727,N_6206);
or U8272 (N_8272,N_7494,N_6045);
nand U8273 (N_8273,N_7255,N_6664);
or U8274 (N_8274,N_5288,N_5310);
xor U8275 (N_8275,N_6614,N_7239);
nor U8276 (N_8276,N_6597,N_6911);
nor U8277 (N_8277,N_7248,N_6163);
nor U8278 (N_8278,N_7167,N_5720);
nand U8279 (N_8279,N_6868,N_5303);
or U8280 (N_8280,N_7486,N_5058);
xor U8281 (N_8281,N_6453,N_7321);
and U8282 (N_8282,N_5432,N_5778);
and U8283 (N_8283,N_6601,N_5480);
xnor U8284 (N_8284,N_5140,N_7358);
or U8285 (N_8285,N_6060,N_6900);
xnor U8286 (N_8286,N_5889,N_7426);
nor U8287 (N_8287,N_5001,N_6676);
and U8288 (N_8288,N_7225,N_7264);
or U8289 (N_8289,N_5026,N_5566);
or U8290 (N_8290,N_5364,N_6897);
or U8291 (N_8291,N_6280,N_6155);
or U8292 (N_8292,N_5233,N_7088);
nor U8293 (N_8293,N_5627,N_5212);
nand U8294 (N_8294,N_6528,N_5743);
or U8295 (N_8295,N_7213,N_5393);
xnor U8296 (N_8296,N_5080,N_6832);
xor U8297 (N_8297,N_6562,N_7395);
xor U8298 (N_8298,N_6972,N_7123);
xnor U8299 (N_8299,N_5036,N_5624);
nor U8300 (N_8300,N_7161,N_5828);
and U8301 (N_8301,N_5268,N_5369);
xor U8302 (N_8302,N_5659,N_6636);
or U8303 (N_8303,N_5552,N_5931);
nand U8304 (N_8304,N_5015,N_7276);
xor U8305 (N_8305,N_5429,N_5594);
nor U8306 (N_8306,N_6356,N_5134);
nand U8307 (N_8307,N_7043,N_6785);
xor U8308 (N_8308,N_6951,N_6298);
xor U8309 (N_8309,N_5317,N_6883);
or U8310 (N_8310,N_5439,N_5956);
nor U8311 (N_8311,N_5567,N_7310);
and U8312 (N_8312,N_6735,N_5753);
or U8313 (N_8313,N_7118,N_6169);
nand U8314 (N_8314,N_5902,N_6726);
xor U8315 (N_8315,N_7173,N_6297);
nor U8316 (N_8316,N_5122,N_6643);
or U8317 (N_8317,N_6435,N_6220);
xnor U8318 (N_8318,N_7326,N_6542);
xnor U8319 (N_8319,N_6711,N_7050);
nand U8320 (N_8320,N_7153,N_7141);
and U8321 (N_8321,N_5394,N_5247);
xnor U8322 (N_8322,N_7144,N_5769);
and U8323 (N_8323,N_7179,N_5916);
xnor U8324 (N_8324,N_6450,N_5706);
xnor U8325 (N_8325,N_5886,N_6130);
nor U8326 (N_8326,N_5236,N_5752);
nand U8327 (N_8327,N_6892,N_6464);
nand U8328 (N_8328,N_5656,N_5618);
and U8329 (N_8329,N_5678,N_5511);
nand U8330 (N_8330,N_5403,N_5046);
nor U8331 (N_8331,N_5245,N_7475);
nand U8332 (N_8332,N_5485,N_6624);
nand U8333 (N_8333,N_6419,N_5936);
nand U8334 (N_8334,N_5836,N_6346);
nor U8335 (N_8335,N_6232,N_5373);
or U8336 (N_8336,N_6022,N_6323);
and U8337 (N_8337,N_6117,N_6103);
xnor U8338 (N_8338,N_5234,N_5150);
or U8339 (N_8339,N_5671,N_7265);
nand U8340 (N_8340,N_6467,N_5728);
and U8341 (N_8341,N_6487,N_6699);
or U8342 (N_8342,N_6148,N_6355);
and U8343 (N_8343,N_6368,N_7195);
nor U8344 (N_8344,N_6260,N_6079);
nand U8345 (N_8345,N_6714,N_6820);
nand U8346 (N_8346,N_5098,N_6115);
xor U8347 (N_8347,N_6623,N_5103);
nor U8348 (N_8348,N_6398,N_6000);
xnor U8349 (N_8349,N_6741,N_5841);
xnor U8350 (N_8350,N_6994,N_5279);
xor U8351 (N_8351,N_7110,N_5277);
and U8352 (N_8352,N_7442,N_6823);
xor U8353 (N_8353,N_6953,N_5357);
nand U8354 (N_8354,N_6001,N_6567);
xnor U8355 (N_8355,N_5294,N_7334);
xor U8356 (N_8356,N_6858,N_5729);
or U8357 (N_8357,N_6396,N_6162);
xnor U8358 (N_8358,N_5986,N_6709);
xor U8359 (N_8359,N_6010,N_6889);
nor U8360 (N_8360,N_7284,N_5847);
nand U8361 (N_8361,N_6269,N_5849);
nor U8362 (N_8362,N_6957,N_6416);
nand U8363 (N_8363,N_6877,N_5390);
xnor U8364 (N_8364,N_7049,N_5945);
or U8365 (N_8365,N_5984,N_5038);
and U8366 (N_8366,N_6292,N_6652);
or U8367 (N_8367,N_6509,N_7066);
and U8368 (N_8368,N_6807,N_5228);
xor U8369 (N_8369,N_5308,N_6478);
and U8370 (N_8370,N_5725,N_7040);
nand U8371 (N_8371,N_6669,N_6691);
nor U8372 (N_8372,N_5183,N_6518);
nand U8373 (N_8373,N_5314,N_5571);
or U8374 (N_8374,N_7277,N_5264);
nor U8375 (N_8375,N_6216,N_5781);
nor U8376 (N_8376,N_6880,N_6606);
or U8377 (N_8377,N_6849,N_7245);
or U8378 (N_8378,N_5059,N_5443);
nor U8379 (N_8379,N_5533,N_6454);
or U8380 (N_8380,N_6268,N_5083);
or U8381 (N_8381,N_5100,N_7297);
nor U8382 (N_8382,N_6967,N_5376);
nand U8383 (N_8383,N_5465,N_5101);
and U8384 (N_8384,N_5967,N_5772);
nor U8385 (N_8385,N_6290,N_5756);
nor U8386 (N_8386,N_6332,N_7220);
and U8387 (N_8387,N_6881,N_6873);
nor U8388 (N_8388,N_5406,N_6933);
xnor U8389 (N_8389,N_5538,N_5748);
or U8390 (N_8390,N_5592,N_5957);
xnor U8391 (N_8391,N_5660,N_7460);
or U8392 (N_8392,N_5030,N_7496);
or U8393 (N_8393,N_5074,N_6775);
xnor U8394 (N_8394,N_5775,N_6698);
and U8395 (N_8395,N_7198,N_5717);
nand U8396 (N_8396,N_5289,N_7386);
nand U8397 (N_8397,N_6621,N_6437);
nor U8398 (N_8398,N_6511,N_5541);
nor U8399 (N_8399,N_5291,N_5617);
xor U8400 (N_8400,N_5738,N_5504);
xor U8401 (N_8401,N_5191,N_6526);
nor U8402 (N_8402,N_6451,N_6402);
xor U8403 (N_8403,N_5263,N_6722);
nand U8404 (N_8404,N_7441,N_5958);
nand U8405 (N_8405,N_5893,N_5607);
xnor U8406 (N_8406,N_6330,N_5350);
and U8407 (N_8407,N_7452,N_5915);
nor U8408 (N_8408,N_7412,N_6369);
and U8409 (N_8409,N_6246,N_6388);
nor U8410 (N_8410,N_6530,N_7499);
or U8411 (N_8411,N_6801,N_5217);
and U8412 (N_8412,N_5767,N_5253);
xnor U8413 (N_8413,N_7260,N_5734);
nand U8414 (N_8414,N_5724,N_5326);
nand U8415 (N_8415,N_7335,N_5180);
nor U8416 (N_8416,N_7238,N_7459);
xor U8417 (N_8417,N_6320,N_7382);
or U8418 (N_8418,N_6740,N_6113);
and U8419 (N_8419,N_6937,N_6684);
and U8420 (N_8420,N_5750,N_5324);
xnor U8421 (N_8421,N_5132,N_5271);
xnor U8422 (N_8422,N_5136,N_7029);
xor U8423 (N_8423,N_6956,N_5675);
and U8424 (N_8424,N_6170,N_6647);
or U8425 (N_8425,N_5124,N_6692);
nand U8426 (N_8426,N_6053,N_7381);
nor U8427 (N_8427,N_5733,N_5490);
nor U8428 (N_8428,N_5337,N_7485);
xnor U8429 (N_8429,N_7204,N_5099);
or U8430 (N_8430,N_7004,N_5489);
and U8431 (N_8431,N_7048,N_6515);
nor U8432 (N_8432,N_7271,N_6787);
or U8433 (N_8433,N_5374,N_7362);
and U8434 (N_8434,N_5475,N_5020);
xor U8435 (N_8435,N_6899,N_7012);
or U8436 (N_8436,N_5241,N_6178);
or U8437 (N_8437,N_7354,N_7159);
nor U8438 (N_8438,N_5726,N_7446);
nand U8439 (N_8439,N_7117,N_5092);
nand U8440 (N_8440,N_6970,N_6637);
nand U8441 (N_8441,N_6240,N_6629);
nand U8442 (N_8442,N_5949,N_6713);
xor U8443 (N_8443,N_6466,N_6882);
nor U8444 (N_8444,N_6007,N_5448);
nor U8445 (N_8445,N_6504,N_6543);
xnor U8446 (N_8446,N_5405,N_7266);
xnor U8447 (N_8447,N_6724,N_5365);
nor U8448 (N_8448,N_6315,N_6299);
nand U8449 (N_8449,N_5704,N_6675);
nor U8450 (N_8450,N_5621,N_6096);
nand U8451 (N_8451,N_5400,N_5203);
nand U8452 (N_8452,N_6704,N_6776);
xnor U8453 (N_8453,N_5186,N_6850);
xor U8454 (N_8454,N_6655,N_5895);
or U8455 (N_8455,N_5351,N_5202);
and U8456 (N_8456,N_5740,N_5569);
or U8457 (N_8457,N_5932,N_5848);
nor U8458 (N_8458,N_6383,N_6457);
xnor U8459 (N_8459,N_6086,N_5142);
nor U8460 (N_8460,N_7149,N_5380);
xor U8461 (N_8461,N_6705,N_5662);
nor U8462 (N_8462,N_5128,N_6918);
nor U8463 (N_8463,N_6571,N_7254);
xnor U8464 (N_8464,N_6657,N_7089);
xor U8465 (N_8465,N_5089,N_7251);
xnor U8466 (N_8466,N_6968,N_6421);
nand U8467 (N_8467,N_5168,N_7361);
nand U8468 (N_8468,N_5974,N_6831);
xor U8469 (N_8469,N_5304,N_5000);
nor U8470 (N_8470,N_7111,N_5663);
nor U8471 (N_8471,N_6764,N_6127);
nor U8472 (N_8472,N_6088,N_5757);
or U8473 (N_8473,N_6590,N_5379);
nor U8474 (N_8474,N_7187,N_6012);
and U8475 (N_8475,N_6152,N_7010);
xor U8476 (N_8476,N_7497,N_7071);
nor U8477 (N_8477,N_5777,N_5946);
nor U8478 (N_8478,N_5440,N_5978);
nand U8479 (N_8479,N_7453,N_6358);
and U8480 (N_8480,N_6090,N_7274);
and U8481 (N_8481,N_5492,N_5923);
xor U8482 (N_8482,N_7203,N_5068);
nand U8483 (N_8483,N_7116,N_5461);
or U8484 (N_8484,N_6934,N_5160);
nand U8485 (N_8485,N_6603,N_5396);
and U8486 (N_8486,N_5764,N_5773);
nor U8487 (N_8487,N_5224,N_5043);
nor U8488 (N_8488,N_5417,N_7484);
or U8489 (N_8489,N_6066,N_7233);
and U8490 (N_8490,N_6650,N_5187);
nand U8491 (N_8491,N_5214,N_7414);
xnor U8492 (N_8492,N_7286,N_6498);
xor U8493 (N_8493,N_5009,N_7147);
nand U8494 (N_8494,N_6549,N_5900);
or U8495 (N_8495,N_5152,N_7053);
and U8496 (N_8496,N_5257,N_7023);
nor U8497 (N_8497,N_5145,N_6434);
xnor U8498 (N_8498,N_6523,N_6448);
and U8499 (N_8499,N_5411,N_7372);
nor U8500 (N_8500,N_5787,N_5114);
xnor U8501 (N_8501,N_6626,N_5248);
nand U8502 (N_8502,N_5322,N_5372);
and U8503 (N_8503,N_5339,N_6288);
nor U8504 (N_8504,N_6732,N_6097);
or U8505 (N_8505,N_5039,N_7132);
xor U8506 (N_8506,N_5018,N_5909);
or U8507 (N_8507,N_6166,N_5189);
nand U8508 (N_8508,N_6075,N_5021);
xnor U8509 (N_8509,N_6395,N_5184);
or U8510 (N_8510,N_5530,N_6928);
and U8511 (N_8511,N_7114,N_7170);
or U8512 (N_8512,N_6903,N_5330);
or U8513 (N_8513,N_7492,N_6084);
nor U8514 (N_8514,N_6476,N_6063);
nor U8515 (N_8515,N_6233,N_7397);
nor U8516 (N_8516,N_6520,N_5472);
nand U8517 (N_8517,N_7042,N_6855);
and U8518 (N_8518,N_6008,N_5031);
nand U8519 (N_8519,N_6494,N_5462);
nor U8520 (N_8520,N_5913,N_6328);
nand U8521 (N_8521,N_6879,N_5532);
nand U8522 (N_8522,N_7263,N_7316);
and U8523 (N_8523,N_6296,N_5933);
nor U8524 (N_8524,N_6508,N_6795);
nand U8525 (N_8525,N_6659,N_5463);
nor U8526 (N_8526,N_6991,N_7059);
xor U8527 (N_8527,N_7024,N_7479);
nor U8528 (N_8528,N_5983,N_6370);
nor U8529 (N_8529,N_5384,N_7013);
and U8530 (N_8530,N_7112,N_6065);
nand U8531 (N_8531,N_5542,N_5185);
xor U8532 (N_8532,N_5296,N_7085);
or U8533 (N_8533,N_5888,N_5702);
nand U8534 (N_8534,N_6262,N_5206);
and U8535 (N_8535,N_6067,N_6708);
nor U8536 (N_8536,N_7369,N_7183);
or U8537 (N_8537,N_5521,N_5014);
nor U8538 (N_8538,N_6550,N_5832);
nor U8539 (N_8539,N_5563,N_5370);
nor U8540 (N_8540,N_6146,N_5598);
xor U8541 (N_8541,N_5544,N_5270);
xnor U8542 (N_8542,N_6759,N_7291);
nand U8543 (N_8543,N_7340,N_5073);
or U8544 (N_8544,N_5067,N_5868);
or U8545 (N_8545,N_6334,N_6341);
nand U8546 (N_8546,N_5071,N_6111);
or U8547 (N_8547,N_5306,N_7221);
or U8548 (N_8548,N_5654,N_5896);
and U8549 (N_8549,N_5620,N_6980);
nand U8550 (N_8550,N_7392,N_7399);
and U8551 (N_8551,N_7227,N_6374);
or U8552 (N_8552,N_5237,N_5672);
nand U8553 (N_8553,N_5506,N_7350);
nand U8554 (N_8554,N_7490,N_7325);
xor U8555 (N_8555,N_5109,N_6662);
and U8556 (N_8556,N_5166,N_7246);
and U8557 (N_8557,N_6971,N_6114);
nor U8558 (N_8558,N_5027,N_5822);
and U8559 (N_8559,N_6512,N_6073);
nand U8560 (N_8560,N_6648,N_6506);
xor U8561 (N_8561,N_5845,N_6199);
or U8562 (N_8562,N_6758,N_5774);
xor U8563 (N_8563,N_6204,N_7470);
and U8564 (N_8564,N_5003,N_5313);
nand U8565 (N_8565,N_6139,N_6977);
nor U8566 (N_8566,N_5172,N_6257);
xnor U8567 (N_8567,N_5658,N_5269);
and U8568 (N_8568,N_5951,N_7032);
nor U8569 (N_8569,N_6619,N_5006);
and U8570 (N_8570,N_6471,N_6887);
nand U8571 (N_8571,N_6219,N_7352);
and U8572 (N_8572,N_5254,N_6547);
nand U8573 (N_8573,N_5469,N_6695);
or U8574 (N_8574,N_6289,N_7035);
or U8575 (N_8575,N_7339,N_6575);
or U8576 (N_8576,N_5545,N_6444);
and U8577 (N_8577,N_5826,N_5319);
or U8578 (N_8578,N_6553,N_5048);
nor U8579 (N_8579,N_5171,N_6048);
xnor U8580 (N_8580,N_5193,N_7206);
xor U8581 (N_8581,N_6488,N_6459);
or U8582 (N_8582,N_7398,N_6441);
and U8583 (N_8583,N_6916,N_5819);
or U8584 (N_8584,N_5425,N_5954);
or U8585 (N_8585,N_6417,N_5404);
nor U8586 (N_8586,N_6095,N_7056);
and U8587 (N_8587,N_6984,N_7016);
xnor U8588 (N_8588,N_5135,N_6382);
or U8589 (N_8589,N_5399,N_5898);
xnor U8590 (N_8590,N_5095,N_5053);
nand U8591 (N_8591,N_5977,N_5574);
or U8592 (N_8592,N_6366,N_5353);
nor U8593 (N_8593,N_6377,N_6753);
nand U8594 (N_8594,N_5266,N_6141);
or U8595 (N_8595,N_7365,N_5513);
nor U8596 (N_8596,N_6821,N_5925);
nor U8597 (N_8597,N_5751,N_6876);
or U8598 (N_8598,N_7473,N_5763);
nand U8599 (N_8599,N_5197,N_5464);
xor U8600 (N_8600,N_5858,N_7288);
xor U8601 (N_8601,N_5669,N_6247);
or U8602 (N_8602,N_6908,N_6051);
xor U8603 (N_8603,N_5996,N_5803);
or U8604 (N_8604,N_5792,N_5491);
xor U8605 (N_8605,N_6716,N_5086);
nand U8606 (N_8606,N_6578,N_7299);
xor U8607 (N_8607,N_5870,N_5459);
or U8608 (N_8608,N_7101,N_6004);
xnor U8609 (N_8609,N_6287,N_7482);
or U8610 (N_8610,N_5534,N_5719);
and U8611 (N_8611,N_7351,N_5297);
nor U8612 (N_8612,N_7073,N_6812);
and U8613 (N_8613,N_7440,N_6901);
or U8614 (N_8614,N_5867,N_6077);
nand U8615 (N_8615,N_5514,N_7055);
nor U8616 (N_8616,N_5629,N_5349);
xnor U8617 (N_8617,N_5572,N_6056);
and U8618 (N_8618,N_5047,N_7185);
or U8619 (N_8619,N_5587,N_7181);
nand U8620 (N_8620,N_6817,N_7278);
nor U8621 (N_8621,N_6105,N_5024);
nand U8622 (N_8622,N_7168,N_6640);
or U8623 (N_8623,N_6179,N_6796);
xnor U8624 (N_8624,N_6389,N_5904);
and U8625 (N_8625,N_6147,N_7377);
xor U8626 (N_8626,N_5453,N_5960);
nand U8627 (N_8627,N_6182,N_7047);
xnor U8628 (N_8628,N_5997,N_6895);
xor U8629 (N_8629,N_5300,N_5231);
or U8630 (N_8630,N_6747,N_5079);
nor U8631 (N_8631,N_5635,N_5029);
xnor U8632 (N_8632,N_6797,N_5102);
nor U8633 (N_8633,N_7279,N_5382);
nor U8634 (N_8634,N_5428,N_7102);
nand U8635 (N_8635,N_7387,N_5267);
or U8636 (N_8636,N_6445,N_7303);
or U8637 (N_8637,N_6631,N_5890);
nor U8638 (N_8638,N_6586,N_5362);
nor U8639 (N_8639,N_5281,N_6122);
xor U8640 (N_8640,N_5676,N_5012);
xor U8641 (N_8641,N_5293,N_5295);
and U8642 (N_8642,N_6221,N_7370);
nand U8643 (N_8643,N_5762,N_6404);
nand U8644 (N_8644,N_7008,N_6949);
or U8645 (N_8645,N_6326,N_6554);
nand U8646 (N_8646,N_5455,N_6237);
nor U8647 (N_8647,N_6738,N_6259);
xnor U8648 (N_8648,N_5922,N_6340);
xnor U8649 (N_8649,N_7422,N_6524);
nor U8650 (N_8650,N_7357,N_6074);
nand U8651 (N_8651,N_6305,N_6278);
and U8652 (N_8652,N_6189,N_5760);
and U8653 (N_8653,N_5941,N_5878);
and U8654 (N_8654,N_7498,N_7379);
nand U8655 (N_8655,N_6312,N_6473);
xor U8656 (N_8656,N_6565,N_5177);
and U8657 (N_8657,N_6184,N_6167);
nor U8658 (N_8658,N_7005,N_5022);
and U8659 (N_8659,N_6425,N_5045);
and U8660 (N_8660,N_7298,N_6569);
and U8661 (N_8661,N_6944,N_5696);
or U8662 (N_8662,N_6535,N_6666);
nand U8663 (N_8663,N_5987,N_5352);
nand U8664 (N_8664,N_5084,N_5407);
and U8665 (N_8665,N_5718,N_7091);
or U8666 (N_8666,N_6959,N_7356);
and U8667 (N_8667,N_6035,N_6458);
or U8668 (N_8668,N_6731,N_6616);
nand U8669 (N_8669,N_5882,N_6266);
or U8670 (N_8670,N_6427,N_5600);
nor U8671 (N_8671,N_5219,N_5908);
nor U8672 (N_8672,N_6023,N_5063);
nand U8673 (N_8673,N_5096,N_5779);
xnor U8674 (N_8674,N_5194,N_5227);
nand U8675 (N_8675,N_7456,N_6181);
xor U8676 (N_8676,N_6976,N_5523);
and U8677 (N_8677,N_6029,N_7120);
xnor U8678 (N_8678,N_5714,N_6078);
nor U8679 (N_8679,N_5558,N_7160);
nand U8680 (N_8680,N_6430,N_7435);
xnor U8681 (N_8681,N_7389,N_6771);
or U8682 (N_8682,N_5139,N_5421);
and U8683 (N_8683,N_6864,N_5387);
xnor U8684 (N_8684,N_5450,N_7061);
or U8685 (N_8685,N_6945,N_7197);
or U8686 (N_8686,N_6884,N_5588);
nor U8687 (N_8687,N_6677,N_6890);
and U8688 (N_8688,N_6217,N_7404);
or U8689 (N_8689,N_7098,N_6600);
and U8690 (N_8690,N_5979,N_5041);
xor U8691 (N_8691,N_6057,N_6104);
nor U8692 (N_8692,N_5446,N_6479);
or U8693 (N_8693,N_5546,N_6568);
xnor U8694 (N_8694,N_7174,N_6491);
and U8695 (N_8695,N_6436,N_6810);
xnor U8696 (N_8696,N_6284,N_7447);
xnor U8697 (N_8697,N_6475,N_6816);
nor U8698 (N_8698,N_6950,N_6100);
nor U8699 (N_8699,N_6277,N_6134);
nand U8700 (N_8700,N_6409,N_5551);
nand U8701 (N_8701,N_7421,N_5860);
nor U8702 (N_8702,N_7128,N_6641);
or U8703 (N_8703,N_6739,N_6338);
and U8704 (N_8704,N_5235,N_7176);
nand U8705 (N_8705,N_5968,N_5243);
xor U8706 (N_8706,N_6426,N_6517);
or U8707 (N_8707,N_6774,N_6131);
nand U8708 (N_8708,N_7322,N_6806);
xnor U8709 (N_8709,N_6183,N_7129);
nor U8710 (N_8710,N_7072,N_5876);
or U8711 (N_8711,N_7253,N_7165);
and U8712 (N_8712,N_5415,N_6132);
xnor U8713 (N_8713,N_5175,N_5727);
xor U8714 (N_8714,N_5700,N_6999);
and U8715 (N_8715,N_5712,N_6274);
nand U8716 (N_8716,N_6610,N_6316);
xor U8717 (N_8717,N_5106,N_6069);
or U8718 (N_8718,N_5613,N_6791);
or U8719 (N_8719,N_5378,N_5344);
xnor U8720 (N_8720,N_6281,N_5582);
and U8721 (N_8721,N_6026,N_6306);
or U8722 (N_8722,N_5409,N_7068);
nor U8723 (N_8723,N_5301,N_7281);
nor U8724 (N_8724,N_5786,N_7099);
and U8725 (N_8725,N_5599,N_6519);
and U8726 (N_8726,N_6948,N_5249);
xor U8727 (N_8727,N_5273,N_5060);
or U8728 (N_8728,N_6337,N_5438);
nor U8729 (N_8729,N_7346,N_7436);
nand U8730 (N_8730,N_6846,N_6943);
nand U8731 (N_8731,N_6861,N_7345);
and U8732 (N_8732,N_6124,N_6833);
or U8733 (N_8733,N_5331,N_5953);
or U8734 (N_8734,N_5927,N_7336);
nand U8735 (N_8735,N_7307,N_5677);
xor U8736 (N_8736,N_6372,N_5971);
nand U8737 (N_8737,N_7124,N_7491);
xor U8738 (N_8738,N_7039,N_5470);
nor U8739 (N_8739,N_5553,N_5255);
nor U8740 (N_8740,N_6052,N_7092);
xor U8741 (N_8741,N_5441,N_6544);
xnor U8742 (N_8742,N_6223,N_5343);
or U8743 (N_8743,N_5389,N_5991);
and U8744 (N_8744,N_6351,N_5419);
or U8745 (N_8745,N_7469,N_6062);
nor U8746 (N_8746,N_5315,N_6906);
nand U8747 (N_8747,N_5161,N_7192);
xnor U8748 (N_8748,N_6371,N_5920);
and U8749 (N_8749,N_5383,N_6594);
xor U8750 (N_8750,N_7360,N_6344);
and U8751 (N_8751,N_5229,N_6726);
nand U8752 (N_8752,N_6904,N_5813);
or U8753 (N_8753,N_7255,N_5262);
xor U8754 (N_8754,N_5694,N_5752);
nand U8755 (N_8755,N_5146,N_6279);
or U8756 (N_8756,N_5154,N_5128);
or U8757 (N_8757,N_6272,N_7472);
and U8758 (N_8758,N_5624,N_5312);
xnor U8759 (N_8759,N_6119,N_5159);
xor U8760 (N_8760,N_5097,N_5321);
or U8761 (N_8761,N_7275,N_6041);
nor U8762 (N_8762,N_6255,N_7280);
xor U8763 (N_8763,N_5855,N_5646);
nand U8764 (N_8764,N_5737,N_7342);
or U8765 (N_8765,N_7243,N_6934);
xor U8766 (N_8766,N_6354,N_6029);
or U8767 (N_8767,N_7490,N_6134);
nor U8768 (N_8768,N_7132,N_7456);
nor U8769 (N_8769,N_6922,N_6283);
xnor U8770 (N_8770,N_5114,N_5614);
xnor U8771 (N_8771,N_5658,N_6329);
and U8772 (N_8772,N_6411,N_7147);
nand U8773 (N_8773,N_6836,N_6533);
or U8774 (N_8774,N_6146,N_6068);
nand U8775 (N_8775,N_5451,N_6146);
xnor U8776 (N_8776,N_7497,N_7258);
or U8777 (N_8777,N_7497,N_5256);
or U8778 (N_8778,N_7306,N_5641);
nor U8779 (N_8779,N_5909,N_5955);
nand U8780 (N_8780,N_7353,N_5993);
or U8781 (N_8781,N_5813,N_6502);
nand U8782 (N_8782,N_6962,N_6333);
and U8783 (N_8783,N_5148,N_5198);
or U8784 (N_8784,N_6655,N_5857);
or U8785 (N_8785,N_5052,N_5835);
nor U8786 (N_8786,N_5476,N_6525);
or U8787 (N_8787,N_6528,N_6859);
nand U8788 (N_8788,N_7270,N_5980);
and U8789 (N_8789,N_7199,N_7222);
and U8790 (N_8790,N_5138,N_7092);
or U8791 (N_8791,N_5422,N_5703);
and U8792 (N_8792,N_7200,N_7053);
xnor U8793 (N_8793,N_7317,N_5520);
and U8794 (N_8794,N_7293,N_5887);
xnor U8795 (N_8795,N_6659,N_6643);
nor U8796 (N_8796,N_5266,N_5894);
xnor U8797 (N_8797,N_7165,N_6387);
nand U8798 (N_8798,N_5488,N_5061);
nor U8799 (N_8799,N_7438,N_5319);
and U8800 (N_8800,N_5119,N_6349);
nor U8801 (N_8801,N_5048,N_6111);
nand U8802 (N_8802,N_6960,N_7428);
and U8803 (N_8803,N_5958,N_5326);
or U8804 (N_8804,N_7333,N_6860);
nor U8805 (N_8805,N_5797,N_5491);
or U8806 (N_8806,N_6477,N_5499);
and U8807 (N_8807,N_5796,N_5527);
nor U8808 (N_8808,N_6571,N_6330);
xor U8809 (N_8809,N_6826,N_7463);
xnor U8810 (N_8810,N_5532,N_6624);
and U8811 (N_8811,N_5008,N_7072);
nor U8812 (N_8812,N_6743,N_6411);
nor U8813 (N_8813,N_5082,N_5156);
or U8814 (N_8814,N_5727,N_6454);
xor U8815 (N_8815,N_6528,N_5210);
xnor U8816 (N_8816,N_5002,N_6140);
xnor U8817 (N_8817,N_5982,N_6093);
xor U8818 (N_8818,N_6171,N_5103);
and U8819 (N_8819,N_5869,N_7488);
xnor U8820 (N_8820,N_5498,N_6265);
nor U8821 (N_8821,N_6484,N_6471);
xor U8822 (N_8822,N_5893,N_5757);
xor U8823 (N_8823,N_5995,N_6760);
nor U8824 (N_8824,N_5534,N_7243);
or U8825 (N_8825,N_7309,N_5472);
or U8826 (N_8826,N_5312,N_6485);
and U8827 (N_8827,N_5160,N_5941);
xor U8828 (N_8828,N_6058,N_6471);
nand U8829 (N_8829,N_5454,N_5274);
nand U8830 (N_8830,N_5742,N_5590);
nand U8831 (N_8831,N_5899,N_7102);
or U8832 (N_8832,N_5467,N_7399);
nor U8833 (N_8833,N_5400,N_6740);
nor U8834 (N_8834,N_5965,N_5372);
xor U8835 (N_8835,N_5475,N_5924);
xor U8836 (N_8836,N_7213,N_6718);
and U8837 (N_8837,N_6294,N_5150);
and U8838 (N_8838,N_6692,N_7421);
and U8839 (N_8839,N_5126,N_6989);
nor U8840 (N_8840,N_6942,N_7449);
or U8841 (N_8841,N_7037,N_6820);
and U8842 (N_8842,N_7035,N_7190);
nand U8843 (N_8843,N_6039,N_7491);
and U8844 (N_8844,N_6760,N_5589);
or U8845 (N_8845,N_6143,N_6695);
nor U8846 (N_8846,N_7065,N_5595);
xnor U8847 (N_8847,N_6784,N_5249);
and U8848 (N_8848,N_6010,N_5134);
xnor U8849 (N_8849,N_7197,N_7287);
and U8850 (N_8850,N_6419,N_7487);
xnor U8851 (N_8851,N_5009,N_7351);
nand U8852 (N_8852,N_6701,N_5382);
and U8853 (N_8853,N_6923,N_6236);
nor U8854 (N_8854,N_6003,N_5168);
and U8855 (N_8855,N_7436,N_6661);
nand U8856 (N_8856,N_7161,N_7127);
or U8857 (N_8857,N_6256,N_5159);
nor U8858 (N_8858,N_5755,N_7456);
and U8859 (N_8859,N_5505,N_5759);
and U8860 (N_8860,N_5915,N_5660);
and U8861 (N_8861,N_6945,N_6295);
xnor U8862 (N_8862,N_5706,N_6030);
xor U8863 (N_8863,N_6474,N_6850);
xor U8864 (N_8864,N_5653,N_6172);
nor U8865 (N_8865,N_7344,N_6665);
or U8866 (N_8866,N_5359,N_5705);
nand U8867 (N_8867,N_7059,N_5774);
or U8868 (N_8868,N_5825,N_5440);
nand U8869 (N_8869,N_6257,N_5438);
nand U8870 (N_8870,N_5911,N_6158);
and U8871 (N_8871,N_5975,N_5370);
xnor U8872 (N_8872,N_5874,N_7096);
xnor U8873 (N_8873,N_5621,N_6055);
or U8874 (N_8874,N_6886,N_5259);
nand U8875 (N_8875,N_7343,N_5575);
xor U8876 (N_8876,N_6049,N_7384);
nand U8877 (N_8877,N_7040,N_5581);
and U8878 (N_8878,N_5588,N_5595);
nand U8879 (N_8879,N_6018,N_5572);
xnor U8880 (N_8880,N_6356,N_5916);
nor U8881 (N_8881,N_5595,N_7045);
xor U8882 (N_8882,N_6267,N_5807);
nand U8883 (N_8883,N_5956,N_6182);
xor U8884 (N_8884,N_6841,N_6831);
nor U8885 (N_8885,N_7201,N_6148);
xor U8886 (N_8886,N_6157,N_5638);
nor U8887 (N_8887,N_6714,N_5297);
or U8888 (N_8888,N_6109,N_5520);
xnor U8889 (N_8889,N_6196,N_5711);
nand U8890 (N_8890,N_6607,N_5991);
xor U8891 (N_8891,N_5885,N_5990);
xnor U8892 (N_8892,N_6809,N_6269);
nor U8893 (N_8893,N_7257,N_5921);
nor U8894 (N_8894,N_7088,N_7231);
and U8895 (N_8895,N_7478,N_6032);
xor U8896 (N_8896,N_7475,N_5051);
xnor U8897 (N_8897,N_7164,N_6480);
xor U8898 (N_8898,N_6413,N_7031);
nand U8899 (N_8899,N_6714,N_5273);
or U8900 (N_8900,N_5839,N_6110);
nand U8901 (N_8901,N_7079,N_5672);
xnor U8902 (N_8902,N_6045,N_6884);
nand U8903 (N_8903,N_6732,N_5543);
nand U8904 (N_8904,N_5695,N_5204);
and U8905 (N_8905,N_6129,N_6096);
nand U8906 (N_8906,N_5613,N_5800);
nor U8907 (N_8907,N_7126,N_5435);
and U8908 (N_8908,N_6356,N_6739);
nand U8909 (N_8909,N_6619,N_6632);
nand U8910 (N_8910,N_7103,N_5871);
nand U8911 (N_8911,N_7044,N_5316);
nand U8912 (N_8912,N_5028,N_5564);
or U8913 (N_8913,N_5057,N_5654);
or U8914 (N_8914,N_6668,N_5209);
nor U8915 (N_8915,N_7487,N_5306);
nand U8916 (N_8916,N_6133,N_5224);
xnor U8917 (N_8917,N_6671,N_7076);
xor U8918 (N_8918,N_6777,N_5122);
and U8919 (N_8919,N_6496,N_5429);
and U8920 (N_8920,N_5010,N_5999);
nand U8921 (N_8921,N_6654,N_7252);
xor U8922 (N_8922,N_7150,N_6571);
xnor U8923 (N_8923,N_7373,N_5565);
xor U8924 (N_8924,N_5201,N_6826);
or U8925 (N_8925,N_6114,N_7159);
and U8926 (N_8926,N_5396,N_7213);
xnor U8927 (N_8927,N_6105,N_5414);
xor U8928 (N_8928,N_7151,N_7024);
xor U8929 (N_8929,N_5320,N_5802);
nor U8930 (N_8930,N_7439,N_6085);
nand U8931 (N_8931,N_7121,N_6584);
and U8932 (N_8932,N_5274,N_7431);
nand U8933 (N_8933,N_6930,N_5768);
nand U8934 (N_8934,N_7331,N_5048);
xnor U8935 (N_8935,N_6892,N_7001);
nor U8936 (N_8936,N_6821,N_5516);
xnor U8937 (N_8937,N_5603,N_7147);
nand U8938 (N_8938,N_6399,N_7493);
or U8939 (N_8939,N_7237,N_6724);
or U8940 (N_8940,N_5492,N_6251);
nand U8941 (N_8941,N_7057,N_6374);
nor U8942 (N_8942,N_5941,N_5179);
and U8943 (N_8943,N_7269,N_7234);
nor U8944 (N_8944,N_5730,N_5590);
and U8945 (N_8945,N_6857,N_5599);
nand U8946 (N_8946,N_5602,N_6692);
and U8947 (N_8947,N_6499,N_7434);
and U8948 (N_8948,N_6949,N_6762);
and U8949 (N_8949,N_6696,N_7279);
nand U8950 (N_8950,N_6987,N_7293);
nand U8951 (N_8951,N_5675,N_5776);
or U8952 (N_8952,N_5576,N_5349);
or U8953 (N_8953,N_5931,N_7086);
and U8954 (N_8954,N_5584,N_5232);
or U8955 (N_8955,N_5091,N_6075);
nand U8956 (N_8956,N_6133,N_5417);
nor U8957 (N_8957,N_6178,N_6690);
nor U8958 (N_8958,N_6516,N_6926);
nor U8959 (N_8959,N_6827,N_6006);
nand U8960 (N_8960,N_5783,N_5056);
or U8961 (N_8961,N_5159,N_5166);
and U8962 (N_8962,N_6643,N_6232);
or U8963 (N_8963,N_6674,N_6590);
and U8964 (N_8964,N_5886,N_6565);
or U8965 (N_8965,N_5930,N_5291);
xnor U8966 (N_8966,N_5414,N_7186);
and U8967 (N_8967,N_5259,N_6126);
and U8968 (N_8968,N_5726,N_7423);
or U8969 (N_8969,N_6169,N_5066);
nand U8970 (N_8970,N_5473,N_5450);
nand U8971 (N_8971,N_6259,N_6703);
xnor U8972 (N_8972,N_7455,N_5887);
and U8973 (N_8973,N_5350,N_6126);
or U8974 (N_8974,N_5394,N_5161);
or U8975 (N_8975,N_5451,N_7224);
nand U8976 (N_8976,N_6222,N_6183);
nand U8977 (N_8977,N_6894,N_5873);
nor U8978 (N_8978,N_5148,N_5924);
xnor U8979 (N_8979,N_7229,N_6670);
xnor U8980 (N_8980,N_5836,N_5365);
or U8981 (N_8981,N_6715,N_5927);
or U8982 (N_8982,N_6327,N_7110);
nand U8983 (N_8983,N_5802,N_5089);
nor U8984 (N_8984,N_5126,N_6808);
or U8985 (N_8985,N_7499,N_7297);
nor U8986 (N_8986,N_5522,N_7401);
xnor U8987 (N_8987,N_6535,N_5895);
nor U8988 (N_8988,N_6856,N_6093);
and U8989 (N_8989,N_5748,N_5006);
nor U8990 (N_8990,N_5633,N_6971);
or U8991 (N_8991,N_5087,N_7280);
xor U8992 (N_8992,N_6728,N_6771);
nor U8993 (N_8993,N_6008,N_6187);
or U8994 (N_8994,N_6206,N_6292);
nor U8995 (N_8995,N_5701,N_6412);
nor U8996 (N_8996,N_5940,N_6823);
or U8997 (N_8997,N_6643,N_5393);
or U8998 (N_8998,N_6006,N_5854);
and U8999 (N_8999,N_5809,N_5263);
xor U9000 (N_9000,N_7104,N_6376);
or U9001 (N_9001,N_5737,N_6237);
or U9002 (N_9002,N_6134,N_7073);
xor U9003 (N_9003,N_6865,N_5950);
and U9004 (N_9004,N_5201,N_5485);
nand U9005 (N_9005,N_6681,N_5275);
nand U9006 (N_9006,N_5581,N_7119);
nand U9007 (N_9007,N_5673,N_5023);
and U9008 (N_9008,N_5045,N_5956);
xnor U9009 (N_9009,N_6479,N_5928);
or U9010 (N_9010,N_5583,N_5209);
or U9011 (N_9011,N_5100,N_5145);
nand U9012 (N_9012,N_7183,N_6294);
xor U9013 (N_9013,N_7402,N_5964);
or U9014 (N_9014,N_6493,N_7021);
nand U9015 (N_9015,N_5927,N_5742);
and U9016 (N_9016,N_7242,N_6145);
or U9017 (N_9017,N_5383,N_5774);
or U9018 (N_9018,N_6602,N_5042);
and U9019 (N_9019,N_6077,N_5417);
and U9020 (N_9020,N_6983,N_5865);
or U9021 (N_9021,N_6618,N_5448);
xor U9022 (N_9022,N_5430,N_7265);
xnor U9023 (N_9023,N_5723,N_5926);
nand U9024 (N_9024,N_5284,N_6433);
nor U9025 (N_9025,N_5602,N_6793);
nand U9026 (N_9026,N_6025,N_7134);
xnor U9027 (N_9027,N_6695,N_5935);
xnor U9028 (N_9028,N_6346,N_6974);
xor U9029 (N_9029,N_6772,N_6123);
nand U9030 (N_9030,N_6550,N_7122);
and U9031 (N_9031,N_7169,N_6324);
nor U9032 (N_9032,N_7498,N_7275);
nor U9033 (N_9033,N_6807,N_7426);
and U9034 (N_9034,N_6270,N_6126);
and U9035 (N_9035,N_6633,N_5349);
nor U9036 (N_9036,N_6599,N_5938);
xnor U9037 (N_9037,N_6951,N_7037);
nor U9038 (N_9038,N_6108,N_5164);
and U9039 (N_9039,N_6238,N_6337);
or U9040 (N_9040,N_6309,N_6761);
or U9041 (N_9041,N_5876,N_7041);
xnor U9042 (N_9042,N_6826,N_6022);
or U9043 (N_9043,N_5573,N_6432);
nand U9044 (N_9044,N_6288,N_5337);
xnor U9045 (N_9045,N_5680,N_6646);
or U9046 (N_9046,N_7163,N_5685);
and U9047 (N_9047,N_5048,N_5825);
nor U9048 (N_9048,N_5815,N_6993);
xnor U9049 (N_9049,N_5070,N_5277);
nand U9050 (N_9050,N_5738,N_6931);
xnor U9051 (N_9051,N_6479,N_5198);
or U9052 (N_9052,N_7235,N_6158);
and U9053 (N_9053,N_6296,N_6640);
nor U9054 (N_9054,N_7488,N_7129);
or U9055 (N_9055,N_5725,N_6509);
xnor U9056 (N_9056,N_5394,N_5374);
xnor U9057 (N_9057,N_6400,N_5794);
xor U9058 (N_9058,N_5980,N_6934);
nor U9059 (N_9059,N_6765,N_5557);
xnor U9060 (N_9060,N_6900,N_5016);
and U9061 (N_9061,N_7497,N_5228);
nor U9062 (N_9062,N_6331,N_7250);
and U9063 (N_9063,N_5714,N_5363);
or U9064 (N_9064,N_6252,N_7342);
nand U9065 (N_9065,N_6325,N_6376);
nor U9066 (N_9066,N_6861,N_6239);
and U9067 (N_9067,N_5484,N_5086);
nand U9068 (N_9068,N_7463,N_7445);
and U9069 (N_9069,N_5906,N_5974);
and U9070 (N_9070,N_5420,N_6123);
or U9071 (N_9071,N_5298,N_6498);
or U9072 (N_9072,N_6233,N_6729);
xor U9073 (N_9073,N_6545,N_6422);
nor U9074 (N_9074,N_5402,N_7309);
nand U9075 (N_9075,N_6233,N_6188);
xnor U9076 (N_9076,N_5930,N_6448);
xnor U9077 (N_9077,N_6295,N_6436);
or U9078 (N_9078,N_6736,N_6876);
and U9079 (N_9079,N_5448,N_5115);
xnor U9080 (N_9080,N_7036,N_7094);
and U9081 (N_9081,N_6096,N_5233);
xor U9082 (N_9082,N_5488,N_5163);
and U9083 (N_9083,N_7041,N_6504);
xnor U9084 (N_9084,N_6084,N_5781);
xor U9085 (N_9085,N_6605,N_6004);
and U9086 (N_9086,N_5463,N_6189);
and U9087 (N_9087,N_5367,N_5517);
nor U9088 (N_9088,N_6713,N_5250);
and U9089 (N_9089,N_6280,N_6108);
and U9090 (N_9090,N_6279,N_6462);
or U9091 (N_9091,N_5619,N_6519);
or U9092 (N_9092,N_5983,N_7405);
xnor U9093 (N_9093,N_6035,N_5202);
xnor U9094 (N_9094,N_5700,N_7198);
nor U9095 (N_9095,N_5558,N_6833);
and U9096 (N_9096,N_5017,N_7014);
nor U9097 (N_9097,N_7436,N_6853);
xnor U9098 (N_9098,N_6496,N_5439);
xnor U9099 (N_9099,N_5068,N_5713);
xnor U9100 (N_9100,N_7001,N_5505);
and U9101 (N_9101,N_7201,N_5075);
and U9102 (N_9102,N_5133,N_5762);
or U9103 (N_9103,N_7085,N_7274);
xor U9104 (N_9104,N_5103,N_5864);
nand U9105 (N_9105,N_5663,N_7133);
nand U9106 (N_9106,N_7440,N_5507);
and U9107 (N_9107,N_6672,N_6970);
and U9108 (N_9108,N_6297,N_5173);
nand U9109 (N_9109,N_5254,N_7354);
xnor U9110 (N_9110,N_7308,N_7043);
and U9111 (N_9111,N_6918,N_6904);
and U9112 (N_9112,N_5781,N_5360);
and U9113 (N_9113,N_5876,N_7212);
xnor U9114 (N_9114,N_6379,N_6098);
xor U9115 (N_9115,N_6706,N_6271);
or U9116 (N_9116,N_5835,N_6914);
nand U9117 (N_9117,N_6291,N_7355);
nand U9118 (N_9118,N_7100,N_5949);
nor U9119 (N_9119,N_5518,N_6979);
and U9120 (N_9120,N_6452,N_7480);
or U9121 (N_9121,N_5879,N_5731);
and U9122 (N_9122,N_6240,N_5137);
and U9123 (N_9123,N_6846,N_6121);
and U9124 (N_9124,N_6412,N_5316);
nor U9125 (N_9125,N_6234,N_6466);
nor U9126 (N_9126,N_5667,N_6368);
xor U9127 (N_9127,N_7355,N_5616);
and U9128 (N_9128,N_7158,N_6129);
nand U9129 (N_9129,N_5342,N_6243);
nand U9130 (N_9130,N_7455,N_7494);
nor U9131 (N_9131,N_5279,N_6164);
xor U9132 (N_9132,N_5135,N_5768);
nand U9133 (N_9133,N_7321,N_5392);
nor U9134 (N_9134,N_7403,N_7260);
xnor U9135 (N_9135,N_5612,N_6223);
or U9136 (N_9136,N_7482,N_5058);
nor U9137 (N_9137,N_7154,N_7360);
and U9138 (N_9138,N_5407,N_6916);
or U9139 (N_9139,N_6053,N_6701);
and U9140 (N_9140,N_6855,N_5303);
nor U9141 (N_9141,N_5312,N_5378);
xnor U9142 (N_9142,N_6483,N_5182);
nand U9143 (N_9143,N_5168,N_6965);
nor U9144 (N_9144,N_6146,N_6918);
nor U9145 (N_9145,N_7082,N_7145);
and U9146 (N_9146,N_5125,N_6585);
or U9147 (N_9147,N_6363,N_7151);
nand U9148 (N_9148,N_6974,N_6120);
xnor U9149 (N_9149,N_6143,N_5858);
nor U9150 (N_9150,N_7058,N_5399);
nand U9151 (N_9151,N_5885,N_5913);
xnor U9152 (N_9152,N_5986,N_6455);
nor U9153 (N_9153,N_6884,N_5876);
and U9154 (N_9154,N_7085,N_7069);
nor U9155 (N_9155,N_5495,N_5236);
nor U9156 (N_9156,N_5987,N_5508);
xnor U9157 (N_9157,N_5195,N_5866);
nor U9158 (N_9158,N_7222,N_6080);
nor U9159 (N_9159,N_7448,N_6081);
nor U9160 (N_9160,N_6613,N_7045);
xnor U9161 (N_9161,N_7264,N_5113);
nor U9162 (N_9162,N_5049,N_5174);
nor U9163 (N_9163,N_5739,N_5873);
and U9164 (N_9164,N_6679,N_7314);
nand U9165 (N_9165,N_5900,N_5363);
and U9166 (N_9166,N_6111,N_6620);
and U9167 (N_9167,N_6749,N_6341);
and U9168 (N_9168,N_5057,N_6527);
nor U9169 (N_9169,N_5515,N_6184);
nor U9170 (N_9170,N_5632,N_6975);
or U9171 (N_9171,N_6687,N_5473);
or U9172 (N_9172,N_5514,N_6063);
nand U9173 (N_9173,N_5722,N_5122);
and U9174 (N_9174,N_5291,N_5942);
and U9175 (N_9175,N_6213,N_5741);
or U9176 (N_9176,N_6306,N_6428);
nor U9177 (N_9177,N_7494,N_5999);
nor U9178 (N_9178,N_5538,N_5796);
nor U9179 (N_9179,N_6021,N_7044);
nor U9180 (N_9180,N_7287,N_5075);
nor U9181 (N_9181,N_5266,N_7463);
nand U9182 (N_9182,N_5112,N_7498);
and U9183 (N_9183,N_7153,N_5684);
or U9184 (N_9184,N_5723,N_7152);
nand U9185 (N_9185,N_6479,N_5017);
and U9186 (N_9186,N_7140,N_5158);
nand U9187 (N_9187,N_6436,N_6958);
or U9188 (N_9188,N_6633,N_5593);
nand U9189 (N_9189,N_6454,N_5913);
nand U9190 (N_9190,N_6610,N_6667);
nor U9191 (N_9191,N_5239,N_6699);
nor U9192 (N_9192,N_5850,N_7088);
and U9193 (N_9193,N_7405,N_5125);
nor U9194 (N_9194,N_5912,N_5134);
nand U9195 (N_9195,N_5970,N_6105);
or U9196 (N_9196,N_6439,N_5444);
nor U9197 (N_9197,N_5762,N_5888);
xnor U9198 (N_9198,N_7392,N_6806);
xor U9199 (N_9199,N_6692,N_5669);
xnor U9200 (N_9200,N_6768,N_6307);
nor U9201 (N_9201,N_6419,N_5097);
and U9202 (N_9202,N_7215,N_5734);
nand U9203 (N_9203,N_5315,N_7095);
nand U9204 (N_9204,N_5296,N_5847);
or U9205 (N_9205,N_5783,N_5424);
nor U9206 (N_9206,N_5414,N_5032);
nand U9207 (N_9207,N_6848,N_7262);
xnor U9208 (N_9208,N_5282,N_5553);
nand U9209 (N_9209,N_7461,N_7349);
and U9210 (N_9210,N_5413,N_5660);
xor U9211 (N_9211,N_7288,N_7317);
nor U9212 (N_9212,N_6528,N_6280);
or U9213 (N_9213,N_5331,N_6346);
xor U9214 (N_9214,N_7423,N_5337);
nand U9215 (N_9215,N_6375,N_6357);
and U9216 (N_9216,N_6540,N_6805);
nor U9217 (N_9217,N_6484,N_6569);
nand U9218 (N_9218,N_6414,N_6328);
nor U9219 (N_9219,N_5364,N_7215);
and U9220 (N_9220,N_6949,N_7335);
nor U9221 (N_9221,N_5394,N_6261);
nor U9222 (N_9222,N_5211,N_5052);
nand U9223 (N_9223,N_6283,N_5911);
xnor U9224 (N_9224,N_6862,N_6080);
and U9225 (N_9225,N_5515,N_6666);
nor U9226 (N_9226,N_5280,N_6864);
xnor U9227 (N_9227,N_5533,N_5092);
or U9228 (N_9228,N_5106,N_6662);
nand U9229 (N_9229,N_6280,N_6393);
nand U9230 (N_9230,N_5153,N_5782);
nand U9231 (N_9231,N_6616,N_5825);
xor U9232 (N_9232,N_6153,N_7119);
nand U9233 (N_9233,N_7298,N_6232);
nand U9234 (N_9234,N_6730,N_5109);
nand U9235 (N_9235,N_5836,N_6972);
xor U9236 (N_9236,N_6539,N_6669);
and U9237 (N_9237,N_6998,N_7405);
or U9238 (N_9238,N_6032,N_5068);
and U9239 (N_9239,N_5090,N_6853);
nand U9240 (N_9240,N_5937,N_7373);
xor U9241 (N_9241,N_5663,N_6774);
nand U9242 (N_9242,N_7178,N_6233);
or U9243 (N_9243,N_5423,N_5510);
nor U9244 (N_9244,N_7274,N_7050);
and U9245 (N_9245,N_5469,N_5782);
nand U9246 (N_9246,N_6525,N_5021);
xor U9247 (N_9247,N_6610,N_6249);
xor U9248 (N_9248,N_6897,N_5774);
nand U9249 (N_9249,N_6914,N_5594);
and U9250 (N_9250,N_6371,N_5727);
and U9251 (N_9251,N_5545,N_5863);
nor U9252 (N_9252,N_5721,N_5208);
nand U9253 (N_9253,N_6150,N_5992);
and U9254 (N_9254,N_5175,N_5570);
and U9255 (N_9255,N_6233,N_6241);
nor U9256 (N_9256,N_6658,N_5862);
nand U9257 (N_9257,N_5531,N_6915);
nor U9258 (N_9258,N_6720,N_6110);
and U9259 (N_9259,N_5173,N_5712);
nand U9260 (N_9260,N_6797,N_7150);
or U9261 (N_9261,N_6916,N_6846);
or U9262 (N_9262,N_5835,N_6515);
xor U9263 (N_9263,N_5269,N_5385);
nand U9264 (N_9264,N_6283,N_5291);
xnor U9265 (N_9265,N_5989,N_5169);
nand U9266 (N_9266,N_7261,N_7351);
xor U9267 (N_9267,N_7442,N_5087);
and U9268 (N_9268,N_5288,N_6597);
nor U9269 (N_9269,N_5463,N_5403);
and U9270 (N_9270,N_6962,N_5015);
nand U9271 (N_9271,N_5618,N_5210);
nand U9272 (N_9272,N_5211,N_6273);
nand U9273 (N_9273,N_6467,N_6465);
xor U9274 (N_9274,N_6283,N_6059);
or U9275 (N_9275,N_5416,N_7236);
nand U9276 (N_9276,N_6790,N_5732);
nand U9277 (N_9277,N_6321,N_6867);
nor U9278 (N_9278,N_5565,N_5517);
nand U9279 (N_9279,N_7284,N_5041);
or U9280 (N_9280,N_5568,N_5818);
or U9281 (N_9281,N_7481,N_7434);
nor U9282 (N_9282,N_7402,N_7085);
or U9283 (N_9283,N_6501,N_7013);
nor U9284 (N_9284,N_5140,N_6236);
nand U9285 (N_9285,N_5106,N_5033);
or U9286 (N_9286,N_6139,N_7341);
xor U9287 (N_9287,N_6924,N_6991);
nor U9288 (N_9288,N_6828,N_6317);
xor U9289 (N_9289,N_7387,N_7174);
xor U9290 (N_9290,N_5869,N_7039);
or U9291 (N_9291,N_7005,N_6737);
or U9292 (N_9292,N_5226,N_6627);
or U9293 (N_9293,N_6679,N_7191);
xnor U9294 (N_9294,N_6564,N_7338);
and U9295 (N_9295,N_6923,N_7265);
nand U9296 (N_9296,N_5323,N_6012);
nand U9297 (N_9297,N_6511,N_5345);
xor U9298 (N_9298,N_6063,N_6445);
nand U9299 (N_9299,N_7449,N_6643);
xnor U9300 (N_9300,N_5771,N_5156);
and U9301 (N_9301,N_6069,N_7345);
or U9302 (N_9302,N_7342,N_6715);
nand U9303 (N_9303,N_6465,N_5978);
xnor U9304 (N_9304,N_6238,N_5598);
nor U9305 (N_9305,N_6280,N_5389);
or U9306 (N_9306,N_5545,N_7005);
nor U9307 (N_9307,N_5897,N_7375);
nor U9308 (N_9308,N_6076,N_5943);
xor U9309 (N_9309,N_5187,N_7430);
nor U9310 (N_9310,N_6241,N_5479);
and U9311 (N_9311,N_6771,N_5091);
nor U9312 (N_9312,N_6152,N_5717);
nand U9313 (N_9313,N_7301,N_6005);
nand U9314 (N_9314,N_6678,N_6759);
xor U9315 (N_9315,N_5749,N_7092);
nand U9316 (N_9316,N_7358,N_6875);
and U9317 (N_9317,N_5575,N_6328);
nor U9318 (N_9318,N_5908,N_6642);
and U9319 (N_9319,N_6220,N_5485);
and U9320 (N_9320,N_7268,N_5491);
xor U9321 (N_9321,N_5397,N_7181);
xor U9322 (N_9322,N_6759,N_6150);
xor U9323 (N_9323,N_6464,N_5893);
nor U9324 (N_9324,N_7239,N_6401);
or U9325 (N_9325,N_5886,N_6048);
and U9326 (N_9326,N_6422,N_6075);
xnor U9327 (N_9327,N_6497,N_7195);
xnor U9328 (N_9328,N_6945,N_7307);
nand U9329 (N_9329,N_6634,N_6401);
xor U9330 (N_9330,N_6784,N_7115);
nand U9331 (N_9331,N_6470,N_5350);
nor U9332 (N_9332,N_6599,N_5730);
and U9333 (N_9333,N_7251,N_5380);
xnor U9334 (N_9334,N_5838,N_5670);
and U9335 (N_9335,N_7345,N_5853);
nand U9336 (N_9336,N_7019,N_5116);
xor U9337 (N_9337,N_5676,N_7260);
or U9338 (N_9338,N_6361,N_6292);
xor U9339 (N_9339,N_5761,N_5815);
or U9340 (N_9340,N_6218,N_6454);
or U9341 (N_9341,N_6031,N_5057);
nor U9342 (N_9342,N_5439,N_7424);
xnor U9343 (N_9343,N_5016,N_6809);
or U9344 (N_9344,N_5019,N_6626);
and U9345 (N_9345,N_7311,N_5412);
nor U9346 (N_9346,N_6643,N_6434);
or U9347 (N_9347,N_6957,N_5526);
or U9348 (N_9348,N_5403,N_7292);
nor U9349 (N_9349,N_5861,N_5164);
nor U9350 (N_9350,N_6376,N_6163);
xor U9351 (N_9351,N_5957,N_5733);
xor U9352 (N_9352,N_6596,N_7464);
and U9353 (N_9353,N_6044,N_5525);
or U9354 (N_9354,N_5485,N_5937);
nand U9355 (N_9355,N_6776,N_6386);
xor U9356 (N_9356,N_5660,N_5859);
or U9357 (N_9357,N_7132,N_7324);
xor U9358 (N_9358,N_7247,N_5033);
nand U9359 (N_9359,N_7458,N_6901);
and U9360 (N_9360,N_6301,N_5155);
nand U9361 (N_9361,N_5961,N_6722);
xor U9362 (N_9362,N_6067,N_6327);
nand U9363 (N_9363,N_6387,N_6475);
xnor U9364 (N_9364,N_6311,N_6722);
xor U9365 (N_9365,N_5837,N_5155);
or U9366 (N_9366,N_6560,N_7315);
and U9367 (N_9367,N_5232,N_7217);
nand U9368 (N_9368,N_6893,N_6245);
xor U9369 (N_9369,N_6786,N_6074);
nor U9370 (N_9370,N_7181,N_7187);
xor U9371 (N_9371,N_6056,N_6972);
nand U9372 (N_9372,N_5295,N_5978);
nand U9373 (N_9373,N_7292,N_7137);
and U9374 (N_9374,N_6155,N_7224);
and U9375 (N_9375,N_5624,N_6481);
nand U9376 (N_9376,N_5764,N_7227);
xor U9377 (N_9377,N_5508,N_6722);
nor U9378 (N_9378,N_5824,N_6469);
nor U9379 (N_9379,N_5971,N_6082);
nor U9380 (N_9380,N_7383,N_6651);
and U9381 (N_9381,N_7185,N_6192);
nand U9382 (N_9382,N_7052,N_7005);
and U9383 (N_9383,N_5399,N_6655);
nor U9384 (N_9384,N_5773,N_6322);
xnor U9385 (N_9385,N_6010,N_5856);
xnor U9386 (N_9386,N_7091,N_5950);
and U9387 (N_9387,N_6180,N_6329);
xnor U9388 (N_9388,N_7157,N_5601);
and U9389 (N_9389,N_5468,N_7087);
nand U9390 (N_9390,N_5562,N_5623);
xor U9391 (N_9391,N_5815,N_7462);
nor U9392 (N_9392,N_6249,N_5826);
nand U9393 (N_9393,N_6531,N_7107);
xor U9394 (N_9394,N_5628,N_5845);
or U9395 (N_9395,N_7388,N_7049);
and U9396 (N_9396,N_5116,N_5853);
or U9397 (N_9397,N_5632,N_6494);
xor U9398 (N_9398,N_5461,N_6983);
nand U9399 (N_9399,N_6585,N_5631);
and U9400 (N_9400,N_7044,N_7458);
and U9401 (N_9401,N_7432,N_6244);
nand U9402 (N_9402,N_6754,N_6006);
nand U9403 (N_9403,N_6461,N_6704);
nand U9404 (N_9404,N_6283,N_6604);
xor U9405 (N_9405,N_6948,N_6979);
and U9406 (N_9406,N_7118,N_6449);
or U9407 (N_9407,N_5159,N_6088);
and U9408 (N_9408,N_5969,N_7244);
xor U9409 (N_9409,N_5650,N_5764);
or U9410 (N_9410,N_7194,N_6886);
xnor U9411 (N_9411,N_5582,N_5160);
nand U9412 (N_9412,N_5385,N_6133);
nor U9413 (N_9413,N_6424,N_5807);
nand U9414 (N_9414,N_6783,N_6570);
or U9415 (N_9415,N_5810,N_6621);
xnor U9416 (N_9416,N_5193,N_6002);
nand U9417 (N_9417,N_7297,N_5609);
nand U9418 (N_9418,N_5859,N_5279);
xnor U9419 (N_9419,N_5673,N_6988);
xor U9420 (N_9420,N_7139,N_7000);
or U9421 (N_9421,N_6075,N_6353);
nor U9422 (N_9422,N_7131,N_5742);
or U9423 (N_9423,N_5566,N_5147);
or U9424 (N_9424,N_7305,N_5119);
nor U9425 (N_9425,N_5602,N_6404);
nor U9426 (N_9426,N_5895,N_5005);
and U9427 (N_9427,N_5771,N_5817);
nor U9428 (N_9428,N_7190,N_5348);
xnor U9429 (N_9429,N_7424,N_5723);
and U9430 (N_9430,N_6935,N_5417);
nand U9431 (N_9431,N_7358,N_5640);
xnor U9432 (N_9432,N_5008,N_5158);
nor U9433 (N_9433,N_6352,N_7485);
nor U9434 (N_9434,N_6779,N_7289);
xor U9435 (N_9435,N_6553,N_6619);
xnor U9436 (N_9436,N_7443,N_7054);
xnor U9437 (N_9437,N_5985,N_7008);
and U9438 (N_9438,N_5144,N_6115);
and U9439 (N_9439,N_6833,N_5384);
and U9440 (N_9440,N_6897,N_7301);
or U9441 (N_9441,N_6927,N_5794);
and U9442 (N_9442,N_5542,N_5475);
nor U9443 (N_9443,N_5149,N_5742);
nor U9444 (N_9444,N_6116,N_5976);
nand U9445 (N_9445,N_5164,N_5191);
and U9446 (N_9446,N_6312,N_7251);
xnor U9447 (N_9447,N_7278,N_6340);
and U9448 (N_9448,N_5414,N_5520);
or U9449 (N_9449,N_6798,N_5613);
xnor U9450 (N_9450,N_6504,N_6758);
xor U9451 (N_9451,N_6443,N_6750);
and U9452 (N_9452,N_6121,N_5922);
and U9453 (N_9453,N_6629,N_7390);
xnor U9454 (N_9454,N_7277,N_5313);
and U9455 (N_9455,N_7196,N_7094);
nand U9456 (N_9456,N_5669,N_5166);
or U9457 (N_9457,N_5066,N_5171);
nor U9458 (N_9458,N_5323,N_5047);
or U9459 (N_9459,N_6857,N_7030);
and U9460 (N_9460,N_7401,N_5961);
or U9461 (N_9461,N_5331,N_6140);
and U9462 (N_9462,N_5239,N_6514);
and U9463 (N_9463,N_6956,N_5689);
nor U9464 (N_9464,N_7144,N_5742);
xnor U9465 (N_9465,N_5799,N_6536);
or U9466 (N_9466,N_6494,N_7350);
xor U9467 (N_9467,N_7416,N_6649);
xnor U9468 (N_9468,N_6249,N_5620);
nor U9469 (N_9469,N_6425,N_6494);
and U9470 (N_9470,N_5549,N_5480);
nor U9471 (N_9471,N_6738,N_6225);
xnor U9472 (N_9472,N_6218,N_5437);
nor U9473 (N_9473,N_5579,N_5263);
nand U9474 (N_9474,N_6717,N_6448);
xnor U9475 (N_9475,N_6001,N_5982);
xnor U9476 (N_9476,N_7432,N_7347);
and U9477 (N_9477,N_5068,N_6835);
or U9478 (N_9478,N_6544,N_6036);
nand U9479 (N_9479,N_6544,N_6549);
nor U9480 (N_9480,N_5746,N_5616);
nand U9481 (N_9481,N_7027,N_5513);
nor U9482 (N_9482,N_5511,N_6664);
or U9483 (N_9483,N_6453,N_6244);
and U9484 (N_9484,N_5647,N_6147);
nand U9485 (N_9485,N_6340,N_6675);
or U9486 (N_9486,N_6228,N_6989);
nor U9487 (N_9487,N_6543,N_6429);
and U9488 (N_9488,N_7070,N_5310);
nor U9489 (N_9489,N_5677,N_7174);
and U9490 (N_9490,N_5902,N_6541);
or U9491 (N_9491,N_7171,N_7499);
and U9492 (N_9492,N_5777,N_6142);
or U9493 (N_9493,N_6667,N_7315);
xor U9494 (N_9494,N_7125,N_5723);
and U9495 (N_9495,N_7286,N_5172);
xnor U9496 (N_9496,N_5555,N_7466);
xnor U9497 (N_9497,N_5978,N_7395);
or U9498 (N_9498,N_6655,N_5152);
nor U9499 (N_9499,N_5337,N_5785);
and U9500 (N_9500,N_6333,N_5758);
or U9501 (N_9501,N_6613,N_5896);
and U9502 (N_9502,N_6097,N_5589);
xor U9503 (N_9503,N_7033,N_6717);
and U9504 (N_9504,N_5704,N_7399);
nand U9505 (N_9505,N_5521,N_7085);
and U9506 (N_9506,N_6204,N_7376);
xor U9507 (N_9507,N_7466,N_5027);
and U9508 (N_9508,N_5268,N_5765);
and U9509 (N_9509,N_6671,N_6736);
nand U9510 (N_9510,N_7197,N_6216);
nor U9511 (N_9511,N_6459,N_5210);
nand U9512 (N_9512,N_6525,N_5781);
or U9513 (N_9513,N_6185,N_7181);
and U9514 (N_9514,N_6300,N_5355);
or U9515 (N_9515,N_6077,N_6797);
xnor U9516 (N_9516,N_5803,N_5076);
and U9517 (N_9517,N_6171,N_5634);
and U9518 (N_9518,N_5223,N_6837);
and U9519 (N_9519,N_7155,N_7065);
xor U9520 (N_9520,N_6411,N_6403);
xor U9521 (N_9521,N_5048,N_7198);
nand U9522 (N_9522,N_6663,N_6348);
and U9523 (N_9523,N_5124,N_5281);
and U9524 (N_9524,N_5147,N_6752);
or U9525 (N_9525,N_7283,N_5951);
and U9526 (N_9526,N_6240,N_5730);
and U9527 (N_9527,N_5607,N_5735);
nor U9528 (N_9528,N_6247,N_6657);
nand U9529 (N_9529,N_5878,N_6449);
xor U9530 (N_9530,N_6394,N_6981);
xor U9531 (N_9531,N_7040,N_6966);
and U9532 (N_9532,N_6110,N_5133);
xor U9533 (N_9533,N_6166,N_7281);
and U9534 (N_9534,N_5425,N_6144);
or U9535 (N_9535,N_6780,N_5474);
xor U9536 (N_9536,N_7340,N_6377);
xor U9537 (N_9537,N_5469,N_6256);
or U9538 (N_9538,N_5598,N_6572);
nor U9539 (N_9539,N_5600,N_7389);
xnor U9540 (N_9540,N_7410,N_6219);
xor U9541 (N_9541,N_6010,N_5674);
nor U9542 (N_9542,N_5350,N_7385);
nand U9543 (N_9543,N_7466,N_6294);
nor U9544 (N_9544,N_6044,N_7373);
and U9545 (N_9545,N_5226,N_6852);
and U9546 (N_9546,N_5694,N_6474);
nor U9547 (N_9547,N_7203,N_5945);
xor U9548 (N_9548,N_7124,N_5017);
and U9549 (N_9549,N_5786,N_6918);
and U9550 (N_9550,N_5656,N_5750);
nand U9551 (N_9551,N_5010,N_7488);
or U9552 (N_9552,N_5071,N_7425);
nand U9553 (N_9553,N_6548,N_7052);
nor U9554 (N_9554,N_6749,N_7170);
xor U9555 (N_9555,N_5084,N_6356);
xor U9556 (N_9556,N_7139,N_6697);
nand U9557 (N_9557,N_6964,N_7036);
xor U9558 (N_9558,N_6901,N_5998);
or U9559 (N_9559,N_7078,N_5420);
and U9560 (N_9560,N_5219,N_6916);
nor U9561 (N_9561,N_6858,N_5437);
and U9562 (N_9562,N_7207,N_5217);
and U9563 (N_9563,N_5475,N_7233);
nand U9564 (N_9564,N_7425,N_6122);
nand U9565 (N_9565,N_6432,N_7223);
or U9566 (N_9566,N_6763,N_5641);
and U9567 (N_9567,N_6091,N_6662);
nand U9568 (N_9568,N_5654,N_6006);
or U9569 (N_9569,N_6987,N_6215);
and U9570 (N_9570,N_6141,N_5896);
or U9571 (N_9571,N_5996,N_5965);
and U9572 (N_9572,N_6734,N_6690);
and U9573 (N_9573,N_6373,N_6126);
xnor U9574 (N_9574,N_7023,N_7219);
xor U9575 (N_9575,N_5360,N_6753);
nand U9576 (N_9576,N_6823,N_6255);
and U9577 (N_9577,N_5776,N_6228);
or U9578 (N_9578,N_6960,N_6859);
nor U9579 (N_9579,N_7239,N_7005);
or U9580 (N_9580,N_6937,N_5283);
or U9581 (N_9581,N_5661,N_5289);
xnor U9582 (N_9582,N_6996,N_6883);
xor U9583 (N_9583,N_6408,N_5841);
or U9584 (N_9584,N_5077,N_7387);
and U9585 (N_9585,N_7302,N_7212);
nand U9586 (N_9586,N_6175,N_7257);
nor U9587 (N_9587,N_5372,N_5775);
and U9588 (N_9588,N_6342,N_5196);
or U9589 (N_9589,N_5640,N_6004);
nand U9590 (N_9590,N_5084,N_5647);
and U9591 (N_9591,N_6993,N_7086);
or U9592 (N_9592,N_5734,N_6748);
nand U9593 (N_9593,N_5293,N_7015);
nor U9594 (N_9594,N_5490,N_5476);
and U9595 (N_9595,N_6453,N_5748);
xnor U9596 (N_9596,N_5966,N_5245);
or U9597 (N_9597,N_5297,N_7386);
or U9598 (N_9598,N_6539,N_5810);
xnor U9599 (N_9599,N_6649,N_6452);
nand U9600 (N_9600,N_5802,N_5496);
xnor U9601 (N_9601,N_6006,N_6175);
xnor U9602 (N_9602,N_6263,N_5589);
xor U9603 (N_9603,N_6177,N_6291);
or U9604 (N_9604,N_5812,N_5728);
or U9605 (N_9605,N_6197,N_5314);
nand U9606 (N_9606,N_5111,N_5747);
xnor U9607 (N_9607,N_6752,N_5521);
xor U9608 (N_9608,N_7252,N_5381);
nand U9609 (N_9609,N_6976,N_6196);
nor U9610 (N_9610,N_5531,N_6266);
and U9611 (N_9611,N_7351,N_6998);
and U9612 (N_9612,N_6057,N_5313);
nor U9613 (N_9613,N_5948,N_5191);
nor U9614 (N_9614,N_5827,N_5344);
and U9615 (N_9615,N_7384,N_6786);
xnor U9616 (N_9616,N_6442,N_6101);
nand U9617 (N_9617,N_6069,N_5868);
nand U9618 (N_9618,N_7092,N_5334);
nand U9619 (N_9619,N_6493,N_6678);
xnor U9620 (N_9620,N_5173,N_7036);
and U9621 (N_9621,N_5596,N_5052);
and U9622 (N_9622,N_7443,N_6488);
xor U9623 (N_9623,N_7259,N_6799);
nor U9624 (N_9624,N_6800,N_6975);
nand U9625 (N_9625,N_5805,N_6765);
and U9626 (N_9626,N_6306,N_6527);
or U9627 (N_9627,N_6880,N_5286);
and U9628 (N_9628,N_6621,N_7346);
nand U9629 (N_9629,N_6158,N_6535);
xnor U9630 (N_9630,N_6391,N_6354);
xor U9631 (N_9631,N_6709,N_6276);
or U9632 (N_9632,N_6484,N_6489);
and U9633 (N_9633,N_6875,N_5822);
nand U9634 (N_9634,N_7039,N_7175);
and U9635 (N_9635,N_6579,N_5476);
nor U9636 (N_9636,N_6487,N_6896);
and U9637 (N_9637,N_7248,N_6584);
xnor U9638 (N_9638,N_5979,N_5386);
xnor U9639 (N_9639,N_5598,N_5952);
xor U9640 (N_9640,N_5679,N_5376);
and U9641 (N_9641,N_7354,N_6010);
or U9642 (N_9642,N_5987,N_5202);
and U9643 (N_9643,N_6582,N_6831);
and U9644 (N_9644,N_5200,N_6302);
and U9645 (N_9645,N_6690,N_5224);
or U9646 (N_9646,N_7182,N_6561);
nor U9647 (N_9647,N_5883,N_7291);
or U9648 (N_9648,N_5639,N_5046);
and U9649 (N_9649,N_5886,N_7439);
and U9650 (N_9650,N_6811,N_5456);
and U9651 (N_9651,N_6232,N_6451);
and U9652 (N_9652,N_7152,N_7411);
and U9653 (N_9653,N_5506,N_5219);
and U9654 (N_9654,N_7408,N_5854);
or U9655 (N_9655,N_5413,N_5692);
nor U9656 (N_9656,N_6150,N_5335);
xnor U9657 (N_9657,N_6094,N_6589);
nor U9658 (N_9658,N_7154,N_6818);
and U9659 (N_9659,N_5545,N_5694);
nor U9660 (N_9660,N_5679,N_5280);
xnor U9661 (N_9661,N_5008,N_5763);
nand U9662 (N_9662,N_7472,N_7471);
and U9663 (N_9663,N_6004,N_5317);
xnor U9664 (N_9664,N_5902,N_5583);
xnor U9665 (N_9665,N_5044,N_6746);
and U9666 (N_9666,N_6233,N_5590);
and U9667 (N_9667,N_5414,N_5351);
or U9668 (N_9668,N_7353,N_5753);
and U9669 (N_9669,N_5686,N_5007);
nand U9670 (N_9670,N_5332,N_6992);
or U9671 (N_9671,N_5527,N_6031);
or U9672 (N_9672,N_5079,N_5518);
xnor U9673 (N_9673,N_6723,N_5342);
xnor U9674 (N_9674,N_7443,N_6360);
nor U9675 (N_9675,N_5792,N_5276);
nand U9676 (N_9676,N_5491,N_5589);
and U9677 (N_9677,N_5194,N_5447);
and U9678 (N_9678,N_6931,N_6234);
xnor U9679 (N_9679,N_6918,N_5065);
or U9680 (N_9680,N_6477,N_5968);
and U9681 (N_9681,N_6814,N_6253);
xnor U9682 (N_9682,N_5901,N_7386);
nor U9683 (N_9683,N_6962,N_6998);
and U9684 (N_9684,N_5341,N_5174);
xor U9685 (N_9685,N_7050,N_5196);
and U9686 (N_9686,N_7353,N_7333);
or U9687 (N_9687,N_6053,N_6441);
nand U9688 (N_9688,N_6078,N_6551);
nand U9689 (N_9689,N_5534,N_7448);
nand U9690 (N_9690,N_6070,N_7192);
nor U9691 (N_9691,N_6389,N_5832);
or U9692 (N_9692,N_7494,N_5823);
nand U9693 (N_9693,N_5313,N_6232);
xor U9694 (N_9694,N_7110,N_5628);
or U9695 (N_9695,N_6083,N_6717);
nor U9696 (N_9696,N_5379,N_5765);
nand U9697 (N_9697,N_7387,N_7118);
or U9698 (N_9698,N_6565,N_6610);
xnor U9699 (N_9699,N_6712,N_6083);
nand U9700 (N_9700,N_7369,N_6057);
nor U9701 (N_9701,N_5812,N_6554);
nand U9702 (N_9702,N_6131,N_6510);
and U9703 (N_9703,N_5367,N_7417);
and U9704 (N_9704,N_6177,N_7105);
and U9705 (N_9705,N_5497,N_7314);
nand U9706 (N_9706,N_7181,N_6608);
and U9707 (N_9707,N_7037,N_6585);
or U9708 (N_9708,N_7187,N_7203);
nor U9709 (N_9709,N_5246,N_5863);
xor U9710 (N_9710,N_5254,N_6745);
xor U9711 (N_9711,N_5382,N_5899);
nand U9712 (N_9712,N_6878,N_5924);
or U9713 (N_9713,N_6709,N_6662);
or U9714 (N_9714,N_6216,N_6455);
xnor U9715 (N_9715,N_6638,N_6561);
nand U9716 (N_9716,N_5767,N_6467);
or U9717 (N_9717,N_5408,N_5450);
and U9718 (N_9718,N_7314,N_6484);
nand U9719 (N_9719,N_7404,N_5697);
or U9720 (N_9720,N_7240,N_5207);
nand U9721 (N_9721,N_6808,N_5184);
xnor U9722 (N_9722,N_6915,N_7178);
nor U9723 (N_9723,N_6861,N_5119);
nor U9724 (N_9724,N_5223,N_5619);
and U9725 (N_9725,N_7352,N_6932);
xnor U9726 (N_9726,N_5862,N_7208);
nand U9727 (N_9727,N_7333,N_5437);
or U9728 (N_9728,N_5889,N_5988);
or U9729 (N_9729,N_6798,N_5619);
nand U9730 (N_9730,N_5188,N_5490);
nand U9731 (N_9731,N_7076,N_5209);
nor U9732 (N_9732,N_5541,N_6003);
xor U9733 (N_9733,N_6050,N_5038);
nand U9734 (N_9734,N_7278,N_5505);
and U9735 (N_9735,N_7007,N_6974);
or U9736 (N_9736,N_6651,N_7172);
xnor U9737 (N_9737,N_5689,N_5084);
nand U9738 (N_9738,N_5469,N_6208);
and U9739 (N_9739,N_7392,N_6796);
nor U9740 (N_9740,N_5260,N_7461);
xnor U9741 (N_9741,N_6436,N_5908);
or U9742 (N_9742,N_5937,N_7264);
and U9743 (N_9743,N_5280,N_5415);
or U9744 (N_9744,N_7113,N_5187);
nor U9745 (N_9745,N_6317,N_6435);
xnor U9746 (N_9746,N_6217,N_5360);
and U9747 (N_9747,N_5465,N_5273);
and U9748 (N_9748,N_6829,N_5258);
nor U9749 (N_9749,N_5866,N_5857);
nor U9750 (N_9750,N_6048,N_7274);
and U9751 (N_9751,N_7235,N_6692);
xnor U9752 (N_9752,N_6765,N_6721);
xor U9753 (N_9753,N_5259,N_6516);
xor U9754 (N_9754,N_6865,N_5315);
xnor U9755 (N_9755,N_7432,N_6696);
nand U9756 (N_9756,N_7400,N_5116);
nand U9757 (N_9757,N_6816,N_5460);
or U9758 (N_9758,N_6921,N_7381);
or U9759 (N_9759,N_6400,N_6819);
xor U9760 (N_9760,N_6331,N_6698);
or U9761 (N_9761,N_6884,N_5467);
nor U9762 (N_9762,N_6796,N_5447);
xor U9763 (N_9763,N_5117,N_5842);
xor U9764 (N_9764,N_6072,N_6172);
and U9765 (N_9765,N_6470,N_5054);
or U9766 (N_9766,N_5270,N_5501);
nand U9767 (N_9767,N_7141,N_6542);
xnor U9768 (N_9768,N_6260,N_6243);
nor U9769 (N_9769,N_6860,N_6934);
nand U9770 (N_9770,N_7070,N_6496);
xnor U9771 (N_9771,N_7238,N_6579);
or U9772 (N_9772,N_5844,N_6810);
xnor U9773 (N_9773,N_5064,N_5218);
or U9774 (N_9774,N_6448,N_7132);
or U9775 (N_9775,N_5950,N_5776);
nor U9776 (N_9776,N_6166,N_6776);
nor U9777 (N_9777,N_5854,N_5782);
and U9778 (N_9778,N_7207,N_5129);
nand U9779 (N_9779,N_6813,N_6663);
xor U9780 (N_9780,N_7457,N_6204);
or U9781 (N_9781,N_7442,N_7113);
nor U9782 (N_9782,N_6669,N_6436);
or U9783 (N_9783,N_6187,N_7151);
nor U9784 (N_9784,N_6192,N_6611);
nand U9785 (N_9785,N_5927,N_5593);
nand U9786 (N_9786,N_7358,N_7323);
or U9787 (N_9787,N_5889,N_6527);
nor U9788 (N_9788,N_5565,N_6754);
xnor U9789 (N_9789,N_5259,N_7077);
or U9790 (N_9790,N_5207,N_6351);
xor U9791 (N_9791,N_5771,N_5159);
nand U9792 (N_9792,N_5451,N_5901);
or U9793 (N_9793,N_6042,N_7358);
or U9794 (N_9794,N_7168,N_5688);
and U9795 (N_9795,N_6245,N_7327);
nor U9796 (N_9796,N_5180,N_6983);
nor U9797 (N_9797,N_6444,N_6238);
nor U9798 (N_9798,N_5204,N_6486);
and U9799 (N_9799,N_5954,N_5470);
and U9800 (N_9800,N_7349,N_5399);
or U9801 (N_9801,N_6935,N_6708);
xor U9802 (N_9802,N_5821,N_6239);
or U9803 (N_9803,N_5843,N_6468);
or U9804 (N_9804,N_7190,N_6191);
nand U9805 (N_9805,N_6408,N_7287);
xor U9806 (N_9806,N_7492,N_7326);
nand U9807 (N_9807,N_5677,N_7071);
or U9808 (N_9808,N_6651,N_7454);
nand U9809 (N_9809,N_5884,N_6549);
or U9810 (N_9810,N_5050,N_6763);
xnor U9811 (N_9811,N_7078,N_5880);
or U9812 (N_9812,N_5537,N_5212);
and U9813 (N_9813,N_7386,N_5194);
xnor U9814 (N_9814,N_7309,N_5702);
xor U9815 (N_9815,N_6290,N_6738);
or U9816 (N_9816,N_7207,N_7247);
or U9817 (N_9817,N_7256,N_6669);
nor U9818 (N_9818,N_6788,N_5650);
xor U9819 (N_9819,N_6938,N_5684);
nor U9820 (N_9820,N_5566,N_5365);
or U9821 (N_9821,N_5664,N_5161);
and U9822 (N_9822,N_7348,N_7241);
and U9823 (N_9823,N_7250,N_7358);
nor U9824 (N_9824,N_5189,N_5168);
or U9825 (N_9825,N_7005,N_5334);
and U9826 (N_9826,N_5268,N_7180);
nor U9827 (N_9827,N_5764,N_7322);
or U9828 (N_9828,N_6544,N_5781);
and U9829 (N_9829,N_6497,N_6404);
or U9830 (N_9830,N_5414,N_6003);
xor U9831 (N_9831,N_6568,N_6747);
xnor U9832 (N_9832,N_6325,N_7472);
or U9833 (N_9833,N_5147,N_6445);
and U9834 (N_9834,N_6865,N_7016);
and U9835 (N_9835,N_5112,N_6837);
and U9836 (N_9836,N_7024,N_6077);
or U9837 (N_9837,N_6864,N_7171);
nor U9838 (N_9838,N_5417,N_6932);
nor U9839 (N_9839,N_6635,N_5664);
and U9840 (N_9840,N_6935,N_5755);
nor U9841 (N_9841,N_5549,N_6458);
xnor U9842 (N_9842,N_6038,N_5046);
xnor U9843 (N_9843,N_5865,N_6603);
nand U9844 (N_9844,N_5087,N_5041);
or U9845 (N_9845,N_7059,N_6765);
xor U9846 (N_9846,N_5930,N_6933);
or U9847 (N_9847,N_7295,N_5649);
nand U9848 (N_9848,N_5812,N_6016);
and U9849 (N_9849,N_5320,N_6915);
nand U9850 (N_9850,N_6877,N_6722);
and U9851 (N_9851,N_5252,N_6480);
nand U9852 (N_9852,N_6574,N_6245);
and U9853 (N_9853,N_7486,N_5662);
or U9854 (N_9854,N_5548,N_6252);
nand U9855 (N_9855,N_5585,N_5203);
nand U9856 (N_9856,N_6841,N_6809);
and U9857 (N_9857,N_5319,N_6026);
and U9858 (N_9858,N_6018,N_5987);
or U9859 (N_9859,N_5607,N_6417);
or U9860 (N_9860,N_5785,N_7460);
nor U9861 (N_9861,N_5686,N_5111);
xor U9862 (N_9862,N_5211,N_6603);
nor U9863 (N_9863,N_7079,N_5348);
and U9864 (N_9864,N_7374,N_7114);
nor U9865 (N_9865,N_5714,N_6049);
xnor U9866 (N_9866,N_5466,N_6947);
and U9867 (N_9867,N_5108,N_5822);
and U9868 (N_9868,N_5966,N_5347);
nand U9869 (N_9869,N_5642,N_6037);
xnor U9870 (N_9870,N_6906,N_5911);
and U9871 (N_9871,N_7066,N_6486);
and U9872 (N_9872,N_7394,N_7285);
nor U9873 (N_9873,N_7196,N_6939);
or U9874 (N_9874,N_6938,N_6698);
xor U9875 (N_9875,N_6263,N_6926);
or U9876 (N_9876,N_6500,N_6139);
xor U9877 (N_9877,N_7162,N_6572);
and U9878 (N_9878,N_6261,N_6919);
nor U9879 (N_9879,N_5761,N_6345);
xnor U9880 (N_9880,N_6859,N_5589);
nand U9881 (N_9881,N_6657,N_5548);
nor U9882 (N_9882,N_7447,N_6427);
nor U9883 (N_9883,N_6750,N_5843);
and U9884 (N_9884,N_5618,N_7229);
nor U9885 (N_9885,N_5314,N_6230);
and U9886 (N_9886,N_6329,N_6876);
nand U9887 (N_9887,N_6998,N_6484);
and U9888 (N_9888,N_6243,N_6974);
nand U9889 (N_9889,N_6525,N_7251);
and U9890 (N_9890,N_5011,N_5149);
or U9891 (N_9891,N_6201,N_5292);
or U9892 (N_9892,N_5515,N_6281);
or U9893 (N_9893,N_5944,N_6928);
and U9894 (N_9894,N_7378,N_6862);
and U9895 (N_9895,N_5804,N_7232);
and U9896 (N_9896,N_5977,N_5267);
nand U9897 (N_9897,N_5084,N_5436);
nor U9898 (N_9898,N_6888,N_6837);
nor U9899 (N_9899,N_6515,N_7052);
xnor U9900 (N_9900,N_6477,N_5310);
and U9901 (N_9901,N_5669,N_6863);
nor U9902 (N_9902,N_5341,N_6582);
and U9903 (N_9903,N_5183,N_6700);
or U9904 (N_9904,N_5162,N_6169);
or U9905 (N_9905,N_6230,N_5020);
or U9906 (N_9906,N_6015,N_6029);
or U9907 (N_9907,N_6502,N_6930);
xor U9908 (N_9908,N_5681,N_6838);
or U9909 (N_9909,N_6783,N_6654);
and U9910 (N_9910,N_6565,N_6856);
nand U9911 (N_9911,N_6560,N_5236);
nand U9912 (N_9912,N_7212,N_5366);
xnor U9913 (N_9913,N_5565,N_6719);
and U9914 (N_9914,N_6788,N_5370);
and U9915 (N_9915,N_6978,N_5103);
or U9916 (N_9916,N_7402,N_5308);
nor U9917 (N_9917,N_6648,N_5283);
nand U9918 (N_9918,N_5887,N_7324);
and U9919 (N_9919,N_5433,N_5403);
and U9920 (N_9920,N_5416,N_7016);
and U9921 (N_9921,N_5068,N_6346);
nor U9922 (N_9922,N_7292,N_5138);
nand U9923 (N_9923,N_6152,N_5091);
nand U9924 (N_9924,N_7416,N_6739);
nand U9925 (N_9925,N_7457,N_5863);
or U9926 (N_9926,N_7370,N_6344);
or U9927 (N_9927,N_5115,N_5426);
or U9928 (N_9928,N_5757,N_5200);
and U9929 (N_9929,N_5054,N_6173);
nand U9930 (N_9930,N_6953,N_5117);
or U9931 (N_9931,N_7227,N_5337);
or U9932 (N_9932,N_7072,N_5985);
nand U9933 (N_9933,N_5292,N_6646);
nand U9934 (N_9934,N_6334,N_6232);
nand U9935 (N_9935,N_6790,N_6112);
nor U9936 (N_9936,N_7293,N_5104);
xor U9937 (N_9937,N_5441,N_5746);
or U9938 (N_9938,N_7126,N_6438);
nor U9939 (N_9939,N_5853,N_5512);
xnor U9940 (N_9940,N_6526,N_7042);
or U9941 (N_9941,N_5484,N_6606);
or U9942 (N_9942,N_6067,N_6246);
nor U9943 (N_9943,N_7069,N_7481);
nor U9944 (N_9944,N_5177,N_7065);
or U9945 (N_9945,N_6270,N_5189);
or U9946 (N_9946,N_5525,N_5066);
xor U9947 (N_9947,N_7471,N_5863);
nand U9948 (N_9948,N_6498,N_5654);
and U9949 (N_9949,N_5091,N_5266);
xor U9950 (N_9950,N_6480,N_6812);
or U9951 (N_9951,N_5336,N_6945);
or U9952 (N_9952,N_7157,N_6792);
nor U9953 (N_9953,N_6273,N_5584);
xor U9954 (N_9954,N_7445,N_7253);
nor U9955 (N_9955,N_6229,N_7231);
or U9956 (N_9956,N_6416,N_6301);
nand U9957 (N_9957,N_5328,N_6743);
or U9958 (N_9958,N_6975,N_7028);
nand U9959 (N_9959,N_7012,N_6005);
nor U9960 (N_9960,N_6695,N_6503);
nor U9961 (N_9961,N_5440,N_5587);
nand U9962 (N_9962,N_6571,N_5119);
xor U9963 (N_9963,N_5363,N_6753);
nor U9964 (N_9964,N_7165,N_6812);
or U9965 (N_9965,N_5727,N_6473);
nor U9966 (N_9966,N_5809,N_7035);
nand U9967 (N_9967,N_5855,N_6627);
xor U9968 (N_9968,N_6065,N_7433);
nand U9969 (N_9969,N_7110,N_5978);
or U9970 (N_9970,N_7244,N_5283);
nand U9971 (N_9971,N_5787,N_5067);
nor U9972 (N_9972,N_6418,N_6123);
and U9973 (N_9973,N_7282,N_7061);
and U9974 (N_9974,N_5114,N_5790);
nor U9975 (N_9975,N_5104,N_5143);
nand U9976 (N_9976,N_6753,N_6972);
xor U9977 (N_9977,N_5431,N_7140);
xor U9978 (N_9978,N_6248,N_7211);
nor U9979 (N_9979,N_5960,N_6610);
or U9980 (N_9980,N_5534,N_7390);
nor U9981 (N_9981,N_5894,N_7060);
nor U9982 (N_9982,N_6747,N_5228);
and U9983 (N_9983,N_6780,N_6605);
and U9984 (N_9984,N_6756,N_5142);
nor U9985 (N_9985,N_7294,N_5541);
or U9986 (N_9986,N_7476,N_5709);
nor U9987 (N_9987,N_7177,N_7056);
and U9988 (N_9988,N_7290,N_6761);
or U9989 (N_9989,N_5321,N_6470);
nor U9990 (N_9990,N_5667,N_5468);
nor U9991 (N_9991,N_6531,N_5185);
xnor U9992 (N_9992,N_5932,N_5714);
nand U9993 (N_9993,N_7102,N_5405);
nor U9994 (N_9994,N_6310,N_6458);
nand U9995 (N_9995,N_7470,N_6668);
and U9996 (N_9996,N_5732,N_5951);
nand U9997 (N_9997,N_5318,N_5288);
and U9998 (N_9998,N_5561,N_6983);
nor U9999 (N_9999,N_5932,N_5810);
xor UO_0 (O_0,N_9315,N_9109);
or UO_1 (O_1,N_8144,N_9081);
and UO_2 (O_2,N_8729,N_7620);
nor UO_3 (O_3,N_8514,N_9686);
xor UO_4 (O_4,N_9875,N_8964);
nor UO_5 (O_5,N_7529,N_9764);
nand UO_6 (O_6,N_9526,N_9171);
nor UO_7 (O_7,N_7834,N_9520);
and UO_8 (O_8,N_9303,N_8907);
xnor UO_9 (O_9,N_7976,N_9126);
nand UO_10 (O_10,N_9298,N_7953);
nand UO_11 (O_11,N_8105,N_8091);
or UO_12 (O_12,N_8647,N_9196);
nand UO_13 (O_13,N_9436,N_8842);
and UO_14 (O_14,N_7954,N_9593);
nor UO_15 (O_15,N_9967,N_8324);
nor UO_16 (O_16,N_8624,N_8449);
or UO_17 (O_17,N_8423,N_9037);
xor UO_18 (O_18,N_8009,N_9955);
xnor UO_19 (O_19,N_7669,N_9750);
and UO_20 (O_20,N_8222,N_8694);
nor UO_21 (O_21,N_7527,N_7764);
nor UO_22 (O_22,N_8262,N_8915);
xor UO_23 (O_23,N_7896,N_9505);
and UO_24 (O_24,N_7651,N_8470);
nor UO_25 (O_25,N_7504,N_8456);
nand UO_26 (O_26,N_8741,N_9355);
xnor UO_27 (O_27,N_8497,N_9842);
nand UO_28 (O_28,N_7857,N_7972);
nand UO_29 (O_29,N_8448,N_9963);
or UO_30 (O_30,N_8788,N_9388);
or UO_31 (O_31,N_9926,N_9840);
nand UO_32 (O_32,N_8180,N_7913);
and UO_33 (O_33,N_8780,N_8162);
or UO_34 (O_34,N_7705,N_8601);
and UO_35 (O_35,N_7926,N_9628);
nor UO_36 (O_36,N_8755,N_7945);
or UO_37 (O_37,N_8905,N_8159);
nand UO_38 (O_38,N_7961,N_8765);
and UO_39 (O_39,N_9155,N_7829);
nor UO_40 (O_40,N_7995,N_8848);
or UO_41 (O_41,N_8465,N_9683);
nor UO_42 (O_42,N_8068,N_9542);
nand UO_43 (O_43,N_8975,N_9787);
nor UO_44 (O_44,N_7747,N_9825);
and UO_45 (O_45,N_8256,N_9134);
and UO_46 (O_46,N_8434,N_9713);
xor UO_47 (O_47,N_9739,N_7664);
nor UO_48 (O_48,N_9027,N_7964);
and UO_49 (O_49,N_8223,N_9437);
xnor UO_50 (O_50,N_9264,N_8045);
or UO_51 (O_51,N_7724,N_8752);
nor UO_52 (O_52,N_9491,N_8948);
and UO_53 (O_53,N_9814,N_8220);
nor UO_54 (O_54,N_7791,N_7606);
nand UO_55 (O_55,N_8409,N_9152);
nand UO_56 (O_56,N_8711,N_8730);
and UO_57 (O_57,N_8827,N_8316);
xnor UO_58 (O_58,N_7854,N_8749);
nand UO_59 (O_59,N_9177,N_8475);
or UO_60 (O_60,N_9116,N_9668);
or UO_61 (O_61,N_9891,N_8268);
nor UO_62 (O_62,N_8861,N_9295);
xor UO_63 (O_63,N_7503,N_9577);
xor UO_64 (O_64,N_7978,N_9404);
nor UO_65 (O_65,N_8230,N_8295);
xor UO_66 (O_66,N_9680,N_8330);
xnor UO_67 (O_67,N_7958,N_8961);
nand UO_68 (O_68,N_9993,N_9103);
nor UO_69 (O_69,N_9884,N_9775);
nor UO_70 (O_70,N_9416,N_8480);
and UO_71 (O_71,N_9465,N_9267);
and UO_72 (O_72,N_8306,N_8996);
nand UO_73 (O_73,N_8175,N_8691);
xor UO_74 (O_74,N_9689,N_8642);
or UO_75 (O_75,N_8745,N_7649);
xor UO_76 (O_76,N_8547,N_8705);
nor UO_77 (O_77,N_8696,N_9205);
xor UO_78 (O_78,N_7956,N_9531);
nand UO_79 (O_79,N_7540,N_9794);
nand UO_80 (O_80,N_9877,N_7973);
nand UO_81 (O_81,N_9914,N_8061);
and UO_82 (O_82,N_9943,N_9497);
nor UO_83 (O_83,N_7563,N_8002);
and UO_84 (O_84,N_9788,N_9307);
and UO_85 (O_85,N_7640,N_8777);
nor UO_86 (O_86,N_8797,N_8196);
xor UO_87 (O_87,N_8543,N_9864);
nand UO_88 (O_88,N_8687,N_8633);
nand UO_89 (O_89,N_7979,N_8927);
and UO_90 (O_90,N_9507,N_9031);
nand UO_91 (O_91,N_7681,N_9682);
nor UO_92 (O_92,N_8972,N_8431);
or UO_93 (O_93,N_8999,N_8962);
and UO_94 (O_94,N_9795,N_9285);
nor UO_95 (O_95,N_8513,N_9965);
xor UO_96 (O_96,N_9957,N_8454);
or UO_97 (O_97,N_7610,N_9612);
xor UO_98 (O_98,N_9151,N_7536);
nor UO_99 (O_99,N_9895,N_7952);
nand UO_100 (O_100,N_8899,N_9816);
xnor UO_101 (O_101,N_7888,N_8488);
or UO_102 (O_102,N_9170,N_8496);
nor UO_103 (O_103,N_7862,N_7505);
nand UO_104 (O_104,N_9589,N_7611);
and UO_105 (O_105,N_8122,N_7615);
xor UO_106 (O_106,N_7641,N_9799);
and UO_107 (O_107,N_8243,N_7673);
and UO_108 (O_108,N_9930,N_8479);
or UO_109 (O_109,N_7562,N_8791);
and UO_110 (O_110,N_8461,N_9278);
or UO_111 (O_111,N_7583,N_8548);
xnor UO_112 (O_112,N_7515,N_8918);
and UO_113 (O_113,N_8618,N_7553);
and UO_114 (O_114,N_9880,N_8892);
nor UO_115 (O_115,N_8864,N_8049);
xor UO_116 (O_116,N_9405,N_8081);
nor UO_117 (O_117,N_9075,N_7831);
nand UO_118 (O_118,N_7692,N_9079);
xor UO_119 (O_119,N_8874,N_8327);
or UO_120 (O_120,N_9472,N_8212);
nor UO_121 (O_121,N_9654,N_7839);
nand UO_122 (O_122,N_7604,N_7548);
nor UO_123 (O_123,N_8527,N_9870);
or UO_124 (O_124,N_7512,N_9883);
or UO_125 (O_125,N_8870,N_9874);
and UO_126 (O_126,N_7866,N_7818);
nor UO_127 (O_127,N_9857,N_9136);
xnor UO_128 (O_128,N_8151,N_9362);
or UO_129 (O_129,N_9546,N_9956);
or UO_130 (O_130,N_9178,N_9025);
nand UO_131 (O_131,N_9016,N_9083);
nand UO_132 (O_132,N_9624,N_9928);
nor UO_133 (O_133,N_8845,N_9694);
and UO_134 (O_134,N_9143,N_9435);
xor UO_135 (O_135,N_9474,N_9559);
or UO_136 (O_136,N_9499,N_9919);
xor UO_137 (O_137,N_9467,N_7689);
nand UO_138 (O_138,N_8373,N_9020);
nor UO_139 (O_139,N_9731,N_9233);
and UO_140 (O_140,N_9476,N_9541);
or UO_141 (O_141,N_9516,N_8377);
and UO_142 (O_142,N_7549,N_8690);
and UO_143 (O_143,N_9906,N_7694);
and UO_144 (O_144,N_8176,N_8013);
and UO_145 (O_145,N_8652,N_8519);
nor UO_146 (O_146,N_8440,N_8047);
xnor UO_147 (O_147,N_8406,N_8900);
or UO_148 (O_148,N_7977,N_9420);
xnor UO_149 (O_149,N_9270,N_9304);
and UO_150 (O_150,N_9243,N_9064);
or UO_151 (O_151,N_9294,N_9661);
nand UO_152 (O_152,N_9157,N_9970);
nor UO_153 (O_153,N_9718,N_8312);
nor UO_154 (O_154,N_9801,N_9346);
nor UO_155 (O_155,N_8979,N_7612);
nor UO_156 (O_156,N_8700,N_8878);
and UO_157 (O_157,N_8552,N_8883);
xnor UO_158 (O_158,N_9466,N_8202);
xor UO_159 (O_159,N_9872,N_7573);
xnor UO_160 (O_160,N_8005,N_8632);
xnor UO_161 (O_161,N_9826,N_8984);
nand UO_162 (O_162,N_8364,N_7766);
nor UO_163 (O_163,N_9123,N_9754);
nand UO_164 (O_164,N_8404,N_9184);
nand UO_165 (O_165,N_7723,N_8492);
nor UO_166 (O_166,N_9836,N_8796);
and UO_167 (O_167,N_8795,N_9937);
and UO_168 (O_168,N_9591,N_9832);
or UO_169 (O_169,N_8494,N_9700);
nand UO_170 (O_170,N_9940,N_9827);
nor UO_171 (O_171,N_8171,N_9746);
nand UO_172 (O_172,N_8334,N_9063);
nor UO_173 (O_173,N_8909,N_9908);
nor UO_174 (O_174,N_7805,N_7628);
nand UO_175 (O_175,N_8048,N_8375);
and UO_176 (O_176,N_9334,N_9815);
and UO_177 (O_177,N_7859,N_8981);
nand UO_178 (O_178,N_8693,N_9250);
nand UO_179 (O_179,N_8289,N_7630);
or UO_180 (O_180,N_8123,N_8060);
xnor UO_181 (O_181,N_7517,N_9637);
xor UO_182 (O_182,N_7927,N_9649);
xnor UO_183 (O_183,N_7579,N_7833);
and UO_184 (O_184,N_7544,N_7986);
or UO_185 (O_185,N_9108,N_8390);
xnor UO_186 (O_186,N_8075,N_9481);
or UO_187 (O_187,N_9949,N_9479);
nor UO_188 (O_188,N_7974,N_7777);
nor UO_189 (O_189,N_7572,N_8750);
or UO_190 (O_190,N_7537,N_9089);
nor UO_191 (O_191,N_9732,N_9777);
or UO_192 (O_192,N_7781,N_9318);
and UO_193 (O_193,N_9458,N_7545);
nor UO_194 (O_194,N_7883,N_9810);
nand UO_195 (O_195,N_9087,N_8712);
nand UO_196 (O_196,N_9807,N_9978);
nand UO_197 (O_197,N_8567,N_7653);
nand UO_198 (O_198,N_8623,N_8681);
and UO_199 (O_199,N_7775,N_9973);
or UO_200 (O_200,N_9859,N_9129);
nand UO_201 (O_201,N_8916,N_8634);
nand UO_202 (O_202,N_8432,N_7812);
xor UO_203 (O_203,N_8043,N_7750);
or UO_204 (O_204,N_9246,N_7917);
nand UO_205 (O_205,N_8142,N_7982);
xnor UO_206 (O_206,N_9347,N_8938);
or UO_207 (O_207,N_9770,N_9008);
and UO_208 (O_208,N_9256,N_9399);
xnor UO_209 (O_209,N_8239,N_7817);
nor UO_210 (O_210,N_9641,N_7752);
nor UO_211 (O_211,N_9805,N_8779);
nand UO_212 (O_212,N_9569,N_7696);
xnor UO_213 (O_213,N_8393,N_8355);
and UO_214 (O_214,N_9340,N_8310);
and UO_215 (O_215,N_9525,N_8811);
or UO_216 (O_216,N_7707,N_9962);
nor UO_217 (O_217,N_8871,N_9773);
nor UO_218 (O_218,N_8433,N_9968);
and UO_219 (O_219,N_9708,N_8912);
nand UO_220 (O_220,N_7746,N_9371);
xor UO_221 (O_221,N_8638,N_9696);
nor UO_222 (O_222,N_7571,N_8235);
or UO_223 (O_223,N_8088,N_8774);
nor UO_224 (O_224,N_9677,N_8704);
nor UO_225 (O_225,N_9760,N_8130);
nor UO_226 (O_226,N_8588,N_8258);
or UO_227 (O_227,N_7999,N_7867);
nand UO_228 (O_228,N_9780,N_9976);
and UO_229 (O_229,N_9176,N_9321);
nand UO_230 (O_230,N_8149,N_8302);
nand UO_231 (O_231,N_8341,N_9287);
nand UO_232 (O_232,N_8879,N_7959);
nor UO_233 (O_233,N_9735,N_8391);
nand UO_234 (O_234,N_9092,N_9581);
and UO_235 (O_235,N_9900,N_8085);
nor UO_236 (O_236,N_7555,N_8935);
or UO_237 (O_237,N_9600,N_8993);
xnor UO_238 (O_238,N_9161,N_8007);
and UO_239 (O_239,N_9301,N_8438);
nand UO_240 (O_240,N_9488,N_9232);
xor UO_241 (O_241,N_9084,N_8904);
nand UO_242 (O_242,N_9980,N_9172);
and UO_243 (O_243,N_9158,N_7909);
nor UO_244 (O_244,N_8453,N_8771);
or UO_245 (O_245,N_9284,N_8034);
xor UO_246 (O_246,N_8739,N_8619);
xor UO_247 (O_247,N_8221,N_7645);
xor UO_248 (O_248,N_9942,N_8669);
nand UO_249 (O_249,N_9858,N_8246);
xor UO_250 (O_250,N_9240,N_9360);
xor UO_251 (O_251,N_7756,N_8402);
nand UO_252 (O_252,N_7558,N_9005);
or UO_253 (O_253,N_9596,N_7785);
or UO_254 (O_254,N_9571,N_8857);
xor UO_255 (O_255,N_9691,N_7969);
nand UO_256 (O_256,N_9761,N_8555);
nand UO_257 (O_257,N_9998,N_9389);
or UO_258 (O_258,N_7672,N_7758);
and UO_259 (O_259,N_7970,N_8836);
or UO_260 (O_260,N_8509,N_9055);
or UO_261 (O_261,N_8491,N_9644);
and UO_262 (O_262,N_9021,N_8420);
xnor UO_263 (O_263,N_7815,N_7789);
nand UO_264 (O_264,N_8169,N_8291);
xor UO_265 (O_265,N_8792,N_9131);
or UO_266 (O_266,N_8510,N_7835);
or UO_267 (O_267,N_8775,N_8150);
nand UO_268 (O_268,N_9165,N_8512);
and UO_269 (O_269,N_9663,N_8401);
or UO_270 (O_270,N_7726,N_9580);
nand UO_271 (O_271,N_8668,N_8133);
xnor UO_272 (O_272,N_8279,N_8216);
nor UO_273 (O_273,N_8666,N_7698);
or UO_274 (O_274,N_7703,N_8462);
and UO_275 (O_275,N_9395,N_7626);
or UO_276 (O_276,N_8766,N_8111);
or UO_277 (O_277,N_8228,N_8217);
and UO_278 (O_278,N_8374,N_7784);
nor UO_279 (O_279,N_7535,N_8102);
or UO_280 (O_280,N_9623,N_8953);
xnor UO_281 (O_281,N_8004,N_8400);
nor UO_282 (O_282,N_8641,N_9527);
xor UO_283 (O_283,N_8969,N_8337);
nor UO_284 (O_284,N_9975,N_9168);
or UO_285 (O_285,N_9633,N_9440);
xnor UO_286 (O_286,N_9626,N_9583);
and UO_287 (O_287,N_9227,N_9769);
nor UO_288 (O_288,N_7621,N_9582);
nand UO_289 (O_289,N_9394,N_7680);
nor UO_290 (O_290,N_8658,N_7871);
nand UO_291 (O_291,N_8020,N_9709);
nor UO_292 (O_292,N_8264,N_9019);
nor UO_293 (O_293,N_9100,N_8551);
and UO_294 (O_294,N_8825,N_7714);
or UO_295 (O_295,N_8833,N_9515);
nor UO_296 (O_296,N_8192,N_8053);
nor UO_297 (O_297,N_8155,N_9164);
nor UO_298 (O_298,N_8136,N_9557);
or UO_299 (O_299,N_9763,N_9049);
nand UO_300 (O_300,N_9255,N_9945);
nor UO_301 (O_301,N_7518,N_8080);
or UO_302 (O_302,N_8959,N_8054);
or UO_303 (O_303,N_9309,N_7910);
or UO_304 (O_304,N_9793,N_7912);
nor UO_305 (O_305,N_8482,N_8683);
and UO_306 (O_306,N_9621,N_9707);
or UO_307 (O_307,N_8742,N_8466);
nand UO_308 (O_308,N_9122,N_8835);
and UO_309 (O_309,N_7605,N_9785);
or UO_310 (O_310,N_7638,N_8106);
nor UO_311 (O_311,N_8824,N_8326);
and UO_312 (O_312,N_9114,N_8358);
xor UO_313 (O_313,N_7780,N_7711);
and UO_314 (O_314,N_9283,N_8985);
nor UO_315 (O_315,N_8347,N_9345);
nor UO_316 (O_316,N_7666,N_8017);
and UO_317 (O_317,N_9265,N_8224);
or UO_318 (O_318,N_7807,N_8773);
and UO_319 (O_319,N_9473,N_9230);
nor UO_320 (O_320,N_8182,N_9209);
nand UO_321 (O_321,N_8037,N_8506);
nor UO_322 (O_322,N_9915,N_7836);
or UO_323 (O_323,N_8349,N_9979);
nor UO_324 (O_324,N_8903,N_8472);
nor UO_325 (O_325,N_9838,N_7801);
and UO_326 (O_326,N_9705,N_9206);
or UO_327 (O_327,N_9030,N_7845);
nand UO_328 (O_328,N_8022,N_9819);
and UO_329 (O_329,N_9625,N_8052);
or UO_330 (O_330,N_9572,N_8782);
xor UO_331 (O_331,N_7670,N_8701);
xnor UO_332 (O_332,N_8338,N_9349);
nor UO_333 (O_333,N_7613,N_8876);
nand UO_334 (O_334,N_8101,N_7588);
nand UO_335 (O_335,N_9464,N_7892);
xnor UO_336 (O_336,N_7884,N_9077);
nand UO_337 (O_337,N_9720,N_9556);
nor UO_338 (O_338,N_8132,N_8158);
nor UO_339 (O_339,N_9638,N_9385);
nor UO_340 (O_340,N_9927,N_9809);
nand UO_341 (O_341,N_7510,N_8096);
or UO_342 (O_342,N_7656,N_9128);
xnor UO_343 (O_343,N_8332,N_8625);
nand UO_344 (O_344,N_8914,N_7542);
or UO_345 (O_345,N_7797,N_9828);
and UO_346 (O_346,N_9017,N_8826);
or UO_347 (O_347,N_9426,N_9043);
nor UO_348 (O_348,N_8441,N_8850);
and UO_349 (O_349,N_8671,N_7924);
and UO_350 (O_350,N_9193,N_8604);
nand UO_351 (O_351,N_9470,N_8630);
nand UO_352 (O_352,N_7879,N_8757);
xor UO_353 (O_353,N_8181,N_8923);
xor UO_354 (O_354,N_8397,N_7864);
and UO_355 (O_355,N_7509,N_9563);
nor UO_356 (O_356,N_8376,N_7753);
nand UO_357 (O_357,N_8887,N_8902);
nand UO_358 (O_358,N_9174,N_9549);
xor UO_359 (O_359,N_8645,N_9590);
nand UO_360 (O_360,N_9118,N_7849);
nor UO_361 (O_361,N_8134,N_8098);
xnor UO_362 (O_362,N_8413,N_9459);
or UO_363 (O_363,N_9221,N_8934);
xor UO_364 (O_364,N_9702,N_9598);
nor UO_365 (O_365,N_9144,N_9802);
and UO_366 (O_366,N_8010,N_8906);
and UO_367 (O_367,N_8145,N_9575);
nor UO_368 (O_368,N_9540,N_9640);
nor UO_369 (O_369,N_9886,N_9292);
xnor UO_370 (O_370,N_7962,N_9276);
or UO_371 (O_371,N_8897,N_8362);
nor UO_372 (O_372,N_8713,N_9873);
xor UO_373 (O_373,N_9511,N_9441);
nor UO_374 (O_374,N_8858,N_8895);
nor UO_375 (O_375,N_9220,N_9489);
xor UO_376 (O_376,N_9052,N_9153);
and UO_377 (O_377,N_7901,N_8637);
xnor UO_378 (O_378,N_9410,N_8852);
nor UO_379 (O_379,N_7916,N_8317);
and UO_380 (O_380,N_7826,N_7985);
and UO_381 (O_381,N_7902,N_8946);
and UO_382 (O_382,N_8304,N_9237);
and UO_383 (O_383,N_9939,N_9185);
nor UO_384 (O_384,N_9982,N_9796);
nor UO_385 (O_385,N_8398,N_9163);
and UO_386 (O_386,N_9905,N_7650);
xor UO_387 (O_387,N_9190,N_7687);
and UO_388 (O_388,N_8129,N_8354);
nor UO_389 (O_389,N_9024,N_9258);
nand UO_390 (O_390,N_9681,N_7660);
or UO_391 (O_391,N_7551,N_8550);
and UO_392 (O_392,N_8227,N_8951);
nand UO_393 (O_393,N_8225,N_8185);
and UO_394 (O_394,N_9584,N_8352);
nand UO_395 (O_395,N_8076,N_8571);
xnor UO_396 (O_396,N_8501,N_9071);
xor UO_397 (O_397,N_7994,N_8763);
nor UO_398 (O_398,N_8089,N_7809);
nand UO_399 (O_399,N_9698,N_9747);
and UO_400 (O_400,N_9194,N_8890);
or UO_401 (O_401,N_7806,N_9999);
nor UO_402 (O_402,N_9881,N_9667);
nor UO_403 (O_403,N_9837,N_7811);
nand UO_404 (O_404,N_7998,N_7798);
or UO_405 (O_405,N_7800,N_8649);
xnor UO_406 (O_406,N_8884,N_9182);
and UO_407 (O_407,N_8605,N_9647);
and UO_408 (O_408,N_7602,N_9703);
and UO_409 (O_409,N_9188,N_9811);
nor UO_410 (O_410,N_9379,N_8793);
or UO_411 (O_411,N_7772,N_9715);
nand UO_412 (O_412,N_9719,N_9393);
nor UO_413 (O_413,N_9833,N_9888);
nor UO_414 (O_414,N_9959,N_8573);
or UO_415 (O_415,N_9411,N_9291);
nor UO_416 (O_416,N_9972,N_8410);
xnor UO_417 (O_417,N_9197,N_7730);
or UO_418 (O_418,N_8919,N_8515);
nor UO_419 (O_419,N_8273,N_8989);
or UO_420 (O_420,N_8939,N_8813);
and UO_421 (O_421,N_9851,N_9482);
xor UO_422 (O_422,N_8115,N_8810);
and UO_423 (O_423,N_7821,N_9282);
nor UO_424 (O_424,N_9313,N_8800);
or UO_425 (O_425,N_9086,N_9533);
nor UO_426 (O_426,N_9931,N_9145);
and UO_427 (O_427,N_7850,N_9768);
nand UO_428 (O_428,N_9512,N_8925);
or UO_429 (O_429,N_9106,N_9358);
nand UO_430 (O_430,N_8271,N_9224);
xnor UO_431 (O_431,N_9018,N_8566);
nor UO_432 (O_432,N_9532,N_7686);
or UO_433 (O_433,N_8275,N_8847);
nor UO_434 (O_434,N_8533,N_7713);
and UO_435 (O_435,N_9803,N_8976);
nor UO_436 (O_436,N_9069,N_8342);
nand UO_437 (O_437,N_9726,N_9800);
nand UO_438 (O_438,N_9124,N_7556);
or UO_439 (O_439,N_8293,N_8365);
nand UO_440 (O_440,N_8849,N_8917);
and UO_441 (O_441,N_8767,N_7508);
xnor UO_442 (O_442,N_9317,N_9852);
nor UO_443 (O_443,N_9279,N_8025);
nor UO_444 (O_444,N_7869,N_8417);
or UO_445 (O_445,N_9297,N_8209);
xnor UO_446 (O_446,N_7591,N_8100);
or UO_447 (O_447,N_8173,N_8877);
and UO_448 (O_448,N_8655,N_8331);
nor UO_449 (O_449,N_7662,N_9879);
or UO_450 (O_450,N_9257,N_9697);
nor UO_451 (O_451,N_9091,N_9894);
and UO_452 (O_452,N_8261,N_8529);
xnor UO_453 (O_453,N_8255,N_7841);
xor UO_454 (O_454,N_9062,N_9609);
and UO_455 (O_455,N_7943,N_8487);
nand UO_456 (O_456,N_9766,N_7759);
nand UO_457 (O_457,N_8523,N_8574);
nor UO_458 (O_458,N_8179,N_8803);
and UO_459 (O_459,N_7599,N_9632);
nor UO_460 (O_460,N_9409,N_8965);
and UO_461 (O_461,N_8908,N_9645);
nand UO_462 (O_462,N_8992,N_9863);
and UO_463 (O_463,N_8591,N_8485);
xnor UO_464 (O_464,N_9314,N_7941);
or UO_465 (O_465,N_8815,N_8654);
nand UO_466 (O_466,N_8517,N_9740);
xor UO_467 (O_467,N_9444,N_9566);
nand UO_468 (O_468,N_9365,N_9186);
xnor UO_469 (O_469,N_9755,N_8280);
or UO_470 (O_470,N_9722,N_8971);
nand UO_471 (O_471,N_9305,N_9994);
and UO_472 (O_472,N_9651,N_9669);
nor UO_473 (O_473,N_8041,N_8039);
and UO_474 (O_474,N_7574,N_8772);
or UO_475 (O_475,N_8926,N_7617);
nor UO_476 (O_476,N_8277,N_8190);
nand UO_477 (O_477,N_9348,N_7722);
nand UO_478 (O_478,N_8036,N_7898);
xnor UO_479 (O_479,N_9280,N_8477);
nand UO_480 (O_480,N_9611,N_9223);
and UO_481 (O_481,N_7987,N_7949);
nor UO_482 (O_482,N_8594,N_7708);
nand UO_483 (O_483,N_8561,N_8403);
or UO_484 (O_484,N_9138,N_9203);
nor UO_485 (O_485,N_8640,N_8819);
nand UO_486 (O_486,N_9610,N_9372);
nand UO_487 (O_487,N_9460,N_8720);
xnor UO_488 (O_488,N_8534,N_9784);
and UO_489 (O_489,N_7802,N_9180);
and UO_490 (O_490,N_9862,N_8886);
xnor UO_491 (O_491,N_9202,N_8955);
nor UO_492 (O_492,N_7937,N_8814);
or UO_493 (O_493,N_9322,N_8042);
nand UO_494 (O_494,N_9869,N_8611);
xor UO_495 (O_495,N_9783,N_9293);
or UO_496 (O_496,N_9534,N_7914);
or UO_497 (O_497,N_9074,N_7861);
or UO_498 (O_498,N_9995,N_7830);
xnor UO_499 (O_499,N_9727,N_9944);
or UO_500 (O_500,N_7648,N_8458);
nand UO_501 (O_501,N_8165,N_9808);
or UO_502 (O_502,N_9160,N_8430);
and UO_503 (O_503,N_9462,N_7838);
and UO_504 (O_504,N_9781,N_9748);
nor UO_505 (O_505,N_8535,N_8808);
nor UO_506 (O_506,N_7567,N_8667);
and UO_507 (O_507,N_9226,N_9023);
nor UO_508 (O_508,N_8659,N_9117);
xor UO_509 (O_509,N_7771,N_8270);
nor UO_510 (O_510,N_9288,N_9015);
nor UO_511 (O_511,N_8234,N_8753);
and UO_512 (O_512,N_8298,N_9311);
and UO_513 (O_513,N_8673,N_8307);
and UO_514 (O_514,N_9095,N_9933);
nor UO_515 (O_515,N_8284,N_9300);
xnor UO_516 (O_516,N_9150,N_9387);
and UO_517 (O_517,N_8853,N_9323);
xor UO_518 (O_518,N_9710,N_9588);
or UO_519 (O_519,N_7552,N_9920);
nor UO_520 (O_520,N_9350,N_9113);
or UO_521 (O_521,N_9854,N_8988);
and UO_522 (O_522,N_8073,N_8356);
xor UO_523 (O_523,N_7674,N_9627);
and UO_524 (O_524,N_8760,N_8357);
xor UO_525 (O_525,N_7846,N_9119);
nand UO_526 (O_526,N_7633,N_7968);
nor UO_527 (O_527,N_8718,N_8072);
nor UO_528 (O_528,N_8931,N_8074);
nor UO_529 (O_529,N_7940,N_8094);
nand UO_530 (O_530,N_8560,N_7848);
or UO_531 (O_531,N_8493,N_9048);
xor UO_532 (O_532,N_9234,N_8503);
and UO_533 (O_533,N_8941,N_8481);
or UO_534 (O_534,N_8412,N_9342);
and UO_535 (O_535,N_7890,N_8582);
xnor UO_536 (O_536,N_7655,N_7623);
nor UO_537 (O_537,N_7684,N_8930);
nand UO_538 (O_538,N_9038,N_8875);
nand UO_539 (O_539,N_9363,N_9361);
xor UO_540 (O_540,N_7930,N_8205);
xor UO_541 (O_541,N_7715,N_8266);
xnor UO_542 (O_542,N_7526,N_8056);
xnor UO_543 (O_543,N_7589,N_9790);
xnor UO_544 (O_544,N_9774,N_8860);
xor UO_545 (O_545,N_9675,N_8429);
nor UO_546 (O_546,N_9548,N_8469);
nor UO_547 (O_547,N_8125,N_9094);
and UO_548 (O_548,N_7614,N_9208);
nand UO_549 (O_549,N_9357,N_8621);
and UO_550 (O_550,N_9181,N_9951);
or UO_551 (O_551,N_8735,N_8473);
xnor UO_552 (O_552,N_9985,N_8674);
or UO_553 (O_553,N_9759,N_8544);
or UO_554 (O_554,N_8361,N_8436);
or UO_555 (O_555,N_9929,N_9014);
or UO_556 (O_556,N_8636,N_9758);
nor UO_557 (O_557,N_8051,N_8881);
and UO_558 (O_558,N_7559,N_9080);
nand UO_559 (O_559,N_7538,N_8723);
xor UO_560 (O_560,N_9723,N_9306);
nand UO_561 (O_561,N_9871,N_9742);
or UO_562 (O_562,N_9222,N_9539);
xor UO_563 (O_563,N_8790,N_8252);
xnor UO_564 (O_564,N_8421,N_8077);
xor UO_565 (O_565,N_8950,N_8751);
and UO_566 (O_566,N_7847,N_7719);
or UO_567 (O_567,N_8383,N_9946);
or UO_568 (O_568,N_9910,N_7925);
xnor UO_569 (O_569,N_8977,N_8038);
nand UO_570 (O_570,N_9034,N_8556);
nor UO_571 (O_571,N_8558,N_9898);
nor UO_572 (O_572,N_8059,N_9111);
and UO_573 (O_573,N_9107,N_9391);
nor UO_574 (O_574,N_8958,N_8418);
nor UO_575 (O_575,N_9954,N_8064);
or UO_576 (O_576,N_7765,N_9530);
or UO_577 (O_577,N_8267,N_7717);
xnor UO_578 (O_578,N_9260,N_8015);
or UO_579 (O_579,N_7595,N_8526);
and UO_580 (O_580,N_8344,N_8734);
nor UO_581 (O_581,N_9585,N_9187);
nor UO_582 (O_582,N_8963,N_9417);
or UO_583 (O_583,N_8922,N_8119);
and UO_584 (O_584,N_8380,N_9339);
or UO_585 (O_585,N_9449,N_8569);
nand UO_586 (O_586,N_9932,N_9238);
or UO_587 (O_587,N_7868,N_9554);
nor UO_588 (O_588,N_8957,N_7646);
or UO_589 (O_589,N_7870,N_9146);
and UO_590 (O_590,N_9952,N_8954);
nor UO_591 (O_591,N_8980,N_9261);
nor UO_592 (O_592,N_7804,N_8783);
nand UO_593 (O_593,N_8381,N_7819);
nor UO_594 (O_594,N_8023,N_7682);
nor UO_595 (O_595,N_8880,N_9961);
and UO_596 (O_596,N_8898,N_8936);
and UO_597 (O_597,N_9480,N_8451);
nand UO_598 (O_598,N_8872,N_8118);
and UO_599 (O_599,N_8568,N_9606);
xnor UO_600 (O_600,N_9736,N_8762);
or UO_601 (O_601,N_8756,N_9402);
or UO_602 (O_602,N_9855,N_8660);
nor UO_603 (O_603,N_9921,N_8389);
or UO_604 (O_604,N_7561,N_9899);
or UO_605 (O_605,N_9835,N_9045);
and UO_606 (O_606,N_7887,N_9659);
and UO_607 (O_607,N_9053,N_8807);
nand UO_608 (O_608,N_8913,N_8686);
or UO_609 (O_609,N_9121,N_8442);
or UO_610 (O_610,N_7795,N_9263);
xor UO_611 (O_611,N_8554,N_9678);
nand UO_612 (O_612,N_8109,N_8070);
nor UO_613 (O_613,N_7824,N_9848);
nor UO_614 (O_614,N_7587,N_9059);
xor UO_615 (O_615,N_7683,N_9376);
or UO_616 (O_616,N_8371,N_7546);
xor UO_617 (O_617,N_7677,N_7786);
nand UO_618 (O_618,N_9110,N_9782);
or UO_619 (O_619,N_8570,N_8924);
nor UO_620 (O_620,N_7644,N_9564);
xnor UO_621 (O_621,N_8539,N_9701);
or UO_622 (O_622,N_7950,N_8616);
nor UO_623 (O_623,N_8785,N_7904);
and UO_624 (O_624,N_8249,N_8006);
xnor UO_625 (O_625,N_7743,N_9890);
xnor UO_626 (O_626,N_9451,N_8956);
and UO_627 (O_627,N_9104,N_9909);
or UO_628 (O_628,N_8709,N_7566);
or UO_629 (O_629,N_8540,N_8104);
nor UO_630 (O_630,N_9918,N_7643);
and UO_631 (O_631,N_7814,N_8942);
and UO_632 (O_632,N_8678,N_7825);
and UO_633 (O_633,N_8698,N_8282);
or UO_634 (O_634,N_8387,N_9607);
and UO_635 (O_635,N_7731,N_8820);
and UO_636 (O_636,N_9341,N_7593);
and UO_637 (O_637,N_9212,N_8086);
and UO_638 (O_638,N_9331,N_8161);
nand UO_639 (O_639,N_7729,N_9594);
or UO_640 (O_640,N_8587,N_8615);
or UO_641 (O_641,N_7921,N_7939);
xor UO_642 (O_642,N_9274,N_7894);
nor UO_643 (O_643,N_9199,N_9456);
xnor UO_644 (O_644,N_9969,N_9538);
and UO_645 (O_645,N_9149,N_8761);
and UO_646 (O_646,N_7629,N_9028);
nand UO_647 (O_647,N_9078,N_9039);
or UO_648 (O_648,N_7516,N_9088);
nand UO_649 (O_649,N_9922,N_9620);
or UO_650 (O_650,N_9996,N_8520);
and UO_651 (O_651,N_9912,N_9893);
xnor UO_652 (O_652,N_8203,N_8003);
nor UO_653 (O_653,N_7793,N_9252);
and UO_654 (O_654,N_8112,N_9007);
xnor UO_655 (O_655,N_7679,N_8559);
nand UO_656 (O_656,N_9729,N_7749);
or UO_657 (O_657,N_8259,N_9866);
xor UO_658 (O_658,N_9308,N_8817);
nor UO_659 (O_659,N_9660,N_9630);
nor UO_660 (O_660,N_8684,N_7774);
and UO_661 (O_661,N_9508,N_7738);
or UO_662 (O_662,N_9818,N_9536);
nand UO_663 (O_663,N_9162,N_8399);
xor UO_664 (O_664,N_7522,N_7891);
nand UO_665 (O_665,N_9639,N_9457);
nor UO_666 (O_666,N_9446,N_9235);
nand UO_667 (O_667,N_8524,N_8478);
or UO_668 (O_668,N_8592,N_7842);
xor UO_669 (O_669,N_8346,N_9629);
and UO_670 (O_670,N_8490,N_8450);
xnor UO_671 (O_671,N_7893,N_9504);
or UO_672 (O_672,N_9772,N_8350);
nand UO_673 (O_673,N_7736,N_8001);
nor UO_674 (O_674,N_7575,N_9498);
nand UO_675 (O_675,N_9445,N_9989);
xor UO_676 (O_676,N_8318,N_9013);
xor UO_677 (O_677,N_7665,N_8308);
nor UO_678 (O_678,N_7667,N_9725);
nand UO_679 (O_679,N_8590,N_8184);
nor UO_680 (O_680,N_9535,N_8862);
or UO_681 (O_681,N_8367,N_8799);
xor UO_682 (O_682,N_8536,N_8812);
nand UO_683 (O_683,N_7594,N_9776);
nor UO_684 (O_684,N_8549,N_9439);
xor UO_685 (O_685,N_8062,N_8117);
xnor UO_686 (O_686,N_8340,N_9634);
xor UO_687 (O_687,N_7874,N_7938);
xor UO_688 (O_688,N_9398,N_8411);
nor UO_689 (O_689,N_7865,N_9407);
or UO_690 (O_690,N_9442,N_8281);
nor UO_691 (O_691,N_9421,N_9422);
and UO_692 (O_692,N_8834,N_8829);
or UO_693 (O_693,N_8283,N_9453);
or UO_694 (O_694,N_9135,N_7762);
nand UO_695 (O_695,N_9378,N_9960);
and UO_696 (O_696,N_9427,N_9861);
nor UO_697 (O_697,N_8809,N_9562);
nand UO_698 (O_698,N_7773,N_8831);
xnor UO_699 (O_699,N_9455,N_7733);
xnor UO_700 (O_700,N_8237,N_7908);
xor UO_701 (O_701,N_7790,N_9882);
xor UO_702 (O_702,N_8315,N_8994);
xnor UO_703 (O_703,N_8147,N_8581);
nand UO_704 (O_704,N_8736,N_8575);
nand UO_705 (O_705,N_8031,N_8321);
nor UO_706 (O_706,N_7577,N_8882);
or UO_707 (O_707,N_9381,N_8830);
or UO_708 (O_708,N_8866,N_9765);
xnor UO_709 (O_709,N_9797,N_9844);
and UO_710 (O_710,N_9139,N_8888);
nand UO_711 (O_711,N_8565,N_7699);
nor UO_712 (O_712,N_9500,N_7769);
nand UO_713 (O_713,N_7582,N_8040);
xnor UO_714 (O_714,N_8272,N_9159);
and UO_715 (O_715,N_9406,N_7900);
and UO_716 (O_716,N_8484,N_9452);
xnor UO_717 (O_717,N_9175,N_9617);
xor UO_718 (O_718,N_8388,N_9964);
and UO_719 (O_719,N_8541,N_9547);
xnor UO_720 (O_720,N_9065,N_8627);
or UO_721 (O_721,N_9646,N_7585);
nand UO_722 (O_722,N_9241,N_9817);
nor UO_723 (O_723,N_9724,N_8427);
nor UO_724 (O_724,N_8084,N_9242);
or UO_725 (O_725,N_8986,N_9514);
and UO_726 (O_726,N_9679,N_8511);
nor UO_727 (O_727,N_8768,N_8468);
nand UO_728 (O_728,N_7928,N_8786);
and UO_729 (O_729,N_8416,N_8839);
xnor UO_730 (O_730,N_7760,N_8428);
nor UO_731 (O_731,N_7678,N_8314);
or UO_732 (O_732,N_7622,N_7539);
or UO_733 (O_733,N_9528,N_8675);
or UO_734 (O_734,N_7963,N_9408);
and UO_735 (O_735,N_7632,N_8854);
nand UO_736 (O_736,N_9767,N_7727);
and UO_737 (O_737,N_7601,N_8018);
nor UO_738 (O_738,N_7547,N_7757);
nand UO_739 (O_739,N_9192,N_7702);
nand UO_740 (O_740,N_7965,N_9685);
nor UO_741 (O_741,N_8522,N_7931);
or UO_742 (O_742,N_8606,N_9517);
nor UO_743 (O_743,N_8855,N_7837);
nor UO_744 (O_744,N_7603,N_9428);
or UO_745 (O_745,N_8032,N_9384);
xnor UO_746 (O_746,N_8065,N_9006);
nor UO_747 (O_747,N_7616,N_8928);
and UO_748 (O_748,N_9253,N_9553);
nand UO_749 (O_749,N_9734,N_8024);
nor UO_750 (O_750,N_8748,N_9642);
nand UO_751 (O_751,N_9036,N_8949);
xor UO_752 (O_752,N_9213,N_7635);
xnor UO_753 (O_753,N_8608,N_9218);
xnor UO_754 (O_754,N_7652,N_8679);
or UO_755 (O_755,N_8128,N_8137);
nor UO_756 (O_756,N_8206,N_9984);
nand UO_757 (O_757,N_9396,N_7709);
nand UO_758 (O_758,N_8557,N_7541);
and UO_759 (O_759,N_8483,N_8586);
or UO_760 (O_760,N_9026,N_8743);
and UO_761 (O_761,N_8665,N_9000);
and UO_762 (O_762,N_8183,N_7794);
nand UO_763 (O_763,N_8607,N_8754);
nor UO_764 (O_764,N_8274,N_9127);
nor UO_765 (O_765,N_8467,N_8596);
nand UO_766 (O_766,N_8648,N_9509);
nand UO_767 (O_767,N_8443,N_9831);
xnor UO_768 (O_768,N_7530,N_9798);
xnor UO_769 (O_769,N_8725,N_7876);
xor UO_770 (O_770,N_8978,N_9657);
or UO_771 (O_771,N_9492,N_7856);
and UO_772 (O_772,N_8300,N_8901);
nand UO_773 (O_773,N_7521,N_8082);
nand UO_774 (O_774,N_7920,N_9483);
nand UO_775 (O_775,N_8265,N_8885);
nand UO_776 (O_776,N_9741,N_9690);
xnor UO_777 (O_777,N_8164,N_8987);
xor UO_778 (O_778,N_7768,N_8372);
and UO_779 (O_779,N_9664,N_9737);
and UO_780 (O_780,N_9105,N_8584);
xnor UO_781 (O_781,N_8286,N_7895);
nor UO_782 (O_782,N_8662,N_8828);
nand UO_783 (O_783,N_7631,N_7966);
nand UO_784 (O_784,N_8507,N_8460);
and UO_785 (O_785,N_8093,N_7608);
nand UO_786 (O_786,N_8199,N_9496);
nor UO_787 (O_787,N_8532,N_8294);
nor UO_788 (O_788,N_7500,N_9383);
and UO_789 (O_789,N_9454,N_9115);
nor UO_790 (O_790,N_8937,N_8167);
xor UO_791 (O_791,N_8617,N_9551);
nand UO_792 (O_792,N_9834,N_8240);
nor UO_793 (O_793,N_8335,N_7624);
nor UO_794 (O_794,N_8055,N_7636);
nand UO_795 (O_795,N_9599,N_9132);
nand UO_796 (O_796,N_7525,N_8945);
nand UO_797 (O_797,N_9359,N_7889);
xnor UO_798 (O_798,N_9463,N_9616);
nand UO_799 (O_799,N_8612,N_8229);
nor UO_800 (O_800,N_8092,N_9953);
or UO_801 (O_801,N_9397,N_7951);
and UO_802 (O_802,N_8160,N_9191);
nand UO_803 (O_803,N_7799,N_7875);
xnor UO_804 (O_804,N_9622,N_9413);
or UO_805 (O_805,N_7813,N_9666);
nand UO_806 (O_806,N_7507,N_8035);
or UO_807 (O_807,N_7984,N_8863);
or UO_808 (O_808,N_8546,N_8027);
and UO_809 (O_809,N_9568,N_8733);
or UO_810 (O_810,N_9120,N_7693);
nor UO_811 (O_811,N_9050,N_8966);
or UO_812 (O_812,N_8309,N_9592);
nand UO_813 (O_813,N_8787,N_8688);
nor UO_814 (O_814,N_7820,N_8794);
xnor UO_815 (O_815,N_7543,N_9447);
nand UO_816 (O_816,N_9351,N_7728);
nor UO_817 (O_817,N_9839,N_7688);
or UO_818 (O_818,N_8489,N_9068);
xor UO_819 (O_819,N_9820,N_7997);
and UO_820 (O_820,N_8537,N_7627);
nor UO_821 (O_821,N_7691,N_9183);
nand UO_822 (O_822,N_9916,N_9570);
xnor UO_823 (O_823,N_8726,N_9268);
xor UO_824 (O_824,N_8000,N_8174);
and UO_825 (O_825,N_8345,N_8706);
and UO_826 (O_826,N_9392,N_8069);
nor UO_827 (O_827,N_9433,N_9887);
nor UO_828 (O_828,N_8593,N_9545);
or UO_829 (O_829,N_7501,N_7767);
and UO_830 (O_830,N_8329,N_9042);
or UO_831 (O_831,N_8120,N_9333);
or UO_832 (O_832,N_8822,N_7991);
xnor UO_833 (O_833,N_8057,N_8804);
or UO_834 (O_834,N_8746,N_8531);
or UO_835 (O_835,N_7533,N_9983);
xor UO_836 (O_836,N_9099,N_8896);
nor UO_837 (O_837,N_7748,N_8211);
nand UO_838 (O_838,N_8113,N_9179);
and UO_839 (O_839,N_7761,N_9878);
and UO_840 (O_840,N_8463,N_8322);
xnor UO_841 (O_841,N_9502,N_9419);
and UO_842 (O_842,N_9430,N_9981);
and UO_843 (O_843,N_7568,N_8439);
nor UO_844 (O_844,N_8333,N_7701);
or UO_845 (O_845,N_9332,N_9056);
or UO_846 (O_846,N_9524,N_8285);
xor UO_847 (O_847,N_9733,N_7737);
or UO_848 (O_848,N_7852,N_7739);
xor UO_849 (O_849,N_8707,N_9239);
and UO_850 (O_850,N_8437,N_9368);
nand UO_851 (O_851,N_9275,N_9745);
xnor UO_852 (O_852,N_9415,N_8798);
nand UO_853 (O_853,N_9259,N_8090);
and UO_854 (O_854,N_8471,N_8747);
nand UO_855 (O_855,N_7534,N_8646);
or UO_856 (O_856,N_8805,N_9490);
nand UO_857 (O_857,N_8670,N_9749);
nand UO_858 (O_858,N_8495,N_9823);
nand UO_859 (O_859,N_8030,N_9484);
xor UO_860 (O_860,N_7851,N_8585);
nand UO_861 (O_861,N_9712,N_8769);
or UO_862 (O_862,N_9438,N_8692);
nand UO_863 (O_863,N_9004,N_7751);
xor UO_864 (O_864,N_8251,N_7955);
nor UO_865 (O_865,N_9353,N_7975);
nor UO_866 (O_866,N_9673,N_7741);
xnor UO_867 (O_867,N_9169,N_7929);
or UO_868 (O_868,N_8297,N_9125);
and UO_869 (O_869,N_8353,N_9901);
xnor UO_870 (O_870,N_9738,N_8126);
and UO_871 (O_871,N_9414,N_9141);
nor UO_872 (O_872,N_8991,N_8008);
nor UO_873 (O_873,N_7755,N_9228);
nor UO_874 (O_874,N_8865,N_8651);
nor UO_875 (O_875,N_8702,N_8516);
nor UO_876 (O_876,N_9636,N_8528);
and UO_877 (O_877,N_7980,N_8066);
nor UO_878 (O_878,N_9716,N_7877);
nor UO_879 (O_879,N_8187,N_7906);
nor UO_880 (O_880,N_9147,N_8614);
nor UO_881 (O_881,N_7740,N_9011);
nand UO_882 (O_882,N_7960,N_8682);
nor UO_883 (O_883,N_9771,N_8207);
nor UO_884 (O_884,N_8740,N_7514);
nor UO_885 (O_885,N_8198,N_7506);
nor UO_886 (O_886,N_8737,N_8770);
and UO_887 (O_887,N_8445,N_7827);
xor UO_888 (O_888,N_9867,N_8629);
nor UO_889 (O_889,N_7989,N_7915);
and UO_890 (O_890,N_7578,N_8518);
or UO_891 (O_891,N_9236,N_7596);
or UO_892 (O_892,N_8816,N_8385);
nor UO_893 (O_893,N_7988,N_8572);
and UO_894 (O_894,N_7779,N_9073);
nand UO_895 (O_895,N_8639,N_7881);
and UO_896 (O_896,N_9762,N_8257);
nor UO_897 (O_897,N_8233,N_9448);
xnor UO_898 (O_898,N_9167,N_9166);
or UO_899 (O_899,N_8806,N_8500);
and UO_900 (O_900,N_7668,N_9902);
nand UO_901 (O_901,N_7519,N_7782);
xor UO_902 (O_902,N_7947,N_9544);
or UO_903 (O_903,N_8238,N_8622);
nand UO_904 (O_904,N_9214,N_8343);
nand UO_905 (O_905,N_8689,N_8644);
or UO_906 (O_906,N_9215,N_8982);
nand UO_907 (O_907,N_9373,N_8368);
or UO_908 (O_908,N_8363,N_9974);
nand UO_909 (O_909,N_8452,N_9653);
and UO_910 (O_910,N_8135,N_7502);
nor UO_911 (O_911,N_8457,N_8973);
xnor UO_912 (O_912,N_7796,N_8172);
nand UO_913 (O_913,N_7808,N_9434);
nor UO_914 (O_914,N_9076,N_8685);
and UO_915 (O_915,N_8613,N_8635);
xor UO_916 (O_916,N_8110,N_9003);
nor UO_917 (O_917,N_9041,N_9728);
and UO_918 (O_918,N_7744,N_8486);
or UO_919 (O_919,N_9751,N_9010);
nor UO_920 (O_920,N_9338,N_8379);
or UO_921 (O_921,N_8014,N_7905);
xor UO_922 (O_922,N_7992,N_9478);
nand UO_923 (O_923,N_9843,N_8276);
and UO_924 (O_924,N_7832,N_8143);
nor UO_925 (O_925,N_8044,N_8553);
and UO_926 (O_926,N_8841,N_9936);
nor UO_927 (O_927,N_8029,N_8395);
nand UO_928 (O_928,N_9148,N_7592);
nor UO_929 (O_929,N_7720,N_7957);
xor UO_930 (O_930,N_9829,N_9792);
xor UO_931 (O_931,N_7788,N_9061);
nand UO_932 (O_932,N_8103,N_8840);
nand UO_933 (O_933,N_9684,N_9354);
nor UO_934 (O_934,N_9990,N_9791);
nand UO_935 (O_935,N_8677,N_7619);
and UO_936 (O_936,N_7897,N_8021);
xnor UO_937 (O_937,N_8821,N_8303);
nor UO_938 (O_938,N_8168,N_9156);
or UO_939 (O_939,N_7946,N_9671);
nor UO_940 (O_940,N_9613,N_9991);
and UO_941 (O_941,N_9941,N_8856);
and UO_942 (O_942,N_9469,N_7642);
xnor UO_943 (O_943,N_8370,N_7828);
or UO_944 (O_944,N_8154,N_8643);
nor UO_945 (O_945,N_8562,N_9868);
nor UO_946 (O_946,N_8894,N_7685);
or UO_947 (O_947,N_8050,N_9281);
and UO_948 (O_948,N_8250,N_7783);
xor UO_949 (O_949,N_9997,N_7647);
or UO_950 (O_950,N_7598,N_8823);
nand UO_951 (O_951,N_8699,N_8576);
and UO_952 (O_952,N_7700,N_8254);
or UO_953 (O_953,N_8530,N_8366);
or UO_954 (O_954,N_7967,N_8672);
nand UO_955 (O_955,N_7858,N_9320);
nor UO_956 (O_956,N_8396,N_7922);
and UO_957 (O_957,N_9066,N_8578);
and UO_958 (O_958,N_8844,N_7570);
nor UO_959 (O_959,N_8138,N_8933);
nand UO_960 (O_960,N_7840,N_8932);
or UO_961 (O_961,N_8609,N_9850);
xor UO_962 (O_962,N_9513,N_9587);
nor UO_963 (O_963,N_8580,N_9904);
nand UO_964 (O_964,N_8405,N_8288);
nor UO_965 (O_965,N_8929,N_9386);
or UO_966 (O_966,N_9779,N_8710);
nand UO_967 (O_967,N_9366,N_7907);
and UO_968 (O_968,N_9142,N_9082);
nand UO_969 (O_969,N_9009,N_9216);
xor UO_970 (O_970,N_7787,N_7554);
nand UO_971 (O_971,N_8889,N_8943);
nand UO_972 (O_972,N_8292,N_8435);
and UO_973 (O_973,N_7878,N_9245);
and UO_974 (O_974,N_9493,N_8046);
nand UO_975 (O_975,N_9555,N_8157);
and UO_976 (O_976,N_8408,N_8657);
xor UO_977 (O_977,N_9204,N_8078);
nor UO_978 (O_978,N_8764,N_9521);
and UO_979 (O_979,N_9475,N_7885);
and UO_980 (O_980,N_8121,N_8873);
or UO_981 (O_981,N_9876,N_8407);
nor UO_982 (O_982,N_8504,N_9695);
nor UO_983 (O_983,N_8141,N_8990);
or UO_984 (O_984,N_9201,N_8464);
and UO_985 (O_985,N_9643,N_8631);
nand UO_986 (O_986,N_8998,N_8447);
xor UO_987 (O_987,N_7899,N_9752);
or UO_988 (O_988,N_7584,N_9704);
xor UO_989 (O_989,N_9327,N_7671);
nor UO_990 (O_990,N_9090,N_9595);
nand UO_991 (O_991,N_8231,N_9558);
or UO_992 (O_992,N_9786,N_9601);
xnor UO_993 (O_993,N_8177,N_9578);
xor UO_994 (O_994,N_8087,N_8253);
xor UO_995 (O_995,N_9717,N_8508);
nand UO_996 (O_996,N_7742,N_8626);
nand UO_997 (O_997,N_8603,N_8983);
nand UO_998 (O_998,N_9846,N_8425);
and UO_999 (O_999,N_9198,N_9518);
nand UO_1000 (O_1000,N_7971,N_8208);
xnor UO_1001 (O_1001,N_8583,N_8444);
and UO_1002 (O_1002,N_8215,N_8920);
nand UO_1003 (O_1003,N_9714,N_9917);
and UO_1004 (O_1004,N_9743,N_8204);
nor UO_1005 (O_1005,N_9207,N_8837);
xor UO_1006 (O_1006,N_8545,N_8278);
xnor UO_1007 (O_1007,N_7618,N_8940);
or UO_1008 (O_1008,N_8589,N_9608);
or UO_1009 (O_1009,N_9249,N_9650);
nor UO_1010 (O_1010,N_8714,N_8801);
nand UO_1011 (O_1011,N_8600,N_8716);
and UO_1012 (O_1012,N_8459,N_7886);
xor UO_1013 (O_1013,N_7770,N_7725);
or UO_1014 (O_1014,N_8995,N_8369);
and UO_1015 (O_1015,N_7675,N_9096);
or UO_1016 (O_1016,N_7532,N_9744);
nand UO_1017 (O_1017,N_8579,N_9597);
nand UO_1018 (O_1018,N_9806,N_7823);
nand UO_1019 (O_1019,N_8016,N_9335);
and UO_1020 (O_1020,N_8116,N_8260);
xnor UO_1021 (O_1021,N_9219,N_8191);
and UO_1022 (O_1022,N_8719,N_9370);
nand UO_1023 (O_1023,N_9674,N_9382);
xnor UO_1024 (O_1024,N_8124,N_8832);
or UO_1025 (O_1025,N_7658,N_9821);
nand UO_1026 (O_1026,N_9485,N_8148);
and UO_1027 (O_1027,N_9130,N_8563);
nor UO_1028 (O_1028,N_8099,N_8577);
and UO_1029 (O_1029,N_9652,N_8012);
xor UO_1030 (O_1030,N_9753,N_9098);
nor UO_1031 (O_1031,N_8628,N_7565);
and UO_1032 (O_1032,N_9966,N_9033);
and UO_1033 (O_1033,N_9231,N_8602);
or UO_1034 (O_1034,N_8200,N_9986);
nand UO_1035 (O_1035,N_7911,N_9377);
xnor UO_1036 (O_1036,N_9431,N_7710);
nand UO_1037 (O_1037,N_8188,N_9477);
nor UO_1038 (O_1038,N_8248,N_9522);
xor UO_1039 (O_1039,N_8967,N_8026);
or UO_1040 (O_1040,N_9400,N_8867);
nand UO_1041 (O_1041,N_9044,N_9461);
or UO_1042 (O_1042,N_8394,N_9841);
nand UO_1043 (O_1043,N_9692,N_9097);
or UO_1044 (O_1044,N_8156,N_8759);
nor UO_1045 (O_1045,N_7654,N_9618);
or UO_1046 (O_1046,N_7695,N_9665);
nand UO_1047 (O_1047,N_9468,N_8498);
and UO_1048 (O_1048,N_8721,N_8214);
xor UO_1049 (O_1049,N_9364,N_8656);
xor UO_1050 (O_1050,N_9845,N_7919);
and UO_1051 (O_1051,N_7564,N_9523);
nand UO_1052 (O_1052,N_9847,N_8717);
nand UO_1053 (O_1053,N_9262,N_9380);
and UO_1054 (O_1054,N_8843,N_9529);
xnor UO_1055 (O_1055,N_9356,N_8505);
xnor UO_1056 (O_1056,N_9586,N_9938);
nand UO_1057 (O_1057,N_7581,N_8287);
nand UO_1058 (O_1058,N_9375,N_8296);
and UO_1059 (O_1059,N_9550,N_8219);
and UO_1060 (O_1060,N_8218,N_7659);
nor UO_1061 (O_1061,N_9510,N_9310);
or UO_1062 (O_1062,N_9247,N_8232);
xor UO_1063 (O_1063,N_8197,N_8028);
xor UO_1064 (O_1064,N_8778,N_9853);
xor UO_1065 (O_1065,N_7872,N_9537);
xor UO_1066 (O_1066,N_9988,N_8189);
or UO_1067 (O_1067,N_8226,N_7569);
xnor UO_1068 (O_1068,N_7903,N_7625);
or UO_1069 (O_1069,N_8146,N_9619);
and UO_1070 (O_1070,N_8163,N_8195);
or UO_1071 (O_1071,N_9324,N_9352);
xor UO_1072 (O_1072,N_9070,N_8328);
nor UO_1073 (O_1073,N_9302,N_9051);
nor UO_1074 (O_1074,N_9757,N_9102);
nand UO_1075 (O_1075,N_9101,N_7528);
nand UO_1076 (O_1076,N_8695,N_7657);
xnor UO_1077 (O_1077,N_9687,N_8319);
nor UO_1078 (O_1078,N_8802,N_8727);
nor UO_1079 (O_1079,N_8063,N_8851);
or UO_1080 (O_1080,N_7816,N_9824);
or UO_1081 (O_1081,N_8838,N_8384);
nand UO_1082 (O_1082,N_9849,N_8186);
nand UO_1083 (O_1083,N_9699,N_9604);
nand UO_1084 (O_1084,N_9057,N_7918);
and UO_1085 (O_1085,N_9603,N_8114);
nor UO_1086 (O_1086,N_8351,N_8728);
or UO_1087 (O_1087,N_9200,N_9032);
and UO_1088 (O_1088,N_7803,N_7933);
and UO_1089 (O_1089,N_8320,N_9987);
nor UO_1090 (O_1090,N_8236,N_9093);
xor UO_1091 (O_1091,N_8290,N_7810);
and UO_1092 (O_1092,N_7520,N_7981);
xnor UO_1093 (O_1093,N_8426,N_8891);
nand UO_1094 (O_1094,N_9277,N_8178);
or UO_1095 (O_1095,N_7863,N_9248);
or UO_1096 (O_1096,N_9896,N_8194);
xnor UO_1097 (O_1097,N_7734,N_8139);
nand UO_1098 (O_1098,N_9225,N_8419);
xnor UO_1099 (O_1099,N_9137,N_9286);
xor UO_1100 (O_1100,N_9865,N_8947);
or UO_1101 (O_1101,N_7524,N_9085);
and UO_1102 (O_1102,N_7944,N_9133);
nand UO_1103 (O_1103,N_7822,N_9112);
xor UO_1104 (O_1104,N_8680,N_9561);
xnor UO_1105 (O_1105,N_9254,N_9658);
nand UO_1106 (O_1106,N_9412,N_9576);
and UO_1107 (O_1107,N_9140,N_9035);
nand UO_1108 (O_1108,N_9519,N_8598);
or UO_1109 (O_1109,N_9813,N_7607);
xor UO_1110 (O_1110,N_8722,N_8974);
xor UO_1111 (O_1111,N_9977,N_8960);
and UO_1112 (O_1112,N_9046,N_8715);
xnor UO_1113 (O_1113,N_7513,N_9721);
nand UO_1114 (O_1114,N_7600,N_7712);
nand UO_1115 (O_1115,N_9067,N_8952);
and UO_1116 (O_1116,N_7586,N_8392);
xor UO_1117 (O_1117,N_9325,N_9635);
nor UO_1118 (O_1118,N_9072,N_9495);
and UO_1119 (O_1119,N_7948,N_9672);
nor UO_1120 (O_1120,N_9602,N_8140);
xnor UO_1121 (O_1121,N_8859,N_7704);
xor UO_1122 (O_1122,N_8201,N_9923);
or UO_1123 (O_1123,N_7732,N_7590);
and UO_1124 (O_1124,N_7843,N_9778);
or UO_1125 (O_1125,N_9329,N_9029);
nand UO_1126 (O_1126,N_8131,N_7763);
or UO_1127 (O_1127,N_7993,N_8703);
nand UO_1128 (O_1128,N_8650,N_7576);
nand UO_1129 (O_1129,N_9574,N_9662);
nor UO_1130 (O_1130,N_7932,N_8676);
or UO_1131 (O_1131,N_7936,N_9266);
nand UO_1132 (O_1132,N_8732,N_8011);
xnor UO_1133 (O_1133,N_7560,N_9950);
nor UO_1134 (O_1134,N_9326,N_9173);
nand UO_1135 (O_1135,N_8269,N_7609);
nor UO_1136 (O_1136,N_8910,N_7855);
nor UO_1137 (O_1137,N_8127,N_8359);
or UO_1138 (O_1138,N_8968,N_8360);
or UO_1139 (O_1139,N_8108,N_9907);
and UO_1140 (O_1140,N_7718,N_9418);
and UO_1141 (O_1141,N_9885,N_8311);
nand UO_1142 (O_1142,N_9211,N_8564);
nand UO_1143 (O_1143,N_9424,N_8071);
xnor UO_1144 (O_1144,N_9860,N_7934);
or UO_1145 (O_1145,N_9934,N_9486);
xnor UO_1146 (O_1146,N_9312,N_7639);
or UO_1147 (O_1147,N_9897,N_7531);
nand UO_1148 (O_1148,N_8301,N_7523);
and UO_1149 (O_1149,N_7690,N_9022);
or UO_1150 (O_1150,N_9503,N_9316);
nand UO_1151 (O_1151,N_9911,N_8153);
or UO_1152 (O_1152,N_7935,N_8386);
xnor UO_1153 (O_1153,N_9925,N_9935);
nor UO_1154 (O_1154,N_8170,N_9789);
xor UO_1155 (O_1155,N_9060,N_7634);
and UO_1156 (O_1156,N_7754,N_7663);
xor UO_1157 (O_1157,N_9830,N_9403);
or UO_1158 (O_1158,N_8348,N_9648);
nand UO_1159 (O_1159,N_9328,N_8664);
nand UO_1160 (O_1160,N_8323,N_9047);
or UO_1161 (O_1161,N_7983,N_9688);
nor UO_1162 (O_1162,N_9501,N_9367);
nor UO_1163 (O_1163,N_9605,N_9947);
xor UO_1164 (O_1164,N_8424,N_8776);
and UO_1165 (O_1165,N_9343,N_8893);
and UO_1166 (O_1166,N_8097,N_9012);
and UO_1167 (O_1167,N_7778,N_9631);
nor UO_1168 (O_1168,N_7942,N_9337);
or UO_1169 (O_1169,N_8033,N_9290);
nand UO_1170 (O_1170,N_8868,N_8339);
or UO_1171 (O_1171,N_9374,N_8414);
xnor UO_1172 (O_1172,N_8305,N_8083);
xor UO_1173 (O_1173,N_9730,N_9579);
or UO_1174 (O_1174,N_9429,N_9693);
xor UO_1175 (O_1175,N_8818,N_9390);
nand UO_1176 (O_1176,N_9506,N_8944);
nand UO_1177 (O_1177,N_7716,N_7550);
and UO_1178 (O_1178,N_9058,N_9401);
nor UO_1179 (O_1179,N_8789,N_8299);
nor UO_1180 (O_1180,N_9804,N_9565);
nand UO_1181 (O_1181,N_8784,N_8538);
and UO_1182 (O_1182,N_8245,N_9369);
nor UO_1183 (O_1183,N_9567,N_7923);
xor UO_1184 (O_1184,N_8620,N_8244);
xor UO_1185 (O_1185,N_7735,N_9924);
nor UO_1186 (O_1186,N_9289,N_9450);
and UO_1187 (O_1187,N_9229,N_8067);
or UO_1188 (O_1188,N_9614,N_7597);
and UO_1189 (O_1189,N_8970,N_8313);
nand UO_1190 (O_1190,N_9992,N_8336);
and UO_1191 (O_1191,N_9189,N_7996);
or UO_1192 (O_1192,N_8781,N_8663);
xnor UO_1193 (O_1193,N_8152,N_9040);
nand UO_1194 (O_1194,N_9676,N_8247);
nand UO_1195 (O_1195,N_8058,N_9272);
nor UO_1196 (O_1196,N_9543,N_8166);
xnor UO_1197 (O_1197,N_8525,N_8921);
nor UO_1198 (O_1198,N_7706,N_9706);
or UO_1199 (O_1199,N_9244,N_8653);
or UO_1200 (O_1200,N_9856,N_9494);
nor UO_1201 (O_1201,N_9269,N_9330);
xnor UO_1202 (O_1202,N_7580,N_9892);
xor UO_1203 (O_1203,N_8455,N_8744);
xor UO_1204 (O_1204,N_8378,N_8193);
nand UO_1205 (O_1205,N_8738,N_9271);
nand UO_1206 (O_1206,N_8079,N_9273);
and UO_1207 (O_1207,N_9913,N_8661);
nor UO_1208 (O_1208,N_9319,N_9573);
xnor UO_1209 (O_1209,N_7880,N_8997);
nand UO_1210 (O_1210,N_8502,N_9756);
xnor UO_1211 (O_1211,N_7661,N_7844);
or UO_1212 (O_1212,N_7721,N_9336);
nor UO_1213 (O_1213,N_8597,N_9560);
or UO_1214 (O_1214,N_9251,N_8724);
or UO_1215 (O_1215,N_8107,N_9655);
xor UO_1216 (O_1216,N_8415,N_9217);
nor UO_1217 (O_1217,N_8263,N_8595);
xnor UO_1218 (O_1218,N_8499,N_9299);
xor UO_1219 (O_1219,N_8610,N_9443);
nor UO_1220 (O_1220,N_9487,N_8325);
nor UO_1221 (O_1221,N_9903,N_7990);
and UO_1222 (O_1222,N_7557,N_9971);
nor UO_1223 (O_1223,N_9344,N_9670);
xor UO_1224 (O_1224,N_7697,N_9822);
and UO_1225 (O_1225,N_9889,N_9432);
or UO_1226 (O_1226,N_9001,N_7637);
or UO_1227 (O_1227,N_7745,N_8213);
and UO_1228 (O_1228,N_7882,N_9296);
or UO_1229 (O_1229,N_9552,N_8846);
or UO_1230 (O_1230,N_7676,N_8095);
xnor UO_1231 (O_1231,N_9195,N_8382);
or UO_1232 (O_1232,N_8731,N_9958);
xor UO_1233 (O_1233,N_8697,N_7860);
nor UO_1234 (O_1234,N_9054,N_8474);
or UO_1235 (O_1235,N_8019,N_9812);
xnor UO_1236 (O_1236,N_7873,N_8241);
or UO_1237 (O_1237,N_9471,N_9154);
or UO_1238 (O_1238,N_7776,N_8446);
xnor UO_1239 (O_1239,N_9002,N_9711);
xor UO_1240 (O_1240,N_8869,N_8911);
xor UO_1241 (O_1241,N_7511,N_9210);
nand UO_1242 (O_1242,N_8599,N_8476);
nand UO_1243 (O_1243,N_8758,N_9948);
nor UO_1244 (O_1244,N_7792,N_8542);
xnor UO_1245 (O_1245,N_9656,N_9423);
or UO_1246 (O_1246,N_8521,N_8242);
nand UO_1247 (O_1247,N_8422,N_9425);
nand UO_1248 (O_1248,N_9615,N_7853);
xnor UO_1249 (O_1249,N_8708,N_8210);
or UO_1250 (O_1250,N_8039,N_8904);
nor UO_1251 (O_1251,N_8279,N_8383);
or UO_1252 (O_1252,N_9405,N_8526);
nand UO_1253 (O_1253,N_8404,N_9349);
and UO_1254 (O_1254,N_7723,N_9745);
nor UO_1255 (O_1255,N_7624,N_8422);
or UO_1256 (O_1256,N_9622,N_9519);
nand UO_1257 (O_1257,N_7586,N_7665);
nor UO_1258 (O_1258,N_9855,N_9741);
or UO_1259 (O_1259,N_8922,N_9377);
xnor UO_1260 (O_1260,N_8200,N_9553);
or UO_1261 (O_1261,N_8520,N_9015);
or UO_1262 (O_1262,N_9351,N_8296);
nand UO_1263 (O_1263,N_9413,N_9781);
xnor UO_1264 (O_1264,N_7938,N_9234);
nand UO_1265 (O_1265,N_8812,N_9349);
xor UO_1266 (O_1266,N_8790,N_8046);
and UO_1267 (O_1267,N_7680,N_9891);
nor UO_1268 (O_1268,N_8334,N_9622);
and UO_1269 (O_1269,N_7627,N_8867);
nor UO_1270 (O_1270,N_9365,N_8810);
nand UO_1271 (O_1271,N_9743,N_9420);
nor UO_1272 (O_1272,N_9245,N_9210);
nor UO_1273 (O_1273,N_8862,N_8651);
nand UO_1274 (O_1274,N_8802,N_9100);
and UO_1275 (O_1275,N_9701,N_8306);
nor UO_1276 (O_1276,N_8772,N_8661);
and UO_1277 (O_1277,N_9830,N_9926);
nor UO_1278 (O_1278,N_9601,N_9529);
nor UO_1279 (O_1279,N_9762,N_7744);
nor UO_1280 (O_1280,N_7899,N_9374);
nand UO_1281 (O_1281,N_9521,N_8682);
or UO_1282 (O_1282,N_8497,N_9982);
nor UO_1283 (O_1283,N_9787,N_7970);
nor UO_1284 (O_1284,N_7700,N_8588);
nor UO_1285 (O_1285,N_8214,N_9603);
xnor UO_1286 (O_1286,N_9883,N_8406);
xor UO_1287 (O_1287,N_9033,N_9967);
nand UO_1288 (O_1288,N_9043,N_9665);
nand UO_1289 (O_1289,N_9794,N_8683);
nand UO_1290 (O_1290,N_8097,N_8189);
nor UO_1291 (O_1291,N_8042,N_9032);
or UO_1292 (O_1292,N_8598,N_9505);
and UO_1293 (O_1293,N_7801,N_8078);
or UO_1294 (O_1294,N_9348,N_8798);
nand UO_1295 (O_1295,N_7794,N_8590);
nand UO_1296 (O_1296,N_8303,N_8500);
nor UO_1297 (O_1297,N_7554,N_8867);
nor UO_1298 (O_1298,N_8591,N_7586);
nor UO_1299 (O_1299,N_8228,N_9261);
nor UO_1300 (O_1300,N_9275,N_9565);
xor UO_1301 (O_1301,N_8519,N_7518);
xor UO_1302 (O_1302,N_7623,N_7601);
nand UO_1303 (O_1303,N_9823,N_8490);
or UO_1304 (O_1304,N_7590,N_9102);
nor UO_1305 (O_1305,N_7853,N_8604);
xor UO_1306 (O_1306,N_7773,N_9766);
nor UO_1307 (O_1307,N_7662,N_8163);
nor UO_1308 (O_1308,N_9990,N_7989);
nor UO_1309 (O_1309,N_7516,N_9815);
xnor UO_1310 (O_1310,N_7948,N_8095);
or UO_1311 (O_1311,N_9466,N_9291);
and UO_1312 (O_1312,N_8380,N_8816);
or UO_1313 (O_1313,N_8082,N_9635);
xor UO_1314 (O_1314,N_8726,N_8530);
xor UO_1315 (O_1315,N_9204,N_9901);
or UO_1316 (O_1316,N_9493,N_9219);
xnor UO_1317 (O_1317,N_9833,N_9504);
xnor UO_1318 (O_1318,N_8123,N_8701);
nand UO_1319 (O_1319,N_7920,N_8810);
and UO_1320 (O_1320,N_9855,N_7838);
nand UO_1321 (O_1321,N_9934,N_9006);
and UO_1322 (O_1322,N_9116,N_8771);
and UO_1323 (O_1323,N_9968,N_9072);
xor UO_1324 (O_1324,N_9328,N_8753);
nand UO_1325 (O_1325,N_9659,N_9837);
xnor UO_1326 (O_1326,N_7936,N_8425);
or UO_1327 (O_1327,N_8572,N_8656);
and UO_1328 (O_1328,N_7632,N_8677);
and UO_1329 (O_1329,N_9255,N_9980);
xnor UO_1330 (O_1330,N_8092,N_9469);
and UO_1331 (O_1331,N_9883,N_7731);
or UO_1332 (O_1332,N_7510,N_8795);
nand UO_1333 (O_1333,N_9141,N_8945);
nand UO_1334 (O_1334,N_8793,N_8327);
nand UO_1335 (O_1335,N_7713,N_7881);
xnor UO_1336 (O_1336,N_9813,N_9216);
and UO_1337 (O_1337,N_9938,N_7838);
nor UO_1338 (O_1338,N_8858,N_7534);
or UO_1339 (O_1339,N_8057,N_8566);
xor UO_1340 (O_1340,N_7782,N_8197);
xnor UO_1341 (O_1341,N_7788,N_9422);
nor UO_1342 (O_1342,N_9627,N_8361);
and UO_1343 (O_1343,N_8888,N_8587);
nand UO_1344 (O_1344,N_9963,N_8329);
nor UO_1345 (O_1345,N_8017,N_8793);
or UO_1346 (O_1346,N_8581,N_7785);
xor UO_1347 (O_1347,N_9444,N_8028);
or UO_1348 (O_1348,N_8789,N_8969);
xnor UO_1349 (O_1349,N_8658,N_8520);
nand UO_1350 (O_1350,N_9132,N_8055);
nand UO_1351 (O_1351,N_7980,N_9426);
nand UO_1352 (O_1352,N_8352,N_9272);
nand UO_1353 (O_1353,N_8609,N_8935);
nor UO_1354 (O_1354,N_7570,N_9931);
or UO_1355 (O_1355,N_9368,N_7798);
or UO_1356 (O_1356,N_9076,N_9245);
xor UO_1357 (O_1357,N_9305,N_9498);
nand UO_1358 (O_1358,N_8868,N_7778);
xor UO_1359 (O_1359,N_9437,N_8432);
and UO_1360 (O_1360,N_9906,N_9554);
nor UO_1361 (O_1361,N_7666,N_9550);
or UO_1362 (O_1362,N_7812,N_8321);
and UO_1363 (O_1363,N_8437,N_8562);
xnor UO_1364 (O_1364,N_9589,N_7647);
nand UO_1365 (O_1365,N_9070,N_8425);
nand UO_1366 (O_1366,N_9397,N_9969);
nand UO_1367 (O_1367,N_8054,N_9389);
and UO_1368 (O_1368,N_9528,N_8938);
nand UO_1369 (O_1369,N_9712,N_9394);
xnor UO_1370 (O_1370,N_8819,N_9620);
or UO_1371 (O_1371,N_8347,N_8463);
and UO_1372 (O_1372,N_8195,N_9167);
or UO_1373 (O_1373,N_8122,N_9707);
and UO_1374 (O_1374,N_7642,N_7712);
xor UO_1375 (O_1375,N_7920,N_7735);
nand UO_1376 (O_1376,N_7538,N_8152);
nor UO_1377 (O_1377,N_8172,N_8827);
nor UO_1378 (O_1378,N_8995,N_7882);
nand UO_1379 (O_1379,N_9489,N_8106);
nor UO_1380 (O_1380,N_7753,N_8298);
nand UO_1381 (O_1381,N_8885,N_8242);
nand UO_1382 (O_1382,N_7793,N_9549);
or UO_1383 (O_1383,N_9906,N_7635);
nand UO_1384 (O_1384,N_9287,N_9086);
nor UO_1385 (O_1385,N_9108,N_9218);
and UO_1386 (O_1386,N_9042,N_9138);
or UO_1387 (O_1387,N_8699,N_8424);
nand UO_1388 (O_1388,N_8891,N_8194);
nor UO_1389 (O_1389,N_9335,N_9854);
nor UO_1390 (O_1390,N_9548,N_8362);
nor UO_1391 (O_1391,N_8911,N_9654);
nand UO_1392 (O_1392,N_7696,N_7783);
and UO_1393 (O_1393,N_9162,N_9564);
nand UO_1394 (O_1394,N_9444,N_9633);
xnor UO_1395 (O_1395,N_8454,N_8185);
nor UO_1396 (O_1396,N_9587,N_7592);
or UO_1397 (O_1397,N_8930,N_7683);
xor UO_1398 (O_1398,N_8737,N_8253);
and UO_1399 (O_1399,N_7672,N_8438);
xnor UO_1400 (O_1400,N_9076,N_7704);
and UO_1401 (O_1401,N_8966,N_9905);
or UO_1402 (O_1402,N_7905,N_8367);
or UO_1403 (O_1403,N_9834,N_9682);
nor UO_1404 (O_1404,N_8152,N_8673);
nand UO_1405 (O_1405,N_9898,N_9419);
or UO_1406 (O_1406,N_7893,N_8751);
xor UO_1407 (O_1407,N_7552,N_9376);
xnor UO_1408 (O_1408,N_8685,N_8472);
or UO_1409 (O_1409,N_9269,N_8235);
nor UO_1410 (O_1410,N_9930,N_7580);
or UO_1411 (O_1411,N_9653,N_9181);
nand UO_1412 (O_1412,N_7772,N_9628);
and UO_1413 (O_1413,N_8911,N_7713);
or UO_1414 (O_1414,N_8357,N_9795);
and UO_1415 (O_1415,N_8277,N_7551);
and UO_1416 (O_1416,N_9618,N_7916);
nand UO_1417 (O_1417,N_7805,N_8112);
nand UO_1418 (O_1418,N_9652,N_7665);
nand UO_1419 (O_1419,N_9859,N_8880);
or UO_1420 (O_1420,N_8795,N_9900);
or UO_1421 (O_1421,N_9936,N_9595);
nand UO_1422 (O_1422,N_7566,N_7523);
nand UO_1423 (O_1423,N_9901,N_8617);
and UO_1424 (O_1424,N_8642,N_8221);
nor UO_1425 (O_1425,N_9835,N_9934);
nor UO_1426 (O_1426,N_9503,N_9423);
nand UO_1427 (O_1427,N_9308,N_9918);
and UO_1428 (O_1428,N_7804,N_8972);
xor UO_1429 (O_1429,N_9158,N_8059);
nand UO_1430 (O_1430,N_7628,N_8511);
or UO_1431 (O_1431,N_9054,N_7936);
and UO_1432 (O_1432,N_8484,N_8735);
nand UO_1433 (O_1433,N_8466,N_8396);
nand UO_1434 (O_1434,N_7628,N_7642);
xor UO_1435 (O_1435,N_7512,N_9339);
nand UO_1436 (O_1436,N_9385,N_9476);
or UO_1437 (O_1437,N_7767,N_9859);
and UO_1438 (O_1438,N_8037,N_7642);
nor UO_1439 (O_1439,N_8582,N_8003);
nor UO_1440 (O_1440,N_7801,N_7996);
and UO_1441 (O_1441,N_7845,N_8886);
and UO_1442 (O_1442,N_9759,N_8429);
nand UO_1443 (O_1443,N_8689,N_8526);
nand UO_1444 (O_1444,N_9518,N_9132);
xnor UO_1445 (O_1445,N_8804,N_8459);
nand UO_1446 (O_1446,N_9323,N_7940);
nor UO_1447 (O_1447,N_8027,N_9150);
xor UO_1448 (O_1448,N_7505,N_8301);
or UO_1449 (O_1449,N_8631,N_9629);
or UO_1450 (O_1450,N_8699,N_8834);
xnor UO_1451 (O_1451,N_9228,N_8828);
nand UO_1452 (O_1452,N_9468,N_9975);
or UO_1453 (O_1453,N_9734,N_7588);
xnor UO_1454 (O_1454,N_8888,N_9493);
xor UO_1455 (O_1455,N_8287,N_9728);
nand UO_1456 (O_1456,N_9133,N_9173);
xnor UO_1457 (O_1457,N_7879,N_8841);
and UO_1458 (O_1458,N_8131,N_8672);
or UO_1459 (O_1459,N_9354,N_8364);
nand UO_1460 (O_1460,N_8502,N_8691);
xnor UO_1461 (O_1461,N_9201,N_8442);
and UO_1462 (O_1462,N_9813,N_7827);
and UO_1463 (O_1463,N_9390,N_8297);
xor UO_1464 (O_1464,N_9001,N_9497);
or UO_1465 (O_1465,N_9607,N_7890);
nor UO_1466 (O_1466,N_7805,N_7528);
nor UO_1467 (O_1467,N_8339,N_9840);
nor UO_1468 (O_1468,N_9598,N_9621);
nor UO_1469 (O_1469,N_8979,N_8981);
nor UO_1470 (O_1470,N_9167,N_8009);
and UO_1471 (O_1471,N_8333,N_8416);
and UO_1472 (O_1472,N_9261,N_9486);
and UO_1473 (O_1473,N_9013,N_8782);
nor UO_1474 (O_1474,N_7858,N_8533);
nand UO_1475 (O_1475,N_7811,N_8137);
nor UO_1476 (O_1476,N_8232,N_9116);
nand UO_1477 (O_1477,N_8797,N_8025);
nand UO_1478 (O_1478,N_9501,N_8527);
and UO_1479 (O_1479,N_9381,N_8443);
nor UO_1480 (O_1480,N_7629,N_8313);
or UO_1481 (O_1481,N_9527,N_8148);
nor UO_1482 (O_1482,N_9577,N_8120);
nand UO_1483 (O_1483,N_8003,N_8263);
and UO_1484 (O_1484,N_8866,N_8447);
and UO_1485 (O_1485,N_8962,N_9398);
nand UO_1486 (O_1486,N_9483,N_9537);
or UO_1487 (O_1487,N_9382,N_9419);
nand UO_1488 (O_1488,N_8230,N_8171);
xnor UO_1489 (O_1489,N_7962,N_8911);
nand UO_1490 (O_1490,N_7732,N_8149);
nor UO_1491 (O_1491,N_9901,N_9054);
nand UO_1492 (O_1492,N_8718,N_7513);
nor UO_1493 (O_1493,N_8257,N_8041);
nor UO_1494 (O_1494,N_9946,N_8541);
and UO_1495 (O_1495,N_8006,N_7913);
or UO_1496 (O_1496,N_9125,N_9472);
nand UO_1497 (O_1497,N_8200,N_7976);
or UO_1498 (O_1498,N_8510,N_8851);
nand UO_1499 (O_1499,N_8531,N_9532);
endmodule