module basic_2500_25000_3000_100_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_2396,In_912);
and U1 (N_1,In_887,In_1368);
nand U2 (N_2,In_1265,In_1065);
or U3 (N_3,In_1603,In_1191);
nand U4 (N_4,In_2476,In_545);
nand U5 (N_5,In_125,In_1294);
nor U6 (N_6,In_1116,In_1559);
nand U7 (N_7,In_480,In_5);
nor U8 (N_8,In_1066,In_2091);
nor U9 (N_9,In_72,In_90);
xor U10 (N_10,In_614,In_1822);
or U11 (N_11,In_2159,In_2236);
xnor U12 (N_12,In_306,In_1354);
xnor U13 (N_13,In_1879,In_2481);
nor U14 (N_14,In_670,In_376);
or U15 (N_15,In_2232,In_487);
or U16 (N_16,In_560,In_1496);
and U17 (N_17,In_1119,In_1159);
xnor U18 (N_18,In_2062,In_463);
nand U19 (N_19,In_536,In_707);
or U20 (N_20,In_1273,In_1322);
or U21 (N_21,In_2467,In_158);
nor U22 (N_22,In_394,In_1769);
nor U23 (N_23,In_2187,In_2449);
nor U24 (N_24,In_1490,In_289);
nand U25 (N_25,In_797,In_593);
xnor U26 (N_26,In_613,In_1782);
nor U27 (N_27,In_984,In_246);
nor U28 (N_28,In_1804,In_419);
nand U29 (N_29,In_1149,In_83);
nand U30 (N_30,In_1777,In_1564);
or U31 (N_31,In_553,In_1009);
or U32 (N_32,In_335,In_1724);
and U33 (N_33,In_1300,In_2233);
and U34 (N_34,In_227,In_2344);
nor U35 (N_35,In_546,In_464);
and U36 (N_36,In_492,In_2147);
and U37 (N_37,In_1403,In_1834);
and U38 (N_38,In_2371,In_1378);
nor U39 (N_39,In_95,In_2193);
and U40 (N_40,In_1685,In_247);
nor U41 (N_41,In_2443,In_819);
nand U42 (N_42,In_344,In_2409);
nand U43 (N_43,In_1594,In_347);
and U44 (N_44,In_368,In_273);
nand U45 (N_45,In_589,In_2380);
nor U46 (N_46,In_1121,In_652);
xor U47 (N_47,In_407,In_1589);
nor U48 (N_48,In_115,In_1889);
and U49 (N_49,In_1142,In_513);
xor U50 (N_50,In_2411,In_1721);
nor U51 (N_51,In_937,In_333);
and U52 (N_52,In_2199,In_2336);
and U53 (N_53,In_11,In_506);
nor U54 (N_54,In_216,In_688);
xor U55 (N_55,In_1468,In_1506);
nand U56 (N_56,In_1775,In_2305);
xnor U57 (N_57,In_1420,In_734);
or U58 (N_58,In_811,In_1745);
and U59 (N_59,In_638,In_1931);
nand U60 (N_60,In_1946,In_1276);
nor U61 (N_61,In_387,In_2417);
and U62 (N_62,In_565,In_1209);
xnor U63 (N_63,In_99,In_2494);
nor U64 (N_64,In_918,In_1023);
nand U65 (N_65,In_852,In_1076);
nor U66 (N_66,In_1038,In_1759);
and U67 (N_67,In_2266,In_2331);
nand U68 (N_68,In_214,In_980);
nand U69 (N_69,In_906,In_2247);
xnor U70 (N_70,In_346,In_436);
or U71 (N_71,In_1188,In_1874);
or U72 (N_72,In_2402,In_1047);
xnor U73 (N_73,In_1622,In_1366);
nand U74 (N_74,In_1839,In_1585);
xnor U75 (N_75,In_1351,In_1082);
nand U76 (N_76,In_1958,In_1203);
nor U77 (N_77,In_1825,In_1566);
nor U78 (N_78,In_1174,In_975);
or U79 (N_79,In_248,In_371);
nand U80 (N_80,In_1957,In_1591);
nor U81 (N_81,In_2095,In_2017);
and U82 (N_82,In_1990,In_1331);
or U83 (N_83,In_1906,In_988);
and U84 (N_84,In_1033,In_2030);
or U85 (N_85,In_2073,In_29);
or U86 (N_86,In_1155,In_266);
nand U87 (N_87,In_1270,In_1424);
xnor U88 (N_88,In_2262,In_1080);
or U89 (N_89,In_1233,In_233);
and U90 (N_90,In_1667,In_449);
or U91 (N_91,In_2210,In_26);
and U92 (N_92,In_2018,In_1676);
nand U93 (N_93,In_448,In_1752);
or U94 (N_94,In_1445,In_1235);
nand U95 (N_95,In_1211,In_1079);
xor U96 (N_96,In_524,In_1637);
nand U97 (N_97,In_2157,In_2106);
nor U98 (N_98,In_2016,In_2052);
nor U99 (N_99,In_869,In_610);
or U100 (N_100,In_821,In_178);
xnor U101 (N_101,In_615,In_1458);
nand U102 (N_102,In_262,In_1640);
nand U103 (N_103,In_786,In_1212);
or U104 (N_104,In_804,In_1588);
and U105 (N_105,In_213,In_129);
and U106 (N_106,In_114,In_2067);
nand U107 (N_107,In_986,In_2351);
nor U108 (N_108,In_1706,In_588);
nor U109 (N_109,In_2303,In_679);
nand U110 (N_110,In_1720,In_102);
nand U111 (N_111,In_1465,In_663);
or U112 (N_112,In_1198,In_1753);
and U113 (N_113,In_2107,In_894);
or U114 (N_114,In_1476,In_2403);
nor U115 (N_115,In_1395,In_2288);
and U116 (N_116,In_1578,In_417);
or U117 (N_117,In_1840,In_2113);
and U118 (N_118,In_2181,In_82);
xor U119 (N_119,In_101,In_2272);
xor U120 (N_120,In_1884,In_1606);
or U121 (N_121,In_330,In_951);
nor U122 (N_122,In_279,In_2466);
nor U123 (N_123,In_985,In_633);
xnor U124 (N_124,In_677,In_2340);
or U125 (N_125,In_369,In_559);
nor U126 (N_126,In_594,In_2094);
or U127 (N_127,In_1538,In_1166);
xor U128 (N_128,In_1767,In_1976);
xnor U129 (N_129,In_1678,In_2065);
nand U130 (N_130,In_1671,In_1213);
nor U131 (N_131,In_1712,In_2369);
nor U132 (N_132,In_37,In_982);
xnor U133 (N_133,In_2333,In_1916);
nand U134 (N_134,In_1050,In_1519);
xnor U135 (N_135,In_789,In_162);
xor U136 (N_136,In_85,In_56);
xor U137 (N_137,In_1075,In_923);
xor U138 (N_138,In_310,In_1470);
nor U139 (N_139,In_485,In_317);
nor U140 (N_140,In_1197,In_1857);
nor U141 (N_141,In_699,In_32);
xor U142 (N_142,In_359,In_2455);
xor U143 (N_143,In_622,In_2381);
or U144 (N_144,In_1972,In_1117);
and U145 (N_145,In_2156,In_1224);
and U146 (N_146,In_584,In_378);
and U147 (N_147,In_254,In_733);
or U148 (N_148,In_98,In_1450);
and U149 (N_149,In_2472,In_864);
nor U150 (N_150,In_1711,In_1567);
nand U151 (N_151,In_899,In_857);
nand U152 (N_152,In_2451,In_316);
or U153 (N_153,In_1878,In_1434);
nor U154 (N_154,In_2043,In_851);
xnor U155 (N_155,In_399,In_1120);
nor U156 (N_156,In_483,In_785);
nand U157 (N_157,In_2424,In_1865);
nor U158 (N_158,In_278,In_1995);
or U159 (N_159,In_805,In_49);
nor U160 (N_160,In_2061,In_1391);
and U161 (N_161,In_1560,In_2273);
and U162 (N_162,In_1126,In_2454);
nor U163 (N_163,In_2323,In_1245);
or U164 (N_164,In_61,In_1094);
nand U165 (N_165,In_2141,In_1084);
nand U166 (N_166,In_598,In_2002);
or U167 (N_167,In_1828,In_1305);
xor U168 (N_168,In_653,In_184);
nor U169 (N_169,In_1702,In_916);
nand U170 (N_170,In_146,In_166);
or U171 (N_171,In_1493,In_211);
nor U172 (N_172,In_625,In_2335);
xnor U173 (N_173,In_435,In_837);
nor U174 (N_174,In_323,In_2475);
or U175 (N_175,In_2037,In_1697);
xnor U176 (N_176,In_1859,In_1230);
and U177 (N_177,In_2484,In_462);
xor U178 (N_178,In_1337,In_277);
xor U179 (N_179,In_958,In_749);
and U180 (N_180,In_430,In_1202);
or U181 (N_181,In_2050,In_640);
and U182 (N_182,In_36,In_1272);
and U183 (N_183,In_960,In_282);
nand U184 (N_184,In_511,In_1993);
and U185 (N_185,In_2020,In_2346);
xnor U186 (N_186,In_533,In_840);
xor U187 (N_187,In_401,In_1815);
xor U188 (N_188,In_603,In_1456);
and U189 (N_189,In_1217,In_2469);
nor U190 (N_190,In_798,In_697);
nor U191 (N_191,In_2334,In_484);
and U192 (N_192,In_2308,In_68);
nor U193 (N_193,In_2418,In_2122);
nand U194 (N_194,In_2332,In_1442);
nor U195 (N_195,In_2234,In_1801);
and U196 (N_196,In_1500,In_41);
and U197 (N_197,In_2006,In_1784);
and U198 (N_198,In_1414,In_2063);
or U199 (N_199,In_362,In_1162);
and U200 (N_200,In_104,In_2169);
nand U201 (N_201,In_966,In_1572);
nand U202 (N_202,In_1242,In_826);
xor U203 (N_203,In_2230,In_2040);
nor U204 (N_204,In_1048,In_2162);
nand U205 (N_205,In_1817,In_1942);
and U206 (N_206,In_885,In_744);
nand U207 (N_207,In_915,In_1021);
nand U208 (N_208,In_1809,In_1133);
xor U209 (N_209,In_949,In_1997);
xor U210 (N_210,In_2220,In_926);
xnor U211 (N_211,In_1173,In_1694);
nand U212 (N_212,In_507,In_2263);
nand U213 (N_213,In_1415,In_1365);
and U214 (N_214,In_2450,In_551);
nor U215 (N_215,In_2367,In_212);
and U216 (N_216,In_1948,In_1803);
and U217 (N_217,In_1228,In_2176);
or U218 (N_218,In_1737,In_1317);
nand U219 (N_219,In_1798,In_757);
nand U220 (N_220,In_2019,In_291);
xnor U221 (N_221,In_1347,In_538);
nand U222 (N_222,In_205,In_2049);
and U223 (N_223,In_1900,In_1915);
xor U224 (N_224,In_112,In_1912);
xor U225 (N_225,In_909,In_249);
xor U226 (N_226,In_1306,In_220);
nand U227 (N_227,In_1432,In_1200);
nand U228 (N_228,In_1169,In_1604);
and U229 (N_229,In_421,In_2183);
or U230 (N_230,In_2201,In_735);
nor U231 (N_231,In_111,In_1841);
xnor U232 (N_232,In_2286,In_2491);
or U233 (N_233,In_1049,In_658);
nor U234 (N_234,In_2296,In_694);
nor U235 (N_235,In_2120,In_929);
nor U236 (N_236,In_1304,In_1123);
and U237 (N_237,In_1639,In_952);
and U238 (N_238,In_1073,In_2311);
or U239 (N_239,In_157,In_1967);
xor U240 (N_240,In_1507,In_423);
and U241 (N_241,In_1708,In_324);
or U242 (N_242,In_2459,In_763);
and U243 (N_243,In_1582,In_428);
nand U244 (N_244,In_1316,In_1619);
nand U245 (N_245,In_606,In_6);
and U246 (N_246,In_2393,In_1569);
nand U247 (N_247,In_1428,In_2100);
xnor U248 (N_248,In_2027,In_8);
nor U249 (N_249,In_534,In_139);
and U250 (N_250,In_1014,In_1314);
xor U251 (N_251,N_185,In_1945);
xor U252 (N_252,In_2190,In_126);
nand U253 (N_253,In_1182,In_1805);
nand U254 (N_254,In_396,In_119);
nor U255 (N_255,In_2170,N_22);
xnor U256 (N_256,In_1446,In_74);
nand U257 (N_257,In_877,In_1590);
nand U258 (N_258,In_1218,In_1061);
nand U259 (N_259,In_683,In_835);
or U260 (N_260,In_1486,In_2322);
and U261 (N_261,In_645,In_1747);
nor U262 (N_262,In_1959,In_81);
or U263 (N_263,In_2026,In_1894);
or U264 (N_264,In_669,In_2284);
nor U265 (N_265,In_71,In_1430);
or U266 (N_266,In_1729,In_742);
nand U267 (N_267,In_1779,N_89);
nand U268 (N_268,In_758,In_176);
nor U269 (N_269,In_451,In_294);
nand U270 (N_270,In_1345,In_2225);
xnor U271 (N_271,In_1029,In_1616);
nand U272 (N_272,In_1373,In_712);
or U273 (N_273,N_60,In_107);
or U274 (N_274,N_178,In_1105);
xnor U275 (N_275,In_860,In_202);
xnor U276 (N_276,In_833,In_849);
nand U277 (N_277,In_1516,In_1277);
and U278 (N_278,In_561,In_526);
and U279 (N_279,N_235,In_1215);
nor U280 (N_280,In_341,In_2434);
and U281 (N_281,N_224,In_935);
xnor U282 (N_282,In_179,N_82);
xnor U283 (N_283,N_138,In_285);
nand U284 (N_284,In_2138,In_321);
nand U285 (N_285,In_1668,In_1342);
or U286 (N_286,In_1303,In_2264);
and U287 (N_287,In_716,N_113);
xnor U288 (N_288,In_1013,In_263);
nand U289 (N_289,In_2196,In_1835);
xor U290 (N_290,In_940,In_818);
or U291 (N_291,In_802,In_732);
xnor U292 (N_292,In_1515,In_2300);
xor U293 (N_293,N_26,In_2295);
nand U294 (N_294,In_838,N_62);
or U295 (N_295,In_1248,In_384);
or U296 (N_296,In_1576,In_1307);
nor U297 (N_297,In_365,In_635);
nand U298 (N_298,In_180,In_810);
nor U299 (N_299,In_741,In_1106);
xnor U300 (N_300,In_1006,In_1214);
and U301 (N_301,In_468,In_1689);
and U302 (N_302,In_259,In_327);
xnor U303 (N_303,In_412,In_236);
nor U304 (N_304,N_100,In_9);
nor U305 (N_305,In_895,In_116);
nand U306 (N_306,In_34,In_163);
nor U307 (N_307,In_1330,In_1807);
and U308 (N_308,In_238,In_1164);
and U309 (N_309,In_1963,N_226);
nor U310 (N_310,In_1943,In_1960);
nand U311 (N_311,N_114,In_284);
or U312 (N_312,In_972,N_165);
nor U313 (N_313,In_1249,In_1707);
xor U314 (N_314,In_2143,In_499);
xor U315 (N_315,In_1498,In_928);
or U316 (N_316,N_131,In_2306);
nor U317 (N_317,In_1356,In_557);
xor U318 (N_318,In_1362,In_1986);
nor U319 (N_319,In_491,In_1101);
nand U320 (N_320,In_2109,In_2146);
xnor U321 (N_321,In_1260,In_2289);
and U322 (N_322,In_2088,In_1229);
nand U323 (N_323,In_340,N_55);
and U324 (N_324,In_2310,In_2128);
nor U325 (N_325,In_400,In_772);
nand U326 (N_326,In_1573,In_2328);
or U327 (N_327,In_320,In_824);
nand U328 (N_328,In_634,N_48);
or U329 (N_329,In_2205,In_908);
nand U330 (N_330,In_67,In_2123);
or U331 (N_331,In_1624,In_188);
or U332 (N_332,In_1687,N_161);
nand U333 (N_333,In_1544,In_914);
or U334 (N_334,In_866,In_977);
nor U335 (N_335,In_1978,In_1222);
xnor U336 (N_336,N_32,N_85);
xor U337 (N_337,In_1469,In_2487);
or U338 (N_338,In_173,In_1238);
nor U339 (N_339,In_1231,In_2389);
xnor U340 (N_340,N_162,In_135);
nor U341 (N_341,In_121,In_486);
xor U342 (N_342,In_1757,N_180);
or U343 (N_343,In_2226,In_1453);
nor U344 (N_344,In_1172,In_1971);
xnor U345 (N_345,In_1291,In_2250);
nand U346 (N_346,In_275,In_1413);
nand U347 (N_347,In_207,In_2330);
xnor U348 (N_348,In_1298,N_140);
and U349 (N_349,In_383,In_611);
xor U350 (N_350,In_717,In_631);
nand U351 (N_351,In_905,In_309);
xor U352 (N_352,N_78,In_1299);
or U353 (N_353,In_1384,In_444);
xor U354 (N_354,In_2244,N_188);
nor U355 (N_355,In_1041,In_1400);
and U356 (N_356,In_2421,In_968);
nor U357 (N_357,In_608,In_825);
xnor U358 (N_358,In_1151,In_252);
and U359 (N_359,In_2337,In_39);
nand U360 (N_360,In_1633,In_527);
and U361 (N_361,In_1359,In_1241);
nand U362 (N_362,In_1353,In_1856);
or U363 (N_363,In_2066,In_1389);
xor U364 (N_364,In_1081,N_73);
or U365 (N_365,In_702,In_358);
and U366 (N_366,In_239,In_1657);
or U367 (N_367,In_1367,In_2178);
nor U368 (N_368,N_119,In_1071);
or U369 (N_369,In_1137,In_953);
xnor U370 (N_370,In_2203,N_7);
or U371 (N_371,N_237,In_865);
nor U372 (N_372,In_411,In_1929);
or U373 (N_373,In_2252,N_47);
xnor U374 (N_374,In_172,In_846);
or U375 (N_375,In_2212,In_427);
xnor U376 (N_376,In_1695,In_801);
and U377 (N_377,In_1053,In_1794);
or U378 (N_378,In_145,In_2297);
xnor U379 (N_379,In_404,In_1054);
and U380 (N_380,In_1800,In_222);
and U381 (N_381,In_841,In_2057);
xor U382 (N_382,In_1766,In_646);
xnor U383 (N_383,In_1148,N_77);
and U384 (N_384,In_1332,In_1600);
nor U385 (N_385,In_1692,In_2285);
nor U386 (N_386,N_171,In_676);
xor U387 (N_387,In_1964,In_446);
and U388 (N_388,In_2348,In_675);
nand U389 (N_389,In_662,In_2327);
nand U390 (N_390,In_2082,N_44);
nand U391 (N_391,In_1275,In_142);
or U392 (N_392,In_1321,N_49);
xor U393 (N_393,In_1909,In_2111);
nand U394 (N_394,In_872,In_965);
nor U395 (N_395,In_52,In_47);
nand U396 (N_396,N_191,In_87);
and U397 (N_397,In_1930,In_410);
or U398 (N_398,In_547,N_193);
and U399 (N_399,In_2011,In_1833);
nor U400 (N_400,In_265,In_1472);
or U401 (N_401,In_1717,In_153);
and U402 (N_402,In_1181,In_1927);
and U403 (N_403,In_217,In_1672);
and U404 (N_404,In_2188,In_1141);
xor U405 (N_405,In_433,In_1765);
and U406 (N_406,In_1178,In_1495);
xnor U407 (N_407,In_2189,In_2084);
nor U408 (N_408,In_2268,In_979);
xor U409 (N_409,In_2426,In_503);
and U410 (N_410,In_1998,In_1962);
and U411 (N_411,In_1240,In_1683);
and U412 (N_412,In_2116,In_504);
or U413 (N_413,In_567,In_947);
or U414 (N_414,In_1327,In_1966);
nor U415 (N_415,In_693,In_1393);
or U416 (N_416,In_779,In_445);
or U417 (N_417,In_151,In_1301);
and U418 (N_418,In_1131,In_437);
xnor U419 (N_419,In_727,In_1183);
nor U420 (N_420,N_1,In_815);
nor U421 (N_421,In_592,In_2153);
xnor U422 (N_422,In_493,In_454);
nor U423 (N_423,In_16,In_1280);
xor U424 (N_424,In_570,In_1690);
nor U425 (N_425,In_475,In_164);
and U426 (N_426,In_1501,In_1858);
nand U427 (N_427,N_247,In_1074);
or U428 (N_428,In_1187,In_175);
nor U429 (N_429,In_4,In_1411);
or U430 (N_430,In_2053,In_1713);
and U431 (N_431,In_50,In_1550);
or U432 (N_432,In_2179,In_692);
nor U433 (N_433,In_2208,In_1190);
or U434 (N_434,In_1237,In_1487);
and U435 (N_435,In_269,In_373);
xnor U436 (N_436,N_220,In_245);
xor U437 (N_437,N_132,In_1620);
or U438 (N_438,In_2241,In_1044);
or U439 (N_439,In_1263,In_1919);
nor U440 (N_440,In_1226,In_1602);
nor U441 (N_441,In_1661,In_1677);
and U442 (N_442,In_1019,In_1264);
nand U443 (N_443,In_1644,In_1059);
or U444 (N_444,N_167,In_2145);
nor U445 (N_445,In_230,In_1360);
xor U446 (N_446,In_1449,In_124);
and U447 (N_447,In_1768,In_349);
xnor U448 (N_448,In_1004,In_1503);
xnor U449 (N_449,In_1246,In_256);
nor U450 (N_450,In_1455,In_1095);
nand U451 (N_451,In_374,In_709);
xor U452 (N_452,In_2152,In_1091);
or U453 (N_453,In_264,In_505);
nor U454 (N_454,In_2461,In_60);
or U455 (N_455,In_495,In_1103);
and U456 (N_456,In_2001,N_5);
nor U457 (N_457,In_432,In_1781);
xor U458 (N_458,In_1176,In_1999);
or U459 (N_459,In_1823,In_2407);
xnor U460 (N_460,N_81,In_2090);
nand U461 (N_461,In_209,In_260);
nor U462 (N_462,In_889,In_1087);
and U463 (N_463,In_1611,In_668);
or U464 (N_464,In_2173,In_1529);
or U465 (N_465,In_719,In_876);
nor U466 (N_466,In_1466,In_2445);
or U467 (N_467,In_1489,In_1494);
xor U468 (N_468,In_2240,In_2320);
nand U469 (N_469,In_1189,In_2359);
xnor U470 (N_470,In_600,N_65);
xnor U471 (N_471,In_2379,In_2175);
nor U472 (N_472,In_1666,In_415);
and U473 (N_473,In_1205,In_408);
nand U474 (N_474,In_429,In_1016);
and U475 (N_475,N_205,In_2126);
or U476 (N_476,In_1113,N_108);
nor U477 (N_477,In_957,In_1583);
xnor U478 (N_478,In_1135,N_186);
or U479 (N_479,In_1975,In_59);
and U480 (N_480,In_2495,In_1742);
and U481 (N_481,In_2114,N_66);
and U482 (N_482,In_1813,In_568);
and U483 (N_483,In_453,In_1847);
or U484 (N_484,In_2158,N_18);
or U485 (N_485,N_39,In_791);
and U486 (N_486,In_2474,In_2185);
nand U487 (N_487,In_460,N_8);
nand U488 (N_488,In_1089,N_51);
nor U489 (N_489,In_878,In_1836);
xor U490 (N_490,In_353,In_440);
nor U491 (N_491,In_1531,N_166);
and U492 (N_492,In_155,In_235);
xnor U493 (N_493,In_2343,In_258);
nand U494 (N_494,In_1398,In_542);
and U495 (N_495,In_808,In_2161);
nor U496 (N_496,In_1618,In_2204);
and U497 (N_497,In_1920,In_131);
nor U498 (N_498,In_2257,In_416);
nor U499 (N_499,N_120,In_579);
nand U500 (N_500,In_2243,In_711);
nor U501 (N_501,In_1227,N_347);
and U502 (N_502,In_1905,In_2197);
nor U503 (N_503,In_1001,N_143);
and U504 (N_504,In_186,In_689);
or U505 (N_505,N_245,In_736);
nand U506 (N_506,In_1743,In_470);
and U507 (N_507,N_12,In_1848);
nor U508 (N_508,N_345,N_295);
nor U509 (N_509,In_1281,In_386);
or U510 (N_510,N_472,In_969);
nor U511 (N_511,In_1820,In_1705);
and U512 (N_512,In_686,N_266);
nor U513 (N_513,In_2290,N_197);
nand U514 (N_514,In_234,N_462);
and U515 (N_515,N_71,In_1612);
nand U516 (N_516,In_1419,In_1508);
nor U517 (N_517,In_389,N_152);
nor U518 (N_518,In_1534,N_84);
xor U519 (N_519,In_739,In_1402);
nor U520 (N_520,In_893,In_1027);
and U521 (N_521,N_11,In_1568);
and U522 (N_522,In_2293,In_192);
or U523 (N_523,In_1448,In_954);
nand U524 (N_524,In_2039,In_1150);
nor U525 (N_525,In_515,In_992);
nand U526 (N_526,In_1541,In_2214);
and U527 (N_527,In_612,In_14);
xnor U528 (N_528,N_377,In_51);
xor U529 (N_529,In_1806,In_671);
and U530 (N_530,In_2267,In_2355);
nor U531 (N_531,N_398,N_335);
nand U532 (N_532,In_932,In_1830);
nand U533 (N_533,In_1436,In_2042);
and U534 (N_534,In_1899,In_1130);
and U535 (N_535,In_1429,In_1372);
nor U536 (N_536,In_927,N_305);
and U537 (N_537,In_587,In_1554);
nor U538 (N_538,In_44,In_363);
nand U539 (N_539,In_2438,In_1882);
nand U540 (N_540,In_601,In_2352);
nand U541 (N_541,N_499,In_2465);
or U542 (N_542,In_73,In_974);
nand U543 (N_543,In_1532,N_225);
and U544 (N_544,In_331,In_1870);
and U545 (N_545,In_620,In_590);
nor U546 (N_546,In_1326,In_1463);
xnor U547 (N_547,In_2433,In_406);
nand U548 (N_548,In_117,In_334);
and U549 (N_549,In_2081,In_618);
and U550 (N_550,In_762,In_1952);
nand U551 (N_551,In_725,In_1947);
nor U552 (N_552,N_149,In_1621);
or U553 (N_553,In_2075,In_226);
xnor U554 (N_554,In_2304,In_641);
xnor U555 (N_555,In_143,In_1158);
nand U556 (N_556,In_150,In_760);
nand U557 (N_557,N_83,N_471);
nand U558 (N_558,In_1346,In_197);
nand U559 (N_559,N_470,In_619);
nor U560 (N_560,In_65,In_883);
nor U561 (N_561,In_842,N_336);
or U562 (N_562,In_1871,N_323);
nand U563 (N_563,In_200,In_1867);
xor U564 (N_564,In_1147,N_111);
or U565 (N_565,In_1736,In_170);
nor U566 (N_566,In_1787,In_704);
nand U567 (N_567,N_413,In_75);
nand U568 (N_568,In_286,In_1934);
nor U569 (N_569,In_783,In_1908);
or U570 (N_570,N_133,In_1850);
nor U571 (N_571,In_628,N_151);
xor U572 (N_572,In_86,In_1669);
nand U573 (N_573,In_1545,N_391);
nand U574 (N_574,In_575,N_268);
or U575 (N_575,In_1996,In_1634);
xnor U576 (N_576,In_1156,In_1040);
xnor U577 (N_577,In_1379,In_223);
or U578 (N_578,In_723,In_2416);
xor U579 (N_579,In_766,N_277);
and U580 (N_580,In_2350,In_2047);
nor U581 (N_581,In_1396,N_194);
and U582 (N_582,In_409,In_133);
and U583 (N_583,In_474,In_1427);
nand U584 (N_584,N_182,In_2054);
nor U585 (N_585,In_2098,In_1649);
or U586 (N_586,N_289,In_2253);
xor U587 (N_587,N_353,In_183);
or U588 (N_588,N_374,In_301);
and U589 (N_589,In_1407,In_759);
nand U590 (N_590,In_701,In_288);
or U591 (N_591,In_2174,N_362);
xnor U592 (N_592,In_420,In_1517);
xor U593 (N_593,In_2388,N_414);
and U594 (N_594,In_2238,In_1987);
and U595 (N_595,In_447,N_256);
nand U596 (N_596,In_1112,N_38);
and U597 (N_597,N_80,In_1361);
nor U598 (N_598,In_198,In_1723);
nor U599 (N_599,In_1570,In_1928);
xor U600 (N_600,In_946,In_1864);
nand U601 (N_601,N_361,In_2014);
or U602 (N_602,N_418,N_179);
and U603 (N_603,In_995,N_204);
and U604 (N_604,In_1623,N_358);
xor U605 (N_605,In_1063,In_2420);
nand U606 (N_606,In_830,In_1923);
nor U607 (N_607,In_647,In_2093);
or U608 (N_608,N_96,In_461);
or U609 (N_609,In_1898,In_2423);
nor U610 (N_610,In_1881,In_1981);
nor U611 (N_611,In_1153,In_544);
or U612 (N_612,In_1730,N_33);
nor U613 (N_613,In_2432,In_1286);
and U614 (N_614,In_576,N_246);
xor U615 (N_615,In_2021,In_70);
or U616 (N_616,In_721,In_1308);
nand U617 (N_617,In_599,In_1944);
nand U618 (N_618,In_745,In_514);
xor U619 (N_619,In_581,In_2033);
xor U620 (N_620,N_468,In_731);
nor U621 (N_621,N_206,In_2029);
and U622 (N_622,In_750,In_1399);
nand U623 (N_623,In_1510,In_2485);
xnor U624 (N_624,In_438,In_1002);
xnor U625 (N_625,N_433,In_1418);
nand U626 (N_626,N_259,In_1645);
and U627 (N_627,In_1108,In_244);
xor U628 (N_628,In_1579,In_2307);
or U629 (N_629,In_1785,N_285);
nor U630 (N_630,N_387,In_1557);
xor U631 (N_631,In_970,N_463);
xor U632 (N_632,N_300,N_415);
nand U633 (N_633,N_292,In_580);
xnor U634 (N_634,N_208,In_1334);
nor U635 (N_635,In_512,In_1271);
and U636 (N_636,In_397,In_1447);
or U637 (N_637,In_516,N_331);
nand U638 (N_638,N_200,N_69);
nor U639 (N_639,In_1643,In_398);
or U640 (N_640,N_407,N_190);
and U641 (N_641,In_2319,N_322);
xnor U642 (N_642,In_103,In_1581);
nand U643 (N_643,In_1526,In_528);
nand U644 (N_644,N_192,N_341);
nand U645 (N_645,In_1390,In_1175);
nor U646 (N_646,In_998,In_1844);
and U647 (N_647,In_1363,In_1406);
nand U648 (N_648,N_442,In_1292);
nand U649 (N_649,N_283,N_213);
nor U650 (N_650,In_1994,In_767);
or U651 (N_651,In_1979,In_890);
nand U652 (N_652,In_1461,In_521);
and U653 (N_653,In_535,In_1780);
nor U654 (N_654,In_78,In_469);
nand U655 (N_655,In_270,In_299);
nand U656 (N_656,In_775,N_352);
or U657 (N_657,In_636,In_1253);
and U658 (N_658,In_2256,In_1911);
nand U659 (N_659,In_403,In_1816);
xnor U660 (N_660,In_1225,In_1970);
xnor U661 (N_661,In_1134,In_687);
xnor U662 (N_662,In_1058,N_37);
nor U663 (N_663,In_122,N_464);
or U664 (N_664,N_242,N_492);
or U665 (N_665,In_232,In_439);
xnor U666 (N_666,In_1686,In_2104);
and U667 (N_667,In_1549,In_1208);
nand U668 (N_668,In_769,In_1348);
nand U669 (N_669,N_371,In_621);
xnor U670 (N_670,In_1323,In_1481);
and U671 (N_671,N_31,In_654);
or U672 (N_672,In_1017,In_1344);
and U673 (N_673,In_1680,In_1656);
nor U674 (N_674,In_1206,In_1262);
nor U675 (N_675,In_459,In_706);
nand U676 (N_676,In_2397,In_2038);
xor U677 (N_677,In_1132,In_191);
nand U678 (N_678,N_394,N_209);
nor U679 (N_679,In_1479,In_1746);
and U680 (N_680,In_473,N_455);
and U681 (N_681,In_2492,In_814);
xnor U682 (N_682,In_267,N_373);
or U683 (N_683,N_129,In_481);
or U684 (N_684,In_1845,In_990);
or U685 (N_685,In_1954,In_181);
xnor U686 (N_686,In_754,In_2480);
or U687 (N_687,In_2194,In_639);
and U688 (N_688,In_1732,In_1937);
xor U689 (N_689,In_123,N_339);
nor U690 (N_690,N_260,N_426);
or U691 (N_691,In_1437,In_2068);
nor U692 (N_692,In_2326,In_917);
or U693 (N_693,In_298,N_489);
xnor U694 (N_694,In_1552,In_2059);
or U695 (N_695,In_728,In_2493);
xnor U696 (N_696,In_2276,In_1851);
and U697 (N_697,In_168,In_2324);
or U698 (N_698,In_859,N_284);
or U699 (N_699,N_153,N_301);
xor U700 (N_700,In_2048,In_2406);
or U701 (N_701,In_1247,In_1145);
or U702 (N_702,In_756,In_2374);
nand U703 (N_703,In_1821,In_868);
or U704 (N_704,In_1922,In_2349);
and U705 (N_705,In_962,In_185);
and U706 (N_706,In_53,In_1630);
and U707 (N_707,In_690,N_447);
and U708 (N_708,In_944,In_1558);
xor U709 (N_709,In_2209,In_167);
nor U710 (N_710,In_160,In_0);
and U711 (N_711,In_1735,In_2237);
nand U712 (N_712,N_482,In_2488);
and U713 (N_713,In_691,In_569);
xnor U714 (N_714,N_404,In_1778);
xnor U715 (N_715,In_2118,In_1122);
and U716 (N_716,N_264,In_318);
nor U717 (N_717,In_1868,In_1693);
or U718 (N_718,In_1764,In_2136);
or U719 (N_719,In_1802,In_1528);
xnor U720 (N_720,In_782,In_2121);
or U721 (N_721,In_2012,In_2294);
or U722 (N_722,In_2182,In_1163);
xor U723 (N_723,N_431,N_118);
and U724 (N_724,In_1154,In_1170);
and U725 (N_725,In_770,In_271);
nor U726 (N_726,In_159,In_2092);
xnor U727 (N_727,In_1477,In_1381);
xor U728 (N_728,In_1797,In_891);
xnor U729 (N_729,In_963,In_1636);
xnor U730 (N_730,N_357,N_249);
nand U731 (N_731,In_605,N_170);
nor U732 (N_732,In_790,In_747);
nand U733 (N_733,In_708,In_792);
or U734 (N_734,In_596,In_1386);
and U735 (N_735,In_2004,In_660);
nand U736 (N_736,In_356,In_1941);
nand U737 (N_737,In_1042,In_1938);
nand U738 (N_738,N_380,In_1674);
xor U739 (N_739,N_173,In_1926);
or U740 (N_740,In_981,N_479);
and U741 (N_741,In_1290,In_1914);
xor U742 (N_742,In_1110,In_2132);
nor U743 (N_743,In_2497,In_920);
nor U744 (N_744,In_1796,In_2404);
nand U745 (N_745,N_104,In_2435);
nor U746 (N_746,In_1977,N_435);
nor U747 (N_747,N_320,N_223);
nor U748 (N_748,In_623,In_15);
and U749 (N_749,In_276,N_313);
nor U750 (N_750,In_1654,In_888);
nand U751 (N_751,In_740,N_746);
xor U752 (N_752,In_2382,In_1547);
and U753 (N_753,In_391,In_1548);
and U754 (N_754,In_360,In_566);
and U755 (N_755,In_1635,N_396);
nor U756 (N_756,N_702,In_1614);
or U757 (N_757,In_1625,N_325);
or U758 (N_758,In_154,N_98);
nor U759 (N_759,In_1497,In_304);
xnor U760 (N_760,In_1282,In_2456);
and U761 (N_761,In_18,In_1223);
nor U762 (N_762,N_465,In_405);
and U763 (N_763,In_1641,In_1056);
or U764 (N_764,N_139,N_551);
or U765 (N_765,In_1725,In_1030);
xor U766 (N_766,N_544,In_2395);
xnor U767 (N_767,In_1514,In_1255);
nand U768 (N_768,In_1936,In_366);
nand U769 (N_769,In_2140,In_1374);
and U770 (N_770,In_1460,In_1935);
and U771 (N_771,N_24,N_16);
nor U772 (N_772,In_2287,In_2058);
and U773 (N_773,In_1340,In_229);
nor U774 (N_774,N_265,N_685);
or U775 (N_775,N_267,In_77);
nor U776 (N_776,In_1293,In_897);
xor U777 (N_777,N_717,N_660);
and U778 (N_778,In_466,In_2154);
and U779 (N_779,In_934,In_650);
and U780 (N_780,N_282,N_488);
and U781 (N_781,N_692,In_2164);
nor U782 (N_782,N_737,N_724);
and U783 (N_783,In_482,In_1201);
nor U784 (N_784,N_662,N_439);
and U785 (N_785,N_422,In_203);
xor U786 (N_786,In_283,In_1257);
and U787 (N_787,In_999,In_377);
xor U788 (N_788,In_812,In_171);
nor U789 (N_789,N_20,In_1258);
nand U790 (N_790,N_262,N_368);
and U791 (N_791,In_1599,In_293);
xor U792 (N_792,In_1026,N_728);
nor U793 (N_793,In_2329,In_1907);
and U794 (N_794,In_1741,N_696);
nand U795 (N_795,N_695,N_593);
nor U796 (N_796,N_272,In_1086);
xor U797 (N_797,N_23,In_983);
xnor U798 (N_798,In_637,N_523);
nor U799 (N_799,N_704,In_773);
xor U800 (N_800,In_1774,In_255);
nor U801 (N_801,In_2315,In_221);
xnor U802 (N_802,In_1259,N_667);
xnor U803 (N_803,In_455,In_1571);
xor U804 (N_804,In_1595,In_1733);
or U805 (N_805,In_563,In_1580);
and U806 (N_806,In_393,In_2361);
nor U807 (N_807,N_416,In_1003);
and U808 (N_808,In_1933,N_681);
xor U809 (N_809,N_70,N_560);
nand U810 (N_810,In_2227,In_136);
nand U811 (N_811,In_2207,In_2448);
and U812 (N_812,In_2453,N_579);
or U813 (N_813,In_2171,N_258);
xnor U814 (N_814,N_533,In_395);
or U815 (N_815,In_661,In_931);
nor U816 (N_816,In_2139,N_713);
and U817 (N_817,In_870,N_508);
nor U818 (N_818,In_1903,In_2215);
nand U819 (N_819,In_1837,In_414);
nor U820 (N_820,In_147,In_319);
or U821 (N_821,In_795,N_437);
and U822 (N_822,In_1055,N_734);
nor U823 (N_823,In_643,In_2372);
xor U824 (N_824,In_1315,In_1504);
nor U825 (N_825,In_375,N_672);
or U826 (N_826,N_564,In_1409);
or U827 (N_827,N_270,In_1715);
nand U828 (N_828,In_604,In_1662);
or U829 (N_829,N_747,In_2117);
nand U830 (N_830,N_164,N_609);
xor U831 (N_831,N_572,In_134);
and U832 (N_832,In_84,In_2281);
and U833 (N_833,In_541,N_626);
or U834 (N_834,In_472,In_2007);
and U835 (N_835,N_516,In_1219);
xnor U836 (N_836,In_2462,In_1698);
xnor U837 (N_837,In_1011,N_513);
nor U838 (N_838,In_2239,N_279);
and U839 (N_839,N_555,N_715);
xnor U840 (N_840,In_1115,In_806);
nand U841 (N_841,In_118,N_27);
or U842 (N_842,In_290,In_2429);
nand U843 (N_843,N_280,In_1297);
nor U844 (N_844,N_742,N_169);
nor U845 (N_845,N_21,In_2384);
xnor U846 (N_846,In_753,N_101);
xor U847 (N_847,In_959,In_1118);
and U848 (N_848,N_574,In_169);
and U849 (N_849,In_2313,In_925);
and U850 (N_850,N_351,N_744);
nor U851 (N_851,In_2127,In_137);
nand U852 (N_852,N_567,N_566);
xor U853 (N_853,In_2269,In_110);
and U854 (N_854,In_2460,In_761);
and U855 (N_855,In_1234,In_1575);
xor U856 (N_856,N_378,In_1888);
or U857 (N_857,N_606,In_332);
nand U858 (N_858,In_1296,In_1818);
nor U859 (N_859,In_219,In_867);
nand U860 (N_860,In_315,In_1536);
or U861 (N_861,N_446,In_199);
nand U862 (N_862,N_102,N_547);
nor U863 (N_863,In_343,In_700);
xor U864 (N_864,N_52,N_434);
or U865 (N_865,N_497,In_1193);
and U866 (N_866,N_72,In_1338);
and U867 (N_867,N_229,N_304);
and U868 (N_868,N_46,N_631);
or U869 (N_869,In_1111,N_134);
nor U870 (N_870,In_1462,In_1716);
nand U871 (N_871,N_158,In_880);
and U872 (N_872,N_87,In_2347);
xor U873 (N_873,In_2364,N_628);
and U874 (N_874,N_324,N_177);
or U875 (N_875,In_2055,N_6);
nor U876 (N_876,In_996,In_141);
or U877 (N_877,N_669,N_142);
or U878 (N_878,In_355,In_1953);
and U879 (N_879,In_388,N_590);
or U880 (N_880,In_1267,N_595);
xor U881 (N_881,In_1160,N_2);
nor U882 (N_882,N_607,In_1763);
and U883 (N_883,In_1336,N_548);
or U884 (N_884,In_97,N_599);
nand U885 (N_885,In_1617,N_61);
or U886 (N_886,N_400,In_467);
or U887 (N_887,In_632,N_573);
nor U888 (N_888,N_299,In_1440);
xor U889 (N_889,N_271,In_64);
or U890 (N_890,N_321,In_350);
nor U891 (N_891,In_1647,N_333);
xnor U892 (N_892,N_326,In_1615);
nor U893 (N_893,In_2318,In_7);
xor U894 (N_894,In_345,N_491);
and U895 (N_895,N_160,N_412);
nand U896 (N_896,In_1387,N_302);
nand U897 (N_897,N_86,In_681);
nor U898 (N_898,In_2216,N_565);
nand U899 (N_899,N_602,In_20);
and U900 (N_900,N_556,In_2078);
xnor U901 (N_901,N_730,N_504);
xnor U902 (N_902,In_1375,In_1444);
xnor U903 (N_903,In_976,N_286);
and U904 (N_904,N_736,N_549);
nand U905 (N_905,In_1875,In_678);
nor U906 (N_906,In_1663,In_1855);
nor U907 (N_907,In_31,N_474);
nand U908 (N_908,In_1744,In_1877);
nor U909 (N_909,In_1385,N_233);
and U910 (N_910,In_1527,In_2363);
nor U911 (N_911,In_2005,In_1826);
xnor U912 (N_912,N_582,In_961);
nor U913 (N_913,In_1704,N_346);
and U914 (N_914,N_343,N_199);
nand U915 (N_915,N_290,N_350);
and U916 (N_916,N_615,N_706);
xnor U917 (N_917,N_676,In_517);
nand U918 (N_918,N_727,In_933);
and U919 (N_919,In_1416,In_152);
nand U920 (N_920,N_424,N_329);
xnor U921 (N_921,In_108,In_2087);
nand U922 (N_922,In_2248,In_2277);
xnor U923 (N_923,N_634,In_853);
xnor U924 (N_924,N_148,In_1031);
nand U925 (N_925,In_874,In_1464);
or U926 (N_926,In_2015,In_1691);
and U927 (N_927,In_425,In_1426);
nand U928 (N_928,In_1653,N_436);
xnor U929 (N_929,In_385,In_94);
or U930 (N_930,In_69,In_1239);
or U931 (N_931,N_622,In_2398);
xor U932 (N_932,N_645,In_43);
nand U933 (N_933,In_672,In_2202);
xor U934 (N_934,In_206,N_195);
nor U935 (N_935,In_2400,N_174);
nand U936 (N_936,In_2314,In_1404);
or U937 (N_937,In_1261,In_994);
and U938 (N_938,In_2260,In_1136);
xnor U939 (N_939,In_1854,In_1484);
xnor U940 (N_940,N_230,In_1207);
nor U941 (N_941,N_19,In_1358);
or U942 (N_942,N_17,In_2166);
nor U943 (N_943,N_15,N_571);
and U944 (N_944,In_919,N_215);
nor U945 (N_945,In_2439,In_148);
or U946 (N_946,In_295,N_740);
nand U947 (N_947,In_875,In_1518);
xor U948 (N_948,N_478,In_109);
or U949 (N_949,In_2206,In_2022);
nor U950 (N_950,In_488,N_116);
or U951 (N_951,In_2115,N_707);
nand U952 (N_952,In_1714,In_2186);
or U953 (N_953,N_344,N_312);
and U954 (N_954,In_573,In_1628);
or U955 (N_955,In_55,N_598);
or U956 (N_956,N_147,N_456);
xnor U957 (N_957,N_308,N_216);
nor U958 (N_958,N_583,In_1045);
xnor U959 (N_959,In_752,In_626);
nor U960 (N_960,In_737,N_269);
nor U961 (N_961,In_478,In_1505);
nor U962 (N_962,In_1435,In_1083);
xnor U963 (N_963,In_649,In_1985);
or U964 (N_964,In_62,N_376);
xnor U965 (N_965,In_210,In_2103);
nor U966 (N_966,In_755,In_978);
or U967 (N_967,In_1007,In_939);
xor U968 (N_968,In_602,In_1488);
nand U969 (N_969,N_614,In_1980);
or U970 (N_970,In_381,In_1521);
and U971 (N_971,N_212,In_938);
and U972 (N_972,In_1010,In_2408);
and U973 (N_973,N_722,In_788);
nor U974 (N_974,N_732,In_1098);
nor U975 (N_975,In_1457,In_1204);
or U976 (N_976,In_268,N_128);
nor U977 (N_977,In_1984,In_2412);
xnor U978 (N_978,In_1961,In_494);
nand U979 (N_979,N_473,In_562);
nand U980 (N_980,In_1184,In_2150);
xnor U981 (N_981,In_2028,N_745);
and U982 (N_982,N_518,In_458);
and U983 (N_983,In_156,In_1254);
nand U984 (N_984,In_648,In_856);
xnor U985 (N_985,N_630,N_691);
xor U986 (N_986,N_653,In_1232);
nor U987 (N_987,In_844,In_2254);
nor U988 (N_988,N_291,In_776);
nor U989 (N_989,N_240,In_1750);
nand U990 (N_990,In_1863,In_964);
nand U991 (N_991,N_420,In_816);
and U992 (N_992,In_2457,N_3);
and U993 (N_993,N_592,In_21);
and U994 (N_994,N_405,In_1563);
nor U995 (N_995,In_2072,In_1186);
or U996 (N_996,In_1295,In_911);
xnor U997 (N_997,N_619,N_135);
nand U998 (N_998,In_1613,N_146);
xor U999 (N_999,In_1380,In_2071);
or U1000 (N_1000,In_257,N_130);
xnor U1001 (N_1001,N_647,In_2023);
or U1002 (N_1002,In_715,N_810);
nand U1003 (N_1003,In_497,N_125);
or U1004 (N_1004,N_91,N_475);
nor U1005 (N_1005,N_873,N_364);
or U1006 (N_1006,N_409,In_1088);
xor U1007 (N_1007,N_616,In_900);
nand U1008 (N_1008,N_721,N_600);
nor U1009 (N_1009,In_46,In_1673);
or U1010 (N_1010,In_243,N_712);
nor U1011 (N_1011,N_821,N_568);
and U1012 (N_1012,In_348,In_781);
nand U1013 (N_1013,In_2368,In_1883);
nand U1014 (N_1014,N_503,In_1339);
nand U1015 (N_1015,In_532,N_807);
nand U1016 (N_1016,In_1324,In_2373);
and U1017 (N_1017,N_937,N_956);
nand U1018 (N_1018,N_757,N_858);
and U1019 (N_1019,In_1165,N_580);
or U1020 (N_1020,N_505,In_1382);
nand U1021 (N_1021,In_1762,In_1598);
and U1022 (N_1022,In_1886,In_144);
nor U1023 (N_1023,In_2302,In_2473);
nand U1024 (N_1024,In_2108,N_512);
nor U1025 (N_1025,N_793,N_806);
and U1026 (N_1026,N_689,N_528);
or U1027 (N_1027,In_91,N_782);
nor U1028 (N_1028,N_115,In_695);
and U1029 (N_1029,In_2224,In_987);
and U1030 (N_1030,In_2003,N_35);
xor U1031 (N_1031,In_2219,N_430);
nor U1032 (N_1032,In_1287,In_656);
nand U1033 (N_1033,N_92,In_836);
xor U1034 (N_1034,N_239,In_1177);
or U1035 (N_1035,In_88,N_236);
nand U1036 (N_1036,In_1710,In_1310);
nor U1037 (N_1037,N_778,N_823);
nor U1038 (N_1038,N_900,In_496);
nand U1039 (N_1039,In_2375,N_176);
nand U1040 (N_1040,In_941,In_2056);
nor U1041 (N_1041,In_215,N_585);
nor U1042 (N_1042,N_664,In_549);
nand U1043 (N_1043,N_348,In_195);
nand U1044 (N_1044,N_862,In_2112);
and U1045 (N_1045,In_1285,In_442);
nand U1046 (N_1046,In_1651,N_370);
xor U1047 (N_1047,In_392,In_738);
xnor U1048 (N_1048,N_578,N_826);
or U1049 (N_1049,N_210,In_1739);
xor U1050 (N_1050,In_1320,In_1012);
nor U1051 (N_1051,In_778,N_992);
or U1052 (N_1052,N_981,N_74);
and U1053 (N_1053,N_844,N_841);
xor U1054 (N_1054,In_921,In_1376);
and U1055 (N_1055,N_124,N_755);
nor U1056 (N_1056,In_174,N_121);
xnor U1057 (N_1057,N_485,In_231);
nor U1058 (N_1058,In_1099,In_518);
nand U1059 (N_1059,In_942,In_27);
nor U1060 (N_1060,N_515,N_356);
xnor U1061 (N_1061,In_907,In_881);
nand U1062 (N_1062,N_933,In_529);
and U1063 (N_1063,In_1349,In_1700);
xnor U1064 (N_1064,In_1,N_501);
nand U1065 (N_1065,In_1070,In_525);
nor U1066 (N_1066,N_976,N_725);
nand U1067 (N_1067,In_1509,N_686);
or U1068 (N_1068,In_1846,In_1412);
and U1069 (N_1069,In_490,In_242);
nor U1070 (N_1070,In_2399,In_2013);
xor U1071 (N_1071,N_553,N_586);
and U1072 (N_1072,In_665,In_1025);
xnor U1073 (N_1073,N_654,N_784);
xor U1074 (N_1074,In_1140,N_765);
nor U1075 (N_1075,N_659,In_1284);
nand U1076 (N_1076,In_1530,N_918);
xnor U1077 (N_1077,In_2245,In_1910);
or U1078 (N_1078,In_1537,In_54);
xnor U1079 (N_1079,In_1266,In_2440);
and U1080 (N_1080,In_1788,N_34);
xor U1081 (N_1081,In_1335,N_808);
or U1082 (N_1082,In_2031,N_527);
or U1083 (N_1083,In_2437,In_591);
nand U1084 (N_1084,N_931,In_973);
or U1085 (N_1085,In_2486,In_380);
xnor U1086 (N_1086,In_1703,In_326);
xor U1087 (N_1087,In_1194,In_2134);
and U1088 (N_1088,In_898,In_1562);
or U1089 (N_1089,In_2085,In_578);
xnor U1090 (N_1090,N_817,N_445);
xnor U1091 (N_1091,N_309,In_1832);
xnor U1092 (N_1092,In_1842,N_452);
nand U1093 (N_1093,In_2000,In_1035);
nand U1094 (N_1094,In_1535,In_803);
xnor U1095 (N_1095,In_2124,In_552);
nand U1096 (N_1096,N_633,In_743);
nand U1097 (N_1097,N_769,N_738);
xor U1098 (N_1098,N_701,N_314);
nor U1099 (N_1099,In_1422,N_145);
nand U1100 (N_1100,N_795,In_1371);
or U1101 (N_1101,N_947,In_886);
xnor U1102 (N_1102,N_763,In_2167);
or U1103 (N_1103,In_1791,In_1555);
nand U1104 (N_1104,In_1480,In_1236);
xnor U1105 (N_1105,In_38,N_537);
and U1106 (N_1106,N_869,In_1022);
nand U1107 (N_1107,In_1853,N_909);
nor U1108 (N_1108,N_154,N_675);
xnor U1109 (N_1109,N_867,In_718);
xor U1110 (N_1110,In_240,In_1664);
xnor U1111 (N_1111,N_604,In_696);
or U1112 (N_1112,In_1565,N_964);
or U1113 (N_1113,In_300,In_1392);
nand U1114 (N_1114,N_611,In_354);
nor U1115 (N_1115,N_261,N_849);
or U1116 (N_1116,In_2099,N_438);
and U1117 (N_1117,N_929,In_1925);
nor U1118 (N_1118,N_729,N_942);
nor U1119 (N_1119,In_274,N_157);
xor U1120 (N_1120,In_1471,In_2479);
or U1121 (N_1121,In_2496,In_2425);
and U1122 (N_1122,N_794,N_735);
nor U1123 (N_1123,N_612,N_853);
nor U1124 (N_1124,In_2499,In_1533);
or U1125 (N_1125,N_940,In_1608);
nand U1126 (N_1126,In_2261,In_586);
and U1127 (N_1127,N_288,N_584);
and U1128 (N_1128,In_1872,In_1244);
and U1129 (N_1129,In_1069,In_2032);
and U1130 (N_1130,N_666,N_550);
nor U1131 (N_1131,In_1474,N_543);
nor U1132 (N_1132,N_53,N_926);
nand U1133 (N_1133,N_41,In_113);
and U1134 (N_1134,In_1540,In_1352);
nand U1135 (N_1135,In_177,In_2415);
nor U1136 (N_1136,In_2394,In_913);
or U1137 (N_1137,N_293,In_2101);
nor U1138 (N_1138,In_1138,In_1652);
or U1139 (N_1139,In_2477,N_891);
and U1140 (N_1140,In_564,N_786);
xor U1141 (N_1141,N_768,In_1196);
or U1142 (N_1142,N_76,In_224);
nand U1143 (N_1143,In_2231,N_594);
or U1144 (N_1144,N_835,In_1161);
nand U1145 (N_1145,In_1433,In_936);
nor U1146 (N_1146,In_1318,In_2410);
xor U1147 (N_1147,N_913,In_510);
xnor U1148 (N_1148,In_2431,In_120);
nand U1149 (N_1149,N_796,In_79);
nand U1150 (N_1150,N_950,N_804);
or U1151 (N_1151,In_312,N_832);
xor U1152 (N_1152,In_12,In_854);
nand U1153 (N_1153,In_1740,In_2024);
xnor U1154 (N_1154,In_796,N_502);
nand U1155 (N_1155,N_375,In_1482);
xor U1156 (N_1156,In_1289,N_652);
nor U1157 (N_1157,In_861,In_1655);
or U1158 (N_1158,In_1068,N_974);
or U1159 (N_1159,N_524,In_2151);
and U1160 (N_1160,N_517,N_906);
or U1161 (N_1161,In_140,In_1605);
and U1162 (N_1162,N_903,In_328);
nor U1163 (N_1163,In_1092,In_1388);
xnor U1164 (N_1164,In_1000,In_253);
or U1165 (N_1165,In_1799,N_753);
or U1166 (N_1166,In_1288,N_448);
and U1167 (N_1167,N_934,In_501);
nand U1168 (N_1168,N_972,N_899);
or U1169 (N_1169,In_1543,In_1955);
or U1170 (N_1170,N_854,In_1250);
nor U1171 (N_1171,N_791,In_1660);
or U1172 (N_1172,In_128,N_658);
nor U1173 (N_1173,In_2105,In_30);
and U1174 (N_1174,In_1102,In_1924);
nor U1175 (N_1175,In_471,N_294);
and U1176 (N_1176,In_1586,N_476);
xor U1177 (N_1177,In_1659,N_307);
and U1178 (N_1178,In_1597,In_1755);
and U1179 (N_1179,In_1789,In_22);
nor U1180 (N_1180,In_904,N_865);
nor U1181 (N_1181,N_901,N_369);
xnor U1182 (N_1182,N_895,N_562);
xor U1183 (N_1183,N_805,N_510);
xnor U1184 (N_1184,N_649,N_920);
or U1185 (N_1185,In_370,In_800);
nand U1186 (N_1186,In_1838,N_802);
or U1187 (N_1187,N_917,In_991);
nor U1188 (N_1188,N_202,In_1688);
nor U1189 (N_1189,N_519,In_25);
or U1190 (N_1190,In_2064,N_156);
or U1191 (N_1191,N_500,In_1195);
nand U1192 (N_1192,In_1921,N_958);
nand U1193 (N_1193,In_1758,N_110);
nand U1194 (N_1194,N_591,N_946);
nand U1195 (N_1195,In_93,In_338);
nor U1196 (N_1196,N_117,N_908);
xor U1197 (N_1197,N_419,N_385);
nand U1198 (N_1198,N_75,In_96);
or U1199 (N_1199,N_487,N_962);
xnor U1200 (N_1200,In_2044,In_1152);
nand U1201 (N_1201,In_2229,N_105);
nand U1202 (N_1202,In_1638,In_1369);
xor U1203 (N_1203,In_2251,In_1168);
nor U1204 (N_1204,N_813,In_1607);
and U1205 (N_1205,N_635,In_2278);
and U1206 (N_1206,N_682,In_1028);
xnor U1207 (N_1207,In_746,In_1220);
nand U1208 (N_1208,In_674,N_542);
nand U1209 (N_1209,N_818,N_627);
and U1210 (N_1210,In_201,In_2168);
nor U1211 (N_1211,In_2470,N_965);
and U1212 (N_1212,N_575,N_833);
nand U1213 (N_1213,In_426,In_2218);
or U1214 (N_1214,In_1312,In_1251);
and U1215 (N_1215,In_1417,In_1278);
or U1216 (N_1216,In_1650,N_183);
nor U1217 (N_1217,In_2325,N_951);
xor U1218 (N_1218,In_583,N_184);
nor U1219 (N_1219,N_30,In_571);
nand U1220 (N_1220,In_1609,N_687);
xnor U1221 (N_1221,N_916,In_724);
nor U1222 (N_1222,N_207,In_871);
nand U1223 (N_1223,N_948,In_193);
xnor U1224 (N_1224,N_984,In_730);
or U1225 (N_1225,N_714,In_1726);
nor U1226 (N_1226,N_175,N_569);
and U1227 (N_1227,In_705,N_811);
and U1228 (N_1228,N_318,In_2228);
or U1229 (N_1229,In_58,In_1421);
or U1230 (N_1230,In_311,In_1015);
nor U1231 (N_1231,N_871,N_756);
or U1232 (N_1232,In_862,N_68);
or U1233 (N_1233,N_234,In_1852);
nand U1234 (N_1234,N_88,In_1756);
or U1235 (N_1235,N_941,In_550);
xnor U1236 (N_1236,In_1754,In_308);
or U1237 (N_1237,In_292,In_685);
xor U1238 (N_1238,In_1684,In_2131);
nor U1239 (N_1239,In_1032,N_316);
or U1240 (N_1240,N_790,In_76);
xnor U1241 (N_1241,N_363,In_2069);
xnor U1242 (N_1242,In_1553,In_1761);
and U1243 (N_1243,N_529,In_218);
or U1244 (N_1244,In_574,N_935);
and U1245 (N_1245,In_903,In_489);
xor U1246 (N_1246,In_1992,N_927);
or U1247 (N_1247,N_787,N_231);
and U1248 (N_1248,In_1891,In_657);
xor U1249 (N_1249,N_610,In_1425);
nand U1250 (N_1250,In_2463,N_274);
nand U1251 (N_1251,N_1059,N_1080);
xor U1252 (N_1252,N_1089,N_1058);
nand U1253 (N_1253,N_1244,In_1039);
or U1254 (N_1254,N_94,In_703);
nor U1255 (N_1255,N_79,In_2441);
xnor U1256 (N_1256,In_2353,In_1973);
nor U1257 (N_1257,N_1113,N_952);
or U1258 (N_1258,N_1204,N_243);
nor U1259 (N_1259,N_1157,N_1226);
nand U1260 (N_1260,In_1829,In_1902);
nand U1261 (N_1261,N_509,In_456);
xnor U1262 (N_1262,N_25,N_772);
or U1263 (N_1263,N_774,N_172);
nand U1264 (N_1264,N_449,In_1885);
xor U1265 (N_1265,In_2060,N_719);
or U1266 (N_1266,N_986,In_629);
or U1267 (N_1267,N_122,In_659);
nor U1268 (N_1268,In_2427,N_953);
or U1269 (N_1269,In_2299,In_1542);
nand U1270 (N_1270,N_393,In_1892);
xor U1271 (N_1271,In_1097,N_460);
xor U1272 (N_1272,N_944,N_1029);
nand U1273 (N_1273,N_359,In_314);
and U1274 (N_1274,N_777,In_1005);
xnor U1275 (N_1275,In_2386,N_816);
and U1276 (N_1276,In_698,N_496);
xor U1277 (N_1277,N_997,N_1206);
xor U1278 (N_1278,N_1193,N_1225);
or U1279 (N_1279,In_194,In_1485);
xnor U1280 (N_1280,N_67,N_855);
nand U1281 (N_1281,In_1072,N_988);
nor U1282 (N_1282,N_392,N_1117);
and U1283 (N_1283,In_627,In_2180);
xnor U1284 (N_1284,N_1105,N_315);
and U1285 (N_1285,In_2490,In_1037);
and U1286 (N_1286,In_1873,N_311);
and U1287 (N_1287,In_1749,In_92);
nor U1288 (N_1288,N_603,N_1164);
nand U1289 (N_1289,N_1159,In_1626);
nor U1290 (N_1290,In_1556,In_2471);
nor U1291 (N_1291,In_597,In_822);
and U1292 (N_1292,In_1574,N_1088);
nand U1293 (N_1293,N_636,N_648);
nor U1294 (N_1294,N_1071,In_1210);
and U1295 (N_1295,In_1679,In_2283);
nand U1296 (N_1296,N_1019,In_305);
nand U1297 (N_1297,N_828,In_1896);
xnor U1298 (N_1298,In_132,In_2316);
xor U1299 (N_1299,N_705,N_1102);
nand U1300 (N_1300,N_1200,In_1377);
nand U1301 (N_1301,In_873,N_1228);
nand U1302 (N_1302,N_1123,In_1808);
or U1303 (N_1303,N_868,N_877);
nand U1304 (N_1304,N_1153,In_1968);
nand U1305 (N_1305,In_1475,N_874);
nor U1306 (N_1306,In_522,N_970);
nand U1307 (N_1307,N_690,In_834);
nor U1308 (N_1308,N_860,In_2291);
and U1309 (N_1309,N_809,N_1135);
or U1310 (N_1310,In_1283,N_514);
or U1311 (N_1311,N_978,N_1236);
nor U1312 (N_1312,In_2213,In_2097);
nor U1313 (N_1313,In_682,In_799);
xnor U1314 (N_1314,N_1069,N_881);
or U1315 (N_1315,N_303,In_2110);
nor U1316 (N_1316,In_204,In_1988);
nand U1317 (N_1317,N_238,In_1020);
or U1318 (N_1318,N_897,In_2279);
xnor U1319 (N_1319,In_1051,In_1646);
or U1320 (N_1320,N_1018,N_621);
or U1321 (N_1321,N_150,N_552);
nor U1322 (N_1322,N_406,In_1539);
xor U1323 (N_1323,N_1179,In_2155);
nand U1324 (N_1324,N_112,In_823);
nand U1325 (N_1325,In_2282,N_1074);
nor U1326 (N_1326,N_827,N_349);
xnor U1327 (N_1327,N_876,N_665);
nand U1328 (N_1328,In_1728,N_1098);
nor U1329 (N_1329,N_1021,In_1451);
xnor U1330 (N_1330,N_752,N_776);
nor U1331 (N_1331,In_1394,N_1161);
nor U1332 (N_1332,N_698,In_2270);
or U1333 (N_1333,N_1147,N_936);
nand U1334 (N_1334,N_1171,In_225);
nor U1335 (N_1335,N_1062,In_847);
xor U1336 (N_1336,In_1974,N_887);
xor U1337 (N_1337,N_250,N_1091);
nand U1338 (N_1338,In_714,In_901);
xnor U1339 (N_1339,N_1144,N_1217);
xnor U1340 (N_1340,N_928,N_1242);
and U1341 (N_1341,N_541,N_1082);
and U1342 (N_1342,In_1104,In_1401);
xor U1343 (N_1343,N_998,In_839);
nor U1344 (N_1344,In_2089,In_577);
xnor U1345 (N_1345,In_2125,In_372);
or U1346 (N_1346,N_850,N_1106);
and U1347 (N_1347,N_1215,In_1096);
nor U1348 (N_1348,N_581,In_1587);
or U1349 (N_1349,In_196,In_1467);
xor U1350 (N_1350,N_1249,In_768);
nand U1351 (N_1351,N_673,In_325);
or U1352 (N_1352,N_1122,In_80);
nor U1353 (N_1353,N_620,In_664);
nand U1354 (N_1354,N_613,N_677);
xor U1355 (N_1355,N_671,In_2458);
and U1356 (N_1356,N_1086,N_1205);
or U1357 (N_1357,N_1224,In_624);
nand U1358 (N_1358,In_2036,N_748);
nand U1359 (N_1359,N_1227,In_2096);
or U1360 (N_1360,N_641,In_1057);
and U1361 (N_1361,N_1057,N_775);
xor U1362 (N_1362,N_694,In_2365);
xor U1363 (N_1363,In_902,N_90);
xnor U1364 (N_1364,N_863,In_1439);
nand U1365 (N_1365,In_1052,N_1104);
xnor U1366 (N_1366,N_425,N_1051);
or U1367 (N_1367,In_45,In_272);
and U1368 (N_1368,N_241,In_882);
nor U1369 (N_1369,In_2133,N_949);
nor U1370 (N_1370,N_1151,In_2377);
or U1371 (N_1371,N_1008,N_189);
or U1372 (N_1372,In_1956,N_884);
nand U1373 (N_1373,N_390,In_1525);
and U1374 (N_1374,N_367,N_486);
or U1375 (N_1375,N_743,In_280);
xor U1376 (N_1376,N_1190,N_1137);
or U1377 (N_1377,N_650,In_303);
xor U1378 (N_1378,In_57,In_879);
and U1379 (N_1379,N_819,N_388);
nand U1380 (N_1380,N_969,N_939);
xor U1381 (N_1381,N_838,N_864);
xnor U1382 (N_1382,In_1681,N_1050);
nor U1383 (N_1383,In_2274,N_847);
and U1384 (N_1384,In_2195,N_880);
or U1385 (N_1385,N_1110,N_643);
nor U1386 (N_1386,N_882,In_554);
and U1387 (N_1387,N_1044,N_1043);
or U1388 (N_1388,N_379,N_1119);
or U1389 (N_1389,N_95,N_217);
nor U1390 (N_1390,In_1772,N_54);
and U1391 (N_1391,N_642,In_2341);
and U1392 (N_1392,In_655,In_1991);
nand U1393 (N_1393,In_1511,In_1551);
xnor U1394 (N_1394,N_839,N_655);
nand U1395 (N_1395,In_130,In_1090);
or U1396 (N_1396,N_668,N_683);
and U1397 (N_1397,N_589,N_366);
xnor U1398 (N_1398,N_1136,N_837);
nand U1399 (N_1399,In_1499,In_1932);
or U1400 (N_1400,N_441,In_1513);
nand U1401 (N_1401,N_251,In_2249);
nor U1402 (N_1402,In_2298,N_1176);
xor U1403 (N_1403,N_13,N_959);
nand U1404 (N_1404,In_1216,N_1076);
or U1405 (N_1405,In_539,In_2074);
or U1406 (N_1406,In_100,N_975);
and U1407 (N_1407,N_1028,In_1610);
xnor U1408 (N_1408,N_1196,N_1003);
xor U1409 (N_1409,N_803,N_1195);
nand U1410 (N_1410,In_2008,N_1191);
xor U1411 (N_1411,N_1124,In_2390);
and U1412 (N_1412,N_423,N_1031);
xnor U1413 (N_1413,N_846,N_330);
xor U1414 (N_1414,N_1014,In_2401);
nor U1415 (N_1415,N_893,N_203);
xnor U1416 (N_1416,In_2376,N_429);
and U1417 (N_1417,In_2165,In_892);
nor U1418 (N_1418,In_2357,N_617);
xnor U1419 (N_1419,N_912,In_313);
xnor U1420 (N_1420,In_884,In_33);
xor U1421 (N_1421,N_836,In_896);
or U1422 (N_1422,N_963,N_319);
and U1423 (N_1423,N_198,N_663);
xor U1424 (N_1424,In_794,In_2235);
nor U1425 (N_1425,N_1232,In_66);
nor U1426 (N_1426,N_825,In_1341);
nand U1427 (N_1427,N_866,In_2321);
nand U1428 (N_1428,N_1120,In_2149);
xnor U1429 (N_1429,N_490,In_1522);
xnor U1430 (N_1430,N_557,In_1329);
nand U1431 (N_1431,N_1099,N_1075);
nor U1432 (N_1432,In_40,In_1256);
nor U1433 (N_1433,N_1108,N_875);
xnor U1434 (N_1434,In_1776,In_2265);
or U1435 (N_1435,N_798,N_14);
nand U1436 (N_1436,In_667,In_1950);
xnor U1437 (N_1437,In_607,In_751);
or U1438 (N_1438,N_365,In_2392);
or U1439 (N_1439,In_2489,N_1235);
nor U1440 (N_1440,In_1333,N_904);
nand U1441 (N_1441,In_2366,N_731);
nor U1442 (N_1442,In_2385,In_1139);
and U1443 (N_1443,N_355,N_1126);
xor U1444 (N_1444,N_1053,In_1067);
xor U1445 (N_1445,In_1364,In_241);
xor U1446 (N_1446,N_536,In_1913);
xnor U1447 (N_1447,In_1124,In_1951);
nor U1448 (N_1448,In_2221,In_422);
and U1449 (N_1449,In_1408,N_297);
or U1450 (N_1450,N_1245,N_1040);
xnor U1451 (N_1451,In_2413,In_127);
nor U1452 (N_1452,In_843,N_1246);
xor U1453 (N_1453,N_1133,N_1007);
or U1454 (N_1454,N_780,In_452);
and U1455 (N_1455,N_1177,In_1109);
or U1456 (N_1456,N_498,In_329);
nor U1457 (N_1457,N_1035,In_1814);
xor U1458 (N_1458,N_993,In_1274);
xnor U1459 (N_1459,N_1081,N_930);
nor U1460 (N_1460,N_1234,N_994);
nor U1461 (N_1461,In_1520,In_1443);
and U1462 (N_1462,In_339,N_859);
xnor U1463 (N_1463,In_1502,In_850);
or U1464 (N_1464,In_2275,N_878);
nor U1465 (N_1465,In_105,N_1241);
and U1466 (N_1466,N_896,N_1032);
and U1467 (N_1467,In_379,In_42);
or U1468 (N_1468,N_403,In_1748);
xnor U1469 (N_1469,In_971,In_1771);
nand U1470 (N_1470,N_219,N_922);
xnor U1471 (N_1471,N_1239,N_382);
nand U1472 (N_1472,N_9,In_2148);
or U1473 (N_1473,In_2447,In_382);
xnor U1474 (N_1474,N_1011,N_1010);
xnor U1475 (N_1475,N_1223,N_196);
nor U1476 (N_1476,In_1062,In_1731);
nand U1477 (N_1477,In_1893,N_824);
or U1478 (N_1478,N_1026,N_1038);
nand U1479 (N_1479,N_1013,In_955);
or U1480 (N_1480,In_182,In_2391);
or U1481 (N_1481,In_89,N_432);
nand U1482 (N_1482,In_945,N_1233);
xnor U1483 (N_1483,N_1212,N_443);
xor U1484 (N_1484,N_834,N_945);
nor U1485 (N_1485,In_2342,N_1129);
nand U1486 (N_1486,N_1181,In_2360);
or U1487 (N_1487,In_434,In_777);
and U1488 (N_1488,N_1143,In_630);
nor U1489 (N_1489,N_480,N_1248);
xnor U1490 (N_1490,N_494,N_1178);
xnor U1491 (N_1491,In_3,N_1203);
and U1492 (N_1492,N_954,N_1237);
or U1493 (N_1493,In_1397,N_1103);
and U1494 (N_1494,In_2119,In_1350);
xor U1495 (N_1495,N_1107,In_1722);
nand U1496 (N_1496,In_1592,In_1064);
nand U1497 (N_1497,N_1023,N_484);
nor U1498 (N_1498,In_848,N_711);
or U1499 (N_1499,N_1015,N_1045);
and U1500 (N_1500,N_410,N_187);
and U1501 (N_1501,In_2312,N_454);
nor U1502 (N_1502,N_1022,In_1790);
xor U1503 (N_1503,N_639,In_774);
nor U1504 (N_1504,N_771,N_1398);
nor U1505 (N_1505,In_1043,In_1410);
or U1506 (N_1506,N_535,N_1002);
or U1507 (N_1507,N_1275,In_2129);
nand U1508 (N_1508,N_1027,N_1453);
or U1509 (N_1509,N_1309,In_1157);
or U1510 (N_1510,N_526,In_1524);
or U1511 (N_1511,N_1175,N_1396);
nand U1512 (N_1512,N_644,N_1459);
xor U1513 (N_1513,In_2387,N_1168);
nor U1514 (N_1514,N_1261,N_1240);
or U1515 (N_1515,N_1378,In_832);
nand U1516 (N_1516,In_2041,In_498);
or U1517 (N_1517,N_1406,N_1194);
nand U1518 (N_1518,N_1455,N_1183);
xnor U1519 (N_1519,N_1490,In_1904);
or U1520 (N_1520,In_477,In_1939);
or U1521 (N_1521,N_214,N_428);
xnor U1522 (N_1522,N_815,In_1268);
and U1523 (N_1523,N_1121,In_2076);
xnor U1524 (N_1524,N_987,N_1348);
nor U1525 (N_1525,N_1095,N_1302);
and U1526 (N_1526,N_1047,N_1338);
nor U1527 (N_1527,N_1446,N_1295);
or U1528 (N_1528,N_1428,In_2135);
xnor U1529 (N_1529,N_1265,In_582);
or U1530 (N_1530,N_453,In_1171);
nand U1531 (N_1531,N_558,N_401);
and U1532 (N_1532,In_1760,N_1413);
and U1533 (N_1533,N_1250,N_342);
and U1534 (N_1534,In_261,In_2442);
nand U1535 (N_1535,N_1219,N_1304);
nor U1536 (N_1536,N_1410,N_1314);
xor U1537 (N_1537,In_780,N_1380);
and U1538 (N_1538,In_1309,N_1473);
or U1539 (N_1539,N_310,N_1426);
nor U1540 (N_1540,In_1313,N_1201);
nand U1541 (N_1541,N_521,In_1199);
and U1542 (N_1542,In_1631,In_713);
or U1543 (N_1543,In_726,In_1701);
xnor U1544 (N_1544,In_1983,In_1880);
or U1545 (N_1545,In_651,N_1485);
xnor U1546 (N_1546,N_1373,N_1369);
or U1547 (N_1547,N_1155,In_720);
and U1548 (N_1548,N_520,In_2009);
nand U1549 (N_1549,N_408,In_161);
xor U1550 (N_1550,N_56,N_1333);
nand U1551 (N_1551,In_1018,N_1247);
xnor U1552 (N_1552,N_1462,In_1454);
nand U1553 (N_1553,In_1512,N_466);
or U1554 (N_1554,In_476,N_1041);
or U1555 (N_1555,N_1327,In_924);
nor U1556 (N_1556,N_872,N_1127);
nor U1557 (N_1557,N_1128,In_500);
nor U1558 (N_1558,N_1416,In_1423);
xnor U1559 (N_1559,In_2362,N_1495);
nand U1560 (N_1560,N_1141,N_894);
nor U1561 (N_1561,In_2077,N_1184);
or U1562 (N_1562,N_227,In_1357);
or U1563 (N_1563,N_1229,N_63);
and U1564 (N_1564,In_910,In_502);
xor U1565 (N_1565,N_1278,N_1263);
nand U1566 (N_1566,In_149,N_923);
nand U1567 (N_1567,In_450,N_1405);
xor U1568 (N_1568,N_29,N_163);
or U1569 (N_1569,N_1262,In_1473);
xnor U1570 (N_1570,In_1355,N_1192);
and U1571 (N_1571,In_1849,N_703);
nand U1572 (N_1572,N_932,N_1366);
and U1573 (N_1573,In_19,N_57);
or U1574 (N_1574,In_807,In_2223);
or U1575 (N_1575,In_2051,In_281);
and U1576 (N_1576,In_2142,In_1561);
xor U1577 (N_1577,In_237,N_1006);
xnor U1578 (N_1578,N_257,In_2137);
nand U1579 (N_1579,In_337,N_656);
xnor U1580 (N_1580,N_545,N_1440);
xnor U1581 (N_1581,In_251,N_1387);
or U1582 (N_1582,In_1866,N_1149);
nand U1583 (N_1583,N_1491,N_507);
and U1584 (N_1584,In_828,N_417);
and U1585 (N_1585,In_322,N_1470);
xnor U1586 (N_1586,N_298,N_106);
nand U1587 (N_1587,In_1279,N_477);
xor U1588 (N_1588,In_2035,N_1042);
or U1589 (N_1589,N_618,N_1434);
nand U1590 (N_1590,N_338,In_1827);
nor U1591 (N_1591,N_749,N_1303);
and U1592 (N_1592,N_814,N_1052);
xor U1593 (N_1593,N_1484,N_1496);
or U1594 (N_1594,In_1751,In_748);
xnor U1595 (N_1595,N_1368,N_1005);
nand U1596 (N_1596,In_1036,In_595);
and U1597 (N_1597,In_2414,N_1342);
and U1598 (N_1598,In_784,In_948);
nor U1599 (N_1599,N_1436,N_1297);
and U1600 (N_1600,N_1097,In_1441);
nand U1601 (N_1601,N_851,In_1786);
or U1602 (N_1602,In_1601,In_1792);
and U1603 (N_1603,N_306,In_1783);
nand U1604 (N_1604,In_187,In_35);
nand U1605 (N_1605,N_444,In_765);
xnor U1606 (N_1606,N_1180,In_1869);
and U1607 (N_1607,In_190,In_1718);
and U1608 (N_1608,N_1442,In_572);
nand U1609 (N_1609,In_1682,N_1474);
xor U1610 (N_1610,In_1709,N_1188);
nor U1611 (N_1611,In_855,N_421);
nand U1612 (N_1612,N_1376,In_1810);
xnor U1613 (N_1613,In_2177,N_1158);
nand U1614 (N_1614,In_993,N_1087);
nor U1615 (N_1615,N_1307,N_459);
and U1616 (N_1616,In_342,N_222);
and U1617 (N_1617,N_327,N_910);
nor U1618 (N_1618,In_2405,N_1025);
or U1619 (N_1619,N_1390,N_1340);
and U1620 (N_1620,N_1377,N_1475);
xnor U1621 (N_1621,N_1372,N_1383);
and U1622 (N_1622,In_813,N_451);
nor U1623 (N_1623,In_2280,In_302);
nor U1624 (N_1624,N_1170,In_1862);
xor U1625 (N_1625,N_1169,In_307);
nand U1626 (N_1626,N_921,N_830);
and U1627 (N_1627,N_1477,N_842);
nand U1628 (N_1628,In_1438,In_2428);
or U1629 (N_1629,N_576,In_1629);
xnor U1630 (N_1630,In_1311,In_530);
nor U1631 (N_1631,N_383,N_1429);
nor U1632 (N_1632,N_1187,In_2217);
nand U1633 (N_1633,In_296,N_554);
xnor U1634 (N_1634,N_534,N_1068);
xor U1635 (N_1635,N_1039,In_922);
and U1636 (N_1636,In_1670,In_1770);
and U1637 (N_1637,N_1357,N_493);
nor U1638 (N_1638,N_733,N_254);
and U1639 (N_1639,In_1824,In_2498);
and U1640 (N_1640,N_840,In_457);
nor U1641 (N_1641,In_540,N_42);
xnor U1642 (N_1642,N_1370,In_1192);
xnor U1643 (N_1643,N_1465,N_991);
nand U1644 (N_1644,N_1070,N_275);
xor U1645 (N_1645,N_1111,N_1489);
or U1646 (N_1646,In_680,N_1300);
nand U1647 (N_1647,In_48,N_1100);
or U1648 (N_1648,N_532,N_1315);
nor U1649 (N_1649,N_781,N_1415);
and U1650 (N_1650,In_23,N_961);
and U1651 (N_1651,In_1024,N_0);
or U1652 (N_1652,N_1347,N_1146);
and U1653 (N_1653,N_1270,N_1063);
nor U1654 (N_1654,N_1167,N_1360);
nand U1655 (N_1655,In_1811,N_1324);
nand U1656 (N_1656,N_966,In_1949);
nor U1657 (N_1657,N_1037,N_255);
xnor U1658 (N_1658,N_925,N_483);
nand U1659 (N_1659,N_1065,N_1310);
nand U1660 (N_1660,N_1284,N_1024);
and U1661 (N_1661,N_1173,In_956);
or U1662 (N_1662,N_919,In_1008);
and U1663 (N_1663,N_1389,In_24);
and U1664 (N_1664,N_1397,N_1049);
nor U1665 (N_1665,N_1480,N_1101);
or U1666 (N_1666,In_1252,N_678);
and U1667 (N_1667,In_1060,N_1375);
nand U1668 (N_1668,In_556,N_137);
nand U1669 (N_1669,N_856,N_1054);
nand U1670 (N_1670,N_1145,N_938);
xnor U1671 (N_1671,N_1404,N_1441);
xor U1672 (N_1672,N_1139,In_1843);
and U1673 (N_1673,In_2246,N_1209);
and U1674 (N_1674,N_1391,N_1273);
nand U1675 (N_1675,N_783,N_898);
nand U1676 (N_1676,N_211,N_1116);
nor U1677 (N_1677,N_458,N_1331);
and U1678 (N_1678,N_1482,N_481);
and U1679 (N_1679,In_1328,N_646);
nor U1680 (N_1680,In_402,N_1437);
and U1681 (N_1681,N_328,N_1140);
and U1682 (N_1682,In_2339,N_1494);
nor U1683 (N_1683,N_1418,In_523);
or U1684 (N_1684,In_787,N_587);
nor U1685 (N_1685,N_1386,In_1918);
xor U1686 (N_1686,N_1379,In_1034);
nand U1687 (N_1687,N_1222,N_1345);
nor U1688 (N_1688,N_1162,In_367);
xor U1689 (N_1689,N_97,N_450);
nand U1690 (N_1690,In_1269,In_228);
xor U1691 (N_1691,N_181,N_1276);
nor U1692 (N_1692,N_561,N_1457);
nor U1693 (N_1693,N_797,N_495);
nor U1694 (N_1694,N_1142,N_1432);
nor U1695 (N_1695,N_1401,In_2378);
nor U1696 (N_1696,N_1337,In_2222);
nand U1697 (N_1697,N_1207,N_1419);
or U1698 (N_1698,N_973,In_2);
nor U1699 (N_1699,N_1084,N_1362);
xnor U1700 (N_1700,In_364,In_1100);
or U1701 (N_1701,N_999,In_2464);
nand U1702 (N_1702,N_996,In_2259);
nor U1703 (N_1703,In_2160,N_843);
or U1704 (N_1704,N_1264,In_1632);
nand U1705 (N_1705,N_680,In_2211);
nor U1706 (N_1706,N_1096,In_729);
or U1707 (N_1707,In_2163,N_332);
and U1708 (N_1708,N_1443,N_1308);
xor U1709 (N_1709,In_2010,In_845);
nor U1710 (N_1710,N_40,N_1486);
nor U1711 (N_1711,N_1444,N_1363);
xnor U1712 (N_1712,N_1271,N_1385);
or U1713 (N_1713,N_1399,N_1323);
or U1714 (N_1714,N_983,In_1077);
xor U1715 (N_1715,In_1897,N_601);
nand U1716 (N_1716,In_771,In_1876);
nor U1717 (N_1717,N_1061,N_461);
nand U1718 (N_1718,In_508,N_1427);
and U1719 (N_1719,N_1286,N_1451);
nor U1720 (N_1720,N_1318,N_563);
nor U1721 (N_1721,N_58,N_1055);
xor U1722 (N_1722,N_985,N_822);
and U1723 (N_1723,N_979,N_45);
nand U1724 (N_1724,N_1417,N_1483);
nand U1725 (N_1725,N_726,In_722);
and U1726 (N_1726,N_657,N_1352);
nor U1727 (N_1727,N_253,N_596);
and U1728 (N_1728,N_977,In_2045);
xnor U1729 (N_1729,In_1128,N_36);
nor U1730 (N_1730,In_930,N_1293);
and U1731 (N_1731,N_723,N_1424);
xnor U1732 (N_1732,N_773,In_967);
xnor U1733 (N_1733,N_1210,In_1144);
or U1734 (N_1734,N_1468,N_159);
xor U1735 (N_1735,N_960,N_59);
nand U1736 (N_1736,N_792,In_1221);
nand U1737 (N_1737,N_762,In_809);
or U1738 (N_1738,N_1364,In_2419);
nand U1739 (N_1739,In_443,N_1138);
nor U1740 (N_1740,N_1257,N_1487);
nand U1741 (N_1741,N_1322,N_1090);
nor U1742 (N_1742,N_539,N_1384);
xor U1743 (N_1743,N_1132,N_469);
nor U1744 (N_1744,N_1020,In_336);
and U1745 (N_1745,N_1447,In_829);
and U1746 (N_1746,N_1312,N_943);
nor U1747 (N_1747,N_605,N_354);
or U1748 (N_1748,N_1471,N_64);
xnor U1749 (N_1749,N_1492,N_395);
or U1750 (N_1750,In_2370,In_2198);
nor U1751 (N_1751,N_1513,N_1677);
and U1752 (N_1752,In_1627,In_1383);
or U1753 (N_1753,In_2184,N_1439);
nand U1754 (N_1754,In_2422,N_1328);
and U1755 (N_1755,N_1725,N_1703);
nand U1756 (N_1756,In_2482,N_1326);
xor U1757 (N_1757,In_441,N_1534);
xnor U1758 (N_1758,N_1606,N_1651);
nor U1759 (N_1759,N_1431,N_1706);
or U1760 (N_1760,In_357,N_758);
nand U1761 (N_1761,N_559,N_1652);
and U1762 (N_1762,N_982,N_467);
xor U1763 (N_1763,N_1605,N_252);
nor U1764 (N_1764,N_1593,N_1610);
and U1765 (N_1765,N_684,N_623);
nor U1766 (N_1766,N_1572,N_788);
nand U1767 (N_1767,N_1532,In_1860);
nor U1768 (N_1768,N_1679,N_1678);
xnor U1769 (N_1769,N_1564,N_1559);
or U1770 (N_1770,N_1628,N_1291);
nor U1771 (N_1771,N_870,N_709);
and U1772 (N_1772,N_457,N_1672);
nand U1773 (N_1773,N_1092,N_386);
xor U1774 (N_1774,N_1717,N_1422);
nand U1775 (N_1775,In_710,In_1129);
xor U1776 (N_1776,N_1734,In_1675);
or U1777 (N_1777,N_1518,N_1695);
nand U1778 (N_1778,N_1356,In_1127);
or U1779 (N_1779,N_1464,N_1512);
xnor U1780 (N_1780,N_1596,N_1715);
nor U1781 (N_1781,N_989,N_1085);
nor U1782 (N_1782,N_1619,In_1125);
nand U1783 (N_1783,In_1584,N_760);
or U1784 (N_1784,N_1629,N_1115);
and U1785 (N_1785,N_1269,N_1198);
or U1786 (N_1786,In_1343,N_1301);
xor U1787 (N_1787,N_263,N_1305);
nor U1788 (N_1788,N_1287,N_1573);
and U1789 (N_1789,In_431,N_1346);
or U1790 (N_1790,N_767,N_1319);
or U1791 (N_1791,N_1587,N_1668);
xnor U1792 (N_1792,N_1230,In_2242);
nor U1793 (N_1793,N_1118,N_1067);
nand U1794 (N_1794,N_1561,N_1266);
xnor U1795 (N_1795,N_1634,N_1714);
xnor U1796 (N_1796,N_799,N_1435);
or U1797 (N_1797,N_360,N_1726);
xnor U1798 (N_1798,N_1639,In_548);
nand U1799 (N_1799,N_1742,N_1077);
nand U1800 (N_1800,In_1890,N_1732);
nor U1801 (N_1801,N_857,In_2046);
or U1802 (N_1802,N_1430,N_1371);
nand U1803 (N_1803,N_971,N_1000);
xnor U1804 (N_1804,In_585,N_1612);
and U1805 (N_1805,N_1691,N_1637);
nand U1806 (N_1806,N_718,N_995);
or U1807 (N_1807,In_1452,In_1085);
and U1808 (N_1808,N_540,In_2356);
xnor U1809 (N_1809,N_915,N_892);
xor U1810 (N_1810,In_2271,N_1553);
nand U1811 (N_1811,N_1538,N_1216);
nor U1812 (N_1812,N_699,N_1339);
or U1813 (N_1813,N_902,N_1577);
xor U1814 (N_1814,N_1306,In_1093);
nand U1815 (N_1815,N_879,In_858);
or U1816 (N_1816,N_905,N_296);
and U1817 (N_1817,N_334,N_1199);
nand U1818 (N_1818,N_751,In_189);
xor U1819 (N_1819,N_1298,N_1558);
and U1820 (N_1820,N_1289,N_1609);
xnor U1821 (N_1821,N_389,N_1526);
or U1822 (N_1822,N_597,N_624);
or U1823 (N_1823,N_1591,N_1670);
xor U1824 (N_1824,N_1671,N_911);
and U1825 (N_1825,N_1282,N_1571);
or U1826 (N_1826,N_852,N_1601);
xor U1827 (N_1827,N_889,N_741);
nand U1828 (N_1828,N_831,N_136);
nand U1829 (N_1829,N_1630,N_287);
xnor U1830 (N_1830,N_1114,In_1719);
and U1831 (N_1831,N_1584,N_1461);
or U1832 (N_1832,In_1795,N_1560);
nand U1833 (N_1833,N_1653,N_1663);
nor U1834 (N_1834,N_1531,N_1580);
xnor U1835 (N_1835,In_2383,N_1197);
and U1836 (N_1836,N_1274,In_1546);
and U1837 (N_1837,N_1697,N_522);
nor U1838 (N_1838,N_750,N_1072);
xor U1839 (N_1839,N_1638,N_1001);
and U1840 (N_1840,N_1361,N_1353);
or U1841 (N_1841,N_1625,N_1516);
nor U1842 (N_1842,N_1673,N_1438);
and U1843 (N_1843,N_1646,N_1355);
nand U1844 (N_1844,N_411,In_17);
xor U1845 (N_1845,In_413,N_1567);
xor U1846 (N_1846,N_1615,N_1208);
or U1847 (N_1847,In_351,In_617);
or U1848 (N_1848,In_1734,N_1592);
nor U1849 (N_1849,N_1623,N_1720);
xor U1850 (N_1850,N_688,N_1220);
and U1851 (N_1851,N_766,In_2086);
or U1852 (N_1852,N_1174,N_1066);
nor U1853 (N_1853,N_820,N_1566);
or U1854 (N_1854,N_1613,N_1258);
xor U1855 (N_1855,N_1565,N_1519);
xor U1856 (N_1856,In_1658,N_1256);
nor U1857 (N_1857,N_1288,N_1211);
xor U1858 (N_1858,In_673,In_543);
and U1859 (N_1859,N_812,N_372);
xor U1860 (N_1860,N_1662,In_1243);
nand U1861 (N_1861,N_1009,In_2338);
xnor U1862 (N_1862,N_126,N_801);
and U1863 (N_1863,N_883,N_1414);
nand U1864 (N_1864,In_297,In_684);
or U1865 (N_1865,N_1739,N_317);
or U1866 (N_1866,N_577,N_1400);
or U1867 (N_1867,N_1616,N_1506);
and U1868 (N_1868,N_1724,N_1449);
or U1869 (N_1869,N_779,N_1705);
xor U1870 (N_1870,In_165,N_1680);
nand U1871 (N_1871,N_1525,N_1719);
nand U1872 (N_1872,N_1669,N_1150);
nor U1873 (N_1873,N_1746,N_1551);
nand U1874 (N_1874,N_1165,In_13);
xor U1875 (N_1875,N_1277,N_1109);
or U1876 (N_1876,In_558,In_2301);
nand U1877 (N_1877,N_1574,N_1656);
nor U1878 (N_1878,N_248,N_1598);
xor U1879 (N_1879,N_1701,N_588);
nand U1880 (N_1880,In_1114,N_1589);
or U1881 (N_1881,N_1454,In_2345);
or U1882 (N_1882,In_1969,In_1302);
or U1883 (N_1883,N_1641,N_4);
nand U1884 (N_1884,N_1621,N_218);
xnor U1885 (N_1885,In_1901,N_1479);
and U1886 (N_1886,N_1493,N_1412);
nor U1887 (N_1887,N_1349,N_1648);
xnor U1888 (N_1888,N_1694,N_1500);
and U1889 (N_1889,N_506,N_770);
or U1890 (N_1890,N_1334,N_1093);
xnor U1891 (N_1891,N_1620,In_424);
nand U1892 (N_1892,N_1030,N_1214);
xnor U1893 (N_1893,N_1469,N_1599);
or U1894 (N_1894,N_427,In_1491);
and U1895 (N_1895,N_1730,N_924);
xor U1896 (N_1896,N_1524,N_144);
nand U1897 (N_1897,In_28,N_1570);
or U1898 (N_1898,N_1700,N_1299);
xor U1899 (N_1899,N_221,N_1320);
or U1900 (N_1900,N_1537,N_1655);
or U1901 (N_1901,N_1657,N_1556);
nand U1902 (N_1902,N_1460,N_1336);
nor U1903 (N_1903,N_1685,N_1218);
nor U1904 (N_1904,In_950,N_1520);
nor U1905 (N_1905,N_1604,N_1330);
nor U1906 (N_1906,N_789,N_1733);
xor U1907 (N_1907,N_761,N_1568);
nand U1908 (N_1908,N_1721,N_848);
or U1909 (N_1909,N_1499,N_1702);
xor U1910 (N_1910,N_538,N_1543);
nand U1911 (N_1911,In_418,N_168);
and U1912 (N_1912,N_693,N_1476);
and U1913 (N_1913,N_1505,In_820);
nand U1914 (N_1914,N_1450,N_1736);
nor U1915 (N_1915,In_644,N_1131);
nor U1916 (N_1916,N_1394,N_1544);
or U1917 (N_1917,In_642,N_384);
nor U1918 (N_1918,N_1707,In_2200);
and U1919 (N_1919,In_764,N_1329);
nand U1920 (N_1920,N_381,N_1654);
nor U1921 (N_1921,In_555,N_109);
nor U1922 (N_1922,N_1148,N_1272);
and U1923 (N_1923,N_1213,N_1632);
and U1924 (N_1924,N_1664,N_674);
xnor U1925 (N_1925,N_1403,N_1501);
or U1926 (N_1926,In_352,N_1729);
xnor U1927 (N_1927,In_2444,N_1521);
nand U1928 (N_1928,N_1642,N_1614);
nor U1929 (N_1929,N_632,N_1533);
and U1930 (N_1930,N_759,In_106);
nand U1931 (N_1931,In_250,N_1421);
nand U1932 (N_1932,In_1831,In_2144);
and U1933 (N_1933,N_1527,In_831);
and U1934 (N_1934,In_2292,N_1351);
or U1935 (N_1935,N_1231,In_2192);
nand U1936 (N_1936,In_2436,N_1557);
or U1937 (N_1937,N_1711,N_1420);
nor U1938 (N_1938,N_1073,N_914);
xor U1939 (N_1939,N_1738,In_793);
nor U1940 (N_1940,N_1575,In_1179);
and U1941 (N_1941,N_1684,In_2102);
nor U1942 (N_1942,N_1238,N_1665);
nand U1943 (N_1943,N_1341,N_1292);
nand U1944 (N_1944,N_785,N_1036);
xor U1945 (N_1945,N_1325,N_1251);
nor U1946 (N_1946,N_1466,N_531);
nand U1947 (N_1947,N_754,N_1504);
xor U1948 (N_1948,In_361,N_1687);
xnor U1949 (N_1949,In_10,In_1861);
xor U1950 (N_1950,N_1709,N_955);
nand U1951 (N_1951,N_980,In_1459);
nand U1952 (N_1952,In_1696,In_1319);
nand U1953 (N_1953,N_640,In_943);
or U1954 (N_1954,N_1467,N_608);
or U1955 (N_1955,N_1134,In_666);
or U1956 (N_1956,N_1698,N_1636);
nor U1957 (N_1957,N_1358,N_1727);
xnor U1958 (N_1958,N_1034,N_1658);
xnor U1959 (N_1959,N_1381,In_2255);
and U1960 (N_1960,N_1594,N_1458);
xnor U1961 (N_1961,N_1686,In_1046);
nor U1962 (N_1962,N_1125,N_1317);
xor U1963 (N_1963,In_1917,N_1529);
xor U1964 (N_1964,N_1578,In_63);
or U1965 (N_1965,N_1409,N_1644);
or U1966 (N_1966,N_845,In_2070);
nand U1967 (N_1967,N_1624,N_1448);
nor U1968 (N_1968,N_661,N_1488);
xor U1969 (N_1969,In_1167,N_276);
and U1970 (N_1970,In_1738,N_967);
or U1971 (N_1971,N_1692,In_1370);
xnor U1972 (N_1972,N_1423,In_2452);
and U1973 (N_1973,N_1618,In_2130);
nand U1974 (N_1974,N_1185,In_1492);
nor U1975 (N_1975,N_1745,N_1350);
nor U1976 (N_1976,N_1740,N_1731);
nand U1977 (N_1977,N_1713,In_2191);
nor U1978 (N_1978,N_990,N_1595);
xnor U1979 (N_1979,N_1530,N_907);
and U1980 (N_1980,N_1452,N_397);
or U1981 (N_1981,N_1535,N_1411);
nor U1982 (N_1982,N_1374,N_1017);
and U1983 (N_1983,N_1704,N_1741);
xnor U1984 (N_1984,N_1743,N_1546);
or U1985 (N_1985,N_1622,N_1064);
and U1986 (N_1986,N_1267,N_1283);
nor U1987 (N_1987,In_2446,In_989);
nor U1988 (N_1988,N_1254,N_625);
or U1989 (N_1989,N_1688,N_1569);
xnor U1990 (N_1990,N_1255,In_1642);
xnor U1991 (N_1991,N_1536,N_1748);
xor U1992 (N_1992,N_1737,N_1555);
nand U1993 (N_1993,In_609,N_1033);
nor U1994 (N_1994,N_1456,In_531);
and U1995 (N_1995,N_1712,N_1243);
nand U1996 (N_1996,N_1549,N_1600);
and U1997 (N_1997,N_530,In_2258);
xor U1998 (N_1998,N_337,N_1649);
nand U1999 (N_1999,N_1675,N_1563);
nor U2000 (N_2000,N_1895,N_1723);
nand U2001 (N_2001,N_1786,In_1819);
nor U2002 (N_2002,N_957,N_1834);
nor U2003 (N_2003,N_1995,N_1757);
xor U2004 (N_2004,N_1617,N_1582);
xor U2005 (N_2005,N_1862,N_1689);
nor U2006 (N_2006,N_1880,N_1994);
nor U2007 (N_2007,N_1899,N_720);
xor U2008 (N_2008,N_1972,N_1252);
and U2009 (N_2009,In_1523,N_1777);
nor U2010 (N_2010,N_1873,N_1902);
and U2011 (N_2011,N_1964,N_1784);
xor U2012 (N_2012,N_1588,N_1968);
or U2013 (N_2013,N_1918,N_1809);
nor U2014 (N_2014,N_1947,N_1048);
xnor U2015 (N_2015,N_1844,N_1750);
and U2016 (N_2016,N_1976,N_1957);
xor U2017 (N_2017,N_1645,N_1763);
nand U2018 (N_2018,N_525,In_479);
xor U2019 (N_2019,N_1650,N_1152);
xnor U2020 (N_2020,N_43,N_670);
nand U2021 (N_2021,In_1940,N_1907);
nand U2022 (N_2022,N_155,In_2025);
xor U2023 (N_2023,N_1785,N_1382);
xor U2024 (N_2024,N_1961,N_1926);
nand U2025 (N_2025,N_1798,N_1911);
nor U2026 (N_2026,N_1764,N_1833);
nor U2027 (N_2027,N_1989,N_1765);
nor U2028 (N_2028,N_1843,In_2468);
and U2029 (N_2029,N_1912,N_1888);
or U2030 (N_2030,N_1906,N_1502);
xnor U2031 (N_2031,N_1640,N_1796);
nor U2032 (N_2032,N_1294,N_1835);
and U2033 (N_2033,N_1975,N_127);
xnor U2034 (N_2034,N_1548,N_1869);
and U2035 (N_2035,N_1881,N_829);
xnor U2036 (N_2036,N_1296,N_1761);
xor U2037 (N_2037,N_716,N_1160);
nand U2038 (N_2038,N_1774,N_1202);
nand U2039 (N_2039,In_519,N_1056);
and U2040 (N_2040,N_1808,N_1507);
nor U2041 (N_2041,N_1759,N_1872);
xnor U2042 (N_2042,N_1953,N_1930);
or U2043 (N_2043,N_1253,N_1004);
nor U2044 (N_2044,N_1260,N_1945);
and U2045 (N_2045,In_1648,N_1913);
and U2046 (N_2046,N_1767,N_1280);
xnor U2047 (N_2047,In_817,N_1259);
nor U2048 (N_2048,N_1581,N_1779);
nor U2049 (N_2049,N_1012,N_1949);
or U2050 (N_2050,In_1431,N_700);
xor U2051 (N_2051,N_1603,N_1890);
nand U2052 (N_2052,N_1631,N_1079);
nand U2053 (N_2053,In_1989,N_1758);
xor U2054 (N_2054,N_1762,N_1946);
xor U2055 (N_2055,N_1916,N_1850);
nor U2056 (N_2056,N_1990,N_1936);
xor U2057 (N_2057,N_1801,N_1407);
xnor U2058 (N_2058,N_1562,N_1497);
nor U2059 (N_2059,N_1884,N_1805);
nand U2060 (N_2060,N_281,N_1928);
nand U2061 (N_2061,N_10,N_1182);
xnor U2062 (N_2062,N_1921,In_2172);
and U2063 (N_2063,N_1510,N_1819);
nand U2064 (N_2064,N_1980,N_1987);
or U2065 (N_2065,N_50,N_1931);
or U2066 (N_2066,In_2309,N_1523);
xnor U2067 (N_2067,In_1078,N_1517);
xnor U2068 (N_2068,In_2317,In_2478);
nor U2069 (N_2069,N_1978,N_1954);
nand U2070 (N_2070,N_1221,N_1772);
and U2071 (N_2071,In_1483,N_1973);
and U2072 (N_2072,N_1959,N_1935);
nor U2073 (N_2073,N_1878,N_1163);
and U2074 (N_2074,N_1579,N_1951);
or U2075 (N_2075,N_1965,N_1778);
nor U2076 (N_2076,N_1923,N_1794);
or U2077 (N_2077,N_1824,N_1856);
xor U2078 (N_2078,N_1539,N_1755);
or U2079 (N_2079,N_1799,N_93);
nor U2080 (N_2080,In_1596,N_885);
or U2081 (N_2081,N_1552,N_1335);
nand U2082 (N_2082,N_1955,In_1180);
and U2083 (N_2083,N_1367,N_99);
nand U2084 (N_2084,N_1332,N_1917);
or U2085 (N_2085,N_1789,N_1863);
nand U2086 (N_2086,N_1979,In_2358);
and U2087 (N_2087,N_1842,N_1866);
or U2088 (N_2088,In_1146,N_1909);
xnor U2089 (N_2089,N_1861,In_1405);
xnor U2090 (N_2090,N_1920,In_1699);
nand U2091 (N_2091,N_1392,N_340);
or U2092 (N_2092,N_1359,N_1666);
and U2093 (N_2093,N_1771,N_1722);
and U2094 (N_2094,N_1826,N_1969);
nor U2095 (N_2095,N_1635,N_710);
or U2096 (N_2096,N_1845,N_1849);
xor U2097 (N_2097,N_1971,N_1611);
nand U2098 (N_2098,N_1633,N_1597);
xnor U2099 (N_2099,N_1905,In_509);
and U2100 (N_2100,N_1815,N_1586);
or U2101 (N_2101,N_1892,N_1886);
xor U2102 (N_2102,N_1887,N_1832);
and U2103 (N_2103,N_1806,N_1402);
nand U2104 (N_2104,N_141,N_1768);
and U2105 (N_2105,N_1365,N_1927);
or U2106 (N_2106,In_1143,N_1667);
nand U2107 (N_2107,N_1682,N_1901);
and U2108 (N_2108,N_651,N_1781);
or U2109 (N_2109,N_1311,N_1780);
and U2110 (N_2110,N_1481,N_1172);
and U2111 (N_2111,N_511,In_1887);
xnor U2112 (N_2112,N_1822,N_1966);
xnor U2113 (N_2113,N_1718,N_1811);
nor U2114 (N_2114,N_1130,N_1983);
or U2115 (N_2115,N_1857,N_764);
and U2116 (N_2116,N_546,N_1770);
xor U2117 (N_2117,N_1851,N_1016);
or U2118 (N_2118,N_1751,In_520);
or U2119 (N_2119,N_1841,N_1313);
xnor U2120 (N_2120,N_1992,In_1727);
and U2121 (N_2121,N_1478,In_2430);
nor U2122 (N_2122,N_861,N_1950);
xor U2123 (N_2123,N_1867,N_1837);
nor U2124 (N_2124,N_1879,N_1773);
or U2125 (N_2125,N_1607,N_1997);
nand U2126 (N_2126,N_1585,N_1699);
nand U2127 (N_2127,N_1993,In_1593);
nand U2128 (N_2128,N_1425,N_1854);
nor U2129 (N_2129,N_1690,N_1776);
xor U2130 (N_2130,In_287,In_2080);
xor U2131 (N_2131,N_1710,N_708);
nand U2132 (N_2132,N_1967,N_1823);
or U2133 (N_2133,N_228,N_890);
and U2134 (N_2134,N_399,N_402);
nor U2135 (N_2135,N_1816,N_1820);
nor U2136 (N_2136,N_1590,N_1528);
or U2137 (N_2137,N_1864,N_1919);
nor U2138 (N_2138,N_1940,N_1828);
and U2139 (N_2139,N_1942,In_208);
nor U2140 (N_2140,N_1756,In_2034);
or U2141 (N_2141,N_1814,N_1848);
and U2142 (N_2142,In_863,N_1875);
and U2143 (N_2143,N_1891,N_1509);
nand U2144 (N_2144,N_1154,N_1830);
nor U2145 (N_2145,N_1716,N_1354);
xnor U2146 (N_2146,N_1511,N_1281);
nor U2147 (N_2147,N_1393,N_1793);
xnor U2148 (N_2148,N_1840,N_1515);
and U2149 (N_2149,N_638,N_1974);
or U2150 (N_2150,N_201,N_1626);
nand U2151 (N_2151,N_1803,N_1883);
and U2152 (N_2152,N_1802,N_1885);
or U2153 (N_2153,In_2483,N_1960);
or U2154 (N_2154,N_1602,N_886);
or U2155 (N_2155,N_1112,N_1186);
nor U2156 (N_2156,N_1962,N_1608);
nand U2157 (N_2157,N_1893,N_637);
xor U2158 (N_2158,N_28,N_1977);
xnor U2159 (N_2159,N_1999,N_1708);
and U2160 (N_2160,N_679,N_1749);
nor U2161 (N_2161,N_1817,N_629);
and U2162 (N_2162,N_1952,N_1752);
nand U2163 (N_2163,N_1550,N_1922);
and U2164 (N_2164,N_1627,N_1915);
nor U2165 (N_2165,N_1735,N_1445);
or U2166 (N_2166,N_123,N_1831);
xnor U2167 (N_2167,N_1728,N_1316);
and U2168 (N_2168,In_1812,N_1847);
and U2169 (N_2169,N_1948,In_616);
nand U2170 (N_2170,N_1941,N_968);
nor U2171 (N_2171,N_1939,N_1782);
xnor U2172 (N_2172,N_273,N_1753);
and U2173 (N_2173,N_1838,N_1813);
nor U2174 (N_2174,N_1825,In_537);
or U2175 (N_2175,N_1898,N_1897);
or U2176 (N_2176,N_1855,N_1910);
and U2177 (N_2177,N_1433,N_1870);
or U2178 (N_2178,In_390,N_1839);
xor U2179 (N_2179,In_1325,N_1889);
or U2180 (N_2180,N_1958,N_1791);
nand U2181 (N_2181,N_1943,N_1285);
xor U2182 (N_2182,N_1388,N_1189);
or U2183 (N_2183,In_1478,N_1934);
nand U2184 (N_2184,N_1981,N_1795);
nand U2185 (N_2185,N_1882,N_278);
nand U2186 (N_2186,N_1744,In_1185);
or U2187 (N_2187,N_1060,N_1865);
nand U2188 (N_2188,N_1166,In_465);
and U2189 (N_2189,N_1925,N_1982);
nor U2190 (N_2190,N_1094,N_1858);
nand U2191 (N_2191,N_1821,In_1107);
and U2192 (N_2192,N_244,N_1268);
and U2193 (N_2193,N_1783,N_1541);
xor U2194 (N_2194,In_1793,N_1853);
or U2195 (N_2195,N_1932,N_1643);
and U2196 (N_2196,N_1395,N_1996);
nand U2197 (N_2197,N_1514,In_1895);
or U2198 (N_2198,N_1924,N_1829);
nand U2199 (N_2199,N_1661,N_1788);
xor U2200 (N_2200,N_1908,N_1985);
and U2201 (N_2201,In_827,N_1938);
or U2202 (N_2202,N_1540,In_1665);
and U2203 (N_2203,N_1792,N_1775);
and U2204 (N_2204,N_1542,N_1846);
xnor U2205 (N_2205,N_1472,N_1876);
or U2206 (N_2206,N_1681,N_1676);
or U2207 (N_2207,N_1818,In_997);
or U2208 (N_2208,N_1522,N_800);
nor U2209 (N_2209,N_1290,N_107);
nand U2210 (N_2210,N_1903,N_1984);
nand U2211 (N_2211,N_1904,N_1463);
nand U2212 (N_2212,N_1583,N_1508);
nor U2213 (N_2213,N_1321,N_1860);
nor U2214 (N_2214,N_1693,N_103);
nor U2215 (N_2215,N_1078,N_1859);
xor U2216 (N_2216,N_1929,N_1871);
and U2217 (N_2217,N_1797,In_138);
or U2218 (N_2218,N_232,N_1852);
xnor U2219 (N_2219,N_1344,N_1547);
xor U2220 (N_2220,N_1576,N_1804);
nor U2221 (N_2221,N_1970,N_1696);
nand U2222 (N_2222,N_1498,N_1956);
or U2223 (N_2223,N_1877,N_1279);
nand U2224 (N_2224,N_1986,N_1836);
nor U2225 (N_2225,In_1577,N_1933);
nand U2226 (N_2226,N_1408,N_1503);
or U2227 (N_2227,N_1343,N_1900);
nor U2228 (N_2228,N_739,N_1754);
or U2229 (N_2229,N_1046,N_1963);
xnor U2230 (N_2230,N_1760,N_1914);
nor U2231 (N_2231,N_1674,N_1156);
or U2232 (N_2232,N_1894,N_888);
and U2233 (N_2233,N_1545,N_1937);
and U2234 (N_2234,N_1554,N_570);
or U2235 (N_2235,N_1827,N_1660);
nand U2236 (N_2236,N_1787,N_1683);
nor U2237 (N_2237,In_1965,N_1747);
nand U2238 (N_2238,N_1998,In_2083);
nand U2239 (N_2239,N_1790,N_1988);
or U2240 (N_2240,N_1766,N_1874);
nor U2241 (N_2241,N_1083,N_1647);
nor U2242 (N_2242,In_1773,In_1982);
or U2243 (N_2243,N_440,N_1659);
xor U2244 (N_2244,N_1991,N_1769);
xnor U2245 (N_2245,In_2079,N_1896);
nand U2246 (N_2246,In_2354,N_1810);
nor U2247 (N_2247,N_1944,N_1868);
xor U2248 (N_2248,N_1800,N_1812);
and U2249 (N_2249,N_1807,N_697);
nand U2250 (N_2250,N_2061,N_2115);
xor U2251 (N_2251,N_2141,N_2173);
nand U2252 (N_2252,N_2021,N_2006);
nor U2253 (N_2253,N_2122,N_2192);
nand U2254 (N_2254,N_2187,N_2209);
nor U2255 (N_2255,N_2167,N_2128);
xnor U2256 (N_2256,N_2155,N_2005);
xor U2257 (N_2257,N_2139,N_2009);
and U2258 (N_2258,N_2012,N_2233);
xnor U2259 (N_2259,N_2180,N_2184);
or U2260 (N_2260,N_2015,N_2077);
or U2261 (N_2261,N_2046,N_2050);
or U2262 (N_2262,N_2095,N_2004);
nand U2263 (N_2263,N_2037,N_2189);
or U2264 (N_2264,N_2071,N_2121);
and U2265 (N_2265,N_2048,N_2099);
xnor U2266 (N_2266,N_2160,N_2244);
xor U2267 (N_2267,N_2178,N_2162);
nand U2268 (N_2268,N_2133,N_2204);
nor U2269 (N_2269,N_2080,N_2194);
xnor U2270 (N_2270,N_2241,N_2148);
or U2271 (N_2271,N_2117,N_2097);
nor U2272 (N_2272,N_2055,N_2172);
nor U2273 (N_2273,N_2216,N_2054);
nor U2274 (N_2274,N_2168,N_2103);
nor U2275 (N_2275,N_2223,N_2056);
and U2276 (N_2276,N_2034,N_2145);
xor U2277 (N_2277,N_2074,N_2063);
nand U2278 (N_2278,N_2066,N_2016);
nand U2279 (N_2279,N_2076,N_2164);
xor U2280 (N_2280,N_2235,N_2142);
xor U2281 (N_2281,N_2199,N_2230);
or U2282 (N_2282,N_2082,N_2035);
nor U2283 (N_2283,N_2070,N_2222);
nand U2284 (N_2284,N_2247,N_2123);
nand U2285 (N_2285,N_2040,N_2088);
or U2286 (N_2286,N_2206,N_2146);
xnor U2287 (N_2287,N_2085,N_2246);
nor U2288 (N_2288,N_2105,N_2170);
nor U2289 (N_2289,N_2190,N_2089);
and U2290 (N_2290,N_2042,N_2157);
xnor U2291 (N_2291,N_2093,N_2113);
nand U2292 (N_2292,N_2159,N_2079);
and U2293 (N_2293,N_2226,N_2182);
nand U2294 (N_2294,N_2196,N_2013);
or U2295 (N_2295,N_2132,N_2130);
and U2296 (N_2296,N_2202,N_2051);
or U2297 (N_2297,N_2098,N_2120);
nor U2298 (N_2298,N_2165,N_2240);
or U2299 (N_2299,N_2210,N_2108);
and U2300 (N_2300,N_2062,N_2030);
xor U2301 (N_2301,N_2221,N_2001);
nand U2302 (N_2302,N_2023,N_2140);
and U2303 (N_2303,N_2101,N_2134);
nand U2304 (N_2304,N_2043,N_2090);
xor U2305 (N_2305,N_2198,N_2067);
and U2306 (N_2306,N_2059,N_2245);
and U2307 (N_2307,N_2144,N_2129);
or U2308 (N_2308,N_2110,N_2169);
and U2309 (N_2309,N_2188,N_2249);
or U2310 (N_2310,N_2242,N_2011);
xnor U2311 (N_2311,N_2237,N_2220);
xor U2312 (N_2312,N_2086,N_2003);
or U2313 (N_2313,N_2143,N_2008);
xor U2314 (N_2314,N_2191,N_2124);
nor U2315 (N_2315,N_2078,N_2248);
nor U2316 (N_2316,N_2064,N_2131);
and U2317 (N_2317,N_2214,N_2068);
xnor U2318 (N_2318,N_2147,N_2243);
or U2319 (N_2319,N_2019,N_2083);
nand U2320 (N_2320,N_2096,N_2150);
or U2321 (N_2321,N_2065,N_2031);
or U2322 (N_2322,N_2002,N_2020);
nor U2323 (N_2323,N_2044,N_2022);
or U2324 (N_2324,N_2177,N_2018);
nand U2325 (N_2325,N_2036,N_2239);
xnor U2326 (N_2326,N_2116,N_2236);
or U2327 (N_2327,N_2215,N_2014);
nand U2328 (N_2328,N_2084,N_2137);
nor U2329 (N_2329,N_2111,N_2026);
and U2330 (N_2330,N_2017,N_2126);
nor U2331 (N_2331,N_2234,N_2218);
and U2332 (N_2332,N_2029,N_2156);
or U2333 (N_2333,N_2112,N_2038);
and U2334 (N_2334,N_2060,N_2114);
nor U2335 (N_2335,N_2053,N_2197);
xnor U2336 (N_2336,N_2109,N_2028);
nor U2337 (N_2337,N_2049,N_2201);
or U2338 (N_2338,N_2175,N_2224);
and U2339 (N_2339,N_2207,N_2045);
and U2340 (N_2340,N_2152,N_2024);
or U2341 (N_2341,N_2231,N_2125);
and U2342 (N_2342,N_2213,N_2104);
or U2343 (N_2343,N_2158,N_2195);
nor U2344 (N_2344,N_2163,N_2229);
nor U2345 (N_2345,N_2047,N_2052);
or U2346 (N_2346,N_2010,N_2039);
and U2347 (N_2347,N_2136,N_2208);
nand U2348 (N_2348,N_2149,N_2100);
xnor U2349 (N_2349,N_2091,N_2183);
and U2350 (N_2350,N_2227,N_2219);
or U2351 (N_2351,N_2193,N_2107);
or U2352 (N_2352,N_2154,N_2000);
or U2353 (N_2353,N_2138,N_2166);
nand U2354 (N_2354,N_2228,N_2032);
xor U2355 (N_2355,N_2161,N_2135);
and U2356 (N_2356,N_2087,N_2238);
nand U2357 (N_2357,N_2094,N_2176);
or U2358 (N_2358,N_2203,N_2069);
or U2359 (N_2359,N_2119,N_2186);
nor U2360 (N_2360,N_2225,N_2171);
nor U2361 (N_2361,N_2153,N_2212);
xnor U2362 (N_2362,N_2211,N_2200);
and U2363 (N_2363,N_2072,N_2057);
or U2364 (N_2364,N_2151,N_2033);
and U2365 (N_2365,N_2118,N_2181);
and U2366 (N_2366,N_2058,N_2092);
or U2367 (N_2367,N_2007,N_2179);
nand U2368 (N_2368,N_2185,N_2174);
or U2369 (N_2369,N_2217,N_2205);
xnor U2370 (N_2370,N_2041,N_2025);
and U2371 (N_2371,N_2106,N_2232);
or U2372 (N_2372,N_2102,N_2081);
or U2373 (N_2373,N_2127,N_2075);
and U2374 (N_2374,N_2027,N_2073);
xor U2375 (N_2375,N_2203,N_2086);
nor U2376 (N_2376,N_2069,N_2060);
nand U2377 (N_2377,N_2014,N_2194);
nor U2378 (N_2378,N_2128,N_2208);
or U2379 (N_2379,N_2181,N_2203);
nand U2380 (N_2380,N_2101,N_2010);
or U2381 (N_2381,N_2040,N_2242);
and U2382 (N_2382,N_2132,N_2111);
xnor U2383 (N_2383,N_2121,N_2245);
nand U2384 (N_2384,N_2225,N_2058);
xnor U2385 (N_2385,N_2135,N_2099);
or U2386 (N_2386,N_2195,N_2084);
xnor U2387 (N_2387,N_2088,N_2241);
xor U2388 (N_2388,N_2227,N_2085);
nor U2389 (N_2389,N_2209,N_2133);
xnor U2390 (N_2390,N_2172,N_2129);
or U2391 (N_2391,N_2140,N_2065);
nand U2392 (N_2392,N_2214,N_2164);
nor U2393 (N_2393,N_2115,N_2106);
nand U2394 (N_2394,N_2080,N_2118);
xnor U2395 (N_2395,N_2205,N_2207);
nor U2396 (N_2396,N_2235,N_2215);
and U2397 (N_2397,N_2230,N_2241);
nor U2398 (N_2398,N_2021,N_2097);
nor U2399 (N_2399,N_2070,N_2238);
nor U2400 (N_2400,N_2047,N_2026);
xnor U2401 (N_2401,N_2090,N_2042);
nor U2402 (N_2402,N_2084,N_2191);
xnor U2403 (N_2403,N_2030,N_2031);
and U2404 (N_2404,N_2240,N_2179);
xnor U2405 (N_2405,N_2108,N_2051);
and U2406 (N_2406,N_2229,N_2107);
nand U2407 (N_2407,N_2074,N_2058);
xnor U2408 (N_2408,N_2230,N_2144);
and U2409 (N_2409,N_2218,N_2024);
or U2410 (N_2410,N_2052,N_2133);
and U2411 (N_2411,N_2248,N_2199);
xor U2412 (N_2412,N_2162,N_2059);
or U2413 (N_2413,N_2049,N_2138);
and U2414 (N_2414,N_2137,N_2138);
nand U2415 (N_2415,N_2014,N_2048);
nand U2416 (N_2416,N_2020,N_2007);
nor U2417 (N_2417,N_2172,N_2037);
and U2418 (N_2418,N_2075,N_2114);
or U2419 (N_2419,N_2017,N_2074);
and U2420 (N_2420,N_2236,N_2073);
and U2421 (N_2421,N_2220,N_2138);
nor U2422 (N_2422,N_2033,N_2022);
nand U2423 (N_2423,N_2027,N_2106);
nor U2424 (N_2424,N_2065,N_2056);
nand U2425 (N_2425,N_2010,N_2171);
and U2426 (N_2426,N_2028,N_2232);
or U2427 (N_2427,N_2162,N_2047);
nand U2428 (N_2428,N_2152,N_2233);
nor U2429 (N_2429,N_2145,N_2102);
nor U2430 (N_2430,N_2158,N_2228);
and U2431 (N_2431,N_2012,N_2195);
nand U2432 (N_2432,N_2183,N_2169);
xor U2433 (N_2433,N_2243,N_2248);
and U2434 (N_2434,N_2041,N_2245);
and U2435 (N_2435,N_2035,N_2018);
nand U2436 (N_2436,N_2242,N_2050);
xor U2437 (N_2437,N_2140,N_2121);
nand U2438 (N_2438,N_2053,N_2115);
and U2439 (N_2439,N_2054,N_2146);
nor U2440 (N_2440,N_2188,N_2179);
nand U2441 (N_2441,N_2172,N_2192);
or U2442 (N_2442,N_2187,N_2161);
nor U2443 (N_2443,N_2094,N_2220);
nor U2444 (N_2444,N_2074,N_2206);
and U2445 (N_2445,N_2034,N_2215);
xnor U2446 (N_2446,N_2165,N_2147);
nor U2447 (N_2447,N_2229,N_2241);
nor U2448 (N_2448,N_2187,N_2045);
nand U2449 (N_2449,N_2182,N_2082);
xor U2450 (N_2450,N_2242,N_2059);
or U2451 (N_2451,N_2052,N_2153);
or U2452 (N_2452,N_2186,N_2049);
or U2453 (N_2453,N_2239,N_2206);
and U2454 (N_2454,N_2157,N_2195);
nand U2455 (N_2455,N_2179,N_2105);
or U2456 (N_2456,N_2228,N_2156);
or U2457 (N_2457,N_2041,N_2160);
or U2458 (N_2458,N_2059,N_2194);
nor U2459 (N_2459,N_2003,N_2048);
or U2460 (N_2460,N_2184,N_2047);
or U2461 (N_2461,N_2060,N_2180);
nand U2462 (N_2462,N_2188,N_2194);
xor U2463 (N_2463,N_2125,N_2154);
nand U2464 (N_2464,N_2038,N_2040);
nor U2465 (N_2465,N_2123,N_2026);
and U2466 (N_2466,N_2237,N_2009);
nand U2467 (N_2467,N_2149,N_2013);
and U2468 (N_2468,N_2033,N_2106);
nand U2469 (N_2469,N_2069,N_2032);
nand U2470 (N_2470,N_2234,N_2169);
nor U2471 (N_2471,N_2173,N_2089);
nand U2472 (N_2472,N_2091,N_2249);
nand U2473 (N_2473,N_2027,N_2178);
or U2474 (N_2474,N_2092,N_2013);
or U2475 (N_2475,N_2060,N_2230);
and U2476 (N_2476,N_2093,N_2141);
xnor U2477 (N_2477,N_2140,N_2208);
nand U2478 (N_2478,N_2109,N_2057);
nand U2479 (N_2479,N_2169,N_2019);
and U2480 (N_2480,N_2028,N_2182);
nand U2481 (N_2481,N_2131,N_2049);
xnor U2482 (N_2482,N_2033,N_2155);
nor U2483 (N_2483,N_2136,N_2048);
xor U2484 (N_2484,N_2245,N_2210);
and U2485 (N_2485,N_2197,N_2150);
and U2486 (N_2486,N_2124,N_2231);
or U2487 (N_2487,N_2087,N_2188);
nand U2488 (N_2488,N_2021,N_2151);
and U2489 (N_2489,N_2173,N_2142);
and U2490 (N_2490,N_2244,N_2221);
or U2491 (N_2491,N_2093,N_2123);
and U2492 (N_2492,N_2104,N_2182);
nor U2493 (N_2493,N_2218,N_2163);
xnor U2494 (N_2494,N_2089,N_2042);
xnor U2495 (N_2495,N_2025,N_2225);
or U2496 (N_2496,N_2198,N_2149);
nor U2497 (N_2497,N_2083,N_2047);
nand U2498 (N_2498,N_2175,N_2032);
xnor U2499 (N_2499,N_2147,N_2056);
and U2500 (N_2500,N_2306,N_2444);
or U2501 (N_2501,N_2370,N_2256);
and U2502 (N_2502,N_2482,N_2434);
xor U2503 (N_2503,N_2255,N_2339);
or U2504 (N_2504,N_2469,N_2372);
or U2505 (N_2505,N_2353,N_2377);
and U2506 (N_2506,N_2304,N_2374);
or U2507 (N_2507,N_2293,N_2442);
xnor U2508 (N_2508,N_2410,N_2390);
nand U2509 (N_2509,N_2385,N_2498);
and U2510 (N_2510,N_2458,N_2396);
xnor U2511 (N_2511,N_2365,N_2425);
nor U2512 (N_2512,N_2398,N_2317);
xor U2513 (N_2513,N_2429,N_2294);
and U2514 (N_2514,N_2481,N_2470);
and U2515 (N_2515,N_2344,N_2438);
nor U2516 (N_2516,N_2412,N_2364);
or U2517 (N_2517,N_2300,N_2287);
or U2518 (N_2518,N_2310,N_2460);
nor U2519 (N_2519,N_2435,N_2312);
xor U2520 (N_2520,N_2457,N_2318);
or U2521 (N_2521,N_2266,N_2269);
xor U2522 (N_2522,N_2309,N_2290);
nand U2523 (N_2523,N_2424,N_2328);
or U2524 (N_2524,N_2314,N_2267);
or U2525 (N_2525,N_2325,N_2378);
nor U2526 (N_2526,N_2348,N_2295);
nand U2527 (N_2527,N_2291,N_2368);
or U2528 (N_2528,N_2386,N_2416);
nor U2529 (N_2529,N_2433,N_2268);
nand U2530 (N_2530,N_2260,N_2452);
nand U2531 (N_2531,N_2430,N_2451);
xor U2532 (N_2532,N_2487,N_2395);
xnor U2533 (N_2533,N_2375,N_2413);
and U2534 (N_2534,N_2338,N_2330);
nand U2535 (N_2535,N_2308,N_2379);
or U2536 (N_2536,N_2384,N_2358);
and U2537 (N_2537,N_2285,N_2273);
nor U2538 (N_2538,N_2278,N_2337);
xor U2539 (N_2539,N_2381,N_2321);
nand U2540 (N_2540,N_2371,N_2406);
and U2541 (N_2541,N_2419,N_2261);
or U2542 (N_2542,N_2329,N_2391);
xor U2543 (N_2543,N_2263,N_2454);
and U2544 (N_2544,N_2292,N_2490);
nand U2545 (N_2545,N_2251,N_2362);
nor U2546 (N_2546,N_2288,N_2252);
or U2547 (N_2547,N_2483,N_2352);
and U2548 (N_2548,N_2316,N_2376);
and U2549 (N_2549,N_2408,N_2473);
and U2550 (N_2550,N_2280,N_2389);
xnor U2551 (N_2551,N_2305,N_2356);
nand U2552 (N_2552,N_2404,N_2296);
or U2553 (N_2553,N_2421,N_2476);
or U2554 (N_2554,N_2415,N_2427);
nand U2555 (N_2555,N_2367,N_2271);
nor U2556 (N_2556,N_2258,N_2496);
and U2557 (N_2557,N_2281,N_2467);
xor U2558 (N_2558,N_2313,N_2324);
and U2559 (N_2559,N_2422,N_2491);
nand U2560 (N_2560,N_2387,N_2439);
nand U2561 (N_2561,N_2488,N_2259);
xnor U2562 (N_2562,N_2453,N_2354);
or U2563 (N_2563,N_2382,N_2462);
xor U2564 (N_2564,N_2445,N_2326);
xnor U2565 (N_2565,N_2493,N_2409);
and U2566 (N_2566,N_2264,N_2345);
nand U2567 (N_2567,N_2283,N_2274);
or U2568 (N_2568,N_2361,N_2414);
xor U2569 (N_2569,N_2399,N_2340);
and U2570 (N_2570,N_2357,N_2363);
xor U2571 (N_2571,N_2299,N_2342);
nor U2572 (N_2572,N_2405,N_2322);
and U2573 (N_2573,N_2286,N_2347);
nor U2574 (N_2574,N_2298,N_2349);
or U2575 (N_2575,N_2254,N_2284);
and U2576 (N_2576,N_2277,N_2383);
nand U2577 (N_2577,N_2323,N_2455);
nor U2578 (N_2578,N_2449,N_2475);
or U2579 (N_2579,N_2464,N_2388);
and U2580 (N_2580,N_2411,N_2486);
and U2581 (N_2581,N_2463,N_2297);
nor U2582 (N_2582,N_2436,N_2289);
nand U2583 (N_2583,N_2336,N_2447);
xnor U2584 (N_2584,N_2393,N_2332);
xnor U2585 (N_2585,N_2495,N_2450);
nand U2586 (N_2586,N_2343,N_2279);
xor U2587 (N_2587,N_2275,N_2466);
nand U2588 (N_2588,N_2400,N_2392);
or U2589 (N_2589,N_2335,N_2333);
and U2590 (N_2590,N_2446,N_2485);
nand U2591 (N_2591,N_2423,N_2428);
or U2592 (N_2592,N_2471,N_2319);
or U2593 (N_2593,N_2468,N_2403);
nor U2594 (N_2594,N_2474,N_2461);
xor U2595 (N_2595,N_2253,N_2373);
nand U2596 (N_2596,N_2303,N_2426);
or U2597 (N_2597,N_2407,N_2331);
or U2598 (N_2598,N_2489,N_2262);
xnor U2599 (N_2599,N_2437,N_2459);
nand U2600 (N_2600,N_2478,N_2350);
and U2601 (N_2601,N_2394,N_2497);
xor U2602 (N_2602,N_2441,N_2443);
xor U2603 (N_2603,N_2355,N_2472);
and U2604 (N_2604,N_2380,N_2270);
xnor U2605 (N_2605,N_2359,N_2418);
and U2606 (N_2606,N_2351,N_2272);
nand U2607 (N_2607,N_2302,N_2315);
nand U2608 (N_2608,N_2257,N_2499);
or U2609 (N_2609,N_2456,N_2341);
and U2610 (N_2610,N_2307,N_2402);
or U2611 (N_2611,N_2448,N_2250);
or U2612 (N_2612,N_2282,N_2366);
xnor U2613 (N_2613,N_2484,N_2465);
and U2614 (N_2614,N_2311,N_2417);
nand U2615 (N_2615,N_2401,N_2440);
nand U2616 (N_2616,N_2397,N_2265);
or U2617 (N_2617,N_2477,N_2494);
and U2618 (N_2618,N_2301,N_2432);
and U2619 (N_2619,N_2276,N_2327);
nand U2620 (N_2620,N_2492,N_2479);
nor U2621 (N_2621,N_2420,N_2334);
nand U2622 (N_2622,N_2431,N_2320);
or U2623 (N_2623,N_2346,N_2369);
and U2624 (N_2624,N_2360,N_2480);
and U2625 (N_2625,N_2370,N_2455);
nand U2626 (N_2626,N_2464,N_2305);
nand U2627 (N_2627,N_2427,N_2385);
xnor U2628 (N_2628,N_2359,N_2449);
or U2629 (N_2629,N_2443,N_2379);
nand U2630 (N_2630,N_2484,N_2491);
or U2631 (N_2631,N_2399,N_2394);
nand U2632 (N_2632,N_2377,N_2444);
or U2633 (N_2633,N_2326,N_2380);
or U2634 (N_2634,N_2482,N_2444);
or U2635 (N_2635,N_2341,N_2464);
and U2636 (N_2636,N_2276,N_2439);
nor U2637 (N_2637,N_2309,N_2465);
or U2638 (N_2638,N_2460,N_2396);
and U2639 (N_2639,N_2297,N_2437);
and U2640 (N_2640,N_2402,N_2392);
nand U2641 (N_2641,N_2464,N_2371);
and U2642 (N_2642,N_2324,N_2470);
and U2643 (N_2643,N_2268,N_2347);
nand U2644 (N_2644,N_2311,N_2454);
xnor U2645 (N_2645,N_2287,N_2376);
and U2646 (N_2646,N_2476,N_2372);
nor U2647 (N_2647,N_2290,N_2269);
nand U2648 (N_2648,N_2391,N_2348);
and U2649 (N_2649,N_2472,N_2405);
nor U2650 (N_2650,N_2450,N_2274);
and U2651 (N_2651,N_2399,N_2342);
nand U2652 (N_2652,N_2451,N_2443);
or U2653 (N_2653,N_2327,N_2432);
and U2654 (N_2654,N_2321,N_2477);
or U2655 (N_2655,N_2291,N_2475);
xor U2656 (N_2656,N_2262,N_2455);
and U2657 (N_2657,N_2294,N_2421);
and U2658 (N_2658,N_2358,N_2411);
nand U2659 (N_2659,N_2290,N_2302);
and U2660 (N_2660,N_2304,N_2339);
and U2661 (N_2661,N_2380,N_2363);
nor U2662 (N_2662,N_2476,N_2405);
or U2663 (N_2663,N_2471,N_2487);
xor U2664 (N_2664,N_2440,N_2478);
nand U2665 (N_2665,N_2412,N_2344);
nand U2666 (N_2666,N_2252,N_2350);
xor U2667 (N_2667,N_2406,N_2420);
nand U2668 (N_2668,N_2305,N_2373);
nor U2669 (N_2669,N_2320,N_2299);
nand U2670 (N_2670,N_2276,N_2470);
xnor U2671 (N_2671,N_2393,N_2354);
xor U2672 (N_2672,N_2460,N_2259);
xor U2673 (N_2673,N_2383,N_2251);
nand U2674 (N_2674,N_2407,N_2432);
or U2675 (N_2675,N_2362,N_2413);
xnor U2676 (N_2676,N_2267,N_2308);
xor U2677 (N_2677,N_2289,N_2302);
nand U2678 (N_2678,N_2436,N_2265);
or U2679 (N_2679,N_2295,N_2423);
or U2680 (N_2680,N_2302,N_2499);
and U2681 (N_2681,N_2332,N_2370);
xnor U2682 (N_2682,N_2381,N_2331);
and U2683 (N_2683,N_2375,N_2261);
nor U2684 (N_2684,N_2294,N_2442);
nand U2685 (N_2685,N_2324,N_2284);
and U2686 (N_2686,N_2468,N_2493);
nor U2687 (N_2687,N_2331,N_2413);
nand U2688 (N_2688,N_2273,N_2467);
and U2689 (N_2689,N_2308,N_2263);
nand U2690 (N_2690,N_2432,N_2458);
or U2691 (N_2691,N_2437,N_2450);
and U2692 (N_2692,N_2483,N_2383);
nor U2693 (N_2693,N_2331,N_2498);
xor U2694 (N_2694,N_2308,N_2352);
xnor U2695 (N_2695,N_2411,N_2284);
xor U2696 (N_2696,N_2464,N_2293);
nand U2697 (N_2697,N_2497,N_2456);
and U2698 (N_2698,N_2461,N_2396);
nor U2699 (N_2699,N_2462,N_2472);
xor U2700 (N_2700,N_2286,N_2365);
nand U2701 (N_2701,N_2373,N_2399);
or U2702 (N_2702,N_2323,N_2499);
and U2703 (N_2703,N_2335,N_2401);
nand U2704 (N_2704,N_2358,N_2261);
xnor U2705 (N_2705,N_2257,N_2311);
or U2706 (N_2706,N_2380,N_2335);
nor U2707 (N_2707,N_2446,N_2473);
nor U2708 (N_2708,N_2465,N_2279);
xnor U2709 (N_2709,N_2251,N_2293);
xnor U2710 (N_2710,N_2295,N_2327);
nor U2711 (N_2711,N_2356,N_2405);
and U2712 (N_2712,N_2309,N_2448);
or U2713 (N_2713,N_2348,N_2480);
and U2714 (N_2714,N_2353,N_2255);
and U2715 (N_2715,N_2307,N_2376);
and U2716 (N_2716,N_2299,N_2443);
nor U2717 (N_2717,N_2332,N_2438);
or U2718 (N_2718,N_2475,N_2328);
and U2719 (N_2719,N_2280,N_2437);
nor U2720 (N_2720,N_2363,N_2479);
xnor U2721 (N_2721,N_2457,N_2353);
nor U2722 (N_2722,N_2357,N_2424);
or U2723 (N_2723,N_2411,N_2436);
nor U2724 (N_2724,N_2463,N_2372);
or U2725 (N_2725,N_2283,N_2317);
and U2726 (N_2726,N_2442,N_2447);
xnor U2727 (N_2727,N_2369,N_2324);
or U2728 (N_2728,N_2346,N_2459);
xnor U2729 (N_2729,N_2428,N_2269);
and U2730 (N_2730,N_2473,N_2394);
nand U2731 (N_2731,N_2498,N_2405);
nor U2732 (N_2732,N_2382,N_2335);
nand U2733 (N_2733,N_2494,N_2294);
or U2734 (N_2734,N_2492,N_2330);
nand U2735 (N_2735,N_2396,N_2456);
nand U2736 (N_2736,N_2398,N_2343);
and U2737 (N_2737,N_2458,N_2292);
xor U2738 (N_2738,N_2482,N_2462);
and U2739 (N_2739,N_2307,N_2269);
or U2740 (N_2740,N_2393,N_2389);
nor U2741 (N_2741,N_2360,N_2315);
xnor U2742 (N_2742,N_2329,N_2361);
or U2743 (N_2743,N_2387,N_2429);
or U2744 (N_2744,N_2455,N_2372);
nand U2745 (N_2745,N_2455,N_2490);
nand U2746 (N_2746,N_2421,N_2437);
or U2747 (N_2747,N_2487,N_2273);
nand U2748 (N_2748,N_2325,N_2412);
nand U2749 (N_2749,N_2377,N_2450);
or U2750 (N_2750,N_2500,N_2593);
and U2751 (N_2751,N_2559,N_2552);
or U2752 (N_2752,N_2725,N_2659);
xor U2753 (N_2753,N_2691,N_2657);
xor U2754 (N_2754,N_2640,N_2608);
xnor U2755 (N_2755,N_2623,N_2699);
xnor U2756 (N_2756,N_2545,N_2674);
nor U2757 (N_2757,N_2537,N_2600);
and U2758 (N_2758,N_2558,N_2653);
nor U2759 (N_2759,N_2508,N_2630);
or U2760 (N_2760,N_2643,N_2717);
and U2761 (N_2761,N_2732,N_2745);
nor U2762 (N_2762,N_2727,N_2512);
nor U2763 (N_2763,N_2567,N_2681);
or U2764 (N_2764,N_2566,N_2531);
or U2765 (N_2765,N_2724,N_2604);
nand U2766 (N_2766,N_2532,N_2549);
or U2767 (N_2767,N_2562,N_2599);
xor U2768 (N_2768,N_2527,N_2580);
or U2769 (N_2769,N_2716,N_2603);
and U2770 (N_2770,N_2694,N_2633);
xor U2771 (N_2771,N_2597,N_2718);
and U2772 (N_2772,N_2707,N_2510);
xor U2773 (N_2773,N_2607,N_2733);
or U2774 (N_2774,N_2652,N_2726);
nand U2775 (N_2775,N_2561,N_2649);
nor U2776 (N_2776,N_2719,N_2587);
or U2777 (N_2777,N_2679,N_2555);
nor U2778 (N_2778,N_2686,N_2617);
or U2779 (N_2779,N_2620,N_2598);
nand U2780 (N_2780,N_2706,N_2668);
nor U2781 (N_2781,N_2589,N_2517);
and U2782 (N_2782,N_2737,N_2525);
nor U2783 (N_2783,N_2667,N_2504);
and U2784 (N_2784,N_2722,N_2648);
and U2785 (N_2785,N_2601,N_2611);
and U2786 (N_2786,N_2502,N_2646);
nor U2787 (N_2787,N_2538,N_2635);
nor U2788 (N_2788,N_2588,N_2728);
and U2789 (N_2789,N_2557,N_2516);
nand U2790 (N_2790,N_2582,N_2542);
xor U2791 (N_2791,N_2696,N_2610);
nand U2792 (N_2792,N_2678,N_2625);
nand U2793 (N_2793,N_2569,N_2735);
xnor U2794 (N_2794,N_2581,N_2505);
nor U2795 (N_2795,N_2594,N_2535);
or U2796 (N_2796,N_2677,N_2613);
or U2797 (N_2797,N_2683,N_2606);
xnor U2798 (N_2798,N_2536,N_2528);
or U2799 (N_2799,N_2628,N_2574);
and U2800 (N_2800,N_2539,N_2665);
and U2801 (N_2801,N_2746,N_2688);
or U2802 (N_2802,N_2669,N_2742);
or U2803 (N_2803,N_2615,N_2583);
and U2804 (N_2804,N_2655,N_2738);
and U2805 (N_2805,N_2710,N_2642);
or U2806 (N_2806,N_2698,N_2689);
xnor U2807 (N_2807,N_2663,N_2743);
or U2808 (N_2808,N_2627,N_2687);
xnor U2809 (N_2809,N_2543,N_2529);
nand U2810 (N_2810,N_2656,N_2704);
nand U2811 (N_2811,N_2634,N_2629);
nand U2812 (N_2812,N_2618,N_2711);
nand U2813 (N_2813,N_2697,N_2546);
or U2814 (N_2814,N_2730,N_2513);
and U2815 (N_2815,N_2602,N_2612);
xnor U2816 (N_2816,N_2712,N_2523);
or U2817 (N_2817,N_2556,N_2700);
and U2818 (N_2818,N_2585,N_2739);
and U2819 (N_2819,N_2644,N_2553);
and U2820 (N_2820,N_2564,N_2541);
and U2821 (N_2821,N_2636,N_2650);
and U2822 (N_2822,N_2720,N_2721);
xnor U2823 (N_2823,N_2747,N_2572);
and U2824 (N_2824,N_2664,N_2637);
nor U2825 (N_2825,N_2501,N_2560);
nor U2826 (N_2826,N_2590,N_2736);
and U2827 (N_2827,N_2748,N_2509);
nor U2828 (N_2828,N_2519,N_2596);
and U2829 (N_2829,N_2544,N_2575);
xor U2830 (N_2830,N_2714,N_2661);
xnor U2831 (N_2831,N_2565,N_2616);
nand U2832 (N_2832,N_2548,N_2507);
and U2833 (N_2833,N_2530,N_2568);
or U2834 (N_2834,N_2658,N_2676);
nand U2835 (N_2835,N_2662,N_2708);
xor U2836 (N_2836,N_2550,N_2723);
and U2837 (N_2837,N_2684,N_2547);
xnor U2838 (N_2838,N_2702,N_2563);
or U2839 (N_2839,N_2654,N_2647);
nor U2840 (N_2840,N_2503,N_2534);
and U2841 (N_2841,N_2540,N_2692);
nand U2842 (N_2842,N_2595,N_2631);
and U2843 (N_2843,N_2605,N_2690);
and U2844 (N_2844,N_2639,N_2632);
and U2845 (N_2845,N_2705,N_2713);
or U2846 (N_2846,N_2666,N_2573);
nand U2847 (N_2847,N_2577,N_2680);
xnor U2848 (N_2848,N_2675,N_2554);
xnor U2849 (N_2849,N_2524,N_2571);
or U2850 (N_2850,N_2609,N_2621);
nand U2851 (N_2851,N_2715,N_2520);
xor U2852 (N_2852,N_2506,N_2522);
nor U2853 (N_2853,N_2729,N_2682);
and U2854 (N_2854,N_2685,N_2570);
nor U2855 (N_2855,N_2671,N_2709);
nor U2856 (N_2856,N_2514,N_2703);
xor U2857 (N_2857,N_2584,N_2660);
xnor U2858 (N_2858,N_2672,N_2624);
and U2859 (N_2859,N_2511,N_2579);
and U2860 (N_2860,N_2626,N_2638);
xnor U2861 (N_2861,N_2576,N_2521);
or U2862 (N_2862,N_2622,N_2741);
and U2863 (N_2863,N_2695,N_2591);
and U2864 (N_2864,N_2619,N_2614);
xor U2865 (N_2865,N_2731,N_2749);
or U2866 (N_2866,N_2526,N_2578);
xor U2867 (N_2867,N_2533,N_2518);
and U2868 (N_2868,N_2515,N_2551);
xor U2869 (N_2869,N_2670,N_2641);
and U2870 (N_2870,N_2701,N_2673);
or U2871 (N_2871,N_2651,N_2645);
and U2872 (N_2872,N_2740,N_2744);
xor U2873 (N_2873,N_2586,N_2693);
or U2874 (N_2874,N_2592,N_2734);
and U2875 (N_2875,N_2579,N_2593);
nand U2876 (N_2876,N_2590,N_2673);
or U2877 (N_2877,N_2720,N_2679);
nand U2878 (N_2878,N_2509,N_2580);
or U2879 (N_2879,N_2679,N_2517);
and U2880 (N_2880,N_2621,N_2640);
or U2881 (N_2881,N_2591,N_2521);
nor U2882 (N_2882,N_2674,N_2551);
nand U2883 (N_2883,N_2529,N_2699);
and U2884 (N_2884,N_2664,N_2520);
or U2885 (N_2885,N_2635,N_2597);
nor U2886 (N_2886,N_2654,N_2622);
nor U2887 (N_2887,N_2517,N_2578);
and U2888 (N_2888,N_2513,N_2550);
or U2889 (N_2889,N_2614,N_2721);
nor U2890 (N_2890,N_2714,N_2691);
and U2891 (N_2891,N_2612,N_2692);
and U2892 (N_2892,N_2543,N_2509);
and U2893 (N_2893,N_2701,N_2689);
xnor U2894 (N_2894,N_2624,N_2506);
xnor U2895 (N_2895,N_2653,N_2668);
nor U2896 (N_2896,N_2715,N_2575);
nor U2897 (N_2897,N_2520,N_2737);
nor U2898 (N_2898,N_2648,N_2609);
and U2899 (N_2899,N_2673,N_2554);
or U2900 (N_2900,N_2565,N_2655);
and U2901 (N_2901,N_2534,N_2674);
xor U2902 (N_2902,N_2644,N_2715);
and U2903 (N_2903,N_2733,N_2663);
nand U2904 (N_2904,N_2632,N_2621);
or U2905 (N_2905,N_2658,N_2584);
or U2906 (N_2906,N_2682,N_2706);
and U2907 (N_2907,N_2658,N_2665);
or U2908 (N_2908,N_2612,N_2620);
xnor U2909 (N_2909,N_2704,N_2509);
xnor U2910 (N_2910,N_2580,N_2650);
nor U2911 (N_2911,N_2698,N_2709);
nor U2912 (N_2912,N_2651,N_2556);
or U2913 (N_2913,N_2633,N_2698);
nand U2914 (N_2914,N_2541,N_2591);
and U2915 (N_2915,N_2736,N_2632);
xor U2916 (N_2916,N_2656,N_2651);
nor U2917 (N_2917,N_2558,N_2588);
nor U2918 (N_2918,N_2608,N_2528);
nand U2919 (N_2919,N_2554,N_2660);
and U2920 (N_2920,N_2515,N_2677);
and U2921 (N_2921,N_2572,N_2743);
and U2922 (N_2922,N_2572,N_2540);
xor U2923 (N_2923,N_2573,N_2531);
nor U2924 (N_2924,N_2569,N_2734);
nor U2925 (N_2925,N_2511,N_2615);
nor U2926 (N_2926,N_2708,N_2727);
and U2927 (N_2927,N_2556,N_2542);
nor U2928 (N_2928,N_2519,N_2724);
or U2929 (N_2929,N_2709,N_2536);
xnor U2930 (N_2930,N_2557,N_2720);
xnor U2931 (N_2931,N_2511,N_2748);
nand U2932 (N_2932,N_2629,N_2536);
and U2933 (N_2933,N_2523,N_2711);
nand U2934 (N_2934,N_2702,N_2515);
nand U2935 (N_2935,N_2534,N_2712);
xor U2936 (N_2936,N_2563,N_2679);
xor U2937 (N_2937,N_2749,N_2725);
nand U2938 (N_2938,N_2529,N_2660);
or U2939 (N_2939,N_2612,N_2553);
nand U2940 (N_2940,N_2700,N_2694);
nor U2941 (N_2941,N_2500,N_2647);
xor U2942 (N_2942,N_2704,N_2539);
and U2943 (N_2943,N_2685,N_2585);
or U2944 (N_2944,N_2520,N_2554);
or U2945 (N_2945,N_2506,N_2681);
xor U2946 (N_2946,N_2637,N_2707);
nand U2947 (N_2947,N_2597,N_2585);
and U2948 (N_2948,N_2510,N_2537);
or U2949 (N_2949,N_2637,N_2727);
or U2950 (N_2950,N_2542,N_2701);
or U2951 (N_2951,N_2524,N_2564);
and U2952 (N_2952,N_2646,N_2737);
and U2953 (N_2953,N_2504,N_2570);
and U2954 (N_2954,N_2509,N_2582);
and U2955 (N_2955,N_2690,N_2663);
xnor U2956 (N_2956,N_2716,N_2581);
or U2957 (N_2957,N_2586,N_2647);
and U2958 (N_2958,N_2739,N_2695);
xor U2959 (N_2959,N_2537,N_2506);
or U2960 (N_2960,N_2725,N_2675);
and U2961 (N_2961,N_2522,N_2627);
nand U2962 (N_2962,N_2621,N_2675);
or U2963 (N_2963,N_2628,N_2616);
nand U2964 (N_2964,N_2547,N_2641);
nor U2965 (N_2965,N_2720,N_2546);
and U2966 (N_2966,N_2550,N_2592);
nand U2967 (N_2967,N_2647,N_2576);
xnor U2968 (N_2968,N_2633,N_2512);
nor U2969 (N_2969,N_2727,N_2526);
and U2970 (N_2970,N_2504,N_2731);
and U2971 (N_2971,N_2735,N_2655);
or U2972 (N_2972,N_2658,N_2529);
nand U2973 (N_2973,N_2616,N_2740);
xor U2974 (N_2974,N_2580,N_2713);
nand U2975 (N_2975,N_2639,N_2638);
nand U2976 (N_2976,N_2581,N_2745);
nand U2977 (N_2977,N_2519,N_2613);
nand U2978 (N_2978,N_2704,N_2712);
nor U2979 (N_2979,N_2570,N_2642);
xnor U2980 (N_2980,N_2729,N_2736);
or U2981 (N_2981,N_2529,N_2680);
or U2982 (N_2982,N_2613,N_2525);
xnor U2983 (N_2983,N_2502,N_2656);
nor U2984 (N_2984,N_2647,N_2638);
nor U2985 (N_2985,N_2516,N_2645);
and U2986 (N_2986,N_2730,N_2749);
nand U2987 (N_2987,N_2641,N_2720);
or U2988 (N_2988,N_2581,N_2701);
nor U2989 (N_2989,N_2732,N_2557);
nor U2990 (N_2990,N_2624,N_2562);
and U2991 (N_2991,N_2623,N_2721);
and U2992 (N_2992,N_2563,N_2667);
xor U2993 (N_2993,N_2610,N_2691);
and U2994 (N_2994,N_2548,N_2600);
or U2995 (N_2995,N_2735,N_2530);
xnor U2996 (N_2996,N_2692,N_2530);
or U2997 (N_2997,N_2618,N_2631);
and U2998 (N_2998,N_2511,N_2735);
nor U2999 (N_2999,N_2722,N_2596);
xor U3000 (N_3000,N_2902,N_2851);
xnor U3001 (N_3001,N_2929,N_2819);
and U3002 (N_3002,N_2756,N_2903);
and U3003 (N_3003,N_2783,N_2925);
nand U3004 (N_3004,N_2838,N_2958);
xnor U3005 (N_3005,N_2764,N_2824);
nand U3006 (N_3006,N_2750,N_2916);
xnor U3007 (N_3007,N_2897,N_2922);
nand U3008 (N_3008,N_2804,N_2955);
nand U3009 (N_3009,N_2842,N_2927);
and U3010 (N_3010,N_2844,N_2928);
xnor U3011 (N_3011,N_2785,N_2891);
nand U3012 (N_3012,N_2846,N_2776);
or U3013 (N_3013,N_2939,N_2966);
and U3014 (N_3014,N_2949,N_2875);
nand U3015 (N_3015,N_2768,N_2962);
xnor U3016 (N_3016,N_2866,N_2912);
or U3017 (N_3017,N_2934,N_2946);
or U3018 (N_3018,N_2970,N_2983);
or U3019 (N_3019,N_2930,N_2992);
and U3020 (N_3020,N_2877,N_2938);
nand U3021 (N_3021,N_2861,N_2818);
xnor U3022 (N_3022,N_2863,N_2885);
xor U3023 (N_3023,N_2780,N_2799);
nand U3024 (N_3024,N_2829,N_2919);
or U3025 (N_3025,N_2926,N_2917);
nor U3026 (N_3026,N_2835,N_2880);
and U3027 (N_3027,N_2883,N_2920);
nor U3028 (N_3028,N_2820,N_2801);
and U3029 (N_3029,N_2759,N_2986);
and U3030 (N_3030,N_2900,N_2810);
and U3031 (N_3031,N_2763,N_2839);
xor U3032 (N_3032,N_2832,N_2967);
or U3033 (N_3033,N_2855,N_2947);
and U3034 (N_3034,N_2760,N_2961);
and U3035 (N_3035,N_2753,N_2813);
and U3036 (N_3036,N_2836,N_2795);
or U3037 (N_3037,N_2867,N_2936);
nand U3038 (N_3038,N_2815,N_2797);
and U3039 (N_3039,N_2881,N_2860);
nor U3040 (N_3040,N_2789,N_2940);
and U3041 (N_3041,N_2879,N_2808);
nand U3042 (N_3042,N_2889,N_2796);
nand U3043 (N_3043,N_2887,N_2911);
xnor U3044 (N_3044,N_2847,N_2972);
xor U3045 (N_3045,N_2784,N_2859);
and U3046 (N_3046,N_2843,N_2850);
or U3047 (N_3047,N_2809,N_2905);
xor U3048 (N_3048,N_2996,N_2841);
nor U3049 (N_3049,N_2886,N_2980);
nor U3050 (N_3050,N_2893,N_2876);
xor U3051 (N_3051,N_2908,N_2869);
nand U3052 (N_3052,N_2770,N_2909);
nor U3053 (N_3053,N_2952,N_2800);
xnor U3054 (N_3054,N_2901,N_2791);
nand U3055 (N_3055,N_2817,N_2769);
or U3056 (N_3056,N_2807,N_2772);
xor U3057 (N_3057,N_2811,N_2971);
or U3058 (N_3058,N_2982,N_2907);
nor U3059 (N_3059,N_2994,N_2787);
and U3060 (N_3060,N_2812,N_2872);
and U3061 (N_3061,N_2805,N_2977);
nand U3062 (N_3062,N_2782,N_2774);
nand U3063 (N_3063,N_2884,N_2822);
and U3064 (N_3064,N_2969,N_2775);
or U3065 (N_3065,N_2948,N_2981);
or U3066 (N_3066,N_2935,N_2874);
xnor U3067 (N_3067,N_2845,N_2921);
nand U3068 (N_3068,N_2899,N_2823);
xor U3069 (N_3069,N_2762,N_2798);
or U3070 (N_3070,N_2894,N_2906);
or U3071 (N_3071,N_2932,N_2904);
xnor U3072 (N_3072,N_2828,N_2840);
and U3073 (N_3073,N_2959,N_2993);
or U3074 (N_3074,N_2975,N_2816);
and U3075 (N_3075,N_2895,N_2924);
nand U3076 (N_3076,N_2802,N_2771);
xor U3077 (N_3077,N_2913,N_2945);
xor U3078 (N_3078,N_2790,N_2755);
nor U3079 (N_3079,N_2892,N_2778);
and U3080 (N_3080,N_2852,N_2960);
xor U3081 (N_3081,N_2777,N_2976);
or U3082 (N_3082,N_2825,N_2856);
nand U3083 (N_3083,N_2773,N_2923);
nor U3084 (N_3084,N_2752,N_2918);
nand U3085 (N_3085,N_2849,N_2765);
nand U3086 (N_3086,N_2833,N_2995);
nor U3087 (N_3087,N_2793,N_2956);
or U3088 (N_3088,N_2830,N_2814);
nor U3089 (N_3089,N_2827,N_2984);
or U3090 (N_3090,N_2803,N_2857);
and U3091 (N_3091,N_2950,N_2826);
nand U3092 (N_3092,N_2871,N_2751);
or U3093 (N_3093,N_2758,N_2794);
nand U3094 (N_3094,N_2868,N_2862);
or U3095 (N_3095,N_2933,N_2985);
and U3096 (N_3096,N_2989,N_2987);
nand U3097 (N_3097,N_2888,N_2974);
or U3098 (N_3098,N_2999,N_2767);
xnor U3099 (N_3099,N_2953,N_2873);
nand U3100 (N_3100,N_2954,N_2757);
nor U3101 (N_3101,N_2898,N_2882);
xnor U3102 (N_3102,N_2754,N_2837);
and U3103 (N_3103,N_2979,N_2944);
or U3104 (N_3104,N_2788,N_2858);
and U3105 (N_3105,N_2831,N_2941);
and U3106 (N_3106,N_2781,N_2865);
and U3107 (N_3107,N_2854,N_2942);
xor U3108 (N_3108,N_2834,N_2973);
nor U3109 (N_3109,N_2991,N_2931);
nand U3110 (N_3110,N_2943,N_2792);
nand U3111 (N_3111,N_2965,N_2951);
xor U3112 (N_3112,N_2957,N_2964);
nand U3113 (N_3113,N_2968,N_2963);
and U3114 (N_3114,N_2853,N_2806);
nor U3115 (N_3115,N_2870,N_2914);
and U3116 (N_3116,N_2978,N_2766);
nand U3117 (N_3117,N_2988,N_2998);
and U3118 (N_3118,N_2878,N_2848);
or U3119 (N_3119,N_2786,N_2779);
nand U3120 (N_3120,N_2890,N_2896);
nand U3121 (N_3121,N_2915,N_2997);
or U3122 (N_3122,N_2990,N_2910);
nand U3123 (N_3123,N_2761,N_2821);
nor U3124 (N_3124,N_2864,N_2937);
nor U3125 (N_3125,N_2948,N_2888);
xor U3126 (N_3126,N_2759,N_2857);
or U3127 (N_3127,N_2945,N_2886);
nand U3128 (N_3128,N_2757,N_2755);
or U3129 (N_3129,N_2752,N_2886);
nor U3130 (N_3130,N_2775,N_2955);
nor U3131 (N_3131,N_2948,N_2999);
nor U3132 (N_3132,N_2936,N_2861);
or U3133 (N_3133,N_2952,N_2821);
or U3134 (N_3134,N_2995,N_2875);
and U3135 (N_3135,N_2881,N_2857);
nor U3136 (N_3136,N_2917,N_2817);
nor U3137 (N_3137,N_2836,N_2762);
nor U3138 (N_3138,N_2835,N_2762);
xnor U3139 (N_3139,N_2751,N_2804);
and U3140 (N_3140,N_2934,N_2844);
or U3141 (N_3141,N_2769,N_2870);
xnor U3142 (N_3142,N_2997,N_2998);
nand U3143 (N_3143,N_2777,N_2943);
nand U3144 (N_3144,N_2863,N_2844);
or U3145 (N_3145,N_2795,N_2934);
nor U3146 (N_3146,N_2818,N_2874);
xnor U3147 (N_3147,N_2786,N_2941);
or U3148 (N_3148,N_2900,N_2797);
xor U3149 (N_3149,N_2812,N_2818);
xnor U3150 (N_3150,N_2921,N_2806);
xor U3151 (N_3151,N_2992,N_2818);
nand U3152 (N_3152,N_2788,N_2812);
or U3153 (N_3153,N_2942,N_2765);
and U3154 (N_3154,N_2832,N_2798);
or U3155 (N_3155,N_2923,N_2786);
nor U3156 (N_3156,N_2987,N_2967);
and U3157 (N_3157,N_2750,N_2948);
or U3158 (N_3158,N_2777,N_2922);
nand U3159 (N_3159,N_2920,N_2922);
and U3160 (N_3160,N_2886,N_2844);
or U3161 (N_3161,N_2944,N_2763);
and U3162 (N_3162,N_2869,N_2794);
or U3163 (N_3163,N_2869,N_2967);
and U3164 (N_3164,N_2771,N_2944);
nand U3165 (N_3165,N_2816,N_2787);
or U3166 (N_3166,N_2870,N_2834);
and U3167 (N_3167,N_2874,N_2793);
nand U3168 (N_3168,N_2871,N_2925);
nand U3169 (N_3169,N_2831,N_2814);
xnor U3170 (N_3170,N_2836,N_2928);
and U3171 (N_3171,N_2892,N_2931);
and U3172 (N_3172,N_2948,N_2772);
nor U3173 (N_3173,N_2895,N_2906);
and U3174 (N_3174,N_2818,N_2934);
or U3175 (N_3175,N_2900,N_2801);
nand U3176 (N_3176,N_2884,N_2958);
nor U3177 (N_3177,N_2755,N_2931);
and U3178 (N_3178,N_2877,N_2811);
nor U3179 (N_3179,N_2764,N_2932);
nand U3180 (N_3180,N_2963,N_2900);
xor U3181 (N_3181,N_2868,N_2798);
nand U3182 (N_3182,N_2971,N_2830);
or U3183 (N_3183,N_2854,N_2943);
nand U3184 (N_3184,N_2972,N_2850);
or U3185 (N_3185,N_2930,N_2964);
nand U3186 (N_3186,N_2857,N_2970);
or U3187 (N_3187,N_2891,N_2767);
or U3188 (N_3188,N_2821,N_2771);
or U3189 (N_3189,N_2856,N_2929);
nor U3190 (N_3190,N_2758,N_2965);
or U3191 (N_3191,N_2923,N_2861);
nand U3192 (N_3192,N_2807,N_2928);
or U3193 (N_3193,N_2907,N_2891);
nand U3194 (N_3194,N_2770,N_2898);
or U3195 (N_3195,N_2963,N_2840);
or U3196 (N_3196,N_2819,N_2780);
nor U3197 (N_3197,N_2778,N_2767);
nand U3198 (N_3198,N_2970,N_2759);
and U3199 (N_3199,N_2956,N_2962);
xor U3200 (N_3200,N_2823,N_2795);
xnor U3201 (N_3201,N_2805,N_2799);
xor U3202 (N_3202,N_2806,N_2928);
nand U3203 (N_3203,N_2918,N_2823);
nor U3204 (N_3204,N_2803,N_2892);
nor U3205 (N_3205,N_2962,N_2982);
nor U3206 (N_3206,N_2989,N_2894);
nand U3207 (N_3207,N_2886,N_2925);
xnor U3208 (N_3208,N_2860,N_2872);
or U3209 (N_3209,N_2799,N_2862);
nor U3210 (N_3210,N_2793,N_2989);
and U3211 (N_3211,N_2891,N_2827);
nor U3212 (N_3212,N_2799,N_2944);
and U3213 (N_3213,N_2780,N_2945);
or U3214 (N_3214,N_2890,N_2894);
xor U3215 (N_3215,N_2850,N_2961);
nor U3216 (N_3216,N_2847,N_2845);
or U3217 (N_3217,N_2904,N_2875);
nor U3218 (N_3218,N_2989,N_2939);
nand U3219 (N_3219,N_2758,N_2987);
and U3220 (N_3220,N_2822,N_2918);
nor U3221 (N_3221,N_2812,N_2755);
or U3222 (N_3222,N_2977,N_2920);
and U3223 (N_3223,N_2847,N_2952);
nor U3224 (N_3224,N_2764,N_2796);
nand U3225 (N_3225,N_2778,N_2815);
nor U3226 (N_3226,N_2816,N_2938);
nand U3227 (N_3227,N_2872,N_2849);
nand U3228 (N_3228,N_2909,N_2941);
and U3229 (N_3229,N_2760,N_2854);
nor U3230 (N_3230,N_2938,N_2770);
and U3231 (N_3231,N_2778,N_2965);
nor U3232 (N_3232,N_2817,N_2915);
nand U3233 (N_3233,N_2989,N_2992);
or U3234 (N_3234,N_2914,N_2973);
or U3235 (N_3235,N_2940,N_2865);
nand U3236 (N_3236,N_2752,N_2962);
xnor U3237 (N_3237,N_2913,N_2848);
nor U3238 (N_3238,N_2793,N_2934);
or U3239 (N_3239,N_2767,N_2994);
nand U3240 (N_3240,N_2788,N_2888);
and U3241 (N_3241,N_2767,N_2785);
or U3242 (N_3242,N_2878,N_2849);
nor U3243 (N_3243,N_2824,N_2839);
xnor U3244 (N_3244,N_2854,N_2753);
nand U3245 (N_3245,N_2938,N_2990);
nand U3246 (N_3246,N_2867,N_2828);
and U3247 (N_3247,N_2819,N_2926);
nor U3248 (N_3248,N_2889,N_2791);
or U3249 (N_3249,N_2892,N_2857);
and U3250 (N_3250,N_3026,N_3099);
xor U3251 (N_3251,N_3045,N_3184);
nand U3252 (N_3252,N_3205,N_3089);
and U3253 (N_3253,N_3206,N_3009);
nor U3254 (N_3254,N_3209,N_3004);
nor U3255 (N_3255,N_3081,N_3215);
xor U3256 (N_3256,N_3113,N_3238);
xor U3257 (N_3257,N_3028,N_3049);
or U3258 (N_3258,N_3104,N_3021);
and U3259 (N_3259,N_3218,N_3135);
nor U3260 (N_3260,N_3235,N_3106);
and U3261 (N_3261,N_3208,N_3245);
nor U3262 (N_3262,N_3037,N_3114);
and U3263 (N_3263,N_3175,N_3234);
xor U3264 (N_3264,N_3074,N_3112);
and U3265 (N_3265,N_3051,N_3195);
xor U3266 (N_3266,N_3212,N_3229);
and U3267 (N_3267,N_3171,N_3164);
and U3268 (N_3268,N_3039,N_3061);
or U3269 (N_3269,N_3134,N_3139);
nand U3270 (N_3270,N_3115,N_3240);
xor U3271 (N_3271,N_3010,N_3050);
nor U3272 (N_3272,N_3202,N_3200);
nand U3273 (N_3273,N_3147,N_3188);
nand U3274 (N_3274,N_3015,N_3110);
or U3275 (N_3275,N_3176,N_3179);
nand U3276 (N_3276,N_3043,N_3020);
and U3277 (N_3277,N_3146,N_3246);
and U3278 (N_3278,N_3007,N_3152);
nand U3279 (N_3279,N_3199,N_3192);
xor U3280 (N_3280,N_3148,N_3088);
or U3281 (N_3281,N_3228,N_3062);
and U3282 (N_3282,N_3125,N_3243);
nor U3283 (N_3283,N_3000,N_3249);
nor U3284 (N_3284,N_3082,N_3219);
and U3285 (N_3285,N_3029,N_3083);
or U3286 (N_3286,N_3034,N_3076);
or U3287 (N_3287,N_3239,N_3144);
or U3288 (N_3288,N_3017,N_3014);
nor U3289 (N_3289,N_3136,N_3003);
xnor U3290 (N_3290,N_3181,N_3221);
or U3291 (N_3291,N_3057,N_3097);
and U3292 (N_3292,N_3047,N_3191);
nor U3293 (N_3293,N_3203,N_3172);
xor U3294 (N_3294,N_3001,N_3040);
nor U3295 (N_3295,N_3052,N_3085);
or U3296 (N_3296,N_3197,N_3054);
or U3297 (N_3297,N_3071,N_3130);
nor U3298 (N_3298,N_3207,N_3162);
xor U3299 (N_3299,N_3247,N_3072);
or U3300 (N_3300,N_3117,N_3189);
nand U3301 (N_3301,N_3158,N_3137);
nor U3302 (N_3302,N_3101,N_3143);
nand U3303 (N_3303,N_3065,N_3103);
and U3304 (N_3304,N_3060,N_3183);
nor U3305 (N_3305,N_3160,N_3180);
nor U3306 (N_3306,N_3107,N_3226);
and U3307 (N_3307,N_3133,N_3005);
nor U3308 (N_3308,N_3236,N_3035);
nand U3309 (N_3309,N_3220,N_3036);
or U3310 (N_3310,N_3124,N_3210);
nand U3311 (N_3311,N_3173,N_3031);
xor U3312 (N_3312,N_3166,N_3230);
and U3313 (N_3313,N_3190,N_3223);
and U3314 (N_3314,N_3041,N_3132);
xnor U3315 (N_3315,N_3157,N_3098);
xnor U3316 (N_3316,N_3193,N_3163);
and U3317 (N_3317,N_3033,N_3142);
or U3318 (N_3318,N_3067,N_3093);
nand U3319 (N_3319,N_3012,N_3027);
or U3320 (N_3320,N_3138,N_3170);
and U3321 (N_3321,N_3187,N_3080);
xor U3322 (N_3322,N_3156,N_3100);
nand U3323 (N_3323,N_3056,N_3222);
and U3324 (N_3324,N_3087,N_3016);
and U3325 (N_3325,N_3237,N_3201);
xor U3326 (N_3326,N_3129,N_3079);
or U3327 (N_3327,N_3120,N_3108);
xor U3328 (N_3328,N_3102,N_3070);
xnor U3329 (N_3329,N_3248,N_3008);
and U3330 (N_3330,N_3042,N_3032);
or U3331 (N_3331,N_3167,N_3105);
or U3332 (N_3332,N_3055,N_3213);
xnor U3333 (N_3333,N_3128,N_3151);
nand U3334 (N_3334,N_3002,N_3058);
nor U3335 (N_3335,N_3121,N_3019);
xor U3336 (N_3336,N_3118,N_3046);
nand U3337 (N_3337,N_3169,N_3231);
xor U3338 (N_3338,N_3196,N_3145);
and U3339 (N_3339,N_3168,N_3069);
nor U3340 (N_3340,N_3214,N_3059);
and U3341 (N_3341,N_3211,N_3217);
xor U3342 (N_3342,N_3116,N_3140);
xnor U3343 (N_3343,N_3177,N_3178);
nand U3344 (N_3344,N_3078,N_3077);
and U3345 (N_3345,N_3091,N_3024);
or U3346 (N_3346,N_3242,N_3241);
or U3347 (N_3347,N_3090,N_3244);
nand U3348 (N_3348,N_3066,N_3025);
and U3349 (N_3349,N_3053,N_3194);
nor U3350 (N_3350,N_3084,N_3204);
nand U3351 (N_3351,N_3063,N_3122);
and U3352 (N_3352,N_3232,N_3131);
or U3353 (N_3353,N_3216,N_3038);
nor U3354 (N_3354,N_3182,N_3198);
or U3355 (N_3355,N_3094,N_3155);
or U3356 (N_3356,N_3044,N_3123);
and U3357 (N_3357,N_3233,N_3225);
nand U3358 (N_3358,N_3068,N_3159);
nand U3359 (N_3359,N_3006,N_3224);
nand U3360 (N_3360,N_3064,N_3073);
or U3361 (N_3361,N_3186,N_3092);
nand U3362 (N_3362,N_3119,N_3227);
nor U3363 (N_3363,N_3023,N_3165);
and U3364 (N_3364,N_3048,N_3096);
nand U3365 (N_3365,N_3185,N_3011);
and U3366 (N_3366,N_3126,N_3153);
nand U3367 (N_3367,N_3174,N_3022);
xor U3368 (N_3368,N_3127,N_3013);
or U3369 (N_3369,N_3149,N_3018);
and U3370 (N_3370,N_3095,N_3154);
xor U3371 (N_3371,N_3075,N_3086);
nand U3372 (N_3372,N_3150,N_3030);
nor U3373 (N_3373,N_3161,N_3109);
xor U3374 (N_3374,N_3111,N_3141);
and U3375 (N_3375,N_3009,N_3130);
nor U3376 (N_3376,N_3133,N_3177);
or U3377 (N_3377,N_3167,N_3026);
nor U3378 (N_3378,N_3048,N_3013);
and U3379 (N_3379,N_3149,N_3240);
or U3380 (N_3380,N_3153,N_3171);
and U3381 (N_3381,N_3219,N_3026);
nor U3382 (N_3382,N_3199,N_3220);
and U3383 (N_3383,N_3066,N_3016);
nor U3384 (N_3384,N_3070,N_3219);
nor U3385 (N_3385,N_3077,N_3127);
nor U3386 (N_3386,N_3189,N_3174);
nor U3387 (N_3387,N_3223,N_3138);
nand U3388 (N_3388,N_3106,N_3054);
nand U3389 (N_3389,N_3189,N_3098);
nor U3390 (N_3390,N_3057,N_3060);
and U3391 (N_3391,N_3224,N_3197);
or U3392 (N_3392,N_3009,N_3072);
nor U3393 (N_3393,N_3002,N_3197);
nand U3394 (N_3394,N_3189,N_3157);
and U3395 (N_3395,N_3185,N_3024);
nand U3396 (N_3396,N_3191,N_3105);
xor U3397 (N_3397,N_3040,N_3187);
and U3398 (N_3398,N_3021,N_3170);
nor U3399 (N_3399,N_3013,N_3152);
xor U3400 (N_3400,N_3170,N_3207);
nor U3401 (N_3401,N_3249,N_3043);
and U3402 (N_3402,N_3247,N_3154);
nand U3403 (N_3403,N_3049,N_3003);
nor U3404 (N_3404,N_3019,N_3007);
nand U3405 (N_3405,N_3023,N_3035);
or U3406 (N_3406,N_3010,N_3198);
or U3407 (N_3407,N_3109,N_3108);
xnor U3408 (N_3408,N_3088,N_3090);
and U3409 (N_3409,N_3229,N_3163);
or U3410 (N_3410,N_3007,N_3055);
nor U3411 (N_3411,N_3033,N_3173);
or U3412 (N_3412,N_3028,N_3226);
or U3413 (N_3413,N_3230,N_3014);
nand U3414 (N_3414,N_3104,N_3138);
nor U3415 (N_3415,N_3016,N_3169);
xnor U3416 (N_3416,N_3243,N_3132);
nand U3417 (N_3417,N_3228,N_3242);
nand U3418 (N_3418,N_3026,N_3111);
and U3419 (N_3419,N_3027,N_3193);
or U3420 (N_3420,N_3233,N_3162);
or U3421 (N_3421,N_3037,N_3160);
xor U3422 (N_3422,N_3117,N_3127);
xor U3423 (N_3423,N_3162,N_3156);
nor U3424 (N_3424,N_3109,N_3142);
nor U3425 (N_3425,N_3188,N_3166);
nor U3426 (N_3426,N_3128,N_3129);
and U3427 (N_3427,N_3170,N_3180);
and U3428 (N_3428,N_3211,N_3075);
nor U3429 (N_3429,N_3144,N_3236);
nor U3430 (N_3430,N_3107,N_3219);
nand U3431 (N_3431,N_3038,N_3203);
or U3432 (N_3432,N_3206,N_3124);
xor U3433 (N_3433,N_3058,N_3201);
nor U3434 (N_3434,N_3239,N_3057);
nand U3435 (N_3435,N_3186,N_3074);
xor U3436 (N_3436,N_3118,N_3042);
nor U3437 (N_3437,N_3167,N_3226);
nor U3438 (N_3438,N_3100,N_3025);
nand U3439 (N_3439,N_3081,N_3073);
and U3440 (N_3440,N_3209,N_3147);
xor U3441 (N_3441,N_3078,N_3005);
xor U3442 (N_3442,N_3196,N_3105);
nand U3443 (N_3443,N_3009,N_3035);
and U3444 (N_3444,N_3201,N_3216);
nor U3445 (N_3445,N_3107,N_3098);
xor U3446 (N_3446,N_3249,N_3114);
nand U3447 (N_3447,N_3123,N_3087);
or U3448 (N_3448,N_3115,N_3134);
nand U3449 (N_3449,N_3209,N_3080);
and U3450 (N_3450,N_3046,N_3088);
or U3451 (N_3451,N_3178,N_3117);
nand U3452 (N_3452,N_3060,N_3219);
or U3453 (N_3453,N_3091,N_3153);
xor U3454 (N_3454,N_3077,N_3167);
and U3455 (N_3455,N_3097,N_3091);
or U3456 (N_3456,N_3190,N_3210);
nand U3457 (N_3457,N_3007,N_3081);
nor U3458 (N_3458,N_3107,N_3000);
nor U3459 (N_3459,N_3117,N_3062);
and U3460 (N_3460,N_3112,N_3167);
nand U3461 (N_3461,N_3171,N_3040);
nand U3462 (N_3462,N_3236,N_3061);
nand U3463 (N_3463,N_3198,N_3185);
nor U3464 (N_3464,N_3218,N_3061);
or U3465 (N_3465,N_3171,N_3147);
nor U3466 (N_3466,N_3178,N_3181);
and U3467 (N_3467,N_3179,N_3100);
and U3468 (N_3468,N_3030,N_3134);
nor U3469 (N_3469,N_3207,N_3244);
xnor U3470 (N_3470,N_3061,N_3105);
or U3471 (N_3471,N_3201,N_3100);
nand U3472 (N_3472,N_3188,N_3193);
nor U3473 (N_3473,N_3075,N_3008);
or U3474 (N_3474,N_3196,N_3224);
nor U3475 (N_3475,N_3138,N_3221);
nor U3476 (N_3476,N_3097,N_3147);
or U3477 (N_3477,N_3158,N_3149);
and U3478 (N_3478,N_3157,N_3198);
or U3479 (N_3479,N_3177,N_3150);
and U3480 (N_3480,N_3062,N_3104);
nor U3481 (N_3481,N_3121,N_3074);
and U3482 (N_3482,N_3144,N_3046);
and U3483 (N_3483,N_3104,N_3246);
nor U3484 (N_3484,N_3087,N_3078);
nor U3485 (N_3485,N_3084,N_3159);
nor U3486 (N_3486,N_3093,N_3122);
or U3487 (N_3487,N_3201,N_3202);
xor U3488 (N_3488,N_3112,N_3062);
and U3489 (N_3489,N_3010,N_3221);
and U3490 (N_3490,N_3149,N_3133);
nor U3491 (N_3491,N_3195,N_3111);
xor U3492 (N_3492,N_3235,N_3125);
nor U3493 (N_3493,N_3033,N_3221);
or U3494 (N_3494,N_3069,N_3140);
or U3495 (N_3495,N_3181,N_3186);
nand U3496 (N_3496,N_3153,N_3116);
nand U3497 (N_3497,N_3099,N_3014);
or U3498 (N_3498,N_3002,N_3085);
or U3499 (N_3499,N_3172,N_3052);
xor U3500 (N_3500,N_3468,N_3370);
or U3501 (N_3501,N_3402,N_3451);
nand U3502 (N_3502,N_3265,N_3405);
and U3503 (N_3503,N_3272,N_3258);
nand U3504 (N_3504,N_3274,N_3276);
nor U3505 (N_3505,N_3484,N_3385);
and U3506 (N_3506,N_3374,N_3356);
xnor U3507 (N_3507,N_3462,N_3477);
or U3508 (N_3508,N_3382,N_3347);
or U3509 (N_3509,N_3263,N_3409);
or U3510 (N_3510,N_3419,N_3390);
or U3511 (N_3511,N_3415,N_3262);
nand U3512 (N_3512,N_3278,N_3449);
and U3513 (N_3513,N_3345,N_3496);
and U3514 (N_3514,N_3487,N_3352);
xnor U3515 (N_3515,N_3351,N_3342);
or U3516 (N_3516,N_3434,N_3321);
or U3517 (N_3517,N_3346,N_3304);
nor U3518 (N_3518,N_3309,N_3421);
or U3519 (N_3519,N_3270,N_3268);
nor U3520 (N_3520,N_3311,N_3429);
and U3521 (N_3521,N_3377,N_3306);
xnor U3522 (N_3522,N_3366,N_3320);
or U3523 (N_3523,N_3373,N_3250);
nor U3524 (N_3524,N_3478,N_3394);
or U3525 (N_3525,N_3444,N_3488);
nand U3526 (N_3526,N_3287,N_3474);
xnor U3527 (N_3527,N_3343,N_3425);
nor U3528 (N_3528,N_3357,N_3486);
nor U3529 (N_3529,N_3294,N_3411);
and U3530 (N_3530,N_3453,N_3393);
and U3531 (N_3531,N_3387,N_3456);
nand U3532 (N_3532,N_3330,N_3426);
xnor U3533 (N_3533,N_3349,N_3441);
or U3534 (N_3534,N_3446,N_3310);
or U3535 (N_3535,N_3398,N_3432);
and U3536 (N_3536,N_3372,N_3489);
xor U3537 (N_3537,N_3261,N_3283);
nand U3538 (N_3538,N_3457,N_3327);
nor U3539 (N_3539,N_3285,N_3436);
or U3540 (N_3540,N_3334,N_3410);
xor U3541 (N_3541,N_3469,N_3348);
nor U3542 (N_3542,N_3389,N_3465);
nand U3543 (N_3543,N_3273,N_3483);
xnor U3544 (N_3544,N_3433,N_3323);
xnor U3545 (N_3545,N_3470,N_3472);
or U3546 (N_3546,N_3255,N_3286);
nand U3547 (N_3547,N_3401,N_3460);
xnor U3548 (N_3548,N_3361,N_3363);
nor U3549 (N_3549,N_3297,N_3284);
nand U3550 (N_3550,N_3467,N_3404);
and U3551 (N_3551,N_3439,N_3466);
xnor U3552 (N_3552,N_3368,N_3391);
xnor U3553 (N_3553,N_3424,N_3314);
nor U3554 (N_3554,N_3379,N_3403);
xor U3555 (N_3555,N_3480,N_3397);
and U3556 (N_3556,N_3281,N_3371);
nor U3557 (N_3557,N_3471,N_3452);
nor U3558 (N_3558,N_3289,N_3337);
nand U3559 (N_3559,N_3406,N_3445);
nor U3560 (N_3560,N_3340,N_3454);
or U3561 (N_3561,N_3443,N_3288);
nand U3562 (N_3562,N_3481,N_3338);
and U3563 (N_3563,N_3324,N_3302);
or U3564 (N_3564,N_3447,N_3279);
and U3565 (N_3565,N_3494,N_3450);
or U3566 (N_3566,N_3335,N_3365);
xor U3567 (N_3567,N_3380,N_3414);
nand U3568 (N_3568,N_3305,N_3381);
nor U3569 (N_3569,N_3359,N_3252);
and U3570 (N_3570,N_3333,N_3355);
and U3571 (N_3571,N_3328,N_3317);
xnor U3572 (N_3572,N_3388,N_3339);
and U3573 (N_3573,N_3308,N_3437);
and U3574 (N_3574,N_3269,N_3296);
or U3575 (N_3575,N_3458,N_3497);
nand U3576 (N_3576,N_3384,N_3275);
nor U3577 (N_3577,N_3461,N_3256);
or U3578 (N_3578,N_3266,N_3319);
and U3579 (N_3579,N_3300,N_3399);
nand U3580 (N_3580,N_3251,N_3463);
nor U3581 (N_3581,N_3264,N_3325);
or U3582 (N_3582,N_3259,N_3312);
xor U3583 (N_3583,N_3495,N_3428);
nand U3584 (N_3584,N_3464,N_3490);
nor U3585 (N_3585,N_3376,N_3291);
xor U3586 (N_3586,N_3344,N_3400);
or U3587 (N_3587,N_3491,N_3440);
nor U3588 (N_3588,N_3431,N_3407);
nand U3589 (N_3589,N_3260,N_3271);
and U3590 (N_3590,N_3492,N_3354);
xnor U3591 (N_3591,N_3331,N_3367);
nand U3592 (N_3592,N_3313,N_3423);
or U3593 (N_3593,N_3299,N_3257);
nor U3594 (N_3594,N_3448,N_3375);
or U3595 (N_3595,N_3318,N_3482);
and U3596 (N_3596,N_3413,N_3280);
or U3597 (N_3597,N_3358,N_3475);
nor U3598 (N_3598,N_3326,N_3369);
and U3599 (N_3599,N_3316,N_3290);
nand U3600 (N_3600,N_3303,N_3418);
nor U3601 (N_3601,N_3430,N_3267);
and U3602 (N_3602,N_3329,N_3455);
xnor U3603 (N_3603,N_3417,N_3473);
nor U3604 (N_3604,N_3416,N_3499);
nand U3605 (N_3605,N_3301,N_3293);
xnor U3606 (N_3606,N_3395,N_3485);
or U3607 (N_3607,N_3493,N_3383);
xor U3608 (N_3608,N_3353,N_3362);
nor U3609 (N_3609,N_3254,N_3442);
or U3610 (N_3610,N_3498,N_3412);
xor U3611 (N_3611,N_3476,N_3341);
and U3612 (N_3612,N_3350,N_3427);
or U3613 (N_3613,N_3459,N_3435);
xnor U3614 (N_3614,N_3332,N_3292);
and U3615 (N_3615,N_3277,N_3386);
or U3616 (N_3616,N_3298,N_3253);
nand U3617 (N_3617,N_3322,N_3378);
nand U3618 (N_3618,N_3360,N_3479);
and U3619 (N_3619,N_3422,N_3315);
or U3620 (N_3620,N_3295,N_3307);
nand U3621 (N_3621,N_3408,N_3282);
and U3622 (N_3622,N_3438,N_3420);
and U3623 (N_3623,N_3392,N_3336);
and U3624 (N_3624,N_3396,N_3364);
nand U3625 (N_3625,N_3289,N_3342);
or U3626 (N_3626,N_3348,N_3467);
and U3627 (N_3627,N_3359,N_3269);
or U3628 (N_3628,N_3408,N_3323);
nand U3629 (N_3629,N_3317,N_3344);
and U3630 (N_3630,N_3367,N_3349);
and U3631 (N_3631,N_3337,N_3332);
nor U3632 (N_3632,N_3401,N_3269);
nor U3633 (N_3633,N_3344,N_3390);
and U3634 (N_3634,N_3330,N_3461);
nand U3635 (N_3635,N_3369,N_3318);
and U3636 (N_3636,N_3300,N_3462);
and U3637 (N_3637,N_3468,N_3404);
nand U3638 (N_3638,N_3368,N_3310);
and U3639 (N_3639,N_3460,N_3458);
or U3640 (N_3640,N_3404,N_3438);
xor U3641 (N_3641,N_3407,N_3367);
nand U3642 (N_3642,N_3341,N_3458);
nand U3643 (N_3643,N_3396,N_3443);
or U3644 (N_3644,N_3496,N_3346);
nand U3645 (N_3645,N_3424,N_3419);
nand U3646 (N_3646,N_3389,N_3278);
xor U3647 (N_3647,N_3439,N_3368);
and U3648 (N_3648,N_3476,N_3425);
nand U3649 (N_3649,N_3431,N_3403);
and U3650 (N_3650,N_3411,N_3296);
or U3651 (N_3651,N_3420,N_3413);
and U3652 (N_3652,N_3423,N_3336);
nand U3653 (N_3653,N_3483,N_3369);
nor U3654 (N_3654,N_3461,N_3454);
nor U3655 (N_3655,N_3341,N_3390);
nor U3656 (N_3656,N_3287,N_3317);
nand U3657 (N_3657,N_3477,N_3303);
xor U3658 (N_3658,N_3421,N_3329);
or U3659 (N_3659,N_3290,N_3466);
nor U3660 (N_3660,N_3481,N_3295);
and U3661 (N_3661,N_3363,N_3265);
xor U3662 (N_3662,N_3383,N_3319);
xor U3663 (N_3663,N_3469,N_3265);
nor U3664 (N_3664,N_3263,N_3482);
and U3665 (N_3665,N_3334,N_3393);
nor U3666 (N_3666,N_3325,N_3445);
nor U3667 (N_3667,N_3474,N_3433);
and U3668 (N_3668,N_3318,N_3408);
nor U3669 (N_3669,N_3316,N_3481);
and U3670 (N_3670,N_3428,N_3262);
xnor U3671 (N_3671,N_3320,N_3456);
nand U3672 (N_3672,N_3443,N_3321);
or U3673 (N_3673,N_3251,N_3484);
nor U3674 (N_3674,N_3482,N_3392);
or U3675 (N_3675,N_3406,N_3415);
or U3676 (N_3676,N_3305,N_3398);
nor U3677 (N_3677,N_3413,N_3383);
xor U3678 (N_3678,N_3260,N_3422);
nand U3679 (N_3679,N_3364,N_3309);
xnor U3680 (N_3680,N_3456,N_3299);
nand U3681 (N_3681,N_3452,N_3318);
xnor U3682 (N_3682,N_3274,N_3446);
or U3683 (N_3683,N_3361,N_3436);
nor U3684 (N_3684,N_3486,N_3449);
xor U3685 (N_3685,N_3288,N_3390);
nor U3686 (N_3686,N_3340,N_3371);
and U3687 (N_3687,N_3287,N_3478);
nor U3688 (N_3688,N_3434,N_3494);
and U3689 (N_3689,N_3495,N_3404);
nor U3690 (N_3690,N_3420,N_3418);
nor U3691 (N_3691,N_3417,N_3387);
or U3692 (N_3692,N_3434,N_3468);
nand U3693 (N_3693,N_3271,N_3269);
and U3694 (N_3694,N_3354,N_3345);
nor U3695 (N_3695,N_3372,N_3363);
or U3696 (N_3696,N_3275,N_3334);
nand U3697 (N_3697,N_3495,N_3372);
nand U3698 (N_3698,N_3398,N_3283);
xor U3699 (N_3699,N_3353,N_3309);
nand U3700 (N_3700,N_3366,N_3387);
nor U3701 (N_3701,N_3346,N_3445);
or U3702 (N_3702,N_3445,N_3487);
nor U3703 (N_3703,N_3357,N_3315);
and U3704 (N_3704,N_3480,N_3318);
nor U3705 (N_3705,N_3266,N_3477);
and U3706 (N_3706,N_3260,N_3283);
nand U3707 (N_3707,N_3361,N_3419);
and U3708 (N_3708,N_3366,N_3431);
or U3709 (N_3709,N_3476,N_3296);
or U3710 (N_3710,N_3256,N_3408);
nor U3711 (N_3711,N_3420,N_3384);
or U3712 (N_3712,N_3254,N_3401);
or U3713 (N_3713,N_3334,N_3356);
xor U3714 (N_3714,N_3412,N_3338);
nand U3715 (N_3715,N_3430,N_3436);
xnor U3716 (N_3716,N_3339,N_3409);
nor U3717 (N_3717,N_3313,N_3253);
xor U3718 (N_3718,N_3481,N_3306);
or U3719 (N_3719,N_3445,N_3301);
and U3720 (N_3720,N_3359,N_3426);
nand U3721 (N_3721,N_3315,N_3355);
nand U3722 (N_3722,N_3274,N_3389);
or U3723 (N_3723,N_3359,N_3295);
xor U3724 (N_3724,N_3401,N_3438);
xor U3725 (N_3725,N_3474,N_3285);
nand U3726 (N_3726,N_3489,N_3353);
nand U3727 (N_3727,N_3340,N_3326);
or U3728 (N_3728,N_3482,N_3354);
or U3729 (N_3729,N_3384,N_3496);
nand U3730 (N_3730,N_3411,N_3450);
nand U3731 (N_3731,N_3361,N_3250);
xnor U3732 (N_3732,N_3382,N_3397);
nor U3733 (N_3733,N_3460,N_3306);
xor U3734 (N_3734,N_3403,N_3418);
and U3735 (N_3735,N_3361,N_3309);
and U3736 (N_3736,N_3369,N_3333);
and U3737 (N_3737,N_3403,N_3451);
and U3738 (N_3738,N_3294,N_3337);
nand U3739 (N_3739,N_3258,N_3354);
and U3740 (N_3740,N_3498,N_3433);
xor U3741 (N_3741,N_3456,N_3310);
nor U3742 (N_3742,N_3284,N_3430);
and U3743 (N_3743,N_3306,N_3401);
or U3744 (N_3744,N_3252,N_3290);
and U3745 (N_3745,N_3321,N_3468);
and U3746 (N_3746,N_3456,N_3265);
nor U3747 (N_3747,N_3372,N_3380);
and U3748 (N_3748,N_3461,N_3485);
and U3749 (N_3749,N_3459,N_3328);
xnor U3750 (N_3750,N_3668,N_3697);
or U3751 (N_3751,N_3733,N_3615);
xnor U3752 (N_3752,N_3694,N_3557);
and U3753 (N_3753,N_3546,N_3690);
nand U3754 (N_3754,N_3587,N_3651);
or U3755 (N_3755,N_3620,N_3722);
and U3756 (N_3756,N_3539,N_3501);
or U3757 (N_3757,N_3602,N_3705);
nor U3758 (N_3758,N_3594,N_3580);
or U3759 (N_3759,N_3653,N_3682);
or U3760 (N_3760,N_3506,N_3718);
nand U3761 (N_3761,N_3563,N_3529);
xor U3762 (N_3762,N_3535,N_3635);
xor U3763 (N_3763,N_3633,N_3622);
nand U3764 (N_3764,N_3619,N_3648);
xor U3765 (N_3765,N_3736,N_3543);
and U3766 (N_3766,N_3695,N_3512);
nand U3767 (N_3767,N_3577,N_3728);
xor U3768 (N_3768,N_3661,N_3672);
and U3769 (N_3769,N_3642,N_3544);
or U3770 (N_3770,N_3646,N_3574);
nand U3771 (N_3771,N_3609,N_3688);
nor U3772 (N_3772,N_3523,N_3590);
nor U3773 (N_3773,N_3737,N_3640);
xnor U3774 (N_3774,N_3547,N_3591);
and U3775 (N_3775,N_3556,N_3745);
xor U3776 (N_3776,N_3606,N_3518);
and U3777 (N_3777,N_3680,N_3702);
and U3778 (N_3778,N_3562,N_3716);
xor U3779 (N_3779,N_3675,N_3656);
nand U3780 (N_3780,N_3638,N_3567);
or U3781 (N_3781,N_3511,N_3558);
and U3782 (N_3782,N_3516,N_3643);
and U3783 (N_3783,N_3720,N_3749);
nand U3784 (N_3784,N_3614,N_3743);
and U3785 (N_3785,N_3571,N_3739);
nor U3786 (N_3786,N_3541,N_3678);
xor U3787 (N_3787,N_3553,N_3578);
or U3788 (N_3788,N_3533,N_3502);
or U3789 (N_3789,N_3579,N_3549);
or U3790 (N_3790,N_3540,N_3669);
xor U3791 (N_3791,N_3537,N_3639);
nor U3792 (N_3792,N_3625,N_3568);
and U3793 (N_3793,N_3664,N_3589);
xnor U3794 (N_3794,N_3674,N_3679);
or U3795 (N_3795,N_3686,N_3671);
and U3796 (N_3796,N_3660,N_3700);
xnor U3797 (N_3797,N_3711,N_3505);
or U3798 (N_3798,N_3717,N_3698);
nor U3799 (N_3799,N_3631,N_3659);
or U3800 (N_3800,N_3724,N_3731);
and U3801 (N_3801,N_3644,N_3605);
or U3802 (N_3802,N_3657,N_3504);
xor U3803 (N_3803,N_3727,N_3707);
and U3804 (N_3804,N_3598,N_3572);
xor U3805 (N_3805,N_3536,N_3517);
and U3806 (N_3806,N_3624,N_3510);
nor U3807 (N_3807,N_3534,N_3706);
nor U3808 (N_3808,N_3647,N_3592);
xor U3809 (N_3809,N_3519,N_3630);
nand U3810 (N_3810,N_3515,N_3600);
nand U3811 (N_3811,N_3617,N_3673);
nand U3812 (N_3812,N_3588,N_3744);
and U3813 (N_3813,N_3611,N_3551);
nand U3814 (N_3814,N_3513,N_3601);
nor U3815 (N_3815,N_3721,N_3608);
and U3816 (N_3816,N_3650,N_3652);
nand U3817 (N_3817,N_3748,N_3564);
nand U3818 (N_3818,N_3747,N_3741);
xor U3819 (N_3819,N_3545,N_3514);
xnor U3820 (N_3820,N_3729,N_3522);
nand U3821 (N_3821,N_3641,N_3735);
nor U3822 (N_3822,N_3696,N_3616);
nor U3823 (N_3823,N_3701,N_3703);
nor U3824 (N_3824,N_3629,N_3526);
nand U3825 (N_3825,N_3654,N_3532);
and U3826 (N_3826,N_3566,N_3725);
nand U3827 (N_3827,N_3637,N_3684);
nand U3828 (N_3828,N_3655,N_3560);
nor U3829 (N_3829,N_3595,N_3584);
xor U3830 (N_3830,N_3746,N_3685);
nor U3831 (N_3831,N_3666,N_3525);
or U3832 (N_3832,N_3667,N_3508);
nand U3833 (N_3833,N_3507,N_3597);
and U3834 (N_3834,N_3708,N_3709);
and U3835 (N_3835,N_3610,N_3527);
xnor U3836 (N_3836,N_3740,N_3612);
nor U3837 (N_3837,N_3704,N_3742);
nor U3838 (N_3838,N_3734,N_3710);
xor U3839 (N_3839,N_3689,N_3604);
xnor U3840 (N_3840,N_3649,N_3663);
nand U3841 (N_3841,N_3714,N_3613);
nor U3842 (N_3842,N_3607,N_3621);
nor U3843 (N_3843,N_3554,N_3576);
nand U3844 (N_3844,N_3538,N_3683);
nand U3845 (N_3845,N_3692,N_3627);
nor U3846 (N_3846,N_3570,N_3687);
nor U3847 (N_3847,N_3712,N_3693);
xor U3848 (N_3848,N_3658,N_3573);
and U3849 (N_3849,N_3632,N_3623);
and U3850 (N_3850,N_3593,N_3503);
nand U3851 (N_3851,N_3662,N_3520);
or U3852 (N_3852,N_3521,N_3561);
nand U3853 (N_3853,N_3552,N_3575);
xor U3854 (N_3854,N_3676,N_3583);
xor U3855 (N_3855,N_3530,N_3730);
nor U3856 (N_3856,N_3582,N_3628);
nand U3857 (N_3857,N_3677,N_3738);
nor U3858 (N_3858,N_3626,N_3691);
or U3859 (N_3859,N_3665,N_3500);
and U3860 (N_3860,N_3509,N_3599);
xor U3861 (N_3861,N_3636,N_3581);
or U3862 (N_3862,N_3670,N_3645);
xnor U3863 (N_3863,N_3585,N_3550);
and U3864 (N_3864,N_3634,N_3531);
and U3865 (N_3865,N_3618,N_3723);
or U3866 (N_3866,N_3524,N_3555);
nor U3867 (N_3867,N_3719,N_3699);
and U3868 (N_3868,N_3569,N_3732);
nor U3869 (N_3869,N_3565,N_3542);
nor U3870 (N_3870,N_3548,N_3596);
and U3871 (N_3871,N_3586,N_3726);
xor U3872 (N_3872,N_3528,N_3559);
nor U3873 (N_3873,N_3603,N_3715);
nor U3874 (N_3874,N_3681,N_3713);
nor U3875 (N_3875,N_3590,N_3629);
xnor U3876 (N_3876,N_3728,N_3663);
and U3877 (N_3877,N_3551,N_3623);
xnor U3878 (N_3878,N_3741,N_3576);
or U3879 (N_3879,N_3577,N_3500);
nor U3880 (N_3880,N_3539,N_3713);
nor U3881 (N_3881,N_3664,N_3669);
nand U3882 (N_3882,N_3581,N_3544);
xnor U3883 (N_3883,N_3636,N_3532);
nor U3884 (N_3884,N_3579,N_3641);
nand U3885 (N_3885,N_3638,N_3511);
nor U3886 (N_3886,N_3663,N_3636);
nor U3887 (N_3887,N_3565,N_3655);
nand U3888 (N_3888,N_3724,N_3641);
xor U3889 (N_3889,N_3729,N_3573);
or U3890 (N_3890,N_3666,N_3733);
xor U3891 (N_3891,N_3537,N_3524);
or U3892 (N_3892,N_3640,N_3608);
or U3893 (N_3893,N_3577,N_3746);
nor U3894 (N_3894,N_3589,N_3525);
or U3895 (N_3895,N_3729,N_3564);
nand U3896 (N_3896,N_3659,N_3643);
or U3897 (N_3897,N_3564,N_3677);
and U3898 (N_3898,N_3569,N_3603);
and U3899 (N_3899,N_3505,N_3621);
and U3900 (N_3900,N_3685,N_3691);
xnor U3901 (N_3901,N_3663,N_3616);
nand U3902 (N_3902,N_3727,N_3531);
or U3903 (N_3903,N_3731,N_3568);
xor U3904 (N_3904,N_3618,N_3547);
xnor U3905 (N_3905,N_3574,N_3693);
nor U3906 (N_3906,N_3559,N_3609);
nor U3907 (N_3907,N_3570,N_3535);
and U3908 (N_3908,N_3662,N_3616);
nor U3909 (N_3909,N_3596,N_3501);
nand U3910 (N_3910,N_3648,N_3588);
xnor U3911 (N_3911,N_3746,N_3571);
and U3912 (N_3912,N_3531,N_3516);
nand U3913 (N_3913,N_3611,N_3586);
or U3914 (N_3914,N_3604,N_3727);
or U3915 (N_3915,N_3714,N_3642);
xor U3916 (N_3916,N_3580,N_3545);
nand U3917 (N_3917,N_3611,N_3719);
nand U3918 (N_3918,N_3500,N_3709);
and U3919 (N_3919,N_3604,N_3556);
nand U3920 (N_3920,N_3684,N_3625);
and U3921 (N_3921,N_3570,N_3575);
nor U3922 (N_3922,N_3674,N_3613);
nor U3923 (N_3923,N_3506,N_3510);
xnor U3924 (N_3924,N_3679,N_3563);
xor U3925 (N_3925,N_3649,N_3634);
xnor U3926 (N_3926,N_3537,N_3712);
xor U3927 (N_3927,N_3646,N_3518);
and U3928 (N_3928,N_3692,N_3508);
xnor U3929 (N_3929,N_3552,N_3623);
nor U3930 (N_3930,N_3651,N_3668);
nor U3931 (N_3931,N_3583,N_3650);
nand U3932 (N_3932,N_3630,N_3701);
and U3933 (N_3933,N_3735,N_3616);
nand U3934 (N_3934,N_3725,N_3570);
nand U3935 (N_3935,N_3732,N_3713);
or U3936 (N_3936,N_3569,N_3662);
nand U3937 (N_3937,N_3721,N_3524);
nand U3938 (N_3938,N_3689,N_3622);
or U3939 (N_3939,N_3603,N_3747);
nor U3940 (N_3940,N_3747,N_3554);
nor U3941 (N_3941,N_3517,N_3713);
nor U3942 (N_3942,N_3725,N_3731);
nand U3943 (N_3943,N_3593,N_3520);
or U3944 (N_3944,N_3616,N_3722);
nand U3945 (N_3945,N_3556,N_3714);
xor U3946 (N_3946,N_3737,N_3562);
or U3947 (N_3947,N_3648,N_3504);
xor U3948 (N_3948,N_3631,N_3680);
nand U3949 (N_3949,N_3707,N_3690);
and U3950 (N_3950,N_3602,N_3664);
nand U3951 (N_3951,N_3579,N_3537);
nand U3952 (N_3952,N_3594,N_3702);
and U3953 (N_3953,N_3606,N_3582);
nand U3954 (N_3954,N_3500,N_3677);
nor U3955 (N_3955,N_3720,N_3592);
nand U3956 (N_3956,N_3731,N_3598);
nor U3957 (N_3957,N_3676,N_3675);
xor U3958 (N_3958,N_3711,N_3640);
xor U3959 (N_3959,N_3664,N_3549);
nor U3960 (N_3960,N_3702,N_3580);
nand U3961 (N_3961,N_3553,N_3577);
and U3962 (N_3962,N_3612,N_3551);
xor U3963 (N_3963,N_3644,N_3732);
nor U3964 (N_3964,N_3647,N_3691);
nand U3965 (N_3965,N_3732,N_3584);
or U3966 (N_3966,N_3729,N_3528);
nand U3967 (N_3967,N_3598,N_3651);
and U3968 (N_3968,N_3630,N_3708);
xor U3969 (N_3969,N_3544,N_3586);
nor U3970 (N_3970,N_3575,N_3711);
nor U3971 (N_3971,N_3718,N_3735);
and U3972 (N_3972,N_3664,N_3523);
and U3973 (N_3973,N_3748,N_3608);
xnor U3974 (N_3974,N_3703,N_3659);
and U3975 (N_3975,N_3716,N_3746);
or U3976 (N_3976,N_3652,N_3629);
and U3977 (N_3977,N_3720,N_3658);
xor U3978 (N_3978,N_3714,N_3732);
xor U3979 (N_3979,N_3710,N_3549);
xor U3980 (N_3980,N_3537,N_3713);
xnor U3981 (N_3981,N_3612,N_3747);
or U3982 (N_3982,N_3668,N_3725);
nand U3983 (N_3983,N_3522,N_3573);
nand U3984 (N_3984,N_3724,N_3694);
xor U3985 (N_3985,N_3718,N_3530);
and U3986 (N_3986,N_3683,N_3551);
xnor U3987 (N_3987,N_3540,N_3526);
or U3988 (N_3988,N_3553,N_3661);
nor U3989 (N_3989,N_3732,N_3535);
nand U3990 (N_3990,N_3565,N_3506);
nand U3991 (N_3991,N_3561,N_3664);
nand U3992 (N_3992,N_3745,N_3736);
xor U3993 (N_3993,N_3532,N_3614);
and U3994 (N_3994,N_3647,N_3655);
xor U3995 (N_3995,N_3516,N_3667);
and U3996 (N_3996,N_3507,N_3659);
and U3997 (N_3997,N_3664,N_3632);
nand U3998 (N_3998,N_3567,N_3622);
or U3999 (N_3999,N_3633,N_3504);
or U4000 (N_4000,N_3803,N_3782);
or U4001 (N_4001,N_3753,N_3877);
or U4002 (N_4002,N_3791,N_3761);
nor U4003 (N_4003,N_3800,N_3994);
nor U4004 (N_4004,N_3856,N_3863);
nor U4005 (N_4005,N_3973,N_3792);
xor U4006 (N_4006,N_3845,N_3983);
nor U4007 (N_4007,N_3965,N_3799);
nor U4008 (N_4008,N_3809,N_3879);
xnor U4009 (N_4009,N_3883,N_3778);
and U4010 (N_4010,N_3843,N_3758);
or U4011 (N_4011,N_3865,N_3752);
and U4012 (N_4012,N_3933,N_3805);
nor U4013 (N_4013,N_3891,N_3899);
or U4014 (N_4014,N_3914,N_3870);
nor U4015 (N_4015,N_3854,N_3806);
or U4016 (N_4016,N_3918,N_3796);
xor U4017 (N_4017,N_3763,N_3882);
nor U4018 (N_4018,N_3884,N_3886);
and U4019 (N_4019,N_3984,N_3903);
nand U4020 (N_4020,N_3954,N_3808);
nand U4021 (N_4021,N_3779,N_3793);
nand U4022 (N_4022,N_3894,N_3975);
xnor U4023 (N_4023,N_3847,N_3757);
xor U4024 (N_4024,N_3940,N_3773);
and U4025 (N_4025,N_3876,N_3905);
and U4026 (N_4026,N_3969,N_3785);
nor U4027 (N_4027,N_3941,N_3974);
xnor U4028 (N_4028,N_3930,N_3978);
xor U4029 (N_4029,N_3935,N_3840);
nand U4030 (N_4030,N_3828,N_3985);
nand U4031 (N_4031,N_3892,N_3948);
xor U4032 (N_4032,N_3767,N_3960);
and U4033 (N_4033,N_3990,N_3772);
xor U4034 (N_4034,N_3762,N_3844);
and U4035 (N_4035,N_3780,N_3812);
or U4036 (N_4036,N_3751,N_3897);
xnor U4037 (N_4037,N_3830,N_3937);
or U4038 (N_4038,N_3966,N_3817);
or U4039 (N_4039,N_3938,N_3825);
or U4040 (N_4040,N_3916,N_3837);
and U4041 (N_4041,N_3839,N_3980);
or U4042 (N_4042,N_3853,N_3971);
and U4043 (N_4043,N_3850,N_3956);
or U4044 (N_4044,N_3928,N_3907);
xnor U4045 (N_4045,N_3864,N_3769);
xor U4046 (N_4046,N_3831,N_3991);
xnor U4047 (N_4047,N_3783,N_3926);
or U4048 (N_4048,N_3776,N_3821);
nor U4049 (N_4049,N_3898,N_3943);
and U4050 (N_4050,N_3921,N_3917);
nor U4051 (N_4051,N_3906,N_3874);
or U4052 (N_4052,N_3992,N_3888);
nor U4053 (N_4053,N_3860,N_3815);
nor U4054 (N_4054,N_3857,N_3873);
nand U4055 (N_4055,N_3922,N_3925);
or U4056 (N_4056,N_3835,N_3827);
xnor U4057 (N_4057,N_3759,N_3887);
and U4058 (N_4058,N_3764,N_3953);
xor U4059 (N_4059,N_3820,N_3775);
and U4060 (N_4060,N_3979,N_3934);
and U4061 (N_4061,N_3755,N_3816);
xor U4062 (N_4062,N_3756,N_3950);
and U4063 (N_4063,N_3833,N_3760);
xor U4064 (N_4064,N_3951,N_3871);
and U4065 (N_4065,N_3855,N_3939);
nor U4066 (N_4066,N_3836,N_3997);
and U4067 (N_4067,N_3765,N_3880);
and U4068 (N_4068,N_3927,N_3964);
and U4069 (N_4069,N_3852,N_3986);
nor U4070 (N_4070,N_3789,N_3962);
or U4071 (N_4071,N_3889,N_3910);
nand U4072 (N_4072,N_3788,N_3861);
or U4073 (N_4073,N_3895,N_3981);
xor U4074 (N_4074,N_3754,N_3790);
and U4075 (N_4075,N_3867,N_3819);
nand U4076 (N_4076,N_3849,N_3885);
xor U4077 (N_4077,N_3968,N_3848);
or U4078 (N_4078,N_3977,N_3766);
or U4079 (N_4079,N_3841,N_3900);
or U4080 (N_4080,N_3909,N_3959);
xnor U4081 (N_4081,N_3967,N_3846);
nand U4082 (N_4082,N_3915,N_3961);
nand U4083 (N_4083,N_3952,N_3822);
or U4084 (N_4084,N_3936,N_3901);
and U4085 (N_4085,N_3750,N_3929);
or U4086 (N_4086,N_3902,N_3878);
or U4087 (N_4087,N_3869,N_3798);
and U4088 (N_4088,N_3777,N_3955);
and U4089 (N_4089,N_3802,N_3813);
nor U4090 (N_4090,N_3811,N_3987);
nor U4091 (N_4091,N_3893,N_3858);
nor U4092 (N_4092,N_3784,N_3807);
nor U4093 (N_4093,N_3963,N_3770);
nand U4094 (N_4094,N_3919,N_3829);
or U4095 (N_4095,N_3768,N_3924);
nand U4096 (N_4096,N_3949,N_3972);
nand U4097 (N_4097,N_3862,N_3931);
and U4098 (N_4098,N_3787,N_3786);
nor U4099 (N_4099,N_3912,N_3794);
nor U4100 (N_4100,N_3896,N_3868);
nand U4101 (N_4101,N_3881,N_3851);
and U4102 (N_4102,N_3996,N_3911);
xnor U4103 (N_4103,N_3823,N_3946);
or U4104 (N_4104,N_3993,N_3958);
nor U4105 (N_4105,N_3947,N_3814);
xor U4106 (N_4106,N_3904,N_3989);
or U4107 (N_4107,N_3944,N_3982);
and U4108 (N_4108,N_3913,N_3801);
xnor U4109 (N_4109,N_3818,N_3872);
nand U4110 (N_4110,N_3957,N_3804);
nand U4111 (N_4111,N_3932,N_3976);
or U4112 (N_4112,N_3942,N_3866);
xnor U4113 (N_4113,N_3842,N_3832);
nand U4114 (N_4114,N_3945,N_3875);
or U4115 (N_4115,N_3781,N_3838);
and U4116 (N_4116,N_3797,N_3920);
and U4117 (N_4117,N_3824,N_3908);
nand U4118 (N_4118,N_3771,N_3795);
nor U4119 (N_4119,N_3995,N_3810);
or U4120 (N_4120,N_3890,N_3999);
nor U4121 (N_4121,N_3923,N_3859);
nor U4122 (N_4122,N_3998,N_3834);
nor U4123 (N_4123,N_3826,N_3988);
xnor U4124 (N_4124,N_3970,N_3774);
nor U4125 (N_4125,N_3906,N_3873);
or U4126 (N_4126,N_3803,N_3770);
xor U4127 (N_4127,N_3896,N_3951);
xnor U4128 (N_4128,N_3755,N_3852);
nand U4129 (N_4129,N_3991,N_3761);
xnor U4130 (N_4130,N_3978,N_3977);
or U4131 (N_4131,N_3794,N_3910);
and U4132 (N_4132,N_3851,N_3958);
or U4133 (N_4133,N_3758,N_3804);
and U4134 (N_4134,N_3944,N_3856);
and U4135 (N_4135,N_3902,N_3831);
nor U4136 (N_4136,N_3917,N_3944);
and U4137 (N_4137,N_3800,N_3910);
or U4138 (N_4138,N_3787,N_3824);
nor U4139 (N_4139,N_3837,N_3925);
nand U4140 (N_4140,N_3883,N_3888);
or U4141 (N_4141,N_3994,N_3973);
nand U4142 (N_4142,N_3858,N_3769);
and U4143 (N_4143,N_3794,N_3959);
and U4144 (N_4144,N_3977,N_3906);
and U4145 (N_4145,N_3755,N_3801);
nand U4146 (N_4146,N_3763,N_3941);
nor U4147 (N_4147,N_3904,N_3794);
or U4148 (N_4148,N_3847,N_3988);
nor U4149 (N_4149,N_3871,N_3756);
or U4150 (N_4150,N_3944,N_3840);
nand U4151 (N_4151,N_3962,N_3761);
xor U4152 (N_4152,N_3977,N_3889);
or U4153 (N_4153,N_3816,N_3752);
nand U4154 (N_4154,N_3868,N_3951);
xnor U4155 (N_4155,N_3959,N_3847);
and U4156 (N_4156,N_3828,N_3874);
and U4157 (N_4157,N_3841,N_3802);
nand U4158 (N_4158,N_3911,N_3842);
nand U4159 (N_4159,N_3927,N_3914);
or U4160 (N_4160,N_3913,N_3951);
nor U4161 (N_4161,N_3962,N_3802);
nor U4162 (N_4162,N_3983,N_3775);
and U4163 (N_4163,N_3828,N_3758);
nand U4164 (N_4164,N_3959,N_3778);
xor U4165 (N_4165,N_3943,N_3921);
xor U4166 (N_4166,N_3855,N_3967);
and U4167 (N_4167,N_3954,N_3802);
and U4168 (N_4168,N_3978,N_3848);
and U4169 (N_4169,N_3924,N_3775);
or U4170 (N_4170,N_3826,N_3940);
and U4171 (N_4171,N_3994,N_3961);
nor U4172 (N_4172,N_3974,N_3813);
nor U4173 (N_4173,N_3894,N_3783);
nand U4174 (N_4174,N_3807,N_3876);
nand U4175 (N_4175,N_3759,N_3797);
xnor U4176 (N_4176,N_3984,N_3924);
nand U4177 (N_4177,N_3784,N_3906);
or U4178 (N_4178,N_3858,N_3806);
xnor U4179 (N_4179,N_3905,N_3758);
or U4180 (N_4180,N_3795,N_3788);
or U4181 (N_4181,N_3996,N_3986);
xnor U4182 (N_4182,N_3875,N_3808);
and U4183 (N_4183,N_3987,N_3983);
nor U4184 (N_4184,N_3813,N_3896);
or U4185 (N_4185,N_3834,N_3857);
or U4186 (N_4186,N_3760,N_3876);
xnor U4187 (N_4187,N_3947,N_3940);
nand U4188 (N_4188,N_3829,N_3950);
nand U4189 (N_4189,N_3862,N_3841);
nand U4190 (N_4190,N_3955,N_3769);
and U4191 (N_4191,N_3759,N_3969);
or U4192 (N_4192,N_3870,N_3907);
nor U4193 (N_4193,N_3963,N_3947);
or U4194 (N_4194,N_3790,N_3917);
xnor U4195 (N_4195,N_3842,N_3886);
or U4196 (N_4196,N_3866,N_3839);
or U4197 (N_4197,N_3762,N_3795);
xor U4198 (N_4198,N_3750,N_3789);
nand U4199 (N_4199,N_3770,N_3968);
or U4200 (N_4200,N_3993,N_3825);
nand U4201 (N_4201,N_3831,N_3797);
nor U4202 (N_4202,N_3788,N_3797);
nor U4203 (N_4203,N_3775,N_3901);
nand U4204 (N_4204,N_3928,N_3775);
nand U4205 (N_4205,N_3800,N_3865);
and U4206 (N_4206,N_3846,N_3750);
xnor U4207 (N_4207,N_3802,N_3923);
nor U4208 (N_4208,N_3867,N_3827);
xor U4209 (N_4209,N_3761,N_3933);
nand U4210 (N_4210,N_3826,N_3836);
or U4211 (N_4211,N_3849,N_3893);
or U4212 (N_4212,N_3901,N_3890);
and U4213 (N_4213,N_3881,N_3994);
nand U4214 (N_4214,N_3788,N_3881);
nand U4215 (N_4215,N_3991,N_3785);
xor U4216 (N_4216,N_3888,N_3847);
and U4217 (N_4217,N_3757,N_3913);
and U4218 (N_4218,N_3789,N_3809);
or U4219 (N_4219,N_3999,N_3979);
or U4220 (N_4220,N_3826,N_3909);
and U4221 (N_4221,N_3863,N_3900);
or U4222 (N_4222,N_3771,N_3909);
xnor U4223 (N_4223,N_3988,N_3777);
nor U4224 (N_4224,N_3886,N_3786);
nand U4225 (N_4225,N_3936,N_3847);
and U4226 (N_4226,N_3758,N_3899);
nor U4227 (N_4227,N_3834,N_3835);
xnor U4228 (N_4228,N_3968,N_3765);
and U4229 (N_4229,N_3941,N_3833);
or U4230 (N_4230,N_3912,N_3759);
and U4231 (N_4231,N_3925,N_3995);
nor U4232 (N_4232,N_3776,N_3803);
and U4233 (N_4233,N_3807,N_3983);
nand U4234 (N_4234,N_3909,N_3818);
or U4235 (N_4235,N_3802,N_3947);
and U4236 (N_4236,N_3823,N_3760);
xnor U4237 (N_4237,N_3798,N_3977);
nand U4238 (N_4238,N_3814,N_3892);
and U4239 (N_4239,N_3944,N_3832);
nor U4240 (N_4240,N_3825,N_3875);
nor U4241 (N_4241,N_3908,N_3782);
or U4242 (N_4242,N_3958,N_3840);
nand U4243 (N_4243,N_3778,N_3750);
xor U4244 (N_4244,N_3812,N_3966);
nor U4245 (N_4245,N_3963,N_3932);
or U4246 (N_4246,N_3909,N_3807);
and U4247 (N_4247,N_3794,N_3759);
nand U4248 (N_4248,N_3947,N_3842);
and U4249 (N_4249,N_3833,N_3956);
nor U4250 (N_4250,N_4028,N_4173);
or U4251 (N_4251,N_4248,N_4197);
xor U4252 (N_4252,N_4154,N_4126);
and U4253 (N_4253,N_4039,N_4165);
or U4254 (N_4254,N_4218,N_4073);
xor U4255 (N_4255,N_4058,N_4199);
xor U4256 (N_4256,N_4157,N_4018);
or U4257 (N_4257,N_4053,N_4227);
nor U4258 (N_4258,N_4177,N_4042);
nand U4259 (N_4259,N_4066,N_4044);
nand U4260 (N_4260,N_4205,N_4178);
or U4261 (N_4261,N_4062,N_4155);
nand U4262 (N_4262,N_4182,N_4083);
nand U4263 (N_4263,N_4085,N_4204);
or U4264 (N_4264,N_4040,N_4070);
xor U4265 (N_4265,N_4153,N_4242);
or U4266 (N_4266,N_4210,N_4176);
nand U4267 (N_4267,N_4110,N_4017);
or U4268 (N_4268,N_4184,N_4198);
xor U4269 (N_4269,N_4164,N_4240);
or U4270 (N_4270,N_4136,N_4012);
and U4271 (N_4271,N_4160,N_4234);
nor U4272 (N_4272,N_4159,N_4119);
and U4273 (N_4273,N_4245,N_4180);
nand U4274 (N_4274,N_4052,N_4141);
nor U4275 (N_4275,N_4191,N_4166);
or U4276 (N_4276,N_4175,N_4217);
xnor U4277 (N_4277,N_4172,N_4023);
nand U4278 (N_4278,N_4093,N_4125);
nand U4279 (N_4279,N_4214,N_4121);
or U4280 (N_4280,N_4067,N_4002);
and U4281 (N_4281,N_4026,N_4037);
or U4282 (N_4282,N_4082,N_4022);
and U4283 (N_4283,N_4167,N_4219);
nor U4284 (N_4284,N_4215,N_4146);
or U4285 (N_4285,N_4031,N_4001);
nor U4286 (N_4286,N_4235,N_4249);
or U4287 (N_4287,N_4105,N_4183);
or U4288 (N_4288,N_4103,N_4003);
or U4289 (N_4289,N_4021,N_4089);
xnor U4290 (N_4290,N_4128,N_4231);
or U4291 (N_4291,N_4161,N_4075);
and U4292 (N_4292,N_4140,N_4096);
or U4293 (N_4293,N_4108,N_4193);
nand U4294 (N_4294,N_4223,N_4056);
nor U4295 (N_4295,N_4013,N_4124);
nor U4296 (N_4296,N_4074,N_4081);
nand U4297 (N_4297,N_4106,N_4221);
nor U4298 (N_4298,N_4060,N_4145);
nand U4299 (N_4299,N_4043,N_4063);
and U4300 (N_4300,N_4079,N_4072);
xor U4301 (N_4301,N_4055,N_4143);
nor U4302 (N_4302,N_4113,N_4115);
nand U4303 (N_4303,N_4051,N_4004);
or U4304 (N_4304,N_4222,N_4226);
and U4305 (N_4305,N_4122,N_4149);
nor U4306 (N_4306,N_4212,N_4048);
or U4307 (N_4307,N_4035,N_4247);
xnor U4308 (N_4308,N_4054,N_4142);
nor U4309 (N_4309,N_4195,N_4187);
xor U4310 (N_4310,N_4008,N_4185);
xnor U4311 (N_4311,N_4220,N_4208);
nor U4312 (N_4312,N_4238,N_4069);
or U4313 (N_4313,N_4030,N_4050);
nand U4314 (N_4314,N_4009,N_4135);
and U4315 (N_4315,N_4131,N_4091);
or U4316 (N_4316,N_4207,N_4020);
and U4317 (N_4317,N_4061,N_4196);
xor U4318 (N_4318,N_4200,N_4077);
and U4319 (N_4319,N_4211,N_4237);
nor U4320 (N_4320,N_4206,N_4011);
or U4321 (N_4321,N_4243,N_4244);
xnor U4322 (N_4322,N_4098,N_4202);
xnor U4323 (N_4323,N_4190,N_4080);
or U4324 (N_4324,N_4036,N_4032);
xnor U4325 (N_4325,N_4151,N_4158);
or U4326 (N_4326,N_4078,N_4156);
nand U4327 (N_4327,N_4049,N_4225);
nor U4328 (N_4328,N_4045,N_4232);
and U4329 (N_4329,N_4209,N_4102);
nor U4330 (N_4330,N_4233,N_4038);
and U4331 (N_4331,N_4117,N_4188);
xor U4332 (N_4332,N_4171,N_4201);
and U4333 (N_4333,N_4094,N_4152);
and U4334 (N_4334,N_4059,N_4229);
nor U4335 (N_4335,N_4150,N_4123);
nor U4336 (N_4336,N_4111,N_4118);
nand U4337 (N_4337,N_4203,N_4120);
or U4338 (N_4338,N_4224,N_4213);
nand U4339 (N_4339,N_4006,N_4130);
and U4340 (N_4340,N_4019,N_4000);
nand U4341 (N_4341,N_4107,N_4170);
and U4342 (N_4342,N_4241,N_4216);
xnor U4343 (N_4343,N_4016,N_4162);
nor U4344 (N_4344,N_4097,N_4186);
nand U4345 (N_4345,N_4101,N_4189);
xnor U4346 (N_4346,N_4064,N_4147);
nor U4347 (N_4347,N_4087,N_4168);
or U4348 (N_4348,N_4114,N_4005);
and U4349 (N_4349,N_4014,N_4139);
nor U4350 (N_4350,N_4127,N_4174);
nor U4351 (N_4351,N_4047,N_4065);
and U4352 (N_4352,N_4076,N_4239);
xnor U4353 (N_4353,N_4236,N_4112);
and U4354 (N_4354,N_4041,N_4129);
or U4355 (N_4355,N_4027,N_4084);
nor U4356 (N_4356,N_4095,N_4169);
xnor U4357 (N_4357,N_4179,N_4246);
and U4358 (N_4358,N_4230,N_4132);
nor U4359 (N_4359,N_4068,N_4088);
xnor U4360 (N_4360,N_4090,N_4148);
and U4361 (N_4361,N_4137,N_4109);
xnor U4362 (N_4362,N_4192,N_4116);
nand U4363 (N_4363,N_4033,N_4138);
and U4364 (N_4364,N_4071,N_4025);
nand U4365 (N_4365,N_4104,N_4029);
nor U4366 (N_4366,N_4100,N_4046);
xnor U4367 (N_4367,N_4034,N_4133);
xor U4368 (N_4368,N_4099,N_4228);
nand U4369 (N_4369,N_4086,N_4092);
nor U4370 (N_4370,N_4144,N_4134);
nand U4371 (N_4371,N_4024,N_4015);
nand U4372 (N_4372,N_4194,N_4057);
nor U4373 (N_4373,N_4007,N_4163);
and U4374 (N_4374,N_4181,N_4010);
and U4375 (N_4375,N_4106,N_4181);
or U4376 (N_4376,N_4236,N_4126);
and U4377 (N_4377,N_4007,N_4177);
xor U4378 (N_4378,N_4028,N_4140);
nor U4379 (N_4379,N_4133,N_4173);
and U4380 (N_4380,N_4079,N_4249);
nor U4381 (N_4381,N_4187,N_4134);
and U4382 (N_4382,N_4220,N_4024);
nand U4383 (N_4383,N_4144,N_4128);
and U4384 (N_4384,N_4092,N_4248);
xnor U4385 (N_4385,N_4171,N_4183);
nor U4386 (N_4386,N_4032,N_4103);
nor U4387 (N_4387,N_4059,N_4239);
xor U4388 (N_4388,N_4001,N_4052);
nand U4389 (N_4389,N_4163,N_4095);
xor U4390 (N_4390,N_4083,N_4102);
xnor U4391 (N_4391,N_4012,N_4193);
xor U4392 (N_4392,N_4172,N_4031);
nand U4393 (N_4393,N_4092,N_4062);
or U4394 (N_4394,N_4035,N_4043);
nor U4395 (N_4395,N_4012,N_4014);
nand U4396 (N_4396,N_4198,N_4150);
xnor U4397 (N_4397,N_4229,N_4014);
nor U4398 (N_4398,N_4163,N_4216);
or U4399 (N_4399,N_4172,N_4018);
nor U4400 (N_4400,N_4102,N_4221);
or U4401 (N_4401,N_4090,N_4229);
and U4402 (N_4402,N_4101,N_4118);
or U4403 (N_4403,N_4249,N_4216);
nand U4404 (N_4404,N_4177,N_4068);
or U4405 (N_4405,N_4116,N_4196);
or U4406 (N_4406,N_4036,N_4052);
and U4407 (N_4407,N_4169,N_4079);
and U4408 (N_4408,N_4156,N_4206);
nand U4409 (N_4409,N_4079,N_4234);
nand U4410 (N_4410,N_4153,N_4125);
nand U4411 (N_4411,N_4214,N_4080);
and U4412 (N_4412,N_4177,N_4087);
and U4413 (N_4413,N_4190,N_4171);
or U4414 (N_4414,N_4176,N_4130);
xnor U4415 (N_4415,N_4146,N_4153);
and U4416 (N_4416,N_4145,N_4226);
or U4417 (N_4417,N_4038,N_4019);
xnor U4418 (N_4418,N_4038,N_4197);
nor U4419 (N_4419,N_4200,N_4160);
and U4420 (N_4420,N_4102,N_4217);
xor U4421 (N_4421,N_4111,N_4154);
nor U4422 (N_4422,N_4191,N_4112);
nand U4423 (N_4423,N_4203,N_4005);
and U4424 (N_4424,N_4047,N_4010);
nand U4425 (N_4425,N_4094,N_4187);
and U4426 (N_4426,N_4218,N_4155);
nor U4427 (N_4427,N_4232,N_4020);
nor U4428 (N_4428,N_4184,N_4163);
nor U4429 (N_4429,N_4075,N_4089);
xor U4430 (N_4430,N_4082,N_4091);
or U4431 (N_4431,N_4231,N_4190);
xor U4432 (N_4432,N_4021,N_4110);
xor U4433 (N_4433,N_4046,N_4248);
nand U4434 (N_4434,N_4117,N_4017);
nor U4435 (N_4435,N_4024,N_4022);
nand U4436 (N_4436,N_4160,N_4033);
nand U4437 (N_4437,N_4204,N_4070);
or U4438 (N_4438,N_4069,N_4072);
nor U4439 (N_4439,N_4199,N_4093);
xor U4440 (N_4440,N_4145,N_4162);
and U4441 (N_4441,N_4139,N_4104);
or U4442 (N_4442,N_4016,N_4177);
nor U4443 (N_4443,N_4248,N_4181);
or U4444 (N_4444,N_4237,N_4047);
xnor U4445 (N_4445,N_4038,N_4104);
nand U4446 (N_4446,N_4154,N_4197);
nor U4447 (N_4447,N_4039,N_4000);
and U4448 (N_4448,N_4031,N_4126);
and U4449 (N_4449,N_4196,N_4058);
nand U4450 (N_4450,N_4003,N_4014);
xnor U4451 (N_4451,N_4220,N_4169);
and U4452 (N_4452,N_4218,N_4198);
nand U4453 (N_4453,N_4113,N_4157);
or U4454 (N_4454,N_4004,N_4242);
nor U4455 (N_4455,N_4110,N_4080);
nand U4456 (N_4456,N_4018,N_4000);
nand U4457 (N_4457,N_4159,N_4021);
nand U4458 (N_4458,N_4143,N_4012);
or U4459 (N_4459,N_4039,N_4123);
nor U4460 (N_4460,N_4051,N_4092);
nor U4461 (N_4461,N_4099,N_4066);
nand U4462 (N_4462,N_4039,N_4095);
nor U4463 (N_4463,N_4194,N_4245);
nor U4464 (N_4464,N_4087,N_4122);
nand U4465 (N_4465,N_4160,N_4040);
xnor U4466 (N_4466,N_4003,N_4204);
or U4467 (N_4467,N_4014,N_4183);
nor U4468 (N_4468,N_4203,N_4162);
nand U4469 (N_4469,N_4161,N_4236);
nand U4470 (N_4470,N_4028,N_4087);
nor U4471 (N_4471,N_4185,N_4019);
nand U4472 (N_4472,N_4076,N_4022);
nor U4473 (N_4473,N_4192,N_4195);
nor U4474 (N_4474,N_4064,N_4173);
nor U4475 (N_4475,N_4047,N_4020);
nand U4476 (N_4476,N_4043,N_4189);
nor U4477 (N_4477,N_4233,N_4031);
nor U4478 (N_4478,N_4010,N_4217);
nor U4479 (N_4479,N_4171,N_4199);
xnor U4480 (N_4480,N_4119,N_4200);
nor U4481 (N_4481,N_4023,N_4213);
or U4482 (N_4482,N_4219,N_4090);
nor U4483 (N_4483,N_4136,N_4117);
nand U4484 (N_4484,N_4035,N_4087);
nand U4485 (N_4485,N_4158,N_4017);
or U4486 (N_4486,N_4001,N_4007);
nor U4487 (N_4487,N_4149,N_4218);
or U4488 (N_4488,N_4236,N_4195);
nand U4489 (N_4489,N_4019,N_4229);
xor U4490 (N_4490,N_4057,N_4246);
xor U4491 (N_4491,N_4111,N_4059);
nor U4492 (N_4492,N_4079,N_4198);
or U4493 (N_4493,N_4144,N_4124);
and U4494 (N_4494,N_4247,N_4232);
and U4495 (N_4495,N_4143,N_4061);
nand U4496 (N_4496,N_4107,N_4206);
and U4497 (N_4497,N_4117,N_4180);
and U4498 (N_4498,N_4201,N_4030);
or U4499 (N_4499,N_4037,N_4098);
nand U4500 (N_4500,N_4416,N_4325);
and U4501 (N_4501,N_4487,N_4351);
nor U4502 (N_4502,N_4410,N_4459);
or U4503 (N_4503,N_4397,N_4262);
and U4504 (N_4504,N_4355,N_4400);
or U4505 (N_4505,N_4476,N_4302);
or U4506 (N_4506,N_4346,N_4404);
and U4507 (N_4507,N_4456,N_4342);
nand U4508 (N_4508,N_4496,N_4253);
xnor U4509 (N_4509,N_4354,N_4465);
and U4510 (N_4510,N_4290,N_4421);
and U4511 (N_4511,N_4449,N_4499);
nand U4512 (N_4512,N_4494,N_4468);
nor U4513 (N_4513,N_4335,N_4424);
nor U4514 (N_4514,N_4357,N_4438);
nand U4515 (N_4515,N_4384,N_4292);
and U4516 (N_4516,N_4329,N_4265);
xor U4517 (N_4517,N_4293,N_4311);
nor U4518 (N_4518,N_4379,N_4339);
and U4519 (N_4519,N_4398,N_4369);
or U4520 (N_4520,N_4442,N_4287);
nor U4521 (N_4521,N_4427,N_4285);
xnor U4522 (N_4522,N_4337,N_4353);
and U4523 (N_4523,N_4446,N_4399);
and U4524 (N_4524,N_4498,N_4394);
xnor U4525 (N_4525,N_4362,N_4288);
nand U4526 (N_4526,N_4386,N_4368);
or U4527 (N_4527,N_4435,N_4323);
and U4528 (N_4528,N_4270,N_4380);
xor U4529 (N_4529,N_4327,N_4305);
xnor U4530 (N_4530,N_4475,N_4412);
xor U4531 (N_4531,N_4331,N_4343);
nand U4532 (N_4532,N_4491,N_4461);
or U4533 (N_4533,N_4291,N_4372);
nor U4534 (N_4534,N_4388,N_4250);
xnor U4535 (N_4535,N_4350,N_4455);
xnor U4536 (N_4536,N_4434,N_4359);
and U4537 (N_4537,N_4352,N_4364);
or U4538 (N_4538,N_4252,N_4425);
nand U4539 (N_4539,N_4382,N_4304);
and U4540 (N_4540,N_4432,N_4445);
or U4541 (N_4541,N_4480,N_4392);
or U4542 (N_4542,N_4276,N_4381);
and U4543 (N_4543,N_4328,N_4486);
nor U4544 (N_4544,N_4467,N_4280);
nor U4545 (N_4545,N_4474,N_4450);
xor U4546 (N_4546,N_4281,N_4439);
xnor U4547 (N_4547,N_4306,N_4300);
and U4548 (N_4548,N_4294,N_4411);
and U4549 (N_4549,N_4460,N_4254);
nand U4550 (N_4550,N_4275,N_4373);
nor U4551 (N_4551,N_4387,N_4279);
nor U4552 (N_4552,N_4395,N_4473);
and U4553 (N_4553,N_4297,N_4308);
or U4554 (N_4554,N_4322,N_4301);
nand U4555 (N_4555,N_4471,N_4433);
and U4556 (N_4556,N_4272,N_4391);
xor U4557 (N_4557,N_4356,N_4436);
nor U4558 (N_4558,N_4454,N_4345);
xnor U4559 (N_4559,N_4361,N_4430);
xnor U4560 (N_4560,N_4371,N_4409);
or U4561 (N_4561,N_4260,N_4336);
and U4562 (N_4562,N_4313,N_4366);
and U4563 (N_4563,N_4413,N_4403);
xnor U4564 (N_4564,N_4451,N_4264);
nor U4565 (N_4565,N_4268,N_4488);
xnor U4566 (N_4566,N_4470,N_4319);
nor U4567 (N_4567,N_4423,N_4481);
nor U4568 (N_4568,N_4495,N_4263);
or U4569 (N_4569,N_4312,N_4375);
xor U4570 (N_4570,N_4278,N_4490);
nand U4571 (N_4571,N_4431,N_4367);
or U4572 (N_4572,N_4377,N_4390);
xor U4573 (N_4573,N_4269,N_4472);
nor U4574 (N_4574,N_4310,N_4296);
nor U4575 (N_4575,N_4447,N_4466);
nand U4576 (N_4576,N_4259,N_4374);
xnor U4577 (N_4577,N_4437,N_4360);
and U4578 (N_4578,N_4358,N_4271);
nor U4579 (N_4579,N_4251,N_4349);
or U4580 (N_4580,N_4370,N_4332);
nand U4581 (N_4581,N_4482,N_4317);
xor U4582 (N_4582,N_4315,N_4378);
and U4583 (N_4583,N_4383,N_4273);
nor U4584 (N_4584,N_4420,N_4258);
nor U4585 (N_4585,N_4396,N_4469);
and U4586 (N_4586,N_4457,N_4277);
and U4587 (N_4587,N_4406,N_4255);
nor U4588 (N_4588,N_4333,N_4334);
and U4589 (N_4589,N_4340,N_4326);
nand U4590 (N_4590,N_4402,N_4330);
nand U4591 (N_4591,N_4483,N_4274);
or U4592 (N_4592,N_4489,N_4295);
nand U4593 (N_4593,N_4365,N_4320);
or U4594 (N_4594,N_4289,N_4448);
and U4595 (N_4595,N_4307,N_4284);
xnor U4596 (N_4596,N_4485,N_4453);
or U4597 (N_4597,N_4385,N_4401);
and U4598 (N_4598,N_4415,N_4422);
and U4599 (N_4599,N_4299,N_4298);
nor U4600 (N_4600,N_4464,N_4428);
or U4601 (N_4601,N_4419,N_4493);
nor U4602 (N_4602,N_4338,N_4478);
or U4603 (N_4603,N_4458,N_4462);
and U4604 (N_4604,N_4347,N_4484);
and U4605 (N_4605,N_4376,N_4479);
nor U4606 (N_4606,N_4429,N_4266);
nor U4607 (N_4607,N_4363,N_4321);
and U4608 (N_4608,N_4408,N_4405);
nand U4609 (N_4609,N_4324,N_4261);
nor U4610 (N_4610,N_4348,N_4267);
or U4611 (N_4611,N_4414,N_4257);
xor U4612 (N_4612,N_4452,N_4393);
or U4613 (N_4613,N_4314,N_4341);
and U4614 (N_4614,N_4303,N_4309);
or U4615 (N_4615,N_4418,N_4318);
or U4616 (N_4616,N_4316,N_4344);
nand U4617 (N_4617,N_4463,N_4282);
nand U4618 (N_4618,N_4389,N_4286);
nor U4619 (N_4619,N_4417,N_4477);
or U4620 (N_4620,N_4492,N_4283);
xnor U4621 (N_4621,N_4443,N_4444);
nor U4622 (N_4622,N_4440,N_4407);
nand U4623 (N_4623,N_4256,N_4441);
nor U4624 (N_4624,N_4497,N_4426);
nor U4625 (N_4625,N_4486,N_4406);
nor U4626 (N_4626,N_4380,N_4250);
xnor U4627 (N_4627,N_4287,N_4356);
nand U4628 (N_4628,N_4441,N_4463);
or U4629 (N_4629,N_4300,N_4457);
nor U4630 (N_4630,N_4495,N_4336);
and U4631 (N_4631,N_4464,N_4303);
nor U4632 (N_4632,N_4489,N_4372);
nor U4633 (N_4633,N_4435,N_4371);
xor U4634 (N_4634,N_4445,N_4323);
nor U4635 (N_4635,N_4416,N_4318);
nor U4636 (N_4636,N_4312,N_4405);
xor U4637 (N_4637,N_4282,N_4280);
nand U4638 (N_4638,N_4298,N_4428);
and U4639 (N_4639,N_4351,N_4458);
nand U4640 (N_4640,N_4412,N_4268);
nor U4641 (N_4641,N_4336,N_4263);
nor U4642 (N_4642,N_4431,N_4330);
nor U4643 (N_4643,N_4384,N_4272);
or U4644 (N_4644,N_4374,N_4343);
and U4645 (N_4645,N_4405,N_4431);
or U4646 (N_4646,N_4381,N_4282);
nor U4647 (N_4647,N_4328,N_4384);
or U4648 (N_4648,N_4277,N_4470);
nor U4649 (N_4649,N_4308,N_4302);
xnor U4650 (N_4650,N_4352,N_4451);
nand U4651 (N_4651,N_4475,N_4374);
and U4652 (N_4652,N_4492,N_4363);
nor U4653 (N_4653,N_4479,N_4339);
and U4654 (N_4654,N_4360,N_4427);
or U4655 (N_4655,N_4328,N_4279);
nor U4656 (N_4656,N_4355,N_4281);
xnor U4657 (N_4657,N_4326,N_4485);
or U4658 (N_4658,N_4478,N_4497);
nand U4659 (N_4659,N_4273,N_4457);
or U4660 (N_4660,N_4279,N_4288);
xor U4661 (N_4661,N_4347,N_4366);
nor U4662 (N_4662,N_4259,N_4434);
xnor U4663 (N_4663,N_4270,N_4365);
and U4664 (N_4664,N_4292,N_4298);
nor U4665 (N_4665,N_4436,N_4444);
or U4666 (N_4666,N_4395,N_4274);
or U4667 (N_4667,N_4339,N_4380);
xor U4668 (N_4668,N_4286,N_4459);
or U4669 (N_4669,N_4349,N_4309);
xnor U4670 (N_4670,N_4458,N_4459);
xor U4671 (N_4671,N_4256,N_4408);
or U4672 (N_4672,N_4360,N_4375);
nand U4673 (N_4673,N_4440,N_4442);
or U4674 (N_4674,N_4474,N_4399);
and U4675 (N_4675,N_4491,N_4453);
xnor U4676 (N_4676,N_4322,N_4495);
nor U4677 (N_4677,N_4406,N_4414);
nand U4678 (N_4678,N_4464,N_4437);
nor U4679 (N_4679,N_4432,N_4461);
nor U4680 (N_4680,N_4492,N_4277);
or U4681 (N_4681,N_4266,N_4396);
xor U4682 (N_4682,N_4440,N_4422);
xnor U4683 (N_4683,N_4339,N_4496);
or U4684 (N_4684,N_4309,N_4301);
nand U4685 (N_4685,N_4269,N_4320);
xor U4686 (N_4686,N_4362,N_4311);
nand U4687 (N_4687,N_4304,N_4443);
or U4688 (N_4688,N_4370,N_4436);
and U4689 (N_4689,N_4335,N_4302);
nand U4690 (N_4690,N_4295,N_4406);
and U4691 (N_4691,N_4269,N_4315);
or U4692 (N_4692,N_4280,N_4353);
or U4693 (N_4693,N_4371,N_4495);
nor U4694 (N_4694,N_4255,N_4466);
xor U4695 (N_4695,N_4360,N_4354);
and U4696 (N_4696,N_4399,N_4414);
nor U4697 (N_4697,N_4376,N_4306);
nand U4698 (N_4698,N_4461,N_4256);
xnor U4699 (N_4699,N_4436,N_4413);
or U4700 (N_4700,N_4268,N_4415);
nand U4701 (N_4701,N_4447,N_4428);
xnor U4702 (N_4702,N_4378,N_4414);
or U4703 (N_4703,N_4342,N_4280);
nor U4704 (N_4704,N_4383,N_4385);
nand U4705 (N_4705,N_4453,N_4331);
nor U4706 (N_4706,N_4435,N_4297);
and U4707 (N_4707,N_4324,N_4292);
or U4708 (N_4708,N_4386,N_4359);
and U4709 (N_4709,N_4444,N_4346);
and U4710 (N_4710,N_4268,N_4267);
xnor U4711 (N_4711,N_4285,N_4417);
nor U4712 (N_4712,N_4451,N_4338);
nor U4713 (N_4713,N_4307,N_4359);
or U4714 (N_4714,N_4341,N_4458);
nand U4715 (N_4715,N_4481,N_4489);
or U4716 (N_4716,N_4362,N_4350);
nor U4717 (N_4717,N_4297,N_4291);
xnor U4718 (N_4718,N_4348,N_4484);
or U4719 (N_4719,N_4490,N_4477);
or U4720 (N_4720,N_4299,N_4303);
and U4721 (N_4721,N_4388,N_4369);
or U4722 (N_4722,N_4443,N_4286);
nor U4723 (N_4723,N_4377,N_4426);
nand U4724 (N_4724,N_4461,N_4458);
nor U4725 (N_4725,N_4359,N_4436);
nand U4726 (N_4726,N_4487,N_4287);
and U4727 (N_4727,N_4256,N_4463);
and U4728 (N_4728,N_4319,N_4342);
or U4729 (N_4729,N_4251,N_4496);
nor U4730 (N_4730,N_4250,N_4467);
nor U4731 (N_4731,N_4437,N_4469);
or U4732 (N_4732,N_4382,N_4424);
nor U4733 (N_4733,N_4320,N_4480);
nand U4734 (N_4734,N_4474,N_4271);
and U4735 (N_4735,N_4472,N_4451);
nor U4736 (N_4736,N_4286,N_4337);
xnor U4737 (N_4737,N_4254,N_4473);
or U4738 (N_4738,N_4402,N_4296);
nor U4739 (N_4739,N_4384,N_4312);
and U4740 (N_4740,N_4289,N_4341);
and U4741 (N_4741,N_4385,N_4476);
nor U4742 (N_4742,N_4326,N_4262);
and U4743 (N_4743,N_4453,N_4353);
nand U4744 (N_4744,N_4460,N_4476);
or U4745 (N_4745,N_4452,N_4474);
and U4746 (N_4746,N_4313,N_4321);
nor U4747 (N_4747,N_4463,N_4415);
xnor U4748 (N_4748,N_4476,N_4422);
nor U4749 (N_4749,N_4466,N_4496);
or U4750 (N_4750,N_4543,N_4540);
and U4751 (N_4751,N_4514,N_4561);
nor U4752 (N_4752,N_4521,N_4707);
or U4753 (N_4753,N_4718,N_4506);
nor U4754 (N_4754,N_4591,N_4530);
and U4755 (N_4755,N_4558,N_4672);
or U4756 (N_4756,N_4713,N_4600);
or U4757 (N_4757,N_4607,N_4578);
xnor U4758 (N_4758,N_4715,N_4692);
xor U4759 (N_4759,N_4532,N_4687);
xor U4760 (N_4760,N_4571,N_4537);
and U4761 (N_4761,N_4716,N_4573);
nor U4762 (N_4762,N_4748,N_4524);
nor U4763 (N_4763,N_4542,N_4701);
or U4764 (N_4764,N_4697,N_4720);
or U4765 (N_4765,N_4722,N_4671);
or U4766 (N_4766,N_4733,N_4717);
xor U4767 (N_4767,N_4628,N_4728);
and U4768 (N_4768,N_4538,N_4659);
xor U4769 (N_4769,N_4550,N_4611);
or U4770 (N_4770,N_4556,N_4545);
nor U4771 (N_4771,N_4566,N_4685);
nor U4772 (N_4772,N_4551,N_4614);
xnor U4773 (N_4773,N_4632,N_4592);
or U4774 (N_4774,N_4652,N_4665);
xor U4775 (N_4775,N_4670,N_4526);
or U4776 (N_4776,N_4554,N_4679);
nand U4777 (N_4777,N_4533,N_4529);
and U4778 (N_4778,N_4518,N_4662);
or U4779 (N_4779,N_4688,N_4702);
and U4780 (N_4780,N_4582,N_4613);
xnor U4781 (N_4781,N_4735,N_4500);
or U4782 (N_4782,N_4503,N_4719);
nand U4783 (N_4783,N_4516,N_4609);
nand U4784 (N_4784,N_4536,N_4653);
or U4785 (N_4785,N_4507,N_4565);
or U4786 (N_4786,N_4563,N_4546);
nor U4787 (N_4787,N_4658,N_4648);
or U4788 (N_4788,N_4657,N_4664);
or U4789 (N_4789,N_4669,N_4605);
or U4790 (N_4790,N_4559,N_4544);
xor U4791 (N_4791,N_4743,N_4705);
and U4792 (N_4792,N_4625,N_4527);
or U4793 (N_4793,N_4636,N_4564);
xnor U4794 (N_4794,N_4531,N_4595);
nand U4795 (N_4795,N_4520,N_4673);
nand U4796 (N_4796,N_4726,N_4570);
xnor U4797 (N_4797,N_4689,N_4642);
nand U4798 (N_4798,N_4721,N_4691);
xor U4799 (N_4799,N_4513,N_4620);
nor U4800 (N_4800,N_4598,N_4647);
or U4801 (N_4801,N_4599,N_4553);
nor U4802 (N_4802,N_4627,N_4700);
nor U4803 (N_4803,N_4637,N_4562);
or U4804 (N_4804,N_4633,N_4712);
nor U4805 (N_4805,N_4575,N_4621);
xor U4806 (N_4806,N_4504,N_4680);
and U4807 (N_4807,N_4731,N_4638);
or U4808 (N_4808,N_4738,N_4698);
xor U4809 (N_4809,N_4547,N_4626);
or U4810 (N_4810,N_4744,N_4668);
nand U4811 (N_4811,N_4683,N_4509);
and U4812 (N_4812,N_4581,N_4615);
nand U4813 (N_4813,N_4624,N_4590);
xor U4814 (N_4814,N_4711,N_4656);
and U4815 (N_4815,N_4661,N_4639);
nand U4816 (N_4816,N_4714,N_4629);
or U4817 (N_4817,N_4696,N_4597);
or U4818 (N_4818,N_4667,N_4522);
or U4819 (N_4819,N_4727,N_4646);
and U4820 (N_4820,N_4616,N_4684);
and U4821 (N_4821,N_4508,N_4552);
and U4822 (N_4822,N_4732,N_4677);
nor U4823 (N_4823,N_4585,N_4724);
nor U4824 (N_4824,N_4706,N_4623);
xnor U4825 (N_4825,N_4539,N_4502);
nor U4826 (N_4826,N_4549,N_4663);
or U4827 (N_4827,N_4630,N_4650);
nand U4828 (N_4828,N_4560,N_4567);
or U4829 (N_4829,N_4501,N_4589);
nor U4830 (N_4830,N_4534,N_4674);
or U4831 (N_4831,N_4675,N_4512);
or U4832 (N_4832,N_4606,N_4736);
or U4833 (N_4833,N_4710,N_4645);
nor U4834 (N_4834,N_4681,N_4517);
xor U4835 (N_4835,N_4525,N_4557);
xor U4836 (N_4836,N_4569,N_4693);
xnor U4837 (N_4837,N_4574,N_4594);
and U4838 (N_4838,N_4709,N_4587);
and U4839 (N_4839,N_4619,N_4643);
nand U4840 (N_4840,N_4519,N_4608);
nand U4841 (N_4841,N_4580,N_4654);
xnor U4842 (N_4842,N_4686,N_4572);
or U4843 (N_4843,N_4737,N_4678);
nand U4844 (N_4844,N_4588,N_4584);
xor U4845 (N_4845,N_4745,N_4666);
nor U4846 (N_4846,N_4610,N_4635);
nand U4847 (N_4847,N_4541,N_4510);
or U4848 (N_4848,N_4548,N_4690);
xor U4849 (N_4849,N_4505,N_4640);
nor U4850 (N_4850,N_4577,N_4703);
nand U4851 (N_4851,N_4602,N_4741);
or U4852 (N_4852,N_4660,N_4746);
nor U4853 (N_4853,N_4695,N_4576);
xnor U4854 (N_4854,N_4644,N_4622);
nor U4855 (N_4855,N_4740,N_4649);
nand U4856 (N_4856,N_4586,N_4604);
and U4857 (N_4857,N_4528,N_4593);
or U4858 (N_4858,N_4739,N_4708);
or U4859 (N_4859,N_4596,N_4634);
nor U4860 (N_4860,N_4704,N_4641);
and U4861 (N_4861,N_4676,N_4617);
nor U4862 (N_4862,N_4618,N_4612);
and U4863 (N_4863,N_4723,N_4631);
nor U4864 (N_4864,N_4729,N_4651);
nor U4865 (N_4865,N_4749,N_4655);
and U4866 (N_4866,N_4730,N_4568);
xor U4867 (N_4867,N_4699,N_4682);
nor U4868 (N_4868,N_4555,N_4583);
nand U4869 (N_4869,N_4725,N_4579);
or U4870 (N_4870,N_4734,N_4535);
xor U4871 (N_4871,N_4523,N_4511);
nor U4872 (N_4872,N_4603,N_4747);
nand U4873 (N_4873,N_4694,N_4601);
nand U4874 (N_4874,N_4515,N_4742);
and U4875 (N_4875,N_4662,N_4680);
nor U4876 (N_4876,N_4730,N_4693);
or U4877 (N_4877,N_4731,N_4747);
or U4878 (N_4878,N_4698,N_4614);
or U4879 (N_4879,N_4502,N_4675);
or U4880 (N_4880,N_4596,N_4716);
or U4881 (N_4881,N_4700,N_4563);
xor U4882 (N_4882,N_4631,N_4568);
or U4883 (N_4883,N_4503,N_4532);
or U4884 (N_4884,N_4744,N_4573);
xor U4885 (N_4885,N_4604,N_4633);
or U4886 (N_4886,N_4624,N_4561);
xor U4887 (N_4887,N_4584,N_4551);
nand U4888 (N_4888,N_4540,N_4532);
nor U4889 (N_4889,N_4746,N_4560);
xnor U4890 (N_4890,N_4517,N_4702);
nand U4891 (N_4891,N_4721,N_4577);
nor U4892 (N_4892,N_4689,N_4692);
and U4893 (N_4893,N_4551,N_4708);
or U4894 (N_4894,N_4733,N_4555);
or U4895 (N_4895,N_4746,N_4569);
or U4896 (N_4896,N_4623,N_4703);
nor U4897 (N_4897,N_4551,N_4586);
xor U4898 (N_4898,N_4664,N_4653);
nand U4899 (N_4899,N_4621,N_4614);
nor U4900 (N_4900,N_4619,N_4676);
and U4901 (N_4901,N_4687,N_4602);
and U4902 (N_4902,N_4580,N_4704);
and U4903 (N_4903,N_4577,N_4511);
or U4904 (N_4904,N_4523,N_4573);
and U4905 (N_4905,N_4531,N_4505);
and U4906 (N_4906,N_4609,N_4671);
nand U4907 (N_4907,N_4592,N_4645);
xor U4908 (N_4908,N_4731,N_4522);
nand U4909 (N_4909,N_4631,N_4635);
or U4910 (N_4910,N_4735,N_4640);
and U4911 (N_4911,N_4644,N_4607);
nor U4912 (N_4912,N_4672,N_4604);
or U4913 (N_4913,N_4548,N_4718);
xnor U4914 (N_4914,N_4690,N_4737);
xnor U4915 (N_4915,N_4720,N_4561);
and U4916 (N_4916,N_4706,N_4545);
and U4917 (N_4917,N_4649,N_4553);
and U4918 (N_4918,N_4506,N_4733);
or U4919 (N_4919,N_4579,N_4632);
and U4920 (N_4920,N_4687,N_4619);
and U4921 (N_4921,N_4683,N_4556);
and U4922 (N_4922,N_4547,N_4555);
nor U4923 (N_4923,N_4562,N_4666);
and U4924 (N_4924,N_4743,N_4696);
and U4925 (N_4925,N_4729,N_4581);
or U4926 (N_4926,N_4597,N_4608);
or U4927 (N_4927,N_4564,N_4600);
or U4928 (N_4928,N_4663,N_4568);
and U4929 (N_4929,N_4571,N_4538);
nor U4930 (N_4930,N_4731,N_4536);
nand U4931 (N_4931,N_4609,N_4653);
nor U4932 (N_4932,N_4655,N_4730);
nand U4933 (N_4933,N_4541,N_4502);
or U4934 (N_4934,N_4714,N_4593);
nand U4935 (N_4935,N_4517,N_4613);
or U4936 (N_4936,N_4635,N_4650);
nand U4937 (N_4937,N_4684,N_4615);
and U4938 (N_4938,N_4586,N_4564);
nand U4939 (N_4939,N_4600,N_4601);
nor U4940 (N_4940,N_4742,N_4651);
nor U4941 (N_4941,N_4619,N_4599);
nor U4942 (N_4942,N_4549,N_4698);
nor U4943 (N_4943,N_4502,N_4623);
and U4944 (N_4944,N_4651,N_4525);
xnor U4945 (N_4945,N_4565,N_4708);
or U4946 (N_4946,N_4650,N_4616);
and U4947 (N_4947,N_4666,N_4654);
nand U4948 (N_4948,N_4695,N_4653);
nand U4949 (N_4949,N_4694,N_4683);
nand U4950 (N_4950,N_4724,N_4580);
and U4951 (N_4951,N_4553,N_4656);
and U4952 (N_4952,N_4581,N_4648);
nand U4953 (N_4953,N_4629,N_4651);
or U4954 (N_4954,N_4655,N_4600);
nand U4955 (N_4955,N_4625,N_4573);
or U4956 (N_4956,N_4686,N_4613);
and U4957 (N_4957,N_4669,N_4659);
xor U4958 (N_4958,N_4587,N_4689);
or U4959 (N_4959,N_4698,N_4711);
and U4960 (N_4960,N_4718,N_4554);
nor U4961 (N_4961,N_4549,N_4517);
nand U4962 (N_4962,N_4622,N_4721);
or U4963 (N_4963,N_4701,N_4646);
xnor U4964 (N_4964,N_4611,N_4571);
or U4965 (N_4965,N_4701,N_4676);
nor U4966 (N_4966,N_4665,N_4613);
or U4967 (N_4967,N_4571,N_4550);
or U4968 (N_4968,N_4659,N_4593);
or U4969 (N_4969,N_4530,N_4627);
xor U4970 (N_4970,N_4584,N_4575);
nor U4971 (N_4971,N_4535,N_4633);
xnor U4972 (N_4972,N_4547,N_4700);
xnor U4973 (N_4973,N_4601,N_4501);
xor U4974 (N_4974,N_4503,N_4504);
and U4975 (N_4975,N_4531,N_4671);
nand U4976 (N_4976,N_4706,N_4571);
nor U4977 (N_4977,N_4685,N_4684);
or U4978 (N_4978,N_4728,N_4608);
xnor U4979 (N_4979,N_4516,N_4667);
or U4980 (N_4980,N_4652,N_4571);
xor U4981 (N_4981,N_4539,N_4710);
xor U4982 (N_4982,N_4687,N_4684);
xnor U4983 (N_4983,N_4511,N_4607);
nand U4984 (N_4984,N_4543,N_4665);
nand U4985 (N_4985,N_4712,N_4693);
or U4986 (N_4986,N_4549,N_4592);
nand U4987 (N_4987,N_4748,N_4618);
nor U4988 (N_4988,N_4584,N_4718);
xor U4989 (N_4989,N_4543,N_4590);
and U4990 (N_4990,N_4532,N_4730);
or U4991 (N_4991,N_4717,N_4586);
nand U4992 (N_4992,N_4591,N_4624);
xor U4993 (N_4993,N_4637,N_4647);
xnor U4994 (N_4994,N_4740,N_4639);
nand U4995 (N_4995,N_4640,N_4564);
nand U4996 (N_4996,N_4633,N_4680);
nor U4997 (N_4997,N_4699,N_4585);
xor U4998 (N_4998,N_4675,N_4653);
or U4999 (N_4999,N_4565,N_4512);
and U5000 (N_5000,N_4862,N_4898);
and U5001 (N_5001,N_4835,N_4901);
nor U5002 (N_5002,N_4857,N_4941);
xnor U5003 (N_5003,N_4895,N_4772);
xor U5004 (N_5004,N_4939,N_4832);
nor U5005 (N_5005,N_4973,N_4969);
nand U5006 (N_5006,N_4871,N_4816);
and U5007 (N_5007,N_4762,N_4882);
nand U5008 (N_5008,N_4866,N_4984);
xnor U5009 (N_5009,N_4810,N_4783);
or U5010 (N_5010,N_4977,N_4915);
or U5011 (N_5011,N_4809,N_4927);
nor U5012 (N_5012,N_4775,N_4983);
or U5013 (N_5013,N_4885,N_4880);
or U5014 (N_5014,N_4753,N_4891);
nor U5015 (N_5015,N_4851,N_4868);
nor U5016 (N_5016,N_4814,N_4801);
nand U5017 (N_5017,N_4834,N_4833);
nand U5018 (N_5018,N_4815,N_4813);
nand U5019 (N_5019,N_4930,N_4959);
or U5020 (N_5020,N_4799,N_4852);
nor U5021 (N_5021,N_4761,N_4933);
or U5022 (N_5022,N_4957,N_4981);
and U5023 (N_5023,N_4844,N_4900);
nor U5024 (N_5024,N_4917,N_4763);
nand U5025 (N_5025,N_4767,N_4796);
or U5026 (N_5026,N_4802,N_4896);
or U5027 (N_5027,N_4926,N_4899);
xnor U5028 (N_5028,N_4911,N_4777);
nor U5029 (N_5029,N_4966,N_4770);
or U5030 (N_5030,N_4924,N_4877);
nand U5031 (N_5031,N_4758,N_4876);
nor U5032 (N_5032,N_4794,N_4902);
xnor U5033 (N_5033,N_4784,N_4993);
or U5034 (N_5034,N_4995,N_4962);
and U5035 (N_5035,N_4764,N_4994);
nand U5036 (N_5036,N_4780,N_4855);
or U5037 (N_5037,N_4823,N_4963);
xor U5038 (N_5038,N_4782,N_4848);
and U5039 (N_5039,N_4918,N_4912);
xor U5040 (N_5040,N_4869,N_4904);
nand U5041 (N_5041,N_4867,N_4890);
and U5042 (N_5042,N_4916,N_4906);
xnor U5043 (N_5043,N_4791,N_4826);
nor U5044 (N_5044,N_4932,N_4800);
or U5045 (N_5045,N_4840,N_4965);
or U5046 (N_5046,N_4831,N_4828);
and U5047 (N_5047,N_4886,N_4953);
xnor U5048 (N_5048,N_4849,N_4980);
xnor U5049 (N_5049,N_4892,N_4845);
nor U5050 (N_5050,N_4944,N_4768);
and U5051 (N_5051,N_4883,N_4946);
nand U5052 (N_5052,N_4818,N_4872);
and U5053 (N_5053,N_4894,N_4888);
nor U5054 (N_5054,N_4803,N_4861);
and U5055 (N_5055,N_4804,N_4884);
and U5056 (N_5056,N_4934,N_4864);
nand U5057 (N_5057,N_4829,N_4875);
xor U5058 (N_5058,N_4914,N_4846);
nor U5059 (N_5059,N_4750,N_4908);
or U5060 (N_5060,N_4893,N_4822);
nand U5061 (N_5061,N_4997,N_4986);
or U5062 (N_5062,N_4757,N_4854);
or U5063 (N_5063,N_4769,N_4942);
nand U5064 (N_5064,N_4931,N_4759);
and U5065 (N_5065,N_4873,N_4805);
or U5066 (N_5066,N_4811,N_4755);
or U5067 (N_5067,N_4935,N_4999);
nand U5068 (N_5068,N_4856,N_4827);
or U5069 (N_5069,N_4964,N_4905);
xnor U5070 (N_5070,N_4787,N_4937);
nand U5071 (N_5071,N_4774,N_4921);
nor U5072 (N_5072,N_4936,N_4853);
xnor U5073 (N_5073,N_4847,N_4863);
nor U5074 (N_5074,N_4878,N_4954);
and U5075 (N_5075,N_4989,N_4760);
nand U5076 (N_5076,N_4889,N_4771);
nor U5077 (N_5077,N_4985,N_4975);
xor U5078 (N_5078,N_4990,N_4788);
xnor U5079 (N_5079,N_4988,N_4991);
or U5080 (N_5080,N_4859,N_4836);
or U5081 (N_5081,N_4843,N_4907);
nand U5082 (N_5082,N_4779,N_4979);
xor U5083 (N_5083,N_4913,N_4909);
xnor U5084 (N_5084,N_4881,N_4830);
or U5085 (N_5085,N_4785,N_4920);
and U5086 (N_5086,N_4879,N_4837);
nor U5087 (N_5087,N_4961,N_4922);
nand U5088 (N_5088,N_4797,N_4955);
nor U5089 (N_5089,N_4978,N_4776);
xor U5090 (N_5090,N_4992,N_4972);
nor U5091 (N_5091,N_4948,N_4943);
and U5092 (N_5092,N_4850,N_4951);
or U5093 (N_5093,N_4968,N_4923);
nor U5094 (N_5094,N_4945,N_4967);
or U5095 (N_5095,N_4919,N_4950);
and U5096 (N_5096,N_4751,N_4765);
nand U5097 (N_5097,N_4971,N_4910);
and U5098 (N_5098,N_4874,N_4903);
and U5099 (N_5099,N_4798,N_4825);
or U5100 (N_5100,N_4938,N_4817);
and U5101 (N_5101,N_4929,N_4806);
nand U5102 (N_5102,N_4841,N_4773);
nor U5103 (N_5103,N_4976,N_4786);
nand U5104 (N_5104,N_4820,N_4858);
xnor U5105 (N_5105,N_4870,N_4789);
and U5106 (N_5106,N_4756,N_4958);
xnor U5107 (N_5107,N_4778,N_4952);
xnor U5108 (N_5108,N_4974,N_4790);
xor U5109 (N_5109,N_4996,N_4860);
and U5110 (N_5110,N_4793,N_4897);
or U5111 (N_5111,N_4819,N_4795);
xor U5112 (N_5112,N_4949,N_4752);
and U5113 (N_5113,N_4998,N_4970);
or U5114 (N_5114,N_4838,N_4839);
xnor U5115 (N_5115,N_4940,N_4766);
and U5116 (N_5116,N_4956,N_4792);
and U5117 (N_5117,N_4865,N_4887);
or U5118 (N_5118,N_4781,N_4821);
xnor U5119 (N_5119,N_4987,N_4960);
or U5120 (N_5120,N_4842,N_4808);
or U5121 (N_5121,N_4947,N_4982);
nor U5122 (N_5122,N_4812,N_4928);
nand U5123 (N_5123,N_4824,N_4807);
or U5124 (N_5124,N_4754,N_4925);
nand U5125 (N_5125,N_4875,N_4911);
and U5126 (N_5126,N_4819,N_4840);
nand U5127 (N_5127,N_4809,N_4821);
and U5128 (N_5128,N_4972,N_4777);
xnor U5129 (N_5129,N_4972,N_4772);
and U5130 (N_5130,N_4928,N_4996);
or U5131 (N_5131,N_4964,N_4920);
nand U5132 (N_5132,N_4879,N_4844);
and U5133 (N_5133,N_4907,N_4997);
nand U5134 (N_5134,N_4920,N_4903);
and U5135 (N_5135,N_4844,N_4875);
and U5136 (N_5136,N_4879,N_4773);
nand U5137 (N_5137,N_4967,N_4881);
or U5138 (N_5138,N_4780,N_4998);
xor U5139 (N_5139,N_4790,N_4809);
xor U5140 (N_5140,N_4987,N_4785);
or U5141 (N_5141,N_4892,N_4937);
xnor U5142 (N_5142,N_4840,N_4872);
or U5143 (N_5143,N_4774,N_4836);
or U5144 (N_5144,N_4822,N_4928);
nor U5145 (N_5145,N_4807,N_4754);
nand U5146 (N_5146,N_4857,N_4958);
and U5147 (N_5147,N_4822,N_4772);
and U5148 (N_5148,N_4864,N_4867);
or U5149 (N_5149,N_4978,N_4917);
nor U5150 (N_5150,N_4895,N_4984);
or U5151 (N_5151,N_4861,N_4947);
and U5152 (N_5152,N_4888,N_4865);
nand U5153 (N_5153,N_4980,N_4869);
xnor U5154 (N_5154,N_4776,N_4870);
nand U5155 (N_5155,N_4882,N_4851);
nand U5156 (N_5156,N_4764,N_4991);
nand U5157 (N_5157,N_4866,N_4761);
xnor U5158 (N_5158,N_4863,N_4924);
nor U5159 (N_5159,N_4785,N_4879);
nand U5160 (N_5160,N_4802,N_4868);
nand U5161 (N_5161,N_4799,N_4859);
or U5162 (N_5162,N_4838,N_4978);
nand U5163 (N_5163,N_4888,N_4780);
nor U5164 (N_5164,N_4851,N_4840);
nor U5165 (N_5165,N_4807,N_4780);
and U5166 (N_5166,N_4917,N_4806);
xor U5167 (N_5167,N_4787,N_4818);
xnor U5168 (N_5168,N_4819,N_4750);
and U5169 (N_5169,N_4949,N_4799);
and U5170 (N_5170,N_4989,N_4776);
or U5171 (N_5171,N_4979,N_4871);
xor U5172 (N_5172,N_4814,N_4875);
and U5173 (N_5173,N_4966,N_4984);
or U5174 (N_5174,N_4902,N_4873);
xnor U5175 (N_5175,N_4936,N_4865);
nand U5176 (N_5176,N_4790,N_4886);
or U5177 (N_5177,N_4928,N_4919);
nor U5178 (N_5178,N_4993,N_4768);
and U5179 (N_5179,N_4853,N_4890);
or U5180 (N_5180,N_4764,N_4932);
and U5181 (N_5181,N_4763,N_4815);
nand U5182 (N_5182,N_4937,N_4872);
nor U5183 (N_5183,N_4793,N_4834);
or U5184 (N_5184,N_4887,N_4848);
xor U5185 (N_5185,N_4913,N_4802);
or U5186 (N_5186,N_4972,N_4799);
nand U5187 (N_5187,N_4969,N_4797);
nand U5188 (N_5188,N_4773,N_4947);
nand U5189 (N_5189,N_4797,N_4979);
nor U5190 (N_5190,N_4858,N_4763);
xor U5191 (N_5191,N_4879,N_4823);
nor U5192 (N_5192,N_4912,N_4781);
nand U5193 (N_5193,N_4983,N_4985);
nor U5194 (N_5194,N_4998,N_4986);
or U5195 (N_5195,N_4983,N_4867);
or U5196 (N_5196,N_4782,N_4910);
or U5197 (N_5197,N_4868,N_4971);
nor U5198 (N_5198,N_4972,N_4790);
and U5199 (N_5199,N_4773,N_4933);
and U5200 (N_5200,N_4932,N_4852);
or U5201 (N_5201,N_4987,N_4963);
xor U5202 (N_5202,N_4832,N_4909);
nand U5203 (N_5203,N_4905,N_4910);
or U5204 (N_5204,N_4752,N_4910);
nand U5205 (N_5205,N_4984,N_4901);
or U5206 (N_5206,N_4997,N_4786);
and U5207 (N_5207,N_4857,N_4756);
nand U5208 (N_5208,N_4967,N_4939);
nor U5209 (N_5209,N_4964,N_4959);
nor U5210 (N_5210,N_4777,N_4951);
and U5211 (N_5211,N_4906,N_4915);
and U5212 (N_5212,N_4778,N_4940);
xnor U5213 (N_5213,N_4932,N_4822);
or U5214 (N_5214,N_4920,N_4796);
nor U5215 (N_5215,N_4771,N_4813);
or U5216 (N_5216,N_4767,N_4858);
xor U5217 (N_5217,N_4990,N_4899);
nor U5218 (N_5218,N_4818,N_4980);
nand U5219 (N_5219,N_4933,N_4944);
and U5220 (N_5220,N_4768,N_4775);
xor U5221 (N_5221,N_4833,N_4917);
or U5222 (N_5222,N_4776,N_4824);
nand U5223 (N_5223,N_4909,N_4888);
or U5224 (N_5224,N_4908,N_4837);
xnor U5225 (N_5225,N_4793,N_4782);
nor U5226 (N_5226,N_4967,N_4812);
or U5227 (N_5227,N_4896,N_4957);
nand U5228 (N_5228,N_4876,N_4902);
nand U5229 (N_5229,N_4765,N_4786);
or U5230 (N_5230,N_4818,N_4938);
and U5231 (N_5231,N_4774,N_4791);
xnor U5232 (N_5232,N_4760,N_4821);
xor U5233 (N_5233,N_4750,N_4820);
nand U5234 (N_5234,N_4889,N_4793);
and U5235 (N_5235,N_4865,N_4794);
xnor U5236 (N_5236,N_4806,N_4800);
xor U5237 (N_5237,N_4927,N_4795);
or U5238 (N_5238,N_4850,N_4856);
and U5239 (N_5239,N_4876,N_4815);
or U5240 (N_5240,N_4916,N_4822);
nand U5241 (N_5241,N_4843,N_4976);
and U5242 (N_5242,N_4888,N_4985);
nor U5243 (N_5243,N_4843,N_4880);
and U5244 (N_5244,N_4790,N_4814);
or U5245 (N_5245,N_4875,N_4982);
or U5246 (N_5246,N_4927,N_4861);
and U5247 (N_5247,N_4928,N_4911);
and U5248 (N_5248,N_4928,N_4784);
or U5249 (N_5249,N_4830,N_4973);
and U5250 (N_5250,N_5074,N_5172);
xnor U5251 (N_5251,N_5020,N_5230);
nand U5252 (N_5252,N_5058,N_5221);
and U5253 (N_5253,N_5076,N_5166);
nand U5254 (N_5254,N_5144,N_5165);
nor U5255 (N_5255,N_5012,N_5003);
or U5256 (N_5256,N_5085,N_5023);
and U5257 (N_5257,N_5130,N_5041);
or U5258 (N_5258,N_5061,N_5121);
xor U5259 (N_5259,N_5186,N_5245);
nor U5260 (N_5260,N_5071,N_5202);
nand U5261 (N_5261,N_5248,N_5086);
or U5262 (N_5262,N_5180,N_5123);
xnor U5263 (N_5263,N_5214,N_5191);
nor U5264 (N_5264,N_5000,N_5001);
or U5265 (N_5265,N_5146,N_5153);
nand U5266 (N_5266,N_5068,N_5196);
and U5267 (N_5267,N_5239,N_5022);
xnor U5268 (N_5268,N_5195,N_5216);
xor U5269 (N_5269,N_5065,N_5060);
and U5270 (N_5270,N_5133,N_5229);
or U5271 (N_5271,N_5181,N_5072);
or U5272 (N_5272,N_5122,N_5155);
or U5273 (N_5273,N_5188,N_5050);
or U5274 (N_5274,N_5114,N_5049);
and U5275 (N_5275,N_5203,N_5167);
nand U5276 (N_5276,N_5128,N_5009);
xor U5277 (N_5277,N_5235,N_5227);
or U5278 (N_5278,N_5150,N_5025);
xor U5279 (N_5279,N_5207,N_5168);
xor U5280 (N_5280,N_5142,N_5113);
and U5281 (N_5281,N_5234,N_5002);
nor U5282 (N_5282,N_5140,N_5206);
and U5283 (N_5283,N_5115,N_5069);
nand U5284 (N_5284,N_5147,N_5097);
and U5285 (N_5285,N_5034,N_5190);
xnor U5286 (N_5286,N_5033,N_5213);
or U5287 (N_5287,N_5127,N_5094);
xor U5288 (N_5288,N_5228,N_5079);
nand U5289 (N_5289,N_5056,N_5212);
nor U5290 (N_5290,N_5151,N_5176);
or U5291 (N_5291,N_5192,N_5178);
nor U5292 (N_5292,N_5028,N_5105);
nor U5293 (N_5293,N_5117,N_5044);
nor U5294 (N_5294,N_5054,N_5047);
or U5295 (N_5295,N_5108,N_5048);
nor U5296 (N_5296,N_5126,N_5057);
nand U5297 (N_5297,N_5204,N_5243);
xor U5298 (N_5298,N_5132,N_5073);
nand U5299 (N_5299,N_5083,N_5030);
or U5300 (N_5300,N_5036,N_5016);
and U5301 (N_5301,N_5184,N_5218);
xor U5302 (N_5302,N_5116,N_5141);
xnor U5303 (N_5303,N_5021,N_5118);
xnor U5304 (N_5304,N_5004,N_5156);
or U5305 (N_5305,N_5055,N_5242);
nand U5306 (N_5306,N_5125,N_5160);
nand U5307 (N_5307,N_5201,N_5032);
nor U5308 (N_5308,N_5019,N_5088);
nor U5309 (N_5309,N_5042,N_5062);
nand U5310 (N_5310,N_5171,N_5075);
xor U5311 (N_5311,N_5200,N_5208);
nor U5312 (N_5312,N_5159,N_5182);
or U5313 (N_5313,N_5026,N_5135);
xor U5314 (N_5314,N_5029,N_5226);
nor U5315 (N_5315,N_5219,N_5194);
nor U5316 (N_5316,N_5015,N_5189);
and U5317 (N_5317,N_5005,N_5149);
and U5318 (N_5318,N_5037,N_5137);
or U5319 (N_5319,N_5090,N_5067);
and U5320 (N_5320,N_5010,N_5110);
and U5321 (N_5321,N_5080,N_5244);
nor U5322 (N_5322,N_5145,N_5222);
or U5323 (N_5323,N_5024,N_5120);
and U5324 (N_5324,N_5119,N_5233);
nand U5325 (N_5325,N_5231,N_5078);
nor U5326 (N_5326,N_5092,N_5082);
nand U5327 (N_5327,N_5236,N_5046);
and U5328 (N_5328,N_5169,N_5193);
xnor U5329 (N_5329,N_5089,N_5014);
and U5330 (N_5330,N_5084,N_5205);
nor U5331 (N_5331,N_5249,N_5102);
or U5332 (N_5332,N_5158,N_5013);
nand U5333 (N_5333,N_5164,N_5098);
or U5334 (N_5334,N_5246,N_5031);
or U5335 (N_5335,N_5209,N_5225);
and U5336 (N_5336,N_5099,N_5104);
nor U5337 (N_5337,N_5087,N_5232);
and U5338 (N_5338,N_5174,N_5198);
nand U5339 (N_5339,N_5011,N_5129);
xor U5340 (N_5340,N_5143,N_5100);
nand U5341 (N_5341,N_5177,N_5138);
nor U5342 (N_5342,N_5109,N_5134);
and U5343 (N_5343,N_5008,N_5240);
nand U5344 (N_5344,N_5101,N_5211);
nand U5345 (N_5345,N_5081,N_5111);
and U5346 (N_5346,N_5106,N_5199);
xnor U5347 (N_5347,N_5224,N_5241);
nand U5348 (N_5348,N_5131,N_5007);
xnor U5349 (N_5349,N_5051,N_5053);
nor U5350 (N_5350,N_5093,N_5043);
or U5351 (N_5351,N_5035,N_5066);
nand U5352 (N_5352,N_5139,N_5170);
and U5353 (N_5353,N_5237,N_5185);
or U5354 (N_5354,N_5157,N_5070);
and U5355 (N_5355,N_5210,N_5238);
nor U5356 (N_5356,N_5173,N_5148);
or U5357 (N_5357,N_5175,N_5027);
xnor U5358 (N_5358,N_5045,N_5040);
nand U5359 (N_5359,N_5161,N_5038);
and U5360 (N_5360,N_5039,N_5152);
or U5361 (N_5361,N_5215,N_5064);
nand U5362 (N_5362,N_5077,N_5247);
xnor U5363 (N_5363,N_5063,N_5103);
xor U5364 (N_5364,N_5136,N_5223);
and U5365 (N_5365,N_5220,N_5197);
nand U5366 (N_5366,N_5124,N_5183);
nand U5367 (N_5367,N_5163,N_5018);
xor U5368 (N_5368,N_5091,N_5006);
nor U5369 (N_5369,N_5107,N_5217);
nor U5370 (N_5370,N_5179,N_5017);
nor U5371 (N_5371,N_5112,N_5154);
and U5372 (N_5372,N_5162,N_5059);
and U5373 (N_5373,N_5096,N_5187);
xor U5374 (N_5374,N_5095,N_5052);
or U5375 (N_5375,N_5222,N_5056);
and U5376 (N_5376,N_5106,N_5056);
or U5377 (N_5377,N_5091,N_5036);
nor U5378 (N_5378,N_5195,N_5115);
or U5379 (N_5379,N_5165,N_5126);
and U5380 (N_5380,N_5245,N_5118);
xor U5381 (N_5381,N_5079,N_5033);
xor U5382 (N_5382,N_5063,N_5023);
xor U5383 (N_5383,N_5183,N_5068);
or U5384 (N_5384,N_5037,N_5033);
or U5385 (N_5385,N_5189,N_5218);
and U5386 (N_5386,N_5192,N_5114);
nor U5387 (N_5387,N_5116,N_5125);
nand U5388 (N_5388,N_5077,N_5184);
and U5389 (N_5389,N_5239,N_5165);
xnor U5390 (N_5390,N_5235,N_5097);
or U5391 (N_5391,N_5122,N_5058);
nand U5392 (N_5392,N_5188,N_5207);
xnor U5393 (N_5393,N_5119,N_5026);
and U5394 (N_5394,N_5210,N_5090);
xnor U5395 (N_5395,N_5185,N_5083);
nand U5396 (N_5396,N_5182,N_5249);
or U5397 (N_5397,N_5066,N_5077);
xor U5398 (N_5398,N_5155,N_5021);
nor U5399 (N_5399,N_5169,N_5239);
nor U5400 (N_5400,N_5206,N_5003);
xor U5401 (N_5401,N_5152,N_5227);
xor U5402 (N_5402,N_5098,N_5102);
xor U5403 (N_5403,N_5069,N_5003);
nor U5404 (N_5404,N_5135,N_5179);
and U5405 (N_5405,N_5179,N_5127);
or U5406 (N_5406,N_5213,N_5026);
and U5407 (N_5407,N_5032,N_5042);
and U5408 (N_5408,N_5169,N_5026);
or U5409 (N_5409,N_5188,N_5093);
nand U5410 (N_5410,N_5227,N_5057);
nor U5411 (N_5411,N_5187,N_5197);
xnor U5412 (N_5412,N_5215,N_5112);
nor U5413 (N_5413,N_5188,N_5143);
xor U5414 (N_5414,N_5092,N_5017);
xor U5415 (N_5415,N_5183,N_5028);
xor U5416 (N_5416,N_5095,N_5132);
nand U5417 (N_5417,N_5132,N_5194);
and U5418 (N_5418,N_5072,N_5076);
nor U5419 (N_5419,N_5160,N_5107);
and U5420 (N_5420,N_5094,N_5170);
or U5421 (N_5421,N_5146,N_5151);
xor U5422 (N_5422,N_5207,N_5014);
and U5423 (N_5423,N_5053,N_5064);
and U5424 (N_5424,N_5090,N_5104);
or U5425 (N_5425,N_5024,N_5022);
nand U5426 (N_5426,N_5161,N_5225);
and U5427 (N_5427,N_5137,N_5048);
and U5428 (N_5428,N_5189,N_5032);
xnor U5429 (N_5429,N_5115,N_5190);
or U5430 (N_5430,N_5210,N_5059);
and U5431 (N_5431,N_5103,N_5153);
xnor U5432 (N_5432,N_5081,N_5097);
and U5433 (N_5433,N_5203,N_5111);
xnor U5434 (N_5434,N_5125,N_5208);
nand U5435 (N_5435,N_5053,N_5241);
and U5436 (N_5436,N_5168,N_5081);
nor U5437 (N_5437,N_5137,N_5093);
nand U5438 (N_5438,N_5058,N_5242);
nand U5439 (N_5439,N_5061,N_5092);
xnor U5440 (N_5440,N_5157,N_5111);
xnor U5441 (N_5441,N_5014,N_5072);
nor U5442 (N_5442,N_5032,N_5071);
nor U5443 (N_5443,N_5207,N_5233);
nor U5444 (N_5444,N_5165,N_5046);
or U5445 (N_5445,N_5172,N_5185);
nor U5446 (N_5446,N_5175,N_5060);
xor U5447 (N_5447,N_5052,N_5235);
and U5448 (N_5448,N_5196,N_5071);
nor U5449 (N_5449,N_5079,N_5198);
xnor U5450 (N_5450,N_5233,N_5204);
nand U5451 (N_5451,N_5207,N_5048);
and U5452 (N_5452,N_5049,N_5098);
or U5453 (N_5453,N_5140,N_5094);
and U5454 (N_5454,N_5126,N_5047);
nor U5455 (N_5455,N_5126,N_5105);
nor U5456 (N_5456,N_5125,N_5242);
nand U5457 (N_5457,N_5099,N_5138);
nor U5458 (N_5458,N_5191,N_5010);
nand U5459 (N_5459,N_5126,N_5006);
nor U5460 (N_5460,N_5241,N_5209);
nand U5461 (N_5461,N_5029,N_5093);
nor U5462 (N_5462,N_5176,N_5136);
and U5463 (N_5463,N_5038,N_5034);
or U5464 (N_5464,N_5219,N_5166);
and U5465 (N_5465,N_5133,N_5172);
xor U5466 (N_5466,N_5070,N_5042);
nor U5467 (N_5467,N_5119,N_5098);
xnor U5468 (N_5468,N_5070,N_5052);
and U5469 (N_5469,N_5035,N_5023);
or U5470 (N_5470,N_5118,N_5146);
xnor U5471 (N_5471,N_5090,N_5036);
xnor U5472 (N_5472,N_5200,N_5221);
nor U5473 (N_5473,N_5214,N_5183);
or U5474 (N_5474,N_5011,N_5186);
xor U5475 (N_5475,N_5137,N_5235);
or U5476 (N_5476,N_5031,N_5068);
nand U5477 (N_5477,N_5214,N_5143);
nand U5478 (N_5478,N_5041,N_5004);
or U5479 (N_5479,N_5076,N_5197);
and U5480 (N_5480,N_5031,N_5102);
or U5481 (N_5481,N_5170,N_5058);
nand U5482 (N_5482,N_5011,N_5175);
xnor U5483 (N_5483,N_5220,N_5012);
xor U5484 (N_5484,N_5041,N_5061);
xor U5485 (N_5485,N_5125,N_5187);
nand U5486 (N_5486,N_5215,N_5167);
or U5487 (N_5487,N_5084,N_5103);
or U5488 (N_5488,N_5080,N_5019);
xnor U5489 (N_5489,N_5176,N_5082);
nor U5490 (N_5490,N_5198,N_5103);
or U5491 (N_5491,N_5009,N_5235);
or U5492 (N_5492,N_5147,N_5221);
and U5493 (N_5493,N_5233,N_5146);
xor U5494 (N_5494,N_5122,N_5148);
nor U5495 (N_5495,N_5078,N_5113);
and U5496 (N_5496,N_5125,N_5077);
and U5497 (N_5497,N_5157,N_5005);
or U5498 (N_5498,N_5073,N_5100);
or U5499 (N_5499,N_5135,N_5037);
and U5500 (N_5500,N_5395,N_5335);
xnor U5501 (N_5501,N_5346,N_5272);
nand U5502 (N_5502,N_5455,N_5258);
and U5503 (N_5503,N_5453,N_5317);
nor U5504 (N_5504,N_5374,N_5494);
nand U5505 (N_5505,N_5408,N_5467);
nand U5506 (N_5506,N_5368,N_5423);
and U5507 (N_5507,N_5431,N_5473);
xor U5508 (N_5508,N_5313,N_5281);
and U5509 (N_5509,N_5273,N_5259);
nand U5510 (N_5510,N_5367,N_5338);
nor U5511 (N_5511,N_5432,N_5369);
xor U5512 (N_5512,N_5268,N_5309);
or U5513 (N_5513,N_5483,N_5470);
and U5514 (N_5514,N_5278,N_5458);
and U5515 (N_5515,N_5400,N_5486);
xor U5516 (N_5516,N_5437,N_5306);
nand U5517 (N_5517,N_5439,N_5420);
nor U5518 (N_5518,N_5255,N_5354);
or U5519 (N_5519,N_5448,N_5436);
nand U5520 (N_5520,N_5305,N_5474);
nor U5521 (N_5521,N_5460,N_5490);
nor U5522 (N_5522,N_5496,N_5330);
or U5523 (N_5523,N_5489,N_5493);
and U5524 (N_5524,N_5347,N_5375);
nand U5525 (N_5525,N_5307,N_5271);
xor U5526 (N_5526,N_5434,N_5397);
and U5527 (N_5527,N_5454,N_5333);
nand U5528 (N_5528,N_5315,N_5343);
or U5529 (N_5529,N_5482,N_5485);
nor U5530 (N_5530,N_5326,N_5320);
or U5531 (N_5531,N_5390,N_5355);
and U5532 (N_5532,N_5344,N_5261);
nand U5533 (N_5533,N_5352,N_5287);
nand U5534 (N_5534,N_5364,N_5481);
nand U5535 (N_5535,N_5282,N_5414);
xor U5536 (N_5536,N_5475,N_5440);
nand U5537 (N_5537,N_5379,N_5464);
or U5538 (N_5538,N_5283,N_5366);
or U5539 (N_5539,N_5331,N_5394);
nor U5540 (N_5540,N_5340,N_5263);
and U5541 (N_5541,N_5457,N_5280);
or U5542 (N_5542,N_5294,N_5362);
nand U5543 (N_5543,N_5363,N_5348);
xnor U5544 (N_5544,N_5292,N_5495);
xnor U5545 (N_5545,N_5372,N_5386);
nand U5546 (N_5546,N_5252,N_5334);
nor U5547 (N_5547,N_5336,N_5266);
or U5548 (N_5548,N_5312,N_5472);
xnor U5549 (N_5549,N_5304,N_5484);
xor U5550 (N_5550,N_5288,N_5446);
or U5551 (N_5551,N_5382,N_5416);
nor U5552 (N_5552,N_5430,N_5498);
or U5553 (N_5553,N_5497,N_5418);
or U5554 (N_5554,N_5279,N_5264);
xnor U5555 (N_5555,N_5341,N_5276);
and U5556 (N_5556,N_5398,N_5396);
or U5557 (N_5557,N_5297,N_5479);
xor U5558 (N_5558,N_5452,N_5492);
xor U5559 (N_5559,N_5303,N_5253);
nor U5560 (N_5560,N_5353,N_5421);
and U5561 (N_5561,N_5403,N_5322);
nor U5562 (N_5562,N_5302,N_5260);
and U5563 (N_5563,N_5441,N_5293);
and U5564 (N_5564,N_5433,N_5257);
nor U5565 (N_5565,N_5373,N_5449);
nand U5566 (N_5566,N_5291,N_5387);
nor U5567 (N_5567,N_5422,N_5314);
nor U5568 (N_5568,N_5357,N_5296);
and U5569 (N_5569,N_5351,N_5356);
nor U5570 (N_5570,N_5383,N_5254);
xnor U5571 (N_5571,N_5413,N_5378);
xnor U5572 (N_5572,N_5465,N_5405);
nand U5573 (N_5573,N_5299,N_5381);
and U5574 (N_5574,N_5274,N_5438);
xnor U5575 (N_5575,N_5251,N_5435);
nand U5576 (N_5576,N_5318,N_5417);
nor U5577 (N_5577,N_5419,N_5447);
xor U5578 (N_5578,N_5319,N_5298);
xnor U5579 (N_5579,N_5345,N_5385);
nor U5580 (N_5580,N_5407,N_5443);
nor U5581 (N_5581,N_5332,N_5342);
nor U5582 (N_5582,N_5462,N_5265);
xnor U5583 (N_5583,N_5262,N_5308);
nor U5584 (N_5584,N_5339,N_5269);
nor U5585 (N_5585,N_5412,N_5286);
xor U5586 (N_5586,N_5456,N_5471);
and U5587 (N_5587,N_5444,N_5337);
nand U5588 (N_5588,N_5327,N_5359);
xnor U5589 (N_5589,N_5350,N_5329);
nand U5590 (N_5590,N_5445,N_5380);
and U5591 (N_5591,N_5415,N_5360);
and U5592 (N_5592,N_5428,N_5476);
and U5593 (N_5593,N_5424,N_5384);
nor U5594 (N_5594,N_5323,N_5451);
nor U5595 (N_5595,N_5404,N_5477);
or U5596 (N_5596,N_5425,N_5411);
xor U5597 (N_5597,N_5328,N_5461);
nor U5598 (N_5598,N_5361,N_5371);
or U5599 (N_5599,N_5488,N_5325);
nand U5600 (N_5600,N_5300,N_5377);
xnor U5601 (N_5601,N_5256,N_5469);
or U5602 (N_5602,N_5402,N_5410);
nor U5603 (N_5603,N_5478,N_5316);
and U5604 (N_5604,N_5285,N_5267);
or U5605 (N_5605,N_5289,N_5376);
and U5606 (N_5606,N_5450,N_5349);
and U5607 (N_5607,N_5391,N_5409);
nand U5608 (N_5608,N_5370,N_5499);
and U5609 (N_5609,N_5310,N_5321);
or U5610 (N_5610,N_5392,N_5284);
or U5611 (N_5611,N_5480,N_5388);
or U5612 (N_5612,N_5277,N_5270);
nor U5613 (N_5613,N_5406,N_5393);
nor U5614 (N_5614,N_5459,N_5301);
nor U5615 (N_5615,N_5358,N_5250);
xor U5616 (N_5616,N_5401,N_5491);
nand U5617 (N_5617,N_5427,N_5365);
xnor U5618 (N_5618,N_5426,N_5389);
nor U5619 (N_5619,N_5429,N_5463);
xnor U5620 (N_5620,N_5468,N_5311);
or U5621 (N_5621,N_5324,N_5290);
or U5622 (N_5622,N_5487,N_5442);
and U5623 (N_5623,N_5466,N_5295);
and U5624 (N_5624,N_5399,N_5275);
nor U5625 (N_5625,N_5287,N_5397);
nor U5626 (N_5626,N_5427,N_5481);
nand U5627 (N_5627,N_5339,N_5377);
or U5628 (N_5628,N_5465,N_5355);
and U5629 (N_5629,N_5274,N_5491);
nand U5630 (N_5630,N_5440,N_5374);
nor U5631 (N_5631,N_5259,N_5370);
and U5632 (N_5632,N_5251,N_5480);
or U5633 (N_5633,N_5314,N_5327);
and U5634 (N_5634,N_5492,N_5423);
nor U5635 (N_5635,N_5283,N_5481);
and U5636 (N_5636,N_5441,N_5287);
or U5637 (N_5637,N_5271,N_5335);
nor U5638 (N_5638,N_5278,N_5481);
nand U5639 (N_5639,N_5297,N_5496);
xor U5640 (N_5640,N_5287,N_5313);
nor U5641 (N_5641,N_5294,N_5485);
or U5642 (N_5642,N_5342,N_5309);
xor U5643 (N_5643,N_5428,N_5250);
nand U5644 (N_5644,N_5403,N_5252);
or U5645 (N_5645,N_5416,N_5362);
and U5646 (N_5646,N_5465,N_5334);
nand U5647 (N_5647,N_5352,N_5464);
xnor U5648 (N_5648,N_5411,N_5460);
or U5649 (N_5649,N_5269,N_5415);
nand U5650 (N_5650,N_5377,N_5331);
nand U5651 (N_5651,N_5427,N_5359);
nand U5652 (N_5652,N_5487,N_5277);
xnor U5653 (N_5653,N_5352,N_5358);
nor U5654 (N_5654,N_5311,N_5338);
or U5655 (N_5655,N_5439,N_5485);
xor U5656 (N_5656,N_5312,N_5284);
or U5657 (N_5657,N_5346,N_5424);
nor U5658 (N_5658,N_5492,N_5298);
xnor U5659 (N_5659,N_5394,N_5344);
and U5660 (N_5660,N_5482,N_5397);
or U5661 (N_5661,N_5356,N_5257);
and U5662 (N_5662,N_5282,N_5296);
nand U5663 (N_5663,N_5337,N_5289);
and U5664 (N_5664,N_5395,N_5330);
and U5665 (N_5665,N_5463,N_5326);
nor U5666 (N_5666,N_5259,N_5409);
xnor U5667 (N_5667,N_5285,N_5284);
or U5668 (N_5668,N_5482,N_5272);
or U5669 (N_5669,N_5416,N_5481);
and U5670 (N_5670,N_5291,N_5463);
or U5671 (N_5671,N_5386,N_5453);
nand U5672 (N_5672,N_5400,N_5477);
xnor U5673 (N_5673,N_5423,N_5496);
xnor U5674 (N_5674,N_5259,N_5381);
nor U5675 (N_5675,N_5320,N_5455);
nor U5676 (N_5676,N_5436,N_5468);
or U5677 (N_5677,N_5254,N_5329);
or U5678 (N_5678,N_5258,N_5337);
nand U5679 (N_5679,N_5324,N_5350);
and U5680 (N_5680,N_5367,N_5422);
nand U5681 (N_5681,N_5318,N_5397);
nor U5682 (N_5682,N_5403,N_5315);
nor U5683 (N_5683,N_5272,N_5366);
nor U5684 (N_5684,N_5256,N_5317);
nor U5685 (N_5685,N_5270,N_5283);
and U5686 (N_5686,N_5254,N_5297);
or U5687 (N_5687,N_5366,N_5342);
or U5688 (N_5688,N_5439,N_5373);
nand U5689 (N_5689,N_5385,N_5422);
and U5690 (N_5690,N_5363,N_5365);
nand U5691 (N_5691,N_5281,N_5260);
nor U5692 (N_5692,N_5282,N_5292);
nor U5693 (N_5693,N_5428,N_5326);
xnor U5694 (N_5694,N_5432,N_5282);
or U5695 (N_5695,N_5376,N_5430);
and U5696 (N_5696,N_5335,N_5305);
nor U5697 (N_5697,N_5357,N_5381);
xnor U5698 (N_5698,N_5381,N_5454);
or U5699 (N_5699,N_5463,N_5431);
nor U5700 (N_5700,N_5261,N_5321);
and U5701 (N_5701,N_5455,N_5374);
xnor U5702 (N_5702,N_5400,N_5280);
or U5703 (N_5703,N_5418,N_5493);
xnor U5704 (N_5704,N_5463,N_5396);
and U5705 (N_5705,N_5352,N_5448);
xnor U5706 (N_5706,N_5288,N_5281);
xnor U5707 (N_5707,N_5358,N_5414);
nand U5708 (N_5708,N_5428,N_5267);
or U5709 (N_5709,N_5369,N_5377);
or U5710 (N_5710,N_5256,N_5325);
xnor U5711 (N_5711,N_5448,N_5466);
or U5712 (N_5712,N_5309,N_5345);
or U5713 (N_5713,N_5403,N_5312);
nand U5714 (N_5714,N_5278,N_5381);
or U5715 (N_5715,N_5278,N_5350);
nand U5716 (N_5716,N_5320,N_5410);
and U5717 (N_5717,N_5429,N_5327);
nand U5718 (N_5718,N_5445,N_5281);
nand U5719 (N_5719,N_5354,N_5479);
nand U5720 (N_5720,N_5367,N_5466);
xnor U5721 (N_5721,N_5316,N_5487);
xnor U5722 (N_5722,N_5291,N_5449);
or U5723 (N_5723,N_5496,N_5497);
nand U5724 (N_5724,N_5301,N_5350);
nand U5725 (N_5725,N_5311,N_5302);
nor U5726 (N_5726,N_5483,N_5276);
nor U5727 (N_5727,N_5295,N_5349);
nor U5728 (N_5728,N_5498,N_5274);
xor U5729 (N_5729,N_5281,N_5497);
or U5730 (N_5730,N_5417,N_5474);
xor U5731 (N_5731,N_5253,N_5483);
nor U5732 (N_5732,N_5477,N_5327);
nor U5733 (N_5733,N_5485,N_5287);
nand U5734 (N_5734,N_5497,N_5273);
nor U5735 (N_5735,N_5358,N_5428);
nand U5736 (N_5736,N_5478,N_5473);
and U5737 (N_5737,N_5265,N_5430);
xnor U5738 (N_5738,N_5370,N_5330);
or U5739 (N_5739,N_5316,N_5350);
nor U5740 (N_5740,N_5303,N_5412);
or U5741 (N_5741,N_5480,N_5296);
and U5742 (N_5742,N_5478,N_5450);
xnor U5743 (N_5743,N_5262,N_5343);
nand U5744 (N_5744,N_5287,N_5435);
nor U5745 (N_5745,N_5300,N_5419);
nor U5746 (N_5746,N_5327,N_5342);
or U5747 (N_5747,N_5465,N_5365);
or U5748 (N_5748,N_5424,N_5297);
and U5749 (N_5749,N_5273,N_5371);
xor U5750 (N_5750,N_5564,N_5555);
and U5751 (N_5751,N_5572,N_5645);
and U5752 (N_5752,N_5718,N_5568);
or U5753 (N_5753,N_5708,N_5730);
or U5754 (N_5754,N_5558,N_5578);
and U5755 (N_5755,N_5683,N_5732);
and U5756 (N_5756,N_5518,N_5616);
xor U5757 (N_5757,N_5501,N_5550);
nor U5758 (N_5758,N_5687,N_5722);
nor U5759 (N_5759,N_5695,N_5570);
xor U5760 (N_5760,N_5562,N_5652);
nor U5761 (N_5761,N_5694,N_5638);
xnor U5762 (N_5762,N_5603,N_5509);
xor U5763 (N_5763,N_5690,N_5736);
nor U5764 (N_5764,N_5662,N_5704);
nand U5765 (N_5765,N_5644,N_5681);
and U5766 (N_5766,N_5677,N_5620);
xnor U5767 (N_5767,N_5686,N_5553);
and U5768 (N_5768,N_5520,N_5716);
and U5769 (N_5769,N_5503,N_5675);
xor U5770 (N_5770,N_5531,N_5549);
and U5771 (N_5771,N_5612,N_5684);
nor U5772 (N_5772,N_5571,N_5559);
and U5773 (N_5773,N_5614,N_5592);
nand U5774 (N_5774,N_5523,N_5532);
xor U5775 (N_5775,N_5679,N_5586);
nand U5776 (N_5776,N_5604,N_5545);
or U5777 (N_5777,N_5726,N_5729);
and U5778 (N_5778,N_5733,N_5670);
nor U5779 (N_5779,N_5575,N_5554);
and U5780 (N_5780,N_5541,N_5655);
or U5781 (N_5781,N_5594,N_5623);
xor U5782 (N_5782,N_5551,N_5714);
xor U5783 (N_5783,N_5715,N_5719);
or U5784 (N_5784,N_5626,N_5691);
or U5785 (N_5785,N_5745,N_5688);
nor U5786 (N_5786,N_5643,N_5622);
or U5787 (N_5787,N_5500,N_5569);
or U5788 (N_5788,N_5513,N_5640);
nand U5789 (N_5789,N_5693,N_5613);
xor U5790 (N_5790,N_5740,N_5560);
or U5791 (N_5791,N_5573,N_5508);
and U5792 (N_5792,N_5649,N_5596);
nand U5793 (N_5793,N_5577,N_5583);
nand U5794 (N_5794,N_5516,N_5534);
nand U5795 (N_5795,N_5672,N_5618);
nand U5796 (N_5796,N_5595,N_5701);
and U5797 (N_5797,N_5741,N_5685);
and U5798 (N_5798,N_5657,N_5746);
nand U5799 (N_5799,N_5666,N_5710);
nor U5800 (N_5800,N_5744,N_5610);
xor U5801 (N_5801,N_5705,N_5642);
xor U5802 (N_5802,N_5712,N_5630);
nand U5803 (N_5803,N_5576,N_5526);
nor U5804 (N_5804,N_5738,N_5661);
xor U5805 (N_5805,N_5692,N_5678);
nor U5806 (N_5806,N_5663,N_5561);
nand U5807 (N_5807,N_5535,N_5632);
xnor U5808 (N_5808,N_5607,N_5689);
nand U5809 (N_5809,N_5742,N_5581);
and U5810 (N_5810,N_5707,N_5627);
or U5811 (N_5811,N_5522,N_5720);
or U5812 (N_5812,N_5566,N_5636);
and U5813 (N_5813,N_5668,N_5665);
xnor U5814 (N_5814,N_5608,N_5533);
and U5815 (N_5815,N_5727,N_5669);
or U5816 (N_5816,N_5739,N_5556);
xor U5817 (N_5817,N_5629,N_5506);
or U5818 (N_5818,N_5599,N_5605);
and U5819 (N_5819,N_5725,N_5749);
and U5820 (N_5820,N_5567,N_5747);
and U5821 (N_5821,N_5624,N_5651);
nand U5822 (N_5822,N_5656,N_5696);
nor U5823 (N_5823,N_5621,N_5593);
or U5824 (N_5824,N_5542,N_5505);
xnor U5825 (N_5825,N_5682,N_5588);
nand U5826 (N_5826,N_5600,N_5552);
nor U5827 (N_5827,N_5667,N_5702);
or U5828 (N_5828,N_5557,N_5734);
nor U5829 (N_5829,N_5584,N_5641);
or U5830 (N_5830,N_5671,N_5680);
xnor U5831 (N_5831,N_5648,N_5524);
or U5832 (N_5832,N_5606,N_5538);
nand U5833 (N_5833,N_5664,N_5658);
nand U5834 (N_5834,N_5619,N_5609);
nand U5835 (N_5835,N_5547,N_5515);
and U5836 (N_5836,N_5543,N_5674);
or U5837 (N_5837,N_5536,N_5717);
xor U5838 (N_5838,N_5529,N_5628);
xor U5839 (N_5839,N_5659,N_5574);
nand U5840 (N_5840,N_5709,N_5580);
and U5841 (N_5841,N_5540,N_5611);
nor U5842 (N_5842,N_5723,N_5527);
or U5843 (N_5843,N_5637,N_5519);
xor U5844 (N_5844,N_5579,N_5582);
and U5845 (N_5845,N_5530,N_5617);
nor U5846 (N_5846,N_5502,N_5563);
nor U5847 (N_5847,N_5512,N_5589);
nor U5848 (N_5848,N_5737,N_5703);
and U5849 (N_5849,N_5521,N_5634);
nand U5850 (N_5850,N_5631,N_5673);
or U5851 (N_5851,N_5615,N_5591);
nand U5852 (N_5852,N_5546,N_5653);
and U5853 (N_5853,N_5700,N_5698);
and U5854 (N_5854,N_5706,N_5625);
and U5855 (N_5855,N_5654,N_5539);
nand U5856 (N_5856,N_5711,N_5504);
nor U5857 (N_5857,N_5528,N_5676);
nand U5858 (N_5858,N_5735,N_5660);
or U5859 (N_5859,N_5514,N_5635);
nand U5860 (N_5860,N_5544,N_5525);
or U5861 (N_5861,N_5507,N_5748);
or U5862 (N_5862,N_5650,N_5743);
or U5863 (N_5863,N_5565,N_5601);
or U5864 (N_5864,N_5699,N_5510);
or U5865 (N_5865,N_5590,N_5517);
nor U5866 (N_5866,N_5731,N_5721);
or U5867 (N_5867,N_5647,N_5598);
xnor U5868 (N_5868,N_5597,N_5713);
and U5869 (N_5869,N_5602,N_5639);
nand U5870 (N_5870,N_5511,N_5548);
xnor U5871 (N_5871,N_5587,N_5697);
nand U5872 (N_5872,N_5633,N_5646);
xor U5873 (N_5873,N_5537,N_5728);
nand U5874 (N_5874,N_5585,N_5724);
nand U5875 (N_5875,N_5603,N_5746);
and U5876 (N_5876,N_5540,N_5621);
nand U5877 (N_5877,N_5682,N_5576);
nand U5878 (N_5878,N_5590,N_5602);
or U5879 (N_5879,N_5599,N_5588);
nor U5880 (N_5880,N_5518,N_5601);
nor U5881 (N_5881,N_5558,N_5530);
xnor U5882 (N_5882,N_5627,N_5639);
nor U5883 (N_5883,N_5513,N_5514);
or U5884 (N_5884,N_5741,N_5573);
and U5885 (N_5885,N_5606,N_5703);
nand U5886 (N_5886,N_5706,N_5650);
nor U5887 (N_5887,N_5746,N_5572);
nand U5888 (N_5888,N_5533,N_5504);
or U5889 (N_5889,N_5627,N_5592);
nand U5890 (N_5890,N_5594,N_5746);
nand U5891 (N_5891,N_5502,N_5537);
nor U5892 (N_5892,N_5703,N_5687);
and U5893 (N_5893,N_5558,N_5710);
nor U5894 (N_5894,N_5501,N_5686);
and U5895 (N_5895,N_5594,N_5516);
or U5896 (N_5896,N_5674,N_5713);
and U5897 (N_5897,N_5554,N_5522);
nand U5898 (N_5898,N_5637,N_5551);
or U5899 (N_5899,N_5519,N_5538);
xor U5900 (N_5900,N_5668,N_5554);
or U5901 (N_5901,N_5500,N_5559);
nand U5902 (N_5902,N_5723,N_5660);
or U5903 (N_5903,N_5534,N_5535);
or U5904 (N_5904,N_5662,N_5649);
or U5905 (N_5905,N_5674,N_5684);
xor U5906 (N_5906,N_5563,N_5640);
or U5907 (N_5907,N_5705,N_5534);
or U5908 (N_5908,N_5668,N_5647);
nor U5909 (N_5909,N_5579,N_5690);
nor U5910 (N_5910,N_5652,N_5520);
xor U5911 (N_5911,N_5601,N_5626);
nor U5912 (N_5912,N_5649,N_5689);
or U5913 (N_5913,N_5706,N_5737);
nand U5914 (N_5914,N_5741,N_5564);
nand U5915 (N_5915,N_5705,N_5748);
nand U5916 (N_5916,N_5740,N_5588);
nor U5917 (N_5917,N_5563,N_5527);
and U5918 (N_5918,N_5571,N_5717);
nand U5919 (N_5919,N_5600,N_5634);
xnor U5920 (N_5920,N_5691,N_5576);
and U5921 (N_5921,N_5617,N_5645);
nand U5922 (N_5922,N_5660,N_5606);
xor U5923 (N_5923,N_5692,N_5631);
nor U5924 (N_5924,N_5703,N_5712);
and U5925 (N_5925,N_5736,N_5696);
xor U5926 (N_5926,N_5717,N_5721);
nor U5927 (N_5927,N_5560,N_5616);
or U5928 (N_5928,N_5731,N_5629);
nor U5929 (N_5929,N_5618,N_5670);
and U5930 (N_5930,N_5596,N_5660);
or U5931 (N_5931,N_5679,N_5538);
nor U5932 (N_5932,N_5527,N_5575);
nor U5933 (N_5933,N_5595,N_5597);
and U5934 (N_5934,N_5603,N_5530);
nand U5935 (N_5935,N_5547,N_5731);
or U5936 (N_5936,N_5556,N_5577);
nand U5937 (N_5937,N_5580,N_5519);
or U5938 (N_5938,N_5622,N_5563);
xnor U5939 (N_5939,N_5740,N_5646);
nand U5940 (N_5940,N_5610,N_5595);
nor U5941 (N_5941,N_5573,N_5568);
nand U5942 (N_5942,N_5565,N_5633);
xnor U5943 (N_5943,N_5694,N_5525);
nor U5944 (N_5944,N_5627,N_5663);
and U5945 (N_5945,N_5630,N_5545);
xor U5946 (N_5946,N_5662,N_5610);
xor U5947 (N_5947,N_5702,N_5565);
nor U5948 (N_5948,N_5641,N_5591);
and U5949 (N_5949,N_5517,N_5697);
nor U5950 (N_5950,N_5648,N_5696);
and U5951 (N_5951,N_5548,N_5704);
nor U5952 (N_5952,N_5743,N_5569);
nor U5953 (N_5953,N_5642,N_5530);
or U5954 (N_5954,N_5524,N_5584);
or U5955 (N_5955,N_5742,N_5584);
and U5956 (N_5956,N_5688,N_5698);
and U5957 (N_5957,N_5528,N_5728);
or U5958 (N_5958,N_5509,N_5504);
xnor U5959 (N_5959,N_5563,N_5611);
or U5960 (N_5960,N_5627,N_5571);
nor U5961 (N_5961,N_5556,N_5579);
nand U5962 (N_5962,N_5630,N_5672);
or U5963 (N_5963,N_5538,N_5545);
or U5964 (N_5964,N_5557,N_5680);
nand U5965 (N_5965,N_5575,N_5743);
nand U5966 (N_5966,N_5678,N_5746);
xnor U5967 (N_5967,N_5597,N_5727);
nor U5968 (N_5968,N_5614,N_5559);
or U5969 (N_5969,N_5626,N_5550);
and U5970 (N_5970,N_5535,N_5723);
nor U5971 (N_5971,N_5527,N_5592);
xnor U5972 (N_5972,N_5608,N_5511);
xnor U5973 (N_5973,N_5518,N_5540);
nand U5974 (N_5974,N_5683,N_5584);
nand U5975 (N_5975,N_5604,N_5521);
or U5976 (N_5976,N_5587,N_5504);
nor U5977 (N_5977,N_5679,N_5646);
or U5978 (N_5978,N_5555,N_5625);
or U5979 (N_5979,N_5719,N_5673);
or U5980 (N_5980,N_5640,N_5578);
xor U5981 (N_5981,N_5731,N_5614);
or U5982 (N_5982,N_5674,N_5733);
or U5983 (N_5983,N_5613,N_5685);
and U5984 (N_5984,N_5507,N_5702);
xor U5985 (N_5985,N_5676,N_5664);
or U5986 (N_5986,N_5544,N_5610);
nor U5987 (N_5987,N_5712,N_5610);
and U5988 (N_5988,N_5706,N_5733);
or U5989 (N_5989,N_5706,N_5599);
nand U5990 (N_5990,N_5653,N_5500);
or U5991 (N_5991,N_5728,N_5651);
nor U5992 (N_5992,N_5524,N_5550);
and U5993 (N_5993,N_5587,N_5618);
or U5994 (N_5994,N_5663,N_5654);
xor U5995 (N_5995,N_5691,N_5603);
nand U5996 (N_5996,N_5578,N_5634);
or U5997 (N_5997,N_5568,N_5626);
nand U5998 (N_5998,N_5608,N_5601);
nand U5999 (N_5999,N_5689,N_5707);
nor U6000 (N_6000,N_5840,N_5860);
or U6001 (N_6001,N_5930,N_5850);
and U6002 (N_6002,N_5969,N_5958);
nor U6003 (N_6003,N_5892,N_5907);
nor U6004 (N_6004,N_5831,N_5982);
nor U6005 (N_6005,N_5875,N_5906);
nand U6006 (N_6006,N_5932,N_5884);
nand U6007 (N_6007,N_5837,N_5825);
nor U6008 (N_6008,N_5876,N_5974);
nor U6009 (N_6009,N_5998,N_5754);
xor U6010 (N_6010,N_5920,N_5894);
and U6011 (N_6011,N_5960,N_5877);
or U6012 (N_6012,N_5781,N_5883);
nand U6013 (N_6013,N_5978,N_5964);
xnor U6014 (N_6014,N_5919,N_5834);
xor U6015 (N_6015,N_5935,N_5971);
nor U6016 (N_6016,N_5983,N_5793);
or U6017 (N_6017,N_5936,N_5939);
nor U6018 (N_6018,N_5921,N_5904);
xor U6019 (N_6019,N_5828,N_5829);
nand U6020 (N_6020,N_5853,N_5918);
xnor U6021 (N_6021,N_5788,N_5776);
nor U6022 (N_6022,N_5959,N_5782);
nand U6023 (N_6023,N_5847,N_5842);
and U6024 (N_6024,N_5815,N_5986);
nand U6025 (N_6025,N_5867,N_5896);
or U6026 (N_6026,N_5845,N_5813);
xnor U6027 (N_6027,N_5942,N_5812);
or U6028 (N_6028,N_5859,N_5796);
nand U6029 (N_6029,N_5862,N_5823);
and U6030 (N_6030,N_5784,N_5945);
and U6031 (N_6031,N_5885,N_5772);
or U6032 (N_6032,N_5928,N_5878);
xnor U6033 (N_6033,N_5756,N_5941);
nand U6034 (N_6034,N_5750,N_5809);
xnor U6035 (N_6035,N_5822,N_5949);
nand U6036 (N_6036,N_5900,N_5800);
nand U6037 (N_6037,N_5799,N_5947);
or U6038 (N_6038,N_5916,N_5880);
or U6039 (N_6039,N_5871,N_5984);
and U6040 (N_6040,N_5777,N_5890);
xor U6041 (N_6041,N_5761,N_5915);
nand U6042 (N_6042,N_5802,N_5855);
xnor U6043 (N_6043,N_5869,N_5752);
xor U6044 (N_6044,N_5786,N_5898);
and U6045 (N_6045,N_5897,N_5925);
and U6046 (N_6046,N_5922,N_5818);
and U6047 (N_6047,N_5775,N_5872);
or U6048 (N_6048,N_5993,N_5902);
and U6049 (N_6049,N_5961,N_5963);
nand U6050 (N_6050,N_5830,N_5950);
xor U6051 (N_6051,N_5765,N_5956);
nor U6052 (N_6052,N_5856,N_5968);
nor U6053 (N_6053,N_5911,N_5773);
or U6054 (N_6054,N_5913,N_5769);
xor U6055 (N_6055,N_5820,N_5865);
nand U6056 (N_6056,N_5927,N_5755);
nor U6057 (N_6057,N_5858,N_5758);
and U6058 (N_6058,N_5843,N_5926);
and U6059 (N_6059,N_5838,N_5912);
nand U6060 (N_6060,N_5962,N_5980);
nor U6061 (N_6061,N_5944,N_5899);
nor U6062 (N_6062,N_5821,N_5990);
and U6063 (N_6063,N_5953,N_5764);
nand U6064 (N_6064,N_5909,N_5891);
xnor U6065 (N_6065,N_5787,N_5934);
or U6066 (N_6066,N_5844,N_5763);
nand U6067 (N_6067,N_5979,N_5937);
and U6068 (N_6068,N_5790,N_5954);
or U6069 (N_6069,N_5996,N_5789);
nor U6070 (N_6070,N_5791,N_5767);
xnor U6071 (N_6071,N_5753,N_5943);
nand U6072 (N_6072,N_5832,N_5768);
xor U6073 (N_6073,N_5914,N_5957);
nand U6074 (N_6074,N_5987,N_5874);
and U6075 (N_6075,N_5895,N_5798);
and U6076 (N_6076,N_5864,N_5888);
nand U6077 (N_6077,N_5785,N_5766);
nand U6078 (N_6078,N_5866,N_5965);
and U6079 (N_6079,N_5863,N_5952);
or U6080 (N_6080,N_5994,N_5903);
nor U6081 (N_6081,N_5975,N_5846);
nand U6082 (N_6082,N_5991,N_5824);
nor U6083 (N_6083,N_5948,N_5835);
nor U6084 (N_6084,N_5999,N_5851);
and U6085 (N_6085,N_5807,N_5774);
xor U6086 (N_6086,N_5985,N_5827);
xor U6087 (N_6087,N_5879,N_5886);
xor U6088 (N_6088,N_5966,N_5908);
and U6089 (N_6089,N_5868,N_5839);
nand U6090 (N_6090,N_5910,N_5870);
nand U6091 (N_6091,N_5751,N_5970);
nand U6092 (N_6092,N_5816,N_5929);
nor U6093 (N_6093,N_5976,N_5792);
or U6094 (N_6094,N_5852,N_5826);
and U6095 (N_6095,N_5995,N_5757);
and U6096 (N_6096,N_5783,N_5811);
nor U6097 (N_6097,N_5794,N_5989);
xnor U6098 (N_6098,N_5992,N_5841);
nand U6099 (N_6099,N_5873,N_5977);
xnor U6100 (N_6100,N_5770,N_5946);
xnor U6101 (N_6101,N_5854,N_5905);
nand U6102 (N_6102,N_5988,N_5848);
nand U6103 (N_6103,N_5967,N_5972);
and U6104 (N_6104,N_5814,N_5887);
or U6105 (N_6105,N_5762,N_5810);
nand U6106 (N_6106,N_5951,N_5808);
nand U6107 (N_6107,N_5819,N_5940);
nor U6108 (N_6108,N_5923,N_5938);
nor U6109 (N_6109,N_5803,N_5759);
and U6110 (N_6110,N_5760,N_5805);
nand U6111 (N_6111,N_5933,N_5973);
or U6112 (N_6112,N_5833,N_5771);
and U6113 (N_6113,N_5857,N_5778);
nand U6114 (N_6114,N_5881,N_5931);
or U6115 (N_6115,N_5806,N_5901);
nor U6116 (N_6116,N_5836,N_5924);
xor U6117 (N_6117,N_5861,N_5817);
nor U6118 (N_6118,N_5797,N_5780);
nor U6119 (N_6119,N_5849,N_5981);
nor U6120 (N_6120,N_5804,N_5955);
nor U6121 (N_6121,N_5889,N_5917);
or U6122 (N_6122,N_5801,N_5997);
xor U6123 (N_6123,N_5882,N_5795);
or U6124 (N_6124,N_5779,N_5893);
or U6125 (N_6125,N_5908,N_5854);
or U6126 (N_6126,N_5947,N_5858);
or U6127 (N_6127,N_5916,N_5780);
nand U6128 (N_6128,N_5996,N_5892);
xnor U6129 (N_6129,N_5823,N_5817);
nand U6130 (N_6130,N_5789,N_5923);
nor U6131 (N_6131,N_5757,N_5784);
nor U6132 (N_6132,N_5933,N_5829);
xnor U6133 (N_6133,N_5805,N_5840);
xor U6134 (N_6134,N_5858,N_5821);
and U6135 (N_6135,N_5886,N_5883);
nand U6136 (N_6136,N_5936,N_5929);
and U6137 (N_6137,N_5964,N_5922);
nor U6138 (N_6138,N_5874,N_5822);
and U6139 (N_6139,N_5890,N_5789);
and U6140 (N_6140,N_5993,N_5943);
and U6141 (N_6141,N_5784,N_5859);
and U6142 (N_6142,N_5783,N_5933);
nand U6143 (N_6143,N_5822,N_5928);
and U6144 (N_6144,N_5828,N_5920);
or U6145 (N_6145,N_5971,N_5768);
and U6146 (N_6146,N_5796,N_5938);
nor U6147 (N_6147,N_5855,N_5838);
nor U6148 (N_6148,N_5763,N_5791);
nor U6149 (N_6149,N_5849,N_5763);
nand U6150 (N_6150,N_5881,N_5839);
and U6151 (N_6151,N_5894,N_5977);
nor U6152 (N_6152,N_5971,N_5829);
and U6153 (N_6153,N_5901,N_5979);
and U6154 (N_6154,N_5978,N_5755);
or U6155 (N_6155,N_5885,N_5994);
nor U6156 (N_6156,N_5900,N_5753);
nand U6157 (N_6157,N_5962,N_5883);
or U6158 (N_6158,N_5903,N_5917);
or U6159 (N_6159,N_5849,N_5824);
or U6160 (N_6160,N_5936,N_5942);
nand U6161 (N_6161,N_5997,N_5921);
nand U6162 (N_6162,N_5955,N_5814);
xnor U6163 (N_6163,N_5810,N_5989);
xor U6164 (N_6164,N_5997,N_5794);
or U6165 (N_6165,N_5827,N_5763);
xor U6166 (N_6166,N_5855,N_5840);
or U6167 (N_6167,N_5784,N_5817);
xor U6168 (N_6168,N_5932,N_5800);
or U6169 (N_6169,N_5986,N_5851);
and U6170 (N_6170,N_5940,N_5785);
nor U6171 (N_6171,N_5799,N_5930);
and U6172 (N_6172,N_5805,N_5905);
and U6173 (N_6173,N_5776,N_5827);
xor U6174 (N_6174,N_5792,N_5813);
nand U6175 (N_6175,N_5912,N_5915);
xnor U6176 (N_6176,N_5848,N_5775);
xnor U6177 (N_6177,N_5861,N_5907);
nand U6178 (N_6178,N_5919,N_5945);
and U6179 (N_6179,N_5797,N_5992);
or U6180 (N_6180,N_5919,N_5761);
and U6181 (N_6181,N_5788,N_5879);
nand U6182 (N_6182,N_5973,N_5961);
or U6183 (N_6183,N_5762,N_5837);
xor U6184 (N_6184,N_5885,N_5863);
or U6185 (N_6185,N_5957,N_5939);
or U6186 (N_6186,N_5878,N_5800);
and U6187 (N_6187,N_5999,N_5882);
and U6188 (N_6188,N_5964,N_5997);
xor U6189 (N_6189,N_5786,N_5879);
and U6190 (N_6190,N_5999,N_5824);
xnor U6191 (N_6191,N_5939,N_5887);
and U6192 (N_6192,N_5991,N_5990);
nand U6193 (N_6193,N_5780,N_5998);
nor U6194 (N_6194,N_5925,N_5860);
nand U6195 (N_6195,N_5922,N_5783);
and U6196 (N_6196,N_5803,N_5923);
or U6197 (N_6197,N_5754,N_5755);
nor U6198 (N_6198,N_5762,N_5858);
and U6199 (N_6199,N_5855,N_5763);
xor U6200 (N_6200,N_5839,N_5751);
xnor U6201 (N_6201,N_5806,N_5771);
nand U6202 (N_6202,N_5839,N_5890);
nand U6203 (N_6203,N_5813,N_5812);
or U6204 (N_6204,N_5929,N_5872);
nor U6205 (N_6205,N_5755,N_5923);
and U6206 (N_6206,N_5900,N_5891);
nor U6207 (N_6207,N_5979,N_5944);
nand U6208 (N_6208,N_5908,N_5921);
nor U6209 (N_6209,N_5751,N_5919);
or U6210 (N_6210,N_5843,N_5917);
nor U6211 (N_6211,N_5805,N_5839);
or U6212 (N_6212,N_5884,N_5757);
nor U6213 (N_6213,N_5957,N_5813);
or U6214 (N_6214,N_5954,N_5809);
nor U6215 (N_6215,N_5979,N_5840);
nand U6216 (N_6216,N_5959,N_5983);
and U6217 (N_6217,N_5779,N_5972);
and U6218 (N_6218,N_5983,N_5809);
and U6219 (N_6219,N_5887,N_5989);
nor U6220 (N_6220,N_5978,N_5876);
nand U6221 (N_6221,N_5897,N_5903);
nor U6222 (N_6222,N_5981,N_5953);
or U6223 (N_6223,N_5842,N_5854);
nor U6224 (N_6224,N_5783,N_5789);
or U6225 (N_6225,N_5892,N_5816);
or U6226 (N_6226,N_5879,N_5939);
xor U6227 (N_6227,N_5839,N_5970);
and U6228 (N_6228,N_5934,N_5799);
nand U6229 (N_6229,N_5889,N_5760);
and U6230 (N_6230,N_5812,N_5932);
xor U6231 (N_6231,N_5880,N_5869);
or U6232 (N_6232,N_5817,N_5812);
xor U6233 (N_6233,N_5895,N_5890);
nor U6234 (N_6234,N_5911,N_5937);
and U6235 (N_6235,N_5875,N_5810);
nand U6236 (N_6236,N_5756,N_5840);
xor U6237 (N_6237,N_5820,N_5933);
xnor U6238 (N_6238,N_5765,N_5927);
and U6239 (N_6239,N_5960,N_5939);
nand U6240 (N_6240,N_5971,N_5920);
nand U6241 (N_6241,N_5798,N_5899);
xnor U6242 (N_6242,N_5812,N_5866);
nor U6243 (N_6243,N_5934,N_5768);
or U6244 (N_6244,N_5922,N_5751);
and U6245 (N_6245,N_5766,N_5978);
and U6246 (N_6246,N_5772,N_5757);
nor U6247 (N_6247,N_5973,N_5778);
xnor U6248 (N_6248,N_5954,N_5755);
and U6249 (N_6249,N_5956,N_5889);
nor U6250 (N_6250,N_6078,N_6186);
nand U6251 (N_6251,N_6201,N_6162);
nand U6252 (N_6252,N_6089,N_6134);
xor U6253 (N_6253,N_6053,N_6199);
and U6254 (N_6254,N_6137,N_6002);
nand U6255 (N_6255,N_6084,N_6048);
xnor U6256 (N_6256,N_6118,N_6046);
or U6257 (N_6257,N_6129,N_6147);
xor U6258 (N_6258,N_6082,N_6063);
xor U6259 (N_6259,N_6206,N_6044);
and U6260 (N_6260,N_6218,N_6023);
or U6261 (N_6261,N_6025,N_6145);
nor U6262 (N_6262,N_6178,N_6144);
nand U6263 (N_6263,N_6071,N_6010);
and U6264 (N_6264,N_6229,N_6116);
or U6265 (N_6265,N_6168,N_6087);
nor U6266 (N_6266,N_6222,N_6183);
or U6267 (N_6267,N_6181,N_6212);
xnor U6268 (N_6268,N_6072,N_6188);
nor U6269 (N_6269,N_6249,N_6031);
xor U6270 (N_6270,N_6146,N_6080);
or U6271 (N_6271,N_6018,N_6111);
xnor U6272 (N_6272,N_6032,N_6180);
and U6273 (N_6273,N_6141,N_6210);
or U6274 (N_6274,N_6047,N_6112);
xnor U6275 (N_6275,N_6193,N_6248);
nand U6276 (N_6276,N_6170,N_6035);
xnor U6277 (N_6277,N_6211,N_6194);
nand U6278 (N_6278,N_6050,N_6090);
and U6279 (N_6279,N_6039,N_6081);
nor U6280 (N_6280,N_6221,N_6200);
and U6281 (N_6281,N_6003,N_6088);
or U6282 (N_6282,N_6175,N_6238);
xnor U6283 (N_6283,N_6156,N_6057);
xor U6284 (N_6284,N_6167,N_6026);
nor U6285 (N_6285,N_6166,N_6065);
nor U6286 (N_6286,N_6066,N_6120);
nand U6287 (N_6287,N_6091,N_6110);
nand U6288 (N_6288,N_6242,N_6030);
nor U6289 (N_6289,N_6171,N_6086);
nor U6290 (N_6290,N_6119,N_6027);
nor U6291 (N_6291,N_6226,N_6219);
nor U6292 (N_6292,N_6244,N_6055);
nor U6293 (N_6293,N_6061,N_6203);
or U6294 (N_6294,N_6138,N_6028);
nand U6295 (N_6295,N_6142,N_6017);
and U6296 (N_6296,N_6069,N_6224);
nor U6297 (N_6297,N_6000,N_6052);
or U6298 (N_6298,N_6140,N_6108);
or U6299 (N_6299,N_6106,N_6241);
and U6300 (N_6300,N_6208,N_6235);
xnor U6301 (N_6301,N_6216,N_6196);
nand U6302 (N_6302,N_6185,N_6041);
nand U6303 (N_6303,N_6165,N_6058);
nand U6304 (N_6304,N_6126,N_6105);
xnor U6305 (N_6305,N_6164,N_6060);
xnor U6306 (N_6306,N_6098,N_6040);
and U6307 (N_6307,N_6240,N_6195);
or U6308 (N_6308,N_6005,N_6093);
xnor U6309 (N_6309,N_6103,N_6109);
xnor U6310 (N_6310,N_6107,N_6095);
nor U6311 (N_6311,N_6092,N_6190);
xor U6312 (N_6312,N_6022,N_6101);
or U6313 (N_6313,N_6076,N_6079);
xnor U6314 (N_6314,N_6013,N_6139);
nand U6315 (N_6315,N_6136,N_6014);
or U6316 (N_6316,N_6127,N_6148);
xor U6317 (N_6317,N_6074,N_6202);
xnor U6318 (N_6318,N_6214,N_6243);
nor U6319 (N_6319,N_6132,N_6024);
nor U6320 (N_6320,N_6124,N_6070);
xnor U6321 (N_6321,N_6045,N_6231);
xor U6322 (N_6322,N_6020,N_6153);
nor U6323 (N_6323,N_6100,N_6239);
nand U6324 (N_6324,N_6004,N_6197);
or U6325 (N_6325,N_6036,N_6054);
nor U6326 (N_6326,N_6143,N_6209);
and U6327 (N_6327,N_6161,N_6245);
and U6328 (N_6328,N_6099,N_6122);
nand U6329 (N_6329,N_6051,N_6007);
and U6330 (N_6330,N_6182,N_6152);
nand U6331 (N_6331,N_6217,N_6228);
xnor U6332 (N_6332,N_6021,N_6192);
nor U6333 (N_6333,N_6177,N_6247);
and U6334 (N_6334,N_6113,N_6029);
nand U6335 (N_6335,N_6172,N_6033);
xor U6336 (N_6336,N_6135,N_6037);
nor U6337 (N_6337,N_6094,N_6097);
nor U6338 (N_6338,N_6001,N_6008);
nor U6339 (N_6339,N_6012,N_6160);
and U6340 (N_6340,N_6233,N_6174);
xnor U6341 (N_6341,N_6184,N_6102);
or U6342 (N_6342,N_6130,N_6151);
nor U6343 (N_6343,N_6230,N_6232);
and U6344 (N_6344,N_6176,N_6154);
and U6345 (N_6345,N_6034,N_6173);
and U6346 (N_6346,N_6067,N_6011);
and U6347 (N_6347,N_6237,N_6049);
and U6348 (N_6348,N_6159,N_6223);
or U6349 (N_6349,N_6042,N_6015);
and U6350 (N_6350,N_6009,N_6149);
nand U6351 (N_6351,N_6179,N_6234);
or U6352 (N_6352,N_6104,N_6207);
and U6353 (N_6353,N_6043,N_6169);
xnor U6354 (N_6354,N_6075,N_6220);
nand U6355 (N_6355,N_6019,N_6096);
nand U6356 (N_6356,N_6150,N_6117);
nand U6357 (N_6357,N_6155,N_6163);
nor U6358 (N_6358,N_6062,N_6157);
or U6359 (N_6359,N_6125,N_6204);
nor U6360 (N_6360,N_6213,N_6225);
xor U6361 (N_6361,N_6123,N_6198);
xor U6362 (N_6362,N_6205,N_6115);
and U6363 (N_6363,N_6059,N_6128);
nor U6364 (N_6364,N_6187,N_6085);
xor U6365 (N_6365,N_6077,N_6227);
nor U6366 (N_6366,N_6121,N_6133);
xor U6367 (N_6367,N_6191,N_6246);
nor U6368 (N_6368,N_6189,N_6073);
nand U6369 (N_6369,N_6038,N_6215);
xnor U6370 (N_6370,N_6064,N_6131);
xor U6371 (N_6371,N_6016,N_6236);
xor U6372 (N_6372,N_6083,N_6068);
and U6373 (N_6373,N_6006,N_6158);
nor U6374 (N_6374,N_6056,N_6114);
or U6375 (N_6375,N_6070,N_6187);
nor U6376 (N_6376,N_6062,N_6041);
or U6377 (N_6377,N_6246,N_6244);
nor U6378 (N_6378,N_6131,N_6241);
nor U6379 (N_6379,N_6057,N_6026);
or U6380 (N_6380,N_6017,N_6028);
nand U6381 (N_6381,N_6160,N_6107);
and U6382 (N_6382,N_6001,N_6245);
nand U6383 (N_6383,N_6118,N_6134);
nor U6384 (N_6384,N_6227,N_6146);
xor U6385 (N_6385,N_6211,N_6201);
nor U6386 (N_6386,N_6019,N_6093);
nand U6387 (N_6387,N_6248,N_6243);
and U6388 (N_6388,N_6123,N_6240);
xnor U6389 (N_6389,N_6109,N_6213);
xor U6390 (N_6390,N_6243,N_6028);
and U6391 (N_6391,N_6054,N_6127);
and U6392 (N_6392,N_6227,N_6095);
xnor U6393 (N_6393,N_6189,N_6152);
and U6394 (N_6394,N_6022,N_6150);
xnor U6395 (N_6395,N_6206,N_6195);
nor U6396 (N_6396,N_6076,N_6144);
and U6397 (N_6397,N_6024,N_6144);
nand U6398 (N_6398,N_6225,N_6239);
xnor U6399 (N_6399,N_6233,N_6243);
or U6400 (N_6400,N_6155,N_6092);
and U6401 (N_6401,N_6105,N_6002);
xor U6402 (N_6402,N_6137,N_6088);
nor U6403 (N_6403,N_6072,N_6030);
nor U6404 (N_6404,N_6180,N_6230);
nor U6405 (N_6405,N_6195,N_6112);
or U6406 (N_6406,N_6239,N_6180);
or U6407 (N_6407,N_6238,N_6094);
xor U6408 (N_6408,N_6217,N_6002);
nor U6409 (N_6409,N_6098,N_6146);
nand U6410 (N_6410,N_6119,N_6237);
nand U6411 (N_6411,N_6143,N_6021);
nand U6412 (N_6412,N_6029,N_6238);
nor U6413 (N_6413,N_6173,N_6184);
nand U6414 (N_6414,N_6223,N_6001);
xnor U6415 (N_6415,N_6025,N_6101);
or U6416 (N_6416,N_6067,N_6161);
or U6417 (N_6417,N_6027,N_6034);
nand U6418 (N_6418,N_6062,N_6039);
or U6419 (N_6419,N_6213,N_6229);
or U6420 (N_6420,N_6047,N_6094);
xnor U6421 (N_6421,N_6175,N_6013);
nand U6422 (N_6422,N_6145,N_6170);
xnor U6423 (N_6423,N_6077,N_6160);
nor U6424 (N_6424,N_6152,N_6007);
and U6425 (N_6425,N_6164,N_6032);
xor U6426 (N_6426,N_6109,N_6106);
and U6427 (N_6427,N_6071,N_6009);
nand U6428 (N_6428,N_6115,N_6040);
and U6429 (N_6429,N_6061,N_6051);
nand U6430 (N_6430,N_6085,N_6000);
nor U6431 (N_6431,N_6032,N_6186);
nand U6432 (N_6432,N_6078,N_6084);
xor U6433 (N_6433,N_6092,N_6182);
and U6434 (N_6434,N_6221,N_6053);
nand U6435 (N_6435,N_6080,N_6055);
xor U6436 (N_6436,N_6007,N_6232);
xnor U6437 (N_6437,N_6003,N_6112);
xor U6438 (N_6438,N_6104,N_6042);
xnor U6439 (N_6439,N_6196,N_6139);
or U6440 (N_6440,N_6154,N_6101);
xor U6441 (N_6441,N_6019,N_6129);
nand U6442 (N_6442,N_6047,N_6149);
xor U6443 (N_6443,N_6129,N_6073);
nand U6444 (N_6444,N_6152,N_6143);
nand U6445 (N_6445,N_6222,N_6153);
and U6446 (N_6446,N_6011,N_6014);
xnor U6447 (N_6447,N_6055,N_6246);
or U6448 (N_6448,N_6107,N_6106);
or U6449 (N_6449,N_6241,N_6047);
xor U6450 (N_6450,N_6101,N_6246);
nand U6451 (N_6451,N_6168,N_6170);
xnor U6452 (N_6452,N_6117,N_6111);
nand U6453 (N_6453,N_6133,N_6053);
or U6454 (N_6454,N_6096,N_6022);
nor U6455 (N_6455,N_6161,N_6225);
nand U6456 (N_6456,N_6053,N_6183);
or U6457 (N_6457,N_6227,N_6012);
and U6458 (N_6458,N_6232,N_6212);
xnor U6459 (N_6459,N_6079,N_6046);
nand U6460 (N_6460,N_6119,N_6006);
nor U6461 (N_6461,N_6089,N_6073);
and U6462 (N_6462,N_6091,N_6098);
nand U6463 (N_6463,N_6095,N_6221);
or U6464 (N_6464,N_6193,N_6042);
nor U6465 (N_6465,N_6188,N_6090);
and U6466 (N_6466,N_6039,N_6202);
xor U6467 (N_6467,N_6236,N_6154);
nand U6468 (N_6468,N_6205,N_6055);
and U6469 (N_6469,N_6078,N_6043);
and U6470 (N_6470,N_6055,N_6166);
or U6471 (N_6471,N_6103,N_6130);
xnor U6472 (N_6472,N_6060,N_6094);
and U6473 (N_6473,N_6009,N_6010);
nand U6474 (N_6474,N_6137,N_6111);
or U6475 (N_6475,N_6014,N_6156);
nand U6476 (N_6476,N_6170,N_6116);
nand U6477 (N_6477,N_6046,N_6159);
nor U6478 (N_6478,N_6035,N_6079);
or U6479 (N_6479,N_6213,N_6145);
nor U6480 (N_6480,N_6185,N_6223);
xor U6481 (N_6481,N_6008,N_6157);
nand U6482 (N_6482,N_6028,N_6211);
or U6483 (N_6483,N_6083,N_6156);
nand U6484 (N_6484,N_6154,N_6054);
nand U6485 (N_6485,N_6159,N_6208);
xor U6486 (N_6486,N_6039,N_6231);
or U6487 (N_6487,N_6064,N_6194);
or U6488 (N_6488,N_6207,N_6019);
or U6489 (N_6489,N_6104,N_6229);
and U6490 (N_6490,N_6077,N_6144);
or U6491 (N_6491,N_6212,N_6213);
and U6492 (N_6492,N_6026,N_6147);
xnor U6493 (N_6493,N_6127,N_6069);
and U6494 (N_6494,N_6229,N_6137);
or U6495 (N_6495,N_6164,N_6180);
nand U6496 (N_6496,N_6124,N_6148);
or U6497 (N_6497,N_6212,N_6033);
nand U6498 (N_6498,N_6115,N_6185);
and U6499 (N_6499,N_6210,N_6112);
or U6500 (N_6500,N_6347,N_6300);
xnor U6501 (N_6501,N_6397,N_6334);
xor U6502 (N_6502,N_6403,N_6484);
nand U6503 (N_6503,N_6423,N_6294);
nor U6504 (N_6504,N_6273,N_6393);
nor U6505 (N_6505,N_6369,N_6394);
and U6506 (N_6506,N_6436,N_6284);
nand U6507 (N_6507,N_6455,N_6461);
or U6508 (N_6508,N_6442,N_6489);
xnor U6509 (N_6509,N_6315,N_6496);
nand U6510 (N_6510,N_6482,N_6278);
nor U6511 (N_6511,N_6493,N_6331);
xnor U6512 (N_6512,N_6299,N_6332);
or U6513 (N_6513,N_6372,N_6324);
nor U6514 (N_6514,N_6430,N_6473);
nor U6515 (N_6515,N_6255,N_6470);
or U6516 (N_6516,N_6379,N_6296);
nor U6517 (N_6517,N_6361,N_6456);
or U6518 (N_6518,N_6398,N_6306);
and U6519 (N_6519,N_6475,N_6349);
nor U6520 (N_6520,N_6320,N_6257);
nand U6521 (N_6521,N_6440,N_6425);
and U6522 (N_6522,N_6271,N_6419);
xnor U6523 (N_6523,N_6437,N_6252);
xor U6524 (N_6524,N_6406,N_6408);
nand U6525 (N_6525,N_6333,N_6363);
nor U6526 (N_6526,N_6365,N_6370);
nor U6527 (N_6527,N_6476,N_6384);
or U6528 (N_6528,N_6356,N_6424);
nor U6529 (N_6529,N_6301,N_6351);
nor U6530 (N_6530,N_6367,N_6358);
xnor U6531 (N_6531,N_6302,N_6413);
and U6532 (N_6532,N_6359,N_6345);
nand U6533 (N_6533,N_6480,N_6499);
nor U6534 (N_6534,N_6486,N_6348);
nand U6535 (N_6535,N_6339,N_6405);
or U6536 (N_6536,N_6410,N_6421);
nand U6537 (N_6537,N_6277,N_6495);
xor U6538 (N_6538,N_6488,N_6481);
xnor U6539 (N_6539,N_6326,N_6313);
nor U6540 (N_6540,N_6281,N_6264);
nand U6541 (N_6541,N_6450,N_6487);
or U6542 (N_6542,N_6328,N_6344);
and U6543 (N_6543,N_6290,N_6311);
or U6544 (N_6544,N_6428,N_6454);
and U6545 (N_6545,N_6375,N_6256);
or U6546 (N_6546,N_6498,N_6389);
nand U6547 (N_6547,N_6402,N_6350);
xnor U6548 (N_6548,N_6411,N_6357);
nand U6549 (N_6549,N_6462,N_6441);
xor U6550 (N_6550,N_6308,N_6265);
and U6551 (N_6551,N_6280,N_6269);
and U6552 (N_6552,N_6383,N_6274);
and U6553 (N_6553,N_6292,N_6459);
nand U6554 (N_6554,N_6352,N_6293);
nand U6555 (N_6555,N_6390,N_6409);
nand U6556 (N_6556,N_6317,N_6483);
and U6557 (N_6557,N_6453,N_6445);
xor U6558 (N_6558,N_6387,N_6270);
nand U6559 (N_6559,N_6282,N_6309);
and U6560 (N_6560,N_6467,N_6378);
nand U6561 (N_6561,N_6435,N_6472);
and U6562 (N_6562,N_6360,N_6283);
nor U6563 (N_6563,N_6429,N_6434);
or U6564 (N_6564,N_6422,N_6287);
nor U6565 (N_6565,N_6376,N_6298);
nor U6566 (N_6566,N_6346,N_6400);
xnor U6567 (N_6567,N_6342,N_6263);
and U6568 (N_6568,N_6285,N_6416);
or U6569 (N_6569,N_6374,N_6254);
xor U6570 (N_6570,N_6318,N_6266);
and U6571 (N_6571,N_6272,N_6340);
or U6572 (N_6572,N_6446,N_6439);
nor U6573 (N_6573,N_6380,N_6362);
or U6574 (N_6574,N_6343,N_6316);
or U6575 (N_6575,N_6432,N_6388);
xor U6576 (N_6576,N_6305,N_6490);
nand U6577 (N_6577,N_6321,N_6417);
or U6578 (N_6578,N_6426,N_6291);
nand U6579 (N_6579,N_6492,N_6449);
or U6580 (N_6580,N_6353,N_6335);
or U6581 (N_6581,N_6338,N_6377);
nand U6582 (N_6582,N_6391,N_6327);
nand U6583 (N_6583,N_6295,N_6494);
or U6584 (N_6584,N_6443,N_6268);
nand U6585 (N_6585,N_6312,N_6262);
and U6586 (N_6586,N_6477,N_6341);
or U6587 (N_6587,N_6431,N_6414);
and U6588 (N_6588,N_6330,N_6322);
xor U6589 (N_6589,N_6364,N_6447);
nand U6590 (N_6590,N_6415,N_6448);
xnor U6591 (N_6591,N_6497,N_6386);
nand U6592 (N_6592,N_6258,N_6276);
and U6593 (N_6593,N_6354,N_6304);
and U6594 (N_6594,N_6392,N_6469);
xnor U6595 (N_6595,N_6418,N_6297);
xor U6596 (N_6596,N_6468,N_6382);
or U6597 (N_6597,N_6381,N_6323);
xnor U6598 (N_6598,N_6463,N_6325);
nor U6599 (N_6599,N_6310,N_6267);
or U6600 (N_6600,N_6458,N_6261);
xor U6601 (N_6601,N_6474,N_6478);
nor U6602 (N_6602,N_6319,N_6433);
or U6603 (N_6603,N_6286,N_6465);
xor U6604 (N_6604,N_6289,N_6407);
nand U6605 (N_6605,N_6464,N_6399);
and U6606 (N_6606,N_6420,N_6337);
xnor U6607 (N_6607,N_6401,N_6412);
nand U6608 (N_6608,N_6471,N_6460);
nor U6609 (N_6609,N_6307,N_6452);
nor U6610 (N_6610,N_6385,N_6438);
and U6611 (N_6611,N_6396,N_6371);
nand U6612 (N_6612,N_6260,N_6485);
nand U6613 (N_6613,N_6279,N_6368);
xor U6614 (N_6614,N_6251,N_6427);
or U6615 (N_6615,N_6275,N_6303);
or U6616 (N_6616,N_6444,N_6479);
nor U6617 (N_6617,N_6253,N_6457);
and U6618 (N_6618,N_6314,N_6451);
nand U6619 (N_6619,N_6336,N_6404);
nor U6620 (N_6620,N_6366,N_6466);
and U6621 (N_6621,N_6355,N_6491);
nand U6622 (N_6622,N_6259,N_6329);
and U6623 (N_6623,N_6250,N_6395);
xnor U6624 (N_6624,N_6373,N_6288);
xnor U6625 (N_6625,N_6390,N_6335);
xor U6626 (N_6626,N_6407,N_6477);
xnor U6627 (N_6627,N_6253,N_6451);
and U6628 (N_6628,N_6359,N_6485);
nand U6629 (N_6629,N_6278,N_6333);
nand U6630 (N_6630,N_6475,N_6430);
nand U6631 (N_6631,N_6475,N_6477);
or U6632 (N_6632,N_6332,N_6359);
and U6633 (N_6633,N_6342,N_6478);
or U6634 (N_6634,N_6492,N_6491);
and U6635 (N_6635,N_6271,N_6350);
nor U6636 (N_6636,N_6255,N_6455);
nand U6637 (N_6637,N_6391,N_6484);
nor U6638 (N_6638,N_6486,N_6421);
and U6639 (N_6639,N_6400,N_6318);
nor U6640 (N_6640,N_6259,N_6401);
xor U6641 (N_6641,N_6432,N_6431);
nor U6642 (N_6642,N_6253,N_6321);
nand U6643 (N_6643,N_6387,N_6310);
xor U6644 (N_6644,N_6429,N_6288);
and U6645 (N_6645,N_6471,N_6331);
nand U6646 (N_6646,N_6258,N_6490);
nor U6647 (N_6647,N_6282,N_6342);
xnor U6648 (N_6648,N_6368,N_6345);
or U6649 (N_6649,N_6286,N_6456);
and U6650 (N_6650,N_6339,N_6375);
nand U6651 (N_6651,N_6453,N_6283);
xnor U6652 (N_6652,N_6461,N_6310);
and U6653 (N_6653,N_6393,N_6268);
or U6654 (N_6654,N_6452,N_6454);
or U6655 (N_6655,N_6398,N_6335);
and U6656 (N_6656,N_6272,N_6441);
xor U6657 (N_6657,N_6491,N_6485);
xor U6658 (N_6658,N_6338,N_6373);
and U6659 (N_6659,N_6414,N_6363);
or U6660 (N_6660,N_6373,N_6313);
and U6661 (N_6661,N_6386,N_6252);
nand U6662 (N_6662,N_6414,N_6281);
nor U6663 (N_6663,N_6415,N_6491);
or U6664 (N_6664,N_6276,N_6310);
xor U6665 (N_6665,N_6298,N_6345);
nor U6666 (N_6666,N_6286,N_6414);
xnor U6667 (N_6667,N_6395,N_6489);
and U6668 (N_6668,N_6285,N_6292);
or U6669 (N_6669,N_6368,N_6260);
or U6670 (N_6670,N_6377,N_6303);
and U6671 (N_6671,N_6481,N_6450);
xnor U6672 (N_6672,N_6407,N_6264);
and U6673 (N_6673,N_6481,N_6308);
nor U6674 (N_6674,N_6484,N_6378);
xnor U6675 (N_6675,N_6442,N_6357);
nand U6676 (N_6676,N_6435,N_6370);
and U6677 (N_6677,N_6300,N_6288);
or U6678 (N_6678,N_6338,N_6281);
or U6679 (N_6679,N_6456,N_6315);
nor U6680 (N_6680,N_6303,N_6338);
or U6681 (N_6681,N_6276,N_6480);
nand U6682 (N_6682,N_6456,N_6281);
nor U6683 (N_6683,N_6286,N_6390);
xnor U6684 (N_6684,N_6282,N_6395);
xor U6685 (N_6685,N_6479,N_6476);
and U6686 (N_6686,N_6435,N_6480);
or U6687 (N_6687,N_6286,N_6346);
nor U6688 (N_6688,N_6297,N_6303);
nor U6689 (N_6689,N_6478,N_6338);
nand U6690 (N_6690,N_6288,N_6420);
and U6691 (N_6691,N_6354,N_6326);
nand U6692 (N_6692,N_6316,N_6290);
xnor U6693 (N_6693,N_6356,N_6252);
nor U6694 (N_6694,N_6407,N_6271);
nor U6695 (N_6695,N_6406,N_6299);
nor U6696 (N_6696,N_6376,N_6325);
nor U6697 (N_6697,N_6416,N_6311);
nand U6698 (N_6698,N_6320,N_6376);
and U6699 (N_6699,N_6367,N_6333);
xnor U6700 (N_6700,N_6426,N_6359);
and U6701 (N_6701,N_6311,N_6280);
nand U6702 (N_6702,N_6463,N_6283);
xor U6703 (N_6703,N_6372,N_6328);
nor U6704 (N_6704,N_6412,N_6457);
xnor U6705 (N_6705,N_6485,N_6469);
nand U6706 (N_6706,N_6421,N_6422);
nor U6707 (N_6707,N_6415,N_6366);
or U6708 (N_6708,N_6341,N_6442);
nor U6709 (N_6709,N_6396,N_6264);
and U6710 (N_6710,N_6499,N_6391);
nor U6711 (N_6711,N_6269,N_6427);
or U6712 (N_6712,N_6327,N_6477);
xor U6713 (N_6713,N_6339,N_6432);
or U6714 (N_6714,N_6420,N_6410);
xnor U6715 (N_6715,N_6356,N_6402);
and U6716 (N_6716,N_6475,N_6393);
nand U6717 (N_6717,N_6491,N_6388);
or U6718 (N_6718,N_6402,N_6366);
or U6719 (N_6719,N_6285,N_6355);
or U6720 (N_6720,N_6375,N_6417);
or U6721 (N_6721,N_6439,N_6261);
nand U6722 (N_6722,N_6412,N_6489);
or U6723 (N_6723,N_6438,N_6253);
nand U6724 (N_6724,N_6472,N_6468);
xor U6725 (N_6725,N_6450,N_6470);
and U6726 (N_6726,N_6475,N_6427);
and U6727 (N_6727,N_6404,N_6285);
nor U6728 (N_6728,N_6422,N_6260);
nor U6729 (N_6729,N_6417,N_6312);
or U6730 (N_6730,N_6493,N_6314);
and U6731 (N_6731,N_6268,N_6437);
or U6732 (N_6732,N_6324,N_6423);
xnor U6733 (N_6733,N_6364,N_6482);
and U6734 (N_6734,N_6317,N_6407);
nand U6735 (N_6735,N_6265,N_6310);
or U6736 (N_6736,N_6278,N_6433);
xor U6737 (N_6737,N_6262,N_6476);
nand U6738 (N_6738,N_6460,N_6412);
nand U6739 (N_6739,N_6319,N_6449);
nand U6740 (N_6740,N_6499,N_6433);
xnor U6741 (N_6741,N_6492,N_6353);
nor U6742 (N_6742,N_6338,N_6351);
or U6743 (N_6743,N_6304,N_6258);
nor U6744 (N_6744,N_6352,N_6467);
or U6745 (N_6745,N_6347,N_6402);
nand U6746 (N_6746,N_6322,N_6376);
or U6747 (N_6747,N_6469,N_6342);
nand U6748 (N_6748,N_6304,N_6375);
xor U6749 (N_6749,N_6324,N_6430);
nor U6750 (N_6750,N_6668,N_6637);
xor U6751 (N_6751,N_6734,N_6695);
and U6752 (N_6752,N_6581,N_6701);
xnor U6753 (N_6753,N_6573,N_6727);
and U6754 (N_6754,N_6541,N_6661);
and U6755 (N_6755,N_6642,N_6656);
xnor U6756 (N_6756,N_6691,N_6548);
and U6757 (N_6757,N_6572,N_6558);
nand U6758 (N_6758,N_6585,N_6561);
and U6759 (N_6759,N_6684,N_6509);
nand U6760 (N_6760,N_6510,N_6749);
nor U6761 (N_6761,N_6711,N_6718);
nor U6762 (N_6762,N_6594,N_6741);
xnor U6763 (N_6763,N_6714,N_6624);
xor U6764 (N_6764,N_6725,N_6644);
nor U6765 (N_6765,N_6640,N_6608);
xnor U6766 (N_6766,N_6702,N_6559);
nand U6767 (N_6767,N_6738,N_6721);
nand U6768 (N_6768,N_6516,N_6690);
and U6769 (N_6769,N_6681,N_6550);
xor U6770 (N_6770,N_6505,N_6658);
nor U6771 (N_6771,N_6523,N_6625);
nor U6772 (N_6772,N_6551,N_6615);
or U6773 (N_6773,N_6515,N_6700);
and U6774 (N_6774,N_6655,N_6612);
xnor U6775 (N_6775,N_6571,N_6586);
xor U6776 (N_6776,N_6611,N_6533);
and U6777 (N_6777,N_6748,N_6710);
nand U6778 (N_6778,N_6588,N_6547);
and U6779 (N_6779,N_6743,N_6745);
or U6780 (N_6780,N_6631,N_6512);
xnor U6781 (N_6781,N_6507,N_6518);
and U6782 (N_6782,N_6660,N_6713);
nor U6783 (N_6783,N_6531,N_6706);
or U6784 (N_6784,N_6705,N_6662);
and U6785 (N_6785,N_6514,N_6526);
or U6786 (N_6786,N_6542,N_6519);
and U6787 (N_6787,N_6715,N_6698);
or U6788 (N_6788,N_6556,N_6545);
or U6789 (N_6789,N_6520,N_6630);
nand U6790 (N_6790,N_6636,N_6595);
and U6791 (N_6791,N_6641,N_6628);
or U6792 (N_6792,N_6600,N_6688);
nand U6793 (N_6793,N_6722,N_6593);
or U6794 (N_6794,N_6685,N_6704);
nor U6795 (N_6795,N_6543,N_6536);
and U6796 (N_6796,N_6579,N_6553);
nor U6797 (N_6797,N_6513,N_6597);
nor U6798 (N_6798,N_6583,N_6564);
or U6799 (N_6799,N_6739,N_6665);
and U6800 (N_6800,N_6546,N_6663);
xor U6801 (N_6801,N_6511,N_6694);
nor U6802 (N_6802,N_6707,N_6563);
or U6803 (N_6803,N_6598,N_6649);
or U6804 (N_6804,N_6610,N_6517);
and U6805 (N_6805,N_6742,N_6746);
xor U6806 (N_6806,N_6549,N_6692);
xnor U6807 (N_6807,N_6678,N_6537);
or U6808 (N_6808,N_6500,N_6724);
xor U6809 (N_6809,N_6577,N_6570);
xnor U6810 (N_6810,N_6635,N_6659);
or U6811 (N_6811,N_6618,N_6651);
nand U6812 (N_6812,N_6667,N_6666);
and U6813 (N_6813,N_6673,N_6530);
xor U6814 (N_6814,N_6647,N_6565);
or U6815 (N_6815,N_6669,N_6538);
and U6816 (N_6816,N_6645,N_6699);
or U6817 (N_6817,N_6508,N_6524);
and U6818 (N_6818,N_6639,N_6535);
nand U6819 (N_6819,N_6560,N_6616);
nor U6820 (N_6820,N_6569,N_6687);
xor U6821 (N_6821,N_6672,N_6590);
xor U6822 (N_6822,N_6719,N_6697);
nand U6823 (N_6823,N_6621,N_6653);
nand U6824 (N_6824,N_6646,N_6629);
and U6825 (N_6825,N_6601,N_6592);
xnor U6826 (N_6826,N_6716,N_6620);
xnor U6827 (N_6827,N_6606,N_6522);
or U6828 (N_6828,N_6696,N_6723);
nand U6829 (N_6829,N_6613,N_6528);
or U6830 (N_6830,N_6557,N_6679);
nor U6831 (N_6831,N_6609,N_6619);
or U6832 (N_6832,N_6554,N_6638);
or U6833 (N_6833,N_6689,N_6584);
nand U6834 (N_6834,N_6632,N_6532);
and U6835 (N_6835,N_6596,N_6575);
and U6836 (N_6836,N_6568,N_6539);
and U6837 (N_6837,N_6604,N_6622);
and U6838 (N_6838,N_6540,N_6708);
xnor U6839 (N_6839,N_6657,N_6671);
and U6840 (N_6840,N_6730,N_6502);
nand U6841 (N_6841,N_6720,N_6728);
xnor U6842 (N_6842,N_6617,N_6626);
nand U6843 (N_6843,N_6562,N_6567);
xnor U6844 (N_6844,N_6693,N_6576);
xnor U6845 (N_6845,N_6623,N_6627);
nand U6846 (N_6846,N_6503,N_6555);
nand U6847 (N_6847,N_6633,N_6574);
xor U6848 (N_6848,N_6740,N_6582);
xor U6849 (N_6849,N_6650,N_6527);
xnor U6850 (N_6850,N_6566,N_6534);
nor U6851 (N_6851,N_6732,N_6735);
nor U6852 (N_6852,N_6709,N_6731);
xnor U6853 (N_6853,N_6726,N_6525);
and U6854 (N_6854,N_6682,N_6552);
xnor U6855 (N_6855,N_6614,N_6736);
nor U6856 (N_6856,N_6544,N_6737);
and U6857 (N_6857,N_6652,N_6521);
or U6858 (N_6858,N_6589,N_6602);
or U6859 (N_6859,N_6648,N_6676);
and U6860 (N_6860,N_6591,N_6664);
xnor U6861 (N_6861,N_6677,N_6501);
nor U6862 (N_6862,N_6605,N_6670);
nor U6863 (N_6863,N_6686,N_6712);
nand U6864 (N_6864,N_6607,N_6703);
nor U6865 (N_6865,N_6747,N_6729);
nor U6866 (N_6866,N_6580,N_6683);
or U6867 (N_6867,N_6506,N_6578);
xor U6868 (N_6868,N_6634,N_6587);
xor U6869 (N_6869,N_6674,N_6733);
and U6870 (N_6870,N_6675,N_6599);
or U6871 (N_6871,N_6680,N_6717);
and U6872 (N_6872,N_6654,N_6529);
nand U6873 (N_6873,N_6744,N_6504);
and U6874 (N_6874,N_6603,N_6643);
and U6875 (N_6875,N_6640,N_6616);
and U6876 (N_6876,N_6540,N_6657);
nand U6877 (N_6877,N_6532,N_6633);
xnor U6878 (N_6878,N_6716,N_6633);
xnor U6879 (N_6879,N_6671,N_6680);
nand U6880 (N_6880,N_6551,N_6700);
or U6881 (N_6881,N_6505,N_6639);
or U6882 (N_6882,N_6651,N_6664);
nor U6883 (N_6883,N_6579,N_6746);
nor U6884 (N_6884,N_6656,N_6501);
and U6885 (N_6885,N_6655,N_6700);
nor U6886 (N_6886,N_6653,N_6595);
nand U6887 (N_6887,N_6550,N_6680);
nand U6888 (N_6888,N_6632,N_6559);
and U6889 (N_6889,N_6723,N_6605);
and U6890 (N_6890,N_6533,N_6535);
nor U6891 (N_6891,N_6531,N_6677);
xor U6892 (N_6892,N_6532,N_6536);
xor U6893 (N_6893,N_6515,N_6576);
nor U6894 (N_6894,N_6509,N_6629);
or U6895 (N_6895,N_6565,N_6623);
and U6896 (N_6896,N_6605,N_6669);
nor U6897 (N_6897,N_6624,N_6604);
nor U6898 (N_6898,N_6673,N_6556);
and U6899 (N_6899,N_6613,N_6500);
nand U6900 (N_6900,N_6706,N_6715);
or U6901 (N_6901,N_6639,N_6664);
or U6902 (N_6902,N_6611,N_6557);
nand U6903 (N_6903,N_6600,N_6662);
xor U6904 (N_6904,N_6735,N_6619);
or U6905 (N_6905,N_6725,N_6704);
and U6906 (N_6906,N_6702,N_6612);
and U6907 (N_6907,N_6721,N_6543);
nor U6908 (N_6908,N_6599,N_6538);
or U6909 (N_6909,N_6717,N_6603);
xnor U6910 (N_6910,N_6684,N_6621);
nor U6911 (N_6911,N_6630,N_6682);
and U6912 (N_6912,N_6561,N_6577);
xor U6913 (N_6913,N_6653,N_6622);
nor U6914 (N_6914,N_6736,N_6543);
and U6915 (N_6915,N_6527,N_6563);
or U6916 (N_6916,N_6694,N_6551);
xnor U6917 (N_6917,N_6505,N_6744);
and U6918 (N_6918,N_6507,N_6557);
nor U6919 (N_6919,N_6684,N_6513);
or U6920 (N_6920,N_6519,N_6621);
nand U6921 (N_6921,N_6591,N_6571);
nand U6922 (N_6922,N_6573,N_6605);
and U6923 (N_6923,N_6544,N_6666);
or U6924 (N_6924,N_6668,N_6611);
or U6925 (N_6925,N_6546,N_6615);
nand U6926 (N_6926,N_6570,N_6509);
xor U6927 (N_6927,N_6551,N_6617);
and U6928 (N_6928,N_6676,N_6726);
nand U6929 (N_6929,N_6593,N_6674);
nor U6930 (N_6930,N_6645,N_6550);
nand U6931 (N_6931,N_6663,N_6573);
xnor U6932 (N_6932,N_6712,N_6571);
or U6933 (N_6933,N_6507,N_6553);
xor U6934 (N_6934,N_6582,N_6554);
or U6935 (N_6935,N_6574,N_6564);
or U6936 (N_6936,N_6705,N_6551);
and U6937 (N_6937,N_6659,N_6732);
xnor U6938 (N_6938,N_6632,N_6531);
nand U6939 (N_6939,N_6731,N_6725);
nor U6940 (N_6940,N_6666,N_6734);
nor U6941 (N_6941,N_6612,N_6581);
or U6942 (N_6942,N_6741,N_6606);
and U6943 (N_6943,N_6722,N_6539);
nand U6944 (N_6944,N_6635,N_6658);
xnor U6945 (N_6945,N_6688,N_6586);
nand U6946 (N_6946,N_6677,N_6523);
nand U6947 (N_6947,N_6589,N_6539);
nor U6948 (N_6948,N_6732,N_6663);
nor U6949 (N_6949,N_6575,N_6645);
xnor U6950 (N_6950,N_6615,N_6548);
or U6951 (N_6951,N_6561,N_6707);
and U6952 (N_6952,N_6623,N_6546);
xor U6953 (N_6953,N_6602,N_6562);
or U6954 (N_6954,N_6681,N_6718);
or U6955 (N_6955,N_6666,N_6632);
and U6956 (N_6956,N_6736,N_6615);
nand U6957 (N_6957,N_6500,N_6515);
or U6958 (N_6958,N_6722,N_6642);
nor U6959 (N_6959,N_6729,N_6563);
nor U6960 (N_6960,N_6626,N_6678);
or U6961 (N_6961,N_6581,N_6585);
and U6962 (N_6962,N_6684,N_6507);
or U6963 (N_6963,N_6603,N_6700);
and U6964 (N_6964,N_6725,N_6576);
xor U6965 (N_6965,N_6709,N_6554);
or U6966 (N_6966,N_6638,N_6594);
or U6967 (N_6967,N_6543,N_6705);
xor U6968 (N_6968,N_6737,N_6608);
xor U6969 (N_6969,N_6685,N_6601);
and U6970 (N_6970,N_6592,N_6633);
nand U6971 (N_6971,N_6582,N_6693);
nor U6972 (N_6972,N_6695,N_6578);
and U6973 (N_6973,N_6634,N_6641);
nor U6974 (N_6974,N_6714,N_6628);
and U6975 (N_6975,N_6544,N_6645);
nand U6976 (N_6976,N_6620,N_6659);
nor U6977 (N_6977,N_6727,N_6513);
or U6978 (N_6978,N_6556,N_6658);
xor U6979 (N_6979,N_6600,N_6671);
xor U6980 (N_6980,N_6556,N_6687);
nand U6981 (N_6981,N_6691,N_6713);
xor U6982 (N_6982,N_6706,N_6552);
and U6983 (N_6983,N_6603,N_6684);
xnor U6984 (N_6984,N_6695,N_6519);
nand U6985 (N_6985,N_6625,N_6655);
and U6986 (N_6986,N_6701,N_6671);
nor U6987 (N_6987,N_6521,N_6644);
nand U6988 (N_6988,N_6694,N_6720);
nor U6989 (N_6989,N_6629,N_6528);
and U6990 (N_6990,N_6675,N_6728);
xor U6991 (N_6991,N_6668,N_6554);
or U6992 (N_6992,N_6564,N_6749);
and U6993 (N_6993,N_6669,N_6680);
or U6994 (N_6994,N_6605,N_6704);
nor U6995 (N_6995,N_6701,N_6604);
nor U6996 (N_6996,N_6613,N_6733);
xnor U6997 (N_6997,N_6697,N_6623);
nand U6998 (N_6998,N_6669,N_6528);
or U6999 (N_6999,N_6586,N_6661);
xnor U7000 (N_7000,N_6800,N_6775);
xor U7001 (N_7001,N_6856,N_6780);
nand U7002 (N_7002,N_6844,N_6877);
nor U7003 (N_7003,N_6833,N_6823);
and U7004 (N_7004,N_6899,N_6771);
and U7005 (N_7005,N_6778,N_6868);
nor U7006 (N_7006,N_6873,N_6924);
and U7007 (N_7007,N_6818,N_6955);
xor U7008 (N_7008,N_6975,N_6754);
or U7009 (N_7009,N_6984,N_6917);
or U7010 (N_7010,N_6822,N_6841);
xor U7011 (N_7011,N_6836,N_6840);
and U7012 (N_7012,N_6895,N_6769);
and U7013 (N_7013,N_6994,N_6908);
and U7014 (N_7014,N_6959,N_6881);
and U7015 (N_7015,N_6811,N_6750);
nor U7016 (N_7016,N_6862,N_6825);
nor U7017 (N_7017,N_6941,N_6947);
xor U7018 (N_7018,N_6831,N_6922);
or U7019 (N_7019,N_6875,N_6968);
nor U7020 (N_7020,N_6808,N_6867);
or U7021 (N_7021,N_6755,N_6952);
and U7022 (N_7022,N_6929,N_6997);
xnor U7023 (N_7023,N_6909,N_6890);
or U7024 (N_7024,N_6795,N_6979);
or U7025 (N_7025,N_6789,N_6886);
nor U7026 (N_7026,N_6946,N_6779);
and U7027 (N_7027,N_6751,N_6765);
nand U7028 (N_7028,N_6853,N_6949);
xor U7029 (N_7029,N_6848,N_6785);
and U7030 (N_7030,N_6813,N_6781);
and U7031 (N_7031,N_6812,N_6900);
xor U7032 (N_7032,N_6992,N_6962);
nor U7033 (N_7033,N_6907,N_6752);
nand U7034 (N_7034,N_6849,N_6784);
and U7035 (N_7035,N_6884,N_6965);
nor U7036 (N_7036,N_6782,N_6887);
xnor U7037 (N_7037,N_6893,N_6869);
nand U7038 (N_7038,N_6816,N_6878);
nor U7039 (N_7039,N_6827,N_6918);
nor U7040 (N_7040,N_6871,N_6933);
and U7041 (N_7041,N_6763,N_6966);
xor U7042 (N_7042,N_6891,N_6806);
nor U7043 (N_7043,N_6989,N_6903);
xnor U7044 (N_7044,N_6961,N_6934);
and U7045 (N_7045,N_6858,N_6936);
nor U7046 (N_7046,N_6972,N_6842);
or U7047 (N_7047,N_6894,N_6896);
or U7048 (N_7048,N_6969,N_6931);
nor U7049 (N_7049,N_6801,N_6912);
nand U7050 (N_7050,N_6993,N_6981);
nand U7051 (N_7051,N_6998,N_6974);
nand U7052 (N_7052,N_6930,N_6817);
or U7053 (N_7053,N_6815,N_6950);
nor U7054 (N_7054,N_6788,N_6857);
and U7055 (N_7055,N_6851,N_6926);
nor U7056 (N_7056,N_6945,N_6938);
xnor U7057 (N_7057,N_6988,N_6980);
nor U7058 (N_7058,N_6939,N_6953);
and U7059 (N_7059,N_6753,N_6935);
nor U7060 (N_7060,N_6843,N_6882);
and U7061 (N_7061,N_6810,N_6995);
and U7062 (N_7062,N_6977,N_6971);
or U7063 (N_7063,N_6872,N_6864);
or U7064 (N_7064,N_6797,N_6940);
and U7065 (N_7065,N_6906,N_6927);
nor U7066 (N_7066,N_6892,N_6824);
nor U7067 (N_7067,N_6913,N_6983);
and U7068 (N_7068,N_6804,N_6866);
nand U7069 (N_7069,N_6865,N_6879);
xor U7070 (N_7070,N_6976,N_6990);
or U7071 (N_7071,N_6796,N_6777);
nor U7072 (N_7072,N_6863,N_6897);
nand U7073 (N_7073,N_6846,N_6803);
nand U7074 (N_7074,N_6957,N_6883);
xnor U7075 (N_7075,N_6898,N_6932);
or U7076 (N_7076,N_6942,N_6854);
nand U7077 (N_7077,N_6986,N_6985);
xor U7078 (N_7078,N_6889,N_6870);
and U7079 (N_7079,N_6855,N_6772);
nand U7080 (N_7080,N_6911,N_6805);
xnor U7081 (N_7081,N_6834,N_6764);
nor U7082 (N_7082,N_6809,N_6910);
xnor U7083 (N_7083,N_6845,N_6814);
nor U7084 (N_7084,N_6821,N_6861);
and U7085 (N_7085,N_6759,N_6919);
nand U7086 (N_7086,N_6991,N_6916);
xor U7087 (N_7087,N_6850,N_6790);
and U7088 (N_7088,N_6960,N_6830);
xor U7089 (N_7089,N_6958,N_6937);
nor U7090 (N_7090,N_6905,N_6786);
and U7091 (N_7091,N_6923,N_6774);
and U7092 (N_7092,N_6928,N_6967);
or U7093 (N_7093,N_6837,N_6920);
or U7094 (N_7094,N_6982,N_6915);
or U7095 (N_7095,N_6847,N_6787);
nand U7096 (N_7096,N_6948,N_6792);
xnor U7097 (N_7097,N_6757,N_6852);
and U7098 (N_7098,N_6888,N_6885);
nand U7099 (N_7099,N_6860,N_6839);
and U7100 (N_7100,N_6859,N_6767);
or U7101 (N_7101,N_6970,N_6838);
nor U7102 (N_7102,N_6880,N_6987);
or U7103 (N_7103,N_6761,N_6762);
xnor U7104 (N_7104,N_6951,N_6826);
xor U7105 (N_7105,N_6791,N_6996);
nor U7106 (N_7106,N_6819,N_6954);
nand U7107 (N_7107,N_6758,N_6921);
or U7108 (N_7108,N_6832,N_6768);
and U7109 (N_7109,N_6876,N_6798);
xor U7110 (N_7110,N_6999,N_6944);
nand U7111 (N_7111,N_6807,N_6799);
nand U7112 (N_7112,N_6963,N_6901);
or U7113 (N_7113,N_6835,N_6828);
xnor U7114 (N_7114,N_6978,N_6973);
or U7115 (N_7115,N_6770,N_6914);
and U7116 (N_7116,N_6756,N_6874);
and U7117 (N_7117,N_6829,N_6793);
or U7118 (N_7118,N_6902,N_6760);
nor U7119 (N_7119,N_6964,N_6802);
nor U7120 (N_7120,N_6820,N_6956);
or U7121 (N_7121,N_6783,N_6904);
or U7122 (N_7122,N_6925,N_6776);
and U7123 (N_7123,N_6773,N_6943);
nand U7124 (N_7124,N_6766,N_6794);
xnor U7125 (N_7125,N_6750,N_6785);
xor U7126 (N_7126,N_6791,N_6926);
or U7127 (N_7127,N_6983,N_6825);
xnor U7128 (N_7128,N_6906,N_6928);
nor U7129 (N_7129,N_6905,N_6964);
nand U7130 (N_7130,N_6951,N_6901);
xor U7131 (N_7131,N_6830,N_6867);
nand U7132 (N_7132,N_6807,N_6886);
or U7133 (N_7133,N_6826,N_6838);
and U7134 (N_7134,N_6790,N_6811);
nor U7135 (N_7135,N_6954,N_6772);
xnor U7136 (N_7136,N_6811,N_6950);
xor U7137 (N_7137,N_6809,N_6987);
xor U7138 (N_7138,N_6883,N_6843);
xnor U7139 (N_7139,N_6980,N_6831);
or U7140 (N_7140,N_6819,N_6991);
nand U7141 (N_7141,N_6843,N_6970);
and U7142 (N_7142,N_6973,N_6972);
xor U7143 (N_7143,N_6767,N_6757);
xor U7144 (N_7144,N_6766,N_6885);
nor U7145 (N_7145,N_6930,N_6851);
nand U7146 (N_7146,N_6856,N_6942);
or U7147 (N_7147,N_6915,N_6952);
nand U7148 (N_7148,N_6758,N_6824);
nor U7149 (N_7149,N_6885,N_6826);
nand U7150 (N_7150,N_6999,N_6822);
xor U7151 (N_7151,N_6788,N_6923);
or U7152 (N_7152,N_6982,N_6847);
nand U7153 (N_7153,N_6780,N_6884);
xnor U7154 (N_7154,N_6853,N_6788);
xor U7155 (N_7155,N_6967,N_6921);
nand U7156 (N_7156,N_6951,N_6961);
or U7157 (N_7157,N_6814,N_6770);
or U7158 (N_7158,N_6919,N_6837);
or U7159 (N_7159,N_6785,N_6825);
and U7160 (N_7160,N_6926,N_6865);
nor U7161 (N_7161,N_6820,N_6816);
or U7162 (N_7162,N_6787,N_6931);
nor U7163 (N_7163,N_6919,N_6814);
or U7164 (N_7164,N_6942,N_6772);
nand U7165 (N_7165,N_6878,N_6834);
nor U7166 (N_7166,N_6896,N_6962);
and U7167 (N_7167,N_6968,N_6928);
xor U7168 (N_7168,N_6755,N_6864);
or U7169 (N_7169,N_6784,N_6965);
and U7170 (N_7170,N_6881,N_6901);
nand U7171 (N_7171,N_6832,N_6997);
and U7172 (N_7172,N_6932,N_6824);
and U7173 (N_7173,N_6758,N_6815);
and U7174 (N_7174,N_6808,N_6766);
or U7175 (N_7175,N_6966,N_6847);
nor U7176 (N_7176,N_6946,N_6764);
xor U7177 (N_7177,N_6806,N_6874);
and U7178 (N_7178,N_6811,N_6942);
xnor U7179 (N_7179,N_6779,N_6943);
nand U7180 (N_7180,N_6909,N_6771);
xnor U7181 (N_7181,N_6999,N_6869);
or U7182 (N_7182,N_6953,N_6823);
or U7183 (N_7183,N_6852,N_6921);
and U7184 (N_7184,N_6918,N_6787);
nand U7185 (N_7185,N_6761,N_6906);
nand U7186 (N_7186,N_6856,N_6866);
and U7187 (N_7187,N_6778,N_6921);
nand U7188 (N_7188,N_6947,N_6885);
xor U7189 (N_7189,N_6999,N_6904);
or U7190 (N_7190,N_6896,N_6902);
nand U7191 (N_7191,N_6783,N_6862);
or U7192 (N_7192,N_6755,N_6862);
nor U7193 (N_7193,N_6869,N_6820);
nor U7194 (N_7194,N_6832,N_6931);
and U7195 (N_7195,N_6779,N_6970);
nand U7196 (N_7196,N_6774,N_6754);
nor U7197 (N_7197,N_6863,N_6850);
or U7198 (N_7198,N_6851,N_6857);
nor U7199 (N_7199,N_6778,N_6886);
or U7200 (N_7200,N_6953,N_6980);
nor U7201 (N_7201,N_6751,N_6786);
nand U7202 (N_7202,N_6856,N_6996);
or U7203 (N_7203,N_6758,N_6853);
or U7204 (N_7204,N_6752,N_6951);
nor U7205 (N_7205,N_6872,N_6924);
nor U7206 (N_7206,N_6934,N_6969);
nand U7207 (N_7207,N_6801,N_6829);
or U7208 (N_7208,N_6753,N_6795);
and U7209 (N_7209,N_6952,N_6825);
and U7210 (N_7210,N_6922,N_6815);
nor U7211 (N_7211,N_6919,N_6933);
xnor U7212 (N_7212,N_6802,N_6839);
nand U7213 (N_7213,N_6798,N_6944);
xor U7214 (N_7214,N_6750,N_6859);
nand U7215 (N_7215,N_6958,N_6984);
nor U7216 (N_7216,N_6790,N_6899);
nor U7217 (N_7217,N_6901,N_6985);
and U7218 (N_7218,N_6954,N_6955);
xor U7219 (N_7219,N_6766,N_6929);
and U7220 (N_7220,N_6909,N_6950);
and U7221 (N_7221,N_6781,N_6807);
nor U7222 (N_7222,N_6769,N_6995);
or U7223 (N_7223,N_6814,N_6826);
and U7224 (N_7224,N_6762,N_6984);
xor U7225 (N_7225,N_6764,N_6817);
or U7226 (N_7226,N_6880,N_6940);
xnor U7227 (N_7227,N_6755,N_6795);
nand U7228 (N_7228,N_6871,N_6962);
nand U7229 (N_7229,N_6984,N_6814);
nor U7230 (N_7230,N_6967,N_6948);
nand U7231 (N_7231,N_6975,N_6920);
or U7232 (N_7232,N_6909,N_6986);
nand U7233 (N_7233,N_6809,N_6758);
xnor U7234 (N_7234,N_6999,N_6952);
nor U7235 (N_7235,N_6858,N_6841);
nor U7236 (N_7236,N_6831,N_6889);
nor U7237 (N_7237,N_6836,N_6796);
nand U7238 (N_7238,N_6911,N_6774);
xor U7239 (N_7239,N_6915,N_6825);
nor U7240 (N_7240,N_6953,N_6765);
nor U7241 (N_7241,N_6894,N_6883);
nand U7242 (N_7242,N_6761,N_6914);
nor U7243 (N_7243,N_6819,N_6818);
nor U7244 (N_7244,N_6941,N_6876);
nand U7245 (N_7245,N_6943,N_6847);
nor U7246 (N_7246,N_6893,N_6970);
xnor U7247 (N_7247,N_6927,N_6980);
and U7248 (N_7248,N_6897,N_6867);
and U7249 (N_7249,N_6801,N_6765);
and U7250 (N_7250,N_7021,N_7046);
or U7251 (N_7251,N_7075,N_7143);
or U7252 (N_7252,N_7040,N_7242);
xor U7253 (N_7253,N_7036,N_7224);
and U7254 (N_7254,N_7200,N_7178);
nor U7255 (N_7255,N_7082,N_7135);
nand U7256 (N_7256,N_7035,N_7227);
xnor U7257 (N_7257,N_7188,N_7017);
or U7258 (N_7258,N_7030,N_7213);
nor U7259 (N_7259,N_7194,N_7151);
nor U7260 (N_7260,N_7105,N_7175);
nor U7261 (N_7261,N_7195,N_7013);
xor U7262 (N_7262,N_7235,N_7187);
nor U7263 (N_7263,N_7064,N_7146);
and U7264 (N_7264,N_7005,N_7083);
or U7265 (N_7265,N_7173,N_7093);
or U7266 (N_7266,N_7184,N_7215);
nand U7267 (N_7267,N_7055,N_7160);
and U7268 (N_7268,N_7069,N_7009);
nand U7269 (N_7269,N_7057,N_7027);
nand U7270 (N_7270,N_7152,N_7060);
and U7271 (N_7271,N_7204,N_7140);
nor U7272 (N_7272,N_7061,N_7050);
nand U7273 (N_7273,N_7123,N_7201);
xnor U7274 (N_7274,N_7206,N_7147);
xor U7275 (N_7275,N_7172,N_7164);
nor U7276 (N_7276,N_7033,N_7232);
xnor U7277 (N_7277,N_7098,N_7159);
nand U7278 (N_7278,N_7216,N_7211);
xor U7279 (N_7279,N_7228,N_7220);
nand U7280 (N_7280,N_7113,N_7192);
and U7281 (N_7281,N_7249,N_7170);
and U7282 (N_7282,N_7053,N_7209);
nor U7283 (N_7283,N_7104,N_7052);
nand U7284 (N_7284,N_7047,N_7189);
nand U7285 (N_7285,N_7071,N_7087);
and U7286 (N_7286,N_7226,N_7106);
and U7287 (N_7287,N_7212,N_7118);
or U7288 (N_7288,N_7205,N_7117);
or U7289 (N_7289,N_7020,N_7028);
nor U7290 (N_7290,N_7086,N_7144);
nor U7291 (N_7291,N_7202,N_7089);
nand U7292 (N_7292,N_7002,N_7092);
nor U7293 (N_7293,N_7121,N_7007);
nor U7294 (N_7294,N_7241,N_7223);
and U7295 (N_7295,N_7230,N_7066);
nor U7296 (N_7296,N_7243,N_7240);
xnor U7297 (N_7297,N_7179,N_7034);
xor U7298 (N_7298,N_7132,N_7122);
xor U7299 (N_7299,N_7088,N_7029);
nand U7300 (N_7300,N_7072,N_7153);
nand U7301 (N_7301,N_7186,N_7039);
nor U7302 (N_7302,N_7207,N_7077);
nor U7303 (N_7303,N_7142,N_7131);
nand U7304 (N_7304,N_7091,N_7129);
or U7305 (N_7305,N_7001,N_7191);
xnor U7306 (N_7306,N_7183,N_7095);
nor U7307 (N_7307,N_7124,N_7246);
and U7308 (N_7308,N_7080,N_7222);
or U7309 (N_7309,N_7141,N_7137);
or U7310 (N_7310,N_7011,N_7081);
xnor U7311 (N_7311,N_7166,N_7058);
and U7312 (N_7312,N_7176,N_7127);
and U7313 (N_7313,N_7218,N_7031);
nand U7314 (N_7314,N_7138,N_7010);
nand U7315 (N_7315,N_7196,N_7062);
nor U7316 (N_7316,N_7169,N_7210);
nand U7317 (N_7317,N_7026,N_7155);
nand U7318 (N_7318,N_7233,N_7168);
nand U7319 (N_7319,N_7162,N_7015);
nand U7320 (N_7320,N_7156,N_7090);
and U7321 (N_7321,N_7024,N_7059);
or U7322 (N_7322,N_7110,N_7041);
nor U7323 (N_7323,N_7076,N_7203);
nand U7324 (N_7324,N_7070,N_7139);
or U7325 (N_7325,N_7000,N_7133);
nand U7326 (N_7326,N_7084,N_7161);
nand U7327 (N_7327,N_7119,N_7073);
nor U7328 (N_7328,N_7180,N_7208);
or U7329 (N_7329,N_7229,N_7044);
and U7330 (N_7330,N_7016,N_7068);
and U7331 (N_7331,N_7217,N_7096);
xor U7332 (N_7332,N_7056,N_7120);
or U7333 (N_7333,N_7219,N_7148);
or U7334 (N_7334,N_7198,N_7103);
nand U7335 (N_7335,N_7145,N_7163);
and U7336 (N_7336,N_7025,N_7149);
nand U7337 (N_7337,N_7126,N_7185);
xor U7338 (N_7338,N_7038,N_7048);
and U7339 (N_7339,N_7023,N_7221);
xnor U7340 (N_7340,N_7049,N_7190);
or U7341 (N_7341,N_7174,N_7125);
nor U7342 (N_7342,N_7004,N_7136);
nand U7343 (N_7343,N_7134,N_7022);
nand U7344 (N_7344,N_7054,N_7157);
nand U7345 (N_7345,N_7158,N_7100);
xnor U7346 (N_7346,N_7003,N_7085);
nand U7347 (N_7347,N_7236,N_7012);
or U7348 (N_7348,N_7079,N_7074);
xnor U7349 (N_7349,N_7182,N_7177);
or U7350 (N_7350,N_7045,N_7101);
and U7351 (N_7351,N_7231,N_7115);
xor U7352 (N_7352,N_7042,N_7193);
or U7353 (N_7353,N_7063,N_7019);
or U7354 (N_7354,N_7006,N_7237);
nor U7355 (N_7355,N_7165,N_7014);
nor U7356 (N_7356,N_7130,N_7065);
and U7357 (N_7357,N_7248,N_7108);
xnor U7358 (N_7358,N_7171,N_7051);
and U7359 (N_7359,N_7109,N_7225);
nor U7360 (N_7360,N_7234,N_7239);
and U7361 (N_7361,N_7094,N_7078);
and U7362 (N_7362,N_7247,N_7097);
or U7363 (N_7363,N_7154,N_7244);
nor U7364 (N_7364,N_7102,N_7197);
nor U7365 (N_7365,N_7116,N_7167);
or U7366 (N_7366,N_7067,N_7111);
nor U7367 (N_7367,N_7107,N_7032);
nand U7368 (N_7368,N_7037,N_7238);
and U7369 (N_7369,N_7008,N_7018);
xor U7370 (N_7370,N_7128,N_7099);
xor U7371 (N_7371,N_7043,N_7114);
or U7372 (N_7372,N_7150,N_7112);
or U7373 (N_7373,N_7214,N_7245);
nor U7374 (N_7374,N_7181,N_7199);
or U7375 (N_7375,N_7245,N_7069);
or U7376 (N_7376,N_7074,N_7168);
or U7377 (N_7377,N_7130,N_7181);
nand U7378 (N_7378,N_7097,N_7042);
nand U7379 (N_7379,N_7123,N_7137);
xnor U7380 (N_7380,N_7061,N_7228);
nand U7381 (N_7381,N_7192,N_7041);
or U7382 (N_7382,N_7003,N_7110);
xnor U7383 (N_7383,N_7132,N_7071);
nor U7384 (N_7384,N_7168,N_7098);
or U7385 (N_7385,N_7219,N_7194);
xor U7386 (N_7386,N_7086,N_7081);
and U7387 (N_7387,N_7170,N_7202);
and U7388 (N_7388,N_7222,N_7129);
nand U7389 (N_7389,N_7077,N_7055);
or U7390 (N_7390,N_7234,N_7186);
nor U7391 (N_7391,N_7238,N_7155);
xnor U7392 (N_7392,N_7072,N_7120);
nand U7393 (N_7393,N_7178,N_7029);
and U7394 (N_7394,N_7094,N_7013);
or U7395 (N_7395,N_7030,N_7072);
or U7396 (N_7396,N_7058,N_7127);
and U7397 (N_7397,N_7054,N_7051);
xor U7398 (N_7398,N_7163,N_7092);
and U7399 (N_7399,N_7205,N_7188);
xnor U7400 (N_7400,N_7080,N_7218);
nand U7401 (N_7401,N_7167,N_7031);
nor U7402 (N_7402,N_7143,N_7169);
or U7403 (N_7403,N_7071,N_7206);
nor U7404 (N_7404,N_7034,N_7027);
xnor U7405 (N_7405,N_7055,N_7017);
and U7406 (N_7406,N_7093,N_7003);
nand U7407 (N_7407,N_7149,N_7043);
nor U7408 (N_7408,N_7197,N_7117);
or U7409 (N_7409,N_7010,N_7091);
or U7410 (N_7410,N_7163,N_7085);
nor U7411 (N_7411,N_7228,N_7109);
xnor U7412 (N_7412,N_7134,N_7025);
and U7413 (N_7413,N_7040,N_7154);
xnor U7414 (N_7414,N_7138,N_7227);
xor U7415 (N_7415,N_7093,N_7105);
nor U7416 (N_7416,N_7175,N_7107);
and U7417 (N_7417,N_7153,N_7082);
xor U7418 (N_7418,N_7046,N_7206);
xor U7419 (N_7419,N_7132,N_7053);
and U7420 (N_7420,N_7222,N_7233);
or U7421 (N_7421,N_7134,N_7157);
or U7422 (N_7422,N_7079,N_7086);
nand U7423 (N_7423,N_7011,N_7077);
and U7424 (N_7424,N_7109,N_7074);
nor U7425 (N_7425,N_7002,N_7039);
nand U7426 (N_7426,N_7041,N_7179);
or U7427 (N_7427,N_7131,N_7103);
nor U7428 (N_7428,N_7036,N_7148);
nor U7429 (N_7429,N_7052,N_7127);
and U7430 (N_7430,N_7095,N_7208);
xnor U7431 (N_7431,N_7202,N_7173);
xnor U7432 (N_7432,N_7207,N_7124);
nand U7433 (N_7433,N_7230,N_7136);
or U7434 (N_7434,N_7197,N_7199);
or U7435 (N_7435,N_7185,N_7053);
or U7436 (N_7436,N_7121,N_7014);
xnor U7437 (N_7437,N_7059,N_7034);
or U7438 (N_7438,N_7141,N_7179);
nor U7439 (N_7439,N_7132,N_7003);
or U7440 (N_7440,N_7161,N_7055);
nor U7441 (N_7441,N_7191,N_7021);
and U7442 (N_7442,N_7130,N_7168);
and U7443 (N_7443,N_7232,N_7193);
nand U7444 (N_7444,N_7077,N_7140);
nor U7445 (N_7445,N_7147,N_7042);
and U7446 (N_7446,N_7004,N_7087);
and U7447 (N_7447,N_7157,N_7211);
and U7448 (N_7448,N_7071,N_7106);
nor U7449 (N_7449,N_7221,N_7150);
xor U7450 (N_7450,N_7022,N_7040);
xnor U7451 (N_7451,N_7119,N_7078);
nand U7452 (N_7452,N_7131,N_7118);
nor U7453 (N_7453,N_7063,N_7240);
xor U7454 (N_7454,N_7002,N_7061);
nor U7455 (N_7455,N_7111,N_7093);
or U7456 (N_7456,N_7170,N_7220);
nand U7457 (N_7457,N_7223,N_7235);
and U7458 (N_7458,N_7224,N_7079);
and U7459 (N_7459,N_7147,N_7214);
or U7460 (N_7460,N_7077,N_7200);
and U7461 (N_7461,N_7028,N_7093);
nor U7462 (N_7462,N_7089,N_7112);
and U7463 (N_7463,N_7093,N_7110);
or U7464 (N_7464,N_7228,N_7219);
or U7465 (N_7465,N_7219,N_7039);
or U7466 (N_7466,N_7182,N_7214);
nor U7467 (N_7467,N_7029,N_7246);
and U7468 (N_7468,N_7070,N_7001);
nand U7469 (N_7469,N_7095,N_7172);
nor U7470 (N_7470,N_7197,N_7146);
nand U7471 (N_7471,N_7101,N_7077);
nor U7472 (N_7472,N_7191,N_7079);
nand U7473 (N_7473,N_7199,N_7184);
or U7474 (N_7474,N_7150,N_7214);
nand U7475 (N_7475,N_7073,N_7122);
nor U7476 (N_7476,N_7021,N_7105);
nand U7477 (N_7477,N_7248,N_7081);
nand U7478 (N_7478,N_7178,N_7106);
xnor U7479 (N_7479,N_7145,N_7056);
and U7480 (N_7480,N_7086,N_7029);
xor U7481 (N_7481,N_7055,N_7165);
and U7482 (N_7482,N_7221,N_7218);
nand U7483 (N_7483,N_7063,N_7101);
and U7484 (N_7484,N_7079,N_7013);
and U7485 (N_7485,N_7064,N_7029);
xnor U7486 (N_7486,N_7088,N_7126);
nand U7487 (N_7487,N_7246,N_7151);
nand U7488 (N_7488,N_7014,N_7190);
nand U7489 (N_7489,N_7023,N_7099);
xor U7490 (N_7490,N_7044,N_7234);
xor U7491 (N_7491,N_7219,N_7193);
nor U7492 (N_7492,N_7042,N_7000);
xnor U7493 (N_7493,N_7235,N_7131);
or U7494 (N_7494,N_7077,N_7144);
nor U7495 (N_7495,N_7043,N_7193);
and U7496 (N_7496,N_7121,N_7235);
and U7497 (N_7497,N_7071,N_7123);
nand U7498 (N_7498,N_7011,N_7197);
nor U7499 (N_7499,N_7040,N_7157);
or U7500 (N_7500,N_7294,N_7465);
or U7501 (N_7501,N_7468,N_7428);
nor U7502 (N_7502,N_7487,N_7474);
nand U7503 (N_7503,N_7331,N_7356);
and U7504 (N_7504,N_7398,N_7414);
xnor U7505 (N_7505,N_7385,N_7288);
nor U7506 (N_7506,N_7390,N_7399);
xnor U7507 (N_7507,N_7381,N_7473);
or U7508 (N_7508,N_7490,N_7302);
nand U7509 (N_7509,N_7289,N_7253);
or U7510 (N_7510,N_7478,N_7342);
xnor U7511 (N_7511,N_7327,N_7433);
or U7512 (N_7512,N_7459,N_7497);
and U7513 (N_7513,N_7306,N_7361);
nand U7514 (N_7514,N_7257,N_7328);
xnor U7515 (N_7515,N_7427,N_7431);
or U7516 (N_7516,N_7282,N_7285);
nor U7517 (N_7517,N_7434,N_7469);
xor U7518 (N_7518,N_7470,N_7362);
or U7519 (N_7519,N_7418,N_7426);
or U7520 (N_7520,N_7295,N_7365);
and U7521 (N_7521,N_7498,N_7326);
nor U7522 (N_7522,N_7379,N_7376);
or U7523 (N_7523,N_7476,N_7348);
nor U7524 (N_7524,N_7271,N_7273);
xor U7525 (N_7525,N_7287,N_7453);
or U7526 (N_7526,N_7401,N_7364);
and U7527 (N_7527,N_7413,N_7318);
xor U7528 (N_7528,N_7296,N_7344);
nor U7529 (N_7529,N_7472,N_7486);
or U7530 (N_7530,N_7353,N_7442);
or U7531 (N_7531,N_7395,N_7304);
nand U7532 (N_7532,N_7264,N_7384);
or U7533 (N_7533,N_7373,N_7281);
and U7534 (N_7534,N_7258,N_7254);
nand U7535 (N_7535,N_7305,N_7340);
xor U7536 (N_7536,N_7492,N_7466);
xor U7537 (N_7537,N_7320,N_7307);
and U7538 (N_7538,N_7443,N_7420);
nand U7539 (N_7539,N_7491,N_7449);
or U7540 (N_7540,N_7280,N_7463);
and U7541 (N_7541,N_7316,N_7485);
xor U7542 (N_7542,N_7338,N_7360);
nand U7543 (N_7543,N_7461,N_7321);
xor U7544 (N_7544,N_7421,N_7341);
and U7545 (N_7545,N_7354,N_7494);
or U7546 (N_7546,N_7496,N_7419);
nand U7547 (N_7547,N_7343,N_7283);
and U7548 (N_7548,N_7475,N_7479);
nor U7549 (N_7549,N_7435,N_7455);
nand U7550 (N_7550,N_7268,N_7436);
nor U7551 (N_7551,N_7299,N_7339);
nor U7552 (N_7552,N_7432,N_7284);
xor U7553 (N_7553,N_7363,N_7383);
xnor U7554 (N_7554,N_7286,N_7368);
xnor U7555 (N_7555,N_7265,N_7448);
and U7556 (N_7556,N_7293,N_7270);
and U7557 (N_7557,N_7392,N_7300);
nand U7558 (N_7558,N_7336,N_7346);
nand U7559 (N_7559,N_7425,N_7409);
nand U7560 (N_7560,N_7489,N_7447);
or U7561 (N_7561,N_7324,N_7255);
nor U7562 (N_7562,N_7349,N_7292);
nand U7563 (N_7563,N_7256,N_7276);
or U7564 (N_7564,N_7404,N_7386);
and U7565 (N_7565,N_7450,N_7329);
or U7566 (N_7566,N_7317,N_7277);
nand U7567 (N_7567,N_7275,N_7488);
xnor U7568 (N_7568,N_7266,N_7400);
and U7569 (N_7569,N_7388,N_7272);
or U7570 (N_7570,N_7355,N_7405);
nand U7571 (N_7571,N_7347,N_7402);
nand U7572 (N_7572,N_7499,N_7345);
nor U7573 (N_7573,N_7462,N_7290);
and U7574 (N_7574,N_7367,N_7484);
nand U7575 (N_7575,N_7279,N_7250);
nor U7576 (N_7576,N_7263,N_7335);
and U7577 (N_7577,N_7359,N_7334);
and U7578 (N_7578,N_7387,N_7325);
xnor U7579 (N_7579,N_7274,N_7482);
nor U7580 (N_7580,N_7262,N_7378);
or U7581 (N_7581,N_7417,N_7471);
xnor U7582 (N_7582,N_7407,N_7410);
and U7583 (N_7583,N_7358,N_7323);
and U7584 (N_7584,N_7456,N_7481);
xnor U7585 (N_7585,N_7445,N_7394);
nor U7586 (N_7586,N_7308,N_7454);
and U7587 (N_7587,N_7429,N_7406);
xor U7588 (N_7588,N_7393,N_7416);
nor U7589 (N_7589,N_7391,N_7333);
or U7590 (N_7590,N_7440,N_7446);
xor U7591 (N_7591,N_7444,N_7350);
xnor U7592 (N_7592,N_7252,N_7441);
xnor U7593 (N_7593,N_7422,N_7439);
nand U7594 (N_7594,N_7389,N_7424);
nand U7595 (N_7595,N_7311,N_7337);
nor U7596 (N_7596,N_7403,N_7467);
nor U7597 (N_7597,N_7313,N_7291);
xor U7598 (N_7598,N_7251,N_7310);
nand U7599 (N_7599,N_7412,N_7480);
or U7600 (N_7600,N_7372,N_7259);
and U7601 (N_7601,N_7303,N_7375);
nor U7602 (N_7602,N_7269,N_7477);
xor U7603 (N_7603,N_7408,N_7458);
and U7604 (N_7604,N_7322,N_7411);
nand U7605 (N_7605,N_7382,N_7493);
nor U7606 (N_7606,N_7301,N_7396);
nand U7607 (N_7607,N_7374,N_7278);
xnor U7608 (N_7608,N_7415,N_7437);
nand U7609 (N_7609,N_7423,N_7366);
xnor U7610 (N_7610,N_7332,N_7451);
or U7611 (N_7611,N_7371,N_7438);
xor U7612 (N_7612,N_7430,N_7312);
nand U7613 (N_7613,N_7483,N_7298);
xnor U7614 (N_7614,N_7261,N_7351);
xor U7615 (N_7615,N_7309,N_7460);
nand U7616 (N_7616,N_7370,N_7330);
or U7617 (N_7617,N_7297,N_7357);
or U7618 (N_7618,N_7377,N_7319);
nor U7619 (N_7619,N_7369,N_7314);
xnor U7620 (N_7620,N_7397,N_7495);
nor U7621 (N_7621,N_7260,N_7452);
nand U7622 (N_7622,N_7457,N_7267);
or U7623 (N_7623,N_7380,N_7315);
and U7624 (N_7624,N_7464,N_7352);
nand U7625 (N_7625,N_7417,N_7357);
or U7626 (N_7626,N_7439,N_7348);
or U7627 (N_7627,N_7432,N_7435);
or U7628 (N_7628,N_7456,N_7273);
nand U7629 (N_7629,N_7480,N_7495);
xor U7630 (N_7630,N_7418,N_7436);
nor U7631 (N_7631,N_7290,N_7388);
nand U7632 (N_7632,N_7254,N_7404);
or U7633 (N_7633,N_7459,N_7433);
nor U7634 (N_7634,N_7484,N_7395);
nand U7635 (N_7635,N_7418,N_7391);
and U7636 (N_7636,N_7444,N_7307);
or U7637 (N_7637,N_7311,N_7406);
nor U7638 (N_7638,N_7455,N_7432);
nor U7639 (N_7639,N_7436,N_7479);
xor U7640 (N_7640,N_7349,N_7311);
or U7641 (N_7641,N_7421,N_7443);
nor U7642 (N_7642,N_7395,N_7298);
nor U7643 (N_7643,N_7468,N_7320);
xnor U7644 (N_7644,N_7280,N_7427);
and U7645 (N_7645,N_7446,N_7268);
nand U7646 (N_7646,N_7482,N_7286);
nor U7647 (N_7647,N_7391,N_7294);
xnor U7648 (N_7648,N_7389,N_7475);
xnor U7649 (N_7649,N_7325,N_7486);
xor U7650 (N_7650,N_7368,N_7303);
nand U7651 (N_7651,N_7496,N_7256);
and U7652 (N_7652,N_7420,N_7467);
or U7653 (N_7653,N_7496,N_7327);
nor U7654 (N_7654,N_7323,N_7451);
xor U7655 (N_7655,N_7328,N_7250);
nor U7656 (N_7656,N_7485,N_7426);
nor U7657 (N_7657,N_7384,N_7493);
and U7658 (N_7658,N_7494,N_7459);
xnor U7659 (N_7659,N_7338,N_7442);
nand U7660 (N_7660,N_7305,N_7496);
nand U7661 (N_7661,N_7325,N_7345);
xor U7662 (N_7662,N_7419,N_7457);
and U7663 (N_7663,N_7349,N_7470);
nor U7664 (N_7664,N_7272,N_7355);
or U7665 (N_7665,N_7351,N_7432);
nor U7666 (N_7666,N_7392,N_7363);
nor U7667 (N_7667,N_7375,N_7464);
or U7668 (N_7668,N_7402,N_7290);
or U7669 (N_7669,N_7470,N_7364);
and U7670 (N_7670,N_7289,N_7432);
or U7671 (N_7671,N_7337,N_7499);
nand U7672 (N_7672,N_7376,N_7271);
xor U7673 (N_7673,N_7339,N_7301);
or U7674 (N_7674,N_7385,N_7278);
nand U7675 (N_7675,N_7468,N_7436);
nand U7676 (N_7676,N_7362,N_7348);
or U7677 (N_7677,N_7268,N_7428);
nor U7678 (N_7678,N_7394,N_7448);
and U7679 (N_7679,N_7392,N_7478);
nor U7680 (N_7680,N_7425,N_7449);
nor U7681 (N_7681,N_7490,N_7337);
and U7682 (N_7682,N_7342,N_7251);
nor U7683 (N_7683,N_7282,N_7312);
xnor U7684 (N_7684,N_7413,N_7287);
nor U7685 (N_7685,N_7452,N_7481);
and U7686 (N_7686,N_7379,N_7368);
nor U7687 (N_7687,N_7400,N_7457);
nand U7688 (N_7688,N_7481,N_7401);
xnor U7689 (N_7689,N_7274,N_7432);
nor U7690 (N_7690,N_7308,N_7279);
and U7691 (N_7691,N_7410,N_7438);
or U7692 (N_7692,N_7335,N_7271);
and U7693 (N_7693,N_7387,N_7349);
nor U7694 (N_7694,N_7298,N_7256);
xnor U7695 (N_7695,N_7339,N_7427);
nor U7696 (N_7696,N_7255,N_7394);
or U7697 (N_7697,N_7352,N_7277);
nand U7698 (N_7698,N_7311,N_7250);
xnor U7699 (N_7699,N_7253,N_7267);
and U7700 (N_7700,N_7271,N_7452);
nor U7701 (N_7701,N_7394,N_7306);
xnor U7702 (N_7702,N_7391,N_7460);
nor U7703 (N_7703,N_7390,N_7382);
or U7704 (N_7704,N_7452,N_7339);
nor U7705 (N_7705,N_7397,N_7412);
or U7706 (N_7706,N_7290,N_7332);
or U7707 (N_7707,N_7470,N_7258);
or U7708 (N_7708,N_7255,N_7448);
nand U7709 (N_7709,N_7446,N_7262);
and U7710 (N_7710,N_7396,N_7430);
and U7711 (N_7711,N_7469,N_7333);
nand U7712 (N_7712,N_7409,N_7347);
or U7713 (N_7713,N_7341,N_7371);
or U7714 (N_7714,N_7297,N_7480);
xnor U7715 (N_7715,N_7389,N_7365);
xor U7716 (N_7716,N_7373,N_7382);
xor U7717 (N_7717,N_7269,N_7474);
nand U7718 (N_7718,N_7369,N_7269);
nor U7719 (N_7719,N_7349,N_7328);
and U7720 (N_7720,N_7488,N_7268);
nor U7721 (N_7721,N_7415,N_7461);
xor U7722 (N_7722,N_7381,N_7398);
or U7723 (N_7723,N_7267,N_7464);
nand U7724 (N_7724,N_7415,N_7439);
and U7725 (N_7725,N_7412,N_7304);
or U7726 (N_7726,N_7480,N_7404);
nor U7727 (N_7727,N_7331,N_7253);
and U7728 (N_7728,N_7439,N_7300);
nand U7729 (N_7729,N_7466,N_7437);
nand U7730 (N_7730,N_7353,N_7301);
nor U7731 (N_7731,N_7499,N_7482);
xor U7732 (N_7732,N_7327,N_7487);
and U7733 (N_7733,N_7428,N_7466);
or U7734 (N_7734,N_7439,N_7317);
xor U7735 (N_7735,N_7441,N_7495);
nand U7736 (N_7736,N_7369,N_7388);
xnor U7737 (N_7737,N_7494,N_7480);
and U7738 (N_7738,N_7410,N_7273);
nor U7739 (N_7739,N_7493,N_7401);
xor U7740 (N_7740,N_7375,N_7347);
nor U7741 (N_7741,N_7312,N_7483);
nor U7742 (N_7742,N_7315,N_7371);
or U7743 (N_7743,N_7293,N_7465);
or U7744 (N_7744,N_7323,N_7332);
nor U7745 (N_7745,N_7392,N_7324);
nor U7746 (N_7746,N_7372,N_7431);
nand U7747 (N_7747,N_7458,N_7460);
xnor U7748 (N_7748,N_7258,N_7438);
or U7749 (N_7749,N_7362,N_7497);
xnor U7750 (N_7750,N_7638,N_7533);
and U7751 (N_7751,N_7613,N_7718);
nor U7752 (N_7752,N_7676,N_7553);
nand U7753 (N_7753,N_7635,N_7597);
or U7754 (N_7754,N_7584,N_7701);
nor U7755 (N_7755,N_7504,N_7721);
nand U7756 (N_7756,N_7747,N_7535);
nor U7757 (N_7757,N_7651,N_7711);
nor U7758 (N_7758,N_7539,N_7598);
nor U7759 (N_7759,N_7709,N_7585);
or U7760 (N_7760,N_7746,N_7736);
and U7761 (N_7761,N_7632,N_7700);
nand U7762 (N_7762,N_7579,N_7655);
or U7763 (N_7763,N_7660,N_7593);
or U7764 (N_7764,N_7591,N_7714);
nor U7765 (N_7765,N_7633,N_7541);
nor U7766 (N_7766,N_7551,N_7626);
xnor U7767 (N_7767,N_7636,N_7732);
nand U7768 (N_7768,N_7534,N_7554);
or U7769 (N_7769,N_7546,N_7657);
nand U7770 (N_7770,N_7666,N_7694);
nand U7771 (N_7771,N_7616,N_7637);
and U7772 (N_7772,N_7744,N_7727);
nand U7773 (N_7773,N_7612,N_7552);
nand U7774 (N_7774,N_7501,N_7658);
or U7775 (N_7775,N_7702,N_7587);
and U7776 (N_7776,N_7514,N_7506);
nor U7777 (N_7777,N_7531,N_7712);
xnor U7778 (N_7778,N_7603,N_7532);
nand U7779 (N_7779,N_7588,N_7629);
or U7780 (N_7780,N_7627,N_7680);
xor U7781 (N_7781,N_7722,N_7735);
nand U7782 (N_7782,N_7621,N_7606);
and U7783 (N_7783,N_7601,N_7716);
and U7784 (N_7784,N_7536,N_7577);
and U7785 (N_7785,N_7668,N_7520);
xnor U7786 (N_7786,N_7557,N_7684);
or U7787 (N_7787,N_7590,N_7681);
nor U7788 (N_7788,N_7625,N_7699);
and U7789 (N_7789,N_7548,N_7595);
xnor U7790 (N_7790,N_7731,N_7592);
nor U7791 (N_7791,N_7697,N_7726);
xor U7792 (N_7792,N_7653,N_7743);
xor U7793 (N_7793,N_7679,N_7696);
xor U7794 (N_7794,N_7540,N_7599);
xnor U7795 (N_7795,N_7510,N_7537);
nand U7796 (N_7796,N_7516,N_7693);
nor U7797 (N_7797,N_7511,N_7508);
and U7798 (N_7798,N_7729,N_7605);
or U7799 (N_7799,N_7708,N_7628);
nor U7800 (N_7800,N_7558,N_7687);
xor U7801 (N_7801,N_7609,N_7674);
nor U7802 (N_7802,N_7705,N_7733);
nand U7803 (N_7803,N_7604,N_7602);
or U7804 (N_7804,N_7656,N_7622);
and U7805 (N_7805,N_7518,N_7525);
xor U7806 (N_7806,N_7503,N_7647);
xnor U7807 (N_7807,N_7739,N_7617);
and U7808 (N_7808,N_7569,N_7582);
nor U7809 (N_7809,N_7563,N_7688);
nand U7810 (N_7810,N_7523,N_7574);
or U7811 (N_7811,N_7704,N_7543);
nand U7812 (N_7812,N_7549,N_7691);
nand U7813 (N_7813,N_7581,N_7724);
nand U7814 (N_7814,N_7538,N_7567);
xnor U7815 (N_7815,N_7524,N_7659);
nand U7816 (N_7816,N_7576,N_7663);
and U7817 (N_7817,N_7644,N_7630);
or U7818 (N_7818,N_7517,N_7678);
nand U7819 (N_7819,N_7620,N_7556);
or U7820 (N_7820,N_7641,N_7689);
nor U7821 (N_7821,N_7619,N_7528);
or U7822 (N_7822,N_7573,N_7741);
nor U7823 (N_7823,N_7728,N_7745);
nand U7824 (N_7824,N_7615,N_7667);
or U7825 (N_7825,N_7652,N_7719);
and U7826 (N_7826,N_7564,N_7645);
nand U7827 (N_7827,N_7748,N_7500);
nand U7828 (N_7828,N_7634,N_7522);
xnor U7829 (N_7829,N_7515,N_7740);
xnor U7830 (N_7830,N_7509,N_7530);
and U7831 (N_7831,N_7671,N_7550);
nand U7832 (N_7832,N_7742,N_7566);
nand U7833 (N_7833,N_7692,N_7570);
xnor U7834 (N_7834,N_7571,N_7648);
and U7835 (N_7835,N_7730,N_7565);
or U7836 (N_7836,N_7586,N_7545);
nand U7837 (N_7837,N_7502,N_7650);
nor U7838 (N_7838,N_7572,N_7610);
nand U7839 (N_7839,N_7738,N_7686);
xnor U7840 (N_7840,N_7560,N_7725);
xor U7841 (N_7841,N_7513,N_7600);
nor U7842 (N_7842,N_7618,N_7527);
and U7843 (N_7843,N_7646,N_7594);
nor U7844 (N_7844,N_7575,N_7555);
nand U7845 (N_7845,N_7639,N_7521);
xor U7846 (N_7846,N_7685,N_7683);
nor U7847 (N_7847,N_7580,N_7649);
or U7848 (N_7848,N_7710,N_7717);
nand U7849 (N_7849,N_7672,N_7690);
nor U7850 (N_7850,N_7529,N_7661);
xnor U7851 (N_7851,N_7578,N_7670);
xor U7852 (N_7852,N_7707,N_7568);
nor U7853 (N_7853,N_7607,N_7631);
nor U7854 (N_7854,N_7669,N_7675);
nand U7855 (N_7855,N_7589,N_7673);
nor U7856 (N_7856,N_7596,N_7544);
nor U7857 (N_7857,N_7706,N_7715);
xor U7858 (N_7858,N_7664,N_7695);
nor U7859 (N_7859,N_7662,N_7723);
or U7860 (N_7860,N_7614,N_7640);
nor U7861 (N_7861,N_7624,N_7559);
nor U7862 (N_7862,N_7562,N_7505);
nand U7863 (N_7863,N_7611,N_7642);
nand U7864 (N_7864,N_7713,N_7583);
nand U7865 (N_7865,N_7519,N_7749);
and U7866 (N_7866,N_7561,N_7682);
and U7867 (N_7867,N_7507,N_7698);
nand U7868 (N_7868,N_7720,N_7526);
xnor U7869 (N_7869,N_7734,N_7703);
xor U7870 (N_7870,N_7643,N_7654);
nor U7871 (N_7871,N_7512,N_7665);
nor U7872 (N_7872,N_7737,N_7547);
nand U7873 (N_7873,N_7677,N_7623);
and U7874 (N_7874,N_7542,N_7608);
nand U7875 (N_7875,N_7646,N_7668);
and U7876 (N_7876,N_7568,N_7698);
and U7877 (N_7877,N_7517,N_7745);
xnor U7878 (N_7878,N_7716,N_7653);
xnor U7879 (N_7879,N_7628,N_7745);
and U7880 (N_7880,N_7542,N_7687);
nand U7881 (N_7881,N_7548,N_7618);
nor U7882 (N_7882,N_7726,N_7576);
xor U7883 (N_7883,N_7576,N_7550);
nor U7884 (N_7884,N_7614,N_7576);
nand U7885 (N_7885,N_7547,N_7735);
nor U7886 (N_7886,N_7580,N_7632);
nand U7887 (N_7887,N_7604,N_7661);
or U7888 (N_7888,N_7652,N_7518);
nand U7889 (N_7889,N_7675,N_7569);
nor U7890 (N_7890,N_7686,N_7708);
xnor U7891 (N_7891,N_7540,N_7695);
nand U7892 (N_7892,N_7520,N_7504);
nor U7893 (N_7893,N_7707,N_7689);
or U7894 (N_7894,N_7606,N_7723);
nor U7895 (N_7895,N_7743,N_7587);
and U7896 (N_7896,N_7609,N_7691);
or U7897 (N_7897,N_7631,N_7719);
nor U7898 (N_7898,N_7632,N_7523);
xnor U7899 (N_7899,N_7526,N_7648);
xnor U7900 (N_7900,N_7647,N_7717);
nor U7901 (N_7901,N_7510,N_7656);
or U7902 (N_7902,N_7687,N_7535);
nor U7903 (N_7903,N_7599,N_7704);
xor U7904 (N_7904,N_7650,N_7580);
or U7905 (N_7905,N_7705,N_7702);
xor U7906 (N_7906,N_7617,N_7630);
or U7907 (N_7907,N_7592,N_7554);
nor U7908 (N_7908,N_7523,N_7708);
nor U7909 (N_7909,N_7642,N_7616);
or U7910 (N_7910,N_7598,N_7707);
nor U7911 (N_7911,N_7745,N_7674);
nor U7912 (N_7912,N_7722,N_7729);
and U7913 (N_7913,N_7749,N_7618);
nand U7914 (N_7914,N_7597,N_7577);
and U7915 (N_7915,N_7632,N_7607);
nor U7916 (N_7916,N_7541,N_7601);
nor U7917 (N_7917,N_7599,N_7725);
nor U7918 (N_7918,N_7639,N_7534);
and U7919 (N_7919,N_7622,N_7563);
nor U7920 (N_7920,N_7547,N_7585);
and U7921 (N_7921,N_7509,N_7729);
and U7922 (N_7922,N_7695,N_7563);
nand U7923 (N_7923,N_7554,N_7693);
xnor U7924 (N_7924,N_7594,N_7650);
or U7925 (N_7925,N_7602,N_7591);
and U7926 (N_7926,N_7743,N_7504);
nor U7927 (N_7927,N_7643,N_7739);
and U7928 (N_7928,N_7560,N_7645);
or U7929 (N_7929,N_7702,N_7653);
or U7930 (N_7930,N_7526,N_7612);
and U7931 (N_7931,N_7744,N_7657);
xor U7932 (N_7932,N_7547,N_7722);
or U7933 (N_7933,N_7586,N_7511);
or U7934 (N_7934,N_7583,N_7564);
and U7935 (N_7935,N_7621,N_7626);
nor U7936 (N_7936,N_7569,N_7706);
and U7937 (N_7937,N_7646,N_7569);
and U7938 (N_7938,N_7606,N_7706);
xor U7939 (N_7939,N_7662,N_7572);
nor U7940 (N_7940,N_7529,N_7511);
xor U7941 (N_7941,N_7501,N_7747);
xnor U7942 (N_7942,N_7525,N_7572);
xnor U7943 (N_7943,N_7746,N_7611);
xor U7944 (N_7944,N_7729,N_7655);
xnor U7945 (N_7945,N_7643,N_7648);
and U7946 (N_7946,N_7529,N_7705);
and U7947 (N_7947,N_7574,N_7693);
nor U7948 (N_7948,N_7500,N_7530);
or U7949 (N_7949,N_7580,N_7525);
or U7950 (N_7950,N_7582,N_7531);
and U7951 (N_7951,N_7744,N_7729);
and U7952 (N_7952,N_7521,N_7735);
nand U7953 (N_7953,N_7727,N_7519);
nand U7954 (N_7954,N_7637,N_7519);
xnor U7955 (N_7955,N_7591,N_7511);
xor U7956 (N_7956,N_7589,N_7555);
and U7957 (N_7957,N_7624,N_7700);
nor U7958 (N_7958,N_7732,N_7517);
nor U7959 (N_7959,N_7682,N_7664);
nor U7960 (N_7960,N_7738,N_7708);
xnor U7961 (N_7961,N_7645,N_7736);
nor U7962 (N_7962,N_7629,N_7687);
nand U7963 (N_7963,N_7582,N_7657);
nand U7964 (N_7964,N_7551,N_7615);
or U7965 (N_7965,N_7727,N_7518);
nor U7966 (N_7966,N_7514,N_7745);
or U7967 (N_7967,N_7524,N_7720);
nand U7968 (N_7968,N_7505,N_7682);
or U7969 (N_7969,N_7709,N_7538);
nand U7970 (N_7970,N_7593,N_7510);
nor U7971 (N_7971,N_7712,N_7580);
and U7972 (N_7972,N_7646,N_7639);
nor U7973 (N_7973,N_7548,N_7537);
nor U7974 (N_7974,N_7574,N_7617);
nand U7975 (N_7975,N_7720,N_7717);
nand U7976 (N_7976,N_7740,N_7679);
nor U7977 (N_7977,N_7683,N_7718);
xnor U7978 (N_7978,N_7618,N_7535);
or U7979 (N_7979,N_7579,N_7607);
and U7980 (N_7980,N_7708,N_7694);
and U7981 (N_7981,N_7563,N_7522);
or U7982 (N_7982,N_7538,N_7613);
nand U7983 (N_7983,N_7725,N_7516);
and U7984 (N_7984,N_7513,N_7612);
xnor U7985 (N_7985,N_7683,N_7529);
or U7986 (N_7986,N_7674,N_7645);
or U7987 (N_7987,N_7510,N_7613);
nand U7988 (N_7988,N_7638,N_7538);
and U7989 (N_7989,N_7536,N_7743);
nand U7990 (N_7990,N_7612,N_7641);
and U7991 (N_7991,N_7637,N_7615);
nand U7992 (N_7992,N_7559,N_7744);
or U7993 (N_7993,N_7697,N_7578);
nor U7994 (N_7994,N_7630,N_7651);
and U7995 (N_7995,N_7713,N_7635);
xnor U7996 (N_7996,N_7631,N_7727);
nand U7997 (N_7997,N_7744,N_7520);
xnor U7998 (N_7998,N_7528,N_7612);
and U7999 (N_7999,N_7742,N_7733);
xor U8000 (N_8000,N_7851,N_7952);
xor U8001 (N_8001,N_7804,N_7847);
and U8002 (N_8002,N_7778,N_7763);
or U8003 (N_8003,N_7974,N_7793);
nor U8004 (N_8004,N_7877,N_7927);
or U8005 (N_8005,N_7968,N_7826);
nor U8006 (N_8006,N_7883,N_7770);
xnor U8007 (N_8007,N_7830,N_7775);
nand U8008 (N_8008,N_7939,N_7756);
nand U8009 (N_8009,N_7882,N_7798);
nand U8010 (N_8010,N_7786,N_7859);
nand U8011 (N_8011,N_7785,N_7755);
nand U8012 (N_8012,N_7867,N_7840);
nor U8013 (N_8013,N_7979,N_7792);
or U8014 (N_8014,N_7779,N_7984);
xnor U8015 (N_8015,N_7889,N_7905);
or U8016 (N_8016,N_7753,N_7926);
xnor U8017 (N_8017,N_7897,N_7922);
and U8018 (N_8018,N_7794,N_7864);
nor U8019 (N_8019,N_7961,N_7946);
xnor U8020 (N_8020,N_7967,N_7869);
nor U8021 (N_8021,N_7916,N_7872);
nor U8022 (N_8022,N_7957,N_7815);
and U8023 (N_8023,N_7782,N_7964);
and U8024 (N_8024,N_7781,N_7904);
nor U8025 (N_8025,N_7949,N_7780);
nor U8026 (N_8026,N_7959,N_7998);
and U8027 (N_8027,N_7978,N_7820);
nand U8028 (N_8028,N_7837,N_7956);
nor U8029 (N_8029,N_7773,N_7777);
nor U8030 (N_8030,N_7907,N_7963);
or U8031 (N_8031,N_7816,N_7824);
xor U8032 (N_8032,N_7865,N_7947);
and U8033 (N_8033,N_7765,N_7923);
xor U8034 (N_8034,N_7898,N_7845);
xor U8035 (N_8035,N_7918,N_7873);
xor U8036 (N_8036,N_7945,N_7915);
and U8037 (N_8037,N_7914,N_7893);
and U8038 (N_8038,N_7989,N_7831);
xor U8039 (N_8039,N_7971,N_7752);
and U8040 (N_8040,N_7875,N_7902);
nor U8041 (N_8041,N_7791,N_7784);
xnor U8042 (N_8042,N_7832,N_7996);
xnor U8043 (N_8043,N_7834,N_7774);
or U8044 (N_8044,N_7888,N_7757);
nor U8045 (N_8045,N_7841,N_7936);
xor U8046 (N_8046,N_7992,N_7766);
and U8047 (N_8047,N_7890,N_7908);
nand U8048 (N_8048,N_7800,N_7894);
nand U8049 (N_8049,N_7919,N_7938);
nor U8050 (N_8050,N_7940,N_7860);
or U8051 (N_8051,N_7958,N_7822);
xor U8052 (N_8052,N_7876,N_7990);
or U8053 (N_8053,N_7892,N_7970);
xnor U8054 (N_8054,N_7814,N_7983);
xnor U8055 (N_8055,N_7828,N_7879);
xor U8056 (N_8056,N_7950,N_7895);
nand U8057 (N_8057,N_7966,N_7759);
xor U8058 (N_8058,N_7891,N_7995);
and U8059 (N_8059,N_7975,N_7795);
nand U8060 (N_8060,N_7987,N_7913);
or U8061 (N_8061,N_7910,N_7776);
or U8062 (N_8062,N_7825,N_7829);
or U8063 (N_8063,N_7976,N_7761);
and U8064 (N_8064,N_7769,N_7880);
nor U8065 (N_8065,N_7930,N_7808);
nand U8066 (N_8066,N_7994,N_7868);
or U8067 (N_8067,N_7886,N_7805);
xnor U8068 (N_8068,N_7874,N_7972);
or U8069 (N_8069,N_7917,N_7861);
nor U8070 (N_8070,N_7758,N_7821);
nand U8071 (N_8071,N_7819,N_7884);
nor U8072 (N_8072,N_7912,N_7948);
nand U8073 (N_8073,N_7899,N_7823);
and U8074 (N_8074,N_7863,N_7817);
or U8075 (N_8075,N_7955,N_7772);
or U8076 (N_8076,N_7937,N_7981);
nand U8077 (N_8077,N_7812,N_7962);
and U8078 (N_8078,N_7943,N_7754);
or U8079 (N_8079,N_7929,N_7856);
or U8080 (N_8080,N_7935,N_7790);
nand U8081 (N_8081,N_7909,N_7811);
nor U8082 (N_8082,N_7928,N_7799);
nor U8083 (N_8083,N_7827,N_7846);
or U8084 (N_8084,N_7911,N_7944);
xor U8085 (N_8085,N_7767,N_7999);
xnor U8086 (N_8086,N_7988,N_7751);
nor U8087 (N_8087,N_7762,N_7810);
nand U8088 (N_8088,N_7787,N_7973);
xnor U8089 (N_8089,N_7942,N_7818);
xor U8090 (N_8090,N_7760,N_7803);
and U8091 (N_8091,N_7997,N_7842);
and U8092 (N_8092,N_7980,N_7796);
and U8093 (N_8093,N_7849,N_7858);
nor U8094 (N_8094,N_7878,N_7960);
and U8095 (N_8095,N_7813,N_7982);
nand U8096 (N_8096,N_7857,N_7887);
nand U8097 (N_8097,N_7932,N_7783);
and U8098 (N_8098,N_7921,N_7870);
nand U8099 (N_8099,N_7809,N_7866);
or U8100 (N_8100,N_7969,N_7941);
and U8101 (N_8101,N_7885,N_7768);
and U8102 (N_8102,N_7771,N_7896);
or U8103 (N_8103,N_7991,N_7931);
and U8104 (N_8104,N_7850,N_7797);
or U8105 (N_8105,N_7854,N_7953);
xnor U8106 (N_8106,N_7848,N_7901);
xnor U8107 (N_8107,N_7789,N_7855);
nand U8108 (N_8108,N_7871,N_7788);
and U8109 (N_8109,N_7920,N_7965);
xor U8110 (N_8110,N_7934,N_7906);
xnor U8111 (N_8111,N_7985,N_7750);
nand U8112 (N_8112,N_7900,N_7801);
xnor U8113 (N_8113,N_7838,N_7951);
and U8114 (N_8114,N_7993,N_7844);
nand U8115 (N_8115,N_7862,N_7924);
nand U8116 (N_8116,N_7933,N_7853);
and U8117 (N_8117,N_7807,N_7833);
nand U8118 (N_8118,N_7835,N_7925);
nand U8119 (N_8119,N_7954,N_7903);
xor U8120 (N_8120,N_7839,N_7836);
nor U8121 (N_8121,N_7802,N_7977);
xnor U8122 (N_8122,N_7806,N_7852);
or U8123 (N_8123,N_7881,N_7843);
and U8124 (N_8124,N_7986,N_7764);
or U8125 (N_8125,N_7783,N_7890);
xnor U8126 (N_8126,N_7937,N_7793);
nand U8127 (N_8127,N_7851,N_7861);
or U8128 (N_8128,N_7874,N_7939);
nand U8129 (N_8129,N_7932,N_7995);
and U8130 (N_8130,N_7797,N_7835);
nand U8131 (N_8131,N_7995,N_7838);
or U8132 (N_8132,N_7845,N_7906);
nand U8133 (N_8133,N_7936,N_7943);
nand U8134 (N_8134,N_7988,N_7952);
or U8135 (N_8135,N_7938,N_7901);
or U8136 (N_8136,N_7974,N_7932);
and U8137 (N_8137,N_7890,N_7766);
nand U8138 (N_8138,N_7930,N_7827);
and U8139 (N_8139,N_7940,N_7776);
xnor U8140 (N_8140,N_7807,N_7929);
nor U8141 (N_8141,N_7755,N_7758);
or U8142 (N_8142,N_7872,N_7899);
nor U8143 (N_8143,N_7847,N_7868);
nand U8144 (N_8144,N_7875,N_7837);
and U8145 (N_8145,N_7764,N_7804);
and U8146 (N_8146,N_7937,N_7883);
nor U8147 (N_8147,N_7804,N_7759);
and U8148 (N_8148,N_7980,N_7849);
and U8149 (N_8149,N_7878,N_7879);
nor U8150 (N_8150,N_7970,N_7948);
nand U8151 (N_8151,N_7898,N_7763);
or U8152 (N_8152,N_7915,N_7902);
and U8153 (N_8153,N_7768,N_7823);
and U8154 (N_8154,N_7822,N_7753);
or U8155 (N_8155,N_7803,N_7960);
xor U8156 (N_8156,N_7845,N_7985);
xor U8157 (N_8157,N_7975,N_7803);
nand U8158 (N_8158,N_7970,N_7985);
and U8159 (N_8159,N_7973,N_7946);
xor U8160 (N_8160,N_7807,N_7915);
xor U8161 (N_8161,N_7916,N_7869);
xor U8162 (N_8162,N_7846,N_7792);
nand U8163 (N_8163,N_7962,N_7887);
nor U8164 (N_8164,N_7939,N_7788);
or U8165 (N_8165,N_7939,N_7975);
nand U8166 (N_8166,N_7818,N_7992);
xnor U8167 (N_8167,N_7964,N_7899);
nor U8168 (N_8168,N_7969,N_7981);
nor U8169 (N_8169,N_7776,N_7927);
nor U8170 (N_8170,N_7970,N_7865);
and U8171 (N_8171,N_7900,N_7771);
xor U8172 (N_8172,N_7753,N_7834);
and U8173 (N_8173,N_7818,N_7877);
nand U8174 (N_8174,N_7966,N_7935);
nand U8175 (N_8175,N_7904,N_7851);
nor U8176 (N_8176,N_7775,N_7897);
nand U8177 (N_8177,N_7872,N_7935);
nor U8178 (N_8178,N_7993,N_7946);
xnor U8179 (N_8179,N_7862,N_7781);
nand U8180 (N_8180,N_7995,N_7883);
and U8181 (N_8181,N_7921,N_7883);
nor U8182 (N_8182,N_7885,N_7918);
and U8183 (N_8183,N_7968,N_7993);
nor U8184 (N_8184,N_7975,N_7908);
nand U8185 (N_8185,N_7885,N_7800);
nand U8186 (N_8186,N_7983,N_7862);
and U8187 (N_8187,N_7894,N_7902);
nor U8188 (N_8188,N_7856,N_7832);
xnor U8189 (N_8189,N_7806,N_7818);
and U8190 (N_8190,N_7875,N_7895);
and U8191 (N_8191,N_7841,N_7764);
nor U8192 (N_8192,N_7788,N_7867);
nor U8193 (N_8193,N_7792,N_7889);
xnor U8194 (N_8194,N_7969,N_7937);
and U8195 (N_8195,N_7825,N_7862);
nor U8196 (N_8196,N_7973,N_7892);
or U8197 (N_8197,N_7997,N_7825);
or U8198 (N_8198,N_7817,N_7766);
nor U8199 (N_8199,N_7849,N_7927);
and U8200 (N_8200,N_7901,N_7784);
xor U8201 (N_8201,N_7948,N_7787);
nand U8202 (N_8202,N_7861,N_7787);
nor U8203 (N_8203,N_7930,N_7954);
or U8204 (N_8204,N_7819,N_7768);
xor U8205 (N_8205,N_7966,N_7889);
xor U8206 (N_8206,N_7953,N_7808);
nand U8207 (N_8207,N_7931,N_7861);
or U8208 (N_8208,N_7788,N_7994);
nand U8209 (N_8209,N_7994,N_7992);
nor U8210 (N_8210,N_7757,N_7850);
xor U8211 (N_8211,N_7997,N_7900);
or U8212 (N_8212,N_7777,N_7962);
or U8213 (N_8213,N_7813,N_7852);
nand U8214 (N_8214,N_7890,N_7913);
and U8215 (N_8215,N_7881,N_7909);
nand U8216 (N_8216,N_7850,N_7760);
xor U8217 (N_8217,N_7769,N_7767);
xor U8218 (N_8218,N_7868,N_7875);
xnor U8219 (N_8219,N_7973,N_7886);
or U8220 (N_8220,N_7837,N_7809);
or U8221 (N_8221,N_7844,N_7842);
and U8222 (N_8222,N_7982,N_7832);
nor U8223 (N_8223,N_7857,N_7862);
and U8224 (N_8224,N_7945,N_7872);
nor U8225 (N_8225,N_7980,N_7817);
and U8226 (N_8226,N_7957,N_7772);
or U8227 (N_8227,N_7948,N_7837);
xnor U8228 (N_8228,N_7838,N_7762);
xnor U8229 (N_8229,N_7785,N_7879);
nor U8230 (N_8230,N_7759,N_7783);
nor U8231 (N_8231,N_7946,N_7916);
xnor U8232 (N_8232,N_7831,N_7813);
and U8233 (N_8233,N_7899,N_7980);
or U8234 (N_8234,N_7896,N_7792);
nand U8235 (N_8235,N_7870,N_7842);
and U8236 (N_8236,N_7980,N_7913);
nand U8237 (N_8237,N_7834,N_7943);
xnor U8238 (N_8238,N_7921,N_7826);
or U8239 (N_8239,N_7791,N_7783);
nor U8240 (N_8240,N_7799,N_7877);
or U8241 (N_8241,N_7943,N_7877);
or U8242 (N_8242,N_7797,N_7928);
nand U8243 (N_8243,N_7786,N_7909);
xor U8244 (N_8244,N_7891,N_7875);
nand U8245 (N_8245,N_7877,N_7803);
and U8246 (N_8246,N_7825,N_7981);
and U8247 (N_8247,N_7984,N_7750);
nand U8248 (N_8248,N_7785,N_7967);
nor U8249 (N_8249,N_7902,N_7886);
and U8250 (N_8250,N_8012,N_8190);
nand U8251 (N_8251,N_8235,N_8127);
nor U8252 (N_8252,N_8003,N_8051);
and U8253 (N_8253,N_8214,N_8196);
nand U8254 (N_8254,N_8061,N_8107);
and U8255 (N_8255,N_8189,N_8146);
or U8256 (N_8256,N_8105,N_8208);
or U8257 (N_8257,N_8064,N_8075);
or U8258 (N_8258,N_8038,N_8004);
xor U8259 (N_8259,N_8162,N_8147);
xnor U8260 (N_8260,N_8066,N_8156);
xnor U8261 (N_8261,N_8157,N_8117);
and U8262 (N_8262,N_8216,N_8089);
nor U8263 (N_8263,N_8129,N_8231);
nand U8264 (N_8264,N_8095,N_8171);
or U8265 (N_8265,N_8232,N_8215);
or U8266 (N_8266,N_8132,N_8010);
nor U8267 (N_8267,N_8062,N_8233);
nand U8268 (N_8268,N_8096,N_8000);
nand U8269 (N_8269,N_8060,N_8218);
nand U8270 (N_8270,N_8238,N_8194);
nor U8271 (N_8271,N_8230,N_8073);
nor U8272 (N_8272,N_8185,N_8212);
nand U8273 (N_8273,N_8183,N_8085);
nand U8274 (N_8274,N_8043,N_8136);
and U8275 (N_8275,N_8020,N_8009);
nor U8276 (N_8276,N_8120,N_8111);
or U8277 (N_8277,N_8188,N_8153);
or U8278 (N_8278,N_8041,N_8145);
nor U8279 (N_8279,N_8101,N_8023);
and U8280 (N_8280,N_8213,N_8143);
xor U8281 (N_8281,N_8170,N_8006);
nand U8282 (N_8282,N_8080,N_8174);
or U8283 (N_8283,N_8052,N_8133);
nand U8284 (N_8284,N_8217,N_8246);
or U8285 (N_8285,N_8021,N_8122);
xnor U8286 (N_8286,N_8109,N_8092);
nor U8287 (N_8287,N_8173,N_8017);
xnor U8288 (N_8288,N_8197,N_8205);
xnor U8289 (N_8289,N_8131,N_8224);
xor U8290 (N_8290,N_8158,N_8201);
xor U8291 (N_8291,N_8001,N_8028);
nand U8292 (N_8292,N_8037,N_8248);
xnor U8293 (N_8293,N_8079,N_8019);
nand U8294 (N_8294,N_8099,N_8139);
nor U8295 (N_8295,N_8053,N_8240);
or U8296 (N_8296,N_8242,N_8039);
nand U8297 (N_8297,N_8106,N_8222);
nor U8298 (N_8298,N_8195,N_8055);
or U8299 (N_8299,N_8093,N_8211);
and U8300 (N_8300,N_8169,N_8124);
nor U8301 (N_8301,N_8031,N_8049);
nand U8302 (N_8302,N_8236,N_8126);
xnor U8303 (N_8303,N_8227,N_8088);
nor U8304 (N_8304,N_8084,N_8177);
nor U8305 (N_8305,N_8022,N_8065);
and U8306 (N_8306,N_8209,N_8058);
xor U8307 (N_8307,N_8172,N_8229);
xnor U8308 (N_8308,N_8239,N_8203);
xnor U8309 (N_8309,N_8057,N_8181);
and U8310 (N_8310,N_8042,N_8030);
nor U8311 (N_8311,N_8115,N_8016);
or U8312 (N_8312,N_8159,N_8138);
and U8313 (N_8313,N_8108,N_8144);
nand U8314 (N_8314,N_8182,N_8068);
xnor U8315 (N_8315,N_8245,N_8063);
and U8316 (N_8316,N_8036,N_8048);
nor U8317 (N_8317,N_8164,N_8098);
nand U8318 (N_8318,N_8210,N_8083);
xor U8319 (N_8319,N_8008,N_8160);
or U8320 (N_8320,N_8130,N_8114);
and U8321 (N_8321,N_8087,N_8168);
nand U8322 (N_8322,N_8237,N_8040);
xor U8323 (N_8323,N_8027,N_8046);
xnor U8324 (N_8324,N_8135,N_8125);
and U8325 (N_8325,N_8202,N_8178);
and U8326 (N_8326,N_8033,N_8206);
xnor U8327 (N_8327,N_8152,N_8082);
nand U8328 (N_8328,N_8176,N_8112);
xnor U8329 (N_8329,N_8163,N_8167);
and U8330 (N_8330,N_8166,N_8024);
and U8331 (N_8331,N_8094,N_8047);
nor U8332 (N_8332,N_8045,N_8228);
and U8333 (N_8333,N_8220,N_8113);
nor U8334 (N_8334,N_8015,N_8186);
nand U8335 (N_8335,N_8011,N_8226);
nor U8336 (N_8336,N_8140,N_8118);
nand U8337 (N_8337,N_8002,N_8070);
and U8338 (N_8338,N_8007,N_8154);
nor U8339 (N_8339,N_8128,N_8241);
nor U8340 (N_8340,N_8249,N_8149);
or U8341 (N_8341,N_8104,N_8221);
nand U8342 (N_8342,N_8076,N_8155);
xor U8343 (N_8343,N_8134,N_8072);
nor U8344 (N_8344,N_8223,N_8077);
nand U8345 (N_8345,N_8110,N_8148);
or U8346 (N_8346,N_8086,N_8198);
and U8347 (N_8347,N_8067,N_8059);
nand U8348 (N_8348,N_8165,N_8029);
and U8349 (N_8349,N_8161,N_8018);
nand U8350 (N_8350,N_8244,N_8179);
xor U8351 (N_8351,N_8100,N_8150);
nand U8352 (N_8352,N_8151,N_8026);
and U8353 (N_8353,N_8069,N_8142);
xor U8354 (N_8354,N_8141,N_8123);
and U8355 (N_8355,N_8014,N_8056);
or U8356 (N_8356,N_8034,N_8137);
nand U8357 (N_8357,N_8243,N_8081);
nand U8358 (N_8358,N_8219,N_8119);
xnor U8359 (N_8359,N_8116,N_8193);
or U8360 (N_8360,N_8184,N_8054);
nor U8361 (N_8361,N_8225,N_8071);
and U8362 (N_8362,N_8121,N_8025);
or U8363 (N_8363,N_8199,N_8175);
or U8364 (N_8364,N_8097,N_8078);
xnor U8365 (N_8365,N_8180,N_8191);
and U8366 (N_8366,N_8044,N_8032);
xor U8367 (N_8367,N_8090,N_8013);
or U8368 (N_8368,N_8091,N_8005);
xor U8369 (N_8369,N_8247,N_8207);
nor U8370 (N_8370,N_8234,N_8200);
nand U8371 (N_8371,N_8192,N_8103);
nand U8372 (N_8372,N_8187,N_8204);
and U8373 (N_8373,N_8102,N_8050);
nor U8374 (N_8374,N_8035,N_8074);
and U8375 (N_8375,N_8162,N_8049);
xnor U8376 (N_8376,N_8185,N_8062);
nand U8377 (N_8377,N_8229,N_8225);
nand U8378 (N_8378,N_8208,N_8159);
or U8379 (N_8379,N_8067,N_8245);
nor U8380 (N_8380,N_8184,N_8221);
nand U8381 (N_8381,N_8103,N_8070);
nand U8382 (N_8382,N_8195,N_8154);
xor U8383 (N_8383,N_8121,N_8230);
and U8384 (N_8384,N_8021,N_8135);
and U8385 (N_8385,N_8117,N_8070);
nand U8386 (N_8386,N_8233,N_8074);
xor U8387 (N_8387,N_8091,N_8103);
or U8388 (N_8388,N_8059,N_8033);
or U8389 (N_8389,N_8127,N_8220);
nor U8390 (N_8390,N_8004,N_8123);
nor U8391 (N_8391,N_8056,N_8004);
and U8392 (N_8392,N_8034,N_8122);
nand U8393 (N_8393,N_8161,N_8189);
nor U8394 (N_8394,N_8202,N_8116);
or U8395 (N_8395,N_8048,N_8237);
xnor U8396 (N_8396,N_8089,N_8102);
and U8397 (N_8397,N_8217,N_8078);
nor U8398 (N_8398,N_8056,N_8108);
or U8399 (N_8399,N_8084,N_8131);
xor U8400 (N_8400,N_8150,N_8066);
or U8401 (N_8401,N_8209,N_8222);
xnor U8402 (N_8402,N_8227,N_8107);
or U8403 (N_8403,N_8173,N_8069);
and U8404 (N_8404,N_8072,N_8206);
nand U8405 (N_8405,N_8211,N_8151);
xnor U8406 (N_8406,N_8033,N_8144);
nor U8407 (N_8407,N_8065,N_8171);
nand U8408 (N_8408,N_8233,N_8063);
xor U8409 (N_8409,N_8011,N_8243);
and U8410 (N_8410,N_8022,N_8044);
or U8411 (N_8411,N_8056,N_8024);
or U8412 (N_8412,N_8184,N_8170);
and U8413 (N_8413,N_8213,N_8086);
and U8414 (N_8414,N_8223,N_8179);
xnor U8415 (N_8415,N_8177,N_8120);
or U8416 (N_8416,N_8231,N_8101);
nor U8417 (N_8417,N_8156,N_8171);
and U8418 (N_8418,N_8225,N_8143);
nor U8419 (N_8419,N_8139,N_8123);
nand U8420 (N_8420,N_8112,N_8017);
nor U8421 (N_8421,N_8212,N_8105);
nand U8422 (N_8422,N_8082,N_8039);
nand U8423 (N_8423,N_8004,N_8170);
or U8424 (N_8424,N_8095,N_8049);
nand U8425 (N_8425,N_8204,N_8195);
or U8426 (N_8426,N_8034,N_8101);
or U8427 (N_8427,N_8249,N_8114);
nand U8428 (N_8428,N_8022,N_8056);
and U8429 (N_8429,N_8208,N_8090);
xnor U8430 (N_8430,N_8019,N_8080);
nand U8431 (N_8431,N_8201,N_8078);
xnor U8432 (N_8432,N_8157,N_8216);
and U8433 (N_8433,N_8195,N_8164);
and U8434 (N_8434,N_8124,N_8039);
xor U8435 (N_8435,N_8084,N_8203);
nand U8436 (N_8436,N_8236,N_8133);
or U8437 (N_8437,N_8161,N_8068);
and U8438 (N_8438,N_8218,N_8223);
xnor U8439 (N_8439,N_8079,N_8045);
or U8440 (N_8440,N_8007,N_8016);
or U8441 (N_8441,N_8248,N_8012);
xor U8442 (N_8442,N_8127,N_8081);
nand U8443 (N_8443,N_8223,N_8182);
or U8444 (N_8444,N_8115,N_8104);
or U8445 (N_8445,N_8049,N_8192);
and U8446 (N_8446,N_8224,N_8173);
nand U8447 (N_8447,N_8165,N_8167);
nand U8448 (N_8448,N_8227,N_8138);
and U8449 (N_8449,N_8099,N_8032);
xnor U8450 (N_8450,N_8227,N_8019);
xnor U8451 (N_8451,N_8082,N_8228);
nor U8452 (N_8452,N_8124,N_8231);
nand U8453 (N_8453,N_8196,N_8009);
nand U8454 (N_8454,N_8051,N_8238);
nor U8455 (N_8455,N_8184,N_8039);
or U8456 (N_8456,N_8223,N_8057);
or U8457 (N_8457,N_8185,N_8121);
and U8458 (N_8458,N_8239,N_8218);
nand U8459 (N_8459,N_8158,N_8047);
nor U8460 (N_8460,N_8017,N_8066);
xor U8461 (N_8461,N_8181,N_8196);
or U8462 (N_8462,N_8182,N_8001);
nand U8463 (N_8463,N_8180,N_8197);
and U8464 (N_8464,N_8238,N_8135);
and U8465 (N_8465,N_8047,N_8106);
xor U8466 (N_8466,N_8019,N_8202);
and U8467 (N_8467,N_8204,N_8051);
xor U8468 (N_8468,N_8126,N_8152);
and U8469 (N_8469,N_8181,N_8039);
xor U8470 (N_8470,N_8149,N_8190);
or U8471 (N_8471,N_8053,N_8026);
nand U8472 (N_8472,N_8037,N_8171);
or U8473 (N_8473,N_8162,N_8114);
nor U8474 (N_8474,N_8234,N_8239);
or U8475 (N_8475,N_8134,N_8157);
nand U8476 (N_8476,N_8154,N_8051);
and U8477 (N_8477,N_8044,N_8046);
and U8478 (N_8478,N_8052,N_8164);
or U8479 (N_8479,N_8068,N_8158);
nor U8480 (N_8480,N_8193,N_8162);
or U8481 (N_8481,N_8180,N_8071);
nor U8482 (N_8482,N_8089,N_8127);
nand U8483 (N_8483,N_8246,N_8125);
nand U8484 (N_8484,N_8079,N_8240);
nand U8485 (N_8485,N_8147,N_8001);
and U8486 (N_8486,N_8243,N_8071);
and U8487 (N_8487,N_8042,N_8200);
xnor U8488 (N_8488,N_8209,N_8141);
and U8489 (N_8489,N_8131,N_8006);
nor U8490 (N_8490,N_8202,N_8209);
nor U8491 (N_8491,N_8192,N_8036);
and U8492 (N_8492,N_8081,N_8085);
and U8493 (N_8493,N_8230,N_8034);
or U8494 (N_8494,N_8171,N_8060);
or U8495 (N_8495,N_8151,N_8230);
nor U8496 (N_8496,N_8244,N_8205);
xnor U8497 (N_8497,N_8079,N_8070);
or U8498 (N_8498,N_8202,N_8181);
nor U8499 (N_8499,N_8169,N_8106);
and U8500 (N_8500,N_8483,N_8342);
and U8501 (N_8501,N_8366,N_8486);
nor U8502 (N_8502,N_8490,N_8260);
nor U8503 (N_8503,N_8421,N_8259);
or U8504 (N_8504,N_8382,N_8328);
or U8505 (N_8505,N_8286,N_8258);
xnor U8506 (N_8506,N_8378,N_8406);
or U8507 (N_8507,N_8475,N_8255);
nand U8508 (N_8508,N_8317,N_8369);
xnor U8509 (N_8509,N_8276,N_8288);
nand U8510 (N_8510,N_8468,N_8325);
or U8511 (N_8511,N_8372,N_8266);
or U8512 (N_8512,N_8389,N_8384);
nand U8513 (N_8513,N_8485,N_8474);
and U8514 (N_8514,N_8261,N_8448);
or U8515 (N_8515,N_8472,N_8411);
or U8516 (N_8516,N_8365,N_8412);
nand U8517 (N_8517,N_8469,N_8352);
or U8518 (N_8518,N_8387,N_8383);
or U8519 (N_8519,N_8481,N_8464);
and U8520 (N_8520,N_8386,N_8357);
and U8521 (N_8521,N_8432,N_8309);
nand U8522 (N_8522,N_8426,N_8457);
and U8523 (N_8523,N_8415,N_8462);
or U8524 (N_8524,N_8435,N_8418);
nand U8525 (N_8525,N_8330,N_8404);
xnor U8526 (N_8526,N_8397,N_8409);
nand U8527 (N_8527,N_8305,N_8262);
nand U8528 (N_8528,N_8381,N_8374);
and U8529 (N_8529,N_8277,N_8497);
nand U8530 (N_8530,N_8287,N_8429);
and U8531 (N_8531,N_8393,N_8430);
nor U8532 (N_8532,N_8375,N_8340);
xor U8533 (N_8533,N_8336,N_8451);
xor U8534 (N_8534,N_8252,N_8269);
and U8535 (N_8535,N_8358,N_8461);
nand U8536 (N_8536,N_8407,N_8280);
nor U8537 (N_8537,N_8494,N_8379);
and U8538 (N_8538,N_8385,N_8360);
or U8539 (N_8539,N_8282,N_8300);
or U8540 (N_8540,N_8450,N_8491);
xor U8541 (N_8541,N_8456,N_8399);
and U8542 (N_8542,N_8298,N_8291);
nor U8543 (N_8543,N_8484,N_8299);
nand U8544 (N_8544,N_8319,N_8463);
xnor U8545 (N_8545,N_8439,N_8422);
nand U8546 (N_8546,N_8416,N_8303);
nor U8547 (N_8547,N_8326,N_8334);
or U8548 (N_8548,N_8493,N_8394);
xnor U8549 (N_8549,N_8272,N_8345);
xnor U8550 (N_8550,N_8445,N_8312);
and U8551 (N_8551,N_8431,N_8293);
nand U8552 (N_8552,N_8473,N_8459);
xor U8553 (N_8553,N_8424,N_8413);
or U8554 (N_8554,N_8353,N_8438);
and U8555 (N_8555,N_8346,N_8477);
and U8556 (N_8556,N_8308,N_8414);
nor U8557 (N_8557,N_8428,N_8443);
nand U8558 (N_8558,N_8437,N_8471);
xor U8559 (N_8559,N_8344,N_8402);
and U8560 (N_8560,N_8351,N_8264);
xnor U8561 (N_8561,N_8489,N_8318);
or U8562 (N_8562,N_8274,N_8256);
nand U8563 (N_8563,N_8400,N_8480);
nor U8564 (N_8564,N_8455,N_8284);
xnor U8565 (N_8565,N_8302,N_8285);
or U8566 (N_8566,N_8337,N_8327);
xnor U8567 (N_8567,N_8495,N_8278);
xor U8568 (N_8568,N_8306,N_8408);
nor U8569 (N_8569,N_8410,N_8403);
or U8570 (N_8570,N_8359,N_8263);
xor U8571 (N_8571,N_8371,N_8447);
and U8572 (N_8572,N_8425,N_8405);
or U8573 (N_8573,N_8388,N_8310);
or U8574 (N_8574,N_8267,N_8396);
and U8575 (N_8575,N_8417,N_8279);
or U8576 (N_8576,N_8391,N_8478);
and U8577 (N_8577,N_8275,N_8301);
and U8578 (N_8578,N_8355,N_8335);
or U8579 (N_8579,N_8440,N_8283);
nand U8580 (N_8580,N_8496,N_8449);
nand U8581 (N_8581,N_8311,N_8434);
nor U8582 (N_8582,N_8356,N_8251);
nand U8583 (N_8583,N_8361,N_8488);
and U8584 (N_8584,N_8290,N_8354);
nor U8585 (N_8585,N_8362,N_8343);
and U8586 (N_8586,N_8442,N_8367);
and U8587 (N_8587,N_8304,N_8271);
or U8588 (N_8588,N_8254,N_8398);
and U8589 (N_8589,N_8467,N_8329);
nor U8590 (N_8590,N_8295,N_8313);
nor U8591 (N_8591,N_8321,N_8270);
and U8592 (N_8592,N_8401,N_8380);
nand U8593 (N_8593,N_8324,N_8420);
xor U8594 (N_8594,N_8349,N_8377);
nor U8595 (N_8595,N_8460,N_8265);
and U8596 (N_8596,N_8368,N_8294);
nor U8597 (N_8597,N_8454,N_8482);
or U8598 (N_8598,N_8350,N_8320);
nand U8599 (N_8599,N_8339,N_8296);
and U8600 (N_8600,N_8392,N_8487);
or U8601 (N_8601,N_8332,N_8470);
xnor U8602 (N_8602,N_8476,N_8273);
nand U8603 (N_8603,N_8370,N_8363);
or U8604 (N_8604,N_8373,N_8250);
xnor U8605 (N_8605,N_8314,N_8333);
or U8606 (N_8606,N_8499,N_8307);
or U8607 (N_8607,N_8419,N_8268);
or U8608 (N_8608,N_8257,N_8253);
or U8609 (N_8609,N_8465,N_8323);
or U8610 (N_8610,N_8436,N_8458);
and U8611 (N_8611,N_8395,N_8289);
or U8612 (N_8612,N_8433,N_8292);
nor U8613 (N_8613,N_8441,N_8341);
nand U8614 (N_8614,N_8331,N_8376);
or U8615 (N_8615,N_8492,N_8466);
and U8616 (N_8616,N_8452,N_8479);
nand U8617 (N_8617,N_8390,N_8498);
nand U8618 (N_8618,N_8322,N_8316);
or U8619 (N_8619,N_8427,N_8347);
nor U8620 (N_8620,N_8364,N_8444);
nand U8621 (N_8621,N_8453,N_8348);
xor U8622 (N_8622,N_8281,N_8423);
and U8623 (N_8623,N_8338,N_8315);
xor U8624 (N_8624,N_8297,N_8446);
or U8625 (N_8625,N_8352,N_8325);
or U8626 (N_8626,N_8377,N_8407);
or U8627 (N_8627,N_8426,N_8316);
and U8628 (N_8628,N_8439,N_8353);
and U8629 (N_8629,N_8387,N_8497);
xor U8630 (N_8630,N_8366,N_8345);
nor U8631 (N_8631,N_8451,N_8330);
nor U8632 (N_8632,N_8433,N_8373);
nand U8633 (N_8633,N_8305,N_8339);
or U8634 (N_8634,N_8302,N_8496);
or U8635 (N_8635,N_8354,N_8288);
nor U8636 (N_8636,N_8356,N_8295);
or U8637 (N_8637,N_8488,N_8300);
or U8638 (N_8638,N_8343,N_8443);
and U8639 (N_8639,N_8368,N_8444);
and U8640 (N_8640,N_8327,N_8411);
nand U8641 (N_8641,N_8436,N_8398);
xor U8642 (N_8642,N_8344,N_8414);
nand U8643 (N_8643,N_8301,N_8493);
and U8644 (N_8644,N_8392,N_8440);
nor U8645 (N_8645,N_8330,N_8419);
xnor U8646 (N_8646,N_8318,N_8374);
nor U8647 (N_8647,N_8377,N_8251);
or U8648 (N_8648,N_8377,N_8381);
xnor U8649 (N_8649,N_8299,N_8461);
xor U8650 (N_8650,N_8429,N_8484);
xor U8651 (N_8651,N_8272,N_8391);
nor U8652 (N_8652,N_8324,N_8489);
or U8653 (N_8653,N_8348,N_8488);
nor U8654 (N_8654,N_8305,N_8413);
nor U8655 (N_8655,N_8294,N_8349);
and U8656 (N_8656,N_8326,N_8437);
or U8657 (N_8657,N_8263,N_8310);
nor U8658 (N_8658,N_8390,N_8337);
or U8659 (N_8659,N_8496,N_8305);
nand U8660 (N_8660,N_8281,N_8331);
nand U8661 (N_8661,N_8492,N_8394);
and U8662 (N_8662,N_8377,N_8486);
nor U8663 (N_8663,N_8307,N_8367);
or U8664 (N_8664,N_8451,N_8280);
or U8665 (N_8665,N_8479,N_8424);
nand U8666 (N_8666,N_8256,N_8418);
and U8667 (N_8667,N_8299,N_8487);
and U8668 (N_8668,N_8357,N_8332);
or U8669 (N_8669,N_8474,N_8460);
nor U8670 (N_8670,N_8488,N_8443);
and U8671 (N_8671,N_8359,N_8427);
and U8672 (N_8672,N_8371,N_8412);
xor U8673 (N_8673,N_8344,N_8342);
nand U8674 (N_8674,N_8341,N_8446);
and U8675 (N_8675,N_8265,N_8279);
and U8676 (N_8676,N_8412,N_8353);
nand U8677 (N_8677,N_8330,N_8486);
xnor U8678 (N_8678,N_8455,N_8372);
nand U8679 (N_8679,N_8372,N_8368);
nand U8680 (N_8680,N_8378,N_8477);
and U8681 (N_8681,N_8384,N_8366);
nor U8682 (N_8682,N_8264,N_8287);
xnor U8683 (N_8683,N_8482,N_8396);
or U8684 (N_8684,N_8327,N_8265);
nor U8685 (N_8685,N_8381,N_8348);
nand U8686 (N_8686,N_8480,N_8298);
and U8687 (N_8687,N_8459,N_8373);
and U8688 (N_8688,N_8465,N_8380);
nor U8689 (N_8689,N_8438,N_8368);
and U8690 (N_8690,N_8349,N_8363);
or U8691 (N_8691,N_8368,N_8303);
nand U8692 (N_8692,N_8320,N_8328);
or U8693 (N_8693,N_8449,N_8402);
nand U8694 (N_8694,N_8373,N_8358);
xnor U8695 (N_8695,N_8431,N_8373);
nor U8696 (N_8696,N_8309,N_8495);
and U8697 (N_8697,N_8402,N_8454);
and U8698 (N_8698,N_8467,N_8325);
nor U8699 (N_8699,N_8463,N_8329);
nand U8700 (N_8700,N_8428,N_8324);
xnor U8701 (N_8701,N_8307,N_8445);
or U8702 (N_8702,N_8395,N_8433);
and U8703 (N_8703,N_8416,N_8410);
or U8704 (N_8704,N_8482,N_8406);
or U8705 (N_8705,N_8414,N_8280);
or U8706 (N_8706,N_8380,N_8440);
nand U8707 (N_8707,N_8445,N_8266);
and U8708 (N_8708,N_8379,N_8462);
nand U8709 (N_8709,N_8291,N_8455);
nand U8710 (N_8710,N_8428,N_8408);
and U8711 (N_8711,N_8353,N_8274);
nor U8712 (N_8712,N_8443,N_8286);
or U8713 (N_8713,N_8484,N_8356);
and U8714 (N_8714,N_8360,N_8303);
or U8715 (N_8715,N_8345,N_8271);
xor U8716 (N_8716,N_8350,N_8404);
nand U8717 (N_8717,N_8412,N_8484);
or U8718 (N_8718,N_8495,N_8376);
and U8719 (N_8719,N_8486,N_8349);
nand U8720 (N_8720,N_8452,N_8286);
and U8721 (N_8721,N_8469,N_8443);
or U8722 (N_8722,N_8440,N_8263);
nand U8723 (N_8723,N_8345,N_8453);
nor U8724 (N_8724,N_8481,N_8448);
or U8725 (N_8725,N_8386,N_8416);
or U8726 (N_8726,N_8258,N_8252);
and U8727 (N_8727,N_8488,N_8413);
and U8728 (N_8728,N_8407,N_8454);
nand U8729 (N_8729,N_8422,N_8351);
xor U8730 (N_8730,N_8483,N_8461);
nand U8731 (N_8731,N_8370,N_8459);
nor U8732 (N_8732,N_8498,N_8305);
nor U8733 (N_8733,N_8491,N_8345);
and U8734 (N_8734,N_8256,N_8400);
and U8735 (N_8735,N_8384,N_8499);
or U8736 (N_8736,N_8419,N_8288);
nor U8737 (N_8737,N_8324,N_8321);
nand U8738 (N_8738,N_8438,N_8397);
and U8739 (N_8739,N_8356,N_8448);
and U8740 (N_8740,N_8445,N_8459);
and U8741 (N_8741,N_8438,N_8428);
xor U8742 (N_8742,N_8264,N_8399);
and U8743 (N_8743,N_8433,N_8421);
nand U8744 (N_8744,N_8393,N_8310);
nor U8745 (N_8745,N_8346,N_8381);
nor U8746 (N_8746,N_8262,N_8434);
nand U8747 (N_8747,N_8455,N_8281);
xor U8748 (N_8748,N_8396,N_8466);
and U8749 (N_8749,N_8282,N_8283);
nand U8750 (N_8750,N_8535,N_8559);
nor U8751 (N_8751,N_8642,N_8521);
or U8752 (N_8752,N_8553,N_8645);
xor U8753 (N_8753,N_8622,N_8671);
nand U8754 (N_8754,N_8627,N_8504);
nor U8755 (N_8755,N_8530,N_8555);
or U8756 (N_8756,N_8603,N_8749);
xor U8757 (N_8757,N_8683,N_8575);
or U8758 (N_8758,N_8510,N_8591);
or U8759 (N_8759,N_8656,N_8515);
xor U8760 (N_8760,N_8501,N_8520);
nand U8761 (N_8761,N_8672,N_8658);
nor U8762 (N_8762,N_8602,N_8560);
xor U8763 (N_8763,N_8505,N_8735);
nor U8764 (N_8764,N_8599,N_8513);
and U8765 (N_8765,N_8579,N_8595);
nor U8766 (N_8766,N_8712,N_8736);
nand U8767 (N_8767,N_8541,N_8666);
or U8768 (N_8768,N_8648,N_8563);
or U8769 (N_8769,N_8681,N_8691);
nand U8770 (N_8770,N_8619,N_8662);
or U8771 (N_8771,N_8634,N_8734);
and U8772 (N_8772,N_8632,N_8650);
nor U8773 (N_8773,N_8682,N_8720);
xnor U8774 (N_8774,N_8611,N_8524);
or U8775 (N_8775,N_8631,N_8721);
or U8776 (N_8776,N_8582,N_8544);
and U8777 (N_8777,N_8674,N_8704);
xor U8778 (N_8778,N_8509,N_8588);
and U8779 (N_8779,N_8739,N_8637);
nor U8780 (N_8780,N_8703,N_8605);
nor U8781 (N_8781,N_8571,N_8639);
nor U8782 (N_8782,N_8557,N_8547);
or U8783 (N_8783,N_8545,N_8701);
nand U8784 (N_8784,N_8686,N_8586);
or U8785 (N_8785,N_8635,N_8731);
nor U8786 (N_8786,N_8742,N_8711);
or U8787 (N_8787,N_8673,N_8694);
or U8788 (N_8788,N_8633,N_8695);
or U8789 (N_8789,N_8710,N_8625);
nand U8790 (N_8790,N_8657,N_8733);
nand U8791 (N_8791,N_8725,N_8743);
nor U8792 (N_8792,N_8716,N_8620);
or U8793 (N_8793,N_8713,N_8518);
nor U8794 (N_8794,N_8536,N_8651);
and U8795 (N_8795,N_8675,N_8727);
nand U8796 (N_8796,N_8665,N_8718);
or U8797 (N_8797,N_8638,N_8717);
and U8798 (N_8798,N_8730,N_8511);
nor U8799 (N_8799,N_8668,N_8534);
or U8800 (N_8800,N_8653,N_8570);
or U8801 (N_8801,N_8542,N_8723);
xor U8802 (N_8802,N_8507,N_8699);
or U8803 (N_8803,N_8550,N_8726);
nor U8804 (N_8804,N_8621,N_8506);
or U8805 (N_8805,N_8549,N_8660);
and U8806 (N_8806,N_8519,N_8641);
and U8807 (N_8807,N_8587,N_8589);
and U8808 (N_8808,N_8585,N_8617);
nand U8809 (N_8809,N_8568,N_8676);
nor U8810 (N_8810,N_8667,N_8548);
or U8811 (N_8811,N_8552,N_8607);
xor U8812 (N_8812,N_8615,N_8577);
nand U8813 (N_8813,N_8689,N_8566);
nor U8814 (N_8814,N_8659,N_8567);
nand U8815 (N_8815,N_8610,N_8594);
nor U8816 (N_8816,N_8606,N_8629);
xnor U8817 (N_8817,N_8700,N_8543);
and U8818 (N_8818,N_8644,N_8612);
xnor U8819 (N_8819,N_8688,N_8598);
and U8820 (N_8820,N_8531,N_8564);
and U8821 (N_8821,N_8546,N_8687);
or U8822 (N_8822,N_8630,N_8628);
nand U8823 (N_8823,N_8540,N_8709);
or U8824 (N_8824,N_8655,N_8643);
nand U8825 (N_8825,N_8590,N_8680);
nand U8826 (N_8826,N_8514,N_8670);
xor U8827 (N_8827,N_8623,N_8702);
xnor U8828 (N_8828,N_8522,N_8604);
xor U8829 (N_8829,N_8729,N_8640);
and U8830 (N_8830,N_8705,N_8609);
nor U8831 (N_8831,N_8741,N_8693);
nor U8832 (N_8832,N_8664,N_8661);
or U8833 (N_8833,N_8618,N_8596);
nand U8834 (N_8834,N_8561,N_8647);
or U8835 (N_8835,N_8584,N_8608);
and U8836 (N_8836,N_8578,N_8685);
xor U8837 (N_8837,N_8669,N_8613);
and U8838 (N_8838,N_8745,N_8574);
and U8839 (N_8839,N_8707,N_8565);
nand U8840 (N_8840,N_8714,N_8706);
nor U8841 (N_8841,N_8500,N_8597);
or U8842 (N_8842,N_8684,N_8740);
nor U8843 (N_8843,N_8539,N_8517);
and U8844 (N_8844,N_8738,N_8747);
xnor U8845 (N_8845,N_8708,N_8724);
nand U8846 (N_8846,N_8715,N_8679);
xnor U8847 (N_8847,N_8551,N_8601);
or U8848 (N_8848,N_8508,N_8593);
nand U8849 (N_8849,N_8558,N_8538);
xnor U8850 (N_8850,N_8529,N_8646);
nor U8851 (N_8851,N_8636,N_8554);
and U8852 (N_8852,N_8624,N_8576);
xor U8853 (N_8853,N_8626,N_8732);
or U8854 (N_8854,N_8502,N_8698);
or U8855 (N_8855,N_8562,N_8654);
or U8856 (N_8856,N_8737,N_8573);
xnor U8857 (N_8857,N_8503,N_8528);
or U8858 (N_8858,N_8649,N_8677);
or U8859 (N_8859,N_8722,N_8516);
and U8860 (N_8860,N_8652,N_8600);
nand U8861 (N_8861,N_8696,N_8746);
and U8862 (N_8862,N_8572,N_8525);
or U8863 (N_8863,N_8728,N_8692);
xor U8864 (N_8864,N_8537,N_8533);
xnor U8865 (N_8865,N_8614,N_8719);
or U8866 (N_8866,N_8527,N_8663);
xor U8867 (N_8867,N_8526,N_8616);
xnor U8868 (N_8868,N_8569,N_8592);
xor U8869 (N_8869,N_8532,N_8678);
nand U8870 (N_8870,N_8523,N_8580);
and U8871 (N_8871,N_8697,N_8581);
xnor U8872 (N_8872,N_8583,N_8690);
or U8873 (N_8873,N_8512,N_8744);
nor U8874 (N_8874,N_8748,N_8556);
and U8875 (N_8875,N_8733,N_8560);
or U8876 (N_8876,N_8559,N_8660);
and U8877 (N_8877,N_8664,N_8570);
nand U8878 (N_8878,N_8592,N_8516);
nor U8879 (N_8879,N_8627,N_8554);
and U8880 (N_8880,N_8612,N_8510);
or U8881 (N_8881,N_8729,N_8686);
or U8882 (N_8882,N_8668,N_8681);
and U8883 (N_8883,N_8681,N_8644);
xor U8884 (N_8884,N_8567,N_8618);
and U8885 (N_8885,N_8639,N_8661);
xor U8886 (N_8886,N_8570,N_8667);
or U8887 (N_8887,N_8665,N_8613);
and U8888 (N_8888,N_8515,N_8626);
nor U8889 (N_8889,N_8628,N_8618);
nand U8890 (N_8890,N_8697,N_8545);
nor U8891 (N_8891,N_8665,N_8729);
nand U8892 (N_8892,N_8626,N_8653);
nor U8893 (N_8893,N_8644,N_8519);
and U8894 (N_8894,N_8562,N_8546);
nand U8895 (N_8895,N_8712,N_8714);
or U8896 (N_8896,N_8729,N_8742);
or U8897 (N_8897,N_8726,N_8673);
xnor U8898 (N_8898,N_8715,N_8505);
nor U8899 (N_8899,N_8564,N_8534);
or U8900 (N_8900,N_8505,N_8579);
nand U8901 (N_8901,N_8739,N_8727);
or U8902 (N_8902,N_8696,N_8502);
nor U8903 (N_8903,N_8669,N_8512);
nand U8904 (N_8904,N_8715,N_8524);
nor U8905 (N_8905,N_8747,N_8598);
nor U8906 (N_8906,N_8644,N_8709);
xnor U8907 (N_8907,N_8692,N_8635);
or U8908 (N_8908,N_8612,N_8687);
xnor U8909 (N_8909,N_8503,N_8651);
or U8910 (N_8910,N_8681,N_8710);
and U8911 (N_8911,N_8623,N_8745);
and U8912 (N_8912,N_8529,N_8649);
or U8913 (N_8913,N_8584,N_8692);
or U8914 (N_8914,N_8711,N_8736);
nand U8915 (N_8915,N_8658,N_8574);
xnor U8916 (N_8916,N_8676,N_8710);
nor U8917 (N_8917,N_8744,N_8534);
nor U8918 (N_8918,N_8694,N_8621);
and U8919 (N_8919,N_8578,N_8724);
or U8920 (N_8920,N_8720,N_8508);
or U8921 (N_8921,N_8511,N_8534);
nor U8922 (N_8922,N_8700,N_8607);
xnor U8923 (N_8923,N_8579,N_8737);
xnor U8924 (N_8924,N_8710,N_8573);
nand U8925 (N_8925,N_8646,N_8500);
xor U8926 (N_8926,N_8679,N_8618);
and U8927 (N_8927,N_8563,N_8630);
xor U8928 (N_8928,N_8742,N_8663);
and U8929 (N_8929,N_8553,N_8577);
xnor U8930 (N_8930,N_8588,N_8520);
xnor U8931 (N_8931,N_8741,N_8747);
and U8932 (N_8932,N_8504,N_8517);
or U8933 (N_8933,N_8697,N_8564);
xor U8934 (N_8934,N_8667,N_8549);
nor U8935 (N_8935,N_8628,N_8702);
nand U8936 (N_8936,N_8749,N_8651);
or U8937 (N_8937,N_8579,N_8615);
nor U8938 (N_8938,N_8642,N_8510);
or U8939 (N_8939,N_8598,N_8713);
or U8940 (N_8940,N_8578,N_8587);
or U8941 (N_8941,N_8528,N_8726);
and U8942 (N_8942,N_8748,N_8605);
or U8943 (N_8943,N_8558,N_8715);
nand U8944 (N_8944,N_8634,N_8717);
or U8945 (N_8945,N_8559,N_8530);
xnor U8946 (N_8946,N_8705,N_8619);
nand U8947 (N_8947,N_8625,N_8702);
nor U8948 (N_8948,N_8544,N_8569);
nor U8949 (N_8949,N_8704,N_8601);
nand U8950 (N_8950,N_8560,N_8749);
nand U8951 (N_8951,N_8510,N_8747);
and U8952 (N_8952,N_8581,N_8741);
nand U8953 (N_8953,N_8742,N_8641);
or U8954 (N_8954,N_8676,N_8529);
xor U8955 (N_8955,N_8538,N_8542);
and U8956 (N_8956,N_8587,N_8547);
or U8957 (N_8957,N_8640,N_8547);
or U8958 (N_8958,N_8600,N_8656);
nand U8959 (N_8959,N_8634,N_8588);
xnor U8960 (N_8960,N_8725,N_8669);
and U8961 (N_8961,N_8616,N_8596);
xor U8962 (N_8962,N_8625,N_8664);
or U8963 (N_8963,N_8539,N_8651);
xor U8964 (N_8964,N_8597,N_8615);
nor U8965 (N_8965,N_8567,N_8713);
nand U8966 (N_8966,N_8672,N_8690);
nand U8967 (N_8967,N_8679,N_8549);
nand U8968 (N_8968,N_8546,N_8617);
or U8969 (N_8969,N_8516,N_8622);
nor U8970 (N_8970,N_8706,N_8592);
nor U8971 (N_8971,N_8569,N_8545);
xor U8972 (N_8972,N_8596,N_8575);
or U8973 (N_8973,N_8664,N_8532);
nor U8974 (N_8974,N_8731,N_8707);
or U8975 (N_8975,N_8661,N_8620);
nor U8976 (N_8976,N_8578,N_8505);
nor U8977 (N_8977,N_8703,N_8604);
nor U8978 (N_8978,N_8595,N_8710);
or U8979 (N_8979,N_8649,N_8558);
and U8980 (N_8980,N_8591,N_8541);
and U8981 (N_8981,N_8594,N_8530);
nand U8982 (N_8982,N_8514,N_8637);
xor U8983 (N_8983,N_8598,N_8551);
or U8984 (N_8984,N_8503,N_8635);
and U8985 (N_8985,N_8564,N_8565);
and U8986 (N_8986,N_8675,N_8582);
xnor U8987 (N_8987,N_8743,N_8534);
xor U8988 (N_8988,N_8670,N_8730);
and U8989 (N_8989,N_8730,N_8718);
nand U8990 (N_8990,N_8688,N_8553);
xnor U8991 (N_8991,N_8740,N_8648);
xnor U8992 (N_8992,N_8716,N_8736);
or U8993 (N_8993,N_8680,N_8503);
or U8994 (N_8994,N_8689,N_8686);
xnor U8995 (N_8995,N_8690,N_8684);
nand U8996 (N_8996,N_8725,N_8590);
or U8997 (N_8997,N_8670,N_8510);
xnor U8998 (N_8998,N_8691,N_8624);
or U8999 (N_8999,N_8545,N_8630);
and U9000 (N_9000,N_8924,N_8995);
and U9001 (N_9001,N_8794,N_8888);
and U9002 (N_9002,N_8841,N_8997);
and U9003 (N_9003,N_8882,N_8805);
or U9004 (N_9004,N_8867,N_8915);
and U9005 (N_9005,N_8777,N_8843);
nor U9006 (N_9006,N_8968,N_8858);
nor U9007 (N_9007,N_8880,N_8821);
or U9008 (N_9008,N_8904,N_8938);
nand U9009 (N_9009,N_8900,N_8866);
or U9010 (N_9010,N_8793,N_8881);
nor U9011 (N_9011,N_8918,N_8790);
nand U9012 (N_9012,N_8943,N_8911);
nor U9013 (N_9013,N_8807,N_8992);
and U9014 (N_9014,N_8934,N_8897);
nor U9015 (N_9015,N_8811,N_8855);
xor U9016 (N_9016,N_8975,N_8874);
or U9017 (N_9017,N_8788,N_8956);
nand U9018 (N_9018,N_8966,N_8906);
xor U9019 (N_9019,N_8871,N_8998);
or U9020 (N_9020,N_8800,N_8981);
nand U9021 (N_9021,N_8856,N_8823);
and U9022 (N_9022,N_8953,N_8809);
and U9023 (N_9023,N_8872,N_8802);
nand U9024 (N_9024,N_8927,N_8849);
xnor U9025 (N_9025,N_8854,N_8772);
nand U9026 (N_9026,N_8842,N_8973);
or U9027 (N_9027,N_8761,N_8864);
or U9028 (N_9028,N_8781,N_8862);
and U9029 (N_9029,N_8891,N_8776);
xor U9030 (N_9030,N_8839,N_8860);
and U9031 (N_9031,N_8758,N_8948);
xnor U9032 (N_9032,N_8806,N_8785);
nand U9033 (N_9033,N_8912,N_8831);
or U9034 (N_9034,N_8914,N_8847);
nand U9035 (N_9035,N_8898,N_8991);
xor U9036 (N_9036,N_8893,N_8869);
and U9037 (N_9037,N_8835,N_8766);
xnor U9038 (N_9038,N_8949,N_8901);
nand U9039 (N_9039,N_8926,N_8764);
nand U9040 (N_9040,N_8762,N_8907);
and U9041 (N_9041,N_8786,N_8894);
and U9042 (N_9042,N_8814,N_8878);
xor U9043 (N_9043,N_8752,N_8851);
or U9044 (N_9044,N_8773,N_8952);
nor U9045 (N_9045,N_8988,N_8917);
and U9046 (N_9046,N_8768,N_8951);
or U9047 (N_9047,N_8834,N_8996);
nor U9048 (N_9048,N_8816,N_8825);
or U9049 (N_9049,N_8852,N_8928);
and U9050 (N_9050,N_8857,N_8868);
xor U9051 (N_9051,N_8879,N_8763);
or U9052 (N_9052,N_8985,N_8950);
and U9053 (N_9053,N_8939,N_8769);
or U9054 (N_9054,N_8982,N_8797);
nor U9055 (N_9055,N_8765,N_8795);
nor U9056 (N_9056,N_8770,N_8941);
nor U9057 (N_9057,N_8885,N_8916);
nand U9058 (N_9058,N_8970,N_8959);
and U9059 (N_9059,N_8824,N_8799);
xor U9060 (N_9060,N_8960,N_8845);
nand U9061 (N_9061,N_8784,N_8962);
and U9062 (N_9062,N_8896,N_8961);
nor U9063 (N_9063,N_8910,N_8853);
or U9064 (N_9064,N_8774,N_8837);
nand U9065 (N_9065,N_8830,N_8993);
and U9066 (N_9066,N_8899,N_8999);
and U9067 (N_9067,N_8930,N_8875);
and U9068 (N_9068,N_8889,N_8944);
or U9069 (N_9069,N_8971,N_8820);
or U9070 (N_9070,N_8919,N_8829);
nor U9071 (N_9071,N_8753,N_8755);
and U9072 (N_9072,N_8945,N_8958);
xnor U9073 (N_9073,N_8801,N_8848);
and U9074 (N_9074,N_8778,N_8932);
xor U9075 (N_9075,N_8771,N_8780);
nor U9076 (N_9076,N_8979,N_8972);
nand U9077 (N_9077,N_8895,N_8832);
nand U9078 (N_9078,N_8873,N_8808);
and U9079 (N_9079,N_8813,N_8908);
nand U9080 (N_9080,N_8756,N_8980);
or U9081 (N_9081,N_8986,N_8990);
xor U9082 (N_9082,N_8886,N_8922);
and U9083 (N_9083,N_8798,N_8957);
and U9084 (N_9084,N_8983,N_8965);
and U9085 (N_9085,N_8810,N_8890);
nand U9086 (N_9086,N_8994,N_8936);
and U9087 (N_9087,N_8978,N_8844);
xnor U9088 (N_9088,N_8977,N_8840);
or U9089 (N_9089,N_8789,N_8779);
and U9090 (N_9090,N_8796,N_8955);
or U9091 (N_9091,N_8850,N_8947);
nand U9092 (N_9092,N_8923,N_8818);
nand U9093 (N_9093,N_8935,N_8940);
xnor U9094 (N_9094,N_8751,N_8876);
and U9095 (N_9095,N_8946,N_8921);
nor U9096 (N_9096,N_8803,N_8887);
and U9097 (N_9097,N_8933,N_8838);
nor U9098 (N_9098,N_8836,N_8937);
or U9099 (N_9099,N_8984,N_8963);
nor U9100 (N_9100,N_8791,N_8759);
nand U9101 (N_9101,N_8792,N_8913);
nor U9102 (N_9102,N_8920,N_8909);
xnor U9103 (N_9103,N_8883,N_8969);
or U9104 (N_9104,N_8767,N_8754);
or U9105 (N_9105,N_8884,N_8833);
nor U9106 (N_9106,N_8757,N_8877);
and U9107 (N_9107,N_8817,N_8815);
and U9108 (N_9108,N_8987,N_8931);
and U9109 (N_9109,N_8905,N_8812);
xor U9110 (N_9110,N_8861,N_8783);
xnor U9111 (N_9111,N_8819,N_8976);
nor U9112 (N_9112,N_8863,N_8826);
nand U9113 (N_9113,N_8967,N_8859);
xnor U9114 (N_9114,N_8828,N_8989);
or U9115 (N_9115,N_8775,N_8925);
or U9116 (N_9116,N_8974,N_8846);
xor U9117 (N_9117,N_8870,N_8750);
nor U9118 (N_9118,N_8827,N_8787);
nand U9119 (N_9119,N_8942,N_8902);
nand U9120 (N_9120,N_8929,N_8964);
and U9121 (N_9121,N_8903,N_8804);
xnor U9122 (N_9122,N_8760,N_8865);
nand U9123 (N_9123,N_8892,N_8782);
xor U9124 (N_9124,N_8822,N_8954);
nand U9125 (N_9125,N_8752,N_8818);
xor U9126 (N_9126,N_8837,N_8997);
and U9127 (N_9127,N_8872,N_8994);
or U9128 (N_9128,N_8855,N_8952);
nor U9129 (N_9129,N_8987,N_8911);
nor U9130 (N_9130,N_8941,N_8787);
or U9131 (N_9131,N_8822,N_8820);
and U9132 (N_9132,N_8769,N_8879);
nand U9133 (N_9133,N_8882,N_8817);
and U9134 (N_9134,N_8899,N_8938);
xor U9135 (N_9135,N_8954,N_8878);
or U9136 (N_9136,N_8873,N_8800);
xnor U9137 (N_9137,N_8813,N_8970);
nand U9138 (N_9138,N_8992,N_8959);
xnor U9139 (N_9139,N_8968,N_8752);
nor U9140 (N_9140,N_8915,N_8837);
and U9141 (N_9141,N_8860,N_8915);
or U9142 (N_9142,N_8805,N_8826);
xnor U9143 (N_9143,N_8877,N_8755);
and U9144 (N_9144,N_8862,N_8941);
or U9145 (N_9145,N_8769,N_8866);
nand U9146 (N_9146,N_8987,N_8777);
or U9147 (N_9147,N_8970,N_8935);
and U9148 (N_9148,N_8764,N_8999);
nor U9149 (N_9149,N_8914,N_8872);
xor U9150 (N_9150,N_8969,N_8977);
nand U9151 (N_9151,N_8817,N_8916);
or U9152 (N_9152,N_8992,N_8924);
xor U9153 (N_9153,N_8766,N_8871);
xor U9154 (N_9154,N_8898,N_8965);
and U9155 (N_9155,N_8780,N_8828);
or U9156 (N_9156,N_8873,N_8838);
or U9157 (N_9157,N_8788,N_8929);
xnor U9158 (N_9158,N_8861,N_8884);
or U9159 (N_9159,N_8884,N_8848);
nand U9160 (N_9160,N_8860,N_8808);
xnor U9161 (N_9161,N_8905,N_8764);
nor U9162 (N_9162,N_8773,N_8903);
and U9163 (N_9163,N_8875,N_8984);
nand U9164 (N_9164,N_8982,N_8993);
and U9165 (N_9165,N_8902,N_8813);
nor U9166 (N_9166,N_8951,N_8978);
and U9167 (N_9167,N_8886,N_8857);
nand U9168 (N_9168,N_8781,N_8810);
nor U9169 (N_9169,N_8861,N_8974);
xnor U9170 (N_9170,N_8852,N_8770);
nor U9171 (N_9171,N_8793,N_8811);
or U9172 (N_9172,N_8908,N_8872);
xor U9173 (N_9173,N_8776,N_8804);
nor U9174 (N_9174,N_8838,N_8772);
nand U9175 (N_9175,N_8988,N_8950);
xnor U9176 (N_9176,N_8914,N_8770);
nand U9177 (N_9177,N_8792,N_8991);
nand U9178 (N_9178,N_8777,N_8828);
xnor U9179 (N_9179,N_8836,N_8764);
or U9180 (N_9180,N_8914,N_8782);
xor U9181 (N_9181,N_8931,N_8973);
nand U9182 (N_9182,N_8943,N_8774);
xnor U9183 (N_9183,N_8988,N_8846);
or U9184 (N_9184,N_8939,N_8782);
and U9185 (N_9185,N_8831,N_8943);
and U9186 (N_9186,N_8968,N_8940);
nand U9187 (N_9187,N_8771,N_8799);
nand U9188 (N_9188,N_8908,N_8825);
or U9189 (N_9189,N_8759,N_8796);
xor U9190 (N_9190,N_8837,N_8938);
nand U9191 (N_9191,N_8925,N_8952);
and U9192 (N_9192,N_8997,N_8797);
nor U9193 (N_9193,N_8851,N_8915);
xor U9194 (N_9194,N_8996,N_8963);
nand U9195 (N_9195,N_8983,N_8951);
xor U9196 (N_9196,N_8880,N_8969);
nand U9197 (N_9197,N_8999,N_8929);
nand U9198 (N_9198,N_8814,N_8931);
xnor U9199 (N_9199,N_8994,N_8966);
xor U9200 (N_9200,N_8784,N_8780);
nand U9201 (N_9201,N_8763,N_8901);
xnor U9202 (N_9202,N_8843,N_8836);
and U9203 (N_9203,N_8900,N_8916);
nand U9204 (N_9204,N_8928,N_8819);
or U9205 (N_9205,N_8913,N_8812);
or U9206 (N_9206,N_8752,N_8754);
or U9207 (N_9207,N_8805,N_8915);
and U9208 (N_9208,N_8990,N_8822);
xnor U9209 (N_9209,N_8792,N_8773);
nand U9210 (N_9210,N_8919,N_8906);
and U9211 (N_9211,N_8899,N_8753);
and U9212 (N_9212,N_8754,N_8801);
or U9213 (N_9213,N_8861,N_8989);
nand U9214 (N_9214,N_8927,N_8993);
nand U9215 (N_9215,N_8928,N_8929);
xor U9216 (N_9216,N_8840,N_8968);
and U9217 (N_9217,N_8810,N_8991);
nand U9218 (N_9218,N_8780,N_8898);
nand U9219 (N_9219,N_8971,N_8816);
nor U9220 (N_9220,N_8924,N_8791);
nand U9221 (N_9221,N_8756,N_8869);
or U9222 (N_9222,N_8772,N_8849);
and U9223 (N_9223,N_8909,N_8893);
xor U9224 (N_9224,N_8910,N_8958);
and U9225 (N_9225,N_8980,N_8952);
nor U9226 (N_9226,N_8908,N_8796);
and U9227 (N_9227,N_8785,N_8935);
nor U9228 (N_9228,N_8765,N_8905);
nand U9229 (N_9229,N_8782,N_8791);
or U9230 (N_9230,N_8829,N_8816);
or U9231 (N_9231,N_8780,N_8835);
or U9232 (N_9232,N_8957,N_8883);
or U9233 (N_9233,N_8874,N_8882);
nor U9234 (N_9234,N_8992,N_8857);
nand U9235 (N_9235,N_8997,N_8894);
nor U9236 (N_9236,N_8779,N_8782);
nor U9237 (N_9237,N_8969,N_8833);
or U9238 (N_9238,N_8754,N_8757);
nor U9239 (N_9239,N_8930,N_8754);
or U9240 (N_9240,N_8965,N_8903);
and U9241 (N_9241,N_8904,N_8790);
and U9242 (N_9242,N_8996,N_8961);
or U9243 (N_9243,N_8995,N_8915);
nor U9244 (N_9244,N_8895,N_8858);
xor U9245 (N_9245,N_8751,N_8942);
or U9246 (N_9246,N_8903,N_8877);
xor U9247 (N_9247,N_8756,N_8918);
nand U9248 (N_9248,N_8942,N_8864);
xor U9249 (N_9249,N_8863,N_8964);
and U9250 (N_9250,N_9231,N_9220);
or U9251 (N_9251,N_9198,N_9014);
nand U9252 (N_9252,N_9227,N_9083);
and U9253 (N_9253,N_9110,N_9242);
xnor U9254 (N_9254,N_9101,N_9208);
or U9255 (N_9255,N_9230,N_9248);
nor U9256 (N_9256,N_9049,N_9059);
nand U9257 (N_9257,N_9028,N_9179);
or U9258 (N_9258,N_9195,N_9247);
nand U9259 (N_9259,N_9181,N_9016);
nor U9260 (N_9260,N_9190,N_9022);
nand U9261 (N_9261,N_9147,N_9001);
nor U9262 (N_9262,N_9152,N_9085);
nor U9263 (N_9263,N_9238,N_9205);
xnor U9264 (N_9264,N_9113,N_9052);
nand U9265 (N_9265,N_9031,N_9019);
or U9266 (N_9266,N_9105,N_9235);
or U9267 (N_9267,N_9011,N_9237);
or U9268 (N_9268,N_9140,N_9005);
nand U9269 (N_9269,N_9174,N_9175);
and U9270 (N_9270,N_9221,N_9162);
or U9271 (N_9271,N_9044,N_9153);
nor U9272 (N_9272,N_9020,N_9056);
xnor U9273 (N_9273,N_9197,N_9021);
and U9274 (N_9274,N_9009,N_9121);
nand U9275 (N_9275,N_9050,N_9201);
nor U9276 (N_9276,N_9004,N_9035);
xnor U9277 (N_9277,N_9047,N_9074);
nand U9278 (N_9278,N_9077,N_9082);
and U9279 (N_9279,N_9106,N_9115);
and U9280 (N_9280,N_9057,N_9128);
xnor U9281 (N_9281,N_9144,N_9245);
nor U9282 (N_9282,N_9088,N_9094);
nor U9283 (N_9283,N_9203,N_9062);
nand U9284 (N_9284,N_9239,N_9224);
nor U9285 (N_9285,N_9109,N_9058);
xor U9286 (N_9286,N_9167,N_9233);
nor U9287 (N_9287,N_9232,N_9145);
xor U9288 (N_9288,N_9182,N_9165);
nand U9289 (N_9289,N_9142,N_9084);
nand U9290 (N_9290,N_9158,N_9071);
and U9291 (N_9291,N_9054,N_9229);
nor U9292 (N_9292,N_9099,N_9169);
nand U9293 (N_9293,N_9068,N_9124);
or U9294 (N_9294,N_9012,N_9129);
xnor U9295 (N_9295,N_9100,N_9200);
and U9296 (N_9296,N_9244,N_9069);
and U9297 (N_9297,N_9075,N_9225);
nor U9298 (N_9298,N_9161,N_9150);
xor U9299 (N_9299,N_9191,N_9055);
nand U9300 (N_9300,N_9163,N_9070);
or U9301 (N_9301,N_9032,N_9051);
xnor U9302 (N_9302,N_9078,N_9234);
nor U9303 (N_9303,N_9199,N_9013);
xor U9304 (N_9304,N_9192,N_9060);
or U9305 (N_9305,N_9146,N_9159);
nor U9306 (N_9306,N_9210,N_9103);
nor U9307 (N_9307,N_9076,N_9039);
and U9308 (N_9308,N_9118,N_9185);
nand U9309 (N_9309,N_9102,N_9137);
nor U9310 (N_9310,N_9092,N_9126);
and U9311 (N_9311,N_9030,N_9127);
and U9312 (N_9312,N_9213,N_9176);
xnor U9313 (N_9313,N_9006,N_9002);
xnor U9314 (N_9314,N_9193,N_9236);
and U9315 (N_9315,N_9148,N_9133);
nand U9316 (N_9316,N_9202,N_9029);
nor U9317 (N_9317,N_9024,N_9061);
nor U9318 (N_9318,N_9108,N_9156);
nand U9319 (N_9319,N_9122,N_9170);
or U9320 (N_9320,N_9041,N_9007);
nor U9321 (N_9321,N_9037,N_9120);
nor U9322 (N_9322,N_9093,N_9164);
nand U9323 (N_9323,N_9160,N_9194);
or U9324 (N_9324,N_9131,N_9135);
or U9325 (N_9325,N_9119,N_9017);
nand U9326 (N_9326,N_9228,N_9080);
or U9327 (N_9327,N_9215,N_9243);
nand U9328 (N_9328,N_9072,N_9114);
and U9329 (N_9329,N_9067,N_9155);
nand U9330 (N_9330,N_9217,N_9036);
or U9331 (N_9331,N_9154,N_9063);
nand U9332 (N_9332,N_9204,N_9218);
nand U9333 (N_9333,N_9151,N_9180);
nor U9334 (N_9334,N_9048,N_9040);
and U9335 (N_9335,N_9089,N_9149);
nor U9336 (N_9336,N_9023,N_9186);
nand U9337 (N_9337,N_9184,N_9177);
and U9338 (N_9338,N_9222,N_9141);
and U9339 (N_9339,N_9206,N_9046);
nor U9340 (N_9340,N_9079,N_9189);
and U9341 (N_9341,N_9064,N_9216);
nand U9342 (N_9342,N_9018,N_9223);
nand U9343 (N_9343,N_9168,N_9132);
xnor U9344 (N_9344,N_9178,N_9095);
nor U9345 (N_9345,N_9015,N_9211);
or U9346 (N_9346,N_9000,N_9171);
or U9347 (N_9347,N_9134,N_9104);
nor U9348 (N_9348,N_9136,N_9246);
nand U9349 (N_9349,N_9065,N_9086);
or U9350 (N_9350,N_9081,N_9045);
nand U9351 (N_9351,N_9173,N_9008);
or U9352 (N_9352,N_9003,N_9025);
or U9353 (N_9353,N_9172,N_9096);
or U9354 (N_9354,N_9196,N_9125);
or U9355 (N_9355,N_9241,N_9112);
or U9356 (N_9356,N_9187,N_9026);
or U9357 (N_9357,N_9066,N_9034);
and U9358 (N_9358,N_9130,N_9053);
xnor U9359 (N_9359,N_9116,N_9107);
xor U9360 (N_9360,N_9033,N_9138);
and U9361 (N_9361,N_9207,N_9157);
xnor U9362 (N_9362,N_9143,N_9212);
or U9363 (N_9363,N_9249,N_9219);
or U9364 (N_9364,N_9139,N_9166);
nand U9365 (N_9365,N_9117,N_9214);
nand U9366 (N_9366,N_9111,N_9043);
nand U9367 (N_9367,N_9027,N_9183);
nor U9368 (N_9368,N_9073,N_9091);
or U9369 (N_9369,N_9226,N_9038);
nand U9370 (N_9370,N_9240,N_9042);
nand U9371 (N_9371,N_9123,N_9188);
and U9372 (N_9372,N_9097,N_9209);
or U9373 (N_9373,N_9087,N_9010);
or U9374 (N_9374,N_9090,N_9098);
xnor U9375 (N_9375,N_9093,N_9039);
nor U9376 (N_9376,N_9163,N_9110);
nand U9377 (N_9377,N_9248,N_9222);
nand U9378 (N_9378,N_9056,N_9088);
nand U9379 (N_9379,N_9119,N_9190);
or U9380 (N_9380,N_9212,N_9113);
nor U9381 (N_9381,N_9211,N_9066);
xnor U9382 (N_9382,N_9094,N_9201);
xor U9383 (N_9383,N_9046,N_9061);
xnor U9384 (N_9384,N_9054,N_9178);
xnor U9385 (N_9385,N_9114,N_9020);
nand U9386 (N_9386,N_9050,N_9030);
nor U9387 (N_9387,N_9061,N_9202);
xnor U9388 (N_9388,N_9106,N_9126);
nand U9389 (N_9389,N_9122,N_9139);
or U9390 (N_9390,N_9138,N_9230);
nand U9391 (N_9391,N_9145,N_9118);
or U9392 (N_9392,N_9063,N_9131);
xnor U9393 (N_9393,N_9241,N_9122);
and U9394 (N_9394,N_9161,N_9167);
xor U9395 (N_9395,N_9094,N_9051);
or U9396 (N_9396,N_9065,N_9042);
xnor U9397 (N_9397,N_9085,N_9101);
or U9398 (N_9398,N_9233,N_9238);
and U9399 (N_9399,N_9207,N_9179);
and U9400 (N_9400,N_9248,N_9106);
xnor U9401 (N_9401,N_9134,N_9056);
nor U9402 (N_9402,N_9002,N_9092);
and U9403 (N_9403,N_9005,N_9129);
xor U9404 (N_9404,N_9199,N_9181);
and U9405 (N_9405,N_9188,N_9105);
xor U9406 (N_9406,N_9222,N_9166);
xor U9407 (N_9407,N_9236,N_9198);
nand U9408 (N_9408,N_9181,N_9154);
and U9409 (N_9409,N_9149,N_9115);
xnor U9410 (N_9410,N_9247,N_9083);
xnor U9411 (N_9411,N_9048,N_9068);
nand U9412 (N_9412,N_9152,N_9162);
nand U9413 (N_9413,N_9022,N_9179);
or U9414 (N_9414,N_9092,N_9115);
xor U9415 (N_9415,N_9037,N_9102);
or U9416 (N_9416,N_9236,N_9177);
nand U9417 (N_9417,N_9016,N_9099);
or U9418 (N_9418,N_9127,N_9080);
nand U9419 (N_9419,N_9018,N_9005);
nand U9420 (N_9420,N_9069,N_9038);
nor U9421 (N_9421,N_9232,N_9212);
xor U9422 (N_9422,N_9000,N_9181);
or U9423 (N_9423,N_9029,N_9170);
and U9424 (N_9424,N_9218,N_9152);
nor U9425 (N_9425,N_9112,N_9246);
and U9426 (N_9426,N_9242,N_9114);
nor U9427 (N_9427,N_9149,N_9153);
xor U9428 (N_9428,N_9159,N_9206);
nand U9429 (N_9429,N_9231,N_9089);
nand U9430 (N_9430,N_9197,N_9115);
and U9431 (N_9431,N_9056,N_9242);
or U9432 (N_9432,N_9089,N_9188);
xor U9433 (N_9433,N_9245,N_9028);
nor U9434 (N_9434,N_9122,N_9073);
nor U9435 (N_9435,N_9134,N_9118);
xnor U9436 (N_9436,N_9134,N_9231);
or U9437 (N_9437,N_9242,N_9023);
nor U9438 (N_9438,N_9141,N_9034);
nand U9439 (N_9439,N_9205,N_9018);
and U9440 (N_9440,N_9178,N_9191);
or U9441 (N_9441,N_9159,N_9044);
nand U9442 (N_9442,N_9181,N_9166);
nor U9443 (N_9443,N_9024,N_9201);
or U9444 (N_9444,N_9174,N_9139);
xnor U9445 (N_9445,N_9135,N_9090);
and U9446 (N_9446,N_9101,N_9216);
nor U9447 (N_9447,N_9032,N_9048);
nor U9448 (N_9448,N_9025,N_9060);
or U9449 (N_9449,N_9028,N_9182);
nor U9450 (N_9450,N_9095,N_9160);
xor U9451 (N_9451,N_9009,N_9010);
nand U9452 (N_9452,N_9228,N_9106);
nand U9453 (N_9453,N_9028,N_9185);
and U9454 (N_9454,N_9177,N_9009);
xor U9455 (N_9455,N_9196,N_9015);
xnor U9456 (N_9456,N_9032,N_9142);
and U9457 (N_9457,N_9108,N_9055);
nor U9458 (N_9458,N_9175,N_9042);
or U9459 (N_9459,N_9065,N_9163);
and U9460 (N_9460,N_9220,N_9091);
and U9461 (N_9461,N_9228,N_9170);
xnor U9462 (N_9462,N_9195,N_9132);
nand U9463 (N_9463,N_9034,N_9101);
xor U9464 (N_9464,N_9240,N_9065);
or U9465 (N_9465,N_9184,N_9097);
nand U9466 (N_9466,N_9056,N_9097);
nand U9467 (N_9467,N_9080,N_9161);
nor U9468 (N_9468,N_9239,N_9083);
xnor U9469 (N_9469,N_9011,N_9073);
nand U9470 (N_9470,N_9170,N_9059);
nand U9471 (N_9471,N_9194,N_9045);
nor U9472 (N_9472,N_9133,N_9097);
and U9473 (N_9473,N_9170,N_9161);
nand U9474 (N_9474,N_9034,N_9155);
or U9475 (N_9475,N_9130,N_9042);
or U9476 (N_9476,N_9191,N_9225);
xnor U9477 (N_9477,N_9010,N_9153);
nor U9478 (N_9478,N_9065,N_9152);
and U9479 (N_9479,N_9134,N_9045);
xor U9480 (N_9480,N_9169,N_9003);
nand U9481 (N_9481,N_9037,N_9129);
nor U9482 (N_9482,N_9209,N_9219);
nand U9483 (N_9483,N_9242,N_9222);
or U9484 (N_9484,N_9115,N_9095);
nand U9485 (N_9485,N_9064,N_9122);
nor U9486 (N_9486,N_9248,N_9247);
xnor U9487 (N_9487,N_9177,N_9103);
nand U9488 (N_9488,N_9249,N_9182);
nand U9489 (N_9489,N_9044,N_9188);
nand U9490 (N_9490,N_9041,N_9010);
and U9491 (N_9491,N_9231,N_9000);
xor U9492 (N_9492,N_9072,N_9172);
and U9493 (N_9493,N_9101,N_9246);
and U9494 (N_9494,N_9185,N_9034);
nand U9495 (N_9495,N_9185,N_9138);
or U9496 (N_9496,N_9239,N_9103);
xnor U9497 (N_9497,N_9210,N_9185);
nand U9498 (N_9498,N_9001,N_9159);
nor U9499 (N_9499,N_9173,N_9244);
nand U9500 (N_9500,N_9410,N_9353);
or U9501 (N_9501,N_9438,N_9429);
nand U9502 (N_9502,N_9315,N_9499);
nor U9503 (N_9503,N_9405,N_9397);
nand U9504 (N_9504,N_9345,N_9275);
or U9505 (N_9505,N_9350,N_9332);
nor U9506 (N_9506,N_9313,N_9450);
nand U9507 (N_9507,N_9372,N_9461);
nor U9508 (N_9508,N_9280,N_9263);
nand U9509 (N_9509,N_9412,N_9423);
or U9510 (N_9510,N_9362,N_9377);
nand U9511 (N_9511,N_9401,N_9347);
nand U9512 (N_9512,N_9383,N_9409);
nor U9513 (N_9513,N_9445,N_9258);
xnor U9514 (N_9514,N_9467,N_9300);
nor U9515 (N_9515,N_9376,N_9355);
xnor U9516 (N_9516,N_9322,N_9305);
and U9517 (N_9517,N_9432,N_9491);
nand U9518 (N_9518,N_9433,N_9308);
and U9519 (N_9519,N_9443,N_9449);
nor U9520 (N_9520,N_9428,N_9329);
and U9521 (N_9521,N_9488,N_9250);
xor U9522 (N_9522,N_9414,N_9320);
and U9523 (N_9523,N_9311,N_9312);
nand U9524 (N_9524,N_9317,N_9382);
nor U9525 (N_9525,N_9498,N_9484);
nand U9526 (N_9526,N_9454,N_9319);
or U9527 (N_9527,N_9289,N_9463);
and U9528 (N_9528,N_9333,N_9442);
nor U9529 (N_9529,N_9477,N_9493);
and U9530 (N_9530,N_9469,N_9371);
or U9531 (N_9531,N_9437,N_9259);
xor U9532 (N_9532,N_9381,N_9490);
and U9533 (N_9533,N_9406,N_9261);
xnor U9534 (N_9534,N_9391,N_9465);
or U9535 (N_9535,N_9394,N_9494);
and U9536 (N_9536,N_9367,N_9393);
or U9537 (N_9537,N_9358,N_9451);
or U9538 (N_9538,N_9257,N_9421);
or U9539 (N_9539,N_9495,N_9361);
and U9540 (N_9540,N_9473,N_9496);
or U9541 (N_9541,N_9339,N_9307);
and U9542 (N_9542,N_9457,N_9277);
nand U9543 (N_9543,N_9349,N_9266);
or U9544 (N_9544,N_9336,N_9483);
nand U9545 (N_9545,N_9486,N_9369);
and U9546 (N_9546,N_9388,N_9286);
and U9547 (N_9547,N_9265,N_9459);
or U9548 (N_9548,N_9373,N_9267);
nand U9549 (N_9549,N_9420,N_9385);
xor U9550 (N_9550,N_9256,N_9447);
nand U9551 (N_9551,N_9400,N_9364);
or U9552 (N_9552,N_9379,N_9341);
nor U9553 (N_9553,N_9416,N_9344);
xor U9554 (N_9554,N_9294,N_9298);
xnor U9555 (N_9555,N_9321,N_9476);
or U9556 (N_9556,N_9368,N_9328);
xnor U9557 (N_9557,N_9310,N_9403);
and U9558 (N_9558,N_9471,N_9268);
and U9559 (N_9559,N_9303,N_9466);
or U9560 (N_9560,N_9431,N_9448);
nand U9561 (N_9561,N_9352,N_9297);
nor U9562 (N_9562,N_9402,N_9331);
xnor U9563 (N_9563,N_9456,N_9276);
xor U9564 (N_9564,N_9482,N_9343);
or U9565 (N_9565,N_9272,N_9470);
xor U9566 (N_9566,N_9478,N_9284);
xor U9567 (N_9567,N_9479,N_9252);
xor U9568 (N_9568,N_9282,N_9422);
nand U9569 (N_9569,N_9292,N_9485);
nor U9570 (N_9570,N_9399,N_9327);
or U9571 (N_9571,N_9301,N_9396);
nand U9572 (N_9572,N_9413,N_9419);
or U9573 (N_9573,N_9338,N_9254);
nor U9574 (N_9574,N_9296,N_9354);
xnor U9575 (N_9575,N_9285,N_9304);
nand U9576 (N_9576,N_9452,N_9475);
nand U9577 (N_9577,N_9489,N_9480);
and U9578 (N_9578,N_9374,N_9440);
nor U9579 (N_9579,N_9323,N_9418);
and U9580 (N_9580,N_9370,N_9337);
and U9581 (N_9581,N_9330,N_9392);
nand U9582 (N_9582,N_9288,N_9404);
nor U9583 (N_9583,N_9444,N_9253);
xnor U9584 (N_9584,N_9434,N_9346);
xnor U9585 (N_9585,N_9407,N_9281);
or U9586 (N_9586,N_9436,N_9264);
nand U9587 (N_9587,N_9424,N_9455);
nor U9588 (N_9588,N_9278,N_9340);
or U9589 (N_9589,N_9441,N_9492);
xor U9590 (N_9590,N_9375,N_9487);
and U9591 (N_9591,N_9464,N_9309);
nand U9592 (N_9592,N_9366,N_9302);
and U9593 (N_9593,N_9415,N_9299);
nand U9594 (N_9594,N_9260,N_9255);
or U9595 (N_9595,N_9318,N_9411);
or U9596 (N_9596,N_9390,N_9386);
and U9597 (N_9597,N_9295,N_9439);
nor U9598 (N_9598,N_9408,N_9481);
nor U9599 (N_9599,N_9417,N_9334);
and U9600 (N_9600,N_9324,N_9293);
xor U9601 (N_9601,N_9497,N_9453);
nor U9602 (N_9602,N_9380,N_9360);
nor U9603 (N_9603,N_9316,N_9291);
or U9604 (N_9604,N_9363,N_9357);
nand U9605 (N_9605,N_9342,N_9306);
and U9606 (N_9606,N_9389,N_9251);
or U9607 (N_9607,N_9274,N_9290);
or U9608 (N_9608,N_9426,N_9270);
nand U9609 (N_9609,N_9359,N_9468);
or U9610 (N_9610,N_9325,N_9326);
and U9611 (N_9611,N_9273,N_9398);
xnor U9612 (N_9612,N_9283,N_9279);
xnor U9613 (N_9613,N_9460,N_9395);
or U9614 (N_9614,N_9348,N_9387);
nand U9615 (N_9615,N_9458,N_9430);
nand U9616 (N_9616,N_9314,N_9271);
xnor U9617 (N_9617,N_9287,N_9435);
and U9618 (N_9618,N_9335,N_9472);
and U9619 (N_9619,N_9446,N_9356);
or U9620 (N_9620,N_9269,N_9427);
xor U9621 (N_9621,N_9262,N_9384);
nor U9622 (N_9622,N_9365,N_9378);
or U9623 (N_9623,N_9462,N_9351);
nor U9624 (N_9624,N_9474,N_9425);
or U9625 (N_9625,N_9389,N_9462);
and U9626 (N_9626,N_9463,N_9327);
and U9627 (N_9627,N_9256,N_9402);
xor U9628 (N_9628,N_9469,N_9296);
nor U9629 (N_9629,N_9473,N_9302);
and U9630 (N_9630,N_9383,N_9482);
nand U9631 (N_9631,N_9388,N_9355);
nand U9632 (N_9632,N_9260,N_9446);
or U9633 (N_9633,N_9358,N_9317);
xnor U9634 (N_9634,N_9280,N_9274);
nor U9635 (N_9635,N_9471,N_9351);
nand U9636 (N_9636,N_9252,N_9453);
nand U9637 (N_9637,N_9477,N_9327);
xnor U9638 (N_9638,N_9446,N_9275);
nand U9639 (N_9639,N_9364,N_9276);
nor U9640 (N_9640,N_9441,N_9372);
nor U9641 (N_9641,N_9422,N_9486);
and U9642 (N_9642,N_9291,N_9432);
nor U9643 (N_9643,N_9330,N_9272);
or U9644 (N_9644,N_9380,N_9424);
and U9645 (N_9645,N_9305,N_9441);
and U9646 (N_9646,N_9469,N_9340);
xor U9647 (N_9647,N_9495,N_9377);
nand U9648 (N_9648,N_9329,N_9339);
or U9649 (N_9649,N_9348,N_9296);
xor U9650 (N_9650,N_9266,N_9296);
and U9651 (N_9651,N_9413,N_9380);
nand U9652 (N_9652,N_9412,N_9269);
xor U9653 (N_9653,N_9285,N_9301);
or U9654 (N_9654,N_9309,N_9381);
or U9655 (N_9655,N_9446,N_9285);
and U9656 (N_9656,N_9401,N_9403);
nor U9657 (N_9657,N_9308,N_9255);
xnor U9658 (N_9658,N_9383,N_9479);
or U9659 (N_9659,N_9338,N_9323);
xnor U9660 (N_9660,N_9293,N_9451);
and U9661 (N_9661,N_9418,N_9436);
or U9662 (N_9662,N_9464,N_9251);
nand U9663 (N_9663,N_9354,N_9449);
xnor U9664 (N_9664,N_9467,N_9437);
nand U9665 (N_9665,N_9315,N_9278);
and U9666 (N_9666,N_9267,N_9449);
xor U9667 (N_9667,N_9283,N_9280);
xor U9668 (N_9668,N_9438,N_9303);
nand U9669 (N_9669,N_9451,N_9294);
nand U9670 (N_9670,N_9271,N_9361);
xor U9671 (N_9671,N_9305,N_9426);
nand U9672 (N_9672,N_9380,N_9377);
nor U9673 (N_9673,N_9283,N_9361);
or U9674 (N_9674,N_9495,N_9426);
and U9675 (N_9675,N_9491,N_9487);
xnor U9676 (N_9676,N_9327,N_9294);
or U9677 (N_9677,N_9340,N_9331);
nor U9678 (N_9678,N_9348,N_9347);
xor U9679 (N_9679,N_9320,N_9453);
nand U9680 (N_9680,N_9393,N_9378);
nor U9681 (N_9681,N_9255,N_9276);
or U9682 (N_9682,N_9327,N_9253);
nand U9683 (N_9683,N_9335,N_9466);
and U9684 (N_9684,N_9389,N_9289);
nor U9685 (N_9685,N_9355,N_9353);
and U9686 (N_9686,N_9485,N_9484);
xor U9687 (N_9687,N_9468,N_9436);
nor U9688 (N_9688,N_9273,N_9299);
xnor U9689 (N_9689,N_9494,N_9472);
nand U9690 (N_9690,N_9276,N_9389);
nand U9691 (N_9691,N_9483,N_9444);
nand U9692 (N_9692,N_9485,N_9353);
or U9693 (N_9693,N_9365,N_9354);
nand U9694 (N_9694,N_9415,N_9418);
and U9695 (N_9695,N_9348,N_9438);
or U9696 (N_9696,N_9405,N_9304);
nor U9697 (N_9697,N_9487,N_9414);
nor U9698 (N_9698,N_9312,N_9440);
or U9699 (N_9699,N_9270,N_9391);
nor U9700 (N_9700,N_9426,N_9402);
xnor U9701 (N_9701,N_9288,N_9395);
xnor U9702 (N_9702,N_9442,N_9254);
xnor U9703 (N_9703,N_9257,N_9280);
nand U9704 (N_9704,N_9391,N_9423);
and U9705 (N_9705,N_9487,N_9388);
and U9706 (N_9706,N_9329,N_9373);
or U9707 (N_9707,N_9310,N_9354);
nor U9708 (N_9708,N_9314,N_9284);
nand U9709 (N_9709,N_9328,N_9285);
and U9710 (N_9710,N_9488,N_9433);
and U9711 (N_9711,N_9364,N_9255);
nand U9712 (N_9712,N_9356,N_9274);
nand U9713 (N_9713,N_9429,N_9347);
and U9714 (N_9714,N_9416,N_9491);
and U9715 (N_9715,N_9320,N_9471);
or U9716 (N_9716,N_9458,N_9411);
xor U9717 (N_9717,N_9427,N_9338);
nor U9718 (N_9718,N_9402,N_9259);
and U9719 (N_9719,N_9373,N_9333);
nor U9720 (N_9720,N_9308,N_9292);
and U9721 (N_9721,N_9269,N_9495);
or U9722 (N_9722,N_9435,N_9425);
and U9723 (N_9723,N_9372,N_9307);
xnor U9724 (N_9724,N_9318,N_9385);
nand U9725 (N_9725,N_9442,N_9252);
xnor U9726 (N_9726,N_9260,N_9480);
xor U9727 (N_9727,N_9328,N_9314);
and U9728 (N_9728,N_9394,N_9253);
nor U9729 (N_9729,N_9483,N_9329);
nand U9730 (N_9730,N_9367,N_9369);
and U9731 (N_9731,N_9277,N_9338);
nor U9732 (N_9732,N_9380,N_9262);
nand U9733 (N_9733,N_9402,N_9270);
nor U9734 (N_9734,N_9309,N_9487);
xor U9735 (N_9735,N_9371,N_9303);
nand U9736 (N_9736,N_9491,N_9471);
or U9737 (N_9737,N_9298,N_9265);
and U9738 (N_9738,N_9324,N_9495);
nand U9739 (N_9739,N_9485,N_9256);
or U9740 (N_9740,N_9484,N_9377);
nand U9741 (N_9741,N_9293,N_9333);
xnor U9742 (N_9742,N_9333,N_9426);
nor U9743 (N_9743,N_9368,N_9350);
or U9744 (N_9744,N_9372,N_9417);
nand U9745 (N_9745,N_9253,N_9378);
xnor U9746 (N_9746,N_9290,N_9401);
nand U9747 (N_9747,N_9455,N_9439);
xnor U9748 (N_9748,N_9331,N_9375);
nand U9749 (N_9749,N_9459,N_9424);
nor U9750 (N_9750,N_9565,N_9728);
and U9751 (N_9751,N_9617,N_9684);
or U9752 (N_9752,N_9574,N_9519);
xnor U9753 (N_9753,N_9676,N_9735);
and U9754 (N_9754,N_9711,N_9545);
xor U9755 (N_9755,N_9616,N_9668);
and U9756 (N_9756,N_9707,N_9725);
or U9757 (N_9757,N_9609,N_9556);
nor U9758 (N_9758,N_9700,N_9723);
nand U9759 (N_9759,N_9720,N_9511);
and U9760 (N_9760,N_9525,N_9583);
and U9761 (N_9761,N_9528,N_9628);
or U9762 (N_9762,N_9693,N_9550);
nor U9763 (N_9763,N_9591,N_9566);
nand U9764 (N_9764,N_9585,N_9548);
and U9765 (N_9765,N_9503,N_9549);
nor U9766 (N_9766,N_9569,N_9655);
or U9767 (N_9767,N_9577,N_9664);
and U9768 (N_9768,N_9680,N_9739);
nand U9769 (N_9769,N_9516,N_9660);
or U9770 (N_9770,N_9532,N_9696);
nand U9771 (N_9771,N_9709,N_9554);
nand U9772 (N_9772,N_9698,N_9636);
xnor U9773 (N_9773,N_9691,N_9702);
or U9774 (N_9774,N_9500,N_9716);
or U9775 (N_9775,N_9612,N_9701);
and U9776 (N_9776,N_9687,N_9634);
nand U9777 (N_9777,N_9527,N_9623);
or U9778 (N_9778,N_9501,N_9593);
or U9779 (N_9779,N_9531,N_9736);
nor U9780 (N_9780,N_9682,N_9544);
or U9781 (N_9781,N_9683,N_9654);
nor U9782 (N_9782,N_9703,N_9604);
nand U9783 (N_9783,N_9598,N_9690);
xnor U9784 (N_9784,N_9620,N_9558);
nor U9785 (N_9785,N_9606,N_9661);
xnor U9786 (N_9786,N_9607,N_9608);
xor U9787 (N_9787,N_9619,N_9637);
xnor U9788 (N_9788,N_9665,N_9656);
or U9789 (N_9789,N_9555,N_9722);
nand U9790 (N_9790,N_9573,N_9602);
nor U9791 (N_9791,N_9539,N_9705);
and U9792 (N_9792,N_9639,N_9650);
xor U9793 (N_9793,N_9713,N_9587);
nand U9794 (N_9794,N_9512,N_9541);
and U9795 (N_9795,N_9670,N_9644);
and U9796 (N_9796,N_9640,N_9621);
xnor U9797 (N_9797,N_9553,N_9746);
and U9798 (N_9798,N_9712,N_9718);
nor U9799 (N_9799,N_9708,N_9748);
xnor U9800 (N_9800,N_9658,N_9572);
nand U9801 (N_9801,N_9570,N_9669);
nor U9802 (N_9802,N_9614,N_9542);
and U9803 (N_9803,N_9633,N_9629);
and U9804 (N_9804,N_9592,N_9729);
nand U9805 (N_9805,N_9505,N_9589);
and U9806 (N_9806,N_9568,N_9529);
nand U9807 (N_9807,N_9625,N_9586);
xnor U9808 (N_9808,N_9595,N_9740);
or U9809 (N_9809,N_9659,N_9695);
xnor U9810 (N_9810,N_9627,N_9653);
nor U9811 (N_9811,N_9559,N_9524);
nor U9812 (N_9812,N_9651,N_9643);
and U9813 (N_9813,N_9534,N_9732);
xor U9814 (N_9814,N_9742,N_9578);
xnor U9815 (N_9815,N_9584,N_9517);
nand U9816 (N_9816,N_9731,N_9611);
nor U9817 (N_9817,N_9560,N_9506);
xor U9818 (N_9818,N_9679,N_9724);
xor U9819 (N_9819,N_9673,N_9557);
and U9820 (N_9820,N_9674,N_9515);
and U9821 (N_9821,N_9518,N_9630);
nor U9822 (N_9822,N_9615,N_9657);
nor U9823 (N_9823,N_9692,N_9538);
nor U9824 (N_9824,N_9710,N_9508);
and U9825 (N_9825,N_9564,N_9743);
or U9826 (N_9826,N_9576,N_9635);
xor U9827 (N_9827,N_9704,N_9719);
nor U9828 (N_9828,N_9678,N_9677);
nor U9829 (N_9829,N_9675,N_9543);
nand U9830 (N_9830,N_9645,N_9561);
and U9831 (N_9831,N_9648,N_9624);
xnor U9832 (N_9832,N_9551,N_9594);
xnor U9833 (N_9833,N_9652,N_9646);
nor U9834 (N_9834,N_9681,N_9596);
xor U9835 (N_9835,N_9744,N_9522);
and U9836 (N_9836,N_9734,N_9613);
nand U9837 (N_9837,N_9738,N_9642);
xnor U9838 (N_9838,N_9714,N_9671);
xor U9839 (N_9839,N_9579,N_9575);
or U9840 (N_9840,N_9730,N_9706);
and U9841 (N_9841,N_9727,N_9697);
nor U9842 (N_9842,N_9649,N_9537);
nor U9843 (N_9843,N_9536,N_9721);
xnor U9844 (N_9844,N_9510,N_9535);
or U9845 (N_9845,N_9638,N_9580);
nor U9846 (N_9846,N_9509,N_9530);
and U9847 (N_9847,N_9523,N_9622);
nor U9848 (N_9848,N_9667,N_9513);
nand U9849 (N_9849,N_9631,N_9526);
or U9850 (N_9850,N_9610,N_9514);
and U9851 (N_9851,N_9552,N_9567);
and U9852 (N_9852,N_9632,N_9588);
or U9853 (N_9853,N_9733,N_9715);
nor U9854 (N_9854,N_9699,N_9686);
xor U9855 (N_9855,N_9747,N_9597);
and U9856 (N_9856,N_9590,N_9672);
or U9857 (N_9857,N_9540,N_9741);
and U9858 (N_9858,N_9694,N_9726);
and U9859 (N_9859,N_9749,N_9737);
xor U9860 (N_9860,N_9521,N_9601);
xor U9861 (N_9861,N_9745,N_9603);
xnor U9862 (N_9862,N_9605,N_9599);
and U9863 (N_9863,N_9689,N_9688);
nand U9864 (N_9864,N_9663,N_9662);
xnor U9865 (N_9865,N_9717,N_9507);
and U9866 (N_9866,N_9647,N_9685);
and U9867 (N_9867,N_9582,N_9504);
nor U9868 (N_9868,N_9533,N_9641);
xor U9869 (N_9869,N_9547,N_9571);
and U9870 (N_9870,N_9618,N_9520);
xnor U9871 (N_9871,N_9502,N_9563);
or U9872 (N_9872,N_9562,N_9600);
xor U9873 (N_9873,N_9626,N_9546);
or U9874 (N_9874,N_9666,N_9581);
or U9875 (N_9875,N_9645,N_9619);
or U9876 (N_9876,N_9573,N_9700);
nand U9877 (N_9877,N_9529,N_9543);
xor U9878 (N_9878,N_9546,N_9550);
and U9879 (N_9879,N_9671,N_9517);
or U9880 (N_9880,N_9663,N_9706);
nand U9881 (N_9881,N_9691,N_9639);
and U9882 (N_9882,N_9673,N_9520);
and U9883 (N_9883,N_9661,N_9577);
xnor U9884 (N_9884,N_9644,N_9737);
and U9885 (N_9885,N_9582,N_9623);
or U9886 (N_9886,N_9577,N_9705);
or U9887 (N_9887,N_9505,N_9658);
nor U9888 (N_9888,N_9632,N_9569);
xor U9889 (N_9889,N_9530,N_9614);
or U9890 (N_9890,N_9503,N_9538);
nor U9891 (N_9891,N_9735,N_9566);
nor U9892 (N_9892,N_9511,N_9712);
nand U9893 (N_9893,N_9709,N_9700);
nand U9894 (N_9894,N_9568,N_9640);
and U9895 (N_9895,N_9714,N_9510);
or U9896 (N_9896,N_9592,N_9531);
or U9897 (N_9897,N_9600,N_9521);
or U9898 (N_9898,N_9537,N_9682);
nor U9899 (N_9899,N_9565,N_9678);
nand U9900 (N_9900,N_9583,N_9536);
nor U9901 (N_9901,N_9748,N_9520);
nor U9902 (N_9902,N_9517,N_9593);
or U9903 (N_9903,N_9509,N_9708);
or U9904 (N_9904,N_9672,N_9633);
or U9905 (N_9905,N_9698,N_9567);
nor U9906 (N_9906,N_9542,N_9507);
xor U9907 (N_9907,N_9625,N_9576);
nor U9908 (N_9908,N_9631,N_9627);
xnor U9909 (N_9909,N_9595,N_9745);
nor U9910 (N_9910,N_9720,N_9647);
nor U9911 (N_9911,N_9644,N_9716);
nor U9912 (N_9912,N_9635,N_9720);
xor U9913 (N_9913,N_9638,N_9589);
xor U9914 (N_9914,N_9725,N_9587);
xor U9915 (N_9915,N_9669,N_9691);
and U9916 (N_9916,N_9547,N_9720);
nand U9917 (N_9917,N_9606,N_9505);
nor U9918 (N_9918,N_9593,N_9743);
nor U9919 (N_9919,N_9611,N_9561);
and U9920 (N_9920,N_9674,N_9721);
nand U9921 (N_9921,N_9531,N_9684);
nor U9922 (N_9922,N_9694,N_9625);
or U9923 (N_9923,N_9747,N_9617);
and U9924 (N_9924,N_9575,N_9604);
or U9925 (N_9925,N_9534,N_9602);
or U9926 (N_9926,N_9643,N_9661);
nor U9927 (N_9927,N_9622,N_9510);
or U9928 (N_9928,N_9734,N_9676);
xnor U9929 (N_9929,N_9618,N_9661);
nor U9930 (N_9930,N_9626,N_9521);
or U9931 (N_9931,N_9649,N_9614);
and U9932 (N_9932,N_9599,N_9512);
xnor U9933 (N_9933,N_9691,N_9603);
xor U9934 (N_9934,N_9691,N_9734);
xor U9935 (N_9935,N_9562,N_9656);
and U9936 (N_9936,N_9651,N_9628);
xor U9937 (N_9937,N_9678,N_9537);
xnor U9938 (N_9938,N_9639,N_9685);
xnor U9939 (N_9939,N_9703,N_9670);
and U9940 (N_9940,N_9716,N_9642);
nand U9941 (N_9941,N_9741,N_9698);
and U9942 (N_9942,N_9714,N_9627);
nor U9943 (N_9943,N_9503,N_9665);
nor U9944 (N_9944,N_9679,N_9509);
xnor U9945 (N_9945,N_9558,N_9657);
nand U9946 (N_9946,N_9712,N_9716);
nor U9947 (N_9947,N_9615,N_9505);
xor U9948 (N_9948,N_9672,N_9660);
xor U9949 (N_9949,N_9728,N_9598);
nand U9950 (N_9950,N_9575,N_9576);
nand U9951 (N_9951,N_9551,N_9687);
and U9952 (N_9952,N_9605,N_9662);
nor U9953 (N_9953,N_9577,N_9671);
or U9954 (N_9954,N_9502,N_9738);
xor U9955 (N_9955,N_9611,N_9565);
nor U9956 (N_9956,N_9552,N_9594);
nand U9957 (N_9957,N_9554,N_9723);
nand U9958 (N_9958,N_9575,N_9562);
nand U9959 (N_9959,N_9585,N_9562);
xor U9960 (N_9960,N_9583,N_9743);
nor U9961 (N_9961,N_9602,N_9671);
xnor U9962 (N_9962,N_9547,N_9697);
nor U9963 (N_9963,N_9546,N_9588);
or U9964 (N_9964,N_9509,N_9711);
nor U9965 (N_9965,N_9719,N_9563);
nand U9966 (N_9966,N_9676,N_9706);
nor U9967 (N_9967,N_9696,N_9647);
and U9968 (N_9968,N_9614,N_9734);
nand U9969 (N_9969,N_9514,N_9650);
and U9970 (N_9970,N_9588,N_9706);
and U9971 (N_9971,N_9632,N_9694);
nor U9972 (N_9972,N_9582,N_9557);
xor U9973 (N_9973,N_9721,N_9611);
nand U9974 (N_9974,N_9552,N_9509);
nor U9975 (N_9975,N_9625,N_9628);
or U9976 (N_9976,N_9670,N_9647);
nor U9977 (N_9977,N_9688,N_9671);
and U9978 (N_9978,N_9749,N_9662);
and U9979 (N_9979,N_9579,N_9744);
and U9980 (N_9980,N_9743,N_9645);
xnor U9981 (N_9981,N_9563,N_9735);
nor U9982 (N_9982,N_9551,N_9643);
or U9983 (N_9983,N_9656,N_9680);
nor U9984 (N_9984,N_9696,N_9653);
nand U9985 (N_9985,N_9539,N_9562);
or U9986 (N_9986,N_9658,N_9581);
or U9987 (N_9987,N_9504,N_9651);
or U9988 (N_9988,N_9507,N_9512);
nand U9989 (N_9989,N_9717,N_9592);
nand U9990 (N_9990,N_9745,N_9726);
nor U9991 (N_9991,N_9569,N_9639);
nand U9992 (N_9992,N_9580,N_9599);
or U9993 (N_9993,N_9651,N_9699);
xnor U9994 (N_9994,N_9670,N_9574);
and U9995 (N_9995,N_9500,N_9690);
and U9996 (N_9996,N_9596,N_9629);
nand U9997 (N_9997,N_9651,N_9596);
xnor U9998 (N_9998,N_9638,N_9717);
and U9999 (N_9999,N_9573,N_9584);
xor U10000 (N_10000,N_9999,N_9851);
and U10001 (N_10001,N_9927,N_9998);
or U10002 (N_10002,N_9835,N_9936);
and U10003 (N_10003,N_9815,N_9890);
or U10004 (N_10004,N_9858,N_9801);
xnor U10005 (N_10005,N_9865,N_9882);
nand U10006 (N_10006,N_9840,N_9976);
xnor U10007 (N_10007,N_9797,N_9867);
or U10008 (N_10008,N_9947,N_9778);
xor U10009 (N_10009,N_9965,N_9839);
nor U10010 (N_10010,N_9769,N_9857);
nand U10011 (N_10011,N_9923,N_9770);
and U10012 (N_10012,N_9940,N_9949);
xor U10013 (N_10013,N_9938,N_9964);
or U10014 (N_10014,N_9791,N_9820);
nor U10015 (N_10015,N_9752,N_9806);
or U10016 (N_10016,N_9765,N_9846);
xor U10017 (N_10017,N_9974,N_9972);
or U10018 (N_10018,N_9982,N_9776);
nand U10019 (N_10019,N_9800,N_9945);
xnor U10020 (N_10020,N_9828,N_9783);
and U10021 (N_10021,N_9794,N_9971);
nand U10022 (N_10022,N_9967,N_9834);
or U10023 (N_10023,N_9939,N_9779);
xor U10024 (N_10024,N_9899,N_9888);
xnor U10025 (N_10025,N_9790,N_9956);
or U10026 (N_10026,N_9980,N_9841);
nor U10027 (N_10027,N_9991,N_9887);
or U10028 (N_10028,N_9996,N_9950);
or U10029 (N_10029,N_9754,N_9994);
and U10030 (N_10030,N_9788,N_9831);
and U10031 (N_10031,N_9863,N_9934);
or U10032 (N_10032,N_9781,N_9931);
nor U10033 (N_10033,N_9786,N_9925);
xnor U10034 (N_10034,N_9808,N_9817);
or U10035 (N_10035,N_9917,N_9914);
xor U10036 (N_10036,N_9963,N_9795);
nand U10037 (N_10037,N_9932,N_9966);
or U10038 (N_10038,N_9958,N_9906);
or U10039 (N_10039,N_9830,N_9916);
nor U10040 (N_10040,N_9983,N_9811);
and U10041 (N_10041,N_9870,N_9960);
and U10042 (N_10042,N_9751,N_9850);
nor U10043 (N_10043,N_9881,N_9922);
and U10044 (N_10044,N_9787,N_9774);
nor U10045 (N_10045,N_9969,N_9883);
and U10046 (N_10046,N_9866,N_9903);
nand U10047 (N_10047,N_9873,N_9951);
nor U10048 (N_10048,N_9847,N_9763);
nand U10049 (N_10049,N_9874,N_9809);
xnor U10050 (N_10050,N_9904,N_9911);
nor U10051 (N_10051,N_9973,N_9818);
and U10052 (N_10052,N_9871,N_9977);
xnor U10053 (N_10053,N_9886,N_9761);
nand U10054 (N_10054,N_9799,N_9946);
or U10055 (N_10055,N_9878,N_9884);
and U10056 (N_10056,N_9913,N_9880);
xnor U10057 (N_10057,N_9920,N_9937);
and U10058 (N_10058,N_9764,N_9756);
xor U10059 (N_10059,N_9814,N_9872);
xor U10060 (N_10060,N_9849,N_9829);
nor U10061 (N_10061,N_9985,N_9944);
nor U10062 (N_10062,N_9796,N_9803);
nand U10063 (N_10063,N_9784,N_9975);
nand U10064 (N_10064,N_9864,N_9984);
and U10065 (N_10065,N_9889,N_9861);
nor U10066 (N_10066,N_9848,N_9772);
and U10067 (N_10067,N_9869,N_9785);
nand U10068 (N_10068,N_9896,N_9876);
nand U10069 (N_10069,N_9968,N_9805);
or U10070 (N_10070,N_9804,N_9792);
nand U10071 (N_10071,N_9902,N_9935);
nand U10072 (N_10072,N_9877,N_9789);
xor U10073 (N_10073,N_9819,N_9928);
nor U10074 (N_10074,N_9900,N_9842);
and U10075 (N_10075,N_9995,N_9898);
nor U10076 (N_10076,N_9875,N_9997);
or U10077 (N_10077,N_9933,N_9986);
nor U10078 (N_10078,N_9859,N_9854);
nor U10079 (N_10079,N_9924,N_9868);
xor U10080 (N_10080,N_9862,N_9909);
and U10081 (N_10081,N_9897,N_9760);
and U10082 (N_10082,N_9827,N_9941);
nand U10083 (N_10083,N_9825,N_9894);
and U10084 (N_10084,N_9855,N_9821);
xor U10085 (N_10085,N_9879,N_9780);
xor U10086 (N_10086,N_9961,N_9978);
nor U10087 (N_10087,N_9942,N_9929);
or U10088 (N_10088,N_9930,N_9852);
or U10089 (N_10089,N_9838,N_9823);
or U10090 (N_10090,N_9832,N_9987);
or U10091 (N_10091,N_9775,N_9816);
or U10092 (N_10092,N_9836,N_9810);
nor U10093 (N_10093,N_9988,N_9766);
or U10094 (N_10094,N_9833,N_9990);
or U10095 (N_10095,N_9753,N_9755);
xor U10096 (N_10096,N_9989,N_9901);
xnor U10097 (N_10097,N_9767,N_9962);
nor U10098 (N_10098,N_9826,N_9912);
xor U10099 (N_10099,N_9822,N_9768);
xor U10100 (N_10100,N_9843,N_9954);
xnor U10101 (N_10101,N_9943,N_9802);
and U10102 (N_10102,N_9895,N_9948);
nor U10103 (N_10103,N_9771,N_9773);
or U10104 (N_10104,N_9905,N_9758);
nand U10105 (N_10105,N_9798,N_9926);
and U10106 (N_10106,N_9893,N_9921);
or U10107 (N_10107,N_9918,N_9782);
nand U10108 (N_10108,N_9981,N_9919);
nand U10109 (N_10109,N_9844,N_9907);
xnor U10110 (N_10110,N_9853,N_9750);
and U10111 (N_10111,N_9915,N_9955);
or U10112 (N_10112,N_9959,N_9957);
and U10113 (N_10113,N_9812,N_9953);
or U10114 (N_10114,N_9979,N_9793);
or U10115 (N_10115,N_9885,N_9845);
and U10116 (N_10116,N_9892,N_9813);
and U10117 (N_10117,N_9762,N_9993);
nor U10118 (N_10118,N_9908,N_9952);
nor U10119 (N_10119,N_9891,N_9910);
and U10120 (N_10120,N_9759,N_9777);
and U10121 (N_10121,N_9757,N_9992);
xnor U10122 (N_10122,N_9807,N_9970);
nor U10123 (N_10123,N_9860,N_9837);
xnor U10124 (N_10124,N_9856,N_9824);
and U10125 (N_10125,N_9810,N_9983);
or U10126 (N_10126,N_9875,N_9895);
or U10127 (N_10127,N_9807,N_9827);
and U10128 (N_10128,N_9879,N_9826);
nand U10129 (N_10129,N_9823,N_9800);
and U10130 (N_10130,N_9813,N_9817);
nand U10131 (N_10131,N_9891,N_9947);
nand U10132 (N_10132,N_9778,N_9764);
nand U10133 (N_10133,N_9787,N_9998);
nor U10134 (N_10134,N_9848,N_9983);
xor U10135 (N_10135,N_9893,N_9830);
and U10136 (N_10136,N_9951,N_9908);
and U10137 (N_10137,N_9977,N_9834);
and U10138 (N_10138,N_9837,N_9863);
or U10139 (N_10139,N_9864,N_9954);
or U10140 (N_10140,N_9852,N_9941);
xor U10141 (N_10141,N_9861,N_9892);
xnor U10142 (N_10142,N_9790,N_9785);
and U10143 (N_10143,N_9870,N_9815);
xnor U10144 (N_10144,N_9825,N_9990);
or U10145 (N_10145,N_9914,N_9994);
and U10146 (N_10146,N_9884,N_9969);
nor U10147 (N_10147,N_9876,N_9843);
and U10148 (N_10148,N_9757,N_9950);
nand U10149 (N_10149,N_9777,N_9807);
or U10150 (N_10150,N_9810,N_9822);
or U10151 (N_10151,N_9790,N_9837);
or U10152 (N_10152,N_9959,N_9912);
nand U10153 (N_10153,N_9845,N_9959);
and U10154 (N_10154,N_9796,N_9845);
and U10155 (N_10155,N_9775,N_9751);
nor U10156 (N_10156,N_9942,N_9891);
nor U10157 (N_10157,N_9940,N_9904);
or U10158 (N_10158,N_9973,N_9982);
nor U10159 (N_10159,N_9921,N_9920);
nor U10160 (N_10160,N_9953,N_9886);
and U10161 (N_10161,N_9845,N_9988);
and U10162 (N_10162,N_9907,N_9765);
nor U10163 (N_10163,N_9899,N_9986);
and U10164 (N_10164,N_9920,N_9924);
nand U10165 (N_10165,N_9862,N_9875);
nand U10166 (N_10166,N_9936,N_9862);
xnor U10167 (N_10167,N_9754,N_9959);
and U10168 (N_10168,N_9766,N_9905);
nand U10169 (N_10169,N_9890,N_9899);
or U10170 (N_10170,N_9855,N_9946);
and U10171 (N_10171,N_9844,N_9796);
and U10172 (N_10172,N_9988,N_9899);
nand U10173 (N_10173,N_9829,N_9809);
nand U10174 (N_10174,N_9948,N_9954);
and U10175 (N_10175,N_9947,N_9979);
xnor U10176 (N_10176,N_9835,N_9891);
xor U10177 (N_10177,N_9846,N_9931);
and U10178 (N_10178,N_9809,N_9758);
xor U10179 (N_10179,N_9951,N_9855);
xnor U10180 (N_10180,N_9807,N_9779);
nor U10181 (N_10181,N_9985,N_9975);
and U10182 (N_10182,N_9897,N_9992);
and U10183 (N_10183,N_9948,N_9759);
nand U10184 (N_10184,N_9921,N_9941);
nand U10185 (N_10185,N_9844,N_9877);
nand U10186 (N_10186,N_9835,N_9912);
xor U10187 (N_10187,N_9935,N_9816);
and U10188 (N_10188,N_9929,N_9907);
nand U10189 (N_10189,N_9828,N_9894);
nand U10190 (N_10190,N_9925,N_9775);
nand U10191 (N_10191,N_9947,N_9899);
xnor U10192 (N_10192,N_9777,N_9871);
xnor U10193 (N_10193,N_9936,N_9892);
nand U10194 (N_10194,N_9920,N_9999);
or U10195 (N_10195,N_9964,N_9941);
xor U10196 (N_10196,N_9953,N_9814);
and U10197 (N_10197,N_9771,N_9917);
or U10198 (N_10198,N_9854,N_9817);
or U10199 (N_10199,N_9852,N_9789);
nor U10200 (N_10200,N_9895,N_9904);
xnor U10201 (N_10201,N_9946,N_9798);
or U10202 (N_10202,N_9990,N_9792);
and U10203 (N_10203,N_9852,N_9843);
nor U10204 (N_10204,N_9846,N_9794);
nand U10205 (N_10205,N_9752,N_9820);
and U10206 (N_10206,N_9784,N_9889);
nor U10207 (N_10207,N_9871,N_9886);
xor U10208 (N_10208,N_9812,N_9838);
nor U10209 (N_10209,N_9949,N_9885);
or U10210 (N_10210,N_9974,N_9759);
or U10211 (N_10211,N_9974,N_9997);
and U10212 (N_10212,N_9838,N_9756);
or U10213 (N_10213,N_9886,N_9813);
xor U10214 (N_10214,N_9931,N_9917);
and U10215 (N_10215,N_9786,N_9965);
xnor U10216 (N_10216,N_9796,N_9822);
nand U10217 (N_10217,N_9884,N_9925);
and U10218 (N_10218,N_9774,N_9934);
and U10219 (N_10219,N_9792,N_9883);
or U10220 (N_10220,N_9893,N_9773);
and U10221 (N_10221,N_9912,N_9998);
xor U10222 (N_10222,N_9765,N_9824);
nand U10223 (N_10223,N_9813,N_9934);
nor U10224 (N_10224,N_9854,N_9820);
nand U10225 (N_10225,N_9783,N_9973);
nand U10226 (N_10226,N_9870,N_9980);
and U10227 (N_10227,N_9933,N_9750);
and U10228 (N_10228,N_9813,N_9842);
xor U10229 (N_10229,N_9965,N_9955);
or U10230 (N_10230,N_9938,N_9930);
or U10231 (N_10231,N_9941,N_9767);
or U10232 (N_10232,N_9854,N_9891);
and U10233 (N_10233,N_9963,N_9778);
and U10234 (N_10234,N_9894,N_9841);
xnor U10235 (N_10235,N_9967,N_9778);
and U10236 (N_10236,N_9876,N_9865);
nand U10237 (N_10237,N_9760,N_9804);
xor U10238 (N_10238,N_9812,N_9859);
xor U10239 (N_10239,N_9800,N_9896);
nand U10240 (N_10240,N_9868,N_9925);
xor U10241 (N_10241,N_9922,N_9937);
xnor U10242 (N_10242,N_9976,N_9933);
xnor U10243 (N_10243,N_9988,N_9791);
and U10244 (N_10244,N_9797,N_9851);
and U10245 (N_10245,N_9822,N_9839);
or U10246 (N_10246,N_9854,N_9809);
nor U10247 (N_10247,N_9791,N_9857);
xor U10248 (N_10248,N_9776,N_9983);
or U10249 (N_10249,N_9764,N_9769);
nand U10250 (N_10250,N_10073,N_10170);
nand U10251 (N_10251,N_10027,N_10030);
nand U10252 (N_10252,N_10057,N_10038);
and U10253 (N_10253,N_10037,N_10187);
xnor U10254 (N_10254,N_10160,N_10232);
nand U10255 (N_10255,N_10195,N_10031);
nand U10256 (N_10256,N_10017,N_10055);
and U10257 (N_10257,N_10196,N_10206);
or U10258 (N_10258,N_10229,N_10070);
or U10259 (N_10259,N_10148,N_10025);
xnor U10260 (N_10260,N_10165,N_10068);
xnor U10261 (N_10261,N_10035,N_10240);
nand U10262 (N_10262,N_10154,N_10210);
and U10263 (N_10263,N_10089,N_10194);
nor U10264 (N_10264,N_10023,N_10242);
nand U10265 (N_10265,N_10149,N_10136);
nor U10266 (N_10266,N_10081,N_10062);
nand U10267 (N_10267,N_10087,N_10107);
or U10268 (N_10268,N_10022,N_10029);
nand U10269 (N_10269,N_10238,N_10010);
and U10270 (N_10270,N_10076,N_10133);
or U10271 (N_10271,N_10114,N_10071);
or U10272 (N_10272,N_10175,N_10225);
xor U10273 (N_10273,N_10122,N_10197);
or U10274 (N_10274,N_10155,N_10167);
nand U10275 (N_10275,N_10101,N_10080);
nor U10276 (N_10276,N_10042,N_10044);
xor U10277 (N_10277,N_10047,N_10054);
nand U10278 (N_10278,N_10235,N_10069);
nor U10279 (N_10279,N_10040,N_10028);
nor U10280 (N_10280,N_10217,N_10103);
or U10281 (N_10281,N_10157,N_10230);
xnor U10282 (N_10282,N_10248,N_10173);
nand U10283 (N_10283,N_10199,N_10059);
and U10284 (N_10284,N_10058,N_10139);
or U10285 (N_10285,N_10088,N_10219);
and U10286 (N_10286,N_10056,N_10128);
nand U10287 (N_10287,N_10012,N_10140);
and U10288 (N_10288,N_10115,N_10245);
xor U10289 (N_10289,N_10168,N_10161);
and U10290 (N_10290,N_10223,N_10061);
nor U10291 (N_10291,N_10241,N_10186);
nor U10292 (N_10292,N_10145,N_10009);
or U10293 (N_10293,N_10171,N_10006);
xor U10294 (N_10294,N_10174,N_10201);
and U10295 (N_10295,N_10099,N_10033);
nand U10296 (N_10296,N_10226,N_10190);
nor U10297 (N_10297,N_10202,N_10118);
nor U10298 (N_10298,N_10112,N_10207);
and U10299 (N_10299,N_10185,N_10036);
or U10300 (N_10300,N_10224,N_10067);
nand U10301 (N_10301,N_10002,N_10172);
or U10302 (N_10302,N_10008,N_10125);
nand U10303 (N_10303,N_10153,N_10105);
nor U10304 (N_10304,N_10227,N_10192);
xnor U10305 (N_10305,N_10050,N_10146);
and U10306 (N_10306,N_10138,N_10191);
nor U10307 (N_10307,N_10106,N_10234);
nand U10308 (N_10308,N_10060,N_10176);
nand U10309 (N_10309,N_10066,N_10082);
nand U10310 (N_10310,N_10046,N_10213);
xor U10311 (N_10311,N_10152,N_10090);
nor U10312 (N_10312,N_10221,N_10239);
nor U10313 (N_10313,N_10236,N_10130);
nor U10314 (N_10314,N_10193,N_10043);
xnor U10315 (N_10315,N_10109,N_10228);
xor U10316 (N_10316,N_10034,N_10003);
nand U10317 (N_10317,N_10124,N_10074);
nand U10318 (N_10318,N_10120,N_10024);
and U10319 (N_10319,N_10110,N_10156);
nand U10320 (N_10320,N_10158,N_10117);
xnor U10321 (N_10321,N_10222,N_10189);
xor U10322 (N_10322,N_10032,N_10111);
nor U10323 (N_10323,N_10097,N_10249);
or U10324 (N_10324,N_10121,N_10244);
or U10325 (N_10325,N_10007,N_10164);
nand U10326 (N_10326,N_10209,N_10095);
xnor U10327 (N_10327,N_10092,N_10104);
nand U10328 (N_10328,N_10123,N_10093);
or U10329 (N_10329,N_10216,N_10065);
and U10330 (N_10330,N_10231,N_10212);
nor U10331 (N_10331,N_10119,N_10000);
and U10332 (N_10332,N_10078,N_10247);
or U10333 (N_10333,N_10098,N_10075);
nor U10334 (N_10334,N_10014,N_10091);
xnor U10335 (N_10335,N_10184,N_10051);
and U10336 (N_10336,N_10214,N_10143);
nor U10337 (N_10337,N_10048,N_10147);
nor U10338 (N_10338,N_10063,N_10129);
and U10339 (N_10339,N_10188,N_10085);
or U10340 (N_10340,N_10001,N_10026);
nor U10341 (N_10341,N_10144,N_10141);
nor U10342 (N_10342,N_10243,N_10108);
or U10343 (N_10343,N_10159,N_10049);
nor U10344 (N_10344,N_10134,N_10021);
xor U10345 (N_10345,N_10211,N_10178);
or U10346 (N_10346,N_10094,N_10041);
and U10347 (N_10347,N_10198,N_10131);
or U10348 (N_10348,N_10116,N_10218);
xnor U10349 (N_10349,N_10150,N_10039);
xor U10350 (N_10350,N_10163,N_10020);
nand U10351 (N_10351,N_10132,N_10127);
and U10352 (N_10352,N_10233,N_10100);
or U10353 (N_10353,N_10246,N_10204);
or U10354 (N_10354,N_10019,N_10181);
and U10355 (N_10355,N_10169,N_10177);
and U10356 (N_10356,N_10166,N_10086);
nor U10357 (N_10357,N_10052,N_10079);
or U10358 (N_10358,N_10179,N_10018);
or U10359 (N_10359,N_10162,N_10013);
xnor U10360 (N_10360,N_10203,N_10016);
or U10361 (N_10361,N_10237,N_10053);
xnor U10362 (N_10362,N_10182,N_10215);
and U10363 (N_10363,N_10220,N_10137);
nor U10364 (N_10364,N_10004,N_10151);
and U10365 (N_10365,N_10142,N_10083);
nand U10366 (N_10366,N_10113,N_10045);
or U10367 (N_10367,N_10096,N_10015);
nor U10368 (N_10368,N_10064,N_10180);
nand U10369 (N_10369,N_10135,N_10126);
or U10370 (N_10370,N_10102,N_10077);
or U10371 (N_10371,N_10205,N_10200);
or U10372 (N_10372,N_10011,N_10208);
xor U10373 (N_10373,N_10005,N_10072);
nand U10374 (N_10374,N_10183,N_10084);
nor U10375 (N_10375,N_10100,N_10077);
nor U10376 (N_10376,N_10118,N_10138);
nand U10377 (N_10377,N_10167,N_10242);
and U10378 (N_10378,N_10002,N_10213);
and U10379 (N_10379,N_10159,N_10075);
xor U10380 (N_10380,N_10077,N_10063);
and U10381 (N_10381,N_10187,N_10004);
xor U10382 (N_10382,N_10124,N_10226);
and U10383 (N_10383,N_10023,N_10064);
xnor U10384 (N_10384,N_10181,N_10011);
nor U10385 (N_10385,N_10042,N_10153);
or U10386 (N_10386,N_10235,N_10105);
nor U10387 (N_10387,N_10241,N_10074);
or U10388 (N_10388,N_10132,N_10138);
xnor U10389 (N_10389,N_10001,N_10013);
and U10390 (N_10390,N_10070,N_10163);
and U10391 (N_10391,N_10024,N_10040);
nor U10392 (N_10392,N_10208,N_10088);
xnor U10393 (N_10393,N_10028,N_10091);
nand U10394 (N_10394,N_10123,N_10217);
nor U10395 (N_10395,N_10092,N_10111);
nor U10396 (N_10396,N_10200,N_10108);
or U10397 (N_10397,N_10179,N_10148);
nor U10398 (N_10398,N_10086,N_10026);
nand U10399 (N_10399,N_10180,N_10161);
or U10400 (N_10400,N_10085,N_10082);
or U10401 (N_10401,N_10228,N_10076);
and U10402 (N_10402,N_10180,N_10098);
nor U10403 (N_10403,N_10015,N_10212);
nor U10404 (N_10404,N_10094,N_10116);
and U10405 (N_10405,N_10225,N_10150);
or U10406 (N_10406,N_10106,N_10133);
nand U10407 (N_10407,N_10188,N_10053);
nor U10408 (N_10408,N_10014,N_10128);
nand U10409 (N_10409,N_10061,N_10173);
and U10410 (N_10410,N_10046,N_10058);
nor U10411 (N_10411,N_10029,N_10210);
nor U10412 (N_10412,N_10162,N_10052);
xnor U10413 (N_10413,N_10100,N_10112);
or U10414 (N_10414,N_10182,N_10026);
nand U10415 (N_10415,N_10098,N_10088);
and U10416 (N_10416,N_10212,N_10233);
nand U10417 (N_10417,N_10010,N_10000);
and U10418 (N_10418,N_10129,N_10033);
nor U10419 (N_10419,N_10220,N_10035);
and U10420 (N_10420,N_10004,N_10144);
nand U10421 (N_10421,N_10162,N_10007);
or U10422 (N_10422,N_10089,N_10039);
and U10423 (N_10423,N_10095,N_10121);
and U10424 (N_10424,N_10112,N_10070);
or U10425 (N_10425,N_10152,N_10037);
nand U10426 (N_10426,N_10168,N_10160);
or U10427 (N_10427,N_10220,N_10163);
and U10428 (N_10428,N_10198,N_10027);
nand U10429 (N_10429,N_10083,N_10192);
nor U10430 (N_10430,N_10014,N_10064);
nor U10431 (N_10431,N_10188,N_10044);
xor U10432 (N_10432,N_10090,N_10164);
nand U10433 (N_10433,N_10038,N_10035);
xnor U10434 (N_10434,N_10112,N_10176);
nand U10435 (N_10435,N_10163,N_10138);
nand U10436 (N_10436,N_10235,N_10025);
nor U10437 (N_10437,N_10137,N_10112);
nand U10438 (N_10438,N_10224,N_10159);
or U10439 (N_10439,N_10028,N_10012);
and U10440 (N_10440,N_10040,N_10091);
and U10441 (N_10441,N_10068,N_10124);
xor U10442 (N_10442,N_10233,N_10025);
or U10443 (N_10443,N_10128,N_10181);
xor U10444 (N_10444,N_10164,N_10202);
nor U10445 (N_10445,N_10156,N_10000);
xor U10446 (N_10446,N_10226,N_10089);
nand U10447 (N_10447,N_10151,N_10187);
xor U10448 (N_10448,N_10231,N_10016);
and U10449 (N_10449,N_10236,N_10197);
nor U10450 (N_10450,N_10173,N_10106);
xnor U10451 (N_10451,N_10161,N_10203);
nand U10452 (N_10452,N_10078,N_10191);
xnor U10453 (N_10453,N_10215,N_10211);
nand U10454 (N_10454,N_10054,N_10189);
nand U10455 (N_10455,N_10175,N_10186);
nor U10456 (N_10456,N_10106,N_10166);
or U10457 (N_10457,N_10065,N_10057);
nand U10458 (N_10458,N_10014,N_10132);
or U10459 (N_10459,N_10068,N_10001);
nor U10460 (N_10460,N_10133,N_10249);
xnor U10461 (N_10461,N_10167,N_10190);
nor U10462 (N_10462,N_10015,N_10225);
and U10463 (N_10463,N_10165,N_10027);
xor U10464 (N_10464,N_10029,N_10053);
nor U10465 (N_10465,N_10011,N_10241);
nor U10466 (N_10466,N_10033,N_10017);
or U10467 (N_10467,N_10159,N_10127);
nor U10468 (N_10468,N_10010,N_10063);
nor U10469 (N_10469,N_10046,N_10012);
xor U10470 (N_10470,N_10190,N_10180);
nor U10471 (N_10471,N_10099,N_10140);
xor U10472 (N_10472,N_10126,N_10023);
nand U10473 (N_10473,N_10120,N_10055);
nor U10474 (N_10474,N_10117,N_10032);
nor U10475 (N_10475,N_10043,N_10111);
nand U10476 (N_10476,N_10238,N_10191);
nor U10477 (N_10477,N_10096,N_10200);
nand U10478 (N_10478,N_10193,N_10191);
xor U10479 (N_10479,N_10096,N_10073);
xor U10480 (N_10480,N_10013,N_10156);
nand U10481 (N_10481,N_10204,N_10236);
nand U10482 (N_10482,N_10221,N_10110);
or U10483 (N_10483,N_10042,N_10036);
xor U10484 (N_10484,N_10139,N_10019);
nand U10485 (N_10485,N_10229,N_10017);
nand U10486 (N_10486,N_10151,N_10198);
nor U10487 (N_10487,N_10078,N_10050);
or U10488 (N_10488,N_10180,N_10077);
and U10489 (N_10489,N_10003,N_10138);
nand U10490 (N_10490,N_10097,N_10098);
xor U10491 (N_10491,N_10246,N_10016);
and U10492 (N_10492,N_10149,N_10148);
nand U10493 (N_10493,N_10152,N_10246);
nor U10494 (N_10494,N_10130,N_10062);
and U10495 (N_10495,N_10196,N_10082);
and U10496 (N_10496,N_10145,N_10167);
or U10497 (N_10497,N_10118,N_10167);
xor U10498 (N_10498,N_10178,N_10075);
nand U10499 (N_10499,N_10160,N_10060);
nand U10500 (N_10500,N_10319,N_10432);
nand U10501 (N_10501,N_10488,N_10364);
xnor U10502 (N_10502,N_10478,N_10369);
and U10503 (N_10503,N_10406,N_10339);
nor U10504 (N_10504,N_10288,N_10382);
and U10505 (N_10505,N_10380,N_10291);
xnor U10506 (N_10506,N_10343,N_10308);
nor U10507 (N_10507,N_10332,N_10395);
or U10508 (N_10508,N_10304,N_10321);
xor U10509 (N_10509,N_10257,N_10347);
or U10510 (N_10510,N_10450,N_10462);
or U10511 (N_10511,N_10325,N_10378);
and U10512 (N_10512,N_10385,N_10476);
and U10513 (N_10513,N_10441,N_10336);
nor U10514 (N_10514,N_10465,N_10252);
or U10515 (N_10515,N_10295,N_10368);
or U10516 (N_10516,N_10397,N_10425);
or U10517 (N_10517,N_10393,N_10453);
nand U10518 (N_10518,N_10373,N_10389);
or U10519 (N_10519,N_10307,N_10250);
xor U10520 (N_10520,N_10322,N_10413);
nand U10521 (N_10521,N_10418,N_10290);
or U10522 (N_10522,N_10374,N_10312);
or U10523 (N_10523,N_10455,N_10485);
nor U10524 (N_10524,N_10261,N_10314);
nor U10525 (N_10525,N_10417,N_10375);
xor U10526 (N_10526,N_10386,N_10349);
and U10527 (N_10527,N_10464,N_10411);
and U10528 (N_10528,N_10387,N_10297);
or U10529 (N_10529,N_10487,N_10424);
and U10530 (N_10530,N_10354,N_10344);
nor U10531 (N_10531,N_10470,N_10443);
xor U10532 (N_10532,N_10444,N_10495);
and U10533 (N_10533,N_10461,N_10340);
and U10534 (N_10534,N_10468,N_10469);
and U10535 (N_10535,N_10271,N_10281);
and U10536 (N_10536,N_10253,N_10346);
nor U10537 (N_10537,N_10458,N_10403);
xnor U10538 (N_10538,N_10482,N_10262);
nor U10539 (N_10539,N_10471,N_10440);
nand U10540 (N_10540,N_10463,N_10422);
or U10541 (N_10541,N_10416,N_10258);
or U10542 (N_10542,N_10268,N_10392);
xnor U10543 (N_10543,N_10251,N_10326);
or U10544 (N_10544,N_10284,N_10279);
and U10545 (N_10545,N_10313,N_10309);
or U10546 (N_10546,N_10415,N_10427);
xor U10547 (N_10547,N_10371,N_10356);
nor U10548 (N_10548,N_10435,N_10494);
or U10549 (N_10549,N_10280,N_10256);
nor U10550 (N_10550,N_10289,N_10275);
or U10551 (N_10551,N_10330,N_10341);
xnor U10552 (N_10552,N_10328,N_10466);
or U10553 (N_10553,N_10404,N_10434);
or U10554 (N_10554,N_10484,N_10260);
nor U10555 (N_10555,N_10263,N_10316);
xor U10556 (N_10556,N_10398,N_10334);
or U10557 (N_10557,N_10451,N_10351);
xor U10558 (N_10558,N_10269,N_10302);
xnor U10559 (N_10559,N_10423,N_10318);
nand U10560 (N_10560,N_10492,N_10479);
and U10561 (N_10561,N_10409,N_10480);
or U10562 (N_10562,N_10396,N_10446);
and U10563 (N_10563,N_10301,N_10477);
and U10564 (N_10564,N_10363,N_10298);
nand U10565 (N_10565,N_10359,N_10272);
or U10566 (N_10566,N_10498,N_10412);
nor U10567 (N_10567,N_10433,N_10442);
nor U10568 (N_10568,N_10497,N_10282);
or U10569 (N_10569,N_10456,N_10419);
nand U10570 (N_10570,N_10445,N_10345);
or U10571 (N_10571,N_10474,N_10329);
and U10572 (N_10572,N_10278,N_10283);
xor U10573 (N_10573,N_10327,N_10454);
nor U10574 (N_10574,N_10266,N_10473);
and U10575 (N_10575,N_10491,N_10431);
xnor U10576 (N_10576,N_10254,N_10310);
nand U10577 (N_10577,N_10475,N_10360);
and U10578 (N_10578,N_10277,N_10390);
nand U10579 (N_10579,N_10358,N_10361);
nand U10580 (N_10580,N_10276,N_10315);
nor U10581 (N_10581,N_10439,N_10426);
nand U10582 (N_10582,N_10366,N_10255);
or U10583 (N_10583,N_10401,N_10459);
nand U10584 (N_10584,N_10481,N_10273);
xnor U10585 (N_10585,N_10323,N_10384);
nand U10586 (N_10586,N_10264,N_10259);
nor U10587 (N_10587,N_10337,N_10400);
and U10588 (N_10588,N_10320,N_10324);
xor U10589 (N_10589,N_10306,N_10429);
and U10590 (N_10590,N_10483,N_10338);
or U10591 (N_10591,N_10287,N_10499);
nor U10592 (N_10592,N_10350,N_10388);
or U10593 (N_10593,N_10299,N_10420);
or U10594 (N_10594,N_10407,N_10293);
nor U10595 (N_10595,N_10342,N_10383);
nor U10596 (N_10596,N_10355,N_10300);
and U10597 (N_10597,N_10452,N_10496);
and U10598 (N_10598,N_10405,N_10489);
or U10599 (N_10599,N_10394,N_10448);
nor U10600 (N_10600,N_10486,N_10437);
nor U10601 (N_10601,N_10331,N_10376);
nor U10602 (N_10602,N_10305,N_10317);
and U10603 (N_10603,N_10377,N_10274);
and U10604 (N_10604,N_10438,N_10367);
nor U10605 (N_10605,N_10493,N_10414);
nand U10606 (N_10606,N_10381,N_10399);
xor U10607 (N_10607,N_10391,N_10410);
xnor U10608 (N_10608,N_10370,N_10365);
nand U10609 (N_10609,N_10285,N_10335);
nor U10610 (N_10610,N_10379,N_10472);
or U10611 (N_10611,N_10436,N_10408);
xor U10612 (N_10612,N_10303,N_10294);
and U10613 (N_10613,N_10348,N_10267);
or U10614 (N_10614,N_10490,N_10286);
nand U10615 (N_10615,N_10292,N_10333);
nand U10616 (N_10616,N_10362,N_10430);
and U10617 (N_10617,N_10372,N_10402);
nand U10618 (N_10618,N_10460,N_10421);
nor U10619 (N_10619,N_10447,N_10352);
and U10620 (N_10620,N_10296,N_10265);
xnor U10621 (N_10621,N_10270,N_10467);
and U10622 (N_10622,N_10449,N_10457);
nand U10623 (N_10623,N_10353,N_10311);
xnor U10624 (N_10624,N_10428,N_10357);
and U10625 (N_10625,N_10404,N_10300);
and U10626 (N_10626,N_10374,N_10418);
nor U10627 (N_10627,N_10478,N_10357);
nor U10628 (N_10628,N_10499,N_10471);
xor U10629 (N_10629,N_10322,N_10261);
and U10630 (N_10630,N_10409,N_10465);
and U10631 (N_10631,N_10323,N_10348);
and U10632 (N_10632,N_10340,N_10470);
nor U10633 (N_10633,N_10380,N_10494);
nand U10634 (N_10634,N_10435,N_10356);
xnor U10635 (N_10635,N_10382,N_10291);
or U10636 (N_10636,N_10344,N_10308);
nand U10637 (N_10637,N_10460,N_10496);
and U10638 (N_10638,N_10261,N_10273);
xnor U10639 (N_10639,N_10343,N_10280);
nor U10640 (N_10640,N_10286,N_10297);
nor U10641 (N_10641,N_10467,N_10381);
nand U10642 (N_10642,N_10468,N_10395);
or U10643 (N_10643,N_10401,N_10383);
nor U10644 (N_10644,N_10441,N_10415);
xnor U10645 (N_10645,N_10449,N_10280);
and U10646 (N_10646,N_10404,N_10426);
and U10647 (N_10647,N_10399,N_10435);
and U10648 (N_10648,N_10432,N_10370);
nand U10649 (N_10649,N_10364,N_10433);
or U10650 (N_10650,N_10393,N_10325);
and U10651 (N_10651,N_10350,N_10439);
and U10652 (N_10652,N_10289,N_10301);
or U10653 (N_10653,N_10279,N_10326);
or U10654 (N_10654,N_10458,N_10398);
nor U10655 (N_10655,N_10336,N_10288);
nand U10656 (N_10656,N_10258,N_10479);
nor U10657 (N_10657,N_10481,N_10277);
nor U10658 (N_10658,N_10318,N_10267);
or U10659 (N_10659,N_10377,N_10416);
and U10660 (N_10660,N_10494,N_10330);
nand U10661 (N_10661,N_10323,N_10431);
nor U10662 (N_10662,N_10481,N_10423);
nand U10663 (N_10663,N_10407,N_10343);
nor U10664 (N_10664,N_10477,N_10311);
nand U10665 (N_10665,N_10367,N_10355);
or U10666 (N_10666,N_10401,N_10497);
or U10667 (N_10667,N_10307,N_10259);
nor U10668 (N_10668,N_10288,N_10322);
xor U10669 (N_10669,N_10325,N_10430);
xnor U10670 (N_10670,N_10412,N_10317);
xnor U10671 (N_10671,N_10318,N_10350);
xor U10672 (N_10672,N_10411,N_10461);
and U10673 (N_10673,N_10497,N_10418);
or U10674 (N_10674,N_10408,N_10472);
or U10675 (N_10675,N_10438,N_10427);
nor U10676 (N_10676,N_10281,N_10357);
or U10677 (N_10677,N_10309,N_10365);
nand U10678 (N_10678,N_10269,N_10274);
or U10679 (N_10679,N_10274,N_10323);
nor U10680 (N_10680,N_10303,N_10319);
nor U10681 (N_10681,N_10315,N_10484);
nand U10682 (N_10682,N_10308,N_10268);
and U10683 (N_10683,N_10284,N_10318);
or U10684 (N_10684,N_10303,N_10349);
or U10685 (N_10685,N_10373,N_10474);
nor U10686 (N_10686,N_10396,N_10294);
and U10687 (N_10687,N_10258,N_10376);
xnor U10688 (N_10688,N_10412,N_10301);
xnor U10689 (N_10689,N_10304,N_10319);
nand U10690 (N_10690,N_10295,N_10436);
or U10691 (N_10691,N_10366,N_10380);
and U10692 (N_10692,N_10380,N_10460);
nor U10693 (N_10693,N_10319,N_10361);
xnor U10694 (N_10694,N_10424,N_10480);
nor U10695 (N_10695,N_10388,N_10405);
and U10696 (N_10696,N_10429,N_10463);
xor U10697 (N_10697,N_10410,N_10327);
or U10698 (N_10698,N_10290,N_10270);
or U10699 (N_10699,N_10252,N_10317);
or U10700 (N_10700,N_10438,N_10259);
or U10701 (N_10701,N_10266,N_10496);
xor U10702 (N_10702,N_10347,N_10282);
nor U10703 (N_10703,N_10283,N_10487);
nor U10704 (N_10704,N_10394,N_10341);
xnor U10705 (N_10705,N_10480,N_10333);
nor U10706 (N_10706,N_10487,N_10346);
or U10707 (N_10707,N_10488,N_10370);
and U10708 (N_10708,N_10343,N_10422);
xor U10709 (N_10709,N_10332,N_10313);
nand U10710 (N_10710,N_10338,N_10474);
and U10711 (N_10711,N_10297,N_10276);
or U10712 (N_10712,N_10311,N_10296);
or U10713 (N_10713,N_10308,N_10262);
or U10714 (N_10714,N_10329,N_10309);
xor U10715 (N_10715,N_10342,N_10337);
and U10716 (N_10716,N_10417,N_10478);
or U10717 (N_10717,N_10414,N_10352);
and U10718 (N_10718,N_10299,N_10423);
nor U10719 (N_10719,N_10334,N_10343);
or U10720 (N_10720,N_10369,N_10468);
and U10721 (N_10721,N_10399,N_10456);
nor U10722 (N_10722,N_10330,N_10323);
nand U10723 (N_10723,N_10451,N_10332);
and U10724 (N_10724,N_10369,N_10281);
and U10725 (N_10725,N_10347,N_10444);
xnor U10726 (N_10726,N_10302,N_10270);
or U10727 (N_10727,N_10453,N_10492);
xnor U10728 (N_10728,N_10324,N_10379);
xor U10729 (N_10729,N_10263,N_10370);
and U10730 (N_10730,N_10426,N_10479);
nor U10731 (N_10731,N_10475,N_10271);
nor U10732 (N_10732,N_10342,N_10468);
nor U10733 (N_10733,N_10286,N_10443);
or U10734 (N_10734,N_10450,N_10291);
and U10735 (N_10735,N_10430,N_10322);
xnor U10736 (N_10736,N_10426,N_10284);
nor U10737 (N_10737,N_10476,N_10293);
nor U10738 (N_10738,N_10376,N_10291);
nor U10739 (N_10739,N_10433,N_10497);
nand U10740 (N_10740,N_10490,N_10385);
and U10741 (N_10741,N_10314,N_10386);
nand U10742 (N_10742,N_10300,N_10382);
nand U10743 (N_10743,N_10259,N_10448);
nand U10744 (N_10744,N_10280,N_10329);
or U10745 (N_10745,N_10495,N_10443);
and U10746 (N_10746,N_10487,N_10320);
xnor U10747 (N_10747,N_10412,N_10367);
or U10748 (N_10748,N_10423,N_10344);
and U10749 (N_10749,N_10279,N_10407);
and U10750 (N_10750,N_10518,N_10675);
or U10751 (N_10751,N_10521,N_10619);
or U10752 (N_10752,N_10536,N_10592);
or U10753 (N_10753,N_10505,N_10574);
and U10754 (N_10754,N_10603,N_10708);
or U10755 (N_10755,N_10690,N_10534);
nand U10756 (N_10756,N_10511,N_10640);
nand U10757 (N_10757,N_10652,N_10528);
nor U10758 (N_10758,N_10571,N_10590);
and U10759 (N_10759,N_10720,N_10577);
nor U10760 (N_10760,N_10558,N_10566);
nand U10761 (N_10761,N_10655,N_10627);
and U10762 (N_10762,N_10615,N_10587);
nand U10763 (N_10763,N_10588,N_10682);
nand U10764 (N_10764,N_10656,N_10556);
xnor U10765 (N_10765,N_10572,N_10614);
nor U10766 (N_10766,N_10749,N_10582);
nand U10767 (N_10767,N_10677,N_10743);
nor U10768 (N_10768,N_10705,N_10621);
xnor U10769 (N_10769,N_10633,N_10601);
and U10770 (N_10770,N_10537,N_10514);
nor U10771 (N_10771,N_10669,N_10575);
xnor U10772 (N_10772,N_10699,N_10706);
nor U10773 (N_10773,N_10728,N_10579);
and U10774 (N_10774,N_10568,N_10507);
and U10775 (N_10775,N_10618,N_10695);
xnor U10776 (N_10776,N_10628,N_10508);
xnor U10777 (N_10777,N_10606,N_10596);
xor U10778 (N_10778,N_10671,N_10510);
xnor U10779 (N_10779,N_10548,N_10676);
and U10780 (N_10780,N_10702,N_10551);
nor U10781 (N_10781,N_10529,N_10597);
xnor U10782 (N_10782,N_10721,N_10623);
and U10783 (N_10783,N_10612,N_10535);
nand U10784 (N_10784,N_10522,N_10745);
xnor U10785 (N_10785,N_10586,N_10642);
xnor U10786 (N_10786,N_10666,N_10608);
and U10787 (N_10787,N_10722,N_10650);
or U10788 (N_10788,N_10717,N_10555);
nand U10789 (N_10789,N_10629,N_10746);
xor U10790 (N_10790,N_10600,N_10689);
xor U10791 (N_10791,N_10658,N_10573);
or U10792 (N_10792,N_10502,N_10515);
xnor U10793 (N_10793,N_10709,N_10638);
or U10794 (N_10794,N_10554,N_10646);
or U10795 (N_10795,N_10530,N_10704);
or U10796 (N_10796,N_10703,N_10609);
and U10797 (N_10797,N_10680,N_10517);
or U10798 (N_10798,N_10581,N_10565);
and U10799 (N_10799,N_10739,N_10538);
and U10800 (N_10800,N_10509,N_10580);
xor U10801 (N_10801,N_10578,N_10672);
or U10802 (N_10802,N_10700,N_10712);
or U10803 (N_10803,N_10540,N_10527);
xnor U10804 (N_10804,N_10732,N_10595);
nor U10805 (N_10805,N_10747,N_10694);
xor U10806 (N_10806,N_10649,N_10626);
and U10807 (N_10807,N_10737,N_10696);
xor U10808 (N_10808,N_10543,N_10516);
nand U10809 (N_10809,N_10567,N_10625);
or U10810 (N_10810,N_10735,N_10532);
or U10811 (N_10811,N_10667,N_10691);
and U10812 (N_10812,N_10500,N_10563);
and U10813 (N_10813,N_10635,N_10594);
nand U10814 (N_10814,N_10653,N_10674);
nand U10815 (N_10815,N_10512,N_10657);
nand U10816 (N_10816,N_10659,N_10553);
or U10817 (N_10817,N_10673,N_10645);
and U10818 (N_10818,N_10665,N_10726);
or U10819 (N_10819,N_10651,N_10670);
and U10820 (N_10820,N_10539,N_10531);
nand U10821 (N_10821,N_10549,N_10620);
xnor U10822 (N_10822,N_10501,N_10533);
nand U10823 (N_10823,N_10641,N_10622);
xnor U10824 (N_10824,N_10683,N_10724);
nand U10825 (N_10825,N_10541,N_10607);
nand U10826 (N_10826,N_10545,N_10599);
and U10827 (N_10827,N_10589,N_10688);
or U10828 (N_10828,N_10678,N_10668);
and U10829 (N_10829,N_10525,N_10637);
nor U10830 (N_10830,N_10584,N_10741);
or U10831 (N_10831,N_10585,N_10730);
or U10832 (N_10832,N_10593,N_10583);
xor U10833 (N_10833,N_10523,N_10685);
and U10834 (N_10834,N_10616,N_10701);
xor U10835 (N_10835,N_10632,N_10644);
or U10836 (N_10836,N_10624,N_10698);
or U10837 (N_10837,N_10604,N_10570);
or U10838 (N_10838,N_10617,N_10552);
nor U10839 (N_10839,N_10569,N_10647);
or U10840 (N_10840,N_10719,N_10727);
nor U10841 (N_10841,N_10550,N_10547);
nor U10842 (N_10842,N_10524,N_10631);
or U10843 (N_10843,N_10714,N_10664);
nand U10844 (N_10844,N_10713,N_10546);
nand U10845 (N_10845,N_10611,N_10602);
xnor U10846 (N_10846,N_10733,N_10562);
nand U10847 (N_10847,N_10520,N_10687);
nand U10848 (N_10848,N_10679,N_10725);
xor U10849 (N_10849,N_10513,N_10723);
nor U10850 (N_10850,N_10636,N_10729);
nand U10851 (N_10851,N_10734,N_10634);
and U10852 (N_10852,N_10564,N_10748);
or U10853 (N_10853,N_10503,N_10557);
xor U10854 (N_10854,N_10648,N_10718);
or U10855 (N_10855,N_10693,N_10710);
or U10856 (N_10856,N_10716,N_10610);
and U10857 (N_10857,N_10506,N_10526);
nand U10858 (N_10858,N_10559,N_10661);
or U10859 (N_10859,N_10639,N_10707);
nor U10860 (N_10860,N_10663,N_10542);
and U10861 (N_10861,N_10740,N_10598);
xnor U10862 (N_10862,N_10662,N_10686);
xor U10863 (N_10863,N_10519,N_10561);
xor U10864 (N_10864,N_10660,N_10697);
xor U10865 (N_10865,N_10613,N_10692);
nor U10866 (N_10866,N_10742,N_10715);
nand U10867 (N_10867,N_10544,N_10643);
nor U10868 (N_10868,N_10684,N_10731);
nor U10869 (N_10869,N_10744,N_10654);
or U10870 (N_10870,N_10630,N_10591);
nand U10871 (N_10871,N_10711,N_10738);
xor U10872 (N_10872,N_10504,N_10681);
nand U10873 (N_10873,N_10736,N_10560);
or U10874 (N_10874,N_10605,N_10576);
and U10875 (N_10875,N_10644,N_10724);
xor U10876 (N_10876,N_10718,N_10688);
nand U10877 (N_10877,N_10618,N_10579);
xnor U10878 (N_10878,N_10542,N_10693);
xnor U10879 (N_10879,N_10743,N_10557);
xor U10880 (N_10880,N_10511,N_10567);
xnor U10881 (N_10881,N_10724,N_10657);
xnor U10882 (N_10882,N_10656,N_10563);
and U10883 (N_10883,N_10725,N_10594);
nand U10884 (N_10884,N_10659,N_10537);
nand U10885 (N_10885,N_10562,N_10731);
and U10886 (N_10886,N_10718,N_10581);
nand U10887 (N_10887,N_10709,N_10697);
xnor U10888 (N_10888,N_10570,N_10550);
nand U10889 (N_10889,N_10588,N_10694);
xor U10890 (N_10890,N_10738,N_10657);
nor U10891 (N_10891,N_10594,N_10667);
nor U10892 (N_10892,N_10554,N_10590);
or U10893 (N_10893,N_10637,N_10664);
xnor U10894 (N_10894,N_10651,N_10703);
nor U10895 (N_10895,N_10587,N_10721);
nor U10896 (N_10896,N_10678,N_10695);
and U10897 (N_10897,N_10739,N_10637);
nand U10898 (N_10898,N_10558,N_10519);
nor U10899 (N_10899,N_10526,N_10565);
or U10900 (N_10900,N_10545,N_10614);
and U10901 (N_10901,N_10723,N_10525);
and U10902 (N_10902,N_10544,N_10555);
xnor U10903 (N_10903,N_10544,N_10505);
and U10904 (N_10904,N_10565,N_10529);
nor U10905 (N_10905,N_10595,N_10601);
xor U10906 (N_10906,N_10512,N_10612);
and U10907 (N_10907,N_10669,N_10672);
nor U10908 (N_10908,N_10704,N_10738);
nand U10909 (N_10909,N_10623,N_10742);
nor U10910 (N_10910,N_10617,N_10605);
and U10911 (N_10911,N_10579,N_10583);
and U10912 (N_10912,N_10692,N_10593);
and U10913 (N_10913,N_10657,N_10728);
nor U10914 (N_10914,N_10594,N_10714);
nor U10915 (N_10915,N_10558,N_10621);
nand U10916 (N_10916,N_10570,N_10690);
or U10917 (N_10917,N_10527,N_10526);
and U10918 (N_10918,N_10646,N_10619);
and U10919 (N_10919,N_10745,N_10593);
nand U10920 (N_10920,N_10703,N_10670);
xor U10921 (N_10921,N_10639,N_10570);
nand U10922 (N_10922,N_10733,N_10523);
nor U10923 (N_10923,N_10726,N_10508);
or U10924 (N_10924,N_10686,N_10609);
and U10925 (N_10925,N_10673,N_10510);
or U10926 (N_10926,N_10559,N_10580);
and U10927 (N_10927,N_10552,N_10564);
and U10928 (N_10928,N_10568,N_10580);
nand U10929 (N_10929,N_10670,N_10734);
nor U10930 (N_10930,N_10511,N_10686);
nor U10931 (N_10931,N_10612,N_10503);
nand U10932 (N_10932,N_10605,N_10723);
nand U10933 (N_10933,N_10636,N_10567);
nand U10934 (N_10934,N_10528,N_10500);
and U10935 (N_10935,N_10681,N_10554);
nor U10936 (N_10936,N_10693,N_10691);
xor U10937 (N_10937,N_10606,N_10716);
nor U10938 (N_10938,N_10670,N_10600);
or U10939 (N_10939,N_10626,N_10623);
and U10940 (N_10940,N_10547,N_10507);
and U10941 (N_10941,N_10602,N_10588);
or U10942 (N_10942,N_10616,N_10520);
nand U10943 (N_10943,N_10582,N_10704);
nor U10944 (N_10944,N_10523,N_10701);
or U10945 (N_10945,N_10573,N_10694);
or U10946 (N_10946,N_10712,N_10647);
or U10947 (N_10947,N_10694,N_10706);
nand U10948 (N_10948,N_10531,N_10712);
or U10949 (N_10949,N_10593,N_10710);
nand U10950 (N_10950,N_10561,N_10621);
nand U10951 (N_10951,N_10695,N_10679);
xnor U10952 (N_10952,N_10502,N_10585);
nor U10953 (N_10953,N_10611,N_10544);
or U10954 (N_10954,N_10534,N_10598);
or U10955 (N_10955,N_10696,N_10686);
xor U10956 (N_10956,N_10743,N_10559);
nand U10957 (N_10957,N_10706,N_10684);
and U10958 (N_10958,N_10747,N_10598);
or U10959 (N_10959,N_10611,N_10534);
or U10960 (N_10960,N_10709,N_10565);
nor U10961 (N_10961,N_10523,N_10505);
or U10962 (N_10962,N_10647,N_10510);
xnor U10963 (N_10963,N_10524,N_10730);
or U10964 (N_10964,N_10670,N_10692);
nor U10965 (N_10965,N_10639,N_10660);
xor U10966 (N_10966,N_10522,N_10660);
or U10967 (N_10967,N_10614,N_10540);
xor U10968 (N_10968,N_10596,N_10738);
nor U10969 (N_10969,N_10525,N_10606);
or U10970 (N_10970,N_10733,N_10508);
xnor U10971 (N_10971,N_10745,N_10679);
and U10972 (N_10972,N_10536,N_10694);
and U10973 (N_10973,N_10622,N_10631);
nand U10974 (N_10974,N_10584,N_10733);
nand U10975 (N_10975,N_10665,N_10613);
or U10976 (N_10976,N_10746,N_10562);
nor U10977 (N_10977,N_10677,N_10632);
and U10978 (N_10978,N_10528,N_10604);
xnor U10979 (N_10979,N_10723,N_10673);
nand U10980 (N_10980,N_10614,N_10667);
nor U10981 (N_10981,N_10570,N_10708);
or U10982 (N_10982,N_10618,N_10607);
xnor U10983 (N_10983,N_10651,N_10546);
nor U10984 (N_10984,N_10597,N_10667);
nand U10985 (N_10985,N_10702,N_10695);
xor U10986 (N_10986,N_10674,N_10547);
and U10987 (N_10987,N_10557,N_10660);
or U10988 (N_10988,N_10637,N_10588);
nand U10989 (N_10989,N_10527,N_10512);
nand U10990 (N_10990,N_10663,N_10520);
nor U10991 (N_10991,N_10504,N_10680);
and U10992 (N_10992,N_10563,N_10534);
nor U10993 (N_10993,N_10691,N_10567);
or U10994 (N_10994,N_10700,N_10537);
and U10995 (N_10995,N_10502,N_10642);
nor U10996 (N_10996,N_10554,N_10675);
and U10997 (N_10997,N_10727,N_10691);
or U10998 (N_10998,N_10686,N_10695);
and U10999 (N_10999,N_10644,N_10687);
or U11000 (N_11000,N_10770,N_10994);
and U11001 (N_11001,N_10879,N_10998);
or U11002 (N_11002,N_10999,N_10936);
nand U11003 (N_11003,N_10774,N_10963);
or U11004 (N_11004,N_10938,N_10803);
nor U11005 (N_11005,N_10754,N_10987);
nor U11006 (N_11006,N_10925,N_10769);
nand U11007 (N_11007,N_10771,N_10810);
nor U11008 (N_11008,N_10832,N_10793);
or U11009 (N_11009,N_10910,N_10966);
nor U11010 (N_11010,N_10797,N_10924);
xor U11011 (N_11011,N_10789,N_10864);
and U11012 (N_11012,N_10929,N_10928);
or U11013 (N_11013,N_10950,N_10990);
xor U11014 (N_11014,N_10772,N_10816);
and U11015 (N_11015,N_10942,N_10927);
or U11016 (N_11016,N_10763,N_10861);
nand U11017 (N_11017,N_10777,N_10996);
nand U11018 (N_11018,N_10775,N_10869);
and U11019 (N_11019,N_10930,N_10886);
and U11020 (N_11020,N_10863,N_10842);
or U11021 (N_11021,N_10962,N_10949);
and U11022 (N_11022,N_10909,N_10898);
and U11023 (N_11023,N_10812,N_10795);
nand U11024 (N_11024,N_10979,N_10752);
or U11025 (N_11025,N_10824,N_10917);
and U11026 (N_11026,N_10857,N_10757);
xnor U11027 (N_11027,N_10884,N_10891);
nor U11028 (N_11028,N_10756,N_10941);
nor U11029 (N_11029,N_10858,N_10843);
or U11030 (N_11030,N_10764,N_10937);
nor U11031 (N_11031,N_10867,N_10953);
xnor U11032 (N_11032,N_10836,N_10922);
or U11033 (N_11033,N_10776,N_10798);
and U11034 (N_11034,N_10888,N_10750);
xnor U11035 (N_11035,N_10915,N_10872);
xnor U11036 (N_11036,N_10782,N_10823);
and U11037 (N_11037,N_10862,N_10956);
nand U11038 (N_11038,N_10830,N_10779);
xor U11039 (N_11039,N_10766,N_10960);
nand U11040 (N_11040,N_10874,N_10762);
nor U11041 (N_11041,N_10838,N_10989);
xor U11042 (N_11042,N_10801,N_10918);
and U11043 (N_11043,N_10903,N_10759);
nor U11044 (N_11044,N_10880,N_10977);
xnor U11045 (N_11045,N_10761,N_10995);
nand U11046 (N_11046,N_10961,N_10947);
nor U11047 (N_11047,N_10984,N_10800);
nand U11048 (N_11048,N_10943,N_10780);
xnor U11049 (N_11049,N_10968,N_10881);
or U11050 (N_11050,N_10852,N_10934);
xor U11051 (N_11051,N_10786,N_10983);
nor U11052 (N_11052,N_10908,N_10844);
nor U11053 (N_11053,N_10846,N_10828);
and U11054 (N_11054,N_10971,N_10818);
xor U11055 (N_11055,N_10975,N_10785);
xor U11056 (N_11056,N_10912,N_10951);
and U11057 (N_11057,N_10760,N_10957);
and U11058 (N_11058,N_10871,N_10964);
xor U11059 (N_11059,N_10856,N_10866);
and U11060 (N_11060,N_10913,N_10976);
xnor U11061 (N_11061,N_10887,N_10940);
and U11062 (N_11062,N_10948,N_10893);
nand U11063 (N_11063,N_10933,N_10821);
nor U11064 (N_11064,N_10973,N_10926);
nor U11065 (N_11065,N_10794,N_10802);
or U11066 (N_11066,N_10847,N_10851);
or U11067 (N_11067,N_10945,N_10952);
or U11068 (N_11068,N_10875,N_10972);
nor U11069 (N_11069,N_10820,N_10905);
nand U11070 (N_11070,N_10923,N_10981);
xor U11071 (N_11071,N_10768,N_10868);
nor U11072 (N_11072,N_10788,N_10982);
xor U11073 (N_11073,N_10767,N_10819);
xnor U11074 (N_11074,N_10817,N_10826);
or U11075 (N_11075,N_10882,N_10865);
and U11076 (N_11076,N_10921,N_10970);
nor U11077 (N_11077,N_10946,N_10758);
nor U11078 (N_11078,N_10799,N_10753);
xnor U11079 (N_11079,N_10958,N_10906);
or U11080 (N_11080,N_10988,N_10877);
and U11081 (N_11081,N_10839,N_10900);
nand U11082 (N_11082,N_10849,N_10831);
nand U11083 (N_11083,N_10791,N_10916);
nor U11084 (N_11084,N_10944,N_10805);
nand U11085 (N_11085,N_10876,N_10809);
and U11086 (N_11086,N_10833,N_10840);
and U11087 (N_11087,N_10787,N_10808);
nand U11088 (N_11088,N_10901,N_10837);
nand U11089 (N_11089,N_10997,N_10784);
and U11090 (N_11090,N_10827,N_10907);
and U11091 (N_11091,N_10811,N_10954);
or U11092 (N_11092,N_10778,N_10781);
nand U11093 (N_11093,N_10878,N_10919);
or U11094 (N_11094,N_10969,N_10792);
xor U11095 (N_11095,N_10902,N_10993);
or U11096 (N_11096,N_10765,N_10755);
and U11097 (N_11097,N_10829,N_10790);
nand U11098 (N_11098,N_10806,N_10895);
and U11099 (N_11099,N_10935,N_10796);
or U11100 (N_11100,N_10897,N_10955);
nand U11101 (N_11101,N_10932,N_10894);
nand U11102 (N_11102,N_10914,N_10889);
nor U11103 (N_11103,N_10822,N_10967);
or U11104 (N_11104,N_10854,N_10773);
xnor U11105 (N_11105,N_10853,N_10992);
nor U11106 (N_11106,N_10848,N_10815);
and U11107 (N_11107,N_10841,N_10890);
xor U11108 (N_11108,N_10985,N_10859);
nand U11109 (N_11109,N_10873,N_10870);
or U11110 (N_11110,N_10899,N_10860);
or U11111 (N_11111,N_10978,N_10845);
and U11112 (N_11112,N_10751,N_10965);
xnor U11113 (N_11113,N_10813,N_10920);
and U11114 (N_11114,N_10783,N_10892);
and U11115 (N_11115,N_10904,N_10911);
nand U11116 (N_11116,N_10991,N_10980);
and U11117 (N_11117,N_10804,N_10986);
nor U11118 (N_11118,N_10834,N_10883);
or U11119 (N_11119,N_10855,N_10896);
nor U11120 (N_11120,N_10814,N_10825);
nor U11121 (N_11121,N_10885,N_10974);
xnor U11122 (N_11122,N_10939,N_10807);
xnor U11123 (N_11123,N_10835,N_10931);
and U11124 (N_11124,N_10959,N_10850);
xor U11125 (N_11125,N_10898,N_10781);
or U11126 (N_11126,N_10885,N_10929);
or U11127 (N_11127,N_10794,N_10777);
nand U11128 (N_11128,N_10949,N_10785);
nand U11129 (N_11129,N_10923,N_10995);
or U11130 (N_11130,N_10971,N_10838);
and U11131 (N_11131,N_10803,N_10905);
and U11132 (N_11132,N_10961,N_10763);
nand U11133 (N_11133,N_10983,N_10788);
nand U11134 (N_11134,N_10836,N_10793);
nand U11135 (N_11135,N_10950,N_10945);
nor U11136 (N_11136,N_10840,N_10850);
xor U11137 (N_11137,N_10776,N_10997);
and U11138 (N_11138,N_10992,N_10985);
and U11139 (N_11139,N_10757,N_10844);
nand U11140 (N_11140,N_10981,N_10757);
or U11141 (N_11141,N_10795,N_10940);
and U11142 (N_11142,N_10951,N_10888);
and U11143 (N_11143,N_10879,N_10947);
and U11144 (N_11144,N_10883,N_10977);
xor U11145 (N_11145,N_10959,N_10808);
and U11146 (N_11146,N_10777,N_10822);
nand U11147 (N_11147,N_10899,N_10927);
and U11148 (N_11148,N_10946,N_10896);
or U11149 (N_11149,N_10884,N_10975);
nand U11150 (N_11150,N_10769,N_10755);
or U11151 (N_11151,N_10974,N_10874);
nand U11152 (N_11152,N_10832,N_10852);
nor U11153 (N_11153,N_10935,N_10757);
xor U11154 (N_11154,N_10854,N_10912);
nand U11155 (N_11155,N_10934,N_10787);
or U11156 (N_11156,N_10854,N_10960);
or U11157 (N_11157,N_10980,N_10886);
xor U11158 (N_11158,N_10823,N_10997);
nand U11159 (N_11159,N_10859,N_10883);
or U11160 (N_11160,N_10785,N_10858);
nor U11161 (N_11161,N_10844,N_10956);
xor U11162 (N_11162,N_10897,N_10960);
and U11163 (N_11163,N_10799,N_10906);
nand U11164 (N_11164,N_10795,N_10822);
nand U11165 (N_11165,N_10913,N_10891);
and U11166 (N_11166,N_10981,N_10916);
and U11167 (N_11167,N_10889,N_10869);
or U11168 (N_11168,N_10769,N_10783);
or U11169 (N_11169,N_10901,N_10752);
xnor U11170 (N_11170,N_10916,N_10815);
and U11171 (N_11171,N_10825,N_10962);
or U11172 (N_11172,N_10813,N_10791);
nor U11173 (N_11173,N_10872,N_10877);
nor U11174 (N_11174,N_10812,N_10823);
or U11175 (N_11175,N_10866,N_10986);
nor U11176 (N_11176,N_10802,N_10814);
xnor U11177 (N_11177,N_10964,N_10802);
and U11178 (N_11178,N_10769,N_10771);
or U11179 (N_11179,N_10750,N_10873);
nand U11180 (N_11180,N_10955,N_10853);
or U11181 (N_11181,N_10962,N_10993);
and U11182 (N_11182,N_10990,N_10765);
or U11183 (N_11183,N_10802,N_10945);
nand U11184 (N_11184,N_10949,N_10763);
or U11185 (N_11185,N_10927,N_10827);
nand U11186 (N_11186,N_10875,N_10936);
or U11187 (N_11187,N_10990,N_10945);
xor U11188 (N_11188,N_10899,N_10987);
xnor U11189 (N_11189,N_10846,N_10899);
and U11190 (N_11190,N_10756,N_10827);
nand U11191 (N_11191,N_10786,N_10958);
nor U11192 (N_11192,N_10837,N_10889);
nand U11193 (N_11193,N_10999,N_10982);
nand U11194 (N_11194,N_10855,N_10885);
nand U11195 (N_11195,N_10783,N_10951);
and U11196 (N_11196,N_10923,N_10800);
nand U11197 (N_11197,N_10947,N_10791);
xor U11198 (N_11198,N_10891,N_10760);
and U11199 (N_11199,N_10798,N_10969);
or U11200 (N_11200,N_10844,N_10843);
nand U11201 (N_11201,N_10947,N_10980);
xor U11202 (N_11202,N_10795,N_10991);
nand U11203 (N_11203,N_10819,N_10964);
nand U11204 (N_11204,N_10980,N_10840);
nand U11205 (N_11205,N_10859,N_10909);
or U11206 (N_11206,N_10877,N_10978);
and U11207 (N_11207,N_10998,N_10903);
xnor U11208 (N_11208,N_10875,N_10938);
nor U11209 (N_11209,N_10806,N_10826);
xnor U11210 (N_11210,N_10765,N_10763);
or U11211 (N_11211,N_10988,N_10980);
and U11212 (N_11212,N_10857,N_10780);
xnor U11213 (N_11213,N_10860,N_10941);
and U11214 (N_11214,N_10838,N_10890);
nand U11215 (N_11215,N_10883,N_10951);
and U11216 (N_11216,N_10794,N_10837);
nand U11217 (N_11217,N_10852,N_10835);
or U11218 (N_11218,N_10822,N_10935);
xnor U11219 (N_11219,N_10786,N_10939);
nand U11220 (N_11220,N_10889,N_10847);
xnor U11221 (N_11221,N_10785,N_10956);
and U11222 (N_11222,N_10855,N_10957);
nor U11223 (N_11223,N_10778,N_10854);
xor U11224 (N_11224,N_10874,N_10872);
nand U11225 (N_11225,N_10884,N_10864);
xor U11226 (N_11226,N_10971,N_10925);
nand U11227 (N_11227,N_10831,N_10794);
and U11228 (N_11228,N_10929,N_10768);
nor U11229 (N_11229,N_10866,N_10835);
or U11230 (N_11230,N_10840,N_10960);
xnor U11231 (N_11231,N_10937,N_10771);
or U11232 (N_11232,N_10821,N_10754);
xor U11233 (N_11233,N_10990,N_10805);
nor U11234 (N_11234,N_10902,N_10932);
xnor U11235 (N_11235,N_10909,N_10789);
nor U11236 (N_11236,N_10879,N_10835);
nand U11237 (N_11237,N_10829,N_10796);
xnor U11238 (N_11238,N_10810,N_10955);
nand U11239 (N_11239,N_10783,N_10931);
and U11240 (N_11240,N_10914,N_10882);
and U11241 (N_11241,N_10983,N_10793);
nand U11242 (N_11242,N_10789,N_10824);
and U11243 (N_11243,N_10933,N_10982);
and U11244 (N_11244,N_10867,N_10949);
nor U11245 (N_11245,N_10901,N_10756);
or U11246 (N_11246,N_10933,N_10825);
xnor U11247 (N_11247,N_10847,N_10965);
xor U11248 (N_11248,N_10844,N_10909);
or U11249 (N_11249,N_10983,N_10826);
nor U11250 (N_11250,N_11008,N_11179);
nand U11251 (N_11251,N_11241,N_11245);
or U11252 (N_11252,N_11076,N_11212);
or U11253 (N_11253,N_11244,N_11223);
or U11254 (N_11254,N_11208,N_11042);
or U11255 (N_11255,N_11003,N_11124);
nand U11256 (N_11256,N_11065,N_11183);
xnor U11257 (N_11257,N_11221,N_11153);
xor U11258 (N_11258,N_11049,N_11031);
xor U11259 (N_11259,N_11155,N_11024);
and U11260 (N_11260,N_11194,N_11072);
xnor U11261 (N_11261,N_11149,N_11226);
and U11262 (N_11262,N_11197,N_11173);
or U11263 (N_11263,N_11112,N_11047);
nand U11264 (N_11264,N_11123,N_11094);
nor U11265 (N_11265,N_11128,N_11106);
or U11266 (N_11266,N_11205,N_11032);
nor U11267 (N_11267,N_11247,N_11063);
nand U11268 (N_11268,N_11014,N_11145);
nand U11269 (N_11269,N_11138,N_11109);
and U11270 (N_11270,N_11136,N_11185);
nor U11271 (N_11271,N_11007,N_11216);
xor U11272 (N_11272,N_11044,N_11019);
and U11273 (N_11273,N_11006,N_11079);
nor U11274 (N_11274,N_11078,N_11059);
or U11275 (N_11275,N_11141,N_11131);
xnor U11276 (N_11276,N_11096,N_11161);
nand U11277 (N_11277,N_11005,N_11229);
xor U11278 (N_11278,N_11175,N_11126);
or U11279 (N_11279,N_11115,N_11129);
and U11280 (N_11280,N_11025,N_11172);
nor U11281 (N_11281,N_11052,N_11061);
nor U11282 (N_11282,N_11043,N_11224);
and U11283 (N_11283,N_11091,N_11217);
nand U11284 (N_11284,N_11240,N_11002);
or U11285 (N_11285,N_11009,N_11162);
or U11286 (N_11286,N_11215,N_11102);
and U11287 (N_11287,N_11133,N_11021);
nor U11288 (N_11288,N_11195,N_11000);
nand U11289 (N_11289,N_11146,N_11236);
nand U11290 (N_11290,N_11062,N_11202);
and U11291 (N_11291,N_11120,N_11068);
nand U11292 (N_11292,N_11203,N_11100);
nand U11293 (N_11293,N_11222,N_11249);
xor U11294 (N_11294,N_11151,N_11142);
nor U11295 (N_11295,N_11054,N_11200);
nor U11296 (N_11296,N_11070,N_11088);
xor U11297 (N_11297,N_11035,N_11103);
nor U11298 (N_11298,N_11191,N_11218);
or U11299 (N_11299,N_11204,N_11225);
or U11300 (N_11300,N_11199,N_11206);
nand U11301 (N_11301,N_11098,N_11234);
nor U11302 (N_11302,N_11028,N_11022);
or U11303 (N_11303,N_11159,N_11227);
nor U11304 (N_11304,N_11140,N_11117);
or U11305 (N_11305,N_11108,N_11015);
nor U11306 (N_11306,N_11132,N_11107);
nand U11307 (N_11307,N_11011,N_11013);
or U11308 (N_11308,N_11119,N_11233);
or U11309 (N_11309,N_11178,N_11087);
xnor U11310 (N_11310,N_11186,N_11080);
nand U11311 (N_11311,N_11093,N_11248);
xnor U11312 (N_11312,N_11198,N_11160);
nand U11313 (N_11313,N_11020,N_11023);
and U11314 (N_11314,N_11125,N_11239);
xnor U11315 (N_11315,N_11097,N_11074);
and U11316 (N_11316,N_11104,N_11127);
and U11317 (N_11317,N_11040,N_11235);
or U11318 (N_11318,N_11134,N_11111);
or U11319 (N_11319,N_11069,N_11148);
xnor U11320 (N_11320,N_11039,N_11037);
nand U11321 (N_11321,N_11150,N_11174);
nand U11322 (N_11322,N_11213,N_11116);
xor U11323 (N_11323,N_11196,N_11018);
nor U11324 (N_11324,N_11114,N_11182);
nand U11325 (N_11325,N_11004,N_11230);
nand U11326 (N_11326,N_11036,N_11164);
nand U11327 (N_11327,N_11056,N_11033);
or U11328 (N_11328,N_11163,N_11077);
nor U11329 (N_11329,N_11167,N_11169);
xnor U11330 (N_11330,N_11110,N_11026);
nor U11331 (N_11331,N_11075,N_11029);
xor U11332 (N_11332,N_11232,N_11053);
and U11333 (N_11333,N_11209,N_11228);
nor U11334 (N_11334,N_11066,N_11084);
nand U11335 (N_11335,N_11176,N_11154);
xnor U11336 (N_11336,N_11030,N_11012);
or U11337 (N_11337,N_11189,N_11089);
and U11338 (N_11338,N_11046,N_11187);
nor U11339 (N_11339,N_11237,N_11242);
nand U11340 (N_11340,N_11058,N_11016);
or U11341 (N_11341,N_11017,N_11055);
and U11342 (N_11342,N_11158,N_11188);
nand U11343 (N_11343,N_11171,N_11207);
nor U11344 (N_11344,N_11211,N_11051);
or U11345 (N_11345,N_11192,N_11214);
nand U11346 (N_11346,N_11081,N_11121);
and U11347 (N_11347,N_11048,N_11034);
xnor U11348 (N_11348,N_11105,N_11010);
and U11349 (N_11349,N_11038,N_11041);
xor U11350 (N_11350,N_11139,N_11190);
xor U11351 (N_11351,N_11181,N_11170);
or U11352 (N_11352,N_11095,N_11118);
xnor U11353 (N_11353,N_11135,N_11156);
or U11354 (N_11354,N_11220,N_11184);
nand U11355 (N_11355,N_11137,N_11219);
xor U11356 (N_11356,N_11165,N_11083);
nor U11357 (N_11357,N_11113,N_11168);
xor U11358 (N_11358,N_11152,N_11166);
or U11359 (N_11359,N_11243,N_11177);
xnor U11360 (N_11360,N_11057,N_11067);
nor U11361 (N_11361,N_11090,N_11045);
nand U11362 (N_11362,N_11050,N_11082);
and U11363 (N_11363,N_11071,N_11238);
and U11364 (N_11364,N_11064,N_11085);
xnor U11365 (N_11365,N_11143,N_11193);
and U11366 (N_11366,N_11246,N_11086);
and U11367 (N_11367,N_11157,N_11060);
and U11368 (N_11368,N_11201,N_11092);
xor U11369 (N_11369,N_11027,N_11122);
nand U11370 (N_11370,N_11101,N_11147);
nand U11371 (N_11371,N_11180,N_11231);
and U11372 (N_11372,N_11210,N_11099);
nor U11373 (N_11373,N_11130,N_11001);
or U11374 (N_11374,N_11073,N_11144);
or U11375 (N_11375,N_11039,N_11141);
nor U11376 (N_11376,N_11013,N_11246);
xnor U11377 (N_11377,N_11029,N_11176);
xnor U11378 (N_11378,N_11173,N_11210);
nand U11379 (N_11379,N_11191,N_11010);
xor U11380 (N_11380,N_11225,N_11121);
or U11381 (N_11381,N_11189,N_11194);
or U11382 (N_11382,N_11002,N_11198);
nand U11383 (N_11383,N_11040,N_11101);
xnor U11384 (N_11384,N_11231,N_11067);
and U11385 (N_11385,N_11098,N_11141);
and U11386 (N_11386,N_11087,N_11213);
and U11387 (N_11387,N_11065,N_11067);
xor U11388 (N_11388,N_11110,N_11149);
nor U11389 (N_11389,N_11001,N_11073);
nor U11390 (N_11390,N_11121,N_11240);
or U11391 (N_11391,N_11007,N_11052);
or U11392 (N_11392,N_11002,N_11059);
nand U11393 (N_11393,N_11091,N_11123);
nand U11394 (N_11394,N_11119,N_11089);
xnor U11395 (N_11395,N_11103,N_11161);
nor U11396 (N_11396,N_11238,N_11081);
xor U11397 (N_11397,N_11005,N_11145);
nor U11398 (N_11398,N_11144,N_11210);
nand U11399 (N_11399,N_11133,N_11071);
nand U11400 (N_11400,N_11137,N_11037);
nor U11401 (N_11401,N_11231,N_11159);
nand U11402 (N_11402,N_11218,N_11133);
nor U11403 (N_11403,N_11122,N_11056);
xor U11404 (N_11404,N_11028,N_11153);
or U11405 (N_11405,N_11182,N_11229);
nor U11406 (N_11406,N_11149,N_11006);
nand U11407 (N_11407,N_11078,N_11098);
nand U11408 (N_11408,N_11213,N_11050);
xor U11409 (N_11409,N_11197,N_11107);
or U11410 (N_11410,N_11230,N_11248);
or U11411 (N_11411,N_11208,N_11117);
or U11412 (N_11412,N_11186,N_11062);
xnor U11413 (N_11413,N_11204,N_11077);
nand U11414 (N_11414,N_11030,N_11241);
and U11415 (N_11415,N_11152,N_11082);
and U11416 (N_11416,N_11006,N_11241);
nand U11417 (N_11417,N_11230,N_11106);
and U11418 (N_11418,N_11021,N_11146);
and U11419 (N_11419,N_11140,N_11030);
or U11420 (N_11420,N_11068,N_11224);
or U11421 (N_11421,N_11228,N_11213);
nand U11422 (N_11422,N_11153,N_11089);
xor U11423 (N_11423,N_11221,N_11186);
and U11424 (N_11424,N_11078,N_11002);
and U11425 (N_11425,N_11076,N_11101);
xnor U11426 (N_11426,N_11167,N_11240);
xor U11427 (N_11427,N_11162,N_11041);
or U11428 (N_11428,N_11197,N_11136);
or U11429 (N_11429,N_11187,N_11057);
nand U11430 (N_11430,N_11194,N_11167);
or U11431 (N_11431,N_11066,N_11053);
and U11432 (N_11432,N_11091,N_11138);
xnor U11433 (N_11433,N_11021,N_11134);
nand U11434 (N_11434,N_11025,N_11184);
and U11435 (N_11435,N_11111,N_11087);
or U11436 (N_11436,N_11207,N_11108);
nand U11437 (N_11437,N_11111,N_11127);
nor U11438 (N_11438,N_11132,N_11110);
or U11439 (N_11439,N_11188,N_11105);
nand U11440 (N_11440,N_11126,N_11157);
or U11441 (N_11441,N_11067,N_11234);
nand U11442 (N_11442,N_11084,N_11248);
nand U11443 (N_11443,N_11114,N_11156);
and U11444 (N_11444,N_11177,N_11159);
nand U11445 (N_11445,N_11095,N_11196);
nand U11446 (N_11446,N_11103,N_11097);
xor U11447 (N_11447,N_11150,N_11065);
nor U11448 (N_11448,N_11237,N_11199);
or U11449 (N_11449,N_11148,N_11094);
nor U11450 (N_11450,N_11011,N_11035);
nor U11451 (N_11451,N_11068,N_11034);
nand U11452 (N_11452,N_11158,N_11202);
and U11453 (N_11453,N_11237,N_11196);
nor U11454 (N_11454,N_11166,N_11126);
nor U11455 (N_11455,N_11187,N_11197);
or U11456 (N_11456,N_11143,N_11134);
nand U11457 (N_11457,N_11170,N_11172);
xor U11458 (N_11458,N_11075,N_11078);
nand U11459 (N_11459,N_11246,N_11003);
and U11460 (N_11460,N_11000,N_11004);
or U11461 (N_11461,N_11088,N_11098);
nor U11462 (N_11462,N_11050,N_11249);
nor U11463 (N_11463,N_11033,N_11044);
xnor U11464 (N_11464,N_11001,N_11220);
nor U11465 (N_11465,N_11108,N_11090);
xnor U11466 (N_11466,N_11006,N_11196);
nor U11467 (N_11467,N_11093,N_11206);
nor U11468 (N_11468,N_11113,N_11080);
xor U11469 (N_11469,N_11198,N_11151);
or U11470 (N_11470,N_11037,N_11239);
and U11471 (N_11471,N_11174,N_11006);
xnor U11472 (N_11472,N_11142,N_11019);
or U11473 (N_11473,N_11068,N_11211);
nand U11474 (N_11474,N_11061,N_11162);
or U11475 (N_11475,N_11116,N_11065);
and U11476 (N_11476,N_11109,N_11163);
nor U11477 (N_11477,N_11248,N_11044);
xor U11478 (N_11478,N_11062,N_11236);
nand U11479 (N_11479,N_11224,N_11197);
xnor U11480 (N_11480,N_11184,N_11133);
or U11481 (N_11481,N_11192,N_11038);
nand U11482 (N_11482,N_11230,N_11175);
and U11483 (N_11483,N_11148,N_11141);
nand U11484 (N_11484,N_11062,N_11013);
xnor U11485 (N_11485,N_11089,N_11120);
nor U11486 (N_11486,N_11197,N_11119);
nor U11487 (N_11487,N_11060,N_11246);
nand U11488 (N_11488,N_11012,N_11122);
nand U11489 (N_11489,N_11117,N_11180);
nand U11490 (N_11490,N_11249,N_11145);
nand U11491 (N_11491,N_11219,N_11238);
nand U11492 (N_11492,N_11060,N_11081);
and U11493 (N_11493,N_11186,N_11143);
nand U11494 (N_11494,N_11012,N_11066);
xnor U11495 (N_11495,N_11190,N_11206);
nor U11496 (N_11496,N_11011,N_11043);
nand U11497 (N_11497,N_11171,N_11068);
or U11498 (N_11498,N_11241,N_11013);
and U11499 (N_11499,N_11244,N_11027);
or U11500 (N_11500,N_11408,N_11251);
nand U11501 (N_11501,N_11498,N_11427);
and U11502 (N_11502,N_11422,N_11256);
nand U11503 (N_11503,N_11428,N_11284);
xnor U11504 (N_11504,N_11357,N_11341);
and U11505 (N_11505,N_11296,N_11454);
nor U11506 (N_11506,N_11295,N_11368);
nand U11507 (N_11507,N_11349,N_11336);
xnor U11508 (N_11508,N_11412,N_11274);
xor U11509 (N_11509,N_11483,N_11437);
and U11510 (N_11510,N_11433,N_11337);
or U11511 (N_11511,N_11384,N_11457);
xnor U11512 (N_11512,N_11345,N_11400);
and U11513 (N_11513,N_11394,N_11312);
nand U11514 (N_11514,N_11405,N_11373);
nor U11515 (N_11515,N_11260,N_11287);
nor U11516 (N_11516,N_11424,N_11329);
xnor U11517 (N_11517,N_11276,N_11436);
or U11518 (N_11518,N_11263,N_11262);
xnor U11519 (N_11519,N_11397,N_11451);
and U11520 (N_11520,N_11320,N_11372);
nor U11521 (N_11521,N_11286,N_11347);
nor U11522 (N_11522,N_11317,N_11448);
xor U11523 (N_11523,N_11315,N_11302);
or U11524 (N_11524,N_11499,N_11406);
nor U11525 (N_11525,N_11378,N_11455);
or U11526 (N_11526,N_11355,N_11361);
xor U11527 (N_11527,N_11362,N_11281);
or U11528 (N_11528,N_11266,N_11356);
and U11529 (N_11529,N_11294,N_11444);
xnor U11530 (N_11530,N_11407,N_11385);
nor U11531 (N_11531,N_11342,N_11461);
or U11532 (N_11532,N_11282,N_11414);
nand U11533 (N_11533,N_11490,N_11478);
nor U11534 (N_11534,N_11321,N_11323);
and U11535 (N_11535,N_11418,N_11253);
xnor U11536 (N_11536,N_11423,N_11370);
nand U11537 (N_11537,N_11460,N_11268);
and U11538 (N_11538,N_11402,N_11421);
xnor U11539 (N_11539,N_11419,N_11261);
or U11540 (N_11540,N_11403,N_11464);
nand U11541 (N_11541,N_11482,N_11279);
xnor U11542 (N_11542,N_11369,N_11495);
nor U11543 (N_11543,N_11270,N_11484);
xnor U11544 (N_11544,N_11365,N_11389);
or U11545 (N_11545,N_11308,N_11469);
xor U11546 (N_11546,N_11387,N_11398);
and U11547 (N_11547,N_11366,N_11364);
or U11548 (N_11548,N_11440,N_11458);
nand U11549 (N_11549,N_11272,N_11360);
or U11550 (N_11550,N_11379,N_11472);
xor U11551 (N_11551,N_11486,N_11380);
nor U11552 (N_11552,N_11273,N_11415);
or U11553 (N_11553,N_11326,N_11447);
or U11554 (N_11554,N_11250,N_11258);
or U11555 (N_11555,N_11333,N_11462);
nor U11556 (N_11556,N_11376,N_11339);
nor U11557 (N_11557,N_11485,N_11453);
or U11558 (N_11558,N_11442,N_11316);
and U11559 (N_11559,N_11393,N_11346);
nor U11560 (N_11560,N_11252,N_11497);
xor U11561 (N_11561,N_11435,N_11471);
nand U11562 (N_11562,N_11374,N_11306);
nand U11563 (N_11563,N_11330,N_11310);
xnor U11564 (N_11564,N_11494,N_11446);
nand U11565 (N_11565,N_11322,N_11354);
and U11566 (N_11566,N_11430,N_11324);
and U11567 (N_11567,N_11409,N_11476);
nand U11568 (N_11568,N_11340,N_11328);
or U11569 (N_11569,N_11488,N_11290);
xor U11570 (N_11570,N_11416,N_11467);
xnor U11571 (N_11571,N_11371,N_11386);
or U11572 (N_11572,N_11283,N_11420);
and U11573 (N_11573,N_11275,N_11265);
nand U11574 (N_11574,N_11410,N_11417);
and U11575 (N_11575,N_11300,N_11363);
nand U11576 (N_11576,N_11277,N_11473);
xor U11577 (N_11577,N_11441,N_11309);
nand U11578 (N_11578,N_11477,N_11289);
xnor U11579 (N_11579,N_11470,N_11267);
xor U11580 (N_11580,N_11381,N_11431);
or U11581 (N_11581,N_11307,N_11313);
xnor U11582 (N_11582,N_11297,N_11429);
and U11583 (N_11583,N_11331,N_11259);
nand U11584 (N_11584,N_11404,N_11311);
nor U11585 (N_11585,N_11450,N_11318);
or U11586 (N_11586,N_11390,N_11353);
xnor U11587 (N_11587,N_11491,N_11487);
nor U11588 (N_11588,N_11280,N_11288);
nor U11589 (N_11589,N_11481,N_11257);
and U11590 (N_11590,N_11375,N_11438);
nand U11591 (N_11591,N_11468,N_11425);
or U11592 (N_11592,N_11350,N_11269);
nand U11593 (N_11593,N_11334,N_11434);
nand U11594 (N_11594,N_11411,N_11474);
xnor U11595 (N_11595,N_11348,N_11399);
nand U11596 (N_11596,N_11383,N_11452);
and U11597 (N_11597,N_11303,N_11352);
xnor U11598 (N_11598,N_11332,N_11396);
nor U11599 (N_11599,N_11278,N_11432);
or U11600 (N_11600,N_11392,N_11382);
or U11601 (N_11601,N_11377,N_11344);
nor U11602 (N_11602,N_11335,N_11314);
xor U11603 (N_11603,N_11271,N_11449);
xnor U11604 (N_11604,N_11298,N_11343);
and U11605 (N_11605,N_11305,N_11254);
xor U11606 (N_11606,N_11463,N_11264);
and U11607 (N_11607,N_11489,N_11475);
or U11608 (N_11608,N_11443,N_11480);
and U11609 (N_11609,N_11319,N_11493);
nand U11610 (N_11610,N_11255,N_11445);
nand U11611 (N_11611,N_11285,N_11388);
xor U11612 (N_11612,N_11395,N_11496);
or U11613 (N_11613,N_11401,N_11359);
nand U11614 (N_11614,N_11338,N_11367);
and U11615 (N_11615,N_11292,N_11291);
nor U11616 (N_11616,N_11492,N_11479);
nand U11617 (N_11617,N_11465,N_11327);
nand U11618 (N_11618,N_11358,N_11301);
or U11619 (N_11619,N_11299,N_11439);
or U11620 (N_11620,N_11456,N_11293);
nand U11621 (N_11621,N_11459,N_11413);
nor U11622 (N_11622,N_11466,N_11325);
nor U11623 (N_11623,N_11304,N_11391);
xnor U11624 (N_11624,N_11351,N_11426);
nor U11625 (N_11625,N_11447,N_11259);
xor U11626 (N_11626,N_11473,N_11422);
xor U11627 (N_11627,N_11478,N_11449);
or U11628 (N_11628,N_11430,N_11420);
or U11629 (N_11629,N_11449,N_11354);
or U11630 (N_11630,N_11404,N_11328);
or U11631 (N_11631,N_11482,N_11335);
nand U11632 (N_11632,N_11383,N_11308);
nand U11633 (N_11633,N_11332,N_11270);
or U11634 (N_11634,N_11497,N_11405);
nor U11635 (N_11635,N_11420,N_11355);
xor U11636 (N_11636,N_11455,N_11309);
nand U11637 (N_11637,N_11394,N_11300);
or U11638 (N_11638,N_11250,N_11294);
nand U11639 (N_11639,N_11256,N_11270);
xnor U11640 (N_11640,N_11362,N_11308);
and U11641 (N_11641,N_11487,N_11281);
nand U11642 (N_11642,N_11463,N_11251);
or U11643 (N_11643,N_11284,N_11431);
xnor U11644 (N_11644,N_11372,N_11381);
and U11645 (N_11645,N_11474,N_11284);
and U11646 (N_11646,N_11302,N_11334);
or U11647 (N_11647,N_11373,N_11317);
and U11648 (N_11648,N_11441,N_11488);
or U11649 (N_11649,N_11476,N_11378);
and U11650 (N_11650,N_11272,N_11495);
nand U11651 (N_11651,N_11419,N_11461);
xor U11652 (N_11652,N_11485,N_11324);
or U11653 (N_11653,N_11404,N_11304);
xor U11654 (N_11654,N_11478,N_11467);
xnor U11655 (N_11655,N_11407,N_11410);
nor U11656 (N_11656,N_11255,N_11310);
nand U11657 (N_11657,N_11325,N_11458);
nor U11658 (N_11658,N_11267,N_11332);
or U11659 (N_11659,N_11424,N_11386);
nand U11660 (N_11660,N_11311,N_11299);
xnor U11661 (N_11661,N_11276,N_11365);
and U11662 (N_11662,N_11306,N_11272);
or U11663 (N_11663,N_11396,N_11392);
nor U11664 (N_11664,N_11362,N_11305);
or U11665 (N_11665,N_11290,N_11371);
nor U11666 (N_11666,N_11371,N_11495);
nor U11667 (N_11667,N_11252,N_11344);
and U11668 (N_11668,N_11458,N_11264);
nor U11669 (N_11669,N_11419,N_11268);
xor U11670 (N_11670,N_11289,N_11308);
xor U11671 (N_11671,N_11371,N_11314);
xnor U11672 (N_11672,N_11446,N_11392);
or U11673 (N_11673,N_11373,N_11447);
or U11674 (N_11674,N_11358,N_11454);
xnor U11675 (N_11675,N_11466,N_11426);
nand U11676 (N_11676,N_11322,N_11478);
nor U11677 (N_11677,N_11254,N_11413);
xor U11678 (N_11678,N_11375,N_11266);
xnor U11679 (N_11679,N_11394,N_11476);
nand U11680 (N_11680,N_11281,N_11345);
and U11681 (N_11681,N_11274,N_11255);
or U11682 (N_11682,N_11410,N_11416);
or U11683 (N_11683,N_11361,N_11400);
nor U11684 (N_11684,N_11401,N_11271);
xor U11685 (N_11685,N_11429,N_11356);
nand U11686 (N_11686,N_11344,N_11385);
and U11687 (N_11687,N_11391,N_11447);
xor U11688 (N_11688,N_11272,N_11493);
xnor U11689 (N_11689,N_11438,N_11431);
xnor U11690 (N_11690,N_11346,N_11331);
and U11691 (N_11691,N_11472,N_11278);
nand U11692 (N_11692,N_11439,N_11270);
or U11693 (N_11693,N_11361,N_11266);
nand U11694 (N_11694,N_11311,N_11360);
nor U11695 (N_11695,N_11426,N_11277);
nand U11696 (N_11696,N_11373,N_11365);
or U11697 (N_11697,N_11349,N_11413);
or U11698 (N_11698,N_11293,N_11362);
or U11699 (N_11699,N_11250,N_11327);
nor U11700 (N_11700,N_11260,N_11317);
and U11701 (N_11701,N_11417,N_11346);
or U11702 (N_11702,N_11283,N_11459);
nand U11703 (N_11703,N_11371,N_11357);
or U11704 (N_11704,N_11372,N_11330);
and U11705 (N_11705,N_11469,N_11411);
and U11706 (N_11706,N_11425,N_11290);
nand U11707 (N_11707,N_11428,N_11389);
or U11708 (N_11708,N_11361,N_11498);
xnor U11709 (N_11709,N_11279,N_11271);
and U11710 (N_11710,N_11355,N_11430);
and U11711 (N_11711,N_11447,N_11338);
or U11712 (N_11712,N_11273,N_11469);
nor U11713 (N_11713,N_11492,N_11461);
nor U11714 (N_11714,N_11465,N_11259);
xor U11715 (N_11715,N_11389,N_11348);
xor U11716 (N_11716,N_11424,N_11412);
nor U11717 (N_11717,N_11377,N_11308);
and U11718 (N_11718,N_11445,N_11394);
xnor U11719 (N_11719,N_11345,N_11279);
nor U11720 (N_11720,N_11487,N_11363);
nor U11721 (N_11721,N_11273,N_11392);
or U11722 (N_11722,N_11328,N_11324);
or U11723 (N_11723,N_11406,N_11279);
nor U11724 (N_11724,N_11342,N_11354);
nand U11725 (N_11725,N_11479,N_11395);
xnor U11726 (N_11726,N_11255,N_11260);
xnor U11727 (N_11727,N_11495,N_11361);
nand U11728 (N_11728,N_11470,N_11465);
nor U11729 (N_11729,N_11373,N_11262);
and U11730 (N_11730,N_11463,N_11347);
xor U11731 (N_11731,N_11463,N_11471);
and U11732 (N_11732,N_11306,N_11316);
nand U11733 (N_11733,N_11293,N_11251);
and U11734 (N_11734,N_11284,N_11482);
and U11735 (N_11735,N_11413,N_11498);
nand U11736 (N_11736,N_11440,N_11496);
nand U11737 (N_11737,N_11448,N_11355);
nand U11738 (N_11738,N_11432,N_11428);
nand U11739 (N_11739,N_11269,N_11495);
or U11740 (N_11740,N_11448,N_11384);
xnor U11741 (N_11741,N_11319,N_11323);
nand U11742 (N_11742,N_11258,N_11416);
xnor U11743 (N_11743,N_11303,N_11275);
nand U11744 (N_11744,N_11447,N_11482);
and U11745 (N_11745,N_11421,N_11317);
nor U11746 (N_11746,N_11426,N_11393);
nor U11747 (N_11747,N_11480,N_11453);
xnor U11748 (N_11748,N_11347,N_11458);
and U11749 (N_11749,N_11336,N_11347);
xnor U11750 (N_11750,N_11579,N_11540);
xor U11751 (N_11751,N_11680,N_11641);
and U11752 (N_11752,N_11590,N_11719);
and U11753 (N_11753,N_11543,N_11520);
xnor U11754 (N_11754,N_11708,N_11621);
or U11755 (N_11755,N_11599,N_11516);
nand U11756 (N_11756,N_11729,N_11630);
nor U11757 (N_11757,N_11613,N_11502);
xor U11758 (N_11758,N_11545,N_11702);
nand U11759 (N_11759,N_11727,N_11669);
and U11760 (N_11760,N_11660,N_11577);
xor U11761 (N_11761,N_11721,N_11527);
nor U11762 (N_11762,N_11512,N_11560);
and U11763 (N_11763,N_11564,N_11732);
or U11764 (N_11764,N_11639,N_11553);
xor U11765 (N_11765,N_11746,N_11651);
xor U11766 (N_11766,N_11503,N_11602);
nor U11767 (N_11767,N_11521,N_11685);
and U11768 (N_11768,N_11723,N_11622);
or U11769 (N_11769,N_11508,N_11556);
or U11770 (N_11770,N_11552,N_11569);
nor U11771 (N_11771,N_11519,N_11698);
and U11772 (N_11772,N_11705,N_11598);
and U11773 (N_11773,N_11734,N_11709);
or U11774 (N_11774,N_11667,N_11584);
and U11775 (N_11775,N_11696,N_11653);
nand U11776 (N_11776,N_11693,N_11506);
and U11777 (N_11777,N_11731,N_11583);
and U11778 (N_11778,N_11593,N_11601);
xor U11779 (N_11779,N_11666,N_11627);
and U11780 (N_11780,N_11715,N_11511);
or U11781 (N_11781,N_11554,N_11718);
xnor U11782 (N_11782,N_11636,N_11739);
nand U11783 (N_11783,N_11532,N_11604);
or U11784 (N_11784,N_11572,N_11624);
nor U11785 (N_11785,N_11657,N_11597);
xnor U11786 (N_11786,N_11720,N_11518);
and U11787 (N_11787,N_11717,N_11534);
and U11788 (N_11788,N_11699,N_11595);
and U11789 (N_11789,N_11672,N_11644);
and U11790 (N_11790,N_11629,N_11513);
and U11791 (N_11791,N_11529,N_11741);
nand U11792 (N_11792,N_11707,N_11634);
or U11793 (N_11793,N_11649,N_11711);
xor U11794 (N_11794,N_11663,N_11500);
nand U11795 (N_11795,N_11716,N_11647);
xnor U11796 (N_11796,N_11738,N_11735);
and U11797 (N_11797,N_11697,N_11524);
and U11798 (N_11798,N_11631,N_11536);
nor U11799 (N_11799,N_11539,N_11625);
nand U11800 (N_11800,N_11571,N_11740);
xnor U11801 (N_11801,N_11588,N_11676);
or U11802 (N_11802,N_11578,N_11736);
nor U11803 (N_11803,N_11606,N_11600);
nor U11804 (N_11804,N_11563,N_11704);
or U11805 (N_11805,N_11550,N_11690);
xor U11806 (N_11806,N_11743,N_11561);
and U11807 (N_11807,N_11677,N_11575);
nor U11808 (N_11808,N_11659,N_11562);
or U11809 (N_11809,N_11632,N_11642);
and U11810 (N_11810,N_11603,N_11558);
xnor U11811 (N_11811,N_11725,N_11522);
or U11812 (N_11812,N_11538,N_11733);
nand U11813 (N_11813,N_11684,N_11713);
or U11814 (N_11814,N_11694,N_11637);
or U11815 (N_11815,N_11565,N_11611);
or U11816 (N_11816,N_11581,N_11594);
or U11817 (N_11817,N_11566,N_11555);
and U11818 (N_11818,N_11635,N_11692);
or U11819 (N_11819,N_11643,N_11510);
xor U11820 (N_11820,N_11744,N_11609);
nand U11821 (N_11821,N_11618,N_11655);
nor U11822 (N_11822,N_11526,N_11547);
nor U11823 (N_11823,N_11724,N_11691);
and U11824 (N_11824,N_11514,N_11530);
nand U11825 (N_11825,N_11658,N_11747);
nor U11826 (N_11826,N_11652,N_11670);
xnor U11827 (N_11827,N_11589,N_11681);
or U11828 (N_11828,N_11714,N_11674);
nor U11829 (N_11829,N_11585,N_11706);
and U11830 (N_11830,N_11608,N_11531);
or U11831 (N_11831,N_11591,N_11537);
or U11832 (N_11832,N_11648,N_11619);
nand U11833 (N_11833,N_11745,N_11712);
xnor U11834 (N_11834,N_11551,N_11682);
nand U11835 (N_11835,N_11504,N_11687);
nand U11836 (N_11836,N_11546,N_11722);
nand U11837 (N_11837,N_11665,N_11749);
or U11838 (N_11838,N_11661,N_11501);
nor U11839 (N_11839,N_11616,N_11615);
or U11840 (N_11840,N_11576,N_11568);
and U11841 (N_11841,N_11626,N_11640);
xor U11842 (N_11842,N_11535,N_11656);
nor U11843 (N_11843,N_11737,N_11573);
nand U11844 (N_11844,N_11528,N_11505);
nand U11845 (N_11845,N_11675,N_11683);
nor U11846 (N_11846,N_11517,N_11596);
xor U11847 (N_11847,N_11668,N_11620);
nand U11848 (N_11848,N_11549,N_11580);
and U11849 (N_11849,N_11662,N_11703);
and U11850 (N_11850,N_11582,N_11525);
nor U11851 (N_11851,N_11650,N_11586);
and U11852 (N_11852,N_11614,N_11567);
xor U11853 (N_11853,N_11507,N_11509);
xnor U11854 (N_11854,N_11574,N_11607);
and U11855 (N_11855,N_11688,N_11592);
nand U11856 (N_11856,N_11617,N_11628);
and U11857 (N_11857,N_11610,N_11664);
xor U11858 (N_11858,N_11689,N_11523);
or U11859 (N_11859,N_11605,N_11559);
and U11860 (N_11860,N_11544,N_11686);
nor U11861 (N_11861,N_11623,N_11515);
nand U11862 (N_11862,N_11679,N_11742);
xnor U11863 (N_11863,N_11678,N_11638);
and U11864 (N_11864,N_11748,N_11673);
nand U11865 (N_11865,N_11728,N_11645);
or U11866 (N_11866,N_11726,N_11587);
nand U11867 (N_11867,N_11700,N_11695);
nor U11868 (N_11868,N_11570,N_11701);
and U11869 (N_11869,N_11533,N_11671);
nand U11870 (N_11870,N_11654,N_11612);
xor U11871 (N_11871,N_11542,N_11710);
and U11872 (N_11872,N_11541,N_11633);
xor U11873 (N_11873,N_11557,N_11646);
nor U11874 (N_11874,N_11730,N_11548);
or U11875 (N_11875,N_11603,N_11587);
and U11876 (N_11876,N_11717,N_11730);
or U11877 (N_11877,N_11736,N_11741);
and U11878 (N_11878,N_11514,N_11644);
xor U11879 (N_11879,N_11674,N_11509);
nor U11880 (N_11880,N_11651,N_11673);
and U11881 (N_11881,N_11567,N_11560);
and U11882 (N_11882,N_11561,N_11642);
nand U11883 (N_11883,N_11664,N_11605);
nor U11884 (N_11884,N_11745,N_11509);
nor U11885 (N_11885,N_11683,N_11712);
or U11886 (N_11886,N_11693,N_11555);
nor U11887 (N_11887,N_11665,N_11530);
nor U11888 (N_11888,N_11523,N_11732);
xor U11889 (N_11889,N_11683,N_11568);
nor U11890 (N_11890,N_11554,N_11709);
xnor U11891 (N_11891,N_11526,N_11590);
xor U11892 (N_11892,N_11677,N_11606);
nor U11893 (N_11893,N_11526,N_11675);
or U11894 (N_11894,N_11583,N_11664);
or U11895 (N_11895,N_11596,N_11566);
nand U11896 (N_11896,N_11704,N_11529);
or U11897 (N_11897,N_11579,N_11595);
and U11898 (N_11898,N_11720,N_11744);
nand U11899 (N_11899,N_11531,N_11627);
and U11900 (N_11900,N_11593,N_11560);
xnor U11901 (N_11901,N_11746,N_11674);
and U11902 (N_11902,N_11534,N_11549);
xnor U11903 (N_11903,N_11559,N_11729);
xor U11904 (N_11904,N_11579,N_11561);
nand U11905 (N_11905,N_11728,N_11737);
or U11906 (N_11906,N_11602,N_11500);
nor U11907 (N_11907,N_11683,N_11690);
and U11908 (N_11908,N_11732,N_11569);
xnor U11909 (N_11909,N_11602,N_11577);
nor U11910 (N_11910,N_11530,N_11575);
nor U11911 (N_11911,N_11640,N_11610);
nand U11912 (N_11912,N_11700,N_11657);
and U11913 (N_11913,N_11621,N_11714);
nor U11914 (N_11914,N_11651,N_11669);
nor U11915 (N_11915,N_11671,N_11511);
nand U11916 (N_11916,N_11558,N_11642);
nand U11917 (N_11917,N_11533,N_11515);
and U11918 (N_11918,N_11527,N_11573);
nor U11919 (N_11919,N_11615,N_11544);
or U11920 (N_11920,N_11724,N_11655);
xnor U11921 (N_11921,N_11711,N_11600);
xnor U11922 (N_11922,N_11626,N_11720);
xnor U11923 (N_11923,N_11540,N_11599);
nor U11924 (N_11924,N_11530,N_11709);
nand U11925 (N_11925,N_11717,N_11710);
nand U11926 (N_11926,N_11535,N_11573);
nand U11927 (N_11927,N_11543,N_11602);
nand U11928 (N_11928,N_11701,N_11722);
xnor U11929 (N_11929,N_11596,N_11634);
nor U11930 (N_11930,N_11749,N_11573);
or U11931 (N_11931,N_11680,N_11571);
xor U11932 (N_11932,N_11691,N_11677);
nor U11933 (N_11933,N_11590,N_11745);
nor U11934 (N_11934,N_11510,N_11527);
and U11935 (N_11935,N_11525,N_11688);
xor U11936 (N_11936,N_11699,N_11719);
nor U11937 (N_11937,N_11746,N_11585);
or U11938 (N_11938,N_11660,N_11746);
nand U11939 (N_11939,N_11525,N_11529);
or U11940 (N_11940,N_11624,N_11582);
xor U11941 (N_11941,N_11747,N_11727);
xor U11942 (N_11942,N_11723,N_11698);
nor U11943 (N_11943,N_11707,N_11708);
and U11944 (N_11944,N_11743,N_11603);
and U11945 (N_11945,N_11641,N_11651);
xor U11946 (N_11946,N_11598,N_11540);
xor U11947 (N_11947,N_11748,N_11745);
and U11948 (N_11948,N_11725,N_11575);
nand U11949 (N_11949,N_11748,N_11678);
or U11950 (N_11950,N_11706,N_11652);
or U11951 (N_11951,N_11518,N_11744);
and U11952 (N_11952,N_11746,N_11583);
xor U11953 (N_11953,N_11711,N_11574);
and U11954 (N_11954,N_11575,N_11706);
and U11955 (N_11955,N_11632,N_11571);
nor U11956 (N_11956,N_11718,N_11704);
or U11957 (N_11957,N_11536,N_11553);
nor U11958 (N_11958,N_11504,N_11580);
nand U11959 (N_11959,N_11634,N_11665);
xor U11960 (N_11960,N_11514,N_11574);
nor U11961 (N_11961,N_11674,N_11527);
xor U11962 (N_11962,N_11511,N_11590);
nor U11963 (N_11963,N_11673,N_11632);
or U11964 (N_11964,N_11592,N_11635);
nand U11965 (N_11965,N_11558,N_11528);
xor U11966 (N_11966,N_11630,N_11542);
and U11967 (N_11967,N_11578,N_11619);
xor U11968 (N_11968,N_11534,N_11683);
or U11969 (N_11969,N_11661,N_11629);
nand U11970 (N_11970,N_11749,N_11540);
xor U11971 (N_11971,N_11561,N_11571);
or U11972 (N_11972,N_11742,N_11739);
nand U11973 (N_11973,N_11680,N_11572);
nand U11974 (N_11974,N_11566,N_11617);
or U11975 (N_11975,N_11592,N_11586);
nor U11976 (N_11976,N_11573,N_11634);
nor U11977 (N_11977,N_11542,N_11599);
nand U11978 (N_11978,N_11656,N_11651);
nand U11979 (N_11979,N_11511,N_11748);
xnor U11980 (N_11980,N_11617,N_11625);
xnor U11981 (N_11981,N_11634,N_11519);
and U11982 (N_11982,N_11586,N_11698);
nand U11983 (N_11983,N_11518,N_11714);
xor U11984 (N_11984,N_11584,N_11652);
nand U11985 (N_11985,N_11519,N_11660);
and U11986 (N_11986,N_11654,N_11589);
or U11987 (N_11987,N_11531,N_11719);
and U11988 (N_11988,N_11575,N_11736);
nand U11989 (N_11989,N_11616,N_11507);
nand U11990 (N_11990,N_11539,N_11723);
xor U11991 (N_11991,N_11648,N_11589);
and U11992 (N_11992,N_11570,N_11687);
nor U11993 (N_11993,N_11745,N_11582);
nand U11994 (N_11994,N_11739,N_11543);
and U11995 (N_11995,N_11735,N_11538);
nor U11996 (N_11996,N_11735,N_11675);
nand U11997 (N_11997,N_11661,N_11512);
and U11998 (N_11998,N_11578,N_11595);
xnor U11999 (N_11999,N_11528,N_11531);
nor U12000 (N_12000,N_11753,N_11770);
and U12001 (N_12001,N_11956,N_11940);
or U12002 (N_12002,N_11835,N_11979);
xnor U12003 (N_12003,N_11988,N_11978);
or U12004 (N_12004,N_11761,N_11769);
nor U12005 (N_12005,N_11793,N_11885);
or U12006 (N_12006,N_11759,N_11865);
nor U12007 (N_12007,N_11965,N_11797);
xnor U12008 (N_12008,N_11851,N_11928);
or U12009 (N_12009,N_11828,N_11839);
or U12010 (N_12010,N_11868,N_11934);
and U12011 (N_12011,N_11813,N_11869);
nor U12012 (N_12012,N_11833,N_11768);
or U12013 (N_12013,N_11888,N_11808);
xnor U12014 (N_12014,N_11872,N_11779);
and U12015 (N_12015,N_11774,N_11765);
xnor U12016 (N_12016,N_11800,N_11908);
xnor U12017 (N_12017,N_11792,N_11817);
xor U12018 (N_12018,N_11931,N_11947);
xnor U12019 (N_12019,N_11789,N_11751);
or U12020 (N_12020,N_11767,N_11829);
nor U12021 (N_12021,N_11998,N_11983);
nor U12022 (N_12022,N_11843,N_11757);
xor U12023 (N_12023,N_11944,N_11857);
and U12024 (N_12024,N_11899,N_11790);
and U12025 (N_12025,N_11805,N_11912);
and U12026 (N_12026,N_11926,N_11943);
and U12027 (N_12027,N_11838,N_11891);
xnor U12028 (N_12028,N_11796,N_11905);
nor U12029 (N_12029,N_11830,N_11989);
and U12030 (N_12030,N_11848,N_11810);
nor U12031 (N_12031,N_11977,N_11860);
nand U12032 (N_12032,N_11879,N_11918);
or U12033 (N_12033,N_11780,N_11952);
or U12034 (N_12034,N_11936,N_11837);
and U12035 (N_12035,N_11787,N_11754);
xnor U12036 (N_12036,N_11875,N_11786);
and U12037 (N_12037,N_11882,N_11795);
or U12038 (N_12038,N_11816,N_11913);
and U12039 (N_12039,N_11844,N_11784);
xor U12040 (N_12040,N_11832,N_11907);
nand U12041 (N_12041,N_11880,N_11971);
nand U12042 (N_12042,N_11929,N_11866);
nor U12043 (N_12043,N_11763,N_11846);
nand U12044 (N_12044,N_11783,N_11871);
nand U12045 (N_12045,N_11893,N_11897);
xor U12046 (N_12046,N_11752,N_11812);
nand U12047 (N_12047,N_11903,N_11930);
and U12048 (N_12048,N_11889,N_11847);
and U12049 (N_12049,N_11982,N_11827);
and U12050 (N_12050,N_11772,N_11775);
xor U12051 (N_12051,N_11996,N_11831);
nand U12052 (N_12052,N_11953,N_11973);
nor U12053 (N_12053,N_11802,N_11821);
and U12054 (N_12054,N_11852,N_11994);
nand U12055 (N_12055,N_11845,N_11886);
nor U12056 (N_12056,N_11840,N_11807);
nand U12057 (N_12057,N_11895,N_11858);
xor U12058 (N_12058,N_11898,N_11777);
nand U12059 (N_12059,N_11937,N_11764);
and U12060 (N_12060,N_11874,N_11932);
xnor U12061 (N_12061,N_11778,N_11966);
nor U12062 (N_12062,N_11986,N_11801);
or U12063 (N_12063,N_11890,N_11924);
nand U12064 (N_12064,N_11750,N_11849);
nor U12065 (N_12065,N_11922,N_11963);
nor U12066 (N_12066,N_11902,N_11993);
nand U12067 (N_12067,N_11948,N_11804);
nor U12068 (N_12068,N_11799,N_11864);
nand U12069 (N_12069,N_11946,N_11818);
and U12070 (N_12070,N_11949,N_11938);
nor U12071 (N_12071,N_11809,N_11856);
xor U12072 (N_12072,N_11758,N_11927);
nor U12073 (N_12073,N_11841,N_11755);
or U12074 (N_12074,N_11883,N_11803);
and U12075 (N_12075,N_11760,N_11788);
nand U12076 (N_12076,N_11798,N_11862);
or U12077 (N_12077,N_11878,N_11962);
nor U12078 (N_12078,N_11811,N_11861);
xnor U12079 (N_12079,N_11776,N_11873);
and U12080 (N_12080,N_11959,N_11853);
nand U12081 (N_12081,N_11781,N_11967);
or U12082 (N_12082,N_11914,N_11990);
and U12083 (N_12083,N_11855,N_11824);
nor U12084 (N_12084,N_11999,N_11911);
and U12085 (N_12085,N_11919,N_11909);
and U12086 (N_12086,N_11773,N_11794);
xnor U12087 (N_12087,N_11976,N_11762);
nor U12088 (N_12088,N_11921,N_11910);
nand U12089 (N_12089,N_11820,N_11863);
and U12090 (N_12090,N_11917,N_11870);
or U12091 (N_12091,N_11819,N_11960);
nand U12092 (N_12092,N_11859,N_11969);
or U12093 (N_12093,N_11854,N_11904);
nor U12094 (N_12094,N_11901,N_11935);
nor U12095 (N_12095,N_11877,N_11997);
nor U12096 (N_12096,N_11925,N_11972);
and U12097 (N_12097,N_11887,N_11964);
nor U12098 (N_12098,N_11942,N_11842);
nor U12099 (N_12099,N_11881,N_11850);
nand U12100 (N_12100,N_11958,N_11991);
and U12101 (N_12101,N_11923,N_11981);
and U12102 (N_12102,N_11980,N_11915);
and U12103 (N_12103,N_11995,N_11834);
xnor U12104 (N_12104,N_11826,N_11815);
nor U12105 (N_12105,N_11876,N_11896);
xor U12106 (N_12106,N_11892,N_11933);
nand U12107 (N_12107,N_11771,N_11791);
nor U12108 (N_12108,N_11825,N_11985);
or U12109 (N_12109,N_11968,N_11955);
nor U12110 (N_12110,N_11984,N_11884);
and U12111 (N_12111,N_11782,N_11785);
and U12112 (N_12112,N_11836,N_11822);
or U12113 (N_12113,N_11950,N_11939);
and U12114 (N_12114,N_11957,N_11941);
xor U12115 (N_12115,N_11900,N_11951);
xor U12116 (N_12116,N_11987,N_11974);
nand U12117 (N_12117,N_11806,N_11970);
xnor U12118 (N_12118,N_11992,N_11945);
or U12119 (N_12119,N_11916,N_11894);
nor U12120 (N_12120,N_11906,N_11961);
and U12121 (N_12121,N_11766,N_11975);
and U12122 (N_12122,N_11814,N_11920);
nor U12123 (N_12123,N_11954,N_11756);
xnor U12124 (N_12124,N_11823,N_11867);
nor U12125 (N_12125,N_11814,N_11939);
nand U12126 (N_12126,N_11897,N_11942);
or U12127 (N_12127,N_11777,N_11976);
or U12128 (N_12128,N_11871,N_11823);
and U12129 (N_12129,N_11952,N_11923);
nor U12130 (N_12130,N_11753,N_11911);
xor U12131 (N_12131,N_11962,N_11795);
xor U12132 (N_12132,N_11892,N_11768);
or U12133 (N_12133,N_11982,N_11879);
and U12134 (N_12134,N_11838,N_11983);
xor U12135 (N_12135,N_11802,N_11990);
or U12136 (N_12136,N_11922,N_11935);
and U12137 (N_12137,N_11923,N_11768);
and U12138 (N_12138,N_11852,N_11982);
and U12139 (N_12139,N_11813,N_11816);
nor U12140 (N_12140,N_11877,N_11843);
and U12141 (N_12141,N_11816,N_11885);
and U12142 (N_12142,N_11786,N_11761);
xnor U12143 (N_12143,N_11920,N_11800);
xnor U12144 (N_12144,N_11811,N_11842);
nor U12145 (N_12145,N_11938,N_11752);
and U12146 (N_12146,N_11792,N_11831);
nor U12147 (N_12147,N_11887,N_11888);
nor U12148 (N_12148,N_11927,N_11970);
nor U12149 (N_12149,N_11811,N_11911);
or U12150 (N_12150,N_11815,N_11823);
nand U12151 (N_12151,N_11851,N_11779);
xnor U12152 (N_12152,N_11883,N_11896);
nor U12153 (N_12153,N_11858,N_11801);
and U12154 (N_12154,N_11763,N_11750);
nand U12155 (N_12155,N_11968,N_11919);
nand U12156 (N_12156,N_11781,N_11825);
nand U12157 (N_12157,N_11799,N_11846);
or U12158 (N_12158,N_11947,N_11914);
nand U12159 (N_12159,N_11822,N_11799);
xnor U12160 (N_12160,N_11977,N_11951);
and U12161 (N_12161,N_11801,N_11883);
or U12162 (N_12162,N_11868,N_11958);
xor U12163 (N_12163,N_11759,N_11935);
xor U12164 (N_12164,N_11899,N_11772);
nand U12165 (N_12165,N_11808,N_11991);
nor U12166 (N_12166,N_11881,N_11792);
xor U12167 (N_12167,N_11783,N_11906);
or U12168 (N_12168,N_11758,N_11944);
nor U12169 (N_12169,N_11791,N_11829);
nand U12170 (N_12170,N_11775,N_11884);
and U12171 (N_12171,N_11772,N_11971);
and U12172 (N_12172,N_11759,N_11962);
xor U12173 (N_12173,N_11777,N_11954);
and U12174 (N_12174,N_11781,N_11834);
nand U12175 (N_12175,N_11887,N_11806);
xnor U12176 (N_12176,N_11929,N_11973);
or U12177 (N_12177,N_11834,N_11964);
nor U12178 (N_12178,N_11997,N_11788);
and U12179 (N_12179,N_11796,N_11834);
nand U12180 (N_12180,N_11882,N_11937);
and U12181 (N_12181,N_11864,N_11840);
xnor U12182 (N_12182,N_11984,N_11826);
xnor U12183 (N_12183,N_11951,N_11856);
nand U12184 (N_12184,N_11857,N_11967);
xor U12185 (N_12185,N_11798,N_11951);
xor U12186 (N_12186,N_11841,N_11968);
or U12187 (N_12187,N_11896,N_11799);
or U12188 (N_12188,N_11898,N_11977);
xor U12189 (N_12189,N_11877,N_11766);
nand U12190 (N_12190,N_11822,N_11888);
nor U12191 (N_12191,N_11934,N_11924);
nor U12192 (N_12192,N_11859,N_11908);
nor U12193 (N_12193,N_11950,N_11911);
nand U12194 (N_12194,N_11772,N_11877);
or U12195 (N_12195,N_11978,N_11981);
xor U12196 (N_12196,N_11894,N_11994);
nor U12197 (N_12197,N_11960,N_11962);
nand U12198 (N_12198,N_11984,N_11765);
nor U12199 (N_12199,N_11861,N_11750);
and U12200 (N_12200,N_11952,N_11906);
nor U12201 (N_12201,N_11768,N_11970);
xor U12202 (N_12202,N_11771,N_11818);
or U12203 (N_12203,N_11928,N_11884);
and U12204 (N_12204,N_11841,N_11986);
xor U12205 (N_12205,N_11798,N_11857);
or U12206 (N_12206,N_11960,N_11874);
xor U12207 (N_12207,N_11912,N_11953);
or U12208 (N_12208,N_11920,N_11906);
or U12209 (N_12209,N_11954,N_11959);
nor U12210 (N_12210,N_11971,N_11893);
nand U12211 (N_12211,N_11976,N_11782);
nor U12212 (N_12212,N_11761,N_11815);
and U12213 (N_12213,N_11922,N_11964);
or U12214 (N_12214,N_11884,N_11942);
nor U12215 (N_12215,N_11994,N_11983);
xnor U12216 (N_12216,N_11928,N_11768);
xnor U12217 (N_12217,N_11979,N_11859);
and U12218 (N_12218,N_11821,N_11811);
and U12219 (N_12219,N_11842,N_11999);
and U12220 (N_12220,N_11994,N_11836);
or U12221 (N_12221,N_11758,N_11940);
nor U12222 (N_12222,N_11909,N_11971);
and U12223 (N_12223,N_11805,N_11797);
nor U12224 (N_12224,N_11964,N_11852);
or U12225 (N_12225,N_11772,N_11837);
or U12226 (N_12226,N_11929,N_11902);
nand U12227 (N_12227,N_11889,N_11893);
nand U12228 (N_12228,N_11750,N_11907);
xnor U12229 (N_12229,N_11961,N_11902);
and U12230 (N_12230,N_11893,N_11821);
xor U12231 (N_12231,N_11834,N_11993);
and U12232 (N_12232,N_11859,N_11840);
nor U12233 (N_12233,N_11876,N_11957);
nor U12234 (N_12234,N_11861,N_11838);
nand U12235 (N_12235,N_11775,N_11789);
nor U12236 (N_12236,N_11981,N_11851);
xor U12237 (N_12237,N_11883,N_11982);
xnor U12238 (N_12238,N_11767,N_11879);
nor U12239 (N_12239,N_11828,N_11989);
xor U12240 (N_12240,N_11963,N_11843);
nand U12241 (N_12241,N_11831,N_11810);
xnor U12242 (N_12242,N_11900,N_11798);
nor U12243 (N_12243,N_11769,N_11771);
xor U12244 (N_12244,N_11948,N_11899);
or U12245 (N_12245,N_11997,N_11863);
and U12246 (N_12246,N_11916,N_11763);
or U12247 (N_12247,N_11785,N_11857);
and U12248 (N_12248,N_11949,N_11998);
and U12249 (N_12249,N_11867,N_11860);
nand U12250 (N_12250,N_12098,N_12221);
nor U12251 (N_12251,N_12132,N_12207);
and U12252 (N_12252,N_12162,N_12151);
and U12253 (N_12253,N_12057,N_12002);
and U12254 (N_12254,N_12133,N_12109);
or U12255 (N_12255,N_12099,N_12239);
or U12256 (N_12256,N_12247,N_12001);
or U12257 (N_12257,N_12120,N_12061);
or U12258 (N_12258,N_12153,N_12148);
xor U12259 (N_12259,N_12198,N_12249);
and U12260 (N_12260,N_12145,N_12228);
or U12261 (N_12261,N_12222,N_12027);
nor U12262 (N_12262,N_12155,N_12178);
or U12263 (N_12263,N_12204,N_12106);
nor U12264 (N_12264,N_12059,N_12067);
nor U12265 (N_12265,N_12058,N_12236);
nand U12266 (N_12266,N_12179,N_12063);
and U12267 (N_12267,N_12248,N_12122);
and U12268 (N_12268,N_12044,N_12140);
nor U12269 (N_12269,N_12097,N_12081);
or U12270 (N_12270,N_12074,N_12226);
xnor U12271 (N_12271,N_12144,N_12124);
and U12272 (N_12272,N_12128,N_12108);
or U12273 (N_12273,N_12232,N_12216);
nor U12274 (N_12274,N_12012,N_12125);
xor U12275 (N_12275,N_12242,N_12009);
nand U12276 (N_12276,N_12079,N_12220);
nand U12277 (N_12277,N_12011,N_12191);
and U12278 (N_12278,N_12215,N_12028);
nand U12279 (N_12279,N_12161,N_12157);
nor U12280 (N_12280,N_12025,N_12233);
nand U12281 (N_12281,N_12101,N_12126);
nand U12282 (N_12282,N_12017,N_12034);
xnor U12283 (N_12283,N_12013,N_12189);
nor U12284 (N_12284,N_12091,N_12150);
or U12285 (N_12285,N_12167,N_12010);
nand U12286 (N_12286,N_12104,N_12203);
xnor U12287 (N_12287,N_12054,N_12165);
xor U12288 (N_12288,N_12187,N_12042);
or U12289 (N_12289,N_12018,N_12168);
xor U12290 (N_12290,N_12114,N_12019);
nand U12291 (N_12291,N_12246,N_12070);
or U12292 (N_12292,N_12209,N_12135);
xor U12293 (N_12293,N_12107,N_12041);
or U12294 (N_12294,N_12053,N_12075);
xor U12295 (N_12295,N_12038,N_12095);
or U12296 (N_12296,N_12181,N_12229);
xnor U12297 (N_12297,N_12142,N_12036);
or U12298 (N_12298,N_12238,N_12100);
nor U12299 (N_12299,N_12152,N_12193);
or U12300 (N_12300,N_12194,N_12078);
nand U12301 (N_12301,N_12048,N_12113);
or U12302 (N_12302,N_12211,N_12050);
xnor U12303 (N_12303,N_12082,N_12139);
nand U12304 (N_12304,N_12062,N_12197);
nand U12305 (N_12305,N_12234,N_12171);
nor U12306 (N_12306,N_12087,N_12088);
nor U12307 (N_12307,N_12093,N_12185);
and U12308 (N_12308,N_12219,N_12068);
xor U12309 (N_12309,N_12066,N_12123);
or U12310 (N_12310,N_12035,N_12000);
nand U12311 (N_12311,N_12031,N_12170);
and U12312 (N_12312,N_12046,N_12173);
xor U12313 (N_12313,N_12083,N_12240);
and U12314 (N_12314,N_12172,N_12092);
nand U12315 (N_12315,N_12130,N_12213);
and U12316 (N_12316,N_12147,N_12024);
nor U12317 (N_12317,N_12014,N_12205);
xnor U12318 (N_12318,N_12201,N_12032);
nor U12319 (N_12319,N_12119,N_12192);
xor U12320 (N_12320,N_12055,N_12177);
and U12321 (N_12321,N_12143,N_12243);
and U12322 (N_12322,N_12129,N_12040);
nand U12323 (N_12323,N_12137,N_12105);
nand U12324 (N_12324,N_12015,N_12127);
nor U12325 (N_12325,N_12073,N_12195);
and U12326 (N_12326,N_12094,N_12005);
nor U12327 (N_12327,N_12188,N_12004);
xor U12328 (N_12328,N_12186,N_12200);
nand U12329 (N_12329,N_12116,N_12118);
nand U12330 (N_12330,N_12245,N_12065);
or U12331 (N_12331,N_12047,N_12111);
xnor U12332 (N_12332,N_12131,N_12069);
xnor U12333 (N_12333,N_12225,N_12149);
xnor U12334 (N_12334,N_12214,N_12023);
or U12335 (N_12335,N_12096,N_12159);
nand U12336 (N_12336,N_12103,N_12235);
nand U12337 (N_12337,N_12208,N_12230);
nor U12338 (N_12338,N_12086,N_12174);
nand U12339 (N_12339,N_12026,N_12085);
nand U12340 (N_12340,N_12180,N_12072);
or U12341 (N_12341,N_12206,N_12182);
nand U12342 (N_12342,N_12064,N_12029);
or U12343 (N_12343,N_12154,N_12084);
or U12344 (N_12344,N_12231,N_12110);
nor U12345 (N_12345,N_12102,N_12089);
nor U12346 (N_12346,N_12056,N_12244);
nor U12347 (N_12347,N_12016,N_12224);
nor U12348 (N_12348,N_12223,N_12164);
and U12349 (N_12349,N_12146,N_12077);
nand U12350 (N_12350,N_12210,N_12022);
xnor U12351 (N_12351,N_12033,N_12212);
xnor U12352 (N_12352,N_12169,N_12166);
nor U12353 (N_12353,N_12196,N_12052);
xnor U12354 (N_12354,N_12136,N_12134);
nor U12355 (N_12355,N_12003,N_12060);
nand U12356 (N_12356,N_12043,N_12080);
nor U12357 (N_12357,N_12020,N_12039);
and U12358 (N_12358,N_12199,N_12202);
or U12359 (N_12359,N_12008,N_12183);
xnor U12360 (N_12360,N_12158,N_12006);
or U12361 (N_12361,N_12076,N_12190);
and U12362 (N_12362,N_12112,N_12115);
nor U12363 (N_12363,N_12141,N_12049);
and U12364 (N_12364,N_12007,N_12176);
and U12365 (N_12365,N_12030,N_12218);
or U12366 (N_12366,N_12184,N_12163);
nor U12367 (N_12367,N_12160,N_12121);
and U12368 (N_12368,N_12071,N_12227);
nand U12369 (N_12369,N_12156,N_12241);
nor U12370 (N_12370,N_12021,N_12217);
and U12371 (N_12371,N_12117,N_12090);
nor U12372 (N_12372,N_12175,N_12037);
nor U12373 (N_12373,N_12237,N_12051);
or U12374 (N_12374,N_12138,N_12045);
or U12375 (N_12375,N_12192,N_12023);
or U12376 (N_12376,N_12174,N_12115);
nand U12377 (N_12377,N_12066,N_12183);
or U12378 (N_12378,N_12168,N_12117);
nor U12379 (N_12379,N_12122,N_12228);
nor U12380 (N_12380,N_12064,N_12105);
xor U12381 (N_12381,N_12023,N_12184);
nand U12382 (N_12382,N_12166,N_12236);
or U12383 (N_12383,N_12070,N_12193);
nor U12384 (N_12384,N_12021,N_12086);
or U12385 (N_12385,N_12012,N_12183);
and U12386 (N_12386,N_12196,N_12121);
and U12387 (N_12387,N_12113,N_12237);
nor U12388 (N_12388,N_12033,N_12167);
nor U12389 (N_12389,N_12240,N_12077);
xor U12390 (N_12390,N_12141,N_12003);
nand U12391 (N_12391,N_12064,N_12013);
and U12392 (N_12392,N_12222,N_12103);
or U12393 (N_12393,N_12240,N_12102);
nand U12394 (N_12394,N_12044,N_12207);
or U12395 (N_12395,N_12074,N_12047);
nor U12396 (N_12396,N_12239,N_12002);
xnor U12397 (N_12397,N_12072,N_12074);
nor U12398 (N_12398,N_12075,N_12184);
and U12399 (N_12399,N_12158,N_12031);
and U12400 (N_12400,N_12011,N_12070);
nor U12401 (N_12401,N_12154,N_12225);
xor U12402 (N_12402,N_12109,N_12208);
or U12403 (N_12403,N_12059,N_12064);
or U12404 (N_12404,N_12193,N_12132);
xnor U12405 (N_12405,N_12157,N_12052);
and U12406 (N_12406,N_12003,N_12138);
and U12407 (N_12407,N_12127,N_12038);
nor U12408 (N_12408,N_12208,N_12202);
xor U12409 (N_12409,N_12241,N_12042);
nor U12410 (N_12410,N_12005,N_12123);
nor U12411 (N_12411,N_12089,N_12199);
or U12412 (N_12412,N_12204,N_12087);
nor U12413 (N_12413,N_12224,N_12135);
or U12414 (N_12414,N_12168,N_12161);
xnor U12415 (N_12415,N_12034,N_12102);
nor U12416 (N_12416,N_12090,N_12194);
nand U12417 (N_12417,N_12232,N_12009);
nand U12418 (N_12418,N_12219,N_12138);
and U12419 (N_12419,N_12028,N_12133);
and U12420 (N_12420,N_12065,N_12145);
nor U12421 (N_12421,N_12139,N_12247);
and U12422 (N_12422,N_12034,N_12109);
nand U12423 (N_12423,N_12049,N_12194);
nor U12424 (N_12424,N_12120,N_12216);
or U12425 (N_12425,N_12092,N_12137);
xnor U12426 (N_12426,N_12055,N_12079);
xnor U12427 (N_12427,N_12016,N_12045);
nand U12428 (N_12428,N_12008,N_12070);
and U12429 (N_12429,N_12085,N_12018);
and U12430 (N_12430,N_12178,N_12089);
and U12431 (N_12431,N_12037,N_12246);
nand U12432 (N_12432,N_12164,N_12200);
nor U12433 (N_12433,N_12022,N_12078);
nand U12434 (N_12434,N_12192,N_12054);
nand U12435 (N_12435,N_12164,N_12054);
xnor U12436 (N_12436,N_12134,N_12118);
nand U12437 (N_12437,N_12069,N_12156);
or U12438 (N_12438,N_12030,N_12067);
or U12439 (N_12439,N_12012,N_12246);
nand U12440 (N_12440,N_12240,N_12243);
xnor U12441 (N_12441,N_12208,N_12081);
and U12442 (N_12442,N_12068,N_12211);
or U12443 (N_12443,N_12067,N_12069);
or U12444 (N_12444,N_12158,N_12063);
nand U12445 (N_12445,N_12229,N_12000);
and U12446 (N_12446,N_12122,N_12042);
or U12447 (N_12447,N_12191,N_12083);
or U12448 (N_12448,N_12104,N_12030);
nor U12449 (N_12449,N_12097,N_12134);
and U12450 (N_12450,N_12213,N_12117);
and U12451 (N_12451,N_12221,N_12067);
and U12452 (N_12452,N_12001,N_12067);
nand U12453 (N_12453,N_12003,N_12171);
or U12454 (N_12454,N_12028,N_12207);
nand U12455 (N_12455,N_12245,N_12068);
or U12456 (N_12456,N_12069,N_12189);
nand U12457 (N_12457,N_12004,N_12223);
or U12458 (N_12458,N_12093,N_12194);
xnor U12459 (N_12459,N_12171,N_12084);
xor U12460 (N_12460,N_12071,N_12069);
or U12461 (N_12461,N_12195,N_12051);
xnor U12462 (N_12462,N_12148,N_12140);
nand U12463 (N_12463,N_12093,N_12212);
or U12464 (N_12464,N_12149,N_12049);
nor U12465 (N_12465,N_12216,N_12005);
and U12466 (N_12466,N_12210,N_12236);
or U12467 (N_12467,N_12025,N_12096);
nor U12468 (N_12468,N_12104,N_12156);
nand U12469 (N_12469,N_12219,N_12046);
nand U12470 (N_12470,N_12066,N_12117);
xor U12471 (N_12471,N_12053,N_12102);
nor U12472 (N_12472,N_12037,N_12181);
and U12473 (N_12473,N_12036,N_12096);
or U12474 (N_12474,N_12239,N_12006);
and U12475 (N_12475,N_12026,N_12087);
and U12476 (N_12476,N_12232,N_12121);
and U12477 (N_12477,N_12112,N_12199);
xnor U12478 (N_12478,N_12055,N_12149);
or U12479 (N_12479,N_12158,N_12164);
or U12480 (N_12480,N_12065,N_12111);
or U12481 (N_12481,N_12026,N_12049);
xnor U12482 (N_12482,N_12168,N_12147);
nor U12483 (N_12483,N_12167,N_12169);
nor U12484 (N_12484,N_12096,N_12151);
xnor U12485 (N_12485,N_12111,N_12248);
nor U12486 (N_12486,N_12013,N_12115);
nand U12487 (N_12487,N_12157,N_12165);
nand U12488 (N_12488,N_12199,N_12224);
or U12489 (N_12489,N_12211,N_12021);
nand U12490 (N_12490,N_12086,N_12033);
xor U12491 (N_12491,N_12160,N_12157);
nor U12492 (N_12492,N_12125,N_12047);
nand U12493 (N_12493,N_12240,N_12193);
and U12494 (N_12494,N_12088,N_12188);
and U12495 (N_12495,N_12105,N_12131);
nor U12496 (N_12496,N_12148,N_12094);
and U12497 (N_12497,N_12134,N_12132);
xnor U12498 (N_12498,N_12169,N_12005);
or U12499 (N_12499,N_12195,N_12049);
or U12500 (N_12500,N_12471,N_12274);
nand U12501 (N_12501,N_12379,N_12383);
or U12502 (N_12502,N_12441,N_12278);
nor U12503 (N_12503,N_12412,N_12391);
or U12504 (N_12504,N_12479,N_12330);
xor U12505 (N_12505,N_12451,N_12254);
nand U12506 (N_12506,N_12499,N_12483);
nor U12507 (N_12507,N_12453,N_12429);
and U12508 (N_12508,N_12469,N_12454);
nor U12509 (N_12509,N_12268,N_12375);
nand U12510 (N_12510,N_12318,N_12283);
nand U12511 (N_12511,N_12310,N_12442);
or U12512 (N_12512,N_12466,N_12365);
or U12513 (N_12513,N_12378,N_12339);
or U12514 (N_12514,N_12397,N_12255);
and U12515 (N_12515,N_12349,N_12486);
and U12516 (N_12516,N_12271,N_12332);
xnor U12517 (N_12517,N_12394,N_12460);
xor U12518 (N_12518,N_12288,N_12298);
nand U12519 (N_12519,N_12273,N_12345);
xnor U12520 (N_12520,N_12449,N_12286);
and U12521 (N_12521,N_12467,N_12348);
xnor U12522 (N_12522,N_12296,N_12389);
nor U12523 (N_12523,N_12494,N_12347);
nor U12524 (N_12524,N_12265,N_12437);
or U12525 (N_12525,N_12300,N_12363);
xor U12526 (N_12526,N_12420,N_12401);
nand U12527 (N_12527,N_12317,N_12481);
nand U12528 (N_12528,N_12251,N_12262);
nand U12529 (N_12529,N_12368,N_12439);
xor U12530 (N_12530,N_12490,N_12353);
xnor U12531 (N_12531,N_12386,N_12455);
xnor U12532 (N_12532,N_12430,N_12484);
xor U12533 (N_12533,N_12334,N_12338);
and U12534 (N_12534,N_12299,N_12470);
nor U12535 (N_12535,N_12281,N_12361);
or U12536 (N_12536,N_12400,N_12417);
xnor U12537 (N_12537,N_12303,N_12457);
and U12538 (N_12538,N_12289,N_12290);
nor U12539 (N_12539,N_12362,N_12293);
nor U12540 (N_12540,N_12392,N_12425);
nand U12541 (N_12541,N_12343,N_12323);
and U12542 (N_12542,N_12277,N_12475);
xor U12543 (N_12543,N_12371,N_12411);
and U12544 (N_12544,N_12450,N_12282);
xnor U12545 (N_12545,N_12419,N_12415);
xor U12546 (N_12546,N_12497,N_12374);
nor U12547 (N_12547,N_12478,N_12344);
and U12548 (N_12548,N_12313,N_12354);
nand U12549 (N_12549,N_12263,N_12301);
and U12550 (N_12550,N_12284,N_12482);
nor U12551 (N_12551,N_12364,N_12459);
nand U12552 (N_12552,N_12440,N_12297);
nand U12553 (N_12553,N_12477,N_12359);
nand U12554 (N_12554,N_12306,N_12285);
nand U12555 (N_12555,N_12385,N_12387);
or U12556 (N_12556,N_12292,N_12452);
xor U12557 (N_12557,N_12433,N_12493);
nor U12558 (N_12558,N_12256,N_12322);
nor U12559 (N_12559,N_12380,N_12464);
nand U12560 (N_12560,N_12473,N_12406);
nor U12561 (N_12561,N_12270,N_12456);
and U12562 (N_12562,N_12404,N_12367);
xor U12563 (N_12563,N_12356,N_12329);
xnor U12564 (N_12564,N_12416,N_12444);
xnor U12565 (N_12565,N_12396,N_12340);
nor U12566 (N_12566,N_12258,N_12408);
nor U12567 (N_12567,N_12461,N_12462);
xor U12568 (N_12568,N_12314,N_12331);
or U12569 (N_12569,N_12266,N_12384);
nor U12570 (N_12570,N_12346,N_12305);
xnor U12571 (N_12571,N_12405,N_12360);
or U12572 (N_12572,N_12259,N_12448);
and U12573 (N_12573,N_12312,N_12370);
and U12574 (N_12574,N_12485,N_12333);
nand U12575 (N_12575,N_12492,N_12381);
nor U12576 (N_12576,N_12491,N_12295);
xor U12577 (N_12577,N_12250,N_12436);
and U12578 (N_12578,N_12434,N_12369);
or U12579 (N_12579,N_12328,N_12341);
xnor U12580 (N_12580,N_12414,N_12324);
and U12581 (N_12581,N_12257,N_12352);
or U12582 (N_12582,N_12319,N_12402);
and U12583 (N_12583,N_12309,N_12327);
nor U12584 (N_12584,N_12468,N_12357);
and U12585 (N_12585,N_12253,N_12432);
or U12586 (N_12586,N_12438,N_12418);
nand U12587 (N_12587,N_12446,N_12428);
nand U12588 (N_12588,N_12315,N_12409);
nand U12589 (N_12589,N_12390,N_12424);
nand U12590 (N_12590,N_12276,N_12373);
nor U12591 (N_12591,N_12423,N_12498);
nand U12592 (N_12592,N_12351,N_12307);
nand U12593 (N_12593,N_12325,N_12465);
nand U12594 (N_12594,N_12337,N_12291);
and U12595 (N_12595,N_12399,N_12311);
nand U12596 (N_12596,N_12316,N_12358);
nor U12597 (N_12597,N_12304,N_12377);
xor U12598 (N_12598,N_12350,N_12435);
nor U12599 (N_12599,N_12280,N_12335);
xor U12600 (N_12600,N_12445,N_12476);
xnor U12601 (N_12601,N_12496,N_12398);
nand U12602 (N_12602,N_12489,N_12407);
or U12603 (N_12603,N_12413,N_12422);
nor U12604 (N_12604,N_12252,N_12443);
nor U12605 (N_12605,N_12463,N_12372);
nor U12606 (N_12606,N_12269,N_12410);
or U12607 (N_12607,N_12487,N_12495);
nor U12608 (N_12608,N_12261,N_12321);
xor U12609 (N_12609,N_12421,N_12447);
nand U12610 (N_12610,N_12488,N_12366);
and U12611 (N_12611,N_12431,N_12260);
nor U12612 (N_12612,N_12272,N_12403);
or U12613 (N_12613,N_12376,N_12474);
and U12614 (N_12614,N_12388,N_12393);
xor U12615 (N_12615,N_12458,N_12320);
xor U12616 (N_12616,N_12275,N_12308);
nand U12617 (N_12617,N_12382,N_12336);
xnor U12618 (N_12618,N_12427,N_12426);
or U12619 (N_12619,N_12355,N_12302);
and U12620 (N_12620,N_12294,N_12287);
or U12621 (N_12621,N_12267,N_12480);
xor U12622 (N_12622,N_12326,N_12264);
xnor U12623 (N_12623,N_12342,N_12279);
or U12624 (N_12624,N_12472,N_12395);
nand U12625 (N_12625,N_12464,N_12310);
xor U12626 (N_12626,N_12343,N_12368);
xnor U12627 (N_12627,N_12300,N_12258);
nor U12628 (N_12628,N_12382,N_12312);
or U12629 (N_12629,N_12467,N_12454);
nand U12630 (N_12630,N_12346,N_12287);
nand U12631 (N_12631,N_12274,N_12255);
and U12632 (N_12632,N_12326,N_12381);
and U12633 (N_12633,N_12370,N_12474);
xor U12634 (N_12634,N_12256,N_12494);
and U12635 (N_12635,N_12269,N_12460);
and U12636 (N_12636,N_12341,N_12293);
nand U12637 (N_12637,N_12475,N_12470);
nand U12638 (N_12638,N_12260,N_12282);
or U12639 (N_12639,N_12347,N_12456);
nand U12640 (N_12640,N_12388,N_12333);
xnor U12641 (N_12641,N_12324,N_12288);
and U12642 (N_12642,N_12270,N_12333);
nor U12643 (N_12643,N_12385,N_12256);
and U12644 (N_12644,N_12345,N_12410);
nand U12645 (N_12645,N_12491,N_12299);
and U12646 (N_12646,N_12330,N_12420);
nand U12647 (N_12647,N_12254,N_12481);
or U12648 (N_12648,N_12406,N_12431);
nand U12649 (N_12649,N_12337,N_12275);
and U12650 (N_12650,N_12408,N_12327);
nor U12651 (N_12651,N_12360,N_12358);
nor U12652 (N_12652,N_12424,N_12291);
nand U12653 (N_12653,N_12349,N_12250);
or U12654 (N_12654,N_12456,N_12388);
and U12655 (N_12655,N_12419,N_12327);
or U12656 (N_12656,N_12356,N_12392);
nand U12657 (N_12657,N_12392,N_12408);
and U12658 (N_12658,N_12295,N_12478);
and U12659 (N_12659,N_12279,N_12419);
xor U12660 (N_12660,N_12472,N_12319);
and U12661 (N_12661,N_12438,N_12309);
nor U12662 (N_12662,N_12381,N_12434);
nand U12663 (N_12663,N_12378,N_12251);
and U12664 (N_12664,N_12356,N_12408);
and U12665 (N_12665,N_12307,N_12258);
or U12666 (N_12666,N_12378,N_12473);
and U12667 (N_12667,N_12348,N_12323);
xnor U12668 (N_12668,N_12317,N_12441);
nor U12669 (N_12669,N_12367,N_12285);
nor U12670 (N_12670,N_12382,N_12479);
nand U12671 (N_12671,N_12411,N_12465);
nand U12672 (N_12672,N_12364,N_12393);
nand U12673 (N_12673,N_12284,N_12297);
xnor U12674 (N_12674,N_12458,N_12383);
and U12675 (N_12675,N_12378,N_12285);
or U12676 (N_12676,N_12251,N_12392);
xor U12677 (N_12677,N_12434,N_12258);
and U12678 (N_12678,N_12466,N_12445);
or U12679 (N_12679,N_12280,N_12271);
or U12680 (N_12680,N_12250,N_12312);
nor U12681 (N_12681,N_12431,N_12350);
or U12682 (N_12682,N_12286,N_12322);
nand U12683 (N_12683,N_12435,N_12474);
and U12684 (N_12684,N_12273,N_12352);
or U12685 (N_12685,N_12326,N_12496);
nor U12686 (N_12686,N_12353,N_12414);
or U12687 (N_12687,N_12255,N_12377);
nor U12688 (N_12688,N_12439,N_12264);
nor U12689 (N_12689,N_12406,N_12459);
xnor U12690 (N_12690,N_12269,N_12371);
or U12691 (N_12691,N_12324,N_12434);
nor U12692 (N_12692,N_12335,N_12305);
xnor U12693 (N_12693,N_12336,N_12437);
nand U12694 (N_12694,N_12337,N_12411);
nand U12695 (N_12695,N_12388,N_12491);
and U12696 (N_12696,N_12379,N_12295);
and U12697 (N_12697,N_12386,N_12494);
or U12698 (N_12698,N_12449,N_12416);
nor U12699 (N_12699,N_12475,N_12340);
nand U12700 (N_12700,N_12328,N_12449);
or U12701 (N_12701,N_12400,N_12438);
nand U12702 (N_12702,N_12277,N_12347);
nand U12703 (N_12703,N_12431,N_12269);
or U12704 (N_12704,N_12262,N_12282);
nor U12705 (N_12705,N_12432,N_12255);
and U12706 (N_12706,N_12398,N_12472);
xnor U12707 (N_12707,N_12466,N_12497);
or U12708 (N_12708,N_12350,N_12334);
xor U12709 (N_12709,N_12410,N_12400);
and U12710 (N_12710,N_12475,N_12420);
nor U12711 (N_12711,N_12468,N_12422);
or U12712 (N_12712,N_12331,N_12393);
xnor U12713 (N_12713,N_12455,N_12474);
or U12714 (N_12714,N_12309,N_12442);
nand U12715 (N_12715,N_12421,N_12411);
nand U12716 (N_12716,N_12393,N_12420);
nor U12717 (N_12717,N_12284,N_12447);
nand U12718 (N_12718,N_12276,N_12372);
or U12719 (N_12719,N_12401,N_12320);
nand U12720 (N_12720,N_12476,N_12352);
xnor U12721 (N_12721,N_12394,N_12455);
or U12722 (N_12722,N_12329,N_12266);
xor U12723 (N_12723,N_12375,N_12489);
nor U12724 (N_12724,N_12409,N_12431);
nand U12725 (N_12725,N_12295,N_12354);
xnor U12726 (N_12726,N_12428,N_12286);
nand U12727 (N_12727,N_12430,N_12432);
nor U12728 (N_12728,N_12495,N_12296);
nor U12729 (N_12729,N_12250,N_12313);
nand U12730 (N_12730,N_12294,N_12443);
xor U12731 (N_12731,N_12486,N_12404);
and U12732 (N_12732,N_12313,N_12492);
and U12733 (N_12733,N_12459,N_12354);
and U12734 (N_12734,N_12326,N_12278);
xnor U12735 (N_12735,N_12314,N_12444);
xnor U12736 (N_12736,N_12328,N_12271);
xnor U12737 (N_12737,N_12382,N_12388);
nand U12738 (N_12738,N_12350,N_12277);
nand U12739 (N_12739,N_12487,N_12298);
nor U12740 (N_12740,N_12270,N_12321);
nor U12741 (N_12741,N_12442,N_12330);
or U12742 (N_12742,N_12389,N_12293);
and U12743 (N_12743,N_12295,N_12439);
or U12744 (N_12744,N_12349,N_12432);
and U12745 (N_12745,N_12452,N_12338);
xnor U12746 (N_12746,N_12383,N_12288);
or U12747 (N_12747,N_12370,N_12473);
or U12748 (N_12748,N_12387,N_12367);
nand U12749 (N_12749,N_12318,N_12413);
or U12750 (N_12750,N_12702,N_12587);
or U12751 (N_12751,N_12692,N_12675);
and U12752 (N_12752,N_12589,N_12636);
and U12753 (N_12753,N_12501,N_12654);
and U12754 (N_12754,N_12632,N_12672);
xnor U12755 (N_12755,N_12720,N_12540);
xor U12756 (N_12756,N_12542,N_12509);
nand U12757 (N_12757,N_12610,N_12717);
or U12758 (N_12758,N_12665,N_12521);
nor U12759 (N_12759,N_12684,N_12531);
or U12760 (N_12760,N_12555,N_12732);
or U12761 (N_12761,N_12549,N_12663);
and U12762 (N_12762,N_12507,N_12627);
nor U12763 (N_12763,N_12749,N_12538);
nand U12764 (N_12764,N_12524,N_12546);
and U12765 (N_12765,N_12686,N_12506);
or U12766 (N_12766,N_12747,N_12646);
xor U12767 (N_12767,N_12705,N_12680);
xnor U12768 (N_12768,N_12709,N_12510);
and U12769 (N_12769,N_12676,N_12593);
nor U12770 (N_12770,N_12631,N_12609);
xnor U12771 (N_12771,N_12508,N_12505);
or U12772 (N_12772,N_12569,N_12607);
nand U12773 (N_12773,N_12550,N_12625);
nand U12774 (N_12774,N_12583,N_12710);
and U12775 (N_12775,N_12635,N_12662);
nor U12776 (N_12776,N_12623,N_12746);
or U12777 (N_12777,N_12580,N_12595);
and U12778 (N_12778,N_12726,N_12643);
xnor U12779 (N_12779,N_12700,N_12500);
and U12780 (N_12780,N_12685,N_12703);
or U12781 (N_12781,N_12577,N_12718);
xor U12782 (N_12782,N_12641,N_12563);
xor U12783 (N_12783,N_12677,N_12669);
and U12784 (N_12784,N_12698,N_12748);
nand U12785 (N_12785,N_12644,N_12565);
or U12786 (N_12786,N_12503,N_12727);
or U12787 (N_12787,N_12708,N_12648);
and U12788 (N_12788,N_12597,N_12733);
and U12789 (N_12789,N_12602,N_12551);
and U12790 (N_12790,N_12659,N_12530);
nor U12791 (N_12791,N_12573,N_12670);
and U12792 (N_12792,N_12539,N_12529);
and U12793 (N_12793,N_12557,N_12712);
or U12794 (N_12794,N_12650,N_12574);
xor U12795 (N_12795,N_12729,N_12624);
nor U12796 (N_12796,N_12516,N_12628);
or U12797 (N_12797,N_12590,N_12598);
and U12798 (N_12798,N_12730,N_12585);
nand U12799 (N_12799,N_12566,N_12601);
xor U12800 (N_12800,N_12608,N_12562);
and U12801 (N_12801,N_12745,N_12515);
nor U12802 (N_12802,N_12679,N_12738);
nand U12803 (N_12803,N_12618,N_12630);
nor U12804 (N_12804,N_12548,N_12527);
and U12805 (N_12805,N_12649,N_12605);
and U12806 (N_12806,N_12570,N_12737);
or U12807 (N_12807,N_12532,N_12525);
and U12808 (N_12808,N_12558,N_12523);
xor U12809 (N_12809,N_12575,N_12547);
nor U12810 (N_12810,N_12504,N_12571);
xor U12811 (N_12811,N_12743,N_12701);
xnor U12812 (N_12812,N_12613,N_12656);
xor U12813 (N_12813,N_12617,N_12731);
and U12814 (N_12814,N_12728,N_12576);
nand U12815 (N_12815,N_12658,N_12689);
nand U12816 (N_12816,N_12704,N_12722);
nor U12817 (N_12817,N_12707,N_12604);
and U12818 (N_12818,N_12713,N_12661);
nand U12819 (N_12819,N_12678,N_12638);
xnor U12820 (N_12820,N_12626,N_12706);
nor U12821 (N_12821,N_12611,N_12652);
nand U12822 (N_12822,N_12572,N_12541);
nand U12823 (N_12823,N_12714,N_12544);
nor U12824 (N_12824,N_12511,N_12647);
or U12825 (N_12825,N_12579,N_12554);
nand U12826 (N_12826,N_12696,N_12581);
and U12827 (N_12827,N_12568,N_12517);
nor U12828 (N_12828,N_12711,N_12616);
nor U12829 (N_12829,N_12526,N_12560);
xnor U12830 (N_12830,N_12543,N_12519);
and U12831 (N_12831,N_12592,N_12674);
xor U12832 (N_12832,N_12619,N_12633);
or U12833 (N_12833,N_12528,N_12629);
nand U12834 (N_12834,N_12584,N_12742);
and U12835 (N_12835,N_12682,N_12596);
xnor U12836 (N_12836,N_12520,N_12578);
xor U12837 (N_12837,N_12673,N_12522);
nand U12838 (N_12838,N_12734,N_12721);
nor U12839 (N_12839,N_12620,N_12561);
or U12840 (N_12840,N_12588,N_12657);
nor U12841 (N_12841,N_12699,N_12645);
xor U12842 (N_12842,N_12668,N_12671);
xnor U12843 (N_12843,N_12683,N_12518);
nand U12844 (N_12844,N_12514,N_12599);
nor U12845 (N_12845,N_12739,N_12655);
and U12846 (N_12846,N_12612,N_12637);
xnor U12847 (N_12847,N_12664,N_12552);
or U12848 (N_12848,N_12639,N_12614);
and U12849 (N_12849,N_12693,N_12735);
or U12850 (N_12850,N_12537,N_12603);
and U12851 (N_12851,N_12513,N_12640);
nor U12852 (N_12852,N_12690,N_12667);
nand U12853 (N_12853,N_12606,N_12688);
xnor U12854 (N_12854,N_12564,N_12559);
xnor U12855 (N_12855,N_12653,N_12694);
and U12856 (N_12856,N_12651,N_12536);
or U12857 (N_12857,N_12586,N_12642);
nand U12858 (N_12858,N_12545,N_12744);
or U12859 (N_12859,N_12533,N_12582);
and U12860 (N_12860,N_12594,N_12621);
nor U12861 (N_12861,N_12622,N_12567);
nor U12862 (N_12862,N_12600,N_12719);
nor U12863 (N_12863,N_12725,N_12591);
xnor U12864 (N_12864,N_12740,N_12534);
and U12865 (N_12865,N_12634,N_12715);
and U12866 (N_12866,N_12553,N_12736);
nand U12867 (N_12867,N_12681,N_12723);
or U12868 (N_12868,N_12512,N_12666);
xor U12869 (N_12869,N_12660,N_12687);
nand U12870 (N_12870,N_12697,N_12724);
nand U12871 (N_12871,N_12691,N_12535);
xor U12872 (N_12872,N_12716,N_12502);
and U12873 (N_12873,N_12741,N_12556);
or U12874 (N_12874,N_12615,N_12695);
xnor U12875 (N_12875,N_12571,N_12586);
nor U12876 (N_12876,N_12551,N_12521);
nor U12877 (N_12877,N_12712,N_12612);
or U12878 (N_12878,N_12576,N_12596);
or U12879 (N_12879,N_12731,N_12641);
and U12880 (N_12880,N_12615,N_12731);
and U12881 (N_12881,N_12744,N_12730);
or U12882 (N_12882,N_12744,N_12542);
xnor U12883 (N_12883,N_12608,N_12705);
and U12884 (N_12884,N_12712,N_12539);
nor U12885 (N_12885,N_12555,N_12659);
xnor U12886 (N_12886,N_12526,N_12638);
nand U12887 (N_12887,N_12542,N_12685);
nor U12888 (N_12888,N_12621,N_12538);
or U12889 (N_12889,N_12538,N_12530);
nand U12890 (N_12890,N_12647,N_12629);
nor U12891 (N_12891,N_12695,N_12525);
or U12892 (N_12892,N_12727,N_12526);
nor U12893 (N_12893,N_12570,N_12537);
nor U12894 (N_12894,N_12656,N_12504);
and U12895 (N_12895,N_12698,N_12559);
nor U12896 (N_12896,N_12709,N_12555);
nor U12897 (N_12897,N_12625,N_12627);
or U12898 (N_12898,N_12511,N_12704);
and U12899 (N_12899,N_12654,N_12719);
or U12900 (N_12900,N_12706,N_12503);
or U12901 (N_12901,N_12608,N_12688);
and U12902 (N_12902,N_12544,N_12505);
nor U12903 (N_12903,N_12664,N_12640);
nor U12904 (N_12904,N_12693,N_12514);
nor U12905 (N_12905,N_12674,N_12668);
or U12906 (N_12906,N_12652,N_12696);
nand U12907 (N_12907,N_12707,N_12586);
nor U12908 (N_12908,N_12619,N_12666);
xor U12909 (N_12909,N_12586,N_12523);
nor U12910 (N_12910,N_12710,N_12659);
xor U12911 (N_12911,N_12635,N_12542);
or U12912 (N_12912,N_12717,N_12604);
xnor U12913 (N_12913,N_12678,N_12674);
nor U12914 (N_12914,N_12629,N_12564);
nand U12915 (N_12915,N_12746,N_12512);
xor U12916 (N_12916,N_12657,N_12713);
nor U12917 (N_12917,N_12677,N_12547);
xnor U12918 (N_12918,N_12667,N_12508);
or U12919 (N_12919,N_12508,N_12719);
nor U12920 (N_12920,N_12559,N_12500);
nor U12921 (N_12921,N_12596,N_12580);
or U12922 (N_12922,N_12592,N_12678);
xnor U12923 (N_12923,N_12645,N_12579);
or U12924 (N_12924,N_12546,N_12624);
or U12925 (N_12925,N_12641,N_12723);
and U12926 (N_12926,N_12627,N_12512);
xnor U12927 (N_12927,N_12581,N_12623);
xor U12928 (N_12928,N_12639,N_12621);
xor U12929 (N_12929,N_12532,N_12598);
nor U12930 (N_12930,N_12683,N_12723);
and U12931 (N_12931,N_12579,N_12667);
or U12932 (N_12932,N_12694,N_12644);
nor U12933 (N_12933,N_12548,N_12748);
nor U12934 (N_12934,N_12659,N_12577);
or U12935 (N_12935,N_12536,N_12512);
or U12936 (N_12936,N_12722,N_12713);
nand U12937 (N_12937,N_12603,N_12688);
nor U12938 (N_12938,N_12708,N_12600);
nor U12939 (N_12939,N_12681,N_12684);
and U12940 (N_12940,N_12553,N_12727);
nor U12941 (N_12941,N_12544,N_12582);
and U12942 (N_12942,N_12577,N_12614);
nand U12943 (N_12943,N_12636,N_12634);
or U12944 (N_12944,N_12513,N_12518);
nand U12945 (N_12945,N_12744,N_12746);
nor U12946 (N_12946,N_12680,N_12615);
or U12947 (N_12947,N_12626,N_12515);
xnor U12948 (N_12948,N_12623,N_12684);
nor U12949 (N_12949,N_12681,N_12589);
xnor U12950 (N_12950,N_12594,N_12550);
nor U12951 (N_12951,N_12700,N_12699);
xnor U12952 (N_12952,N_12574,N_12539);
xnor U12953 (N_12953,N_12501,N_12504);
nor U12954 (N_12954,N_12627,N_12545);
and U12955 (N_12955,N_12610,N_12670);
xnor U12956 (N_12956,N_12712,N_12601);
xor U12957 (N_12957,N_12556,N_12576);
xnor U12958 (N_12958,N_12515,N_12643);
xor U12959 (N_12959,N_12729,N_12684);
or U12960 (N_12960,N_12640,N_12641);
and U12961 (N_12961,N_12644,N_12540);
nand U12962 (N_12962,N_12500,N_12674);
nor U12963 (N_12963,N_12619,N_12531);
or U12964 (N_12964,N_12605,N_12693);
and U12965 (N_12965,N_12574,N_12742);
or U12966 (N_12966,N_12646,N_12637);
or U12967 (N_12967,N_12602,N_12711);
xnor U12968 (N_12968,N_12726,N_12617);
nor U12969 (N_12969,N_12537,N_12580);
and U12970 (N_12970,N_12671,N_12576);
nor U12971 (N_12971,N_12728,N_12704);
nor U12972 (N_12972,N_12631,N_12621);
nand U12973 (N_12973,N_12704,N_12741);
or U12974 (N_12974,N_12705,N_12610);
nand U12975 (N_12975,N_12542,N_12615);
nor U12976 (N_12976,N_12562,N_12628);
or U12977 (N_12977,N_12584,N_12707);
and U12978 (N_12978,N_12532,N_12610);
or U12979 (N_12979,N_12692,N_12731);
and U12980 (N_12980,N_12687,N_12688);
and U12981 (N_12981,N_12590,N_12640);
or U12982 (N_12982,N_12586,N_12628);
nand U12983 (N_12983,N_12710,N_12682);
and U12984 (N_12984,N_12616,N_12625);
xor U12985 (N_12985,N_12595,N_12539);
xnor U12986 (N_12986,N_12595,N_12563);
nand U12987 (N_12987,N_12704,N_12611);
and U12988 (N_12988,N_12579,N_12604);
nor U12989 (N_12989,N_12605,N_12616);
nand U12990 (N_12990,N_12504,N_12578);
or U12991 (N_12991,N_12731,N_12655);
and U12992 (N_12992,N_12591,N_12547);
nand U12993 (N_12993,N_12749,N_12537);
xnor U12994 (N_12994,N_12566,N_12556);
nor U12995 (N_12995,N_12519,N_12639);
nor U12996 (N_12996,N_12749,N_12571);
or U12997 (N_12997,N_12542,N_12663);
nor U12998 (N_12998,N_12694,N_12680);
or U12999 (N_12999,N_12571,N_12746);
and U13000 (N_13000,N_12989,N_12826);
or U13001 (N_13001,N_12787,N_12872);
nor U13002 (N_13002,N_12788,N_12860);
or U13003 (N_13003,N_12897,N_12928);
nand U13004 (N_13004,N_12770,N_12804);
nand U13005 (N_13005,N_12895,N_12923);
nand U13006 (N_13006,N_12870,N_12906);
xor U13007 (N_13007,N_12853,N_12818);
and U13008 (N_13008,N_12988,N_12884);
nor U13009 (N_13009,N_12773,N_12842);
nand U13010 (N_13010,N_12756,N_12807);
or U13011 (N_13011,N_12806,N_12900);
nor U13012 (N_13012,N_12801,N_12789);
nor U13013 (N_13013,N_12793,N_12820);
or U13014 (N_13014,N_12994,N_12968);
or U13015 (N_13015,N_12758,N_12769);
nor U13016 (N_13016,N_12963,N_12930);
or U13017 (N_13017,N_12786,N_12780);
nand U13018 (N_13018,N_12991,N_12812);
nor U13019 (N_13019,N_12799,N_12905);
xor U13020 (N_13020,N_12976,N_12840);
or U13021 (N_13021,N_12848,N_12760);
and U13022 (N_13022,N_12800,N_12847);
and U13023 (N_13023,N_12816,N_12855);
xnor U13024 (N_13024,N_12899,N_12885);
and U13025 (N_13025,N_12782,N_12997);
nand U13026 (N_13026,N_12886,N_12857);
nor U13027 (N_13027,N_12887,N_12859);
nand U13028 (N_13028,N_12829,N_12942);
and U13029 (N_13029,N_12998,N_12992);
nor U13030 (N_13030,N_12843,N_12791);
and U13031 (N_13031,N_12827,N_12817);
nand U13032 (N_13032,N_12766,N_12919);
nor U13033 (N_13033,N_12865,N_12830);
xnor U13034 (N_13034,N_12935,N_12759);
xor U13035 (N_13035,N_12875,N_12888);
nand U13036 (N_13036,N_12783,N_12985);
nor U13037 (N_13037,N_12752,N_12776);
or U13038 (N_13038,N_12951,N_12965);
xnor U13039 (N_13039,N_12937,N_12771);
xor U13040 (N_13040,N_12993,N_12933);
and U13041 (N_13041,N_12784,N_12983);
nand U13042 (N_13042,N_12863,N_12894);
nand U13043 (N_13043,N_12972,N_12819);
or U13044 (N_13044,N_12955,N_12854);
nand U13045 (N_13045,N_12957,N_12938);
xnor U13046 (N_13046,N_12845,N_12889);
nand U13047 (N_13047,N_12896,N_12802);
nand U13048 (N_13048,N_12912,N_12844);
or U13049 (N_13049,N_12798,N_12932);
nand U13050 (N_13050,N_12967,N_12914);
nor U13051 (N_13051,N_12908,N_12765);
xor U13052 (N_13052,N_12809,N_12892);
or U13053 (N_13053,N_12980,N_12846);
and U13054 (N_13054,N_12902,N_12867);
xnor U13055 (N_13055,N_12987,N_12813);
nor U13056 (N_13056,N_12977,N_12757);
xnor U13057 (N_13057,N_12975,N_12946);
nor U13058 (N_13058,N_12768,N_12831);
or U13059 (N_13059,N_12891,N_12861);
and U13060 (N_13060,N_12962,N_12936);
xnor U13061 (N_13061,N_12909,N_12934);
nand U13062 (N_13062,N_12881,N_12856);
or U13063 (N_13063,N_12956,N_12971);
nand U13064 (N_13064,N_12838,N_12918);
or U13065 (N_13065,N_12832,N_12879);
xor U13066 (N_13066,N_12970,N_12949);
xnor U13067 (N_13067,N_12959,N_12915);
nand U13068 (N_13068,N_12778,N_12822);
and U13069 (N_13069,N_12810,N_12940);
nand U13070 (N_13070,N_12903,N_12849);
xor U13071 (N_13071,N_12958,N_12877);
or U13072 (N_13072,N_12767,N_12808);
or U13073 (N_13073,N_12952,N_12961);
nand U13074 (N_13074,N_12753,N_12794);
or U13075 (N_13075,N_12911,N_12834);
nand U13076 (N_13076,N_12871,N_12839);
or U13077 (N_13077,N_12841,N_12969);
nor U13078 (N_13078,N_12796,N_12904);
nor U13079 (N_13079,N_12797,N_12751);
nand U13080 (N_13080,N_12945,N_12907);
or U13081 (N_13081,N_12851,N_12772);
or U13082 (N_13082,N_12823,N_12790);
and U13083 (N_13083,N_12922,N_12775);
or U13084 (N_13084,N_12974,N_12984);
xor U13085 (N_13085,N_12943,N_12835);
or U13086 (N_13086,N_12948,N_12795);
or U13087 (N_13087,N_12837,N_12916);
and U13088 (N_13088,N_12866,N_12755);
or U13089 (N_13089,N_12921,N_12982);
xnor U13090 (N_13090,N_12927,N_12990);
nor U13091 (N_13091,N_12792,N_12939);
nand U13092 (N_13092,N_12876,N_12874);
nor U13093 (N_13093,N_12883,N_12750);
or U13094 (N_13094,N_12805,N_12864);
xor U13095 (N_13095,N_12869,N_12761);
nand U13096 (N_13096,N_12978,N_12890);
nor U13097 (N_13097,N_12996,N_12941);
or U13098 (N_13098,N_12824,N_12777);
or U13099 (N_13099,N_12763,N_12828);
and U13100 (N_13100,N_12858,N_12924);
nand U13101 (N_13101,N_12901,N_12960);
xnor U13102 (N_13102,N_12913,N_12925);
xor U13103 (N_13103,N_12779,N_12815);
or U13104 (N_13104,N_12898,N_12882);
xnor U13105 (N_13105,N_12931,N_12878);
nor U13106 (N_13106,N_12833,N_12814);
nor U13107 (N_13107,N_12917,N_12999);
nor U13108 (N_13108,N_12862,N_12873);
and U13109 (N_13109,N_12986,N_12950);
or U13110 (N_13110,N_12774,N_12852);
or U13111 (N_13111,N_12910,N_12825);
or U13112 (N_13112,N_12821,N_12785);
nor U13113 (N_13113,N_12764,N_12981);
xnor U13114 (N_13114,N_12966,N_12803);
and U13115 (N_13115,N_12920,N_12836);
nor U13116 (N_13116,N_12893,N_12954);
and U13117 (N_13117,N_12868,N_12944);
nor U13118 (N_13118,N_12953,N_12781);
nand U13119 (N_13119,N_12762,N_12754);
nand U13120 (N_13120,N_12964,N_12880);
or U13121 (N_13121,N_12811,N_12995);
xnor U13122 (N_13122,N_12947,N_12850);
nor U13123 (N_13123,N_12926,N_12973);
nand U13124 (N_13124,N_12979,N_12929);
and U13125 (N_13125,N_12787,N_12896);
nand U13126 (N_13126,N_12948,N_12778);
nand U13127 (N_13127,N_12848,N_12927);
nor U13128 (N_13128,N_12940,N_12876);
xor U13129 (N_13129,N_12924,N_12822);
nand U13130 (N_13130,N_12781,N_12925);
xnor U13131 (N_13131,N_12759,N_12920);
or U13132 (N_13132,N_12891,N_12992);
or U13133 (N_13133,N_12896,N_12955);
nor U13134 (N_13134,N_12849,N_12806);
xnor U13135 (N_13135,N_12797,N_12850);
xnor U13136 (N_13136,N_12861,N_12882);
or U13137 (N_13137,N_12788,N_12948);
nor U13138 (N_13138,N_12865,N_12884);
or U13139 (N_13139,N_12865,N_12794);
nor U13140 (N_13140,N_12973,N_12837);
and U13141 (N_13141,N_12929,N_12828);
or U13142 (N_13142,N_12857,N_12763);
xor U13143 (N_13143,N_12911,N_12886);
xor U13144 (N_13144,N_12944,N_12801);
nor U13145 (N_13145,N_12862,N_12992);
nand U13146 (N_13146,N_12813,N_12966);
nand U13147 (N_13147,N_12837,N_12967);
nand U13148 (N_13148,N_12833,N_12821);
and U13149 (N_13149,N_12942,N_12926);
and U13150 (N_13150,N_12794,N_12947);
or U13151 (N_13151,N_12754,N_12994);
and U13152 (N_13152,N_12956,N_12792);
xnor U13153 (N_13153,N_12773,N_12877);
nand U13154 (N_13154,N_12766,N_12812);
and U13155 (N_13155,N_12905,N_12923);
xnor U13156 (N_13156,N_12893,N_12853);
xor U13157 (N_13157,N_12781,N_12878);
and U13158 (N_13158,N_12920,N_12977);
or U13159 (N_13159,N_12901,N_12998);
and U13160 (N_13160,N_12758,N_12890);
and U13161 (N_13161,N_12802,N_12835);
and U13162 (N_13162,N_12804,N_12938);
or U13163 (N_13163,N_12914,N_12779);
nand U13164 (N_13164,N_12768,N_12794);
xnor U13165 (N_13165,N_12925,N_12957);
or U13166 (N_13166,N_12809,N_12951);
xnor U13167 (N_13167,N_12890,N_12908);
xor U13168 (N_13168,N_12880,N_12784);
and U13169 (N_13169,N_12916,N_12832);
xnor U13170 (N_13170,N_12804,N_12840);
nor U13171 (N_13171,N_12978,N_12893);
or U13172 (N_13172,N_12941,N_12836);
or U13173 (N_13173,N_12953,N_12777);
nand U13174 (N_13174,N_12765,N_12861);
nor U13175 (N_13175,N_12768,N_12861);
nor U13176 (N_13176,N_12893,N_12770);
xnor U13177 (N_13177,N_12945,N_12806);
and U13178 (N_13178,N_12879,N_12948);
nor U13179 (N_13179,N_12899,N_12751);
xnor U13180 (N_13180,N_12889,N_12967);
or U13181 (N_13181,N_12945,N_12982);
nand U13182 (N_13182,N_12916,N_12799);
xnor U13183 (N_13183,N_12876,N_12819);
and U13184 (N_13184,N_12852,N_12815);
xor U13185 (N_13185,N_12907,N_12983);
nand U13186 (N_13186,N_12899,N_12994);
nand U13187 (N_13187,N_12912,N_12795);
and U13188 (N_13188,N_12752,N_12923);
or U13189 (N_13189,N_12985,N_12924);
xnor U13190 (N_13190,N_12879,N_12858);
nor U13191 (N_13191,N_12754,N_12953);
nor U13192 (N_13192,N_12893,N_12752);
xnor U13193 (N_13193,N_12833,N_12889);
and U13194 (N_13194,N_12846,N_12875);
or U13195 (N_13195,N_12880,N_12918);
nor U13196 (N_13196,N_12893,N_12791);
and U13197 (N_13197,N_12954,N_12876);
xnor U13198 (N_13198,N_12759,N_12812);
nand U13199 (N_13199,N_12883,N_12757);
nor U13200 (N_13200,N_12858,N_12998);
xor U13201 (N_13201,N_12777,N_12776);
and U13202 (N_13202,N_12978,N_12758);
nor U13203 (N_13203,N_12944,N_12786);
nand U13204 (N_13204,N_12775,N_12971);
xnor U13205 (N_13205,N_12864,N_12794);
and U13206 (N_13206,N_12759,N_12975);
nor U13207 (N_13207,N_12781,N_12831);
nor U13208 (N_13208,N_12872,N_12835);
nand U13209 (N_13209,N_12822,N_12766);
nor U13210 (N_13210,N_12943,N_12782);
or U13211 (N_13211,N_12772,N_12895);
nor U13212 (N_13212,N_12806,N_12938);
nand U13213 (N_13213,N_12801,N_12761);
or U13214 (N_13214,N_12913,N_12906);
or U13215 (N_13215,N_12903,N_12926);
nand U13216 (N_13216,N_12946,N_12926);
and U13217 (N_13217,N_12857,N_12851);
xnor U13218 (N_13218,N_12850,N_12756);
and U13219 (N_13219,N_12810,N_12944);
xnor U13220 (N_13220,N_12934,N_12992);
xor U13221 (N_13221,N_12929,N_12987);
nand U13222 (N_13222,N_12810,N_12771);
and U13223 (N_13223,N_12897,N_12751);
nand U13224 (N_13224,N_12942,N_12880);
nand U13225 (N_13225,N_12904,N_12935);
and U13226 (N_13226,N_12945,N_12926);
nand U13227 (N_13227,N_12896,N_12991);
and U13228 (N_13228,N_12889,N_12974);
and U13229 (N_13229,N_12835,N_12874);
nor U13230 (N_13230,N_12779,N_12859);
or U13231 (N_13231,N_12848,N_12940);
and U13232 (N_13232,N_12962,N_12978);
or U13233 (N_13233,N_12923,N_12872);
and U13234 (N_13234,N_12971,N_12819);
nand U13235 (N_13235,N_12752,N_12797);
nor U13236 (N_13236,N_12997,N_12952);
nand U13237 (N_13237,N_12808,N_12792);
xnor U13238 (N_13238,N_12753,N_12969);
and U13239 (N_13239,N_12959,N_12753);
nand U13240 (N_13240,N_12844,N_12978);
nor U13241 (N_13241,N_12909,N_12782);
nor U13242 (N_13242,N_12783,N_12755);
xor U13243 (N_13243,N_12811,N_12976);
or U13244 (N_13244,N_12915,N_12890);
nand U13245 (N_13245,N_12937,N_12780);
or U13246 (N_13246,N_12936,N_12755);
and U13247 (N_13247,N_12857,N_12906);
nor U13248 (N_13248,N_12766,N_12764);
nor U13249 (N_13249,N_12995,N_12983);
nor U13250 (N_13250,N_13194,N_13192);
xor U13251 (N_13251,N_13066,N_13189);
or U13252 (N_13252,N_13226,N_13090);
and U13253 (N_13253,N_13195,N_13114);
and U13254 (N_13254,N_13115,N_13024);
nand U13255 (N_13255,N_13096,N_13142);
nand U13256 (N_13256,N_13130,N_13073);
nand U13257 (N_13257,N_13235,N_13008);
and U13258 (N_13258,N_13206,N_13244);
xor U13259 (N_13259,N_13182,N_13205);
or U13260 (N_13260,N_13029,N_13001);
and U13261 (N_13261,N_13157,N_13062);
nand U13262 (N_13262,N_13025,N_13187);
xor U13263 (N_13263,N_13148,N_13119);
xor U13264 (N_13264,N_13241,N_13232);
nand U13265 (N_13265,N_13043,N_13067);
and U13266 (N_13266,N_13080,N_13211);
nand U13267 (N_13267,N_13199,N_13221);
nand U13268 (N_13268,N_13028,N_13057);
nand U13269 (N_13269,N_13129,N_13107);
nand U13270 (N_13270,N_13046,N_13230);
nor U13271 (N_13271,N_13179,N_13095);
nor U13272 (N_13272,N_13237,N_13166);
and U13273 (N_13273,N_13003,N_13089);
nand U13274 (N_13274,N_13208,N_13063);
xnor U13275 (N_13275,N_13030,N_13105);
and U13276 (N_13276,N_13151,N_13204);
xnor U13277 (N_13277,N_13200,N_13035);
nor U13278 (N_13278,N_13170,N_13069);
and U13279 (N_13279,N_13156,N_13233);
nand U13280 (N_13280,N_13249,N_13087);
and U13281 (N_13281,N_13054,N_13188);
or U13282 (N_13282,N_13219,N_13123);
xor U13283 (N_13283,N_13047,N_13141);
nand U13284 (N_13284,N_13143,N_13092);
or U13285 (N_13285,N_13122,N_13190);
xor U13286 (N_13286,N_13136,N_13088);
nand U13287 (N_13287,N_13059,N_13071);
nand U13288 (N_13288,N_13017,N_13217);
or U13289 (N_13289,N_13106,N_13239);
or U13290 (N_13290,N_13060,N_13038);
xnor U13291 (N_13291,N_13076,N_13074);
and U13292 (N_13292,N_13197,N_13031);
or U13293 (N_13293,N_13155,N_13091);
nor U13294 (N_13294,N_13004,N_13149);
xnor U13295 (N_13295,N_13049,N_13061);
or U13296 (N_13296,N_13083,N_13150);
xnor U13297 (N_13297,N_13234,N_13118);
nand U13298 (N_13298,N_13011,N_13135);
xnor U13299 (N_13299,N_13174,N_13128);
and U13300 (N_13300,N_13176,N_13227);
xnor U13301 (N_13301,N_13116,N_13094);
nand U13302 (N_13302,N_13140,N_13229);
nand U13303 (N_13303,N_13222,N_13243);
xor U13304 (N_13304,N_13218,N_13099);
and U13305 (N_13305,N_13223,N_13103);
xnor U13306 (N_13306,N_13006,N_13125);
xor U13307 (N_13307,N_13186,N_13220);
or U13308 (N_13308,N_13145,N_13027);
nor U13309 (N_13309,N_13183,N_13042);
xor U13310 (N_13310,N_13064,N_13247);
nand U13311 (N_13311,N_13098,N_13033);
nand U13312 (N_13312,N_13100,N_13133);
and U13313 (N_13313,N_13079,N_13026);
and U13314 (N_13314,N_13065,N_13007);
and U13315 (N_13315,N_13245,N_13172);
nor U13316 (N_13316,N_13044,N_13022);
nand U13317 (N_13317,N_13160,N_13191);
or U13318 (N_13318,N_13154,N_13178);
or U13319 (N_13319,N_13153,N_13162);
and U13320 (N_13320,N_13020,N_13147);
and U13321 (N_13321,N_13146,N_13216);
nor U13322 (N_13322,N_13051,N_13037);
nor U13323 (N_13323,N_13198,N_13055);
nor U13324 (N_13324,N_13039,N_13112);
nand U13325 (N_13325,N_13126,N_13048);
nor U13326 (N_13326,N_13212,N_13132);
nor U13327 (N_13327,N_13165,N_13248);
nor U13328 (N_13328,N_13196,N_13159);
and U13329 (N_13329,N_13019,N_13209);
or U13330 (N_13330,N_13203,N_13109);
nor U13331 (N_13331,N_13131,N_13097);
xnor U13332 (N_13332,N_13181,N_13213);
and U13333 (N_13333,N_13201,N_13193);
nor U13334 (N_13334,N_13000,N_13163);
nand U13335 (N_13335,N_13078,N_13108);
and U13336 (N_13336,N_13127,N_13168);
nand U13337 (N_13337,N_13246,N_13238);
and U13338 (N_13338,N_13075,N_13036);
nor U13339 (N_13339,N_13225,N_13012);
nand U13340 (N_13340,N_13034,N_13040);
xnor U13341 (N_13341,N_13242,N_13158);
nor U13342 (N_13342,N_13185,N_13041);
nand U13343 (N_13343,N_13152,N_13137);
xor U13344 (N_13344,N_13082,N_13010);
nor U13345 (N_13345,N_13032,N_13228);
or U13346 (N_13346,N_13124,N_13139);
nand U13347 (N_13347,N_13093,N_13111);
nand U13348 (N_13348,N_13053,N_13023);
nand U13349 (N_13349,N_13052,N_13173);
xor U13350 (N_13350,N_13144,N_13117);
xnor U13351 (N_13351,N_13215,N_13014);
or U13352 (N_13352,N_13102,N_13171);
nor U13353 (N_13353,N_13016,N_13070);
or U13354 (N_13354,N_13120,N_13005);
and U13355 (N_13355,N_13207,N_13077);
xnor U13356 (N_13356,N_13013,N_13184);
or U13357 (N_13357,N_13085,N_13002);
and U13358 (N_13358,N_13021,N_13101);
nand U13359 (N_13359,N_13134,N_13086);
xnor U13360 (N_13360,N_13202,N_13072);
xnor U13361 (N_13361,N_13121,N_13169);
nand U13362 (N_13362,N_13068,N_13081);
or U13363 (N_13363,N_13240,N_13113);
xnor U13364 (N_13364,N_13236,N_13056);
or U13365 (N_13365,N_13177,N_13161);
xnor U13366 (N_13366,N_13214,N_13167);
nor U13367 (N_13367,N_13015,N_13138);
and U13368 (N_13368,N_13210,N_13104);
or U13369 (N_13369,N_13050,N_13045);
xnor U13370 (N_13370,N_13175,N_13224);
nand U13371 (N_13371,N_13084,N_13180);
nand U13372 (N_13372,N_13058,N_13231);
nand U13373 (N_13373,N_13009,N_13164);
nand U13374 (N_13374,N_13110,N_13018);
or U13375 (N_13375,N_13156,N_13238);
or U13376 (N_13376,N_13128,N_13125);
or U13377 (N_13377,N_13080,N_13143);
nand U13378 (N_13378,N_13220,N_13109);
and U13379 (N_13379,N_13209,N_13180);
nor U13380 (N_13380,N_13083,N_13129);
nand U13381 (N_13381,N_13168,N_13184);
nor U13382 (N_13382,N_13050,N_13026);
xor U13383 (N_13383,N_13042,N_13134);
nor U13384 (N_13384,N_13244,N_13122);
nor U13385 (N_13385,N_13170,N_13135);
xnor U13386 (N_13386,N_13132,N_13196);
and U13387 (N_13387,N_13066,N_13245);
nand U13388 (N_13388,N_13173,N_13229);
nand U13389 (N_13389,N_13130,N_13157);
nand U13390 (N_13390,N_13030,N_13232);
and U13391 (N_13391,N_13195,N_13236);
xor U13392 (N_13392,N_13244,N_13238);
or U13393 (N_13393,N_13047,N_13102);
nor U13394 (N_13394,N_13042,N_13151);
and U13395 (N_13395,N_13136,N_13232);
nor U13396 (N_13396,N_13159,N_13239);
and U13397 (N_13397,N_13245,N_13016);
nor U13398 (N_13398,N_13177,N_13159);
and U13399 (N_13399,N_13149,N_13166);
nor U13400 (N_13400,N_13192,N_13025);
nand U13401 (N_13401,N_13170,N_13092);
nand U13402 (N_13402,N_13079,N_13041);
or U13403 (N_13403,N_13118,N_13012);
nor U13404 (N_13404,N_13080,N_13242);
xnor U13405 (N_13405,N_13107,N_13044);
or U13406 (N_13406,N_13074,N_13228);
nor U13407 (N_13407,N_13006,N_13061);
xnor U13408 (N_13408,N_13098,N_13102);
xnor U13409 (N_13409,N_13147,N_13032);
nand U13410 (N_13410,N_13157,N_13002);
nand U13411 (N_13411,N_13233,N_13226);
and U13412 (N_13412,N_13216,N_13153);
or U13413 (N_13413,N_13184,N_13194);
or U13414 (N_13414,N_13106,N_13235);
nor U13415 (N_13415,N_13115,N_13117);
xor U13416 (N_13416,N_13070,N_13113);
xor U13417 (N_13417,N_13215,N_13247);
xnor U13418 (N_13418,N_13009,N_13001);
xnor U13419 (N_13419,N_13151,N_13248);
nor U13420 (N_13420,N_13211,N_13225);
and U13421 (N_13421,N_13040,N_13136);
nand U13422 (N_13422,N_13022,N_13021);
or U13423 (N_13423,N_13038,N_13023);
xor U13424 (N_13424,N_13019,N_13021);
or U13425 (N_13425,N_13026,N_13078);
nand U13426 (N_13426,N_13168,N_13014);
nor U13427 (N_13427,N_13186,N_13028);
or U13428 (N_13428,N_13117,N_13108);
nand U13429 (N_13429,N_13122,N_13200);
nand U13430 (N_13430,N_13039,N_13207);
and U13431 (N_13431,N_13039,N_13003);
xor U13432 (N_13432,N_13122,N_13192);
xor U13433 (N_13433,N_13131,N_13178);
xor U13434 (N_13434,N_13087,N_13238);
nand U13435 (N_13435,N_13197,N_13071);
and U13436 (N_13436,N_13075,N_13018);
xnor U13437 (N_13437,N_13223,N_13104);
nor U13438 (N_13438,N_13115,N_13125);
and U13439 (N_13439,N_13007,N_13059);
nor U13440 (N_13440,N_13189,N_13103);
nor U13441 (N_13441,N_13202,N_13146);
xor U13442 (N_13442,N_13192,N_13199);
xor U13443 (N_13443,N_13015,N_13206);
nand U13444 (N_13444,N_13193,N_13220);
or U13445 (N_13445,N_13154,N_13240);
nand U13446 (N_13446,N_13109,N_13191);
xnor U13447 (N_13447,N_13080,N_13012);
or U13448 (N_13448,N_13239,N_13062);
and U13449 (N_13449,N_13029,N_13196);
xnor U13450 (N_13450,N_13197,N_13092);
xnor U13451 (N_13451,N_13172,N_13145);
nand U13452 (N_13452,N_13165,N_13082);
or U13453 (N_13453,N_13118,N_13038);
xnor U13454 (N_13454,N_13184,N_13104);
nand U13455 (N_13455,N_13067,N_13176);
xnor U13456 (N_13456,N_13102,N_13105);
nand U13457 (N_13457,N_13004,N_13188);
nand U13458 (N_13458,N_13098,N_13038);
xor U13459 (N_13459,N_13069,N_13065);
xnor U13460 (N_13460,N_13201,N_13182);
xor U13461 (N_13461,N_13077,N_13236);
and U13462 (N_13462,N_13247,N_13087);
or U13463 (N_13463,N_13140,N_13200);
and U13464 (N_13464,N_13030,N_13165);
nand U13465 (N_13465,N_13162,N_13186);
nand U13466 (N_13466,N_13106,N_13053);
nor U13467 (N_13467,N_13092,N_13215);
or U13468 (N_13468,N_13085,N_13138);
nor U13469 (N_13469,N_13087,N_13170);
nand U13470 (N_13470,N_13020,N_13156);
or U13471 (N_13471,N_13242,N_13121);
nand U13472 (N_13472,N_13059,N_13101);
nand U13473 (N_13473,N_13012,N_13214);
or U13474 (N_13474,N_13045,N_13049);
and U13475 (N_13475,N_13031,N_13057);
or U13476 (N_13476,N_13235,N_13197);
nor U13477 (N_13477,N_13034,N_13061);
xnor U13478 (N_13478,N_13210,N_13047);
nand U13479 (N_13479,N_13153,N_13103);
or U13480 (N_13480,N_13007,N_13240);
nor U13481 (N_13481,N_13052,N_13151);
and U13482 (N_13482,N_13083,N_13218);
nor U13483 (N_13483,N_13101,N_13091);
nand U13484 (N_13484,N_13041,N_13170);
nor U13485 (N_13485,N_13247,N_13019);
or U13486 (N_13486,N_13150,N_13214);
nand U13487 (N_13487,N_13014,N_13207);
nand U13488 (N_13488,N_13012,N_13167);
and U13489 (N_13489,N_13203,N_13188);
nor U13490 (N_13490,N_13169,N_13144);
nand U13491 (N_13491,N_13120,N_13246);
nand U13492 (N_13492,N_13171,N_13129);
and U13493 (N_13493,N_13173,N_13109);
nand U13494 (N_13494,N_13021,N_13023);
and U13495 (N_13495,N_13139,N_13224);
and U13496 (N_13496,N_13086,N_13001);
nand U13497 (N_13497,N_13217,N_13141);
nand U13498 (N_13498,N_13219,N_13091);
nor U13499 (N_13499,N_13134,N_13077);
xnor U13500 (N_13500,N_13424,N_13307);
nand U13501 (N_13501,N_13280,N_13378);
or U13502 (N_13502,N_13456,N_13420);
and U13503 (N_13503,N_13435,N_13427);
nor U13504 (N_13504,N_13321,N_13332);
and U13505 (N_13505,N_13309,N_13405);
xnor U13506 (N_13506,N_13319,N_13251);
or U13507 (N_13507,N_13484,N_13411);
or U13508 (N_13508,N_13347,N_13317);
and U13509 (N_13509,N_13440,N_13310);
nand U13510 (N_13510,N_13467,N_13451);
nor U13511 (N_13511,N_13371,N_13489);
nand U13512 (N_13512,N_13461,N_13412);
xor U13513 (N_13513,N_13344,N_13413);
or U13514 (N_13514,N_13318,N_13471);
xor U13515 (N_13515,N_13334,N_13443);
xnor U13516 (N_13516,N_13450,N_13485);
nand U13517 (N_13517,N_13268,N_13491);
and U13518 (N_13518,N_13480,N_13335);
nand U13519 (N_13519,N_13271,N_13483);
and U13520 (N_13520,N_13296,N_13353);
and U13521 (N_13521,N_13281,N_13381);
nand U13522 (N_13522,N_13286,N_13391);
nor U13523 (N_13523,N_13359,N_13430);
nand U13524 (N_13524,N_13322,N_13390);
and U13525 (N_13525,N_13386,N_13294);
or U13526 (N_13526,N_13290,N_13341);
nand U13527 (N_13527,N_13434,N_13358);
or U13528 (N_13528,N_13299,N_13260);
nor U13529 (N_13529,N_13301,N_13306);
xor U13530 (N_13530,N_13432,N_13399);
and U13531 (N_13531,N_13409,N_13361);
and U13532 (N_13532,N_13278,N_13493);
xor U13533 (N_13533,N_13499,N_13472);
or U13534 (N_13534,N_13323,N_13304);
or U13535 (N_13535,N_13262,N_13331);
or U13536 (N_13536,N_13495,N_13292);
nand U13537 (N_13537,N_13368,N_13396);
nor U13538 (N_13538,N_13395,N_13410);
nand U13539 (N_13539,N_13316,N_13473);
nand U13540 (N_13540,N_13452,N_13270);
xor U13541 (N_13541,N_13259,N_13388);
and U13542 (N_13542,N_13453,N_13274);
nand U13543 (N_13543,N_13482,N_13329);
xnor U13544 (N_13544,N_13449,N_13376);
nor U13545 (N_13545,N_13369,N_13345);
xnor U13546 (N_13546,N_13479,N_13404);
nand U13547 (N_13547,N_13422,N_13363);
and U13548 (N_13548,N_13283,N_13282);
nor U13549 (N_13549,N_13367,N_13291);
nor U13550 (N_13550,N_13476,N_13494);
and U13551 (N_13551,N_13464,N_13364);
or U13552 (N_13552,N_13383,N_13406);
xor U13553 (N_13553,N_13387,N_13454);
xor U13554 (N_13554,N_13373,N_13275);
nor U13555 (N_13555,N_13357,N_13448);
or U13556 (N_13556,N_13338,N_13269);
nand U13557 (N_13557,N_13374,N_13298);
nor U13558 (N_13558,N_13255,N_13287);
nor U13559 (N_13559,N_13477,N_13419);
nor U13560 (N_13560,N_13354,N_13402);
xor U13561 (N_13561,N_13415,N_13365);
xnor U13562 (N_13562,N_13349,N_13403);
xor U13563 (N_13563,N_13289,N_13447);
nand U13564 (N_13564,N_13324,N_13377);
nand U13565 (N_13565,N_13328,N_13337);
and U13566 (N_13566,N_13256,N_13394);
nand U13567 (N_13567,N_13469,N_13455);
nand U13568 (N_13568,N_13356,N_13343);
or U13569 (N_13569,N_13492,N_13437);
nor U13570 (N_13570,N_13393,N_13276);
or U13571 (N_13571,N_13490,N_13315);
xnor U13572 (N_13572,N_13408,N_13312);
nor U13573 (N_13573,N_13460,N_13253);
and U13574 (N_13574,N_13407,N_13265);
nand U13575 (N_13575,N_13258,N_13261);
or U13576 (N_13576,N_13284,N_13326);
nor U13577 (N_13577,N_13463,N_13264);
xnor U13578 (N_13578,N_13293,N_13486);
nor U13579 (N_13579,N_13351,N_13433);
and U13580 (N_13580,N_13397,N_13314);
and U13581 (N_13581,N_13257,N_13311);
nand U13582 (N_13582,N_13470,N_13429);
nor U13583 (N_13583,N_13342,N_13300);
nand U13584 (N_13584,N_13439,N_13279);
nand U13585 (N_13585,N_13444,N_13421);
and U13586 (N_13586,N_13325,N_13277);
or U13587 (N_13587,N_13320,N_13487);
and U13588 (N_13588,N_13263,N_13272);
xnor U13589 (N_13589,N_13288,N_13438);
nor U13590 (N_13590,N_13266,N_13392);
and U13591 (N_13591,N_13348,N_13441);
xnor U13592 (N_13592,N_13416,N_13375);
and U13593 (N_13593,N_13423,N_13445);
nor U13594 (N_13594,N_13446,N_13426);
or U13595 (N_13595,N_13379,N_13303);
or U13596 (N_13596,N_13352,N_13425);
nor U13597 (N_13597,N_13382,N_13398);
and U13598 (N_13598,N_13428,N_13340);
nor U13599 (N_13599,N_13400,N_13418);
nand U13600 (N_13600,N_13362,N_13370);
nor U13601 (N_13601,N_13466,N_13465);
or U13602 (N_13602,N_13336,N_13346);
xnor U13603 (N_13603,N_13481,N_13468);
xnor U13604 (N_13604,N_13478,N_13308);
and U13605 (N_13605,N_13389,N_13459);
or U13606 (N_13606,N_13305,N_13462);
or U13607 (N_13607,N_13496,N_13330);
and U13608 (N_13608,N_13417,N_13414);
nor U13609 (N_13609,N_13355,N_13333);
nand U13610 (N_13610,N_13366,N_13285);
nor U13611 (N_13611,N_13385,N_13254);
and U13612 (N_13612,N_13475,N_13250);
and U13613 (N_13613,N_13313,N_13252);
and U13614 (N_13614,N_13474,N_13457);
or U13615 (N_13615,N_13431,N_13295);
or U13616 (N_13616,N_13498,N_13442);
nand U13617 (N_13617,N_13297,N_13497);
and U13618 (N_13618,N_13360,N_13384);
nor U13619 (N_13619,N_13302,N_13350);
or U13620 (N_13620,N_13488,N_13458);
xnor U13621 (N_13621,N_13436,N_13372);
xnor U13622 (N_13622,N_13273,N_13327);
and U13623 (N_13623,N_13401,N_13267);
or U13624 (N_13624,N_13380,N_13339);
nor U13625 (N_13625,N_13480,N_13338);
nor U13626 (N_13626,N_13447,N_13287);
and U13627 (N_13627,N_13275,N_13421);
or U13628 (N_13628,N_13356,N_13379);
nor U13629 (N_13629,N_13280,N_13310);
xor U13630 (N_13630,N_13268,N_13375);
and U13631 (N_13631,N_13304,N_13360);
or U13632 (N_13632,N_13346,N_13417);
or U13633 (N_13633,N_13447,N_13471);
nand U13634 (N_13634,N_13374,N_13406);
xnor U13635 (N_13635,N_13295,N_13256);
or U13636 (N_13636,N_13438,N_13272);
or U13637 (N_13637,N_13336,N_13291);
and U13638 (N_13638,N_13387,N_13276);
xnor U13639 (N_13639,N_13266,N_13480);
and U13640 (N_13640,N_13412,N_13365);
or U13641 (N_13641,N_13459,N_13417);
nor U13642 (N_13642,N_13466,N_13264);
nor U13643 (N_13643,N_13414,N_13314);
nor U13644 (N_13644,N_13477,N_13276);
and U13645 (N_13645,N_13487,N_13273);
xnor U13646 (N_13646,N_13307,N_13462);
nand U13647 (N_13647,N_13282,N_13427);
or U13648 (N_13648,N_13424,N_13355);
nor U13649 (N_13649,N_13413,N_13305);
nand U13650 (N_13650,N_13254,N_13467);
and U13651 (N_13651,N_13251,N_13343);
xnor U13652 (N_13652,N_13466,N_13382);
or U13653 (N_13653,N_13476,N_13429);
xor U13654 (N_13654,N_13339,N_13397);
nand U13655 (N_13655,N_13496,N_13380);
xnor U13656 (N_13656,N_13425,N_13298);
nor U13657 (N_13657,N_13293,N_13286);
nand U13658 (N_13658,N_13313,N_13432);
xnor U13659 (N_13659,N_13418,N_13365);
nor U13660 (N_13660,N_13474,N_13335);
xor U13661 (N_13661,N_13396,N_13316);
nand U13662 (N_13662,N_13493,N_13444);
xor U13663 (N_13663,N_13278,N_13453);
nor U13664 (N_13664,N_13277,N_13273);
xor U13665 (N_13665,N_13382,N_13404);
xor U13666 (N_13666,N_13329,N_13253);
or U13667 (N_13667,N_13381,N_13396);
xnor U13668 (N_13668,N_13389,N_13306);
xor U13669 (N_13669,N_13272,N_13261);
nor U13670 (N_13670,N_13433,N_13484);
xnor U13671 (N_13671,N_13434,N_13442);
nor U13672 (N_13672,N_13290,N_13307);
nand U13673 (N_13673,N_13252,N_13421);
and U13674 (N_13674,N_13423,N_13379);
or U13675 (N_13675,N_13373,N_13485);
nor U13676 (N_13676,N_13469,N_13406);
xor U13677 (N_13677,N_13443,N_13342);
xnor U13678 (N_13678,N_13435,N_13327);
xnor U13679 (N_13679,N_13270,N_13334);
or U13680 (N_13680,N_13386,N_13358);
and U13681 (N_13681,N_13347,N_13423);
xor U13682 (N_13682,N_13452,N_13468);
nand U13683 (N_13683,N_13463,N_13375);
nand U13684 (N_13684,N_13379,N_13342);
or U13685 (N_13685,N_13480,N_13460);
and U13686 (N_13686,N_13344,N_13334);
and U13687 (N_13687,N_13350,N_13423);
or U13688 (N_13688,N_13425,N_13466);
or U13689 (N_13689,N_13280,N_13357);
and U13690 (N_13690,N_13363,N_13251);
xnor U13691 (N_13691,N_13269,N_13363);
xor U13692 (N_13692,N_13438,N_13301);
nand U13693 (N_13693,N_13329,N_13465);
nand U13694 (N_13694,N_13396,N_13459);
or U13695 (N_13695,N_13276,N_13362);
and U13696 (N_13696,N_13443,N_13499);
xnor U13697 (N_13697,N_13298,N_13303);
and U13698 (N_13698,N_13301,N_13251);
xor U13699 (N_13699,N_13292,N_13444);
and U13700 (N_13700,N_13259,N_13321);
and U13701 (N_13701,N_13347,N_13260);
nor U13702 (N_13702,N_13482,N_13339);
nor U13703 (N_13703,N_13399,N_13315);
nand U13704 (N_13704,N_13396,N_13455);
xor U13705 (N_13705,N_13319,N_13268);
xnor U13706 (N_13706,N_13443,N_13315);
nor U13707 (N_13707,N_13281,N_13382);
xor U13708 (N_13708,N_13353,N_13470);
xor U13709 (N_13709,N_13491,N_13385);
and U13710 (N_13710,N_13371,N_13456);
nand U13711 (N_13711,N_13381,N_13378);
xor U13712 (N_13712,N_13299,N_13251);
and U13713 (N_13713,N_13480,N_13383);
xnor U13714 (N_13714,N_13400,N_13438);
xor U13715 (N_13715,N_13328,N_13379);
and U13716 (N_13716,N_13281,N_13267);
nand U13717 (N_13717,N_13356,N_13320);
nand U13718 (N_13718,N_13395,N_13281);
and U13719 (N_13719,N_13315,N_13445);
and U13720 (N_13720,N_13296,N_13291);
xnor U13721 (N_13721,N_13448,N_13483);
or U13722 (N_13722,N_13258,N_13457);
nor U13723 (N_13723,N_13288,N_13286);
xnor U13724 (N_13724,N_13303,N_13269);
nor U13725 (N_13725,N_13275,N_13406);
nand U13726 (N_13726,N_13460,N_13452);
xor U13727 (N_13727,N_13347,N_13318);
nor U13728 (N_13728,N_13411,N_13263);
xor U13729 (N_13729,N_13362,N_13410);
nor U13730 (N_13730,N_13467,N_13341);
and U13731 (N_13731,N_13386,N_13404);
or U13732 (N_13732,N_13357,N_13268);
and U13733 (N_13733,N_13490,N_13459);
and U13734 (N_13734,N_13282,N_13346);
xnor U13735 (N_13735,N_13460,N_13487);
nand U13736 (N_13736,N_13428,N_13284);
nor U13737 (N_13737,N_13459,N_13428);
and U13738 (N_13738,N_13293,N_13300);
nand U13739 (N_13739,N_13343,N_13375);
xnor U13740 (N_13740,N_13257,N_13282);
xnor U13741 (N_13741,N_13270,N_13313);
and U13742 (N_13742,N_13497,N_13438);
nor U13743 (N_13743,N_13272,N_13396);
nand U13744 (N_13744,N_13342,N_13475);
or U13745 (N_13745,N_13294,N_13483);
xnor U13746 (N_13746,N_13484,N_13457);
or U13747 (N_13747,N_13304,N_13322);
nand U13748 (N_13748,N_13389,N_13303);
nand U13749 (N_13749,N_13466,N_13260);
nor U13750 (N_13750,N_13583,N_13641);
or U13751 (N_13751,N_13573,N_13539);
nor U13752 (N_13752,N_13534,N_13572);
and U13753 (N_13753,N_13737,N_13611);
or U13754 (N_13754,N_13739,N_13646);
nand U13755 (N_13755,N_13742,N_13569);
nor U13756 (N_13756,N_13512,N_13616);
nor U13757 (N_13757,N_13650,N_13588);
or U13758 (N_13758,N_13501,N_13651);
xor U13759 (N_13759,N_13718,N_13730);
xor U13760 (N_13760,N_13585,N_13744);
or U13761 (N_13761,N_13595,N_13720);
and U13762 (N_13762,N_13557,N_13500);
nor U13763 (N_13763,N_13552,N_13607);
nand U13764 (N_13764,N_13608,N_13656);
and U13765 (N_13765,N_13580,N_13697);
and U13766 (N_13766,N_13526,N_13635);
or U13767 (N_13767,N_13725,N_13628);
or U13768 (N_13768,N_13639,N_13714);
nor U13769 (N_13769,N_13507,N_13693);
nand U13770 (N_13770,N_13536,N_13627);
xor U13771 (N_13771,N_13565,N_13612);
nor U13772 (N_13772,N_13561,N_13509);
xor U13773 (N_13773,N_13516,N_13642);
or U13774 (N_13774,N_13645,N_13578);
or U13775 (N_13775,N_13553,N_13706);
nor U13776 (N_13776,N_13604,N_13615);
xor U13777 (N_13777,N_13638,N_13674);
xnor U13778 (N_13778,N_13729,N_13688);
nor U13779 (N_13779,N_13506,N_13748);
xnor U13780 (N_13780,N_13547,N_13570);
nand U13781 (N_13781,N_13503,N_13733);
or U13782 (N_13782,N_13576,N_13677);
xnor U13783 (N_13783,N_13738,N_13666);
and U13784 (N_13784,N_13695,N_13568);
and U13785 (N_13785,N_13740,N_13746);
and U13786 (N_13786,N_13529,N_13521);
and U13787 (N_13787,N_13523,N_13712);
xor U13788 (N_13788,N_13590,N_13519);
xnor U13789 (N_13789,N_13532,N_13537);
nor U13790 (N_13790,N_13584,N_13551);
nand U13791 (N_13791,N_13518,N_13571);
xnor U13792 (N_13792,N_13665,N_13597);
and U13793 (N_13793,N_13629,N_13685);
or U13794 (N_13794,N_13726,N_13626);
nand U13795 (N_13795,N_13530,N_13727);
and U13796 (N_13796,N_13579,N_13563);
nand U13797 (N_13797,N_13696,N_13717);
nand U13798 (N_13798,N_13687,N_13566);
or U13799 (N_13799,N_13701,N_13623);
and U13800 (N_13800,N_13619,N_13621);
or U13801 (N_13801,N_13541,N_13510);
and U13802 (N_13802,N_13502,N_13589);
nor U13803 (N_13803,N_13649,N_13524);
and U13804 (N_13804,N_13609,N_13513);
or U13805 (N_13805,N_13653,N_13538);
or U13806 (N_13806,N_13731,N_13515);
nor U13807 (N_13807,N_13648,N_13724);
nor U13808 (N_13808,N_13533,N_13577);
nand U13809 (N_13809,N_13603,N_13617);
nand U13810 (N_13810,N_13594,N_13660);
or U13811 (N_13811,N_13599,N_13620);
nor U13812 (N_13812,N_13741,N_13632);
and U13813 (N_13813,N_13508,N_13736);
nor U13814 (N_13814,N_13544,N_13735);
and U13815 (N_13815,N_13670,N_13644);
or U13816 (N_13816,N_13684,N_13698);
and U13817 (N_13817,N_13633,N_13676);
nor U13818 (N_13818,N_13527,N_13596);
nand U13819 (N_13819,N_13517,N_13722);
or U13820 (N_13820,N_13713,N_13686);
or U13821 (N_13821,N_13587,N_13575);
nand U13822 (N_13822,N_13689,N_13679);
nor U13823 (N_13823,N_13559,N_13668);
and U13824 (N_13824,N_13745,N_13564);
and U13825 (N_13825,N_13636,N_13681);
xor U13826 (N_13826,N_13548,N_13593);
nor U13827 (N_13827,N_13683,N_13630);
nand U13828 (N_13828,N_13669,N_13675);
nand U13829 (N_13829,N_13520,N_13601);
nor U13830 (N_13830,N_13702,N_13647);
and U13831 (N_13831,N_13567,N_13691);
nand U13832 (N_13832,N_13732,N_13558);
nor U13833 (N_13833,N_13582,N_13618);
and U13834 (N_13834,N_13540,N_13622);
xnor U13835 (N_13835,N_13721,N_13662);
or U13836 (N_13836,N_13728,N_13624);
nand U13837 (N_13837,N_13708,N_13574);
nor U13838 (N_13838,N_13600,N_13562);
nand U13839 (N_13839,N_13705,N_13711);
and U13840 (N_13840,N_13598,N_13663);
nor U13841 (N_13841,N_13719,N_13699);
nor U13842 (N_13842,N_13555,N_13709);
xor U13843 (N_13843,N_13749,N_13743);
or U13844 (N_13844,N_13522,N_13586);
nand U13845 (N_13845,N_13700,N_13554);
and U13846 (N_13846,N_13704,N_13667);
or U13847 (N_13847,N_13606,N_13707);
xor U13848 (N_13848,N_13591,N_13543);
nand U13849 (N_13849,N_13592,N_13634);
xnor U13850 (N_13850,N_13657,N_13692);
or U13851 (N_13851,N_13614,N_13525);
nand U13852 (N_13852,N_13694,N_13549);
nand U13853 (N_13853,N_13655,N_13542);
nor U13854 (N_13854,N_13690,N_13581);
nor U13855 (N_13855,N_13545,N_13605);
nand U13856 (N_13856,N_13625,N_13528);
xor U13857 (N_13857,N_13710,N_13631);
and U13858 (N_13858,N_13659,N_13556);
or U13859 (N_13859,N_13703,N_13661);
and U13860 (N_13860,N_13560,N_13682);
nand U13861 (N_13861,N_13658,N_13672);
xor U13862 (N_13862,N_13671,N_13680);
or U13863 (N_13863,N_13747,N_13654);
nor U13864 (N_13864,N_13715,N_13535);
nor U13865 (N_13865,N_13652,N_13511);
or U13866 (N_13866,N_13716,N_13514);
nor U13867 (N_13867,N_13643,N_13664);
xnor U13868 (N_13868,N_13723,N_13504);
xnor U13869 (N_13869,N_13505,N_13734);
and U13870 (N_13870,N_13531,N_13640);
nor U13871 (N_13871,N_13602,N_13678);
xnor U13872 (N_13872,N_13613,N_13637);
xor U13873 (N_13873,N_13673,N_13610);
and U13874 (N_13874,N_13550,N_13546);
nand U13875 (N_13875,N_13699,N_13561);
or U13876 (N_13876,N_13729,N_13613);
xnor U13877 (N_13877,N_13694,N_13744);
nand U13878 (N_13878,N_13507,N_13696);
nand U13879 (N_13879,N_13500,N_13647);
nor U13880 (N_13880,N_13596,N_13677);
and U13881 (N_13881,N_13642,N_13515);
nand U13882 (N_13882,N_13521,N_13653);
nand U13883 (N_13883,N_13520,N_13694);
or U13884 (N_13884,N_13534,N_13565);
or U13885 (N_13885,N_13608,N_13516);
nand U13886 (N_13886,N_13597,N_13711);
nand U13887 (N_13887,N_13691,N_13571);
xor U13888 (N_13888,N_13711,N_13575);
xnor U13889 (N_13889,N_13570,N_13502);
or U13890 (N_13890,N_13509,N_13665);
or U13891 (N_13891,N_13541,N_13536);
and U13892 (N_13892,N_13690,N_13567);
xor U13893 (N_13893,N_13512,N_13525);
nand U13894 (N_13894,N_13505,N_13720);
nand U13895 (N_13895,N_13509,N_13730);
nand U13896 (N_13896,N_13698,N_13521);
xor U13897 (N_13897,N_13703,N_13710);
or U13898 (N_13898,N_13591,N_13514);
xnor U13899 (N_13899,N_13593,N_13521);
xnor U13900 (N_13900,N_13651,N_13690);
nor U13901 (N_13901,N_13745,N_13622);
nor U13902 (N_13902,N_13713,N_13628);
nor U13903 (N_13903,N_13536,N_13648);
xor U13904 (N_13904,N_13680,N_13645);
nand U13905 (N_13905,N_13601,N_13539);
or U13906 (N_13906,N_13566,N_13614);
xor U13907 (N_13907,N_13658,N_13735);
nor U13908 (N_13908,N_13542,N_13614);
or U13909 (N_13909,N_13730,N_13729);
xor U13910 (N_13910,N_13592,N_13706);
or U13911 (N_13911,N_13523,N_13670);
nand U13912 (N_13912,N_13683,N_13718);
xor U13913 (N_13913,N_13573,N_13569);
or U13914 (N_13914,N_13552,N_13703);
nor U13915 (N_13915,N_13589,N_13570);
xor U13916 (N_13916,N_13531,N_13656);
xnor U13917 (N_13917,N_13604,N_13601);
and U13918 (N_13918,N_13576,N_13502);
or U13919 (N_13919,N_13585,N_13626);
xnor U13920 (N_13920,N_13505,N_13701);
nand U13921 (N_13921,N_13508,N_13613);
nand U13922 (N_13922,N_13518,N_13634);
xnor U13923 (N_13923,N_13572,N_13545);
xor U13924 (N_13924,N_13727,N_13739);
and U13925 (N_13925,N_13695,N_13533);
and U13926 (N_13926,N_13713,N_13731);
nand U13927 (N_13927,N_13711,N_13680);
xor U13928 (N_13928,N_13623,N_13554);
and U13929 (N_13929,N_13558,N_13637);
and U13930 (N_13930,N_13532,N_13598);
nor U13931 (N_13931,N_13620,N_13504);
nor U13932 (N_13932,N_13549,N_13723);
or U13933 (N_13933,N_13658,N_13637);
nand U13934 (N_13934,N_13656,N_13676);
nor U13935 (N_13935,N_13700,N_13664);
xor U13936 (N_13936,N_13679,N_13636);
xor U13937 (N_13937,N_13604,N_13677);
nand U13938 (N_13938,N_13524,N_13543);
xor U13939 (N_13939,N_13631,N_13584);
or U13940 (N_13940,N_13671,N_13721);
or U13941 (N_13941,N_13608,N_13693);
and U13942 (N_13942,N_13659,N_13629);
or U13943 (N_13943,N_13500,N_13545);
or U13944 (N_13944,N_13628,N_13656);
nand U13945 (N_13945,N_13725,N_13682);
nor U13946 (N_13946,N_13720,N_13538);
or U13947 (N_13947,N_13620,N_13602);
or U13948 (N_13948,N_13585,N_13670);
xnor U13949 (N_13949,N_13717,N_13636);
or U13950 (N_13950,N_13675,N_13739);
or U13951 (N_13951,N_13743,N_13731);
or U13952 (N_13952,N_13632,N_13625);
and U13953 (N_13953,N_13630,N_13663);
nor U13954 (N_13954,N_13582,N_13545);
xnor U13955 (N_13955,N_13553,N_13652);
xor U13956 (N_13956,N_13711,N_13547);
xor U13957 (N_13957,N_13742,N_13630);
nand U13958 (N_13958,N_13732,N_13657);
nand U13959 (N_13959,N_13573,N_13537);
or U13960 (N_13960,N_13622,N_13635);
and U13961 (N_13961,N_13638,N_13623);
nand U13962 (N_13962,N_13744,N_13736);
xnor U13963 (N_13963,N_13687,N_13623);
nand U13964 (N_13964,N_13639,N_13625);
nor U13965 (N_13965,N_13622,N_13556);
nor U13966 (N_13966,N_13718,N_13658);
or U13967 (N_13967,N_13581,N_13696);
or U13968 (N_13968,N_13568,N_13660);
xnor U13969 (N_13969,N_13569,N_13743);
nor U13970 (N_13970,N_13570,N_13694);
or U13971 (N_13971,N_13639,N_13524);
or U13972 (N_13972,N_13618,N_13737);
nand U13973 (N_13973,N_13610,N_13504);
and U13974 (N_13974,N_13617,N_13739);
nand U13975 (N_13975,N_13740,N_13732);
xnor U13976 (N_13976,N_13611,N_13719);
or U13977 (N_13977,N_13646,N_13728);
or U13978 (N_13978,N_13629,N_13523);
xor U13979 (N_13979,N_13529,N_13684);
and U13980 (N_13980,N_13563,N_13674);
and U13981 (N_13981,N_13666,N_13619);
nor U13982 (N_13982,N_13659,N_13583);
nor U13983 (N_13983,N_13509,N_13620);
nand U13984 (N_13984,N_13690,N_13710);
or U13985 (N_13985,N_13577,N_13683);
nor U13986 (N_13986,N_13739,N_13717);
xnor U13987 (N_13987,N_13662,N_13527);
or U13988 (N_13988,N_13608,N_13530);
nand U13989 (N_13989,N_13687,N_13619);
and U13990 (N_13990,N_13742,N_13654);
and U13991 (N_13991,N_13646,N_13506);
or U13992 (N_13992,N_13705,N_13631);
nand U13993 (N_13993,N_13634,N_13698);
or U13994 (N_13994,N_13620,N_13732);
nand U13995 (N_13995,N_13518,N_13543);
and U13996 (N_13996,N_13556,N_13679);
xnor U13997 (N_13997,N_13537,N_13526);
and U13998 (N_13998,N_13550,N_13512);
or U13999 (N_13999,N_13620,N_13704);
and U14000 (N_14000,N_13768,N_13833);
or U14001 (N_14001,N_13982,N_13953);
nor U14002 (N_14002,N_13775,N_13917);
nand U14003 (N_14003,N_13901,N_13893);
or U14004 (N_14004,N_13834,N_13894);
nand U14005 (N_14005,N_13762,N_13809);
and U14006 (N_14006,N_13884,N_13760);
or U14007 (N_14007,N_13880,N_13767);
or U14008 (N_14008,N_13974,N_13858);
and U14009 (N_14009,N_13877,N_13941);
and U14010 (N_14010,N_13853,N_13875);
and U14011 (N_14011,N_13979,N_13784);
nor U14012 (N_14012,N_13907,N_13992);
and U14013 (N_14013,N_13930,N_13954);
xor U14014 (N_14014,N_13786,N_13755);
and U14015 (N_14015,N_13783,N_13935);
or U14016 (N_14016,N_13859,N_13774);
and U14017 (N_14017,N_13978,N_13920);
or U14018 (N_14018,N_13855,N_13895);
nor U14019 (N_14019,N_13942,N_13812);
nand U14020 (N_14020,N_13932,N_13840);
nand U14021 (N_14021,N_13994,N_13802);
nand U14022 (N_14022,N_13811,N_13928);
xnor U14023 (N_14023,N_13826,N_13863);
xnor U14024 (N_14024,N_13850,N_13951);
nor U14025 (N_14025,N_13921,N_13771);
nor U14026 (N_14026,N_13870,N_13997);
or U14027 (N_14027,N_13909,N_13869);
and U14028 (N_14028,N_13780,N_13881);
or U14029 (N_14029,N_13874,N_13857);
nor U14030 (N_14030,N_13960,N_13757);
and U14031 (N_14031,N_13950,N_13801);
xor U14032 (N_14032,N_13989,N_13830);
or U14033 (N_14033,N_13887,N_13910);
xnor U14034 (N_14034,N_13918,N_13911);
xnor U14035 (N_14035,N_13815,N_13965);
nand U14036 (N_14036,N_13899,N_13946);
and U14037 (N_14037,N_13985,N_13929);
nand U14038 (N_14038,N_13842,N_13821);
xnor U14039 (N_14039,N_13864,N_13959);
and U14040 (N_14040,N_13810,N_13849);
or U14041 (N_14041,N_13862,N_13795);
or U14042 (N_14042,N_13754,N_13898);
nor U14043 (N_14043,N_13940,N_13996);
and U14044 (N_14044,N_13963,N_13751);
or U14045 (N_14045,N_13885,N_13927);
and U14046 (N_14046,N_13818,N_13792);
nor U14047 (N_14047,N_13764,N_13759);
nand U14048 (N_14048,N_13816,N_13817);
and U14049 (N_14049,N_13847,N_13793);
and U14050 (N_14050,N_13876,N_13856);
nand U14051 (N_14051,N_13846,N_13756);
nor U14052 (N_14052,N_13938,N_13914);
nor U14053 (N_14053,N_13808,N_13906);
nand U14054 (N_14054,N_13777,N_13984);
nand U14055 (N_14055,N_13890,N_13990);
or U14056 (N_14056,N_13837,N_13902);
nand U14057 (N_14057,N_13948,N_13966);
nor U14058 (N_14058,N_13913,N_13806);
or U14059 (N_14059,N_13993,N_13972);
nand U14060 (N_14060,N_13831,N_13860);
and U14061 (N_14061,N_13970,N_13976);
xor U14062 (N_14062,N_13763,N_13844);
and U14063 (N_14063,N_13790,N_13839);
and U14064 (N_14064,N_13861,N_13796);
xnor U14065 (N_14065,N_13991,N_13886);
and U14066 (N_14066,N_13813,N_13949);
and U14067 (N_14067,N_13805,N_13883);
and U14068 (N_14068,N_13933,N_13867);
nor U14069 (N_14069,N_13804,N_13820);
xor U14070 (N_14070,N_13843,N_13761);
nor U14071 (N_14071,N_13848,N_13787);
nor U14072 (N_14072,N_13865,N_13905);
or U14073 (N_14073,N_13952,N_13915);
nor U14074 (N_14074,N_13766,N_13934);
and U14075 (N_14075,N_13799,N_13878);
xor U14076 (N_14076,N_13981,N_13971);
and U14077 (N_14077,N_13868,N_13828);
xor U14078 (N_14078,N_13879,N_13785);
xor U14079 (N_14079,N_13791,N_13999);
xor U14080 (N_14080,N_13889,N_13838);
nor U14081 (N_14081,N_13904,N_13931);
xor U14082 (N_14082,N_13937,N_13750);
nand U14083 (N_14083,N_13882,N_13753);
nand U14084 (N_14084,N_13822,N_13967);
nand U14085 (N_14085,N_13945,N_13827);
or U14086 (N_14086,N_13936,N_13975);
nand U14087 (N_14087,N_13947,N_13912);
xnor U14088 (N_14088,N_13851,N_13961);
xnor U14089 (N_14089,N_13969,N_13983);
xor U14090 (N_14090,N_13962,N_13925);
and U14091 (N_14091,N_13926,N_13772);
xor U14092 (N_14092,N_13794,N_13903);
nor U14093 (N_14093,N_13797,N_13824);
nand U14094 (N_14094,N_13980,N_13852);
nand U14095 (N_14095,N_13973,N_13968);
and U14096 (N_14096,N_13788,N_13939);
nor U14097 (N_14097,N_13825,N_13958);
xor U14098 (N_14098,N_13916,N_13919);
nand U14099 (N_14099,N_13986,N_13782);
nand U14100 (N_14100,N_13908,N_13922);
nor U14101 (N_14101,N_13923,N_13789);
or U14102 (N_14102,N_13956,N_13776);
or U14103 (N_14103,N_13832,N_13758);
or U14104 (N_14104,N_13900,N_13819);
or U14105 (N_14105,N_13836,N_13924);
nand U14106 (N_14106,N_13871,N_13823);
nand U14107 (N_14107,N_13814,N_13891);
or U14108 (N_14108,N_13964,N_13835);
xor U14109 (N_14109,N_13866,N_13807);
nand U14110 (N_14110,N_13987,N_13841);
xor U14111 (N_14111,N_13897,N_13845);
xnor U14112 (N_14112,N_13892,N_13800);
nand U14113 (N_14113,N_13769,N_13998);
or U14114 (N_14114,N_13803,N_13854);
nand U14115 (N_14115,N_13896,N_13779);
or U14116 (N_14116,N_13752,N_13995);
xor U14117 (N_14117,N_13781,N_13829);
xnor U14118 (N_14118,N_13888,N_13773);
or U14119 (N_14119,N_13977,N_13765);
nor U14120 (N_14120,N_13943,N_13957);
and U14121 (N_14121,N_13770,N_13873);
nor U14122 (N_14122,N_13944,N_13798);
nor U14123 (N_14123,N_13988,N_13778);
or U14124 (N_14124,N_13872,N_13955);
or U14125 (N_14125,N_13872,N_13855);
or U14126 (N_14126,N_13886,N_13881);
or U14127 (N_14127,N_13772,N_13948);
and U14128 (N_14128,N_13982,N_13972);
or U14129 (N_14129,N_13953,N_13930);
nor U14130 (N_14130,N_13844,N_13856);
nor U14131 (N_14131,N_13783,N_13985);
or U14132 (N_14132,N_13862,N_13908);
and U14133 (N_14133,N_13913,N_13792);
or U14134 (N_14134,N_13889,N_13797);
xnor U14135 (N_14135,N_13811,N_13803);
nor U14136 (N_14136,N_13854,N_13997);
nor U14137 (N_14137,N_13950,N_13966);
xnor U14138 (N_14138,N_13819,N_13767);
nand U14139 (N_14139,N_13930,N_13913);
xnor U14140 (N_14140,N_13898,N_13967);
nand U14141 (N_14141,N_13827,N_13850);
and U14142 (N_14142,N_13861,N_13753);
or U14143 (N_14143,N_13946,N_13905);
nor U14144 (N_14144,N_13914,N_13934);
and U14145 (N_14145,N_13783,N_13762);
and U14146 (N_14146,N_13989,N_13759);
nand U14147 (N_14147,N_13869,N_13944);
or U14148 (N_14148,N_13895,N_13830);
or U14149 (N_14149,N_13861,N_13947);
nand U14150 (N_14150,N_13816,N_13935);
nand U14151 (N_14151,N_13925,N_13940);
xnor U14152 (N_14152,N_13768,N_13987);
nand U14153 (N_14153,N_13784,N_13768);
nand U14154 (N_14154,N_13848,N_13942);
nand U14155 (N_14155,N_13965,N_13779);
xnor U14156 (N_14156,N_13759,N_13853);
or U14157 (N_14157,N_13797,N_13945);
or U14158 (N_14158,N_13858,N_13839);
nor U14159 (N_14159,N_13887,N_13755);
nand U14160 (N_14160,N_13916,N_13961);
nand U14161 (N_14161,N_13878,N_13904);
or U14162 (N_14162,N_13914,N_13927);
nor U14163 (N_14163,N_13934,N_13972);
xor U14164 (N_14164,N_13856,N_13961);
or U14165 (N_14165,N_13763,N_13809);
xnor U14166 (N_14166,N_13846,N_13788);
and U14167 (N_14167,N_13889,N_13841);
or U14168 (N_14168,N_13799,N_13838);
and U14169 (N_14169,N_13981,N_13957);
nand U14170 (N_14170,N_13803,N_13886);
and U14171 (N_14171,N_13825,N_13952);
and U14172 (N_14172,N_13793,N_13897);
nand U14173 (N_14173,N_13954,N_13854);
xnor U14174 (N_14174,N_13834,N_13970);
nor U14175 (N_14175,N_13982,N_13853);
xor U14176 (N_14176,N_13855,N_13762);
and U14177 (N_14177,N_13754,N_13779);
nand U14178 (N_14178,N_13965,N_13883);
xor U14179 (N_14179,N_13885,N_13839);
nand U14180 (N_14180,N_13812,N_13892);
nor U14181 (N_14181,N_13988,N_13895);
xor U14182 (N_14182,N_13761,N_13910);
nor U14183 (N_14183,N_13779,N_13807);
or U14184 (N_14184,N_13996,N_13875);
nor U14185 (N_14185,N_13833,N_13844);
xor U14186 (N_14186,N_13969,N_13755);
nand U14187 (N_14187,N_13981,N_13790);
nor U14188 (N_14188,N_13852,N_13954);
nor U14189 (N_14189,N_13978,N_13878);
nor U14190 (N_14190,N_13927,N_13775);
nor U14191 (N_14191,N_13928,N_13797);
nand U14192 (N_14192,N_13809,N_13953);
nand U14193 (N_14193,N_13876,N_13903);
xor U14194 (N_14194,N_13926,N_13932);
and U14195 (N_14195,N_13822,N_13830);
nand U14196 (N_14196,N_13801,N_13841);
nand U14197 (N_14197,N_13959,N_13837);
xnor U14198 (N_14198,N_13796,N_13777);
and U14199 (N_14199,N_13984,N_13931);
or U14200 (N_14200,N_13857,N_13933);
xor U14201 (N_14201,N_13810,N_13885);
nand U14202 (N_14202,N_13878,N_13983);
nor U14203 (N_14203,N_13998,N_13917);
xor U14204 (N_14204,N_13900,N_13843);
and U14205 (N_14205,N_13999,N_13803);
nor U14206 (N_14206,N_13895,N_13999);
nand U14207 (N_14207,N_13840,N_13922);
nand U14208 (N_14208,N_13769,N_13977);
and U14209 (N_14209,N_13980,N_13796);
xnor U14210 (N_14210,N_13838,N_13934);
and U14211 (N_14211,N_13861,N_13888);
or U14212 (N_14212,N_13956,N_13906);
and U14213 (N_14213,N_13894,N_13791);
xnor U14214 (N_14214,N_13776,N_13925);
or U14215 (N_14215,N_13764,N_13967);
nor U14216 (N_14216,N_13849,N_13917);
and U14217 (N_14217,N_13882,N_13930);
xor U14218 (N_14218,N_13896,N_13795);
and U14219 (N_14219,N_13896,N_13916);
xnor U14220 (N_14220,N_13851,N_13878);
xor U14221 (N_14221,N_13833,N_13923);
and U14222 (N_14222,N_13780,N_13908);
or U14223 (N_14223,N_13906,N_13953);
xor U14224 (N_14224,N_13787,N_13914);
nand U14225 (N_14225,N_13941,N_13952);
xor U14226 (N_14226,N_13958,N_13862);
nand U14227 (N_14227,N_13986,N_13907);
or U14228 (N_14228,N_13779,N_13904);
xnor U14229 (N_14229,N_13945,N_13878);
nor U14230 (N_14230,N_13975,N_13847);
nor U14231 (N_14231,N_13919,N_13788);
nand U14232 (N_14232,N_13834,N_13855);
or U14233 (N_14233,N_13963,N_13971);
nand U14234 (N_14234,N_13777,N_13960);
or U14235 (N_14235,N_13979,N_13846);
xnor U14236 (N_14236,N_13975,N_13797);
and U14237 (N_14237,N_13870,N_13754);
and U14238 (N_14238,N_13987,N_13761);
nand U14239 (N_14239,N_13756,N_13949);
xor U14240 (N_14240,N_13931,N_13960);
or U14241 (N_14241,N_13983,N_13902);
nand U14242 (N_14242,N_13939,N_13834);
and U14243 (N_14243,N_13844,N_13806);
xor U14244 (N_14244,N_13785,N_13789);
nand U14245 (N_14245,N_13854,N_13948);
or U14246 (N_14246,N_13925,N_13964);
xnor U14247 (N_14247,N_13883,N_13945);
or U14248 (N_14248,N_13851,N_13951);
nor U14249 (N_14249,N_13970,N_13937);
or U14250 (N_14250,N_14041,N_14230);
nand U14251 (N_14251,N_14133,N_14206);
xor U14252 (N_14252,N_14062,N_14014);
xor U14253 (N_14253,N_14244,N_14129);
nand U14254 (N_14254,N_14099,N_14142);
and U14255 (N_14255,N_14243,N_14124);
nand U14256 (N_14256,N_14074,N_14120);
and U14257 (N_14257,N_14245,N_14144);
nand U14258 (N_14258,N_14107,N_14180);
and U14259 (N_14259,N_14131,N_14228);
or U14260 (N_14260,N_14079,N_14114);
nand U14261 (N_14261,N_14155,N_14015);
xnor U14262 (N_14262,N_14072,N_14147);
and U14263 (N_14263,N_14196,N_14223);
or U14264 (N_14264,N_14018,N_14138);
or U14265 (N_14265,N_14076,N_14025);
nand U14266 (N_14266,N_14174,N_14017);
nor U14267 (N_14267,N_14088,N_14211);
xor U14268 (N_14268,N_14236,N_14219);
nor U14269 (N_14269,N_14190,N_14140);
and U14270 (N_14270,N_14169,N_14179);
nor U14271 (N_14271,N_14020,N_14004);
nand U14272 (N_14272,N_14069,N_14035);
nor U14273 (N_14273,N_14175,N_14104);
xnor U14274 (N_14274,N_14064,N_14019);
or U14275 (N_14275,N_14216,N_14045);
xor U14276 (N_14276,N_14183,N_14071);
nand U14277 (N_14277,N_14077,N_14086);
or U14278 (N_14278,N_14164,N_14221);
nand U14279 (N_14279,N_14002,N_14146);
nand U14280 (N_14280,N_14052,N_14213);
and U14281 (N_14281,N_14225,N_14172);
and U14282 (N_14282,N_14026,N_14205);
nand U14283 (N_14283,N_14091,N_14151);
nand U14284 (N_14284,N_14003,N_14118);
and U14285 (N_14285,N_14009,N_14115);
or U14286 (N_14286,N_14238,N_14182);
and U14287 (N_14287,N_14160,N_14214);
nor U14288 (N_14288,N_14161,N_14116);
xor U14289 (N_14289,N_14051,N_14049);
and U14290 (N_14290,N_14218,N_14101);
or U14291 (N_14291,N_14029,N_14093);
and U14292 (N_14292,N_14143,N_14148);
or U14293 (N_14293,N_14095,N_14134);
nand U14294 (N_14294,N_14028,N_14229);
nor U14295 (N_14295,N_14001,N_14204);
nand U14296 (N_14296,N_14192,N_14149);
and U14297 (N_14297,N_14123,N_14033);
nand U14298 (N_14298,N_14200,N_14157);
and U14299 (N_14299,N_14013,N_14199);
nor U14300 (N_14300,N_14067,N_14171);
nand U14301 (N_14301,N_14130,N_14234);
or U14302 (N_14302,N_14152,N_14168);
xor U14303 (N_14303,N_14112,N_14178);
xnor U14304 (N_14304,N_14187,N_14040);
xor U14305 (N_14305,N_14121,N_14089);
nand U14306 (N_14306,N_14194,N_14034);
or U14307 (N_14307,N_14209,N_14135);
and U14308 (N_14308,N_14188,N_14094);
nand U14309 (N_14309,N_14184,N_14233);
nand U14310 (N_14310,N_14042,N_14239);
or U14311 (N_14311,N_14201,N_14080);
and U14312 (N_14312,N_14141,N_14105);
nand U14313 (N_14313,N_14007,N_14081);
nor U14314 (N_14314,N_14038,N_14203);
nand U14315 (N_14315,N_14136,N_14006);
or U14316 (N_14316,N_14185,N_14113);
nor U14317 (N_14317,N_14247,N_14159);
nor U14318 (N_14318,N_14240,N_14106);
and U14319 (N_14319,N_14048,N_14231);
nand U14320 (N_14320,N_14224,N_14210);
or U14321 (N_14321,N_14046,N_14153);
xor U14322 (N_14322,N_14032,N_14173);
and U14323 (N_14323,N_14012,N_14158);
nor U14324 (N_14324,N_14082,N_14207);
or U14325 (N_14325,N_14057,N_14132);
and U14326 (N_14326,N_14191,N_14128);
nand U14327 (N_14327,N_14167,N_14037);
or U14328 (N_14328,N_14085,N_14165);
nor U14329 (N_14329,N_14126,N_14202);
and U14330 (N_14330,N_14083,N_14117);
nand U14331 (N_14331,N_14145,N_14139);
xnor U14332 (N_14332,N_14217,N_14031);
and U14333 (N_14333,N_14068,N_14189);
and U14334 (N_14334,N_14154,N_14008);
or U14335 (N_14335,N_14056,N_14109);
and U14336 (N_14336,N_14156,N_14023);
nor U14337 (N_14337,N_14050,N_14226);
nand U14338 (N_14338,N_14170,N_14098);
and U14339 (N_14339,N_14021,N_14103);
xnor U14340 (N_14340,N_14039,N_14054);
and U14341 (N_14341,N_14022,N_14059);
nor U14342 (N_14342,N_14186,N_14122);
xnor U14343 (N_14343,N_14066,N_14215);
or U14344 (N_14344,N_14084,N_14119);
xor U14345 (N_14345,N_14073,N_14092);
nand U14346 (N_14346,N_14176,N_14087);
and U14347 (N_14347,N_14235,N_14011);
nor U14348 (N_14348,N_14108,N_14044);
xnor U14349 (N_14349,N_14127,N_14137);
xor U14350 (N_14350,N_14061,N_14030);
xor U14351 (N_14351,N_14197,N_14163);
nor U14352 (N_14352,N_14063,N_14102);
nor U14353 (N_14353,N_14181,N_14198);
nand U14354 (N_14354,N_14249,N_14065);
nor U14355 (N_14355,N_14212,N_14047);
nand U14356 (N_14356,N_14060,N_14016);
and U14357 (N_14357,N_14220,N_14125);
xor U14358 (N_14358,N_14193,N_14090);
nor U14359 (N_14359,N_14000,N_14043);
or U14360 (N_14360,N_14232,N_14100);
nand U14361 (N_14361,N_14195,N_14070);
nand U14362 (N_14362,N_14162,N_14248);
and U14363 (N_14363,N_14111,N_14110);
or U14364 (N_14364,N_14246,N_14241);
and U14365 (N_14365,N_14150,N_14177);
nor U14366 (N_14366,N_14010,N_14096);
nor U14367 (N_14367,N_14005,N_14237);
xor U14368 (N_14368,N_14097,N_14208);
nor U14369 (N_14369,N_14227,N_14036);
nor U14370 (N_14370,N_14078,N_14055);
or U14371 (N_14371,N_14058,N_14024);
nor U14372 (N_14372,N_14075,N_14242);
or U14373 (N_14373,N_14222,N_14027);
nand U14374 (N_14374,N_14053,N_14166);
and U14375 (N_14375,N_14104,N_14222);
nor U14376 (N_14376,N_14106,N_14177);
or U14377 (N_14377,N_14096,N_14113);
nor U14378 (N_14378,N_14178,N_14176);
or U14379 (N_14379,N_14189,N_14128);
and U14380 (N_14380,N_14126,N_14052);
xor U14381 (N_14381,N_14103,N_14117);
nand U14382 (N_14382,N_14136,N_14028);
and U14383 (N_14383,N_14171,N_14080);
and U14384 (N_14384,N_14113,N_14187);
or U14385 (N_14385,N_14198,N_14002);
or U14386 (N_14386,N_14051,N_14081);
nand U14387 (N_14387,N_14075,N_14123);
nor U14388 (N_14388,N_14075,N_14066);
or U14389 (N_14389,N_14096,N_14129);
nand U14390 (N_14390,N_14183,N_14141);
xor U14391 (N_14391,N_14128,N_14123);
nand U14392 (N_14392,N_14083,N_14220);
and U14393 (N_14393,N_14207,N_14072);
nor U14394 (N_14394,N_14245,N_14246);
nor U14395 (N_14395,N_14134,N_14154);
nand U14396 (N_14396,N_14076,N_14116);
xor U14397 (N_14397,N_14120,N_14026);
nand U14398 (N_14398,N_14114,N_14184);
and U14399 (N_14399,N_14040,N_14248);
and U14400 (N_14400,N_14080,N_14205);
nor U14401 (N_14401,N_14095,N_14220);
xnor U14402 (N_14402,N_14180,N_14113);
nand U14403 (N_14403,N_14009,N_14105);
xor U14404 (N_14404,N_14216,N_14131);
nand U14405 (N_14405,N_14113,N_14134);
nand U14406 (N_14406,N_14196,N_14120);
xnor U14407 (N_14407,N_14073,N_14196);
and U14408 (N_14408,N_14208,N_14184);
nand U14409 (N_14409,N_14044,N_14109);
nor U14410 (N_14410,N_14030,N_14074);
or U14411 (N_14411,N_14151,N_14203);
nor U14412 (N_14412,N_14103,N_14240);
xor U14413 (N_14413,N_14081,N_14223);
xnor U14414 (N_14414,N_14056,N_14098);
nand U14415 (N_14415,N_14017,N_14247);
nor U14416 (N_14416,N_14124,N_14168);
xor U14417 (N_14417,N_14039,N_14105);
nand U14418 (N_14418,N_14106,N_14112);
or U14419 (N_14419,N_14245,N_14002);
or U14420 (N_14420,N_14202,N_14125);
or U14421 (N_14421,N_14175,N_14226);
xor U14422 (N_14422,N_14010,N_14235);
xnor U14423 (N_14423,N_14044,N_14118);
nand U14424 (N_14424,N_14227,N_14138);
and U14425 (N_14425,N_14164,N_14033);
or U14426 (N_14426,N_14191,N_14000);
or U14427 (N_14427,N_14193,N_14132);
nand U14428 (N_14428,N_14027,N_14020);
or U14429 (N_14429,N_14108,N_14185);
xnor U14430 (N_14430,N_14036,N_14126);
or U14431 (N_14431,N_14114,N_14049);
or U14432 (N_14432,N_14020,N_14000);
xor U14433 (N_14433,N_14006,N_14025);
or U14434 (N_14434,N_14218,N_14076);
and U14435 (N_14435,N_14081,N_14135);
xor U14436 (N_14436,N_14054,N_14111);
nor U14437 (N_14437,N_14106,N_14158);
xor U14438 (N_14438,N_14153,N_14011);
and U14439 (N_14439,N_14141,N_14179);
and U14440 (N_14440,N_14199,N_14215);
xor U14441 (N_14441,N_14084,N_14071);
nor U14442 (N_14442,N_14018,N_14201);
nor U14443 (N_14443,N_14204,N_14008);
and U14444 (N_14444,N_14231,N_14025);
and U14445 (N_14445,N_14172,N_14114);
and U14446 (N_14446,N_14063,N_14131);
xor U14447 (N_14447,N_14136,N_14123);
or U14448 (N_14448,N_14206,N_14167);
xnor U14449 (N_14449,N_14069,N_14073);
nand U14450 (N_14450,N_14174,N_14232);
nand U14451 (N_14451,N_14021,N_14091);
xnor U14452 (N_14452,N_14011,N_14018);
and U14453 (N_14453,N_14210,N_14172);
xnor U14454 (N_14454,N_14248,N_14242);
nor U14455 (N_14455,N_14206,N_14029);
or U14456 (N_14456,N_14221,N_14003);
and U14457 (N_14457,N_14117,N_14090);
xnor U14458 (N_14458,N_14106,N_14061);
and U14459 (N_14459,N_14016,N_14237);
nand U14460 (N_14460,N_14110,N_14121);
xnor U14461 (N_14461,N_14092,N_14154);
and U14462 (N_14462,N_14164,N_14123);
or U14463 (N_14463,N_14017,N_14137);
or U14464 (N_14464,N_14148,N_14206);
or U14465 (N_14465,N_14240,N_14007);
nor U14466 (N_14466,N_14013,N_14044);
nor U14467 (N_14467,N_14096,N_14114);
nand U14468 (N_14468,N_14143,N_14165);
nand U14469 (N_14469,N_14109,N_14082);
xor U14470 (N_14470,N_14241,N_14185);
nor U14471 (N_14471,N_14149,N_14203);
or U14472 (N_14472,N_14187,N_14016);
nor U14473 (N_14473,N_14007,N_14113);
nor U14474 (N_14474,N_14177,N_14037);
xnor U14475 (N_14475,N_14210,N_14177);
xnor U14476 (N_14476,N_14103,N_14244);
nor U14477 (N_14477,N_14122,N_14165);
nand U14478 (N_14478,N_14103,N_14203);
or U14479 (N_14479,N_14019,N_14059);
and U14480 (N_14480,N_14010,N_14110);
or U14481 (N_14481,N_14169,N_14045);
nor U14482 (N_14482,N_14085,N_14077);
nor U14483 (N_14483,N_14227,N_14158);
nand U14484 (N_14484,N_14249,N_14106);
xor U14485 (N_14485,N_14022,N_14002);
xnor U14486 (N_14486,N_14037,N_14065);
nand U14487 (N_14487,N_14132,N_14232);
nor U14488 (N_14488,N_14230,N_14236);
or U14489 (N_14489,N_14044,N_14000);
nand U14490 (N_14490,N_14157,N_14000);
xor U14491 (N_14491,N_14163,N_14246);
nor U14492 (N_14492,N_14215,N_14032);
or U14493 (N_14493,N_14016,N_14225);
or U14494 (N_14494,N_14245,N_14214);
or U14495 (N_14495,N_14056,N_14023);
or U14496 (N_14496,N_14208,N_14072);
nand U14497 (N_14497,N_14026,N_14216);
nand U14498 (N_14498,N_14018,N_14089);
xnor U14499 (N_14499,N_14158,N_14180);
nor U14500 (N_14500,N_14381,N_14369);
xnor U14501 (N_14501,N_14270,N_14471);
or U14502 (N_14502,N_14461,N_14467);
or U14503 (N_14503,N_14253,N_14393);
or U14504 (N_14504,N_14304,N_14423);
nor U14505 (N_14505,N_14494,N_14449);
and U14506 (N_14506,N_14269,N_14311);
and U14507 (N_14507,N_14300,N_14496);
and U14508 (N_14508,N_14410,N_14367);
nand U14509 (N_14509,N_14479,N_14464);
and U14510 (N_14510,N_14359,N_14360);
xnor U14511 (N_14511,N_14466,N_14402);
and U14512 (N_14512,N_14411,N_14356);
and U14513 (N_14513,N_14344,N_14440);
xor U14514 (N_14514,N_14303,N_14323);
and U14515 (N_14515,N_14302,N_14256);
and U14516 (N_14516,N_14351,N_14493);
or U14517 (N_14517,N_14366,N_14414);
and U14518 (N_14518,N_14305,N_14388);
and U14519 (N_14519,N_14378,N_14383);
and U14520 (N_14520,N_14294,N_14364);
nor U14521 (N_14521,N_14474,N_14347);
or U14522 (N_14522,N_14463,N_14430);
nor U14523 (N_14523,N_14397,N_14322);
nand U14524 (N_14524,N_14319,N_14385);
nor U14525 (N_14525,N_14485,N_14292);
and U14526 (N_14526,N_14308,N_14408);
nor U14527 (N_14527,N_14379,N_14421);
nand U14528 (N_14528,N_14324,N_14276);
nor U14529 (N_14529,N_14382,N_14442);
nor U14530 (N_14530,N_14403,N_14350);
nand U14531 (N_14531,N_14296,N_14336);
nand U14532 (N_14532,N_14268,N_14437);
nor U14533 (N_14533,N_14441,N_14343);
nand U14534 (N_14534,N_14424,N_14499);
xnor U14535 (N_14535,N_14266,N_14353);
nor U14536 (N_14536,N_14370,N_14390);
xnor U14537 (N_14537,N_14352,N_14457);
nand U14538 (N_14538,N_14258,N_14298);
xor U14539 (N_14539,N_14313,N_14368);
or U14540 (N_14540,N_14425,N_14480);
and U14541 (N_14541,N_14257,N_14401);
and U14542 (N_14542,N_14316,N_14317);
nor U14543 (N_14543,N_14484,N_14272);
xnor U14544 (N_14544,N_14309,N_14492);
and U14545 (N_14545,N_14462,N_14330);
and U14546 (N_14546,N_14404,N_14427);
nor U14547 (N_14547,N_14497,N_14454);
xnor U14548 (N_14548,N_14338,N_14418);
xor U14549 (N_14549,N_14416,N_14291);
nand U14550 (N_14550,N_14419,N_14438);
and U14551 (N_14551,N_14259,N_14262);
xnor U14552 (N_14552,N_14355,N_14475);
and U14553 (N_14553,N_14432,N_14469);
or U14554 (N_14554,N_14282,N_14326);
xor U14555 (N_14555,N_14279,N_14306);
nand U14556 (N_14556,N_14387,N_14341);
nand U14557 (N_14557,N_14371,N_14384);
or U14558 (N_14558,N_14377,N_14498);
nor U14559 (N_14559,N_14358,N_14481);
and U14560 (N_14560,N_14389,N_14301);
and U14561 (N_14561,N_14374,N_14446);
nor U14562 (N_14562,N_14261,N_14349);
xor U14563 (N_14563,N_14287,N_14473);
and U14564 (N_14564,N_14456,N_14478);
xnor U14565 (N_14565,N_14486,N_14288);
nand U14566 (N_14566,N_14284,N_14289);
xnor U14567 (N_14567,N_14398,N_14357);
xor U14568 (N_14568,N_14420,N_14459);
nor U14569 (N_14569,N_14400,N_14375);
nor U14570 (N_14570,N_14495,N_14331);
and U14571 (N_14571,N_14407,N_14405);
or U14572 (N_14572,N_14334,N_14487);
xor U14573 (N_14573,N_14490,N_14345);
and U14574 (N_14574,N_14372,N_14264);
xnor U14575 (N_14575,N_14299,N_14314);
nand U14576 (N_14576,N_14340,N_14468);
and U14577 (N_14577,N_14281,N_14290);
and U14578 (N_14578,N_14277,N_14362);
xnor U14579 (N_14579,N_14391,N_14396);
and U14580 (N_14580,N_14491,N_14482);
nand U14581 (N_14581,N_14477,N_14321);
or U14582 (N_14582,N_14489,N_14285);
xnor U14583 (N_14583,N_14318,N_14394);
nand U14584 (N_14584,N_14453,N_14445);
nand U14585 (N_14585,N_14392,N_14483);
or U14586 (N_14586,N_14451,N_14450);
nand U14587 (N_14587,N_14271,N_14337);
nor U14588 (N_14588,N_14470,N_14422);
nand U14589 (N_14589,N_14332,N_14458);
or U14590 (N_14590,N_14431,N_14325);
and U14591 (N_14591,N_14380,N_14339);
and U14592 (N_14592,N_14275,N_14310);
xnor U14593 (N_14593,N_14472,N_14265);
or U14594 (N_14594,N_14376,N_14328);
nor U14595 (N_14595,N_14412,N_14283);
xnor U14596 (N_14596,N_14267,N_14363);
nand U14597 (N_14597,N_14413,N_14333);
and U14598 (N_14598,N_14409,N_14274);
xnor U14599 (N_14599,N_14251,N_14386);
nand U14600 (N_14600,N_14447,N_14307);
nand U14601 (N_14601,N_14315,N_14444);
nand U14602 (N_14602,N_14434,N_14295);
nand U14603 (N_14603,N_14278,N_14286);
or U14604 (N_14604,N_14436,N_14361);
nand U14605 (N_14605,N_14428,N_14439);
or U14606 (N_14606,N_14280,N_14327);
and U14607 (N_14607,N_14254,N_14293);
or U14608 (N_14608,N_14476,N_14250);
and U14609 (N_14609,N_14320,N_14452);
xnor U14610 (N_14610,N_14335,N_14465);
nand U14611 (N_14611,N_14399,N_14435);
xor U14612 (N_14612,N_14429,N_14395);
nand U14613 (N_14613,N_14406,N_14348);
nand U14614 (N_14614,N_14433,N_14346);
or U14615 (N_14615,N_14455,N_14354);
and U14616 (N_14616,N_14260,N_14448);
xnor U14617 (N_14617,N_14426,N_14488);
nand U14618 (N_14618,N_14373,N_14417);
and U14619 (N_14619,N_14255,N_14297);
nor U14620 (N_14620,N_14329,N_14415);
and U14621 (N_14621,N_14365,N_14443);
or U14622 (N_14622,N_14312,N_14263);
nor U14623 (N_14623,N_14273,N_14342);
xor U14624 (N_14624,N_14460,N_14252);
nand U14625 (N_14625,N_14383,N_14489);
xor U14626 (N_14626,N_14468,N_14277);
and U14627 (N_14627,N_14278,N_14456);
nor U14628 (N_14628,N_14258,N_14496);
nand U14629 (N_14629,N_14469,N_14313);
or U14630 (N_14630,N_14304,N_14403);
nor U14631 (N_14631,N_14384,N_14277);
nand U14632 (N_14632,N_14341,N_14311);
nor U14633 (N_14633,N_14271,N_14498);
and U14634 (N_14634,N_14319,N_14431);
nand U14635 (N_14635,N_14263,N_14308);
nor U14636 (N_14636,N_14487,N_14427);
or U14637 (N_14637,N_14287,N_14259);
nor U14638 (N_14638,N_14292,N_14317);
nand U14639 (N_14639,N_14303,N_14283);
or U14640 (N_14640,N_14419,N_14336);
nand U14641 (N_14641,N_14476,N_14305);
xor U14642 (N_14642,N_14322,N_14435);
xnor U14643 (N_14643,N_14269,N_14433);
xor U14644 (N_14644,N_14302,N_14286);
nor U14645 (N_14645,N_14384,N_14420);
nand U14646 (N_14646,N_14312,N_14324);
xor U14647 (N_14647,N_14318,N_14408);
and U14648 (N_14648,N_14263,N_14395);
or U14649 (N_14649,N_14263,N_14490);
xor U14650 (N_14650,N_14317,N_14269);
or U14651 (N_14651,N_14325,N_14284);
or U14652 (N_14652,N_14424,N_14480);
nor U14653 (N_14653,N_14342,N_14301);
or U14654 (N_14654,N_14434,N_14277);
or U14655 (N_14655,N_14316,N_14331);
or U14656 (N_14656,N_14305,N_14306);
and U14657 (N_14657,N_14378,N_14485);
or U14658 (N_14658,N_14492,N_14310);
nor U14659 (N_14659,N_14421,N_14433);
nand U14660 (N_14660,N_14388,N_14359);
nor U14661 (N_14661,N_14425,N_14486);
and U14662 (N_14662,N_14316,N_14351);
or U14663 (N_14663,N_14275,N_14328);
and U14664 (N_14664,N_14416,N_14312);
xor U14665 (N_14665,N_14425,N_14451);
or U14666 (N_14666,N_14471,N_14277);
xor U14667 (N_14667,N_14301,N_14462);
xnor U14668 (N_14668,N_14421,N_14321);
or U14669 (N_14669,N_14302,N_14271);
or U14670 (N_14670,N_14289,N_14374);
xnor U14671 (N_14671,N_14446,N_14493);
xor U14672 (N_14672,N_14252,N_14409);
and U14673 (N_14673,N_14436,N_14391);
or U14674 (N_14674,N_14293,N_14256);
or U14675 (N_14675,N_14286,N_14383);
or U14676 (N_14676,N_14466,N_14496);
nand U14677 (N_14677,N_14449,N_14391);
nand U14678 (N_14678,N_14408,N_14444);
xnor U14679 (N_14679,N_14429,N_14418);
or U14680 (N_14680,N_14438,N_14290);
or U14681 (N_14681,N_14416,N_14357);
xor U14682 (N_14682,N_14495,N_14366);
xnor U14683 (N_14683,N_14268,N_14337);
nand U14684 (N_14684,N_14457,N_14485);
nor U14685 (N_14685,N_14262,N_14343);
nand U14686 (N_14686,N_14345,N_14296);
nor U14687 (N_14687,N_14290,N_14437);
xor U14688 (N_14688,N_14493,N_14367);
nand U14689 (N_14689,N_14358,N_14425);
nand U14690 (N_14690,N_14497,N_14405);
and U14691 (N_14691,N_14495,N_14309);
nand U14692 (N_14692,N_14251,N_14389);
or U14693 (N_14693,N_14462,N_14256);
nor U14694 (N_14694,N_14275,N_14263);
and U14695 (N_14695,N_14252,N_14485);
nand U14696 (N_14696,N_14453,N_14418);
and U14697 (N_14697,N_14345,N_14496);
and U14698 (N_14698,N_14333,N_14315);
or U14699 (N_14699,N_14352,N_14368);
or U14700 (N_14700,N_14357,N_14367);
xnor U14701 (N_14701,N_14302,N_14270);
nor U14702 (N_14702,N_14440,N_14253);
nand U14703 (N_14703,N_14322,N_14289);
nor U14704 (N_14704,N_14385,N_14394);
or U14705 (N_14705,N_14309,N_14424);
and U14706 (N_14706,N_14486,N_14398);
xnor U14707 (N_14707,N_14254,N_14409);
xor U14708 (N_14708,N_14383,N_14411);
nand U14709 (N_14709,N_14428,N_14278);
nand U14710 (N_14710,N_14269,N_14381);
nor U14711 (N_14711,N_14461,N_14318);
nor U14712 (N_14712,N_14463,N_14462);
nor U14713 (N_14713,N_14450,N_14324);
xnor U14714 (N_14714,N_14342,N_14417);
nor U14715 (N_14715,N_14390,N_14384);
nand U14716 (N_14716,N_14479,N_14347);
and U14717 (N_14717,N_14383,N_14287);
or U14718 (N_14718,N_14282,N_14379);
or U14719 (N_14719,N_14327,N_14380);
nor U14720 (N_14720,N_14268,N_14409);
and U14721 (N_14721,N_14296,N_14398);
and U14722 (N_14722,N_14485,N_14498);
xnor U14723 (N_14723,N_14494,N_14479);
and U14724 (N_14724,N_14297,N_14402);
nand U14725 (N_14725,N_14335,N_14328);
nor U14726 (N_14726,N_14374,N_14297);
xnor U14727 (N_14727,N_14275,N_14341);
nand U14728 (N_14728,N_14272,N_14303);
nor U14729 (N_14729,N_14352,N_14260);
nor U14730 (N_14730,N_14329,N_14383);
or U14731 (N_14731,N_14447,N_14471);
xnor U14732 (N_14732,N_14411,N_14325);
nand U14733 (N_14733,N_14260,N_14291);
and U14734 (N_14734,N_14270,N_14337);
nand U14735 (N_14735,N_14407,N_14451);
or U14736 (N_14736,N_14423,N_14387);
or U14737 (N_14737,N_14473,N_14295);
xnor U14738 (N_14738,N_14453,N_14468);
nor U14739 (N_14739,N_14309,N_14480);
xnor U14740 (N_14740,N_14346,N_14380);
and U14741 (N_14741,N_14407,N_14253);
nor U14742 (N_14742,N_14376,N_14320);
or U14743 (N_14743,N_14395,N_14426);
nor U14744 (N_14744,N_14274,N_14347);
or U14745 (N_14745,N_14477,N_14396);
xnor U14746 (N_14746,N_14277,N_14483);
or U14747 (N_14747,N_14394,N_14486);
xor U14748 (N_14748,N_14326,N_14415);
or U14749 (N_14749,N_14367,N_14286);
nand U14750 (N_14750,N_14710,N_14528);
nor U14751 (N_14751,N_14716,N_14513);
or U14752 (N_14752,N_14664,N_14563);
and U14753 (N_14753,N_14660,N_14674);
or U14754 (N_14754,N_14628,N_14744);
nand U14755 (N_14755,N_14668,N_14666);
nor U14756 (N_14756,N_14593,N_14557);
xor U14757 (N_14757,N_14512,N_14518);
nor U14758 (N_14758,N_14706,N_14638);
xor U14759 (N_14759,N_14629,N_14594);
or U14760 (N_14760,N_14527,N_14611);
and U14761 (N_14761,N_14514,N_14502);
and U14762 (N_14762,N_14555,N_14700);
nand U14763 (N_14763,N_14635,N_14573);
nor U14764 (N_14764,N_14616,N_14617);
and U14765 (N_14765,N_14721,N_14575);
and U14766 (N_14766,N_14578,N_14656);
or U14767 (N_14767,N_14570,N_14579);
nor U14768 (N_14768,N_14724,N_14504);
xnor U14769 (N_14769,N_14548,N_14655);
or U14770 (N_14770,N_14590,N_14620);
or U14771 (N_14771,N_14624,N_14582);
nand U14772 (N_14772,N_14542,N_14622);
or U14773 (N_14773,N_14720,N_14610);
nand U14774 (N_14774,N_14735,N_14659);
nor U14775 (N_14775,N_14729,N_14552);
nand U14776 (N_14776,N_14569,N_14585);
nor U14777 (N_14777,N_14601,N_14583);
and U14778 (N_14778,N_14690,N_14670);
and U14779 (N_14779,N_14529,N_14567);
xor U14780 (N_14780,N_14743,N_14540);
xnor U14781 (N_14781,N_14737,N_14707);
or U14782 (N_14782,N_14517,N_14592);
or U14783 (N_14783,N_14562,N_14701);
nand U14784 (N_14784,N_14653,N_14532);
xnor U14785 (N_14785,N_14534,N_14609);
or U14786 (N_14786,N_14725,N_14525);
and U14787 (N_14787,N_14722,N_14597);
and U14788 (N_14788,N_14539,N_14566);
nor U14789 (N_14789,N_14692,N_14697);
nor U14790 (N_14790,N_14549,N_14565);
nand U14791 (N_14791,N_14627,N_14718);
xnor U14792 (N_14792,N_14554,N_14673);
and U14793 (N_14793,N_14694,N_14682);
nand U14794 (N_14794,N_14665,N_14688);
nor U14795 (N_14795,N_14511,N_14516);
and U14796 (N_14796,N_14731,N_14501);
nor U14797 (N_14797,N_14632,N_14551);
nand U14798 (N_14798,N_14723,N_14714);
xnor U14799 (N_14799,N_14506,N_14553);
xor U14800 (N_14800,N_14580,N_14589);
and U14801 (N_14801,N_14507,N_14615);
and U14802 (N_14802,N_14543,N_14538);
nor U14803 (N_14803,N_14509,N_14685);
and U14804 (N_14804,N_14505,N_14571);
and U14805 (N_14805,N_14625,N_14614);
nand U14806 (N_14806,N_14676,N_14564);
xnor U14807 (N_14807,N_14728,N_14645);
nor U14808 (N_14808,N_14630,N_14727);
nor U14809 (N_14809,N_14623,N_14537);
nor U14810 (N_14810,N_14531,N_14715);
nor U14811 (N_14811,N_14671,N_14577);
nand U14812 (N_14812,N_14675,N_14703);
nand U14813 (N_14813,N_14606,N_14595);
or U14814 (N_14814,N_14524,N_14658);
xor U14815 (N_14815,N_14600,N_14641);
xnor U14816 (N_14816,N_14530,N_14604);
xor U14817 (N_14817,N_14695,N_14717);
xor U14818 (N_14818,N_14602,N_14646);
xnor U14819 (N_14819,N_14608,N_14650);
nor U14820 (N_14820,N_14712,N_14719);
or U14821 (N_14821,N_14515,N_14550);
or U14822 (N_14822,N_14683,N_14533);
nand U14823 (N_14823,N_14702,N_14520);
and U14824 (N_14824,N_14568,N_14734);
xor U14825 (N_14825,N_14708,N_14541);
and U14826 (N_14826,N_14576,N_14672);
or U14827 (N_14827,N_14679,N_14684);
nor U14828 (N_14828,N_14560,N_14733);
or U14829 (N_14829,N_14747,N_14581);
and U14830 (N_14830,N_14603,N_14588);
xnor U14831 (N_14831,N_14640,N_14547);
and U14832 (N_14832,N_14745,N_14545);
and U14833 (N_14833,N_14732,N_14619);
nand U14834 (N_14834,N_14654,N_14503);
and U14835 (N_14835,N_14613,N_14738);
xnor U14836 (N_14836,N_14651,N_14662);
and U14837 (N_14837,N_14693,N_14587);
and U14838 (N_14838,N_14599,N_14698);
or U14839 (N_14839,N_14574,N_14681);
xor U14840 (N_14840,N_14596,N_14510);
nand U14841 (N_14841,N_14643,N_14648);
nand U14842 (N_14842,N_14633,N_14536);
and U14843 (N_14843,N_14704,N_14742);
xor U14844 (N_14844,N_14612,N_14689);
xor U14845 (N_14845,N_14686,N_14748);
or U14846 (N_14846,N_14705,N_14591);
nor U14847 (N_14847,N_14652,N_14667);
nand U14848 (N_14848,N_14559,N_14713);
nor U14849 (N_14849,N_14607,N_14746);
or U14850 (N_14850,N_14642,N_14678);
nor U14851 (N_14851,N_14647,N_14558);
or U14852 (N_14852,N_14730,N_14508);
xnor U14853 (N_14853,N_14634,N_14661);
xor U14854 (N_14854,N_14556,N_14739);
and U14855 (N_14855,N_14726,N_14639);
xor U14856 (N_14856,N_14691,N_14605);
nand U14857 (N_14857,N_14523,N_14637);
nand U14858 (N_14858,N_14621,N_14535);
nand U14859 (N_14859,N_14572,N_14709);
nand U14860 (N_14860,N_14521,N_14522);
nor U14861 (N_14861,N_14687,N_14749);
xnor U14862 (N_14862,N_14740,N_14584);
or U14863 (N_14863,N_14677,N_14561);
or U14864 (N_14864,N_14526,N_14696);
nand U14865 (N_14865,N_14631,N_14711);
and U14866 (N_14866,N_14736,N_14626);
xnor U14867 (N_14867,N_14636,N_14699);
nor U14868 (N_14868,N_14544,N_14669);
nand U14869 (N_14869,N_14618,N_14546);
and U14870 (N_14870,N_14680,N_14663);
and U14871 (N_14871,N_14519,N_14741);
nor U14872 (N_14872,N_14598,N_14586);
nand U14873 (N_14873,N_14500,N_14657);
nand U14874 (N_14874,N_14644,N_14649);
and U14875 (N_14875,N_14527,N_14583);
nor U14876 (N_14876,N_14721,N_14542);
nand U14877 (N_14877,N_14748,N_14632);
and U14878 (N_14878,N_14611,N_14693);
nor U14879 (N_14879,N_14607,N_14628);
xnor U14880 (N_14880,N_14687,N_14573);
xor U14881 (N_14881,N_14720,N_14699);
xor U14882 (N_14882,N_14557,N_14658);
xor U14883 (N_14883,N_14612,N_14738);
xnor U14884 (N_14884,N_14678,N_14588);
nor U14885 (N_14885,N_14505,N_14673);
xor U14886 (N_14886,N_14612,N_14515);
and U14887 (N_14887,N_14531,N_14659);
and U14888 (N_14888,N_14670,N_14586);
nor U14889 (N_14889,N_14554,N_14536);
or U14890 (N_14890,N_14584,N_14561);
nand U14891 (N_14891,N_14604,N_14626);
nand U14892 (N_14892,N_14715,N_14582);
nor U14893 (N_14893,N_14618,N_14512);
and U14894 (N_14894,N_14526,N_14523);
xnor U14895 (N_14895,N_14733,N_14713);
nor U14896 (N_14896,N_14523,N_14580);
or U14897 (N_14897,N_14727,N_14723);
xor U14898 (N_14898,N_14545,N_14546);
or U14899 (N_14899,N_14590,N_14605);
and U14900 (N_14900,N_14526,N_14619);
nand U14901 (N_14901,N_14640,N_14604);
nor U14902 (N_14902,N_14637,N_14636);
or U14903 (N_14903,N_14649,N_14583);
and U14904 (N_14904,N_14567,N_14726);
nand U14905 (N_14905,N_14732,N_14557);
or U14906 (N_14906,N_14747,N_14509);
or U14907 (N_14907,N_14710,N_14747);
or U14908 (N_14908,N_14589,N_14545);
xor U14909 (N_14909,N_14590,N_14749);
and U14910 (N_14910,N_14531,N_14606);
or U14911 (N_14911,N_14547,N_14624);
and U14912 (N_14912,N_14568,N_14713);
or U14913 (N_14913,N_14732,N_14646);
and U14914 (N_14914,N_14620,N_14644);
xor U14915 (N_14915,N_14508,N_14581);
xnor U14916 (N_14916,N_14745,N_14719);
or U14917 (N_14917,N_14602,N_14744);
nor U14918 (N_14918,N_14584,N_14729);
nand U14919 (N_14919,N_14590,N_14570);
and U14920 (N_14920,N_14556,N_14646);
nand U14921 (N_14921,N_14733,N_14645);
or U14922 (N_14922,N_14590,N_14696);
xor U14923 (N_14923,N_14543,N_14648);
nor U14924 (N_14924,N_14642,N_14716);
nor U14925 (N_14925,N_14641,N_14642);
nand U14926 (N_14926,N_14644,N_14710);
or U14927 (N_14927,N_14715,N_14683);
and U14928 (N_14928,N_14648,N_14733);
and U14929 (N_14929,N_14592,N_14714);
xor U14930 (N_14930,N_14531,N_14743);
xnor U14931 (N_14931,N_14735,N_14604);
and U14932 (N_14932,N_14685,N_14626);
xor U14933 (N_14933,N_14744,N_14669);
nor U14934 (N_14934,N_14549,N_14570);
nand U14935 (N_14935,N_14579,N_14745);
or U14936 (N_14936,N_14705,N_14639);
and U14937 (N_14937,N_14746,N_14562);
xor U14938 (N_14938,N_14583,N_14538);
or U14939 (N_14939,N_14651,N_14509);
or U14940 (N_14940,N_14666,N_14505);
or U14941 (N_14941,N_14617,N_14612);
or U14942 (N_14942,N_14537,N_14580);
and U14943 (N_14943,N_14631,N_14571);
xnor U14944 (N_14944,N_14530,N_14578);
or U14945 (N_14945,N_14685,N_14579);
nand U14946 (N_14946,N_14667,N_14517);
and U14947 (N_14947,N_14646,N_14649);
nand U14948 (N_14948,N_14671,N_14744);
xor U14949 (N_14949,N_14591,N_14725);
nand U14950 (N_14950,N_14529,N_14725);
xnor U14951 (N_14951,N_14515,N_14718);
xnor U14952 (N_14952,N_14584,N_14722);
nor U14953 (N_14953,N_14718,N_14733);
xnor U14954 (N_14954,N_14700,N_14592);
or U14955 (N_14955,N_14555,N_14667);
xor U14956 (N_14956,N_14735,N_14652);
nor U14957 (N_14957,N_14573,N_14675);
xnor U14958 (N_14958,N_14537,N_14523);
nor U14959 (N_14959,N_14638,N_14565);
nor U14960 (N_14960,N_14643,N_14580);
xor U14961 (N_14961,N_14504,N_14637);
and U14962 (N_14962,N_14517,N_14616);
and U14963 (N_14963,N_14500,N_14681);
xor U14964 (N_14964,N_14623,N_14749);
or U14965 (N_14965,N_14648,N_14663);
nor U14966 (N_14966,N_14619,N_14684);
or U14967 (N_14967,N_14649,N_14677);
and U14968 (N_14968,N_14736,N_14505);
nand U14969 (N_14969,N_14674,N_14620);
nor U14970 (N_14970,N_14651,N_14513);
and U14971 (N_14971,N_14601,N_14741);
nor U14972 (N_14972,N_14530,N_14513);
or U14973 (N_14973,N_14514,N_14564);
nor U14974 (N_14974,N_14538,N_14746);
xnor U14975 (N_14975,N_14569,N_14679);
and U14976 (N_14976,N_14598,N_14695);
xor U14977 (N_14977,N_14600,N_14643);
xnor U14978 (N_14978,N_14622,N_14627);
and U14979 (N_14979,N_14710,N_14584);
and U14980 (N_14980,N_14658,N_14584);
xnor U14981 (N_14981,N_14740,N_14741);
nand U14982 (N_14982,N_14693,N_14645);
and U14983 (N_14983,N_14594,N_14678);
and U14984 (N_14984,N_14554,N_14565);
and U14985 (N_14985,N_14613,N_14659);
or U14986 (N_14986,N_14730,N_14625);
and U14987 (N_14987,N_14730,N_14616);
xnor U14988 (N_14988,N_14689,N_14562);
nand U14989 (N_14989,N_14601,N_14542);
nor U14990 (N_14990,N_14667,N_14664);
xnor U14991 (N_14991,N_14720,N_14594);
and U14992 (N_14992,N_14514,N_14654);
or U14993 (N_14993,N_14618,N_14654);
nand U14994 (N_14994,N_14554,N_14561);
nor U14995 (N_14995,N_14515,N_14591);
nor U14996 (N_14996,N_14621,N_14514);
xor U14997 (N_14997,N_14616,N_14550);
nand U14998 (N_14998,N_14622,N_14533);
xnor U14999 (N_14999,N_14660,N_14559);
xor U15000 (N_15000,N_14760,N_14901);
and U15001 (N_15001,N_14931,N_14854);
and U15002 (N_15002,N_14956,N_14763);
xnor U15003 (N_15003,N_14769,N_14878);
or U15004 (N_15004,N_14967,N_14975);
nand U15005 (N_15005,N_14885,N_14940);
xnor U15006 (N_15006,N_14987,N_14910);
nand U15007 (N_15007,N_14918,N_14973);
xnor U15008 (N_15008,N_14806,N_14906);
xnor U15009 (N_15009,N_14894,N_14865);
xnor U15010 (N_15010,N_14882,N_14823);
nor U15011 (N_15011,N_14807,N_14771);
nor U15012 (N_15012,N_14884,N_14965);
nor U15013 (N_15013,N_14850,N_14880);
and U15014 (N_15014,N_14876,N_14893);
xor U15015 (N_15015,N_14838,N_14890);
and U15016 (N_15016,N_14934,N_14974);
nand U15017 (N_15017,N_14881,N_14813);
nand U15018 (N_15018,N_14916,N_14820);
xor U15019 (N_15019,N_14919,N_14752);
nor U15020 (N_15020,N_14909,N_14992);
and U15021 (N_15021,N_14946,N_14796);
nor U15022 (N_15022,N_14842,N_14976);
nand U15023 (N_15023,N_14811,N_14913);
nand U15024 (N_15024,N_14791,N_14867);
nand U15025 (N_15025,N_14793,N_14832);
and U15026 (N_15026,N_14907,N_14912);
and U15027 (N_15027,N_14911,N_14799);
or U15028 (N_15028,N_14817,N_14843);
and U15029 (N_15029,N_14874,N_14908);
nand U15030 (N_15030,N_14966,N_14941);
or U15031 (N_15031,N_14824,N_14954);
xor U15032 (N_15032,N_14785,N_14944);
nand U15033 (N_15033,N_14795,N_14750);
nand U15034 (N_15034,N_14939,N_14859);
and U15035 (N_15035,N_14869,N_14979);
and U15036 (N_15036,N_14801,N_14904);
or U15037 (N_15037,N_14831,N_14942);
xnor U15038 (N_15038,N_14856,N_14819);
and U15039 (N_15039,N_14927,N_14822);
xnor U15040 (N_15040,N_14764,N_14937);
nor U15041 (N_15041,N_14778,N_14960);
xnor U15042 (N_15042,N_14922,N_14943);
nand U15043 (N_15043,N_14810,N_14768);
and U15044 (N_15044,N_14905,N_14947);
xnor U15045 (N_15045,N_14929,N_14797);
nor U15046 (N_15046,N_14818,N_14871);
and U15047 (N_15047,N_14920,N_14751);
xor U15048 (N_15048,N_14825,N_14873);
and U15049 (N_15049,N_14926,N_14846);
or U15050 (N_15050,N_14945,N_14892);
and U15051 (N_15051,N_14756,N_14952);
xnor U15052 (N_15052,N_14808,N_14870);
xnor U15053 (N_15053,N_14955,N_14949);
or U15054 (N_15054,N_14816,N_14898);
nor U15055 (N_15055,N_14993,N_14963);
nor U15056 (N_15056,N_14917,N_14784);
nor U15057 (N_15057,N_14962,N_14977);
or U15058 (N_15058,N_14923,N_14789);
xnor U15059 (N_15059,N_14875,N_14803);
nand U15060 (N_15060,N_14950,N_14997);
xor U15061 (N_15061,N_14903,N_14780);
and U15062 (N_15062,N_14996,N_14834);
or U15063 (N_15063,N_14981,N_14897);
xor U15064 (N_15064,N_14775,N_14837);
and U15065 (N_15065,N_14896,N_14852);
nor U15066 (N_15066,N_14957,N_14985);
and U15067 (N_15067,N_14938,N_14936);
nor U15068 (N_15068,N_14921,N_14872);
xnor U15069 (N_15069,N_14829,N_14932);
or U15070 (N_15070,N_14858,N_14899);
and U15071 (N_15071,N_14928,N_14833);
nor U15072 (N_15072,N_14969,N_14847);
nand U15073 (N_15073,N_14781,N_14844);
nor U15074 (N_15074,N_14788,N_14933);
xnor U15075 (N_15075,N_14805,N_14891);
xnor U15076 (N_15076,N_14959,N_14984);
or U15077 (N_15077,N_14887,N_14958);
and U15078 (N_15078,N_14986,N_14830);
and U15079 (N_15079,N_14924,N_14840);
xor U15080 (N_15080,N_14779,N_14988);
nor U15081 (N_15081,N_14828,N_14755);
xor U15082 (N_15082,N_14776,N_14783);
nor U15083 (N_15083,N_14990,N_14868);
nor U15084 (N_15084,N_14895,N_14766);
xnor U15085 (N_15085,N_14777,N_14836);
nand U15086 (N_15086,N_14948,N_14902);
and U15087 (N_15087,N_14982,N_14839);
xor U15088 (N_15088,N_14800,N_14765);
nand U15089 (N_15089,N_14925,N_14970);
xor U15090 (N_15090,N_14862,N_14972);
or U15091 (N_15091,N_14877,N_14857);
xor U15092 (N_15092,N_14802,N_14971);
or U15093 (N_15093,N_14798,N_14761);
and U15094 (N_15094,N_14883,N_14792);
or U15095 (N_15095,N_14851,N_14991);
nand U15096 (N_15096,N_14758,N_14794);
nand U15097 (N_15097,N_14804,N_14964);
nor U15098 (N_15098,N_14812,N_14860);
and U15099 (N_15099,N_14853,N_14827);
or U15100 (N_15100,N_14900,N_14889);
nor U15101 (N_15101,N_14790,N_14773);
or U15102 (N_15102,N_14753,N_14961);
nand U15103 (N_15103,N_14995,N_14914);
xor U15104 (N_15104,N_14762,N_14849);
xor U15105 (N_15105,N_14787,N_14809);
nand U15106 (N_15106,N_14866,N_14951);
nand U15107 (N_15107,N_14855,N_14772);
nor U15108 (N_15108,N_14861,N_14848);
or U15109 (N_15109,N_14770,N_14953);
nor U15110 (N_15110,N_14845,N_14886);
xnor U15111 (N_15111,N_14915,N_14767);
xnor U15112 (N_15112,N_14774,N_14814);
nor U15113 (N_15113,N_14978,N_14826);
or U15114 (N_15114,N_14994,N_14782);
nand U15115 (N_15115,N_14863,N_14757);
or U15116 (N_15116,N_14888,N_14759);
nand U15117 (N_15117,N_14989,N_14864);
xnor U15118 (N_15118,N_14980,N_14815);
xor U15119 (N_15119,N_14754,N_14821);
nor U15120 (N_15120,N_14999,N_14935);
nand U15121 (N_15121,N_14983,N_14841);
nor U15122 (N_15122,N_14998,N_14968);
nor U15123 (N_15123,N_14835,N_14786);
nor U15124 (N_15124,N_14930,N_14879);
or U15125 (N_15125,N_14827,N_14951);
nand U15126 (N_15126,N_14834,N_14944);
or U15127 (N_15127,N_14929,N_14777);
xor U15128 (N_15128,N_14977,N_14778);
or U15129 (N_15129,N_14806,N_14994);
or U15130 (N_15130,N_14896,N_14765);
nor U15131 (N_15131,N_14823,N_14860);
or U15132 (N_15132,N_14769,N_14799);
and U15133 (N_15133,N_14891,N_14840);
and U15134 (N_15134,N_14801,N_14821);
xnor U15135 (N_15135,N_14959,N_14958);
nor U15136 (N_15136,N_14951,N_14974);
nand U15137 (N_15137,N_14981,N_14754);
and U15138 (N_15138,N_14839,N_14856);
or U15139 (N_15139,N_14822,N_14806);
or U15140 (N_15140,N_14967,N_14969);
and U15141 (N_15141,N_14759,N_14763);
xnor U15142 (N_15142,N_14835,N_14769);
xor U15143 (N_15143,N_14754,N_14790);
xnor U15144 (N_15144,N_14827,N_14861);
xnor U15145 (N_15145,N_14766,N_14795);
and U15146 (N_15146,N_14973,N_14827);
xor U15147 (N_15147,N_14958,N_14754);
nor U15148 (N_15148,N_14938,N_14935);
or U15149 (N_15149,N_14845,N_14762);
nand U15150 (N_15150,N_14928,N_14914);
nand U15151 (N_15151,N_14990,N_14785);
nor U15152 (N_15152,N_14923,N_14803);
xnor U15153 (N_15153,N_14923,N_14949);
nor U15154 (N_15154,N_14967,N_14786);
and U15155 (N_15155,N_14756,N_14785);
nor U15156 (N_15156,N_14853,N_14902);
nor U15157 (N_15157,N_14857,N_14786);
xor U15158 (N_15158,N_14864,N_14827);
xor U15159 (N_15159,N_14974,N_14789);
and U15160 (N_15160,N_14993,N_14976);
and U15161 (N_15161,N_14757,N_14819);
xor U15162 (N_15162,N_14924,N_14976);
and U15163 (N_15163,N_14976,N_14757);
nand U15164 (N_15164,N_14897,N_14948);
nor U15165 (N_15165,N_14921,N_14940);
or U15166 (N_15166,N_14902,N_14781);
nor U15167 (N_15167,N_14942,N_14977);
nor U15168 (N_15168,N_14922,N_14803);
or U15169 (N_15169,N_14889,N_14817);
nor U15170 (N_15170,N_14997,N_14920);
nor U15171 (N_15171,N_14940,N_14974);
or U15172 (N_15172,N_14856,N_14776);
or U15173 (N_15173,N_14924,N_14899);
or U15174 (N_15174,N_14866,N_14848);
and U15175 (N_15175,N_14759,N_14940);
xor U15176 (N_15176,N_14930,N_14835);
xnor U15177 (N_15177,N_14844,N_14917);
xor U15178 (N_15178,N_14805,N_14884);
nand U15179 (N_15179,N_14870,N_14811);
and U15180 (N_15180,N_14850,N_14973);
xor U15181 (N_15181,N_14957,N_14898);
or U15182 (N_15182,N_14760,N_14911);
or U15183 (N_15183,N_14863,N_14967);
and U15184 (N_15184,N_14905,N_14934);
and U15185 (N_15185,N_14813,N_14822);
nor U15186 (N_15186,N_14919,N_14848);
xor U15187 (N_15187,N_14761,N_14946);
nand U15188 (N_15188,N_14806,N_14876);
xnor U15189 (N_15189,N_14841,N_14802);
and U15190 (N_15190,N_14784,N_14790);
and U15191 (N_15191,N_14898,N_14941);
or U15192 (N_15192,N_14876,N_14820);
nor U15193 (N_15193,N_14840,N_14910);
nand U15194 (N_15194,N_14783,N_14871);
nor U15195 (N_15195,N_14775,N_14760);
or U15196 (N_15196,N_14995,N_14796);
and U15197 (N_15197,N_14917,N_14995);
and U15198 (N_15198,N_14897,N_14851);
nor U15199 (N_15199,N_14916,N_14878);
nand U15200 (N_15200,N_14827,N_14939);
and U15201 (N_15201,N_14872,N_14780);
nand U15202 (N_15202,N_14893,N_14822);
nor U15203 (N_15203,N_14752,N_14948);
and U15204 (N_15204,N_14926,N_14826);
nand U15205 (N_15205,N_14785,N_14847);
nand U15206 (N_15206,N_14834,N_14973);
xor U15207 (N_15207,N_14979,N_14999);
or U15208 (N_15208,N_14783,N_14788);
or U15209 (N_15209,N_14877,N_14939);
or U15210 (N_15210,N_14793,N_14972);
or U15211 (N_15211,N_14776,N_14839);
nor U15212 (N_15212,N_14915,N_14841);
nand U15213 (N_15213,N_14949,N_14836);
xnor U15214 (N_15214,N_14897,N_14983);
xor U15215 (N_15215,N_14815,N_14989);
nand U15216 (N_15216,N_14814,N_14905);
or U15217 (N_15217,N_14886,N_14998);
nor U15218 (N_15218,N_14869,N_14943);
and U15219 (N_15219,N_14847,N_14817);
xnor U15220 (N_15220,N_14972,N_14863);
xor U15221 (N_15221,N_14823,N_14754);
or U15222 (N_15222,N_14841,N_14966);
and U15223 (N_15223,N_14777,N_14783);
and U15224 (N_15224,N_14894,N_14851);
and U15225 (N_15225,N_14770,N_14773);
xnor U15226 (N_15226,N_14843,N_14750);
nand U15227 (N_15227,N_14797,N_14916);
or U15228 (N_15228,N_14874,N_14850);
nor U15229 (N_15229,N_14921,N_14862);
or U15230 (N_15230,N_14931,N_14997);
nor U15231 (N_15231,N_14775,N_14901);
or U15232 (N_15232,N_14893,N_14953);
xnor U15233 (N_15233,N_14831,N_14885);
nand U15234 (N_15234,N_14931,N_14873);
nor U15235 (N_15235,N_14952,N_14915);
xnor U15236 (N_15236,N_14787,N_14892);
or U15237 (N_15237,N_14988,N_14819);
and U15238 (N_15238,N_14823,N_14784);
xnor U15239 (N_15239,N_14949,N_14966);
nor U15240 (N_15240,N_14837,N_14770);
nand U15241 (N_15241,N_14777,N_14816);
nand U15242 (N_15242,N_14842,N_14965);
nor U15243 (N_15243,N_14905,N_14938);
nand U15244 (N_15244,N_14871,N_14846);
nor U15245 (N_15245,N_14805,N_14776);
nor U15246 (N_15246,N_14964,N_14830);
xor U15247 (N_15247,N_14759,N_14781);
nand U15248 (N_15248,N_14877,N_14875);
or U15249 (N_15249,N_14826,N_14769);
nor U15250 (N_15250,N_15244,N_15049);
xnor U15251 (N_15251,N_15129,N_15139);
xnor U15252 (N_15252,N_15005,N_15219);
or U15253 (N_15253,N_15233,N_15059);
nor U15254 (N_15254,N_15030,N_15141);
and U15255 (N_15255,N_15038,N_15043);
or U15256 (N_15256,N_15164,N_15154);
and U15257 (N_15257,N_15151,N_15065);
nor U15258 (N_15258,N_15101,N_15202);
or U15259 (N_15259,N_15127,N_15185);
nand U15260 (N_15260,N_15207,N_15175);
and U15261 (N_15261,N_15234,N_15144);
or U15262 (N_15262,N_15146,N_15147);
or U15263 (N_15263,N_15203,N_15196);
nand U15264 (N_15264,N_15120,N_15015);
and U15265 (N_15265,N_15078,N_15072);
or U15266 (N_15266,N_15084,N_15089);
nor U15267 (N_15267,N_15247,N_15054);
or U15268 (N_15268,N_15158,N_15083);
and U15269 (N_15269,N_15241,N_15169);
or U15270 (N_15270,N_15042,N_15097);
nand U15271 (N_15271,N_15200,N_15080);
and U15272 (N_15272,N_15240,N_15011);
xor U15273 (N_15273,N_15004,N_15071);
and U15274 (N_15274,N_15021,N_15137);
or U15275 (N_15275,N_15201,N_15070);
or U15276 (N_15276,N_15124,N_15179);
nor U15277 (N_15277,N_15022,N_15152);
and U15278 (N_15278,N_15093,N_15055);
or U15279 (N_15279,N_15012,N_15035);
nand U15280 (N_15280,N_15160,N_15140);
xor U15281 (N_15281,N_15106,N_15232);
or U15282 (N_15282,N_15061,N_15226);
nand U15283 (N_15283,N_15193,N_15047);
nor U15284 (N_15284,N_15216,N_15066);
and U15285 (N_15285,N_15033,N_15103);
nor U15286 (N_15286,N_15192,N_15198);
nand U15287 (N_15287,N_15181,N_15115);
nor U15288 (N_15288,N_15121,N_15003);
nor U15289 (N_15289,N_15117,N_15087);
xnor U15290 (N_15290,N_15224,N_15010);
xor U15291 (N_15291,N_15161,N_15046);
or U15292 (N_15292,N_15039,N_15211);
or U15293 (N_15293,N_15027,N_15095);
xnor U15294 (N_15294,N_15096,N_15057);
xnor U15295 (N_15295,N_15218,N_15090);
nand U15296 (N_15296,N_15183,N_15170);
and U15297 (N_15297,N_15001,N_15116);
or U15298 (N_15298,N_15212,N_15053);
and U15299 (N_15299,N_15168,N_15014);
nor U15300 (N_15300,N_15236,N_15023);
nand U15301 (N_15301,N_15220,N_15032);
nand U15302 (N_15302,N_15111,N_15214);
and U15303 (N_15303,N_15123,N_15159);
xor U15304 (N_15304,N_15017,N_15197);
and U15305 (N_15305,N_15077,N_15237);
or U15306 (N_15306,N_15209,N_15187);
xnor U15307 (N_15307,N_15020,N_15075);
xnor U15308 (N_15308,N_15031,N_15135);
nand U15309 (N_15309,N_15249,N_15045);
nand U15310 (N_15310,N_15007,N_15112);
and U15311 (N_15311,N_15190,N_15081);
nor U15312 (N_15312,N_15025,N_15186);
xor U15313 (N_15313,N_15178,N_15125);
nand U15314 (N_15314,N_15088,N_15091);
or U15315 (N_15315,N_15002,N_15036);
nand U15316 (N_15316,N_15191,N_15060);
nor U15317 (N_15317,N_15056,N_15098);
and U15318 (N_15318,N_15184,N_15136);
or U15319 (N_15319,N_15157,N_15188);
and U15320 (N_15320,N_15165,N_15248);
xor U15321 (N_15321,N_15052,N_15148);
nor U15322 (N_15322,N_15118,N_15199);
and U15323 (N_15323,N_15213,N_15149);
and U15324 (N_15324,N_15040,N_15107);
or U15325 (N_15325,N_15013,N_15051);
or U15326 (N_15326,N_15133,N_15016);
and U15327 (N_15327,N_15063,N_15104);
xor U15328 (N_15328,N_15138,N_15028);
and U15329 (N_15329,N_15108,N_15131);
nand U15330 (N_15330,N_15153,N_15182);
nor U15331 (N_15331,N_15128,N_15222);
or U15332 (N_15332,N_15174,N_15204);
and U15333 (N_15333,N_15074,N_15019);
nor U15334 (N_15334,N_15073,N_15082);
nand U15335 (N_15335,N_15134,N_15150);
nor U15336 (N_15336,N_15243,N_15227);
or U15337 (N_15337,N_15099,N_15092);
nand U15338 (N_15338,N_15119,N_15189);
and U15339 (N_15339,N_15048,N_15210);
nor U15340 (N_15340,N_15126,N_15246);
xor U15341 (N_15341,N_15041,N_15067);
xnor U15342 (N_15342,N_15105,N_15029);
nor U15343 (N_15343,N_15206,N_15102);
or U15344 (N_15344,N_15215,N_15113);
nand U15345 (N_15345,N_15026,N_15062);
or U15346 (N_15346,N_15037,N_15205);
and U15347 (N_15347,N_15069,N_15024);
xnor U15348 (N_15348,N_15034,N_15180);
or U15349 (N_15349,N_15217,N_15235);
nand U15350 (N_15350,N_15195,N_15177);
xnor U15351 (N_15351,N_15044,N_15006);
nor U15352 (N_15352,N_15167,N_15109);
xor U15353 (N_15353,N_15114,N_15221);
xnor U15354 (N_15354,N_15122,N_15000);
xor U15355 (N_15355,N_15172,N_15018);
nor U15356 (N_15356,N_15130,N_15173);
nor U15357 (N_15357,N_15064,N_15155);
nor U15358 (N_15358,N_15132,N_15231);
nand U15359 (N_15359,N_15076,N_15171);
nand U15360 (N_15360,N_15245,N_15156);
and U15361 (N_15361,N_15162,N_15223);
xnor U15362 (N_15362,N_15230,N_15225);
xnor U15363 (N_15363,N_15050,N_15242);
nand U15364 (N_15364,N_15100,N_15194);
nor U15365 (N_15365,N_15085,N_15009);
xor U15366 (N_15366,N_15143,N_15086);
and U15367 (N_15367,N_15166,N_15058);
nand U15368 (N_15368,N_15208,N_15142);
xnor U15369 (N_15369,N_15229,N_15110);
nor U15370 (N_15370,N_15176,N_15094);
xor U15371 (N_15371,N_15228,N_15008);
xor U15372 (N_15372,N_15079,N_15238);
and U15373 (N_15373,N_15068,N_15239);
nor U15374 (N_15374,N_15145,N_15163);
nand U15375 (N_15375,N_15092,N_15088);
or U15376 (N_15376,N_15053,N_15098);
xor U15377 (N_15377,N_15245,N_15187);
and U15378 (N_15378,N_15026,N_15108);
nor U15379 (N_15379,N_15013,N_15112);
or U15380 (N_15380,N_15125,N_15200);
xor U15381 (N_15381,N_15146,N_15116);
or U15382 (N_15382,N_15149,N_15107);
xnor U15383 (N_15383,N_15042,N_15135);
xnor U15384 (N_15384,N_15146,N_15210);
xnor U15385 (N_15385,N_15017,N_15057);
nand U15386 (N_15386,N_15025,N_15041);
and U15387 (N_15387,N_15227,N_15110);
nand U15388 (N_15388,N_15094,N_15247);
or U15389 (N_15389,N_15171,N_15113);
or U15390 (N_15390,N_15079,N_15231);
and U15391 (N_15391,N_15240,N_15024);
nand U15392 (N_15392,N_15247,N_15062);
or U15393 (N_15393,N_15003,N_15241);
and U15394 (N_15394,N_15144,N_15076);
nor U15395 (N_15395,N_15001,N_15232);
or U15396 (N_15396,N_15203,N_15003);
and U15397 (N_15397,N_15170,N_15186);
nand U15398 (N_15398,N_15065,N_15191);
or U15399 (N_15399,N_15010,N_15033);
nand U15400 (N_15400,N_15229,N_15129);
or U15401 (N_15401,N_15220,N_15123);
or U15402 (N_15402,N_15164,N_15005);
nor U15403 (N_15403,N_15021,N_15052);
or U15404 (N_15404,N_15020,N_15171);
or U15405 (N_15405,N_15126,N_15098);
nand U15406 (N_15406,N_15091,N_15245);
or U15407 (N_15407,N_15191,N_15170);
nand U15408 (N_15408,N_15138,N_15223);
nand U15409 (N_15409,N_15073,N_15121);
xnor U15410 (N_15410,N_15090,N_15003);
and U15411 (N_15411,N_15138,N_15063);
nor U15412 (N_15412,N_15045,N_15172);
and U15413 (N_15413,N_15168,N_15004);
xnor U15414 (N_15414,N_15214,N_15100);
xor U15415 (N_15415,N_15050,N_15041);
xnor U15416 (N_15416,N_15222,N_15003);
nand U15417 (N_15417,N_15217,N_15189);
xor U15418 (N_15418,N_15086,N_15000);
xnor U15419 (N_15419,N_15156,N_15191);
xor U15420 (N_15420,N_15219,N_15126);
or U15421 (N_15421,N_15220,N_15158);
and U15422 (N_15422,N_15086,N_15116);
and U15423 (N_15423,N_15079,N_15240);
xnor U15424 (N_15424,N_15144,N_15190);
xor U15425 (N_15425,N_15241,N_15058);
nand U15426 (N_15426,N_15222,N_15100);
xor U15427 (N_15427,N_15097,N_15218);
nand U15428 (N_15428,N_15214,N_15078);
xor U15429 (N_15429,N_15007,N_15003);
nand U15430 (N_15430,N_15049,N_15069);
xor U15431 (N_15431,N_15167,N_15129);
xor U15432 (N_15432,N_15137,N_15022);
and U15433 (N_15433,N_15234,N_15213);
xnor U15434 (N_15434,N_15066,N_15146);
or U15435 (N_15435,N_15200,N_15100);
xor U15436 (N_15436,N_15123,N_15116);
nor U15437 (N_15437,N_15055,N_15004);
and U15438 (N_15438,N_15243,N_15212);
xnor U15439 (N_15439,N_15109,N_15169);
xor U15440 (N_15440,N_15007,N_15149);
xnor U15441 (N_15441,N_15086,N_15208);
or U15442 (N_15442,N_15149,N_15086);
nor U15443 (N_15443,N_15198,N_15062);
nand U15444 (N_15444,N_15084,N_15110);
or U15445 (N_15445,N_15198,N_15163);
and U15446 (N_15446,N_15120,N_15229);
xnor U15447 (N_15447,N_15132,N_15094);
nor U15448 (N_15448,N_15013,N_15146);
nor U15449 (N_15449,N_15014,N_15150);
and U15450 (N_15450,N_15210,N_15124);
xnor U15451 (N_15451,N_15159,N_15216);
and U15452 (N_15452,N_15157,N_15059);
nor U15453 (N_15453,N_15071,N_15134);
xor U15454 (N_15454,N_15221,N_15146);
nand U15455 (N_15455,N_15144,N_15151);
xor U15456 (N_15456,N_15035,N_15083);
nand U15457 (N_15457,N_15015,N_15163);
nor U15458 (N_15458,N_15092,N_15143);
or U15459 (N_15459,N_15005,N_15185);
or U15460 (N_15460,N_15073,N_15051);
xor U15461 (N_15461,N_15113,N_15173);
xor U15462 (N_15462,N_15204,N_15090);
xor U15463 (N_15463,N_15181,N_15040);
xnor U15464 (N_15464,N_15210,N_15110);
or U15465 (N_15465,N_15082,N_15100);
xor U15466 (N_15466,N_15186,N_15140);
nand U15467 (N_15467,N_15238,N_15127);
xnor U15468 (N_15468,N_15066,N_15008);
and U15469 (N_15469,N_15014,N_15100);
nor U15470 (N_15470,N_15009,N_15089);
nand U15471 (N_15471,N_15055,N_15048);
or U15472 (N_15472,N_15152,N_15173);
or U15473 (N_15473,N_15197,N_15039);
xnor U15474 (N_15474,N_15229,N_15214);
or U15475 (N_15475,N_15057,N_15108);
nor U15476 (N_15476,N_15204,N_15083);
xnor U15477 (N_15477,N_15008,N_15247);
or U15478 (N_15478,N_15207,N_15016);
xnor U15479 (N_15479,N_15143,N_15096);
and U15480 (N_15480,N_15034,N_15138);
nor U15481 (N_15481,N_15203,N_15128);
xnor U15482 (N_15482,N_15159,N_15188);
nor U15483 (N_15483,N_15133,N_15142);
nand U15484 (N_15484,N_15223,N_15218);
nand U15485 (N_15485,N_15172,N_15070);
or U15486 (N_15486,N_15120,N_15076);
nand U15487 (N_15487,N_15001,N_15078);
xnor U15488 (N_15488,N_15038,N_15001);
or U15489 (N_15489,N_15153,N_15158);
and U15490 (N_15490,N_15140,N_15178);
nand U15491 (N_15491,N_15051,N_15178);
nor U15492 (N_15492,N_15222,N_15235);
and U15493 (N_15493,N_15171,N_15158);
nor U15494 (N_15494,N_15016,N_15026);
nand U15495 (N_15495,N_15070,N_15182);
nand U15496 (N_15496,N_15167,N_15078);
nor U15497 (N_15497,N_15048,N_15173);
or U15498 (N_15498,N_15166,N_15061);
xor U15499 (N_15499,N_15020,N_15061);
or U15500 (N_15500,N_15283,N_15362);
and U15501 (N_15501,N_15303,N_15302);
nand U15502 (N_15502,N_15356,N_15458);
or U15503 (N_15503,N_15497,N_15288);
or U15504 (N_15504,N_15454,N_15471);
nor U15505 (N_15505,N_15460,N_15420);
nand U15506 (N_15506,N_15263,N_15364);
xnor U15507 (N_15507,N_15482,N_15278);
nor U15508 (N_15508,N_15404,N_15448);
or U15509 (N_15509,N_15439,N_15435);
nor U15510 (N_15510,N_15375,N_15333);
nor U15511 (N_15511,N_15436,N_15256);
xnor U15512 (N_15512,N_15253,N_15255);
nand U15513 (N_15513,N_15279,N_15261);
xnor U15514 (N_15514,N_15277,N_15344);
nor U15515 (N_15515,N_15337,N_15359);
xor U15516 (N_15516,N_15403,N_15257);
or U15517 (N_15517,N_15453,N_15352);
and U15518 (N_15518,N_15341,N_15347);
and U15519 (N_15519,N_15281,N_15293);
xnor U15520 (N_15520,N_15284,N_15473);
or U15521 (N_15521,N_15423,N_15402);
nand U15522 (N_15522,N_15319,N_15465);
nand U15523 (N_15523,N_15455,N_15363);
and U15524 (N_15524,N_15264,N_15373);
nand U15525 (N_15525,N_15414,N_15271);
nor U15526 (N_15526,N_15353,N_15400);
or U15527 (N_15527,N_15289,N_15331);
and U15528 (N_15528,N_15495,N_15450);
or U15529 (N_15529,N_15421,N_15412);
or U15530 (N_15530,N_15346,N_15348);
and U15531 (N_15531,N_15456,N_15317);
or U15532 (N_15532,N_15259,N_15358);
xnor U15533 (N_15533,N_15407,N_15382);
and U15534 (N_15534,N_15260,N_15372);
or U15535 (N_15535,N_15345,N_15472);
or U15536 (N_15536,N_15494,N_15273);
nand U15537 (N_15537,N_15387,N_15441);
and U15538 (N_15538,N_15308,N_15342);
xor U15539 (N_15539,N_15269,N_15286);
nor U15540 (N_15540,N_15469,N_15327);
nor U15541 (N_15541,N_15336,N_15328);
and U15542 (N_15542,N_15468,N_15315);
xor U15543 (N_15543,N_15295,N_15272);
xnor U15544 (N_15544,N_15451,N_15305);
nand U15545 (N_15545,N_15399,N_15434);
xnor U15546 (N_15546,N_15325,N_15300);
xor U15547 (N_15547,N_15401,N_15285);
nor U15548 (N_15548,N_15258,N_15408);
nor U15549 (N_15549,N_15266,N_15498);
or U15550 (N_15550,N_15367,N_15340);
nand U15551 (N_15551,N_15276,N_15318);
xor U15552 (N_15552,N_15416,N_15390);
nor U15553 (N_15553,N_15459,N_15312);
nor U15554 (N_15554,N_15488,N_15475);
nand U15555 (N_15555,N_15486,N_15332);
and U15556 (N_15556,N_15366,N_15313);
nand U15557 (N_15557,N_15395,N_15349);
nand U15558 (N_15558,N_15379,N_15483);
nor U15559 (N_15559,N_15419,N_15424);
nand U15560 (N_15560,N_15485,N_15389);
or U15561 (N_15561,N_15307,N_15357);
nand U15562 (N_15562,N_15368,N_15480);
nand U15563 (N_15563,N_15299,N_15490);
nand U15564 (N_15564,N_15351,N_15462);
nand U15565 (N_15565,N_15397,N_15445);
and U15566 (N_15566,N_15444,N_15426);
nor U15567 (N_15567,N_15323,N_15311);
xnor U15568 (N_15568,N_15374,N_15388);
nand U15569 (N_15569,N_15296,N_15411);
nand U15570 (N_15570,N_15415,N_15304);
xor U15571 (N_15571,N_15287,N_15447);
nor U15572 (N_15572,N_15355,N_15343);
and U15573 (N_15573,N_15291,N_15334);
or U15574 (N_15574,N_15492,N_15487);
nor U15575 (N_15575,N_15481,N_15298);
and U15576 (N_15576,N_15338,N_15437);
and U15577 (N_15577,N_15425,N_15377);
and U15578 (N_15578,N_15409,N_15470);
and U15579 (N_15579,N_15275,N_15282);
nand U15580 (N_15580,N_15392,N_15499);
xor U15581 (N_15581,N_15262,N_15265);
or U15582 (N_15582,N_15326,N_15427);
nor U15583 (N_15583,N_15443,N_15354);
nor U15584 (N_15584,N_15294,N_15383);
nor U15585 (N_15585,N_15446,N_15491);
or U15586 (N_15586,N_15370,N_15452);
nand U15587 (N_15587,N_15478,N_15314);
xnor U15588 (N_15588,N_15376,N_15474);
or U15589 (N_15589,N_15384,N_15385);
or U15590 (N_15590,N_15467,N_15489);
nand U15591 (N_15591,N_15422,N_15316);
and U15592 (N_15592,N_15393,N_15442);
nand U15593 (N_15593,N_15396,N_15496);
nand U15594 (N_15594,N_15322,N_15430);
nand U15595 (N_15595,N_15484,N_15321);
xnor U15596 (N_15596,N_15461,N_15309);
nand U15597 (N_15597,N_15330,N_15290);
xnor U15598 (N_15598,N_15405,N_15386);
xor U15599 (N_15599,N_15252,N_15438);
nand U15600 (N_15600,N_15413,N_15329);
nor U15601 (N_15601,N_15254,N_15274);
nand U15602 (N_15602,N_15350,N_15398);
or U15603 (N_15603,N_15466,N_15310);
and U15604 (N_15604,N_15391,N_15297);
nand U15605 (N_15605,N_15335,N_15464);
nand U15606 (N_15606,N_15250,N_15380);
nor U15607 (N_15607,N_15371,N_15418);
nor U15608 (N_15608,N_15477,N_15268);
and U15609 (N_15609,N_15394,N_15378);
xnor U15610 (N_15610,N_15433,N_15476);
xor U15611 (N_15611,N_15320,N_15428);
and U15612 (N_15612,N_15301,N_15493);
nor U15613 (N_15613,N_15365,N_15280);
and U15614 (N_15614,N_15369,N_15440);
or U15615 (N_15615,N_15292,N_15431);
or U15616 (N_15616,N_15406,N_15324);
nand U15617 (N_15617,N_15479,N_15360);
or U15618 (N_15618,N_15410,N_15381);
xor U15619 (N_15619,N_15449,N_15417);
xnor U15620 (N_15620,N_15429,N_15339);
and U15621 (N_15621,N_15457,N_15306);
nor U15622 (N_15622,N_15267,N_15270);
nand U15623 (N_15623,N_15361,N_15463);
and U15624 (N_15624,N_15432,N_15251);
xnor U15625 (N_15625,N_15361,N_15302);
nand U15626 (N_15626,N_15291,N_15486);
xnor U15627 (N_15627,N_15322,N_15268);
xnor U15628 (N_15628,N_15427,N_15476);
and U15629 (N_15629,N_15281,N_15384);
nor U15630 (N_15630,N_15255,N_15360);
nand U15631 (N_15631,N_15443,N_15481);
or U15632 (N_15632,N_15251,N_15349);
nor U15633 (N_15633,N_15303,N_15349);
xor U15634 (N_15634,N_15447,N_15460);
nand U15635 (N_15635,N_15333,N_15348);
xnor U15636 (N_15636,N_15434,N_15454);
or U15637 (N_15637,N_15258,N_15343);
nand U15638 (N_15638,N_15283,N_15388);
xor U15639 (N_15639,N_15297,N_15474);
nor U15640 (N_15640,N_15419,N_15427);
and U15641 (N_15641,N_15394,N_15319);
nand U15642 (N_15642,N_15416,N_15297);
or U15643 (N_15643,N_15363,N_15463);
and U15644 (N_15644,N_15447,N_15370);
or U15645 (N_15645,N_15468,N_15425);
or U15646 (N_15646,N_15284,N_15267);
or U15647 (N_15647,N_15405,N_15331);
nor U15648 (N_15648,N_15451,N_15338);
nand U15649 (N_15649,N_15286,N_15352);
or U15650 (N_15650,N_15499,N_15373);
nor U15651 (N_15651,N_15475,N_15330);
nor U15652 (N_15652,N_15337,N_15331);
or U15653 (N_15653,N_15351,N_15400);
or U15654 (N_15654,N_15463,N_15404);
xor U15655 (N_15655,N_15264,N_15491);
and U15656 (N_15656,N_15332,N_15450);
xor U15657 (N_15657,N_15478,N_15464);
or U15658 (N_15658,N_15484,N_15256);
nand U15659 (N_15659,N_15358,N_15308);
and U15660 (N_15660,N_15424,N_15316);
nor U15661 (N_15661,N_15306,N_15324);
or U15662 (N_15662,N_15425,N_15319);
and U15663 (N_15663,N_15250,N_15444);
and U15664 (N_15664,N_15419,N_15270);
or U15665 (N_15665,N_15461,N_15467);
xor U15666 (N_15666,N_15462,N_15375);
xnor U15667 (N_15667,N_15489,N_15351);
or U15668 (N_15668,N_15338,N_15334);
xor U15669 (N_15669,N_15259,N_15318);
and U15670 (N_15670,N_15263,N_15475);
nor U15671 (N_15671,N_15293,N_15358);
or U15672 (N_15672,N_15344,N_15359);
nand U15673 (N_15673,N_15423,N_15336);
nand U15674 (N_15674,N_15276,N_15385);
nand U15675 (N_15675,N_15253,N_15314);
xnor U15676 (N_15676,N_15276,N_15336);
xor U15677 (N_15677,N_15257,N_15481);
nand U15678 (N_15678,N_15398,N_15335);
nand U15679 (N_15679,N_15407,N_15351);
and U15680 (N_15680,N_15310,N_15336);
and U15681 (N_15681,N_15365,N_15397);
nor U15682 (N_15682,N_15367,N_15288);
nor U15683 (N_15683,N_15321,N_15309);
and U15684 (N_15684,N_15333,N_15457);
xor U15685 (N_15685,N_15272,N_15322);
and U15686 (N_15686,N_15305,N_15276);
nor U15687 (N_15687,N_15498,N_15422);
or U15688 (N_15688,N_15259,N_15268);
nor U15689 (N_15689,N_15283,N_15327);
xor U15690 (N_15690,N_15427,N_15455);
nand U15691 (N_15691,N_15342,N_15409);
nand U15692 (N_15692,N_15362,N_15487);
nor U15693 (N_15693,N_15483,N_15423);
nand U15694 (N_15694,N_15426,N_15317);
and U15695 (N_15695,N_15417,N_15341);
or U15696 (N_15696,N_15368,N_15414);
nand U15697 (N_15697,N_15371,N_15498);
nor U15698 (N_15698,N_15287,N_15304);
and U15699 (N_15699,N_15470,N_15416);
nor U15700 (N_15700,N_15334,N_15329);
nand U15701 (N_15701,N_15405,N_15371);
and U15702 (N_15702,N_15379,N_15296);
or U15703 (N_15703,N_15402,N_15392);
nor U15704 (N_15704,N_15294,N_15351);
and U15705 (N_15705,N_15377,N_15363);
and U15706 (N_15706,N_15340,N_15298);
nor U15707 (N_15707,N_15465,N_15279);
nand U15708 (N_15708,N_15370,N_15393);
nor U15709 (N_15709,N_15461,N_15364);
nand U15710 (N_15710,N_15290,N_15389);
nand U15711 (N_15711,N_15367,N_15382);
and U15712 (N_15712,N_15398,N_15473);
nor U15713 (N_15713,N_15441,N_15405);
nor U15714 (N_15714,N_15273,N_15257);
and U15715 (N_15715,N_15457,N_15323);
xor U15716 (N_15716,N_15409,N_15272);
xnor U15717 (N_15717,N_15253,N_15451);
nand U15718 (N_15718,N_15287,N_15274);
and U15719 (N_15719,N_15382,N_15335);
or U15720 (N_15720,N_15403,N_15415);
or U15721 (N_15721,N_15462,N_15423);
nand U15722 (N_15722,N_15298,N_15296);
nand U15723 (N_15723,N_15494,N_15405);
or U15724 (N_15724,N_15484,N_15373);
xor U15725 (N_15725,N_15495,N_15256);
xnor U15726 (N_15726,N_15496,N_15422);
nor U15727 (N_15727,N_15432,N_15357);
or U15728 (N_15728,N_15396,N_15287);
nand U15729 (N_15729,N_15259,N_15343);
or U15730 (N_15730,N_15390,N_15267);
nor U15731 (N_15731,N_15353,N_15420);
xor U15732 (N_15732,N_15346,N_15401);
and U15733 (N_15733,N_15470,N_15336);
or U15734 (N_15734,N_15492,N_15458);
or U15735 (N_15735,N_15497,N_15362);
or U15736 (N_15736,N_15397,N_15336);
nand U15737 (N_15737,N_15474,N_15492);
xor U15738 (N_15738,N_15386,N_15410);
xnor U15739 (N_15739,N_15386,N_15284);
nor U15740 (N_15740,N_15478,N_15287);
xor U15741 (N_15741,N_15269,N_15384);
or U15742 (N_15742,N_15449,N_15422);
nand U15743 (N_15743,N_15394,N_15495);
xor U15744 (N_15744,N_15318,N_15381);
and U15745 (N_15745,N_15343,N_15406);
nor U15746 (N_15746,N_15264,N_15450);
nor U15747 (N_15747,N_15447,N_15250);
or U15748 (N_15748,N_15407,N_15253);
nor U15749 (N_15749,N_15272,N_15357);
and U15750 (N_15750,N_15574,N_15652);
nand U15751 (N_15751,N_15658,N_15628);
nand U15752 (N_15752,N_15743,N_15533);
nor U15753 (N_15753,N_15611,N_15716);
nor U15754 (N_15754,N_15728,N_15580);
nor U15755 (N_15755,N_15646,N_15665);
or U15756 (N_15756,N_15571,N_15702);
nor U15757 (N_15757,N_15562,N_15518);
nor U15758 (N_15758,N_15714,N_15503);
xor U15759 (N_15759,N_15729,N_15688);
or U15760 (N_15760,N_15553,N_15519);
nor U15761 (N_15761,N_15620,N_15726);
nor U15762 (N_15762,N_15635,N_15501);
nand U15763 (N_15763,N_15584,N_15661);
nor U15764 (N_15764,N_15520,N_15672);
nor U15765 (N_15765,N_15737,N_15685);
nor U15766 (N_15766,N_15720,N_15730);
and U15767 (N_15767,N_15511,N_15698);
nand U15768 (N_15768,N_15670,N_15565);
and U15769 (N_15769,N_15576,N_15634);
nor U15770 (N_15770,N_15554,N_15722);
xor U15771 (N_15771,N_15724,N_15595);
xor U15772 (N_15772,N_15616,N_15640);
nand U15773 (N_15773,N_15542,N_15594);
and U15774 (N_15774,N_15650,N_15684);
or U15775 (N_15775,N_15683,N_15559);
xor U15776 (N_15776,N_15669,N_15693);
xor U15777 (N_15777,N_15551,N_15596);
nand U15778 (N_15778,N_15514,N_15541);
and U15779 (N_15779,N_15641,N_15675);
and U15780 (N_15780,N_15526,N_15686);
or U15781 (N_15781,N_15626,N_15638);
nor U15782 (N_15782,N_15515,N_15709);
nor U15783 (N_15783,N_15528,N_15599);
nand U15784 (N_15784,N_15648,N_15667);
or U15785 (N_15785,N_15598,N_15746);
nand U15786 (N_15786,N_15593,N_15677);
nand U15787 (N_15787,N_15622,N_15555);
nor U15788 (N_15788,N_15711,N_15703);
nand U15789 (N_15789,N_15549,N_15653);
nor U15790 (N_15790,N_15657,N_15521);
and U15791 (N_15791,N_15681,N_15749);
nand U15792 (N_15792,N_15539,N_15631);
or U15793 (N_15793,N_15727,N_15655);
or U15794 (N_15794,N_15505,N_15673);
xor U15795 (N_15795,N_15609,N_15664);
nor U15796 (N_15796,N_15567,N_15570);
nand U15797 (N_15797,N_15632,N_15668);
nor U15798 (N_15798,N_15605,N_15630);
or U15799 (N_15799,N_15617,N_15556);
nor U15800 (N_15800,N_15610,N_15591);
nand U15801 (N_15801,N_15546,N_15715);
xor U15802 (N_15802,N_15687,N_15557);
and U15803 (N_15803,N_15597,N_15525);
and U15804 (N_15804,N_15608,N_15507);
or U15805 (N_15805,N_15568,N_15659);
or U15806 (N_15806,N_15572,N_15705);
nand U15807 (N_15807,N_15740,N_15625);
and U15808 (N_15808,N_15732,N_15600);
nor U15809 (N_15809,N_15619,N_15624);
and U15810 (N_15810,N_15540,N_15585);
or U15811 (N_15811,N_15569,N_15535);
and U15812 (N_15812,N_15654,N_15536);
nor U15813 (N_15813,N_15586,N_15575);
and U15814 (N_15814,N_15582,N_15679);
nand U15815 (N_15815,N_15723,N_15674);
and U15816 (N_15816,N_15708,N_15721);
or U15817 (N_15817,N_15642,N_15736);
and U15818 (N_15818,N_15629,N_15623);
nand U15819 (N_15819,N_15590,N_15548);
xnor U15820 (N_15820,N_15747,N_15671);
nand U15821 (N_15821,N_15607,N_15508);
nor U15822 (N_15822,N_15742,N_15516);
nand U15823 (N_15823,N_15573,N_15717);
nor U15824 (N_15824,N_15602,N_15500);
xor U15825 (N_15825,N_15697,N_15738);
or U15826 (N_15826,N_15560,N_15510);
xnor U15827 (N_15827,N_15538,N_15627);
and U15828 (N_15828,N_15700,N_15577);
and U15829 (N_15829,N_15731,N_15550);
and U15830 (N_15830,N_15509,N_15660);
nor U15831 (N_15831,N_15618,N_15592);
nand U15832 (N_15832,N_15547,N_15523);
and U15833 (N_15833,N_15601,N_15578);
and U15834 (N_15834,N_15537,N_15522);
xnor U15835 (N_15835,N_15706,N_15643);
nand U15836 (N_15836,N_15707,N_15713);
xnor U15837 (N_15837,N_15682,N_15531);
or U15838 (N_15838,N_15566,N_15695);
and U15839 (N_15839,N_15645,N_15666);
and U15840 (N_15840,N_15699,N_15603);
and U15841 (N_15841,N_15558,N_15587);
xnor U15842 (N_15842,N_15637,N_15636);
or U15843 (N_15843,N_15543,N_15739);
nor U15844 (N_15844,N_15678,N_15502);
nand U15845 (N_15845,N_15690,N_15614);
nand U15846 (N_15846,N_15589,N_15529);
xnor U15847 (N_15847,N_15544,N_15734);
and U15848 (N_15848,N_15725,N_15621);
nand U15849 (N_15849,N_15748,N_15662);
or U15850 (N_15850,N_15689,N_15741);
xor U15851 (N_15851,N_15563,N_15676);
and U15852 (N_15852,N_15692,N_15710);
or U15853 (N_15853,N_15561,N_15581);
or U15854 (N_15854,N_15696,N_15691);
or U15855 (N_15855,N_15588,N_15583);
and U15856 (N_15856,N_15504,N_15649);
nor U15857 (N_15857,N_15656,N_15644);
and U15858 (N_15858,N_15506,N_15647);
nor U15859 (N_15859,N_15534,N_15524);
and U15860 (N_15860,N_15663,N_15704);
or U15861 (N_15861,N_15606,N_15517);
and U15862 (N_15862,N_15633,N_15512);
xor U15863 (N_15863,N_15612,N_15718);
nor U15864 (N_15864,N_15744,N_15530);
nor U15865 (N_15865,N_15639,N_15527);
nor U15866 (N_15866,N_15545,N_15513);
nand U15867 (N_15867,N_15613,N_15615);
nor U15868 (N_15868,N_15680,N_15701);
xor U15869 (N_15869,N_15579,N_15604);
xor U15870 (N_15870,N_15733,N_15745);
nand U15871 (N_15871,N_15694,N_15532);
nand U15872 (N_15872,N_15564,N_15719);
nand U15873 (N_15873,N_15712,N_15735);
or U15874 (N_15874,N_15651,N_15552);
nor U15875 (N_15875,N_15692,N_15724);
xor U15876 (N_15876,N_15626,N_15739);
nand U15877 (N_15877,N_15656,N_15617);
and U15878 (N_15878,N_15738,N_15527);
xnor U15879 (N_15879,N_15553,N_15637);
xnor U15880 (N_15880,N_15655,N_15692);
nand U15881 (N_15881,N_15698,N_15611);
nor U15882 (N_15882,N_15697,N_15544);
nand U15883 (N_15883,N_15692,N_15733);
nand U15884 (N_15884,N_15618,N_15537);
nand U15885 (N_15885,N_15592,N_15732);
or U15886 (N_15886,N_15719,N_15520);
nand U15887 (N_15887,N_15505,N_15715);
xnor U15888 (N_15888,N_15620,N_15574);
or U15889 (N_15889,N_15531,N_15694);
nor U15890 (N_15890,N_15562,N_15560);
nor U15891 (N_15891,N_15655,N_15702);
and U15892 (N_15892,N_15708,N_15704);
nand U15893 (N_15893,N_15718,N_15632);
and U15894 (N_15894,N_15669,N_15642);
and U15895 (N_15895,N_15604,N_15542);
and U15896 (N_15896,N_15639,N_15530);
nand U15897 (N_15897,N_15570,N_15516);
xnor U15898 (N_15898,N_15625,N_15749);
xnor U15899 (N_15899,N_15606,N_15541);
or U15900 (N_15900,N_15736,N_15662);
xnor U15901 (N_15901,N_15557,N_15727);
nor U15902 (N_15902,N_15656,N_15738);
nor U15903 (N_15903,N_15520,N_15572);
nor U15904 (N_15904,N_15630,N_15731);
xnor U15905 (N_15905,N_15642,N_15501);
nand U15906 (N_15906,N_15712,N_15608);
or U15907 (N_15907,N_15650,N_15743);
nand U15908 (N_15908,N_15621,N_15722);
nor U15909 (N_15909,N_15573,N_15726);
xnor U15910 (N_15910,N_15518,N_15640);
nand U15911 (N_15911,N_15694,N_15730);
nor U15912 (N_15912,N_15702,N_15686);
nor U15913 (N_15913,N_15538,N_15658);
or U15914 (N_15914,N_15546,N_15680);
nor U15915 (N_15915,N_15681,N_15645);
nor U15916 (N_15916,N_15674,N_15631);
or U15917 (N_15917,N_15584,N_15586);
nand U15918 (N_15918,N_15557,N_15718);
nand U15919 (N_15919,N_15645,N_15715);
and U15920 (N_15920,N_15719,N_15545);
nor U15921 (N_15921,N_15665,N_15507);
xor U15922 (N_15922,N_15626,N_15624);
nor U15923 (N_15923,N_15697,N_15611);
nor U15924 (N_15924,N_15675,N_15663);
or U15925 (N_15925,N_15523,N_15632);
nand U15926 (N_15926,N_15737,N_15722);
and U15927 (N_15927,N_15747,N_15646);
nor U15928 (N_15928,N_15708,N_15576);
xnor U15929 (N_15929,N_15531,N_15678);
nand U15930 (N_15930,N_15592,N_15696);
nand U15931 (N_15931,N_15530,N_15581);
nand U15932 (N_15932,N_15631,N_15732);
nor U15933 (N_15933,N_15524,N_15509);
nand U15934 (N_15934,N_15720,N_15721);
nor U15935 (N_15935,N_15613,N_15595);
xnor U15936 (N_15936,N_15624,N_15584);
nor U15937 (N_15937,N_15709,N_15608);
and U15938 (N_15938,N_15637,N_15704);
and U15939 (N_15939,N_15516,N_15625);
or U15940 (N_15940,N_15645,N_15530);
and U15941 (N_15941,N_15642,N_15589);
or U15942 (N_15942,N_15510,N_15539);
and U15943 (N_15943,N_15743,N_15675);
xor U15944 (N_15944,N_15647,N_15618);
nand U15945 (N_15945,N_15546,N_15740);
xor U15946 (N_15946,N_15560,N_15670);
and U15947 (N_15947,N_15657,N_15730);
nand U15948 (N_15948,N_15675,N_15519);
or U15949 (N_15949,N_15593,N_15517);
nand U15950 (N_15950,N_15605,N_15662);
nand U15951 (N_15951,N_15551,N_15705);
nand U15952 (N_15952,N_15538,N_15686);
nor U15953 (N_15953,N_15567,N_15689);
nor U15954 (N_15954,N_15743,N_15614);
xor U15955 (N_15955,N_15565,N_15696);
nor U15956 (N_15956,N_15745,N_15528);
xnor U15957 (N_15957,N_15532,N_15518);
xor U15958 (N_15958,N_15687,N_15591);
nand U15959 (N_15959,N_15507,N_15619);
or U15960 (N_15960,N_15686,N_15595);
nand U15961 (N_15961,N_15644,N_15633);
nand U15962 (N_15962,N_15611,N_15706);
nor U15963 (N_15963,N_15655,N_15659);
and U15964 (N_15964,N_15730,N_15710);
or U15965 (N_15965,N_15568,N_15685);
nand U15966 (N_15966,N_15535,N_15675);
xor U15967 (N_15967,N_15601,N_15506);
nand U15968 (N_15968,N_15592,N_15632);
nor U15969 (N_15969,N_15524,N_15705);
nand U15970 (N_15970,N_15583,N_15621);
or U15971 (N_15971,N_15644,N_15647);
and U15972 (N_15972,N_15734,N_15578);
or U15973 (N_15973,N_15724,N_15549);
nand U15974 (N_15974,N_15651,N_15573);
and U15975 (N_15975,N_15562,N_15516);
and U15976 (N_15976,N_15691,N_15605);
nand U15977 (N_15977,N_15520,N_15524);
nand U15978 (N_15978,N_15614,N_15584);
or U15979 (N_15979,N_15512,N_15513);
and U15980 (N_15980,N_15740,N_15731);
or U15981 (N_15981,N_15626,N_15667);
and U15982 (N_15982,N_15512,N_15717);
nor U15983 (N_15983,N_15640,N_15678);
and U15984 (N_15984,N_15529,N_15601);
or U15985 (N_15985,N_15722,N_15693);
nor U15986 (N_15986,N_15502,N_15606);
or U15987 (N_15987,N_15632,N_15570);
or U15988 (N_15988,N_15668,N_15748);
nand U15989 (N_15989,N_15656,N_15634);
or U15990 (N_15990,N_15736,N_15716);
or U15991 (N_15991,N_15738,N_15518);
xnor U15992 (N_15992,N_15565,N_15690);
and U15993 (N_15993,N_15588,N_15514);
xnor U15994 (N_15994,N_15546,N_15627);
and U15995 (N_15995,N_15545,N_15643);
xnor U15996 (N_15996,N_15743,N_15563);
and U15997 (N_15997,N_15743,N_15674);
or U15998 (N_15998,N_15743,N_15623);
and U15999 (N_15999,N_15525,N_15523);
nor U16000 (N_16000,N_15888,N_15829);
nand U16001 (N_16001,N_15795,N_15814);
nor U16002 (N_16002,N_15753,N_15770);
xor U16003 (N_16003,N_15982,N_15916);
or U16004 (N_16004,N_15782,N_15933);
xor U16005 (N_16005,N_15858,N_15867);
and U16006 (N_16006,N_15785,N_15840);
or U16007 (N_16007,N_15882,N_15994);
and U16008 (N_16008,N_15959,N_15799);
and U16009 (N_16009,N_15809,N_15775);
xnor U16010 (N_16010,N_15844,N_15854);
nor U16011 (N_16011,N_15927,N_15750);
nor U16012 (N_16012,N_15804,N_15958);
xor U16013 (N_16013,N_15996,N_15884);
and U16014 (N_16014,N_15957,N_15988);
and U16015 (N_16015,N_15987,N_15922);
nand U16016 (N_16016,N_15903,N_15900);
xor U16017 (N_16017,N_15760,N_15962);
or U16018 (N_16018,N_15848,N_15998);
or U16019 (N_16019,N_15960,N_15792);
nor U16020 (N_16020,N_15909,N_15934);
xor U16021 (N_16021,N_15872,N_15952);
or U16022 (N_16022,N_15920,N_15774);
nand U16023 (N_16023,N_15947,N_15802);
xor U16024 (N_16024,N_15805,N_15978);
or U16025 (N_16025,N_15965,N_15865);
nand U16026 (N_16026,N_15967,N_15945);
nor U16027 (N_16027,N_15949,N_15816);
or U16028 (N_16028,N_15855,N_15779);
and U16029 (N_16029,N_15905,N_15932);
nor U16030 (N_16030,N_15915,N_15863);
and U16031 (N_16031,N_15851,N_15828);
nor U16032 (N_16032,N_15755,N_15917);
xor U16033 (N_16033,N_15820,N_15811);
nor U16034 (N_16034,N_15997,N_15860);
and U16035 (N_16035,N_15800,N_15845);
or U16036 (N_16036,N_15789,N_15861);
and U16037 (N_16037,N_15758,N_15793);
nor U16038 (N_16038,N_15822,N_15798);
xnor U16039 (N_16039,N_15918,N_15853);
nand U16040 (N_16040,N_15846,N_15899);
nand U16041 (N_16041,N_15788,N_15910);
and U16042 (N_16042,N_15810,N_15906);
nor U16043 (N_16043,N_15943,N_15842);
nand U16044 (N_16044,N_15914,N_15875);
xnor U16045 (N_16045,N_15921,N_15951);
nand U16046 (N_16046,N_15904,N_15819);
or U16047 (N_16047,N_15936,N_15847);
xnor U16048 (N_16048,N_15870,N_15826);
or U16049 (N_16049,N_15776,N_15821);
and U16050 (N_16050,N_15874,N_15806);
nand U16051 (N_16051,N_15857,N_15955);
xnor U16052 (N_16052,N_15878,N_15912);
xnor U16053 (N_16053,N_15838,N_15803);
nor U16054 (N_16054,N_15999,N_15834);
or U16055 (N_16055,N_15784,N_15891);
xor U16056 (N_16056,N_15893,N_15754);
xor U16057 (N_16057,N_15931,N_15971);
and U16058 (N_16058,N_15898,N_15954);
nand U16059 (N_16059,N_15963,N_15813);
nand U16060 (N_16060,N_15968,N_15991);
nand U16061 (N_16061,N_15777,N_15969);
or U16062 (N_16062,N_15975,N_15972);
or U16063 (N_16063,N_15825,N_15790);
and U16064 (N_16064,N_15796,N_15924);
and U16065 (N_16065,N_15769,N_15794);
nand U16066 (N_16066,N_15974,N_15923);
xnor U16067 (N_16067,N_15892,N_15946);
xor U16068 (N_16068,N_15977,N_15986);
and U16069 (N_16069,N_15866,N_15895);
xnor U16070 (N_16070,N_15756,N_15817);
nand U16071 (N_16071,N_15877,N_15993);
nand U16072 (N_16072,N_15812,N_15768);
nor U16073 (N_16073,N_15757,N_15856);
or U16074 (N_16074,N_15902,N_15890);
nand U16075 (N_16075,N_15765,N_15979);
xor U16076 (N_16076,N_15983,N_15956);
nand U16077 (N_16077,N_15764,N_15989);
nor U16078 (N_16078,N_15935,N_15752);
nor U16079 (N_16079,N_15911,N_15832);
and U16080 (N_16080,N_15850,N_15873);
xnor U16081 (N_16081,N_15907,N_15767);
xnor U16082 (N_16082,N_15984,N_15852);
nor U16083 (N_16083,N_15885,N_15761);
or U16084 (N_16084,N_15886,N_15980);
nand U16085 (N_16085,N_15849,N_15778);
and U16086 (N_16086,N_15901,N_15837);
and U16087 (N_16087,N_15771,N_15773);
or U16088 (N_16088,N_15781,N_15883);
xnor U16089 (N_16089,N_15880,N_15869);
nor U16090 (N_16090,N_15862,N_15818);
xor U16091 (N_16091,N_15990,N_15889);
nand U16092 (N_16092,N_15876,N_15836);
xnor U16093 (N_16093,N_15926,N_15783);
nand U16094 (N_16094,N_15940,N_15944);
nand U16095 (N_16095,N_15887,N_15808);
nor U16096 (N_16096,N_15827,N_15970);
nor U16097 (N_16097,N_15995,N_15868);
nor U16098 (N_16098,N_15896,N_15928);
nand U16099 (N_16099,N_15937,N_15992);
and U16100 (N_16100,N_15973,N_15823);
or U16101 (N_16101,N_15966,N_15762);
xnor U16102 (N_16102,N_15835,N_15941);
xnor U16103 (N_16103,N_15831,N_15950);
nand U16104 (N_16104,N_15859,N_15791);
or U16105 (N_16105,N_15929,N_15864);
xor U16106 (N_16106,N_15763,N_15985);
or U16107 (N_16107,N_15981,N_15913);
or U16108 (N_16108,N_15879,N_15830);
nand U16109 (N_16109,N_15772,N_15797);
or U16110 (N_16110,N_15787,N_15833);
and U16111 (N_16111,N_15839,N_15801);
xnor U16112 (N_16112,N_15925,N_15897);
nand U16113 (N_16113,N_15964,N_15786);
nand U16114 (N_16114,N_15815,N_15953);
nand U16115 (N_16115,N_15780,N_15824);
and U16116 (N_16116,N_15942,N_15938);
and U16117 (N_16117,N_15759,N_15930);
and U16118 (N_16118,N_15948,N_15919);
or U16119 (N_16119,N_15939,N_15976);
or U16120 (N_16120,N_15751,N_15841);
nor U16121 (N_16121,N_15843,N_15961);
nand U16122 (N_16122,N_15766,N_15908);
and U16123 (N_16123,N_15871,N_15894);
or U16124 (N_16124,N_15807,N_15881);
or U16125 (N_16125,N_15993,N_15961);
and U16126 (N_16126,N_15967,N_15833);
and U16127 (N_16127,N_15938,N_15821);
nand U16128 (N_16128,N_15798,N_15843);
or U16129 (N_16129,N_15863,N_15923);
xnor U16130 (N_16130,N_15823,N_15858);
xnor U16131 (N_16131,N_15809,N_15953);
and U16132 (N_16132,N_15755,N_15946);
nor U16133 (N_16133,N_15841,N_15822);
nor U16134 (N_16134,N_15756,N_15797);
xor U16135 (N_16135,N_15779,N_15845);
or U16136 (N_16136,N_15754,N_15888);
and U16137 (N_16137,N_15771,N_15901);
and U16138 (N_16138,N_15962,N_15967);
nor U16139 (N_16139,N_15975,N_15898);
xor U16140 (N_16140,N_15959,N_15797);
and U16141 (N_16141,N_15950,N_15840);
and U16142 (N_16142,N_15827,N_15930);
nand U16143 (N_16143,N_15983,N_15789);
or U16144 (N_16144,N_15808,N_15881);
and U16145 (N_16145,N_15907,N_15901);
xor U16146 (N_16146,N_15908,N_15786);
and U16147 (N_16147,N_15920,N_15893);
or U16148 (N_16148,N_15796,N_15897);
xnor U16149 (N_16149,N_15996,N_15979);
and U16150 (N_16150,N_15887,N_15834);
nor U16151 (N_16151,N_15795,N_15833);
or U16152 (N_16152,N_15886,N_15910);
or U16153 (N_16153,N_15758,N_15810);
xnor U16154 (N_16154,N_15987,N_15945);
xor U16155 (N_16155,N_15764,N_15886);
nor U16156 (N_16156,N_15828,N_15955);
and U16157 (N_16157,N_15763,N_15902);
nor U16158 (N_16158,N_15811,N_15987);
and U16159 (N_16159,N_15880,N_15876);
nand U16160 (N_16160,N_15830,N_15987);
and U16161 (N_16161,N_15977,N_15946);
xnor U16162 (N_16162,N_15866,N_15928);
xor U16163 (N_16163,N_15808,N_15984);
xnor U16164 (N_16164,N_15872,N_15838);
nand U16165 (N_16165,N_15971,N_15854);
xor U16166 (N_16166,N_15917,N_15776);
xnor U16167 (N_16167,N_15898,N_15921);
and U16168 (N_16168,N_15976,N_15834);
and U16169 (N_16169,N_15916,N_15826);
xor U16170 (N_16170,N_15875,N_15766);
nand U16171 (N_16171,N_15803,N_15872);
nor U16172 (N_16172,N_15990,N_15772);
xor U16173 (N_16173,N_15942,N_15794);
or U16174 (N_16174,N_15836,N_15890);
or U16175 (N_16175,N_15936,N_15962);
xor U16176 (N_16176,N_15922,N_15876);
or U16177 (N_16177,N_15854,N_15950);
nand U16178 (N_16178,N_15900,N_15904);
nor U16179 (N_16179,N_15926,N_15958);
nand U16180 (N_16180,N_15869,N_15936);
and U16181 (N_16181,N_15895,N_15995);
nand U16182 (N_16182,N_15923,N_15801);
and U16183 (N_16183,N_15883,N_15783);
or U16184 (N_16184,N_15795,N_15878);
xnor U16185 (N_16185,N_15898,N_15838);
xor U16186 (N_16186,N_15940,N_15981);
nor U16187 (N_16187,N_15838,N_15815);
xor U16188 (N_16188,N_15799,N_15845);
xnor U16189 (N_16189,N_15889,N_15944);
nand U16190 (N_16190,N_15890,N_15939);
xor U16191 (N_16191,N_15765,N_15912);
xor U16192 (N_16192,N_15951,N_15883);
nand U16193 (N_16193,N_15879,N_15824);
xor U16194 (N_16194,N_15952,N_15871);
or U16195 (N_16195,N_15909,N_15940);
xor U16196 (N_16196,N_15804,N_15781);
nor U16197 (N_16197,N_15922,N_15990);
nor U16198 (N_16198,N_15857,N_15797);
nor U16199 (N_16199,N_15817,N_15980);
nor U16200 (N_16200,N_15978,N_15804);
and U16201 (N_16201,N_15784,N_15792);
nor U16202 (N_16202,N_15980,N_15820);
and U16203 (N_16203,N_15774,N_15824);
nand U16204 (N_16204,N_15833,N_15778);
nor U16205 (N_16205,N_15829,N_15970);
and U16206 (N_16206,N_15974,N_15933);
nand U16207 (N_16207,N_15854,N_15988);
xnor U16208 (N_16208,N_15942,N_15967);
nand U16209 (N_16209,N_15803,N_15841);
nor U16210 (N_16210,N_15994,N_15806);
or U16211 (N_16211,N_15871,N_15758);
nor U16212 (N_16212,N_15995,N_15943);
xor U16213 (N_16213,N_15910,N_15809);
nor U16214 (N_16214,N_15897,N_15818);
or U16215 (N_16215,N_15908,N_15951);
nand U16216 (N_16216,N_15900,N_15977);
nor U16217 (N_16217,N_15893,N_15953);
or U16218 (N_16218,N_15957,N_15900);
or U16219 (N_16219,N_15849,N_15822);
nand U16220 (N_16220,N_15875,N_15994);
xnor U16221 (N_16221,N_15876,N_15797);
nor U16222 (N_16222,N_15936,N_15961);
or U16223 (N_16223,N_15967,N_15768);
or U16224 (N_16224,N_15951,N_15863);
and U16225 (N_16225,N_15854,N_15896);
xnor U16226 (N_16226,N_15924,N_15968);
xnor U16227 (N_16227,N_15882,N_15811);
xor U16228 (N_16228,N_15897,N_15841);
or U16229 (N_16229,N_15914,N_15911);
and U16230 (N_16230,N_15862,N_15918);
or U16231 (N_16231,N_15804,N_15912);
nor U16232 (N_16232,N_15975,N_15754);
xnor U16233 (N_16233,N_15814,N_15871);
nand U16234 (N_16234,N_15994,N_15758);
nand U16235 (N_16235,N_15882,N_15787);
and U16236 (N_16236,N_15872,N_15770);
and U16237 (N_16237,N_15845,N_15863);
or U16238 (N_16238,N_15988,N_15769);
xor U16239 (N_16239,N_15909,N_15886);
nor U16240 (N_16240,N_15770,N_15994);
xor U16241 (N_16241,N_15864,N_15784);
or U16242 (N_16242,N_15750,N_15765);
nor U16243 (N_16243,N_15891,N_15844);
or U16244 (N_16244,N_15841,N_15781);
nor U16245 (N_16245,N_15856,N_15885);
and U16246 (N_16246,N_15904,N_15941);
nand U16247 (N_16247,N_15825,N_15996);
nor U16248 (N_16248,N_15825,N_15856);
nor U16249 (N_16249,N_15753,N_15798);
nor U16250 (N_16250,N_16219,N_16160);
nor U16251 (N_16251,N_16002,N_16006);
nor U16252 (N_16252,N_16070,N_16063);
xor U16253 (N_16253,N_16134,N_16238);
nor U16254 (N_16254,N_16066,N_16192);
and U16255 (N_16255,N_16039,N_16045);
and U16256 (N_16256,N_16012,N_16175);
xnor U16257 (N_16257,N_16051,N_16162);
nor U16258 (N_16258,N_16170,N_16201);
or U16259 (N_16259,N_16044,N_16123);
xor U16260 (N_16260,N_16004,N_16114);
xnor U16261 (N_16261,N_16043,N_16141);
nor U16262 (N_16262,N_16125,N_16229);
xor U16263 (N_16263,N_16231,N_16245);
and U16264 (N_16264,N_16020,N_16092);
nor U16265 (N_16265,N_16139,N_16240);
and U16266 (N_16266,N_16164,N_16237);
xnor U16267 (N_16267,N_16146,N_16111);
and U16268 (N_16268,N_16076,N_16007);
nand U16269 (N_16269,N_16227,N_16163);
nand U16270 (N_16270,N_16143,N_16179);
xnor U16271 (N_16271,N_16084,N_16106);
nor U16272 (N_16272,N_16119,N_16078);
nor U16273 (N_16273,N_16053,N_16195);
nand U16274 (N_16274,N_16133,N_16248);
xor U16275 (N_16275,N_16234,N_16249);
nand U16276 (N_16276,N_16060,N_16048);
or U16277 (N_16277,N_16242,N_16069);
or U16278 (N_16278,N_16176,N_16015);
and U16279 (N_16279,N_16224,N_16103);
or U16280 (N_16280,N_16050,N_16049);
and U16281 (N_16281,N_16117,N_16064);
xor U16282 (N_16282,N_16140,N_16009);
nor U16283 (N_16283,N_16244,N_16135);
and U16284 (N_16284,N_16035,N_16191);
or U16285 (N_16285,N_16096,N_16113);
and U16286 (N_16286,N_16173,N_16216);
xnor U16287 (N_16287,N_16052,N_16230);
nor U16288 (N_16288,N_16079,N_16054);
xnor U16289 (N_16289,N_16088,N_16178);
nand U16290 (N_16290,N_16055,N_16131);
or U16291 (N_16291,N_16110,N_16025);
or U16292 (N_16292,N_16034,N_16129);
nand U16293 (N_16293,N_16213,N_16124);
nor U16294 (N_16294,N_16165,N_16152);
nand U16295 (N_16295,N_16183,N_16174);
nand U16296 (N_16296,N_16190,N_16104);
or U16297 (N_16297,N_16075,N_16217);
and U16298 (N_16298,N_16130,N_16057);
nand U16299 (N_16299,N_16046,N_16072);
nand U16300 (N_16300,N_16067,N_16241);
xnor U16301 (N_16301,N_16225,N_16246);
or U16302 (N_16302,N_16109,N_16065);
or U16303 (N_16303,N_16196,N_16161);
nor U16304 (N_16304,N_16085,N_16108);
and U16305 (N_16305,N_16086,N_16062);
nor U16306 (N_16306,N_16132,N_16040);
or U16307 (N_16307,N_16080,N_16024);
and U16308 (N_16308,N_16013,N_16121);
or U16309 (N_16309,N_16222,N_16107);
nand U16310 (N_16310,N_16159,N_16010);
or U16311 (N_16311,N_16148,N_16014);
nand U16312 (N_16312,N_16029,N_16042);
xor U16313 (N_16313,N_16099,N_16228);
or U16314 (N_16314,N_16027,N_16171);
nand U16315 (N_16315,N_16188,N_16184);
nor U16316 (N_16316,N_16239,N_16037);
nor U16317 (N_16317,N_16221,N_16243);
or U16318 (N_16318,N_16203,N_16095);
nor U16319 (N_16319,N_16207,N_16016);
nor U16320 (N_16320,N_16189,N_16177);
and U16321 (N_16321,N_16137,N_16102);
and U16322 (N_16322,N_16202,N_16199);
or U16323 (N_16323,N_16194,N_16041);
nor U16324 (N_16324,N_16187,N_16157);
nor U16325 (N_16325,N_16021,N_16198);
xor U16326 (N_16326,N_16073,N_16112);
nand U16327 (N_16327,N_16204,N_16122);
or U16328 (N_16328,N_16038,N_16223);
or U16329 (N_16329,N_16033,N_16087);
or U16330 (N_16330,N_16000,N_16200);
xnor U16331 (N_16331,N_16005,N_16147);
xor U16332 (N_16332,N_16182,N_16036);
nand U16333 (N_16333,N_16226,N_16150);
nor U16334 (N_16334,N_16208,N_16149);
and U16335 (N_16335,N_16169,N_16155);
and U16336 (N_16336,N_16186,N_16097);
nor U16337 (N_16337,N_16105,N_16011);
nor U16338 (N_16338,N_16083,N_16215);
and U16339 (N_16339,N_16193,N_16056);
xnor U16340 (N_16340,N_16089,N_16071);
nand U16341 (N_16341,N_16166,N_16082);
xnor U16342 (N_16342,N_16031,N_16094);
xor U16343 (N_16343,N_16017,N_16209);
and U16344 (N_16344,N_16144,N_16077);
nand U16345 (N_16345,N_16059,N_16115);
nand U16346 (N_16346,N_16172,N_16118);
or U16347 (N_16347,N_16185,N_16090);
or U16348 (N_16348,N_16100,N_16003);
or U16349 (N_16349,N_16091,N_16220);
or U16350 (N_16350,N_16058,N_16047);
nor U16351 (N_16351,N_16206,N_16001);
or U16352 (N_16352,N_16120,N_16030);
nor U16353 (N_16353,N_16074,N_16218);
and U16354 (N_16354,N_16032,N_16061);
nor U16355 (N_16355,N_16205,N_16214);
nand U16356 (N_16356,N_16093,N_16151);
or U16357 (N_16357,N_16023,N_16101);
nand U16358 (N_16358,N_16019,N_16235);
and U16359 (N_16359,N_16127,N_16158);
xor U16360 (N_16360,N_16247,N_16098);
and U16361 (N_16361,N_16068,N_16018);
and U16362 (N_16362,N_16145,N_16154);
and U16363 (N_16363,N_16197,N_16210);
or U16364 (N_16364,N_16180,N_16028);
or U16365 (N_16365,N_16212,N_16116);
or U16366 (N_16366,N_16181,N_16153);
or U16367 (N_16367,N_16233,N_16026);
nand U16368 (N_16368,N_16138,N_16156);
or U16369 (N_16369,N_16022,N_16211);
nor U16370 (N_16370,N_16236,N_16008);
xnor U16371 (N_16371,N_16128,N_16081);
nand U16372 (N_16372,N_16142,N_16136);
nor U16373 (N_16373,N_16167,N_16232);
xor U16374 (N_16374,N_16168,N_16126);
nor U16375 (N_16375,N_16142,N_16080);
and U16376 (N_16376,N_16225,N_16137);
or U16377 (N_16377,N_16008,N_16211);
and U16378 (N_16378,N_16120,N_16022);
or U16379 (N_16379,N_16142,N_16189);
nand U16380 (N_16380,N_16028,N_16027);
nand U16381 (N_16381,N_16162,N_16003);
xnor U16382 (N_16382,N_16113,N_16199);
nand U16383 (N_16383,N_16223,N_16118);
or U16384 (N_16384,N_16149,N_16186);
or U16385 (N_16385,N_16175,N_16011);
or U16386 (N_16386,N_16229,N_16073);
or U16387 (N_16387,N_16159,N_16059);
or U16388 (N_16388,N_16031,N_16167);
and U16389 (N_16389,N_16234,N_16210);
and U16390 (N_16390,N_16143,N_16112);
and U16391 (N_16391,N_16199,N_16163);
nor U16392 (N_16392,N_16106,N_16045);
xnor U16393 (N_16393,N_16095,N_16234);
nor U16394 (N_16394,N_16200,N_16025);
and U16395 (N_16395,N_16148,N_16070);
and U16396 (N_16396,N_16209,N_16203);
nor U16397 (N_16397,N_16068,N_16073);
nand U16398 (N_16398,N_16084,N_16148);
or U16399 (N_16399,N_16044,N_16215);
nand U16400 (N_16400,N_16011,N_16073);
or U16401 (N_16401,N_16096,N_16033);
xnor U16402 (N_16402,N_16184,N_16194);
and U16403 (N_16403,N_16031,N_16088);
or U16404 (N_16404,N_16180,N_16060);
nor U16405 (N_16405,N_16004,N_16240);
or U16406 (N_16406,N_16122,N_16091);
xor U16407 (N_16407,N_16125,N_16187);
nor U16408 (N_16408,N_16036,N_16108);
nor U16409 (N_16409,N_16194,N_16220);
nor U16410 (N_16410,N_16178,N_16079);
nor U16411 (N_16411,N_16231,N_16123);
or U16412 (N_16412,N_16120,N_16224);
nand U16413 (N_16413,N_16185,N_16026);
nand U16414 (N_16414,N_16227,N_16002);
xor U16415 (N_16415,N_16089,N_16081);
or U16416 (N_16416,N_16046,N_16216);
nor U16417 (N_16417,N_16225,N_16123);
nor U16418 (N_16418,N_16142,N_16168);
and U16419 (N_16419,N_16189,N_16092);
nand U16420 (N_16420,N_16144,N_16052);
or U16421 (N_16421,N_16109,N_16039);
and U16422 (N_16422,N_16004,N_16140);
nand U16423 (N_16423,N_16026,N_16191);
nor U16424 (N_16424,N_16219,N_16182);
or U16425 (N_16425,N_16197,N_16064);
nor U16426 (N_16426,N_16128,N_16103);
or U16427 (N_16427,N_16123,N_16019);
nand U16428 (N_16428,N_16011,N_16154);
or U16429 (N_16429,N_16066,N_16070);
and U16430 (N_16430,N_16056,N_16179);
xnor U16431 (N_16431,N_16173,N_16050);
nand U16432 (N_16432,N_16098,N_16207);
nor U16433 (N_16433,N_16211,N_16119);
xnor U16434 (N_16434,N_16169,N_16154);
xor U16435 (N_16435,N_16224,N_16093);
nand U16436 (N_16436,N_16247,N_16248);
xor U16437 (N_16437,N_16051,N_16059);
or U16438 (N_16438,N_16078,N_16076);
nor U16439 (N_16439,N_16083,N_16056);
and U16440 (N_16440,N_16172,N_16061);
and U16441 (N_16441,N_16230,N_16041);
nor U16442 (N_16442,N_16102,N_16029);
nor U16443 (N_16443,N_16004,N_16135);
nor U16444 (N_16444,N_16168,N_16178);
or U16445 (N_16445,N_16032,N_16002);
and U16446 (N_16446,N_16046,N_16109);
or U16447 (N_16447,N_16082,N_16188);
xnor U16448 (N_16448,N_16200,N_16238);
nand U16449 (N_16449,N_16243,N_16058);
and U16450 (N_16450,N_16089,N_16208);
and U16451 (N_16451,N_16035,N_16127);
xor U16452 (N_16452,N_16008,N_16240);
nand U16453 (N_16453,N_16123,N_16177);
nor U16454 (N_16454,N_16235,N_16236);
nand U16455 (N_16455,N_16083,N_16003);
and U16456 (N_16456,N_16167,N_16074);
and U16457 (N_16457,N_16030,N_16106);
nand U16458 (N_16458,N_16219,N_16174);
nand U16459 (N_16459,N_16222,N_16115);
or U16460 (N_16460,N_16137,N_16063);
nor U16461 (N_16461,N_16248,N_16015);
nor U16462 (N_16462,N_16147,N_16078);
xor U16463 (N_16463,N_16111,N_16185);
and U16464 (N_16464,N_16014,N_16064);
or U16465 (N_16465,N_16029,N_16025);
xnor U16466 (N_16466,N_16060,N_16174);
nand U16467 (N_16467,N_16236,N_16090);
and U16468 (N_16468,N_16163,N_16134);
or U16469 (N_16469,N_16009,N_16071);
or U16470 (N_16470,N_16003,N_16120);
nor U16471 (N_16471,N_16158,N_16124);
and U16472 (N_16472,N_16053,N_16179);
nand U16473 (N_16473,N_16080,N_16056);
nand U16474 (N_16474,N_16051,N_16054);
nor U16475 (N_16475,N_16008,N_16016);
and U16476 (N_16476,N_16156,N_16128);
nand U16477 (N_16477,N_16023,N_16022);
or U16478 (N_16478,N_16165,N_16071);
or U16479 (N_16479,N_16165,N_16135);
and U16480 (N_16480,N_16194,N_16191);
xor U16481 (N_16481,N_16229,N_16122);
nor U16482 (N_16482,N_16236,N_16147);
nor U16483 (N_16483,N_16096,N_16053);
or U16484 (N_16484,N_16169,N_16033);
or U16485 (N_16485,N_16182,N_16193);
or U16486 (N_16486,N_16040,N_16094);
and U16487 (N_16487,N_16114,N_16156);
xnor U16488 (N_16488,N_16037,N_16117);
nor U16489 (N_16489,N_16162,N_16048);
xor U16490 (N_16490,N_16234,N_16213);
xnor U16491 (N_16491,N_16229,N_16060);
or U16492 (N_16492,N_16073,N_16052);
and U16493 (N_16493,N_16220,N_16126);
xnor U16494 (N_16494,N_16132,N_16167);
xnor U16495 (N_16495,N_16099,N_16186);
xor U16496 (N_16496,N_16108,N_16210);
nor U16497 (N_16497,N_16075,N_16172);
and U16498 (N_16498,N_16009,N_16070);
xnor U16499 (N_16499,N_16062,N_16200);
and U16500 (N_16500,N_16295,N_16371);
or U16501 (N_16501,N_16459,N_16328);
xnor U16502 (N_16502,N_16279,N_16292);
and U16503 (N_16503,N_16323,N_16454);
or U16504 (N_16504,N_16327,N_16337);
and U16505 (N_16505,N_16362,N_16380);
nor U16506 (N_16506,N_16289,N_16453);
or U16507 (N_16507,N_16359,N_16265);
xnor U16508 (N_16508,N_16304,N_16351);
nand U16509 (N_16509,N_16298,N_16273);
and U16510 (N_16510,N_16314,N_16448);
or U16511 (N_16511,N_16449,N_16263);
or U16512 (N_16512,N_16412,N_16435);
xor U16513 (N_16513,N_16319,N_16375);
or U16514 (N_16514,N_16258,N_16305);
and U16515 (N_16515,N_16267,N_16348);
and U16516 (N_16516,N_16290,N_16256);
and U16517 (N_16517,N_16338,N_16408);
nor U16518 (N_16518,N_16301,N_16287);
nor U16519 (N_16519,N_16491,N_16352);
nor U16520 (N_16520,N_16481,N_16428);
xor U16521 (N_16521,N_16311,N_16344);
nand U16522 (N_16522,N_16366,N_16331);
nor U16523 (N_16523,N_16266,N_16442);
and U16524 (N_16524,N_16425,N_16487);
nand U16525 (N_16525,N_16409,N_16452);
nand U16526 (N_16526,N_16413,N_16250);
nor U16527 (N_16527,N_16414,N_16367);
and U16528 (N_16528,N_16294,N_16300);
nand U16529 (N_16529,N_16285,N_16252);
and U16530 (N_16530,N_16355,N_16395);
nor U16531 (N_16531,N_16335,N_16316);
xor U16532 (N_16532,N_16430,N_16418);
xor U16533 (N_16533,N_16334,N_16339);
nor U16534 (N_16534,N_16440,N_16485);
xor U16535 (N_16535,N_16282,N_16272);
nor U16536 (N_16536,N_16464,N_16261);
or U16537 (N_16537,N_16322,N_16492);
xor U16538 (N_16538,N_16404,N_16444);
xnor U16539 (N_16539,N_16499,N_16309);
and U16540 (N_16540,N_16475,N_16370);
nor U16541 (N_16541,N_16403,N_16391);
nor U16542 (N_16542,N_16460,N_16437);
xnor U16543 (N_16543,N_16284,N_16357);
xor U16544 (N_16544,N_16474,N_16293);
nor U16545 (N_16545,N_16317,N_16429);
nand U16546 (N_16546,N_16441,N_16354);
and U16547 (N_16547,N_16443,N_16382);
or U16548 (N_16548,N_16432,N_16490);
nand U16549 (N_16549,N_16251,N_16369);
nand U16550 (N_16550,N_16320,N_16324);
and U16551 (N_16551,N_16423,N_16488);
and U16552 (N_16552,N_16451,N_16426);
nand U16553 (N_16553,N_16381,N_16387);
nand U16554 (N_16554,N_16358,N_16471);
xnor U16555 (N_16555,N_16340,N_16278);
nand U16556 (N_16556,N_16307,N_16439);
nand U16557 (N_16557,N_16419,N_16281);
xor U16558 (N_16558,N_16496,N_16470);
or U16559 (N_16559,N_16483,N_16262);
nand U16560 (N_16560,N_16384,N_16345);
nand U16561 (N_16561,N_16462,N_16479);
nor U16562 (N_16562,N_16275,N_16390);
or U16563 (N_16563,N_16347,N_16325);
or U16564 (N_16564,N_16424,N_16446);
nand U16565 (N_16565,N_16363,N_16310);
nor U16566 (N_16566,N_16353,N_16349);
and U16567 (N_16567,N_16399,N_16473);
and U16568 (N_16568,N_16438,N_16383);
and U16569 (N_16569,N_16257,N_16450);
xor U16570 (N_16570,N_16379,N_16330);
nor U16571 (N_16571,N_16389,N_16260);
xnor U16572 (N_16572,N_16497,N_16478);
nand U16573 (N_16573,N_16388,N_16374);
xnor U16574 (N_16574,N_16299,N_16288);
nor U16575 (N_16575,N_16482,N_16477);
nor U16576 (N_16576,N_16361,N_16465);
nor U16577 (N_16577,N_16378,N_16297);
and U16578 (N_16578,N_16321,N_16494);
xor U16579 (N_16579,N_16360,N_16421);
and U16580 (N_16580,N_16469,N_16291);
xor U16581 (N_16581,N_16264,N_16329);
xnor U16582 (N_16582,N_16394,N_16364);
or U16583 (N_16583,N_16373,N_16255);
nor U16584 (N_16584,N_16466,N_16397);
and U16585 (N_16585,N_16445,N_16302);
or U16586 (N_16586,N_16436,N_16312);
or U16587 (N_16587,N_16377,N_16472);
nor U16588 (N_16588,N_16398,N_16461);
xor U16589 (N_16589,N_16303,N_16417);
xnor U16590 (N_16590,N_16427,N_16495);
nor U16591 (N_16591,N_16498,N_16393);
xor U16592 (N_16592,N_16332,N_16276);
and U16593 (N_16593,N_16480,N_16405);
or U16594 (N_16594,N_16326,N_16341);
nor U16595 (N_16595,N_16368,N_16271);
nor U16596 (N_16596,N_16420,N_16463);
nor U16597 (N_16597,N_16274,N_16277);
and U16598 (N_16598,N_16306,N_16458);
and U16599 (N_16599,N_16422,N_16333);
nor U16600 (N_16600,N_16392,N_16336);
nor U16601 (N_16601,N_16476,N_16385);
nand U16602 (N_16602,N_16407,N_16283);
nand U16603 (N_16603,N_16315,N_16433);
nor U16604 (N_16604,N_16286,N_16269);
or U16605 (N_16605,N_16318,N_16350);
and U16606 (N_16606,N_16467,N_16313);
and U16607 (N_16607,N_16484,N_16431);
and U16608 (N_16608,N_16259,N_16447);
xor U16609 (N_16609,N_16406,N_16254);
or U16610 (N_16610,N_16486,N_16386);
and U16611 (N_16611,N_16376,N_16308);
and U16612 (N_16612,N_16372,N_16457);
or U16613 (N_16613,N_16356,N_16402);
or U16614 (N_16614,N_16416,N_16456);
nor U16615 (N_16615,N_16415,N_16270);
nor U16616 (N_16616,N_16493,N_16396);
and U16617 (N_16617,N_16296,N_16346);
nor U16618 (N_16618,N_16434,N_16280);
nor U16619 (N_16619,N_16365,N_16489);
or U16620 (N_16620,N_16400,N_16342);
or U16621 (N_16621,N_16401,N_16455);
nand U16622 (N_16622,N_16343,N_16410);
nand U16623 (N_16623,N_16468,N_16268);
nand U16624 (N_16624,N_16253,N_16411);
nand U16625 (N_16625,N_16255,N_16479);
or U16626 (N_16626,N_16310,N_16480);
xnor U16627 (N_16627,N_16328,N_16389);
and U16628 (N_16628,N_16499,N_16453);
and U16629 (N_16629,N_16446,N_16279);
nor U16630 (N_16630,N_16331,N_16263);
xor U16631 (N_16631,N_16258,N_16449);
and U16632 (N_16632,N_16320,N_16281);
nand U16633 (N_16633,N_16253,N_16306);
and U16634 (N_16634,N_16335,N_16273);
or U16635 (N_16635,N_16380,N_16322);
nand U16636 (N_16636,N_16413,N_16496);
xnor U16637 (N_16637,N_16368,N_16360);
xnor U16638 (N_16638,N_16360,N_16338);
and U16639 (N_16639,N_16424,N_16395);
nor U16640 (N_16640,N_16477,N_16453);
xnor U16641 (N_16641,N_16384,N_16349);
nor U16642 (N_16642,N_16380,N_16347);
nor U16643 (N_16643,N_16389,N_16397);
nand U16644 (N_16644,N_16446,N_16390);
xnor U16645 (N_16645,N_16467,N_16402);
and U16646 (N_16646,N_16387,N_16339);
or U16647 (N_16647,N_16407,N_16346);
nor U16648 (N_16648,N_16335,N_16429);
nand U16649 (N_16649,N_16447,N_16296);
or U16650 (N_16650,N_16323,N_16460);
or U16651 (N_16651,N_16467,N_16338);
nand U16652 (N_16652,N_16374,N_16370);
nor U16653 (N_16653,N_16437,N_16349);
and U16654 (N_16654,N_16383,N_16490);
nand U16655 (N_16655,N_16499,N_16390);
and U16656 (N_16656,N_16315,N_16368);
and U16657 (N_16657,N_16388,N_16438);
or U16658 (N_16658,N_16372,N_16337);
nor U16659 (N_16659,N_16385,N_16350);
nand U16660 (N_16660,N_16399,N_16418);
xnor U16661 (N_16661,N_16329,N_16488);
or U16662 (N_16662,N_16268,N_16254);
nand U16663 (N_16663,N_16498,N_16403);
or U16664 (N_16664,N_16258,N_16374);
xnor U16665 (N_16665,N_16472,N_16411);
nand U16666 (N_16666,N_16350,N_16302);
or U16667 (N_16667,N_16354,N_16486);
nor U16668 (N_16668,N_16296,N_16487);
xor U16669 (N_16669,N_16284,N_16361);
or U16670 (N_16670,N_16368,N_16365);
nor U16671 (N_16671,N_16350,N_16401);
xor U16672 (N_16672,N_16297,N_16467);
nand U16673 (N_16673,N_16477,N_16495);
and U16674 (N_16674,N_16271,N_16319);
xor U16675 (N_16675,N_16494,N_16478);
xnor U16676 (N_16676,N_16406,N_16271);
nor U16677 (N_16677,N_16324,N_16351);
xor U16678 (N_16678,N_16314,N_16482);
nand U16679 (N_16679,N_16285,N_16454);
nor U16680 (N_16680,N_16255,N_16345);
nor U16681 (N_16681,N_16459,N_16400);
xnor U16682 (N_16682,N_16321,N_16352);
and U16683 (N_16683,N_16394,N_16485);
nor U16684 (N_16684,N_16452,N_16419);
or U16685 (N_16685,N_16298,N_16454);
nor U16686 (N_16686,N_16268,N_16419);
and U16687 (N_16687,N_16349,N_16464);
or U16688 (N_16688,N_16417,N_16424);
nor U16689 (N_16689,N_16262,N_16368);
xnor U16690 (N_16690,N_16309,N_16365);
nand U16691 (N_16691,N_16466,N_16386);
and U16692 (N_16692,N_16307,N_16430);
nor U16693 (N_16693,N_16337,N_16427);
nand U16694 (N_16694,N_16469,N_16389);
nor U16695 (N_16695,N_16443,N_16427);
nand U16696 (N_16696,N_16360,N_16450);
xor U16697 (N_16697,N_16398,N_16303);
nand U16698 (N_16698,N_16364,N_16379);
and U16699 (N_16699,N_16406,N_16389);
and U16700 (N_16700,N_16303,N_16456);
nand U16701 (N_16701,N_16471,N_16349);
or U16702 (N_16702,N_16398,N_16496);
and U16703 (N_16703,N_16490,N_16341);
or U16704 (N_16704,N_16455,N_16421);
or U16705 (N_16705,N_16404,N_16496);
xnor U16706 (N_16706,N_16375,N_16376);
xor U16707 (N_16707,N_16363,N_16324);
or U16708 (N_16708,N_16256,N_16364);
nor U16709 (N_16709,N_16336,N_16285);
xnor U16710 (N_16710,N_16288,N_16399);
or U16711 (N_16711,N_16408,N_16295);
nor U16712 (N_16712,N_16335,N_16361);
xnor U16713 (N_16713,N_16364,N_16278);
nand U16714 (N_16714,N_16439,N_16278);
and U16715 (N_16715,N_16450,N_16464);
nand U16716 (N_16716,N_16402,N_16406);
or U16717 (N_16717,N_16276,N_16273);
or U16718 (N_16718,N_16266,N_16267);
and U16719 (N_16719,N_16496,N_16377);
or U16720 (N_16720,N_16296,N_16492);
xnor U16721 (N_16721,N_16435,N_16332);
xor U16722 (N_16722,N_16307,N_16272);
nand U16723 (N_16723,N_16310,N_16302);
nand U16724 (N_16724,N_16390,N_16265);
and U16725 (N_16725,N_16372,N_16262);
xor U16726 (N_16726,N_16430,N_16349);
nor U16727 (N_16727,N_16270,N_16269);
xnor U16728 (N_16728,N_16478,N_16457);
xor U16729 (N_16729,N_16476,N_16460);
nor U16730 (N_16730,N_16477,N_16372);
nand U16731 (N_16731,N_16252,N_16454);
and U16732 (N_16732,N_16495,N_16364);
nor U16733 (N_16733,N_16446,N_16286);
nand U16734 (N_16734,N_16277,N_16361);
or U16735 (N_16735,N_16342,N_16262);
or U16736 (N_16736,N_16457,N_16279);
nand U16737 (N_16737,N_16338,N_16466);
or U16738 (N_16738,N_16450,N_16274);
and U16739 (N_16739,N_16382,N_16339);
and U16740 (N_16740,N_16482,N_16278);
or U16741 (N_16741,N_16333,N_16445);
or U16742 (N_16742,N_16271,N_16349);
and U16743 (N_16743,N_16390,N_16430);
or U16744 (N_16744,N_16384,N_16324);
and U16745 (N_16745,N_16498,N_16307);
and U16746 (N_16746,N_16388,N_16272);
nor U16747 (N_16747,N_16368,N_16354);
nand U16748 (N_16748,N_16393,N_16386);
nand U16749 (N_16749,N_16306,N_16385);
and U16750 (N_16750,N_16512,N_16663);
and U16751 (N_16751,N_16684,N_16651);
nand U16752 (N_16752,N_16520,N_16664);
xnor U16753 (N_16753,N_16602,N_16588);
or U16754 (N_16754,N_16667,N_16540);
nor U16755 (N_16755,N_16678,N_16586);
nor U16756 (N_16756,N_16747,N_16621);
nor U16757 (N_16757,N_16691,N_16608);
nand U16758 (N_16758,N_16617,N_16701);
and U16759 (N_16759,N_16703,N_16513);
nor U16760 (N_16760,N_16646,N_16706);
and U16761 (N_16761,N_16696,N_16639);
and U16762 (N_16762,N_16628,N_16541);
nor U16763 (N_16763,N_16626,N_16681);
nor U16764 (N_16764,N_16594,N_16519);
or U16765 (N_16765,N_16606,N_16685);
or U16766 (N_16766,N_16702,N_16654);
xor U16767 (N_16767,N_16642,N_16549);
nor U16768 (N_16768,N_16670,N_16571);
nand U16769 (N_16769,N_16563,N_16614);
or U16770 (N_16770,N_16680,N_16649);
or U16771 (N_16771,N_16682,N_16632);
nor U16772 (N_16772,N_16659,N_16592);
or U16773 (N_16773,N_16698,N_16660);
or U16774 (N_16774,N_16542,N_16507);
nand U16775 (N_16775,N_16741,N_16600);
nor U16776 (N_16776,N_16593,N_16689);
nor U16777 (N_16777,N_16648,N_16645);
nor U16778 (N_16778,N_16577,N_16722);
or U16779 (N_16779,N_16616,N_16688);
xor U16780 (N_16780,N_16572,N_16609);
nand U16781 (N_16781,N_16510,N_16625);
nand U16782 (N_16782,N_16717,N_16587);
and U16783 (N_16783,N_16535,N_16575);
xor U16784 (N_16784,N_16735,N_16567);
nand U16785 (N_16785,N_16611,N_16673);
xnor U16786 (N_16786,N_16695,N_16693);
nor U16787 (N_16787,N_16668,N_16718);
nor U16788 (N_16788,N_16509,N_16697);
or U16789 (N_16789,N_16550,N_16662);
nand U16790 (N_16790,N_16551,N_16748);
nand U16791 (N_16791,N_16506,N_16511);
xor U16792 (N_16792,N_16623,N_16525);
and U16793 (N_16793,N_16730,N_16729);
or U16794 (N_16794,N_16707,N_16554);
xnor U16795 (N_16795,N_16643,N_16523);
nand U16796 (N_16796,N_16584,N_16672);
or U16797 (N_16797,N_16676,N_16711);
and U16798 (N_16798,N_16537,N_16508);
nor U16799 (N_16799,N_16545,N_16737);
xor U16800 (N_16800,N_16533,N_16502);
or U16801 (N_16801,N_16522,N_16599);
and U16802 (N_16802,N_16634,N_16650);
and U16803 (N_16803,N_16530,N_16612);
or U16804 (N_16804,N_16607,N_16704);
nand U16805 (N_16805,N_16553,N_16647);
xnor U16806 (N_16806,N_16579,N_16504);
xnor U16807 (N_16807,N_16618,N_16574);
and U16808 (N_16808,N_16610,N_16582);
nand U16809 (N_16809,N_16573,N_16539);
nor U16810 (N_16810,N_16543,N_16677);
or U16811 (N_16811,N_16590,N_16566);
or U16812 (N_16812,N_16658,N_16595);
nand U16813 (N_16813,N_16605,N_16708);
or U16814 (N_16814,N_16633,N_16749);
and U16815 (N_16815,N_16679,N_16524);
xnor U16816 (N_16816,N_16629,N_16630);
and U16817 (N_16817,N_16552,N_16720);
and U16818 (N_16818,N_16734,N_16565);
nand U16819 (N_16819,N_16714,N_16666);
xnor U16820 (N_16820,N_16675,N_16687);
and U16821 (N_16821,N_16517,N_16740);
and U16822 (N_16822,N_16743,N_16656);
and U16823 (N_16823,N_16596,N_16576);
xnor U16824 (N_16824,N_16555,N_16744);
or U16825 (N_16825,N_16518,N_16674);
or U16826 (N_16826,N_16503,N_16739);
and U16827 (N_16827,N_16700,N_16627);
and U16828 (N_16828,N_16640,N_16526);
xor U16829 (N_16829,N_16655,N_16613);
or U16830 (N_16830,N_16683,N_16603);
and U16831 (N_16831,N_16742,N_16516);
xor U16832 (N_16832,N_16569,N_16726);
xor U16833 (N_16833,N_16637,N_16538);
and U16834 (N_16834,N_16638,N_16652);
and U16835 (N_16835,N_16557,N_16568);
nand U16836 (N_16836,N_16745,N_16501);
and U16837 (N_16837,N_16591,N_16721);
nor U16838 (N_16838,N_16694,N_16527);
nor U16839 (N_16839,N_16598,N_16686);
nor U16840 (N_16840,N_16728,N_16635);
nor U16841 (N_16841,N_16746,N_16665);
and U16842 (N_16842,N_16715,N_16716);
xnor U16843 (N_16843,N_16532,N_16514);
nor U16844 (N_16844,N_16705,N_16589);
xnor U16845 (N_16845,N_16657,N_16731);
and U16846 (N_16846,N_16531,N_16581);
and U16847 (N_16847,N_16601,N_16723);
and U16848 (N_16848,N_16536,N_16641);
xnor U16849 (N_16849,N_16521,N_16727);
and U16850 (N_16850,N_16544,N_16597);
or U16851 (N_16851,N_16546,N_16580);
nor U16852 (N_16852,N_16725,N_16515);
or U16853 (N_16853,N_16548,N_16604);
nand U16854 (N_16854,N_16500,N_16570);
and U16855 (N_16855,N_16619,N_16560);
or U16856 (N_16856,N_16615,N_16556);
or U16857 (N_16857,N_16561,N_16699);
nand U16858 (N_16858,N_16505,N_16692);
and U16859 (N_16859,N_16644,N_16559);
or U16860 (N_16860,N_16733,N_16661);
and U16861 (N_16861,N_16738,N_16558);
or U16862 (N_16862,N_16732,N_16622);
xor U16863 (N_16863,N_16631,N_16534);
xnor U16864 (N_16864,N_16585,N_16736);
and U16865 (N_16865,N_16620,N_16528);
or U16866 (N_16866,N_16624,N_16578);
nand U16867 (N_16867,N_16724,N_16713);
nand U16868 (N_16868,N_16690,N_16547);
nor U16869 (N_16869,N_16529,N_16719);
and U16870 (N_16870,N_16669,N_16562);
or U16871 (N_16871,N_16710,N_16564);
and U16872 (N_16872,N_16583,N_16671);
nor U16873 (N_16873,N_16709,N_16712);
and U16874 (N_16874,N_16653,N_16636);
nor U16875 (N_16875,N_16589,N_16603);
nand U16876 (N_16876,N_16703,N_16672);
and U16877 (N_16877,N_16739,N_16745);
xnor U16878 (N_16878,N_16647,N_16511);
nor U16879 (N_16879,N_16747,N_16556);
or U16880 (N_16880,N_16507,N_16613);
and U16881 (N_16881,N_16668,N_16503);
nand U16882 (N_16882,N_16529,N_16601);
xor U16883 (N_16883,N_16626,N_16610);
nor U16884 (N_16884,N_16502,N_16654);
and U16885 (N_16885,N_16721,N_16511);
nand U16886 (N_16886,N_16514,N_16559);
or U16887 (N_16887,N_16682,N_16559);
nor U16888 (N_16888,N_16554,N_16696);
and U16889 (N_16889,N_16557,N_16506);
xnor U16890 (N_16890,N_16680,N_16628);
nand U16891 (N_16891,N_16502,N_16721);
xnor U16892 (N_16892,N_16659,N_16685);
nand U16893 (N_16893,N_16702,N_16680);
xor U16894 (N_16894,N_16611,N_16614);
nand U16895 (N_16895,N_16518,N_16662);
or U16896 (N_16896,N_16685,N_16716);
nor U16897 (N_16897,N_16695,N_16681);
nor U16898 (N_16898,N_16612,N_16515);
nand U16899 (N_16899,N_16683,N_16562);
or U16900 (N_16900,N_16720,N_16624);
xnor U16901 (N_16901,N_16552,N_16639);
and U16902 (N_16902,N_16649,N_16582);
or U16903 (N_16903,N_16688,N_16538);
nand U16904 (N_16904,N_16709,N_16744);
nand U16905 (N_16905,N_16663,N_16598);
nand U16906 (N_16906,N_16534,N_16739);
nand U16907 (N_16907,N_16712,N_16522);
xnor U16908 (N_16908,N_16546,N_16665);
and U16909 (N_16909,N_16609,N_16671);
nor U16910 (N_16910,N_16573,N_16626);
and U16911 (N_16911,N_16574,N_16602);
nand U16912 (N_16912,N_16705,N_16621);
or U16913 (N_16913,N_16642,N_16612);
nand U16914 (N_16914,N_16689,N_16702);
or U16915 (N_16915,N_16644,N_16743);
nand U16916 (N_16916,N_16615,N_16568);
nand U16917 (N_16917,N_16642,N_16728);
nand U16918 (N_16918,N_16633,N_16650);
xnor U16919 (N_16919,N_16692,N_16722);
or U16920 (N_16920,N_16691,N_16643);
xnor U16921 (N_16921,N_16720,N_16701);
nor U16922 (N_16922,N_16734,N_16710);
xnor U16923 (N_16923,N_16663,N_16716);
xor U16924 (N_16924,N_16724,N_16574);
or U16925 (N_16925,N_16540,N_16537);
and U16926 (N_16926,N_16659,N_16615);
xor U16927 (N_16927,N_16741,N_16699);
xnor U16928 (N_16928,N_16524,N_16584);
or U16929 (N_16929,N_16508,N_16674);
nand U16930 (N_16930,N_16721,N_16644);
nor U16931 (N_16931,N_16660,N_16566);
xnor U16932 (N_16932,N_16685,N_16736);
or U16933 (N_16933,N_16505,N_16729);
nor U16934 (N_16934,N_16626,N_16713);
or U16935 (N_16935,N_16672,N_16679);
or U16936 (N_16936,N_16694,N_16741);
or U16937 (N_16937,N_16622,N_16734);
and U16938 (N_16938,N_16609,N_16541);
or U16939 (N_16939,N_16702,N_16727);
or U16940 (N_16940,N_16605,N_16607);
xnor U16941 (N_16941,N_16631,N_16661);
or U16942 (N_16942,N_16556,N_16614);
and U16943 (N_16943,N_16737,N_16621);
xor U16944 (N_16944,N_16736,N_16510);
nor U16945 (N_16945,N_16539,N_16502);
nor U16946 (N_16946,N_16743,N_16548);
nor U16947 (N_16947,N_16502,N_16680);
or U16948 (N_16948,N_16718,N_16582);
or U16949 (N_16949,N_16687,N_16678);
and U16950 (N_16950,N_16560,N_16583);
xnor U16951 (N_16951,N_16671,N_16703);
nand U16952 (N_16952,N_16540,N_16733);
xnor U16953 (N_16953,N_16584,N_16530);
and U16954 (N_16954,N_16561,N_16544);
and U16955 (N_16955,N_16720,N_16722);
or U16956 (N_16956,N_16539,N_16734);
nand U16957 (N_16957,N_16678,N_16680);
nand U16958 (N_16958,N_16553,N_16528);
xor U16959 (N_16959,N_16740,N_16531);
xnor U16960 (N_16960,N_16634,N_16555);
nor U16961 (N_16961,N_16693,N_16666);
and U16962 (N_16962,N_16702,N_16543);
nor U16963 (N_16963,N_16577,N_16708);
nor U16964 (N_16964,N_16661,N_16576);
nor U16965 (N_16965,N_16677,N_16735);
and U16966 (N_16966,N_16593,N_16737);
xnor U16967 (N_16967,N_16678,N_16536);
nand U16968 (N_16968,N_16505,N_16623);
xor U16969 (N_16969,N_16559,N_16527);
nand U16970 (N_16970,N_16687,N_16697);
and U16971 (N_16971,N_16521,N_16572);
or U16972 (N_16972,N_16717,N_16644);
or U16973 (N_16973,N_16507,N_16501);
nor U16974 (N_16974,N_16677,N_16505);
nor U16975 (N_16975,N_16739,N_16545);
nor U16976 (N_16976,N_16683,N_16698);
nand U16977 (N_16977,N_16660,N_16646);
and U16978 (N_16978,N_16628,N_16694);
xor U16979 (N_16979,N_16579,N_16711);
xnor U16980 (N_16980,N_16559,N_16658);
or U16981 (N_16981,N_16525,N_16546);
nand U16982 (N_16982,N_16693,N_16544);
nand U16983 (N_16983,N_16693,N_16529);
nand U16984 (N_16984,N_16692,N_16550);
nand U16985 (N_16985,N_16600,N_16724);
or U16986 (N_16986,N_16749,N_16631);
nor U16987 (N_16987,N_16725,N_16719);
or U16988 (N_16988,N_16698,N_16522);
and U16989 (N_16989,N_16571,N_16593);
xnor U16990 (N_16990,N_16739,N_16612);
nor U16991 (N_16991,N_16662,N_16515);
and U16992 (N_16992,N_16641,N_16690);
nand U16993 (N_16993,N_16560,N_16702);
xor U16994 (N_16994,N_16668,N_16523);
and U16995 (N_16995,N_16623,N_16569);
xnor U16996 (N_16996,N_16658,N_16667);
and U16997 (N_16997,N_16736,N_16711);
nor U16998 (N_16998,N_16704,N_16640);
nand U16999 (N_16999,N_16730,N_16599);
nand U17000 (N_17000,N_16846,N_16837);
and U17001 (N_17001,N_16826,N_16941);
xor U17002 (N_17002,N_16871,N_16834);
nand U17003 (N_17003,N_16879,N_16791);
and U17004 (N_17004,N_16776,N_16841);
or U17005 (N_17005,N_16833,N_16793);
nand U17006 (N_17006,N_16866,N_16929);
or U17007 (N_17007,N_16764,N_16940);
or U17008 (N_17008,N_16818,N_16986);
nor U17009 (N_17009,N_16870,N_16919);
nor U17010 (N_17010,N_16874,N_16798);
or U17011 (N_17011,N_16817,N_16908);
and U17012 (N_17012,N_16880,N_16800);
nand U17013 (N_17013,N_16858,N_16899);
xnor U17014 (N_17014,N_16981,N_16993);
and U17015 (N_17015,N_16814,N_16850);
or U17016 (N_17016,N_16890,N_16877);
or U17017 (N_17017,N_16997,N_16988);
and U17018 (N_17018,N_16914,N_16774);
nor U17019 (N_17019,N_16762,N_16773);
or U17020 (N_17020,N_16944,N_16783);
xnor U17021 (N_17021,N_16958,N_16822);
and U17022 (N_17022,N_16859,N_16875);
and U17023 (N_17023,N_16838,N_16987);
or U17024 (N_17024,N_16765,N_16831);
nand U17025 (N_17025,N_16878,N_16845);
or U17026 (N_17026,N_16970,N_16991);
xnor U17027 (N_17027,N_16998,N_16785);
xor U17028 (N_17028,N_16889,N_16853);
xor U17029 (N_17029,N_16828,N_16759);
nor U17030 (N_17030,N_16862,N_16855);
or U17031 (N_17031,N_16844,N_16868);
xnor U17032 (N_17032,N_16939,N_16901);
or U17033 (N_17033,N_16849,N_16771);
and U17034 (N_17034,N_16961,N_16936);
nand U17035 (N_17035,N_16933,N_16790);
and U17036 (N_17036,N_16915,N_16983);
or U17037 (N_17037,N_16969,N_16968);
nand U17038 (N_17038,N_16792,N_16851);
xnor U17039 (N_17039,N_16956,N_16891);
nor U17040 (N_17040,N_16984,N_16947);
nor U17041 (N_17041,N_16832,N_16766);
nor U17042 (N_17042,N_16836,N_16777);
and U17043 (N_17043,N_16772,N_16852);
xnor U17044 (N_17044,N_16913,N_16861);
nor U17045 (N_17045,N_16918,N_16819);
or U17046 (N_17046,N_16967,N_16995);
nand U17047 (N_17047,N_16917,N_16886);
and U17048 (N_17048,N_16842,N_16750);
nand U17049 (N_17049,N_16989,N_16896);
nor U17050 (N_17050,N_16928,N_16761);
and U17051 (N_17051,N_16910,N_16811);
and U17052 (N_17052,N_16807,N_16904);
nor U17053 (N_17053,N_16885,N_16932);
and U17054 (N_17054,N_16872,N_16769);
or U17055 (N_17055,N_16847,N_16787);
nor U17056 (N_17056,N_16797,N_16802);
or U17057 (N_17057,N_16952,N_16892);
or U17058 (N_17058,N_16955,N_16843);
and U17059 (N_17059,N_16945,N_16900);
xor U17060 (N_17060,N_16840,N_16805);
or U17061 (N_17061,N_16977,N_16821);
xnor U17062 (N_17062,N_16960,N_16951);
or U17063 (N_17063,N_16954,N_16796);
xnor U17064 (N_17064,N_16775,N_16902);
nand U17065 (N_17065,N_16810,N_16789);
nand U17066 (N_17066,N_16905,N_16972);
and U17067 (N_17067,N_16751,N_16781);
xnor U17068 (N_17068,N_16931,N_16959);
or U17069 (N_17069,N_16808,N_16942);
or U17070 (N_17070,N_16760,N_16803);
xnor U17071 (N_17071,N_16927,N_16780);
nand U17072 (N_17072,N_16985,N_16881);
and U17073 (N_17073,N_16921,N_16888);
xor U17074 (N_17074,N_16926,N_16903);
or U17075 (N_17075,N_16950,N_16949);
and U17076 (N_17076,N_16812,N_16999);
nand U17077 (N_17077,N_16895,N_16820);
xor U17078 (N_17078,N_16825,N_16883);
and U17079 (N_17079,N_16971,N_16909);
nand U17080 (N_17080,N_16975,N_16946);
nor U17081 (N_17081,N_16973,N_16911);
nor U17082 (N_17082,N_16799,N_16887);
nand U17083 (N_17083,N_16894,N_16824);
nor U17084 (N_17084,N_16938,N_16835);
xnor U17085 (N_17085,N_16925,N_16864);
and U17086 (N_17086,N_16912,N_16809);
or U17087 (N_17087,N_16964,N_16907);
xnor U17088 (N_17088,N_16794,N_16865);
nand U17089 (N_17089,N_16965,N_16979);
xnor U17090 (N_17090,N_16992,N_16830);
nor U17091 (N_17091,N_16990,N_16996);
or U17092 (N_17092,N_16943,N_16924);
and U17093 (N_17093,N_16854,N_16898);
xor U17094 (N_17094,N_16884,N_16906);
nor U17095 (N_17095,N_16974,N_16758);
xnor U17096 (N_17096,N_16863,N_16829);
or U17097 (N_17097,N_16882,N_16756);
nand U17098 (N_17098,N_16860,N_16753);
and U17099 (N_17099,N_16839,N_16763);
nor U17100 (N_17100,N_16966,N_16920);
nand U17101 (N_17101,N_16897,N_16869);
nand U17102 (N_17102,N_16982,N_16876);
or U17103 (N_17103,N_16916,N_16784);
or U17104 (N_17104,N_16978,N_16893);
or U17105 (N_17105,N_16930,N_16957);
xnor U17106 (N_17106,N_16948,N_16976);
xnor U17107 (N_17107,N_16922,N_16757);
nor U17108 (N_17108,N_16754,N_16923);
nor U17109 (N_17109,N_16788,N_16804);
or U17110 (N_17110,N_16801,N_16782);
or U17111 (N_17111,N_16963,N_16755);
or U17112 (N_17112,N_16962,N_16779);
nor U17113 (N_17113,N_16934,N_16770);
nand U17114 (N_17114,N_16823,N_16786);
and U17115 (N_17115,N_16856,N_16857);
or U17116 (N_17116,N_16848,N_16980);
xnor U17117 (N_17117,N_16752,N_16953);
nor U17118 (N_17118,N_16867,N_16937);
nor U17119 (N_17119,N_16827,N_16816);
xor U17120 (N_17120,N_16994,N_16815);
nand U17121 (N_17121,N_16935,N_16795);
and U17122 (N_17122,N_16813,N_16806);
and U17123 (N_17123,N_16873,N_16768);
nor U17124 (N_17124,N_16767,N_16778);
nor U17125 (N_17125,N_16962,N_16766);
or U17126 (N_17126,N_16999,N_16955);
xor U17127 (N_17127,N_16811,N_16890);
nand U17128 (N_17128,N_16911,N_16895);
and U17129 (N_17129,N_16775,N_16981);
xor U17130 (N_17130,N_16831,N_16753);
or U17131 (N_17131,N_16758,N_16786);
nor U17132 (N_17132,N_16903,N_16847);
nor U17133 (N_17133,N_16975,N_16838);
and U17134 (N_17134,N_16862,N_16841);
nor U17135 (N_17135,N_16997,N_16794);
or U17136 (N_17136,N_16898,N_16831);
nand U17137 (N_17137,N_16831,N_16933);
nor U17138 (N_17138,N_16969,N_16951);
nor U17139 (N_17139,N_16930,N_16798);
xnor U17140 (N_17140,N_16786,N_16773);
or U17141 (N_17141,N_16822,N_16769);
xor U17142 (N_17142,N_16945,N_16921);
and U17143 (N_17143,N_16799,N_16929);
or U17144 (N_17144,N_16848,N_16784);
or U17145 (N_17145,N_16915,N_16871);
and U17146 (N_17146,N_16960,N_16979);
xnor U17147 (N_17147,N_16868,N_16921);
and U17148 (N_17148,N_16953,N_16884);
and U17149 (N_17149,N_16887,N_16861);
xnor U17150 (N_17150,N_16928,N_16807);
nand U17151 (N_17151,N_16931,N_16869);
xor U17152 (N_17152,N_16765,N_16778);
or U17153 (N_17153,N_16759,N_16867);
nor U17154 (N_17154,N_16832,N_16859);
or U17155 (N_17155,N_16947,N_16915);
nand U17156 (N_17156,N_16776,N_16928);
and U17157 (N_17157,N_16823,N_16942);
xor U17158 (N_17158,N_16951,N_16769);
xnor U17159 (N_17159,N_16948,N_16768);
nand U17160 (N_17160,N_16865,N_16842);
and U17161 (N_17161,N_16942,N_16849);
nand U17162 (N_17162,N_16920,N_16852);
and U17163 (N_17163,N_16921,N_16899);
and U17164 (N_17164,N_16871,N_16751);
or U17165 (N_17165,N_16970,N_16765);
and U17166 (N_17166,N_16902,N_16970);
or U17167 (N_17167,N_16789,N_16936);
or U17168 (N_17168,N_16994,N_16759);
nand U17169 (N_17169,N_16893,N_16835);
nor U17170 (N_17170,N_16894,N_16891);
and U17171 (N_17171,N_16754,N_16768);
nand U17172 (N_17172,N_16830,N_16831);
nand U17173 (N_17173,N_16773,N_16805);
nor U17174 (N_17174,N_16892,N_16978);
or U17175 (N_17175,N_16898,N_16786);
xor U17176 (N_17176,N_16920,N_16786);
xor U17177 (N_17177,N_16967,N_16918);
nand U17178 (N_17178,N_16851,N_16935);
or U17179 (N_17179,N_16842,N_16915);
and U17180 (N_17180,N_16901,N_16836);
nor U17181 (N_17181,N_16953,N_16839);
or U17182 (N_17182,N_16881,N_16942);
nand U17183 (N_17183,N_16870,N_16814);
nor U17184 (N_17184,N_16873,N_16851);
nor U17185 (N_17185,N_16890,N_16990);
nand U17186 (N_17186,N_16861,N_16855);
nand U17187 (N_17187,N_16762,N_16897);
nand U17188 (N_17188,N_16811,N_16961);
nor U17189 (N_17189,N_16913,N_16981);
nand U17190 (N_17190,N_16841,N_16780);
or U17191 (N_17191,N_16945,N_16782);
or U17192 (N_17192,N_16925,N_16799);
or U17193 (N_17193,N_16930,N_16979);
xor U17194 (N_17194,N_16999,N_16818);
nand U17195 (N_17195,N_16854,N_16762);
or U17196 (N_17196,N_16819,N_16839);
or U17197 (N_17197,N_16780,N_16831);
and U17198 (N_17198,N_16839,N_16790);
nand U17199 (N_17199,N_16871,N_16855);
nor U17200 (N_17200,N_16920,N_16925);
nand U17201 (N_17201,N_16782,N_16933);
or U17202 (N_17202,N_16991,N_16760);
or U17203 (N_17203,N_16988,N_16755);
or U17204 (N_17204,N_16979,N_16899);
and U17205 (N_17205,N_16869,N_16998);
nor U17206 (N_17206,N_16763,N_16938);
nor U17207 (N_17207,N_16977,N_16970);
or U17208 (N_17208,N_16820,N_16954);
xnor U17209 (N_17209,N_16937,N_16859);
or U17210 (N_17210,N_16784,N_16940);
or U17211 (N_17211,N_16915,N_16887);
or U17212 (N_17212,N_16983,N_16755);
nand U17213 (N_17213,N_16768,N_16856);
xnor U17214 (N_17214,N_16980,N_16841);
xnor U17215 (N_17215,N_16973,N_16763);
nand U17216 (N_17216,N_16759,N_16943);
nand U17217 (N_17217,N_16970,N_16855);
or U17218 (N_17218,N_16838,N_16856);
or U17219 (N_17219,N_16996,N_16781);
nand U17220 (N_17220,N_16907,N_16916);
nor U17221 (N_17221,N_16775,N_16808);
and U17222 (N_17222,N_16812,N_16774);
or U17223 (N_17223,N_16885,N_16874);
nor U17224 (N_17224,N_16883,N_16774);
nor U17225 (N_17225,N_16959,N_16842);
nand U17226 (N_17226,N_16941,N_16897);
xnor U17227 (N_17227,N_16924,N_16977);
or U17228 (N_17228,N_16958,N_16865);
or U17229 (N_17229,N_16878,N_16789);
or U17230 (N_17230,N_16835,N_16929);
nand U17231 (N_17231,N_16750,N_16851);
nor U17232 (N_17232,N_16906,N_16898);
nor U17233 (N_17233,N_16979,N_16832);
xor U17234 (N_17234,N_16897,N_16999);
or U17235 (N_17235,N_16949,N_16955);
xor U17236 (N_17236,N_16771,N_16833);
nor U17237 (N_17237,N_16781,N_16864);
nand U17238 (N_17238,N_16930,N_16843);
nor U17239 (N_17239,N_16901,N_16769);
nor U17240 (N_17240,N_16806,N_16890);
nand U17241 (N_17241,N_16875,N_16987);
and U17242 (N_17242,N_16921,N_16763);
nor U17243 (N_17243,N_16908,N_16971);
nand U17244 (N_17244,N_16802,N_16822);
nand U17245 (N_17245,N_16751,N_16837);
nand U17246 (N_17246,N_16949,N_16893);
nand U17247 (N_17247,N_16776,N_16969);
nand U17248 (N_17248,N_16764,N_16790);
nor U17249 (N_17249,N_16955,N_16995);
or U17250 (N_17250,N_17056,N_17144);
nor U17251 (N_17251,N_17117,N_17195);
xor U17252 (N_17252,N_17223,N_17220);
xnor U17253 (N_17253,N_17017,N_17080);
nand U17254 (N_17254,N_17177,N_17108);
nand U17255 (N_17255,N_17134,N_17218);
nand U17256 (N_17256,N_17210,N_17213);
xor U17257 (N_17257,N_17243,N_17189);
xnor U17258 (N_17258,N_17046,N_17191);
xnor U17259 (N_17259,N_17086,N_17076);
nor U17260 (N_17260,N_17212,N_17111);
and U17261 (N_17261,N_17156,N_17161);
nand U17262 (N_17262,N_17003,N_17152);
nand U17263 (N_17263,N_17138,N_17235);
nand U17264 (N_17264,N_17198,N_17035);
and U17265 (N_17265,N_17181,N_17123);
and U17266 (N_17266,N_17158,N_17162);
and U17267 (N_17267,N_17019,N_17216);
or U17268 (N_17268,N_17055,N_17145);
or U17269 (N_17269,N_17098,N_17120);
nand U17270 (N_17270,N_17060,N_17050);
nor U17271 (N_17271,N_17022,N_17024);
nand U17272 (N_17272,N_17069,N_17178);
or U17273 (N_17273,N_17209,N_17027);
or U17274 (N_17274,N_17190,N_17155);
and U17275 (N_17275,N_17105,N_17200);
or U17276 (N_17276,N_17079,N_17197);
nand U17277 (N_17277,N_17228,N_17031);
nand U17278 (N_17278,N_17103,N_17176);
nor U17279 (N_17279,N_17225,N_17171);
xor U17280 (N_17280,N_17107,N_17160);
xnor U17281 (N_17281,N_17001,N_17217);
xor U17282 (N_17282,N_17203,N_17233);
xnor U17283 (N_17283,N_17124,N_17088);
xor U17284 (N_17284,N_17241,N_17081);
nand U17285 (N_17285,N_17201,N_17073);
or U17286 (N_17286,N_17102,N_17044);
and U17287 (N_17287,N_17175,N_17137);
or U17288 (N_17288,N_17094,N_17059);
nor U17289 (N_17289,N_17174,N_17106);
nand U17290 (N_17290,N_17010,N_17042);
and U17291 (N_17291,N_17149,N_17136);
nand U17292 (N_17292,N_17018,N_17034);
nor U17293 (N_17293,N_17096,N_17015);
and U17294 (N_17294,N_17192,N_17062);
or U17295 (N_17295,N_17025,N_17185);
nor U17296 (N_17296,N_17089,N_17066);
and U17297 (N_17297,N_17002,N_17140);
or U17298 (N_17298,N_17011,N_17004);
nor U17299 (N_17299,N_17077,N_17008);
nand U17300 (N_17300,N_17068,N_17125);
xnor U17301 (N_17301,N_17016,N_17199);
and U17302 (N_17302,N_17238,N_17232);
xor U17303 (N_17303,N_17187,N_17093);
nor U17304 (N_17304,N_17084,N_17104);
nor U17305 (N_17305,N_17070,N_17115);
or U17306 (N_17306,N_17173,N_17170);
and U17307 (N_17307,N_17071,N_17041);
nand U17308 (N_17308,N_17242,N_17006);
or U17309 (N_17309,N_17072,N_17133);
nand U17310 (N_17310,N_17040,N_17248);
or U17311 (N_17311,N_17023,N_17013);
or U17312 (N_17312,N_17039,N_17202);
or U17313 (N_17313,N_17128,N_17148);
nor U17314 (N_17314,N_17032,N_17012);
or U17315 (N_17315,N_17061,N_17240);
and U17316 (N_17316,N_17229,N_17166);
or U17317 (N_17317,N_17051,N_17053);
nand U17318 (N_17318,N_17247,N_17064);
xnor U17319 (N_17319,N_17186,N_17196);
nor U17320 (N_17320,N_17075,N_17026);
or U17321 (N_17321,N_17036,N_17043);
nor U17322 (N_17322,N_17246,N_17249);
or U17323 (N_17323,N_17116,N_17231);
nand U17324 (N_17324,N_17100,N_17097);
xnor U17325 (N_17325,N_17208,N_17009);
and U17326 (N_17326,N_17126,N_17033);
or U17327 (N_17327,N_17095,N_17226);
nor U17328 (N_17328,N_17028,N_17127);
nand U17329 (N_17329,N_17172,N_17163);
nor U17330 (N_17330,N_17038,N_17121);
xor U17331 (N_17331,N_17118,N_17045);
nor U17332 (N_17332,N_17087,N_17007);
and U17333 (N_17333,N_17234,N_17112);
and U17334 (N_17334,N_17049,N_17083);
and U17335 (N_17335,N_17194,N_17165);
nor U17336 (N_17336,N_17244,N_17101);
nor U17337 (N_17337,N_17014,N_17078);
nand U17338 (N_17338,N_17020,N_17143);
nand U17339 (N_17339,N_17179,N_17207);
nor U17340 (N_17340,N_17132,N_17150);
nand U17341 (N_17341,N_17091,N_17221);
nor U17342 (N_17342,N_17215,N_17129);
nand U17343 (N_17343,N_17206,N_17151);
nor U17344 (N_17344,N_17122,N_17054);
xnor U17345 (N_17345,N_17245,N_17169);
and U17346 (N_17346,N_17204,N_17119);
xor U17347 (N_17347,N_17113,N_17021);
nor U17348 (N_17348,N_17065,N_17082);
nand U17349 (N_17349,N_17180,N_17214);
or U17350 (N_17350,N_17090,N_17037);
nor U17351 (N_17351,N_17085,N_17029);
nand U17352 (N_17352,N_17048,N_17153);
xnor U17353 (N_17353,N_17139,N_17058);
xor U17354 (N_17354,N_17131,N_17168);
nor U17355 (N_17355,N_17157,N_17167);
nand U17356 (N_17356,N_17146,N_17110);
nor U17357 (N_17357,N_17237,N_17219);
or U17358 (N_17358,N_17188,N_17230);
and U17359 (N_17359,N_17092,N_17135);
and U17360 (N_17360,N_17109,N_17057);
or U17361 (N_17361,N_17030,N_17141);
nor U17362 (N_17362,N_17130,N_17224);
xor U17363 (N_17363,N_17063,N_17193);
xnor U17364 (N_17364,N_17182,N_17147);
nor U17365 (N_17365,N_17099,N_17052);
nor U17366 (N_17366,N_17236,N_17047);
and U17367 (N_17367,N_17222,N_17154);
xor U17368 (N_17368,N_17000,N_17074);
xnor U17369 (N_17369,N_17205,N_17184);
nor U17370 (N_17370,N_17211,N_17183);
and U17371 (N_17371,N_17227,N_17114);
nor U17372 (N_17372,N_17005,N_17239);
nor U17373 (N_17373,N_17142,N_17164);
and U17374 (N_17374,N_17067,N_17159);
xnor U17375 (N_17375,N_17121,N_17103);
nand U17376 (N_17376,N_17101,N_17212);
nor U17377 (N_17377,N_17123,N_17085);
and U17378 (N_17378,N_17126,N_17080);
or U17379 (N_17379,N_17115,N_17046);
or U17380 (N_17380,N_17153,N_17013);
or U17381 (N_17381,N_17223,N_17243);
xor U17382 (N_17382,N_17025,N_17119);
xnor U17383 (N_17383,N_17209,N_17108);
or U17384 (N_17384,N_17112,N_17191);
xnor U17385 (N_17385,N_17193,N_17103);
nor U17386 (N_17386,N_17036,N_17073);
xor U17387 (N_17387,N_17091,N_17005);
nor U17388 (N_17388,N_17077,N_17191);
or U17389 (N_17389,N_17227,N_17090);
or U17390 (N_17390,N_17012,N_17059);
nor U17391 (N_17391,N_17139,N_17020);
nor U17392 (N_17392,N_17177,N_17068);
and U17393 (N_17393,N_17082,N_17245);
and U17394 (N_17394,N_17154,N_17230);
nand U17395 (N_17395,N_17225,N_17003);
nor U17396 (N_17396,N_17193,N_17238);
nor U17397 (N_17397,N_17183,N_17169);
nand U17398 (N_17398,N_17003,N_17231);
nor U17399 (N_17399,N_17075,N_17192);
and U17400 (N_17400,N_17194,N_17091);
and U17401 (N_17401,N_17112,N_17039);
nor U17402 (N_17402,N_17079,N_17010);
nand U17403 (N_17403,N_17190,N_17218);
nand U17404 (N_17404,N_17074,N_17218);
or U17405 (N_17405,N_17006,N_17056);
nand U17406 (N_17406,N_17248,N_17014);
xnor U17407 (N_17407,N_17100,N_17108);
and U17408 (N_17408,N_17174,N_17194);
nand U17409 (N_17409,N_17122,N_17049);
nor U17410 (N_17410,N_17071,N_17024);
nand U17411 (N_17411,N_17101,N_17144);
nand U17412 (N_17412,N_17016,N_17091);
nor U17413 (N_17413,N_17107,N_17236);
nand U17414 (N_17414,N_17022,N_17099);
or U17415 (N_17415,N_17144,N_17192);
nand U17416 (N_17416,N_17018,N_17099);
nand U17417 (N_17417,N_17034,N_17127);
and U17418 (N_17418,N_17090,N_17244);
and U17419 (N_17419,N_17145,N_17230);
nand U17420 (N_17420,N_17062,N_17025);
nand U17421 (N_17421,N_17202,N_17037);
xor U17422 (N_17422,N_17007,N_17225);
nand U17423 (N_17423,N_17095,N_17126);
or U17424 (N_17424,N_17006,N_17244);
nand U17425 (N_17425,N_17154,N_17066);
xor U17426 (N_17426,N_17016,N_17055);
nor U17427 (N_17427,N_17091,N_17150);
nor U17428 (N_17428,N_17111,N_17107);
and U17429 (N_17429,N_17099,N_17083);
or U17430 (N_17430,N_17016,N_17028);
xor U17431 (N_17431,N_17147,N_17028);
nor U17432 (N_17432,N_17112,N_17216);
xor U17433 (N_17433,N_17140,N_17067);
nor U17434 (N_17434,N_17179,N_17246);
and U17435 (N_17435,N_17044,N_17123);
and U17436 (N_17436,N_17087,N_17033);
nand U17437 (N_17437,N_17111,N_17248);
and U17438 (N_17438,N_17092,N_17158);
xor U17439 (N_17439,N_17156,N_17089);
nand U17440 (N_17440,N_17038,N_17201);
and U17441 (N_17441,N_17228,N_17141);
nand U17442 (N_17442,N_17085,N_17249);
and U17443 (N_17443,N_17087,N_17156);
and U17444 (N_17444,N_17244,N_17069);
nand U17445 (N_17445,N_17047,N_17092);
xor U17446 (N_17446,N_17000,N_17238);
or U17447 (N_17447,N_17103,N_17008);
xnor U17448 (N_17448,N_17215,N_17003);
xor U17449 (N_17449,N_17217,N_17210);
or U17450 (N_17450,N_17222,N_17210);
and U17451 (N_17451,N_17046,N_17065);
and U17452 (N_17452,N_17178,N_17207);
nand U17453 (N_17453,N_17145,N_17054);
and U17454 (N_17454,N_17213,N_17230);
xor U17455 (N_17455,N_17248,N_17133);
nand U17456 (N_17456,N_17098,N_17061);
or U17457 (N_17457,N_17237,N_17141);
and U17458 (N_17458,N_17166,N_17215);
and U17459 (N_17459,N_17213,N_17224);
and U17460 (N_17460,N_17154,N_17127);
xor U17461 (N_17461,N_17067,N_17041);
xor U17462 (N_17462,N_17231,N_17181);
xnor U17463 (N_17463,N_17127,N_17067);
nand U17464 (N_17464,N_17039,N_17009);
or U17465 (N_17465,N_17234,N_17216);
xor U17466 (N_17466,N_17125,N_17109);
and U17467 (N_17467,N_17207,N_17098);
or U17468 (N_17468,N_17177,N_17210);
nand U17469 (N_17469,N_17122,N_17019);
xnor U17470 (N_17470,N_17182,N_17129);
nand U17471 (N_17471,N_17232,N_17050);
nor U17472 (N_17472,N_17208,N_17196);
nand U17473 (N_17473,N_17072,N_17139);
nand U17474 (N_17474,N_17004,N_17200);
xnor U17475 (N_17475,N_17029,N_17100);
nand U17476 (N_17476,N_17046,N_17040);
nand U17477 (N_17477,N_17064,N_17101);
nor U17478 (N_17478,N_17235,N_17180);
and U17479 (N_17479,N_17198,N_17228);
xor U17480 (N_17480,N_17103,N_17164);
xor U17481 (N_17481,N_17089,N_17184);
nand U17482 (N_17482,N_17198,N_17246);
nor U17483 (N_17483,N_17245,N_17085);
or U17484 (N_17484,N_17187,N_17113);
xnor U17485 (N_17485,N_17182,N_17177);
nor U17486 (N_17486,N_17174,N_17160);
or U17487 (N_17487,N_17075,N_17025);
nor U17488 (N_17488,N_17161,N_17207);
nand U17489 (N_17489,N_17071,N_17139);
nor U17490 (N_17490,N_17100,N_17094);
and U17491 (N_17491,N_17151,N_17030);
xor U17492 (N_17492,N_17100,N_17241);
and U17493 (N_17493,N_17000,N_17012);
or U17494 (N_17494,N_17142,N_17092);
nand U17495 (N_17495,N_17034,N_17075);
nand U17496 (N_17496,N_17023,N_17108);
or U17497 (N_17497,N_17227,N_17038);
nor U17498 (N_17498,N_17026,N_17111);
xor U17499 (N_17499,N_17239,N_17108);
and U17500 (N_17500,N_17450,N_17359);
or U17501 (N_17501,N_17288,N_17404);
xnor U17502 (N_17502,N_17340,N_17490);
or U17503 (N_17503,N_17270,N_17266);
and U17504 (N_17504,N_17291,N_17473);
and U17505 (N_17505,N_17397,N_17337);
or U17506 (N_17506,N_17376,N_17495);
and U17507 (N_17507,N_17487,N_17349);
or U17508 (N_17508,N_17371,N_17332);
nand U17509 (N_17509,N_17287,N_17293);
nor U17510 (N_17510,N_17488,N_17427);
or U17511 (N_17511,N_17420,N_17369);
or U17512 (N_17512,N_17400,N_17477);
and U17513 (N_17513,N_17372,N_17381);
xor U17514 (N_17514,N_17446,N_17452);
or U17515 (N_17515,N_17363,N_17407);
nand U17516 (N_17516,N_17358,N_17274);
and U17517 (N_17517,N_17252,N_17442);
or U17518 (N_17518,N_17364,N_17492);
nand U17519 (N_17519,N_17365,N_17254);
nor U17520 (N_17520,N_17464,N_17317);
xnor U17521 (N_17521,N_17290,N_17297);
nor U17522 (N_17522,N_17341,N_17257);
or U17523 (N_17523,N_17405,N_17497);
nor U17524 (N_17524,N_17251,N_17451);
and U17525 (N_17525,N_17258,N_17296);
or U17526 (N_17526,N_17294,N_17449);
and U17527 (N_17527,N_17489,N_17322);
and U17528 (N_17528,N_17467,N_17283);
nand U17529 (N_17529,N_17466,N_17457);
or U17530 (N_17530,N_17289,N_17484);
nor U17531 (N_17531,N_17319,N_17463);
nand U17532 (N_17532,N_17444,N_17267);
nand U17533 (N_17533,N_17391,N_17379);
and U17534 (N_17534,N_17438,N_17327);
nor U17535 (N_17535,N_17282,N_17356);
and U17536 (N_17536,N_17277,N_17494);
nor U17537 (N_17537,N_17261,N_17269);
xor U17538 (N_17538,N_17271,N_17394);
xor U17539 (N_17539,N_17250,N_17308);
xnor U17540 (N_17540,N_17314,N_17279);
and U17541 (N_17541,N_17348,N_17368);
nand U17542 (N_17542,N_17421,N_17302);
and U17543 (N_17543,N_17307,N_17262);
or U17544 (N_17544,N_17309,N_17426);
and U17545 (N_17545,N_17375,N_17284);
or U17546 (N_17546,N_17433,N_17455);
nor U17547 (N_17547,N_17292,N_17469);
nor U17548 (N_17548,N_17280,N_17414);
nand U17549 (N_17549,N_17318,N_17393);
nor U17550 (N_17550,N_17441,N_17324);
nand U17551 (N_17551,N_17483,N_17440);
nand U17552 (N_17552,N_17431,N_17298);
or U17553 (N_17553,N_17498,N_17333);
or U17554 (N_17554,N_17478,N_17499);
or U17555 (N_17555,N_17351,N_17328);
or U17556 (N_17556,N_17265,N_17355);
nand U17557 (N_17557,N_17264,N_17461);
and U17558 (N_17558,N_17462,N_17260);
nand U17559 (N_17559,N_17415,N_17476);
nand U17560 (N_17560,N_17413,N_17485);
nand U17561 (N_17561,N_17326,N_17272);
and U17562 (N_17562,N_17346,N_17361);
xor U17563 (N_17563,N_17417,N_17419);
or U17564 (N_17564,N_17353,N_17479);
nor U17565 (N_17565,N_17447,N_17315);
nand U17566 (N_17566,N_17336,N_17338);
or U17567 (N_17567,N_17387,N_17325);
nor U17568 (N_17568,N_17301,N_17378);
nand U17569 (N_17569,N_17422,N_17275);
and U17570 (N_17570,N_17286,N_17360);
or U17571 (N_17571,N_17395,N_17345);
or U17572 (N_17572,N_17408,N_17295);
or U17573 (N_17573,N_17439,N_17352);
or U17574 (N_17574,N_17278,N_17320);
xnor U17575 (N_17575,N_17475,N_17403);
or U17576 (N_17576,N_17425,N_17418);
xnor U17577 (N_17577,N_17316,N_17386);
and U17578 (N_17578,N_17383,N_17370);
xor U17579 (N_17579,N_17273,N_17263);
and U17580 (N_17580,N_17402,N_17474);
and U17581 (N_17581,N_17334,N_17374);
xor U17582 (N_17582,N_17435,N_17367);
nand U17583 (N_17583,N_17472,N_17330);
nor U17584 (N_17584,N_17411,N_17373);
nand U17585 (N_17585,N_17470,N_17256);
and U17586 (N_17586,N_17434,N_17350);
nor U17587 (N_17587,N_17276,N_17382);
nand U17588 (N_17588,N_17362,N_17313);
nor U17589 (N_17589,N_17305,N_17268);
nand U17590 (N_17590,N_17304,N_17311);
or U17591 (N_17591,N_17259,N_17392);
xnor U17592 (N_17592,N_17357,N_17401);
xor U17593 (N_17593,N_17456,N_17299);
or U17594 (N_17594,N_17335,N_17253);
and U17595 (N_17595,N_17423,N_17453);
nand U17596 (N_17596,N_17459,N_17329);
or U17597 (N_17597,N_17339,N_17412);
nor U17598 (N_17598,N_17432,N_17380);
or U17599 (N_17599,N_17398,N_17312);
nand U17600 (N_17600,N_17437,N_17390);
nand U17601 (N_17601,N_17396,N_17300);
and U17602 (N_17602,N_17406,N_17306);
xnor U17603 (N_17603,N_17343,N_17255);
nand U17604 (N_17604,N_17429,N_17399);
and U17605 (N_17605,N_17460,N_17445);
nor U17606 (N_17606,N_17436,N_17321);
xnor U17607 (N_17607,N_17486,N_17323);
and U17608 (N_17608,N_17331,N_17468);
xor U17609 (N_17609,N_17310,N_17377);
nand U17610 (N_17610,N_17303,N_17342);
nand U17611 (N_17611,N_17443,N_17281);
nor U17612 (N_17612,N_17416,N_17493);
and U17613 (N_17613,N_17424,N_17430);
xnor U17614 (N_17614,N_17471,N_17366);
nor U17615 (N_17615,N_17448,N_17458);
and U17616 (N_17616,N_17409,N_17480);
nand U17617 (N_17617,N_17428,N_17410);
and U17618 (N_17618,N_17454,N_17496);
nor U17619 (N_17619,N_17385,N_17388);
xor U17620 (N_17620,N_17465,N_17354);
or U17621 (N_17621,N_17491,N_17482);
nor U17622 (N_17622,N_17344,N_17481);
nor U17623 (N_17623,N_17285,N_17347);
or U17624 (N_17624,N_17384,N_17389);
nand U17625 (N_17625,N_17410,N_17393);
xnor U17626 (N_17626,N_17369,N_17467);
and U17627 (N_17627,N_17479,N_17450);
xnor U17628 (N_17628,N_17453,N_17461);
or U17629 (N_17629,N_17264,N_17352);
or U17630 (N_17630,N_17321,N_17475);
and U17631 (N_17631,N_17437,N_17395);
or U17632 (N_17632,N_17425,N_17257);
and U17633 (N_17633,N_17330,N_17256);
nand U17634 (N_17634,N_17252,N_17306);
or U17635 (N_17635,N_17449,N_17325);
or U17636 (N_17636,N_17490,N_17435);
or U17637 (N_17637,N_17367,N_17451);
xnor U17638 (N_17638,N_17276,N_17446);
or U17639 (N_17639,N_17440,N_17420);
and U17640 (N_17640,N_17259,N_17362);
xor U17641 (N_17641,N_17465,N_17350);
nor U17642 (N_17642,N_17487,N_17384);
or U17643 (N_17643,N_17468,N_17303);
nand U17644 (N_17644,N_17301,N_17408);
or U17645 (N_17645,N_17427,N_17250);
nor U17646 (N_17646,N_17445,N_17467);
xor U17647 (N_17647,N_17411,N_17260);
xnor U17648 (N_17648,N_17435,N_17483);
nand U17649 (N_17649,N_17458,N_17365);
nand U17650 (N_17650,N_17429,N_17413);
xor U17651 (N_17651,N_17479,N_17433);
and U17652 (N_17652,N_17335,N_17299);
nand U17653 (N_17653,N_17415,N_17279);
nand U17654 (N_17654,N_17261,N_17378);
and U17655 (N_17655,N_17497,N_17410);
or U17656 (N_17656,N_17389,N_17464);
or U17657 (N_17657,N_17465,N_17343);
or U17658 (N_17658,N_17438,N_17381);
and U17659 (N_17659,N_17324,N_17253);
and U17660 (N_17660,N_17481,N_17285);
and U17661 (N_17661,N_17320,N_17412);
and U17662 (N_17662,N_17356,N_17435);
nand U17663 (N_17663,N_17393,N_17445);
or U17664 (N_17664,N_17322,N_17295);
xor U17665 (N_17665,N_17278,N_17289);
nor U17666 (N_17666,N_17280,N_17388);
xnor U17667 (N_17667,N_17462,N_17335);
and U17668 (N_17668,N_17373,N_17299);
nand U17669 (N_17669,N_17273,N_17364);
nand U17670 (N_17670,N_17425,N_17434);
xor U17671 (N_17671,N_17304,N_17336);
or U17672 (N_17672,N_17453,N_17375);
and U17673 (N_17673,N_17286,N_17254);
nand U17674 (N_17674,N_17336,N_17322);
xnor U17675 (N_17675,N_17443,N_17339);
and U17676 (N_17676,N_17302,N_17389);
nor U17677 (N_17677,N_17276,N_17493);
nor U17678 (N_17678,N_17496,N_17463);
or U17679 (N_17679,N_17386,N_17371);
xor U17680 (N_17680,N_17252,N_17498);
or U17681 (N_17681,N_17264,N_17434);
nor U17682 (N_17682,N_17259,N_17366);
or U17683 (N_17683,N_17339,N_17453);
and U17684 (N_17684,N_17434,N_17463);
nand U17685 (N_17685,N_17325,N_17492);
nand U17686 (N_17686,N_17384,N_17499);
xnor U17687 (N_17687,N_17499,N_17476);
nor U17688 (N_17688,N_17282,N_17417);
nand U17689 (N_17689,N_17466,N_17250);
xor U17690 (N_17690,N_17304,N_17348);
xor U17691 (N_17691,N_17383,N_17462);
nor U17692 (N_17692,N_17489,N_17365);
xor U17693 (N_17693,N_17313,N_17467);
or U17694 (N_17694,N_17430,N_17451);
or U17695 (N_17695,N_17260,N_17458);
and U17696 (N_17696,N_17491,N_17332);
and U17697 (N_17697,N_17434,N_17335);
and U17698 (N_17698,N_17283,N_17483);
and U17699 (N_17699,N_17285,N_17271);
xor U17700 (N_17700,N_17277,N_17251);
nand U17701 (N_17701,N_17444,N_17271);
or U17702 (N_17702,N_17416,N_17287);
xor U17703 (N_17703,N_17298,N_17349);
xnor U17704 (N_17704,N_17313,N_17364);
nand U17705 (N_17705,N_17385,N_17372);
or U17706 (N_17706,N_17362,N_17327);
nor U17707 (N_17707,N_17330,N_17314);
nand U17708 (N_17708,N_17497,N_17386);
and U17709 (N_17709,N_17401,N_17261);
nand U17710 (N_17710,N_17255,N_17351);
or U17711 (N_17711,N_17261,N_17275);
and U17712 (N_17712,N_17461,N_17382);
nor U17713 (N_17713,N_17449,N_17424);
or U17714 (N_17714,N_17466,N_17358);
nand U17715 (N_17715,N_17276,N_17427);
xor U17716 (N_17716,N_17465,N_17279);
and U17717 (N_17717,N_17296,N_17287);
and U17718 (N_17718,N_17331,N_17285);
xnor U17719 (N_17719,N_17477,N_17292);
nand U17720 (N_17720,N_17489,N_17415);
and U17721 (N_17721,N_17439,N_17422);
or U17722 (N_17722,N_17283,N_17457);
or U17723 (N_17723,N_17438,N_17282);
nand U17724 (N_17724,N_17365,N_17452);
nor U17725 (N_17725,N_17348,N_17350);
or U17726 (N_17726,N_17443,N_17373);
or U17727 (N_17727,N_17432,N_17491);
xor U17728 (N_17728,N_17385,N_17479);
nand U17729 (N_17729,N_17335,N_17293);
nand U17730 (N_17730,N_17381,N_17469);
nor U17731 (N_17731,N_17364,N_17478);
and U17732 (N_17732,N_17404,N_17348);
nand U17733 (N_17733,N_17459,N_17282);
nand U17734 (N_17734,N_17459,N_17261);
and U17735 (N_17735,N_17366,N_17475);
nand U17736 (N_17736,N_17467,N_17319);
or U17737 (N_17737,N_17478,N_17316);
xnor U17738 (N_17738,N_17475,N_17438);
and U17739 (N_17739,N_17364,N_17366);
or U17740 (N_17740,N_17492,N_17408);
nand U17741 (N_17741,N_17481,N_17253);
or U17742 (N_17742,N_17318,N_17306);
nand U17743 (N_17743,N_17365,N_17414);
xnor U17744 (N_17744,N_17252,N_17460);
nand U17745 (N_17745,N_17417,N_17458);
xnor U17746 (N_17746,N_17363,N_17298);
nand U17747 (N_17747,N_17401,N_17264);
xor U17748 (N_17748,N_17458,N_17333);
xnor U17749 (N_17749,N_17398,N_17434);
and U17750 (N_17750,N_17744,N_17505);
or U17751 (N_17751,N_17624,N_17689);
and U17752 (N_17752,N_17585,N_17661);
and U17753 (N_17753,N_17727,N_17721);
nand U17754 (N_17754,N_17641,N_17679);
or U17755 (N_17755,N_17672,N_17576);
and U17756 (N_17756,N_17587,N_17570);
nand U17757 (N_17757,N_17539,N_17739);
and U17758 (N_17758,N_17725,N_17552);
xnor U17759 (N_17759,N_17710,N_17536);
and U17760 (N_17760,N_17655,N_17559);
and U17761 (N_17761,N_17521,N_17583);
nand U17762 (N_17762,N_17690,N_17514);
xnor U17763 (N_17763,N_17598,N_17632);
nor U17764 (N_17764,N_17662,N_17605);
xnor U17765 (N_17765,N_17577,N_17666);
nor U17766 (N_17766,N_17674,N_17633);
and U17767 (N_17767,N_17664,N_17504);
nor U17768 (N_17768,N_17707,N_17647);
xnor U17769 (N_17769,N_17635,N_17729);
and U17770 (N_17770,N_17522,N_17698);
nor U17771 (N_17771,N_17606,N_17659);
and U17772 (N_17772,N_17665,N_17591);
and U17773 (N_17773,N_17601,N_17733);
xnor U17774 (N_17774,N_17720,N_17555);
nor U17775 (N_17775,N_17676,N_17600);
and U17776 (N_17776,N_17748,N_17611);
nand U17777 (N_17777,N_17584,N_17702);
xor U17778 (N_17778,N_17640,N_17560);
and U17779 (N_17779,N_17506,N_17708);
xor U17780 (N_17780,N_17706,N_17531);
or U17781 (N_17781,N_17718,N_17656);
nand U17782 (N_17782,N_17700,N_17716);
and U17783 (N_17783,N_17714,N_17648);
or U17784 (N_17784,N_17678,N_17630);
nor U17785 (N_17785,N_17609,N_17722);
nor U17786 (N_17786,N_17580,N_17743);
and U17787 (N_17787,N_17503,N_17594);
or U17788 (N_17788,N_17529,N_17623);
nand U17789 (N_17789,N_17534,N_17510);
and U17790 (N_17790,N_17586,N_17533);
xor U17791 (N_17791,N_17596,N_17711);
and U17792 (N_17792,N_17554,N_17651);
and U17793 (N_17793,N_17582,N_17557);
nor U17794 (N_17794,N_17625,N_17681);
xnor U17795 (N_17795,N_17546,N_17592);
and U17796 (N_17796,N_17738,N_17588);
or U17797 (N_17797,N_17513,N_17572);
xnor U17798 (N_17798,N_17613,N_17682);
and U17799 (N_17799,N_17553,N_17564);
nor U17800 (N_17800,N_17525,N_17571);
nand U17801 (N_17801,N_17634,N_17631);
nand U17802 (N_17802,N_17684,N_17516);
nor U17803 (N_17803,N_17565,N_17537);
nand U17804 (N_17804,N_17696,N_17699);
nor U17805 (N_17805,N_17532,N_17701);
and U17806 (N_17806,N_17691,N_17616);
nor U17807 (N_17807,N_17512,N_17567);
nand U17808 (N_17808,N_17603,N_17642);
or U17809 (N_17809,N_17671,N_17535);
nor U17810 (N_17810,N_17740,N_17660);
and U17811 (N_17811,N_17590,N_17541);
nand U17812 (N_17812,N_17734,N_17686);
nand U17813 (N_17813,N_17728,N_17599);
and U17814 (N_17814,N_17717,N_17735);
xor U17815 (N_17815,N_17575,N_17742);
nand U17816 (N_17816,N_17578,N_17500);
xnor U17817 (N_17817,N_17548,N_17747);
xnor U17818 (N_17818,N_17677,N_17704);
and U17819 (N_17819,N_17637,N_17658);
nand U17820 (N_17820,N_17589,N_17629);
nand U17821 (N_17821,N_17502,N_17602);
xnor U17822 (N_17822,N_17610,N_17675);
nor U17823 (N_17823,N_17712,N_17581);
nand U17824 (N_17824,N_17719,N_17593);
nor U17825 (N_17825,N_17526,N_17618);
xnor U17826 (N_17826,N_17524,N_17544);
and U17827 (N_17827,N_17545,N_17643);
nand U17828 (N_17828,N_17668,N_17579);
nand U17829 (N_17829,N_17713,N_17670);
nand U17830 (N_17830,N_17501,N_17741);
nor U17831 (N_17831,N_17680,N_17562);
nor U17832 (N_17832,N_17644,N_17723);
nand U17833 (N_17833,N_17509,N_17694);
and U17834 (N_17834,N_17683,N_17528);
and U17835 (N_17835,N_17550,N_17638);
nand U17836 (N_17836,N_17551,N_17507);
nand U17837 (N_17837,N_17523,N_17566);
and U17838 (N_17838,N_17558,N_17745);
xor U17839 (N_17839,N_17621,N_17703);
or U17840 (N_17840,N_17673,N_17724);
nor U17841 (N_17841,N_17517,N_17732);
or U17842 (N_17842,N_17619,N_17568);
or U17843 (N_17843,N_17607,N_17697);
or U17844 (N_17844,N_17574,N_17604);
xnor U17845 (N_17845,N_17737,N_17622);
nor U17846 (N_17846,N_17620,N_17650);
or U17847 (N_17847,N_17569,N_17573);
and U17848 (N_17848,N_17612,N_17730);
xor U17849 (N_17849,N_17511,N_17547);
nand U17850 (N_17850,N_17692,N_17561);
nand U17851 (N_17851,N_17542,N_17636);
xnor U17852 (N_17852,N_17540,N_17628);
xnor U17853 (N_17853,N_17726,N_17652);
or U17854 (N_17854,N_17687,N_17508);
and U17855 (N_17855,N_17614,N_17688);
nor U17856 (N_17856,N_17654,N_17519);
nand U17857 (N_17857,N_17608,N_17657);
nand U17858 (N_17858,N_17515,N_17595);
or U17859 (N_17859,N_17663,N_17695);
nor U17860 (N_17860,N_17746,N_17669);
nand U17861 (N_17861,N_17538,N_17653);
or U17862 (N_17862,N_17626,N_17646);
or U17863 (N_17863,N_17736,N_17543);
nor U17864 (N_17864,N_17715,N_17749);
and U17865 (N_17865,N_17731,N_17627);
xnor U17866 (N_17866,N_17649,N_17667);
nand U17867 (N_17867,N_17527,N_17563);
or U17868 (N_17868,N_17709,N_17615);
nor U17869 (N_17869,N_17556,N_17518);
and U17870 (N_17870,N_17639,N_17693);
and U17871 (N_17871,N_17597,N_17705);
nand U17872 (N_17872,N_17645,N_17530);
or U17873 (N_17873,N_17685,N_17549);
nand U17874 (N_17874,N_17520,N_17617);
nor U17875 (N_17875,N_17604,N_17659);
and U17876 (N_17876,N_17650,N_17626);
and U17877 (N_17877,N_17535,N_17749);
or U17878 (N_17878,N_17643,N_17592);
xor U17879 (N_17879,N_17727,N_17742);
nor U17880 (N_17880,N_17635,N_17626);
xor U17881 (N_17881,N_17598,N_17688);
or U17882 (N_17882,N_17614,N_17511);
nand U17883 (N_17883,N_17549,N_17635);
or U17884 (N_17884,N_17639,N_17524);
or U17885 (N_17885,N_17705,N_17739);
nand U17886 (N_17886,N_17726,N_17564);
xnor U17887 (N_17887,N_17687,N_17666);
xor U17888 (N_17888,N_17749,N_17694);
nor U17889 (N_17889,N_17553,N_17648);
and U17890 (N_17890,N_17547,N_17526);
and U17891 (N_17891,N_17623,N_17628);
nand U17892 (N_17892,N_17566,N_17630);
nand U17893 (N_17893,N_17703,N_17624);
nand U17894 (N_17894,N_17592,N_17523);
or U17895 (N_17895,N_17665,N_17712);
nand U17896 (N_17896,N_17662,N_17634);
or U17897 (N_17897,N_17517,N_17640);
xnor U17898 (N_17898,N_17736,N_17719);
nand U17899 (N_17899,N_17557,N_17618);
nor U17900 (N_17900,N_17665,N_17558);
nand U17901 (N_17901,N_17565,N_17732);
xor U17902 (N_17902,N_17698,N_17724);
and U17903 (N_17903,N_17623,N_17684);
and U17904 (N_17904,N_17674,N_17540);
xnor U17905 (N_17905,N_17682,N_17675);
xnor U17906 (N_17906,N_17701,N_17636);
and U17907 (N_17907,N_17727,N_17649);
xor U17908 (N_17908,N_17611,N_17573);
and U17909 (N_17909,N_17651,N_17708);
or U17910 (N_17910,N_17571,N_17635);
and U17911 (N_17911,N_17678,N_17704);
nand U17912 (N_17912,N_17656,N_17501);
xor U17913 (N_17913,N_17516,N_17542);
nor U17914 (N_17914,N_17697,N_17614);
or U17915 (N_17915,N_17691,N_17665);
xnor U17916 (N_17916,N_17691,N_17682);
nor U17917 (N_17917,N_17682,N_17610);
nand U17918 (N_17918,N_17551,N_17747);
xor U17919 (N_17919,N_17596,N_17575);
and U17920 (N_17920,N_17527,N_17533);
nor U17921 (N_17921,N_17582,N_17585);
or U17922 (N_17922,N_17699,N_17581);
nand U17923 (N_17923,N_17667,N_17627);
nor U17924 (N_17924,N_17659,N_17522);
xor U17925 (N_17925,N_17588,N_17696);
nand U17926 (N_17926,N_17508,N_17542);
nor U17927 (N_17927,N_17543,N_17696);
or U17928 (N_17928,N_17712,N_17619);
nor U17929 (N_17929,N_17533,N_17561);
nand U17930 (N_17930,N_17530,N_17730);
xor U17931 (N_17931,N_17555,N_17675);
nor U17932 (N_17932,N_17555,N_17525);
nand U17933 (N_17933,N_17707,N_17596);
nand U17934 (N_17934,N_17694,N_17500);
or U17935 (N_17935,N_17578,N_17641);
and U17936 (N_17936,N_17607,N_17510);
xnor U17937 (N_17937,N_17523,N_17706);
and U17938 (N_17938,N_17607,N_17676);
nand U17939 (N_17939,N_17517,N_17507);
or U17940 (N_17940,N_17575,N_17503);
xor U17941 (N_17941,N_17684,N_17598);
and U17942 (N_17942,N_17543,N_17540);
xnor U17943 (N_17943,N_17504,N_17623);
or U17944 (N_17944,N_17596,N_17736);
or U17945 (N_17945,N_17655,N_17515);
or U17946 (N_17946,N_17636,N_17592);
nand U17947 (N_17947,N_17626,N_17618);
or U17948 (N_17948,N_17734,N_17673);
nand U17949 (N_17949,N_17594,N_17718);
and U17950 (N_17950,N_17675,N_17515);
xor U17951 (N_17951,N_17663,N_17680);
xnor U17952 (N_17952,N_17703,N_17738);
nand U17953 (N_17953,N_17651,N_17655);
or U17954 (N_17954,N_17653,N_17639);
xnor U17955 (N_17955,N_17708,N_17720);
nor U17956 (N_17956,N_17666,N_17697);
nand U17957 (N_17957,N_17555,N_17684);
xor U17958 (N_17958,N_17596,N_17700);
or U17959 (N_17959,N_17557,N_17558);
xor U17960 (N_17960,N_17748,N_17628);
nand U17961 (N_17961,N_17508,N_17680);
or U17962 (N_17962,N_17526,N_17558);
nor U17963 (N_17963,N_17602,N_17721);
xnor U17964 (N_17964,N_17615,N_17742);
nand U17965 (N_17965,N_17558,N_17533);
or U17966 (N_17966,N_17701,N_17688);
nor U17967 (N_17967,N_17704,N_17621);
nor U17968 (N_17968,N_17573,N_17509);
xor U17969 (N_17969,N_17645,N_17705);
and U17970 (N_17970,N_17677,N_17601);
and U17971 (N_17971,N_17514,N_17683);
and U17972 (N_17972,N_17715,N_17550);
nor U17973 (N_17973,N_17566,N_17710);
and U17974 (N_17974,N_17656,N_17666);
and U17975 (N_17975,N_17613,N_17510);
nand U17976 (N_17976,N_17734,N_17520);
nand U17977 (N_17977,N_17510,N_17725);
or U17978 (N_17978,N_17503,N_17631);
and U17979 (N_17979,N_17734,N_17566);
or U17980 (N_17980,N_17620,N_17711);
and U17981 (N_17981,N_17680,N_17689);
or U17982 (N_17982,N_17575,N_17628);
and U17983 (N_17983,N_17583,N_17525);
or U17984 (N_17984,N_17747,N_17666);
nand U17985 (N_17985,N_17693,N_17740);
and U17986 (N_17986,N_17512,N_17684);
nand U17987 (N_17987,N_17726,N_17501);
nor U17988 (N_17988,N_17687,N_17513);
and U17989 (N_17989,N_17585,N_17709);
or U17990 (N_17990,N_17574,N_17697);
nor U17991 (N_17991,N_17746,N_17513);
or U17992 (N_17992,N_17662,N_17716);
xnor U17993 (N_17993,N_17652,N_17691);
or U17994 (N_17994,N_17662,N_17562);
or U17995 (N_17995,N_17664,N_17506);
or U17996 (N_17996,N_17555,N_17744);
nor U17997 (N_17997,N_17591,N_17526);
xor U17998 (N_17998,N_17543,N_17662);
or U17999 (N_17999,N_17500,N_17531);
nor U18000 (N_18000,N_17809,N_17850);
xnor U18001 (N_18001,N_17853,N_17756);
and U18002 (N_18002,N_17958,N_17990);
xor U18003 (N_18003,N_17764,N_17901);
nor U18004 (N_18004,N_17861,N_17895);
or U18005 (N_18005,N_17827,N_17769);
or U18006 (N_18006,N_17968,N_17855);
xnor U18007 (N_18007,N_17800,N_17925);
nor U18008 (N_18008,N_17869,N_17902);
and U18009 (N_18009,N_17971,N_17888);
and U18010 (N_18010,N_17911,N_17859);
nand U18011 (N_18011,N_17998,N_17914);
xor U18012 (N_18012,N_17900,N_17808);
xnor U18013 (N_18013,N_17930,N_17829);
xnor U18014 (N_18014,N_17944,N_17819);
xnor U18015 (N_18015,N_17943,N_17908);
or U18016 (N_18016,N_17789,N_17860);
or U18017 (N_18017,N_17757,N_17781);
nand U18018 (N_18018,N_17933,N_17897);
nand U18019 (N_18019,N_17937,N_17843);
xor U18020 (N_18020,N_17976,N_17903);
nor U18021 (N_18021,N_17940,N_17817);
nand U18022 (N_18022,N_17951,N_17836);
and U18023 (N_18023,N_17982,N_17967);
nand U18024 (N_18024,N_17820,N_17913);
nand U18025 (N_18025,N_17934,N_17965);
or U18026 (N_18026,N_17785,N_17847);
xnor U18027 (N_18027,N_17852,N_17771);
xor U18028 (N_18028,N_17985,N_17912);
xor U18029 (N_18029,N_17765,N_17953);
xor U18030 (N_18030,N_17851,N_17961);
or U18031 (N_18031,N_17876,N_17926);
nor U18032 (N_18032,N_17779,N_17891);
nor U18033 (N_18033,N_17833,N_17812);
or U18034 (N_18034,N_17862,N_17773);
nor U18035 (N_18035,N_17882,N_17919);
xnor U18036 (N_18036,N_17793,N_17831);
nor U18037 (N_18037,N_17893,N_17910);
xnor U18038 (N_18038,N_17830,N_17797);
and U18039 (N_18039,N_17999,N_17814);
xor U18040 (N_18040,N_17811,N_17906);
xor U18041 (N_18041,N_17916,N_17865);
nand U18042 (N_18042,N_17794,N_17837);
or U18043 (N_18043,N_17768,N_17766);
and U18044 (N_18044,N_17993,N_17863);
and U18045 (N_18045,N_17981,N_17992);
nand U18046 (N_18046,N_17870,N_17818);
or U18047 (N_18047,N_17890,N_17783);
nand U18048 (N_18048,N_17894,N_17872);
and U18049 (N_18049,N_17755,N_17962);
nor U18050 (N_18050,N_17776,N_17989);
nor U18051 (N_18051,N_17938,N_17883);
nor U18052 (N_18052,N_17871,N_17762);
nor U18053 (N_18053,N_17973,N_17979);
nor U18054 (N_18054,N_17966,N_17777);
xnor U18055 (N_18055,N_17878,N_17884);
xnor U18056 (N_18056,N_17879,N_17824);
or U18057 (N_18057,N_17904,N_17864);
nand U18058 (N_18058,N_17898,N_17774);
nand U18059 (N_18059,N_17942,N_17795);
nand U18060 (N_18060,N_17841,N_17763);
or U18061 (N_18061,N_17828,N_17950);
xor U18062 (N_18062,N_17801,N_17946);
and U18063 (N_18063,N_17972,N_17915);
nand U18064 (N_18064,N_17886,N_17987);
nand U18065 (N_18065,N_17767,N_17846);
and U18066 (N_18066,N_17923,N_17994);
and U18067 (N_18067,N_17881,N_17826);
nor U18068 (N_18068,N_17945,N_17845);
nand U18069 (N_18069,N_17751,N_17821);
and U18070 (N_18070,N_17866,N_17957);
or U18071 (N_18071,N_17935,N_17840);
nor U18072 (N_18072,N_17799,N_17991);
nor U18073 (N_18073,N_17856,N_17835);
nor U18074 (N_18074,N_17932,N_17980);
and U18075 (N_18075,N_17778,N_17752);
nand U18076 (N_18076,N_17970,N_17997);
xnor U18077 (N_18077,N_17917,N_17792);
nor U18078 (N_18078,N_17754,N_17928);
or U18079 (N_18079,N_17813,N_17877);
nand U18080 (N_18080,N_17905,N_17875);
and U18081 (N_18081,N_17995,N_17782);
or U18082 (N_18082,N_17802,N_17924);
or U18083 (N_18083,N_17796,N_17868);
nor U18084 (N_18084,N_17839,N_17758);
and U18085 (N_18085,N_17939,N_17867);
and U18086 (N_18086,N_17874,N_17775);
nand U18087 (N_18087,N_17844,N_17936);
xnor U18088 (N_18088,N_17984,N_17931);
and U18089 (N_18089,N_17803,N_17770);
or U18090 (N_18090,N_17988,N_17963);
nand U18091 (N_18091,N_17947,N_17975);
or U18092 (N_18092,N_17804,N_17909);
and U18093 (N_18093,N_17927,N_17823);
nand U18094 (N_18094,N_17815,N_17996);
or U18095 (N_18095,N_17892,N_17948);
and U18096 (N_18096,N_17873,N_17887);
and U18097 (N_18097,N_17986,N_17952);
or U18098 (N_18098,N_17918,N_17791);
xor U18099 (N_18099,N_17949,N_17806);
and U18100 (N_18100,N_17974,N_17816);
and U18101 (N_18101,N_17822,N_17848);
or U18102 (N_18102,N_17896,N_17920);
or U18103 (N_18103,N_17825,N_17899);
xor U18104 (N_18104,N_17964,N_17955);
nor U18105 (N_18105,N_17842,N_17978);
nand U18106 (N_18106,N_17807,N_17772);
nand U18107 (N_18107,N_17922,N_17929);
xnor U18108 (N_18108,N_17983,N_17805);
xnor U18109 (N_18109,N_17857,N_17788);
or U18110 (N_18110,N_17907,N_17977);
and U18111 (N_18111,N_17810,N_17838);
or U18112 (N_18112,N_17956,N_17780);
and U18113 (N_18113,N_17798,N_17832);
and U18114 (N_18114,N_17959,N_17854);
nand U18115 (N_18115,N_17889,N_17759);
xnor U18116 (N_18116,N_17760,N_17761);
or U18117 (N_18117,N_17790,N_17834);
xnor U18118 (N_18118,N_17969,N_17954);
nor U18119 (N_18119,N_17885,N_17786);
and U18120 (N_18120,N_17787,N_17880);
xnor U18121 (N_18121,N_17921,N_17753);
and U18122 (N_18122,N_17858,N_17960);
or U18123 (N_18123,N_17849,N_17750);
nand U18124 (N_18124,N_17941,N_17784);
and U18125 (N_18125,N_17812,N_17844);
xnor U18126 (N_18126,N_17850,N_17865);
xnor U18127 (N_18127,N_17992,N_17954);
xnor U18128 (N_18128,N_17914,N_17810);
nor U18129 (N_18129,N_17770,N_17856);
xor U18130 (N_18130,N_17958,N_17882);
nor U18131 (N_18131,N_17778,N_17905);
xnor U18132 (N_18132,N_17923,N_17856);
nand U18133 (N_18133,N_17804,N_17850);
nor U18134 (N_18134,N_17880,N_17772);
nand U18135 (N_18135,N_17946,N_17845);
nor U18136 (N_18136,N_17931,N_17904);
or U18137 (N_18137,N_17894,N_17932);
or U18138 (N_18138,N_17851,N_17843);
nor U18139 (N_18139,N_17845,N_17883);
or U18140 (N_18140,N_17917,N_17834);
or U18141 (N_18141,N_17832,N_17963);
nand U18142 (N_18142,N_17780,N_17989);
or U18143 (N_18143,N_17863,N_17953);
xnor U18144 (N_18144,N_17883,N_17779);
xnor U18145 (N_18145,N_17819,N_17762);
nand U18146 (N_18146,N_17879,N_17988);
and U18147 (N_18147,N_17792,N_17964);
nand U18148 (N_18148,N_17838,N_17768);
or U18149 (N_18149,N_17775,N_17841);
nor U18150 (N_18150,N_17787,N_17921);
and U18151 (N_18151,N_17914,N_17813);
and U18152 (N_18152,N_17814,N_17897);
nand U18153 (N_18153,N_17840,N_17774);
nand U18154 (N_18154,N_17823,N_17949);
nor U18155 (N_18155,N_17760,N_17776);
nor U18156 (N_18156,N_17766,N_17891);
xnor U18157 (N_18157,N_17834,N_17991);
and U18158 (N_18158,N_17847,N_17911);
xor U18159 (N_18159,N_17774,N_17783);
xnor U18160 (N_18160,N_17951,N_17840);
nor U18161 (N_18161,N_17997,N_17900);
xor U18162 (N_18162,N_17861,N_17954);
and U18163 (N_18163,N_17929,N_17752);
nand U18164 (N_18164,N_17887,N_17905);
or U18165 (N_18165,N_17923,N_17876);
and U18166 (N_18166,N_17985,N_17995);
nand U18167 (N_18167,N_17828,N_17838);
nor U18168 (N_18168,N_17906,N_17903);
xor U18169 (N_18169,N_17877,N_17976);
nand U18170 (N_18170,N_17758,N_17800);
and U18171 (N_18171,N_17846,N_17834);
nand U18172 (N_18172,N_17807,N_17920);
nor U18173 (N_18173,N_17768,N_17870);
or U18174 (N_18174,N_17978,N_17863);
nand U18175 (N_18175,N_17914,N_17984);
and U18176 (N_18176,N_17914,N_17790);
nor U18177 (N_18177,N_17977,N_17778);
xnor U18178 (N_18178,N_17948,N_17999);
or U18179 (N_18179,N_17991,N_17951);
xnor U18180 (N_18180,N_17771,N_17839);
and U18181 (N_18181,N_17908,N_17768);
nor U18182 (N_18182,N_17881,N_17757);
nand U18183 (N_18183,N_17911,N_17848);
and U18184 (N_18184,N_17786,N_17754);
or U18185 (N_18185,N_17906,N_17963);
nor U18186 (N_18186,N_17853,N_17919);
nand U18187 (N_18187,N_17896,N_17841);
nand U18188 (N_18188,N_17890,N_17981);
nor U18189 (N_18189,N_17767,N_17824);
or U18190 (N_18190,N_17847,N_17838);
nor U18191 (N_18191,N_17979,N_17910);
xor U18192 (N_18192,N_17983,N_17756);
nor U18193 (N_18193,N_17872,N_17959);
nor U18194 (N_18194,N_17751,N_17815);
xor U18195 (N_18195,N_17888,N_17861);
or U18196 (N_18196,N_17825,N_17823);
nand U18197 (N_18197,N_17986,N_17887);
nor U18198 (N_18198,N_17831,N_17822);
and U18199 (N_18199,N_17918,N_17876);
nand U18200 (N_18200,N_17947,N_17759);
nand U18201 (N_18201,N_17990,N_17868);
nor U18202 (N_18202,N_17756,N_17838);
and U18203 (N_18203,N_17768,N_17921);
and U18204 (N_18204,N_17815,N_17960);
nor U18205 (N_18205,N_17969,N_17949);
nand U18206 (N_18206,N_17909,N_17753);
xor U18207 (N_18207,N_17819,N_17832);
and U18208 (N_18208,N_17798,N_17810);
nor U18209 (N_18209,N_17815,N_17841);
or U18210 (N_18210,N_17947,N_17920);
or U18211 (N_18211,N_17826,N_17907);
xor U18212 (N_18212,N_17793,N_17877);
nor U18213 (N_18213,N_17901,N_17779);
xnor U18214 (N_18214,N_17898,N_17927);
or U18215 (N_18215,N_17911,N_17767);
or U18216 (N_18216,N_17792,N_17766);
xnor U18217 (N_18217,N_17751,N_17963);
nor U18218 (N_18218,N_17891,N_17797);
and U18219 (N_18219,N_17829,N_17828);
xnor U18220 (N_18220,N_17767,N_17768);
nand U18221 (N_18221,N_17769,N_17832);
nor U18222 (N_18222,N_17891,N_17903);
nor U18223 (N_18223,N_17974,N_17812);
nand U18224 (N_18224,N_17906,N_17837);
xor U18225 (N_18225,N_17956,N_17850);
or U18226 (N_18226,N_17854,N_17769);
or U18227 (N_18227,N_17884,N_17880);
nand U18228 (N_18228,N_17752,N_17788);
nor U18229 (N_18229,N_17909,N_17828);
and U18230 (N_18230,N_17784,N_17880);
nand U18231 (N_18231,N_17872,N_17865);
or U18232 (N_18232,N_17821,N_17877);
and U18233 (N_18233,N_17907,N_17988);
xor U18234 (N_18234,N_17884,N_17889);
and U18235 (N_18235,N_17986,N_17810);
or U18236 (N_18236,N_17957,N_17953);
and U18237 (N_18237,N_17849,N_17971);
or U18238 (N_18238,N_17984,N_17925);
or U18239 (N_18239,N_17864,N_17891);
and U18240 (N_18240,N_17926,N_17998);
nand U18241 (N_18241,N_17952,N_17886);
or U18242 (N_18242,N_17929,N_17800);
nand U18243 (N_18243,N_17952,N_17972);
and U18244 (N_18244,N_17917,N_17805);
nor U18245 (N_18245,N_17831,N_17857);
and U18246 (N_18246,N_17883,N_17778);
or U18247 (N_18247,N_17991,N_17835);
xnor U18248 (N_18248,N_17834,N_17864);
xnor U18249 (N_18249,N_17904,N_17767);
and U18250 (N_18250,N_18249,N_18163);
and U18251 (N_18251,N_18117,N_18169);
or U18252 (N_18252,N_18122,N_18164);
and U18253 (N_18253,N_18191,N_18020);
or U18254 (N_18254,N_18107,N_18167);
nand U18255 (N_18255,N_18081,N_18067);
xnor U18256 (N_18256,N_18111,N_18057);
and U18257 (N_18257,N_18084,N_18120);
nand U18258 (N_18258,N_18039,N_18037);
and U18259 (N_18259,N_18017,N_18166);
xor U18260 (N_18260,N_18140,N_18233);
nor U18261 (N_18261,N_18152,N_18075);
nor U18262 (N_18262,N_18192,N_18129);
xor U18263 (N_18263,N_18123,N_18068);
and U18264 (N_18264,N_18069,N_18059);
and U18265 (N_18265,N_18098,N_18034);
xor U18266 (N_18266,N_18132,N_18235);
xor U18267 (N_18267,N_18238,N_18156);
nand U18268 (N_18268,N_18145,N_18025);
nand U18269 (N_18269,N_18224,N_18093);
nor U18270 (N_18270,N_18179,N_18199);
nand U18271 (N_18271,N_18147,N_18012);
xor U18272 (N_18272,N_18027,N_18142);
and U18273 (N_18273,N_18110,N_18230);
and U18274 (N_18274,N_18174,N_18097);
nor U18275 (N_18275,N_18205,N_18248);
or U18276 (N_18276,N_18103,N_18089);
nand U18277 (N_18277,N_18058,N_18095);
nor U18278 (N_18278,N_18109,N_18004);
nor U18279 (N_18279,N_18204,N_18134);
xnor U18280 (N_18280,N_18211,N_18241);
and U18281 (N_18281,N_18116,N_18023);
nand U18282 (N_18282,N_18159,N_18065);
or U18283 (N_18283,N_18155,N_18185);
and U18284 (N_18284,N_18055,N_18042);
xnor U18285 (N_18285,N_18050,N_18128);
and U18286 (N_18286,N_18126,N_18106);
or U18287 (N_18287,N_18138,N_18019);
and U18288 (N_18288,N_18146,N_18049);
nand U18289 (N_18289,N_18045,N_18108);
or U18290 (N_18290,N_18150,N_18178);
nor U18291 (N_18291,N_18086,N_18193);
nor U18292 (N_18292,N_18009,N_18130);
xnor U18293 (N_18293,N_18066,N_18112);
or U18294 (N_18294,N_18182,N_18043);
and U18295 (N_18295,N_18143,N_18162);
or U18296 (N_18296,N_18048,N_18018);
and U18297 (N_18297,N_18007,N_18079);
and U18298 (N_18298,N_18061,N_18035);
nand U18299 (N_18299,N_18070,N_18047);
nor U18300 (N_18300,N_18137,N_18113);
xor U18301 (N_18301,N_18209,N_18168);
nand U18302 (N_18302,N_18078,N_18060);
and U18303 (N_18303,N_18215,N_18114);
xnor U18304 (N_18304,N_18160,N_18234);
and U18305 (N_18305,N_18139,N_18076);
nor U18306 (N_18306,N_18006,N_18180);
or U18307 (N_18307,N_18090,N_18104);
xor U18308 (N_18308,N_18008,N_18038);
and U18309 (N_18309,N_18172,N_18206);
or U18310 (N_18310,N_18022,N_18030);
xor U18311 (N_18311,N_18054,N_18127);
and U18312 (N_18312,N_18237,N_18125);
nand U18313 (N_18313,N_18202,N_18198);
nor U18314 (N_18314,N_18197,N_18208);
nand U18315 (N_18315,N_18005,N_18131);
and U18316 (N_18316,N_18212,N_18175);
nand U18317 (N_18317,N_18196,N_18053);
xor U18318 (N_18318,N_18032,N_18165);
xnor U18319 (N_18319,N_18072,N_18223);
nor U18320 (N_18320,N_18136,N_18148);
nor U18321 (N_18321,N_18201,N_18228);
nand U18322 (N_18322,N_18056,N_18176);
and U18323 (N_18323,N_18064,N_18010);
nand U18324 (N_18324,N_18082,N_18216);
or U18325 (N_18325,N_18229,N_18244);
and U18326 (N_18326,N_18195,N_18013);
nand U18327 (N_18327,N_18016,N_18243);
xnor U18328 (N_18328,N_18207,N_18121);
xnor U18329 (N_18329,N_18100,N_18040);
nor U18330 (N_18330,N_18063,N_18170);
xnor U18331 (N_18331,N_18141,N_18015);
nor U18332 (N_18332,N_18231,N_18183);
or U18333 (N_18333,N_18073,N_18135);
xor U18334 (N_18334,N_18221,N_18133);
or U18335 (N_18335,N_18000,N_18033);
xor U18336 (N_18336,N_18083,N_18219);
and U18337 (N_18337,N_18149,N_18203);
xor U18338 (N_18338,N_18115,N_18157);
xnor U18339 (N_18339,N_18220,N_18002);
or U18340 (N_18340,N_18124,N_18003);
nand U18341 (N_18341,N_18080,N_18217);
xor U18342 (N_18342,N_18046,N_18210);
or U18343 (N_18343,N_18052,N_18227);
xnor U18344 (N_18344,N_18181,N_18184);
or U18345 (N_18345,N_18247,N_18190);
nand U18346 (N_18346,N_18099,N_18161);
nand U18347 (N_18347,N_18186,N_18001);
or U18348 (N_18348,N_18077,N_18200);
nand U18349 (N_18349,N_18188,N_18239);
nand U18350 (N_18350,N_18026,N_18213);
and U18351 (N_18351,N_18091,N_18242);
nor U18352 (N_18352,N_18119,N_18173);
and U18353 (N_18353,N_18194,N_18021);
nor U18354 (N_18354,N_18158,N_18101);
nand U18355 (N_18355,N_18088,N_18096);
or U18356 (N_18356,N_18171,N_18085);
xnor U18357 (N_18357,N_18071,N_18029);
or U18358 (N_18358,N_18031,N_18151);
or U18359 (N_18359,N_18218,N_18245);
and U18360 (N_18360,N_18062,N_18222);
xor U18361 (N_18361,N_18225,N_18153);
and U18362 (N_18362,N_18177,N_18051);
nor U18363 (N_18363,N_18226,N_18074);
nand U18364 (N_18364,N_18187,N_18144);
nand U18365 (N_18365,N_18118,N_18041);
and U18366 (N_18366,N_18011,N_18240);
and U18367 (N_18367,N_18092,N_18232);
and U18368 (N_18368,N_18087,N_18028);
and U18369 (N_18369,N_18044,N_18014);
xor U18370 (N_18370,N_18105,N_18214);
or U18371 (N_18371,N_18246,N_18094);
nor U18372 (N_18372,N_18102,N_18154);
nand U18373 (N_18373,N_18236,N_18189);
nor U18374 (N_18374,N_18036,N_18024);
or U18375 (N_18375,N_18213,N_18221);
xnor U18376 (N_18376,N_18152,N_18041);
nor U18377 (N_18377,N_18078,N_18192);
and U18378 (N_18378,N_18137,N_18016);
nor U18379 (N_18379,N_18067,N_18189);
nand U18380 (N_18380,N_18079,N_18011);
or U18381 (N_18381,N_18051,N_18049);
xnor U18382 (N_18382,N_18223,N_18018);
nor U18383 (N_18383,N_18158,N_18202);
and U18384 (N_18384,N_18242,N_18172);
nor U18385 (N_18385,N_18129,N_18002);
nor U18386 (N_18386,N_18135,N_18097);
nor U18387 (N_18387,N_18187,N_18129);
nor U18388 (N_18388,N_18079,N_18189);
or U18389 (N_18389,N_18217,N_18222);
and U18390 (N_18390,N_18101,N_18229);
xor U18391 (N_18391,N_18221,N_18111);
and U18392 (N_18392,N_18062,N_18068);
nor U18393 (N_18393,N_18086,N_18119);
and U18394 (N_18394,N_18145,N_18176);
and U18395 (N_18395,N_18208,N_18183);
or U18396 (N_18396,N_18050,N_18245);
nor U18397 (N_18397,N_18240,N_18132);
xnor U18398 (N_18398,N_18131,N_18157);
nor U18399 (N_18399,N_18106,N_18026);
xnor U18400 (N_18400,N_18121,N_18017);
and U18401 (N_18401,N_18059,N_18244);
nor U18402 (N_18402,N_18170,N_18232);
nand U18403 (N_18403,N_18140,N_18015);
and U18404 (N_18404,N_18019,N_18136);
nor U18405 (N_18405,N_18019,N_18114);
and U18406 (N_18406,N_18106,N_18017);
nand U18407 (N_18407,N_18076,N_18182);
nor U18408 (N_18408,N_18060,N_18065);
nor U18409 (N_18409,N_18234,N_18224);
nand U18410 (N_18410,N_18059,N_18129);
nor U18411 (N_18411,N_18020,N_18009);
and U18412 (N_18412,N_18210,N_18070);
or U18413 (N_18413,N_18211,N_18165);
nand U18414 (N_18414,N_18106,N_18011);
nand U18415 (N_18415,N_18173,N_18147);
or U18416 (N_18416,N_18083,N_18134);
xnor U18417 (N_18417,N_18165,N_18135);
and U18418 (N_18418,N_18051,N_18150);
and U18419 (N_18419,N_18169,N_18190);
and U18420 (N_18420,N_18094,N_18025);
and U18421 (N_18421,N_18096,N_18151);
xnor U18422 (N_18422,N_18227,N_18096);
xnor U18423 (N_18423,N_18063,N_18246);
and U18424 (N_18424,N_18222,N_18135);
nor U18425 (N_18425,N_18180,N_18018);
xnor U18426 (N_18426,N_18194,N_18094);
or U18427 (N_18427,N_18181,N_18105);
and U18428 (N_18428,N_18200,N_18231);
xor U18429 (N_18429,N_18038,N_18145);
or U18430 (N_18430,N_18019,N_18017);
and U18431 (N_18431,N_18122,N_18022);
nand U18432 (N_18432,N_18048,N_18039);
and U18433 (N_18433,N_18169,N_18058);
and U18434 (N_18434,N_18177,N_18214);
nor U18435 (N_18435,N_18065,N_18247);
or U18436 (N_18436,N_18008,N_18136);
nor U18437 (N_18437,N_18107,N_18045);
or U18438 (N_18438,N_18136,N_18216);
and U18439 (N_18439,N_18017,N_18042);
nor U18440 (N_18440,N_18232,N_18000);
nor U18441 (N_18441,N_18132,N_18089);
nor U18442 (N_18442,N_18057,N_18139);
xor U18443 (N_18443,N_18052,N_18053);
nor U18444 (N_18444,N_18103,N_18021);
nand U18445 (N_18445,N_18136,N_18246);
or U18446 (N_18446,N_18111,N_18154);
xnor U18447 (N_18447,N_18060,N_18142);
nor U18448 (N_18448,N_18229,N_18210);
xor U18449 (N_18449,N_18168,N_18240);
nor U18450 (N_18450,N_18024,N_18109);
and U18451 (N_18451,N_18233,N_18006);
and U18452 (N_18452,N_18227,N_18209);
or U18453 (N_18453,N_18095,N_18232);
nor U18454 (N_18454,N_18199,N_18122);
xor U18455 (N_18455,N_18057,N_18219);
or U18456 (N_18456,N_18061,N_18090);
and U18457 (N_18457,N_18018,N_18136);
nor U18458 (N_18458,N_18025,N_18238);
or U18459 (N_18459,N_18192,N_18156);
and U18460 (N_18460,N_18046,N_18164);
and U18461 (N_18461,N_18225,N_18042);
xnor U18462 (N_18462,N_18000,N_18205);
and U18463 (N_18463,N_18225,N_18040);
and U18464 (N_18464,N_18193,N_18129);
nor U18465 (N_18465,N_18169,N_18152);
and U18466 (N_18466,N_18036,N_18111);
and U18467 (N_18467,N_18043,N_18130);
nand U18468 (N_18468,N_18127,N_18112);
and U18469 (N_18469,N_18048,N_18044);
nor U18470 (N_18470,N_18072,N_18011);
nor U18471 (N_18471,N_18222,N_18225);
nor U18472 (N_18472,N_18187,N_18012);
nor U18473 (N_18473,N_18180,N_18119);
xor U18474 (N_18474,N_18185,N_18063);
xor U18475 (N_18475,N_18017,N_18114);
xor U18476 (N_18476,N_18168,N_18166);
or U18477 (N_18477,N_18235,N_18233);
nor U18478 (N_18478,N_18127,N_18247);
nor U18479 (N_18479,N_18065,N_18158);
xnor U18480 (N_18480,N_18051,N_18214);
nand U18481 (N_18481,N_18227,N_18159);
nor U18482 (N_18482,N_18035,N_18164);
nor U18483 (N_18483,N_18003,N_18234);
and U18484 (N_18484,N_18213,N_18222);
nor U18485 (N_18485,N_18148,N_18147);
xnor U18486 (N_18486,N_18204,N_18066);
nand U18487 (N_18487,N_18047,N_18188);
or U18488 (N_18488,N_18123,N_18065);
nand U18489 (N_18489,N_18207,N_18141);
or U18490 (N_18490,N_18026,N_18115);
and U18491 (N_18491,N_18164,N_18076);
or U18492 (N_18492,N_18232,N_18008);
xnor U18493 (N_18493,N_18195,N_18187);
nand U18494 (N_18494,N_18150,N_18038);
xnor U18495 (N_18495,N_18116,N_18033);
nand U18496 (N_18496,N_18061,N_18051);
or U18497 (N_18497,N_18056,N_18004);
nor U18498 (N_18498,N_18077,N_18157);
and U18499 (N_18499,N_18183,N_18134);
or U18500 (N_18500,N_18461,N_18388);
nand U18501 (N_18501,N_18276,N_18292);
and U18502 (N_18502,N_18280,N_18434);
and U18503 (N_18503,N_18382,N_18321);
and U18504 (N_18504,N_18410,N_18486);
xnor U18505 (N_18505,N_18272,N_18497);
and U18506 (N_18506,N_18416,N_18275);
nand U18507 (N_18507,N_18265,N_18438);
or U18508 (N_18508,N_18312,N_18347);
nor U18509 (N_18509,N_18268,N_18444);
nor U18510 (N_18510,N_18267,N_18354);
xnor U18511 (N_18511,N_18291,N_18311);
xnor U18512 (N_18512,N_18339,N_18274);
nor U18513 (N_18513,N_18282,N_18398);
or U18514 (N_18514,N_18258,N_18458);
nor U18515 (N_18515,N_18278,N_18430);
nor U18516 (N_18516,N_18432,N_18447);
or U18517 (N_18517,N_18273,N_18484);
nand U18518 (N_18518,N_18346,N_18426);
xor U18519 (N_18519,N_18331,N_18300);
nor U18520 (N_18520,N_18355,N_18390);
nand U18521 (N_18521,N_18452,N_18489);
nor U18522 (N_18522,N_18492,N_18387);
or U18523 (N_18523,N_18397,N_18304);
nor U18524 (N_18524,N_18361,N_18368);
and U18525 (N_18525,N_18362,N_18270);
xnor U18526 (N_18526,N_18401,N_18257);
nand U18527 (N_18527,N_18456,N_18499);
nor U18528 (N_18528,N_18404,N_18442);
and U18529 (N_18529,N_18472,N_18261);
nor U18530 (N_18530,N_18328,N_18468);
and U18531 (N_18531,N_18356,N_18408);
or U18532 (N_18532,N_18467,N_18310);
xnor U18533 (N_18533,N_18418,N_18476);
and U18534 (N_18534,N_18289,N_18393);
and U18535 (N_18535,N_18365,N_18448);
and U18536 (N_18536,N_18422,N_18303);
or U18537 (N_18537,N_18396,N_18457);
nand U18538 (N_18538,N_18329,N_18378);
or U18539 (N_18539,N_18302,N_18252);
xnor U18540 (N_18540,N_18412,N_18464);
or U18541 (N_18541,N_18419,N_18394);
xnor U18542 (N_18542,N_18478,N_18399);
nor U18543 (N_18543,N_18309,N_18392);
or U18544 (N_18544,N_18322,N_18255);
or U18545 (N_18545,N_18384,N_18470);
or U18546 (N_18546,N_18495,N_18395);
xnor U18547 (N_18547,N_18305,N_18324);
nor U18548 (N_18548,N_18498,N_18315);
xor U18549 (N_18549,N_18420,N_18333);
and U18550 (N_18550,N_18307,N_18443);
nand U18551 (N_18551,N_18294,N_18372);
nor U18552 (N_18552,N_18367,N_18488);
and U18553 (N_18553,N_18423,N_18296);
nand U18554 (N_18554,N_18327,N_18479);
xor U18555 (N_18555,N_18421,N_18440);
nor U18556 (N_18556,N_18415,N_18375);
xnor U18557 (N_18557,N_18451,N_18454);
and U18558 (N_18558,N_18364,N_18407);
and U18559 (N_18559,N_18429,N_18373);
nand U18560 (N_18560,N_18449,N_18259);
xnor U18561 (N_18561,N_18348,N_18370);
nor U18562 (N_18562,N_18334,N_18344);
xor U18563 (N_18563,N_18424,N_18474);
and U18564 (N_18564,N_18316,N_18299);
xnor U18565 (N_18565,N_18301,N_18284);
xnor U18566 (N_18566,N_18250,N_18383);
and U18567 (N_18567,N_18357,N_18330);
xor U18568 (N_18568,N_18379,N_18336);
nand U18569 (N_18569,N_18471,N_18460);
or U18570 (N_18570,N_18369,N_18473);
nor U18571 (N_18571,N_18350,N_18481);
nand U18572 (N_18572,N_18253,N_18260);
nand U18573 (N_18573,N_18343,N_18462);
or U18574 (N_18574,N_18433,N_18437);
xnor U18575 (N_18575,N_18264,N_18459);
nor U18576 (N_18576,N_18431,N_18405);
and U18577 (N_18577,N_18435,N_18288);
nand U18578 (N_18578,N_18279,N_18269);
and U18579 (N_18579,N_18385,N_18493);
xor U18580 (N_18580,N_18469,N_18286);
nand U18581 (N_18581,N_18256,N_18290);
or U18582 (N_18582,N_18446,N_18389);
or U18583 (N_18583,N_18317,N_18323);
nor U18584 (N_18584,N_18381,N_18360);
or U18585 (N_18585,N_18425,N_18358);
or U18586 (N_18586,N_18428,N_18411);
or U18587 (N_18587,N_18337,N_18445);
nand U18588 (N_18588,N_18298,N_18262);
nor U18589 (N_18589,N_18455,N_18340);
and U18590 (N_18590,N_18406,N_18342);
nor U18591 (N_18591,N_18271,N_18487);
xor U18592 (N_18592,N_18313,N_18319);
and U18593 (N_18593,N_18494,N_18453);
nor U18594 (N_18594,N_18482,N_18439);
xnor U18595 (N_18595,N_18293,N_18353);
nand U18596 (N_18596,N_18266,N_18326);
or U18597 (N_18597,N_18281,N_18251);
nand U18598 (N_18598,N_18475,N_18402);
and U18599 (N_18599,N_18436,N_18283);
and U18600 (N_18600,N_18263,N_18254);
nand U18601 (N_18601,N_18485,N_18277);
and U18602 (N_18602,N_18466,N_18349);
and U18603 (N_18603,N_18359,N_18409);
nor U18604 (N_18604,N_18377,N_18376);
and U18605 (N_18605,N_18335,N_18351);
nor U18606 (N_18606,N_18363,N_18374);
and U18607 (N_18607,N_18325,N_18338);
and U18608 (N_18608,N_18318,N_18441);
xnor U18609 (N_18609,N_18491,N_18332);
nand U18610 (N_18610,N_18341,N_18427);
xnor U18611 (N_18611,N_18366,N_18297);
xor U18612 (N_18612,N_18496,N_18391);
and U18613 (N_18613,N_18450,N_18465);
or U18614 (N_18614,N_18483,N_18308);
and U18615 (N_18615,N_18287,N_18463);
nor U18616 (N_18616,N_18320,N_18314);
nand U18617 (N_18617,N_18417,N_18403);
xnor U18618 (N_18618,N_18306,N_18477);
nor U18619 (N_18619,N_18371,N_18285);
xnor U18620 (N_18620,N_18413,N_18414);
xor U18621 (N_18621,N_18490,N_18295);
nand U18622 (N_18622,N_18480,N_18352);
and U18623 (N_18623,N_18380,N_18400);
xnor U18624 (N_18624,N_18386,N_18345);
or U18625 (N_18625,N_18253,N_18498);
xor U18626 (N_18626,N_18480,N_18333);
xor U18627 (N_18627,N_18434,N_18325);
nor U18628 (N_18628,N_18360,N_18385);
nor U18629 (N_18629,N_18321,N_18346);
nor U18630 (N_18630,N_18499,N_18387);
and U18631 (N_18631,N_18494,N_18289);
xor U18632 (N_18632,N_18485,N_18284);
xnor U18633 (N_18633,N_18297,N_18296);
nor U18634 (N_18634,N_18468,N_18341);
xor U18635 (N_18635,N_18333,N_18290);
nand U18636 (N_18636,N_18372,N_18441);
or U18637 (N_18637,N_18418,N_18320);
and U18638 (N_18638,N_18422,N_18260);
xor U18639 (N_18639,N_18372,N_18388);
and U18640 (N_18640,N_18405,N_18445);
and U18641 (N_18641,N_18395,N_18402);
nor U18642 (N_18642,N_18442,N_18346);
xnor U18643 (N_18643,N_18318,N_18413);
nor U18644 (N_18644,N_18299,N_18391);
or U18645 (N_18645,N_18476,N_18424);
nor U18646 (N_18646,N_18435,N_18426);
or U18647 (N_18647,N_18363,N_18357);
and U18648 (N_18648,N_18379,N_18439);
and U18649 (N_18649,N_18284,N_18368);
and U18650 (N_18650,N_18339,N_18300);
nand U18651 (N_18651,N_18473,N_18319);
nand U18652 (N_18652,N_18353,N_18416);
nor U18653 (N_18653,N_18406,N_18381);
and U18654 (N_18654,N_18301,N_18262);
and U18655 (N_18655,N_18360,N_18271);
nand U18656 (N_18656,N_18497,N_18442);
nor U18657 (N_18657,N_18450,N_18378);
and U18658 (N_18658,N_18452,N_18427);
xor U18659 (N_18659,N_18455,N_18361);
nor U18660 (N_18660,N_18468,N_18470);
or U18661 (N_18661,N_18327,N_18359);
or U18662 (N_18662,N_18290,N_18258);
or U18663 (N_18663,N_18487,N_18398);
or U18664 (N_18664,N_18270,N_18402);
nand U18665 (N_18665,N_18471,N_18270);
nor U18666 (N_18666,N_18437,N_18430);
nor U18667 (N_18667,N_18472,N_18311);
and U18668 (N_18668,N_18317,N_18497);
or U18669 (N_18669,N_18377,N_18302);
nor U18670 (N_18670,N_18315,N_18422);
nor U18671 (N_18671,N_18323,N_18390);
nor U18672 (N_18672,N_18413,N_18493);
xnor U18673 (N_18673,N_18405,N_18350);
nand U18674 (N_18674,N_18289,N_18300);
nand U18675 (N_18675,N_18311,N_18400);
nand U18676 (N_18676,N_18400,N_18307);
and U18677 (N_18677,N_18384,N_18252);
nor U18678 (N_18678,N_18456,N_18263);
xnor U18679 (N_18679,N_18280,N_18315);
and U18680 (N_18680,N_18472,N_18316);
nand U18681 (N_18681,N_18379,N_18410);
nor U18682 (N_18682,N_18423,N_18487);
nand U18683 (N_18683,N_18323,N_18327);
xnor U18684 (N_18684,N_18422,N_18370);
nor U18685 (N_18685,N_18289,N_18421);
nor U18686 (N_18686,N_18262,N_18375);
and U18687 (N_18687,N_18473,N_18488);
nor U18688 (N_18688,N_18448,N_18421);
xnor U18689 (N_18689,N_18397,N_18330);
and U18690 (N_18690,N_18332,N_18412);
xnor U18691 (N_18691,N_18321,N_18400);
or U18692 (N_18692,N_18318,N_18436);
and U18693 (N_18693,N_18347,N_18366);
or U18694 (N_18694,N_18271,N_18275);
and U18695 (N_18695,N_18433,N_18392);
nand U18696 (N_18696,N_18377,N_18362);
nand U18697 (N_18697,N_18280,N_18462);
nor U18698 (N_18698,N_18459,N_18442);
nor U18699 (N_18699,N_18432,N_18474);
nand U18700 (N_18700,N_18462,N_18438);
and U18701 (N_18701,N_18379,N_18394);
nand U18702 (N_18702,N_18290,N_18374);
xnor U18703 (N_18703,N_18260,N_18366);
or U18704 (N_18704,N_18410,N_18323);
nor U18705 (N_18705,N_18337,N_18446);
or U18706 (N_18706,N_18329,N_18280);
nand U18707 (N_18707,N_18452,N_18488);
xnor U18708 (N_18708,N_18389,N_18470);
xor U18709 (N_18709,N_18357,N_18380);
xor U18710 (N_18710,N_18488,N_18425);
and U18711 (N_18711,N_18498,N_18471);
xnor U18712 (N_18712,N_18372,N_18288);
xor U18713 (N_18713,N_18289,N_18381);
nor U18714 (N_18714,N_18342,N_18274);
and U18715 (N_18715,N_18445,N_18312);
xor U18716 (N_18716,N_18495,N_18384);
nor U18717 (N_18717,N_18300,N_18303);
nor U18718 (N_18718,N_18323,N_18395);
nand U18719 (N_18719,N_18276,N_18390);
and U18720 (N_18720,N_18419,N_18264);
and U18721 (N_18721,N_18364,N_18373);
nand U18722 (N_18722,N_18403,N_18300);
and U18723 (N_18723,N_18293,N_18415);
nor U18724 (N_18724,N_18383,N_18282);
nand U18725 (N_18725,N_18299,N_18404);
or U18726 (N_18726,N_18405,N_18353);
nand U18727 (N_18727,N_18420,N_18437);
and U18728 (N_18728,N_18393,N_18423);
and U18729 (N_18729,N_18377,N_18450);
or U18730 (N_18730,N_18392,N_18339);
xnor U18731 (N_18731,N_18250,N_18466);
xor U18732 (N_18732,N_18438,N_18338);
nand U18733 (N_18733,N_18411,N_18412);
or U18734 (N_18734,N_18412,N_18341);
and U18735 (N_18735,N_18275,N_18301);
or U18736 (N_18736,N_18344,N_18311);
or U18737 (N_18737,N_18302,N_18371);
or U18738 (N_18738,N_18458,N_18488);
or U18739 (N_18739,N_18459,N_18255);
nand U18740 (N_18740,N_18462,N_18320);
and U18741 (N_18741,N_18422,N_18280);
and U18742 (N_18742,N_18289,N_18438);
and U18743 (N_18743,N_18487,N_18470);
and U18744 (N_18744,N_18481,N_18407);
and U18745 (N_18745,N_18355,N_18414);
and U18746 (N_18746,N_18271,N_18345);
nor U18747 (N_18747,N_18332,N_18325);
nor U18748 (N_18748,N_18327,N_18345);
or U18749 (N_18749,N_18373,N_18286);
or U18750 (N_18750,N_18692,N_18537);
and U18751 (N_18751,N_18703,N_18723);
xnor U18752 (N_18752,N_18727,N_18680);
and U18753 (N_18753,N_18630,N_18637);
nand U18754 (N_18754,N_18544,N_18597);
or U18755 (N_18755,N_18647,N_18601);
nand U18756 (N_18756,N_18657,N_18574);
nand U18757 (N_18757,N_18747,N_18626);
nand U18758 (N_18758,N_18691,N_18594);
or U18759 (N_18759,N_18618,N_18556);
nand U18760 (N_18760,N_18552,N_18560);
and U18761 (N_18761,N_18698,N_18644);
nand U18762 (N_18762,N_18622,N_18721);
nand U18763 (N_18763,N_18681,N_18504);
or U18764 (N_18764,N_18693,N_18683);
and U18765 (N_18765,N_18539,N_18632);
or U18766 (N_18766,N_18638,N_18641);
xor U18767 (N_18767,N_18586,N_18614);
nand U18768 (N_18768,N_18600,N_18513);
and U18769 (N_18769,N_18643,N_18595);
or U18770 (N_18770,N_18717,N_18652);
or U18771 (N_18771,N_18631,N_18547);
and U18772 (N_18772,N_18533,N_18634);
nor U18773 (N_18773,N_18550,N_18628);
nor U18774 (N_18774,N_18659,N_18598);
xor U18775 (N_18775,N_18682,N_18706);
xor U18776 (N_18776,N_18528,N_18540);
or U18777 (N_18777,N_18509,N_18662);
and U18778 (N_18778,N_18635,N_18542);
or U18779 (N_18779,N_18566,N_18596);
nand U18780 (N_18780,N_18579,N_18715);
xnor U18781 (N_18781,N_18599,N_18620);
nor U18782 (N_18782,N_18732,N_18726);
nor U18783 (N_18783,N_18507,N_18714);
or U18784 (N_18784,N_18615,N_18730);
xnor U18785 (N_18785,N_18650,N_18684);
and U18786 (N_18786,N_18688,N_18526);
nor U18787 (N_18787,N_18593,N_18541);
nand U18788 (N_18788,N_18733,N_18705);
or U18789 (N_18789,N_18604,N_18592);
xnor U18790 (N_18790,N_18745,N_18651);
or U18791 (N_18791,N_18608,N_18720);
or U18792 (N_18792,N_18577,N_18633);
or U18793 (N_18793,N_18653,N_18585);
and U18794 (N_18794,N_18664,N_18661);
nand U18795 (N_18795,N_18561,N_18676);
xnor U18796 (N_18796,N_18654,N_18612);
xnor U18797 (N_18797,N_18736,N_18712);
or U18798 (N_18798,N_18667,N_18518);
nor U18799 (N_18799,N_18591,N_18549);
xor U18800 (N_18800,N_18538,N_18602);
or U18801 (N_18801,N_18567,N_18718);
xor U18802 (N_18802,N_18568,N_18607);
and U18803 (N_18803,N_18700,N_18740);
or U18804 (N_18804,N_18558,N_18534);
nand U18805 (N_18805,N_18695,N_18573);
nor U18806 (N_18806,N_18694,N_18742);
nand U18807 (N_18807,N_18514,N_18731);
and U18808 (N_18808,N_18516,N_18749);
or U18809 (N_18809,N_18645,N_18621);
nor U18810 (N_18810,N_18636,N_18666);
nor U18811 (N_18811,N_18503,N_18512);
and U18812 (N_18812,N_18648,N_18679);
or U18813 (N_18813,N_18575,N_18729);
nor U18814 (N_18814,N_18501,N_18570);
or U18815 (N_18815,N_18519,N_18571);
xnor U18816 (N_18816,N_18738,N_18668);
nand U18817 (N_18817,N_18583,N_18511);
nand U18818 (N_18818,N_18646,N_18725);
xnor U18819 (N_18819,N_18576,N_18527);
xor U18820 (N_18820,N_18524,N_18734);
xor U18821 (N_18821,N_18704,N_18505);
xnor U18822 (N_18822,N_18532,N_18529);
nand U18823 (N_18823,N_18649,N_18702);
xor U18824 (N_18824,N_18707,N_18640);
xnor U18825 (N_18825,N_18611,N_18675);
nor U18826 (N_18826,N_18555,N_18674);
or U18827 (N_18827,N_18642,N_18610);
nor U18828 (N_18828,N_18536,N_18500);
nand U18829 (N_18829,N_18521,N_18605);
xnor U18830 (N_18830,N_18710,N_18673);
nand U18831 (N_18831,N_18701,N_18563);
or U18832 (N_18832,N_18578,N_18656);
xnor U18833 (N_18833,N_18690,N_18724);
xor U18834 (N_18834,N_18590,N_18506);
and U18835 (N_18835,N_18554,N_18587);
and U18836 (N_18836,N_18557,N_18699);
or U18837 (N_18837,N_18746,N_18502);
or U18838 (N_18838,N_18546,N_18580);
or U18839 (N_18839,N_18627,N_18686);
nand U18840 (N_18840,N_18739,N_18617);
or U18841 (N_18841,N_18569,N_18543);
or U18842 (N_18842,N_18551,N_18658);
or U18843 (N_18843,N_18671,N_18625);
nor U18844 (N_18844,N_18711,N_18565);
and U18845 (N_18845,N_18629,N_18741);
or U18846 (N_18846,N_18508,N_18677);
nand U18847 (N_18847,N_18589,N_18722);
nor U18848 (N_18848,N_18535,N_18678);
and U18849 (N_18849,N_18517,N_18553);
nor U18850 (N_18850,N_18584,N_18672);
nor U18851 (N_18851,N_18744,N_18665);
and U18852 (N_18852,N_18623,N_18520);
xor U18853 (N_18853,N_18562,N_18639);
and U18854 (N_18854,N_18748,N_18603);
or U18855 (N_18855,N_18525,N_18619);
xnor U18856 (N_18856,N_18581,N_18588);
and U18857 (N_18857,N_18515,N_18697);
and U18858 (N_18858,N_18559,N_18545);
nor U18859 (N_18859,N_18616,N_18670);
or U18860 (N_18860,N_18685,N_18709);
nor U18861 (N_18861,N_18572,N_18548);
xor U18862 (N_18862,N_18743,N_18522);
or U18863 (N_18863,N_18696,N_18564);
and U18864 (N_18864,N_18606,N_18582);
nor U18865 (N_18865,N_18660,N_18716);
and U18866 (N_18866,N_18713,N_18663);
xor U18867 (N_18867,N_18708,N_18523);
nor U18868 (N_18868,N_18624,N_18655);
nand U18869 (N_18869,N_18728,N_18669);
or U18870 (N_18870,N_18687,N_18735);
or U18871 (N_18871,N_18719,N_18689);
nand U18872 (N_18872,N_18737,N_18530);
xnor U18873 (N_18873,N_18531,N_18613);
xor U18874 (N_18874,N_18510,N_18609);
xor U18875 (N_18875,N_18587,N_18551);
nor U18876 (N_18876,N_18657,N_18705);
or U18877 (N_18877,N_18503,N_18626);
xnor U18878 (N_18878,N_18665,N_18583);
nand U18879 (N_18879,N_18533,N_18645);
xor U18880 (N_18880,N_18581,N_18723);
nor U18881 (N_18881,N_18674,N_18723);
xnor U18882 (N_18882,N_18538,N_18673);
and U18883 (N_18883,N_18678,N_18745);
xor U18884 (N_18884,N_18675,N_18727);
or U18885 (N_18885,N_18574,N_18687);
nand U18886 (N_18886,N_18628,N_18610);
or U18887 (N_18887,N_18510,N_18663);
xor U18888 (N_18888,N_18647,N_18730);
and U18889 (N_18889,N_18666,N_18512);
nand U18890 (N_18890,N_18612,N_18710);
and U18891 (N_18891,N_18554,N_18711);
nand U18892 (N_18892,N_18606,N_18528);
and U18893 (N_18893,N_18638,N_18581);
nand U18894 (N_18894,N_18681,N_18643);
or U18895 (N_18895,N_18635,N_18502);
xor U18896 (N_18896,N_18663,N_18693);
xor U18897 (N_18897,N_18644,N_18686);
and U18898 (N_18898,N_18628,N_18703);
or U18899 (N_18899,N_18508,N_18561);
or U18900 (N_18900,N_18676,N_18595);
and U18901 (N_18901,N_18684,N_18712);
or U18902 (N_18902,N_18509,N_18507);
and U18903 (N_18903,N_18591,N_18608);
or U18904 (N_18904,N_18502,N_18521);
nand U18905 (N_18905,N_18519,N_18586);
nor U18906 (N_18906,N_18587,N_18585);
nor U18907 (N_18907,N_18515,N_18710);
or U18908 (N_18908,N_18673,N_18646);
nand U18909 (N_18909,N_18663,N_18732);
nand U18910 (N_18910,N_18592,N_18681);
nor U18911 (N_18911,N_18576,N_18693);
nor U18912 (N_18912,N_18633,N_18658);
nor U18913 (N_18913,N_18578,N_18560);
nand U18914 (N_18914,N_18712,N_18553);
xnor U18915 (N_18915,N_18531,N_18696);
nand U18916 (N_18916,N_18504,N_18654);
and U18917 (N_18917,N_18618,N_18742);
and U18918 (N_18918,N_18657,N_18686);
xnor U18919 (N_18919,N_18512,N_18589);
nand U18920 (N_18920,N_18566,N_18589);
nor U18921 (N_18921,N_18591,N_18670);
and U18922 (N_18922,N_18677,N_18574);
nor U18923 (N_18923,N_18582,N_18720);
xnor U18924 (N_18924,N_18719,N_18746);
and U18925 (N_18925,N_18507,N_18580);
and U18926 (N_18926,N_18546,N_18531);
xor U18927 (N_18927,N_18696,N_18709);
and U18928 (N_18928,N_18667,N_18554);
or U18929 (N_18929,N_18681,N_18715);
or U18930 (N_18930,N_18648,N_18617);
xor U18931 (N_18931,N_18605,N_18721);
nand U18932 (N_18932,N_18739,N_18517);
nand U18933 (N_18933,N_18563,N_18741);
xor U18934 (N_18934,N_18738,N_18549);
nand U18935 (N_18935,N_18718,N_18566);
nor U18936 (N_18936,N_18660,N_18544);
nand U18937 (N_18937,N_18720,N_18639);
nand U18938 (N_18938,N_18573,N_18523);
nand U18939 (N_18939,N_18622,N_18673);
or U18940 (N_18940,N_18747,N_18712);
nand U18941 (N_18941,N_18551,N_18601);
nand U18942 (N_18942,N_18658,N_18597);
and U18943 (N_18943,N_18725,N_18575);
and U18944 (N_18944,N_18560,N_18532);
or U18945 (N_18945,N_18715,N_18539);
and U18946 (N_18946,N_18699,N_18649);
xor U18947 (N_18947,N_18703,N_18547);
or U18948 (N_18948,N_18580,N_18642);
nor U18949 (N_18949,N_18643,N_18727);
nand U18950 (N_18950,N_18739,N_18725);
and U18951 (N_18951,N_18542,N_18687);
and U18952 (N_18952,N_18502,N_18670);
and U18953 (N_18953,N_18705,N_18523);
nor U18954 (N_18954,N_18748,N_18544);
nor U18955 (N_18955,N_18673,N_18595);
nand U18956 (N_18956,N_18713,N_18509);
nor U18957 (N_18957,N_18722,N_18650);
nand U18958 (N_18958,N_18549,N_18727);
xor U18959 (N_18959,N_18597,N_18556);
nand U18960 (N_18960,N_18593,N_18525);
nor U18961 (N_18961,N_18568,N_18732);
nor U18962 (N_18962,N_18651,N_18595);
xor U18963 (N_18963,N_18610,N_18707);
nand U18964 (N_18964,N_18696,N_18538);
xnor U18965 (N_18965,N_18542,N_18739);
or U18966 (N_18966,N_18628,N_18635);
nor U18967 (N_18967,N_18642,N_18664);
nand U18968 (N_18968,N_18559,N_18633);
xor U18969 (N_18969,N_18579,N_18620);
nor U18970 (N_18970,N_18730,N_18517);
or U18971 (N_18971,N_18513,N_18531);
nor U18972 (N_18972,N_18629,N_18611);
or U18973 (N_18973,N_18580,N_18591);
and U18974 (N_18974,N_18500,N_18648);
or U18975 (N_18975,N_18549,N_18621);
and U18976 (N_18976,N_18571,N_18621);
nand U18977 (N_18977,N_18575,N_18714);
xor U18978 (N_18978,N_18708,N_18613);
nor U18979 (N_18979,N_18730,N_18580);
nor U18980 (N_18980,N_18577,N_18613);
xnor U18981 (N_18981,N_18610,N_18650);
nand U18982 (N_18982,N_18516,N_18696);
nor U18983 (N_18983,N_18541,N_18610);
nand U18984 (N_18984,N_18560,N_18735);
xnor U18985 (N_18985,N_18667,N_18578);
and U18986 (N_18986,N_18568,N_18632);
xnor U18987 (N_18987,N_18605,N_18503);
nor U18988 (N_18988,N_18584,N_18613);
or U18989 (N_18989,N_18504,N_18744);
nand U18990 (N_18990,N_18662,N_18642);
and U18991 (N_18991,N_18623,N_18748);
and U18992 (N_18992,N_18731,N_18587);
nor U18993 (N_18993,N_18717,N_18631);
nand U18994 (N_18994,N_18674,N_18718);
xor U18995 (N_18995,N_18700,N_18564);
or U18996 (N_18996,N_18728,N_18723);
or U18997 (N_18997,N_18662,N_18624);
and U18998 (N_18998,N_18624,N_18665);
nand U18999 (N_18999,N_18726,N_18613);
and U19000 (N_19000,N_18850,N_18843);
nand U19001 (N_19001,N_18998,N_18927);
xnor U19002 (N_19002,N_18768,N_18979);
xor U19003 (N_19003,N_18847,N_18967);
and U19004 (N_19004,N_18878,N_18913);
nor U19005 (N_19005,N_18763,N_18750);
nand U19006 (N_19006,N_18833,N_18958);
nand U19007 (N_19007,N_18925,N_18823);
or U19008 (N_19008,N_18759,N_18947);
nand U19009 (N_19009,N_18882,N_18760);
or U19010 (N_19010,N_18810,N_18941);
nand U19011 (N_19011,N_18803,N_18778);
xnor U19012 (N_19012,N_18963,N_18783);
xor U19013 (N_19013,N_18832,N_18859);
nand U19014 (N_19014,N_18920,N_18918);
or U19015 (N_19015,N_18863,N_18877);
and U19016 (N_19016,N_18813,N_18928);
nand U19017 (N_19017,N_18818,N_18975);
and U19018 (N_19018,N_18966,N_18897);
or U19019 (N_19019,N_18846,N_18828);
or U19020 (N_19020,N_18922,N_18819);
nand U19021 (N_19021,N_18989,N_18899);
or U19022 (N_19022,N_18985,N_18923);
or U19023 (N_19023,N_18964,N_18960);
or U19024 (N_19024,N_18921,N_18860);
nand U19025 (N_19025,N_18868,N_18785);
xor U19026 (N_19026,N_18857,N_18904);
or U19027 (N_19027,N_18786,N_18839);
xor U19028 (N_19028,N_18838,N_18757);
nor U19029 (N_19029,N_18872,N_18996);
and U19030 (N_19030,N_18992,N_18875);
xnor U19031 (N_19031,N_18752,N_18852);
xor U19032 (N_19032,N_18796,N_18933);
xor U19033 (N_19033,N_18802,N_18917);
nor U19034 (N_19034,N_18827,N_18885);
nand U19035 (N_19035,N_18936,N_18952);
or U19036 (N_19036,N_18835,N_18829);
nand U19037 (N_19037,N_18761,N_18800);
xor U19038 (N_19038,N_18926,N_18758);
and U19039 (N_19039,N_18995,N_18999);
nand U19040 (N_19040,N_18861,N_18978);
nor U19041 (N_19041,N_18787,N_18901);
or U19042 (N_19042,N_18915,N_18951);
and U19043 (N_19043,N_18815,N_18983);
or U19044 (N_19044,N_18798,N_18816);
and U19045 (N_19045,N_18971,N_18792);
nand U19046 (N_19046,N_18993,N_18883);
or U19047 (N_19047,N_18948,N_18931);
or U19048 (N_19048,N_18934,N_18826);
xor U19049 (N_19049,N_18869,N_18968);
nand U19050 (N_19050,N_18976,N_18977);
and U19051 (N_19051,N_18943,N_18821);
and U19052 (N_19052,N_18893,N_18900);
and U19053 (N_19053,N_18790,N_18889);
xor U19054 (N_19054,N_18990,N_18765);
xnor U19055 (N_19055,N_18820,N_18884);
nand U19056 (N_19056,N_18780,N_18907);
xor U19057 (N_19057,N_18959,N_18892);
nand U19058 (N_19058,N_18811,N_18804);
or U19059 (N_19059,N_18980,N_18837);
nor U19060 (N_19060,N_18937,N_18895);
nor U19061 (N_19061,N_18806,N_18894);
xnor U19062 (N_19062,N_18962,N_18775);
xor U19063 (N_19063,N_18984,N_18781);
nand U19064 (N_19064,N_18848,N_18944);
xnor U19065 (N_19065,N_18956,N_18845);
nor U19066 (N_19066,N_18880,N_18855);
or U19067 (N_19067,N_18911,N_18957);
xor U19068 (N_19068,N_18879,N_18945);
xor U19069 (N_19069,N_18830,N_18817);
nor U19070 (N_19070,N_18791,N_18997);
nand U19071 (N_19071,N_18942,N_18751);
nor U19072 (N_19072,N_18946,N_18881);
nand U19073 (N_19073,N_18905,N_18844);
nand U19074 (N_19074,N_18896,N_18767);
xnor U19075 (N_19075,N_18909,N_18929);
nand U19076 (N_19076,N_18831,N_18908);
nand U19077 (N_19077,N_18753,N_18797);
nor U19078 (N_19078,N_18981,N_18987);
or U19079 (N_19079,N_18988,N_18939);
and U19080 (N_19080,N_18794,N_18777);
nor U19081 (N_19081,N_18961,N_18914);
xnor U19082 (N_19082,N_18779,N_18849);
nand U19083 (N_19083,N_18795,N_18836);
nand U19084 (N_19084,N_18898,N_18808);
nor U19085 (N_19085,N_18784,N_18822);
nand U19086 (N_19086,N_18772,N_18842);
nand U19087 (N_19087,N_18912,N_18874);
nor U19088 (N_19088,N_18953,N_18867);
or U19089 (N_19089,N_18814,N_18807);
nor U19090 (N_19090,N_18886,N_18812);
and U19091 (N_19091,N_18972,N_18876);
nor U19092 (N_19092,N_18910,N_18940);
and U19093 (N_19093,N_18834,N_18965);
nand U19094 (N_19094,N_18870,N_18764);
or U19095 (N_19095,N_18755,N_18871);
nand U19096 (N_19096,N_18902,N_18991);
and U19097 (N_19097,N_18970,N_18754);
or U19098 (N_19098,N_18935,N_18938);
nor U19099 (N_19099,N_18866,N_18851);
nand U19100 (N_19100,N_18854,N_18776);
xnor U19101 (N_19101,N_18762,N_18973);
xor U19102 (N_19102,N_18986,N_18864);
or U19103 (N_19103,N_18793,N_18888);
nand U19104 (N_19104,N_18805,N_18887);
or U19105 (N_19105,N_18856,N_18969);
and U19106 (N_19106,N_18825,N_18891);
xor U19107 (N_19107,N_18771,N_18954);
xor U19108 (N_19108,N_18789,N_18930);
and U19109 (N_19109,N_18799,N_18809);
xnor U19110 (N_19110,N_18994,N_18853);
nor U19111 (N_19111,N_18862,N_18974);
or U19112 (N_19112,N_18858,N_18769);
nand U19113 (N_19113,N_18903,N_18824);
or U19114 (N_19114,N_18801,N_18919);
xnor U19115 (N_19115,N_18906,N_18955);
xnor U19116 (N_19116,N_18782,N_18774);
and U19117 (N_19117,N_18982,N_18840);
and U19118 (N_19118,N_18770,N_18773);
or U19119 (N_19119,N_18932,N_18766);
xor U19120 (N_19120,N_18756,N_18949);
nor U19121 (N_19121,N_18873,N_18916);
and U19122 (N_19122,N_18841,N_18950);
xnor U19123 (N_19123,N_18865,N_18788);
xnor U19124 (N_19124,N_18890,N_18924);
or U19125 (N_19125,N_18883,N_18826);
nand U19126 (N_19126,N_18871,N_18953);
xor U19127 (N_19127,N_18896,N_18919);
and U19128 (N_19128,N_18780,N_18833);
xnor U19129 (N_19129,N_18829,N_18800);
xnor U19130 (N_19130,N_18949,N_18754);
and U19131 (N_19131,N_18995,N_18854);
and U19132 (N_19132,N_18925,N_18891);
or U19133 (N_19133,N_18927,N_18964);
and U19134 (N_19134,N_18881,N_18884);
or U19135 (N_19135,N_18903,N_18759);
and U19136 (N_19136,N_18924,N_18993);
and U19137 (N_19137,N_18888,N_18976);
nor U19138 (N_19138,N_18947,N_18844);
nand U19139 (N_19139,N_18911,N_18826);
xnor U19140 (N_19140,N_18856,N_18839);
and U19141 (N_19141,N_18884,N_18784);
nand U19142 (N_19142,N_18763,N_18943);
or U19143 (N_19143,N_18945,N_18883);
nand U19144 (N_19144,N_18883,N_18848);
and U19145 (N_19145,N_18839,N_18995);
or U19146 (N_19146,N_18831,N_18886);
nor U19147 (N_19147,N_18756,N_18754);
xnor U19148 (N_19148,N_18816,N_18791);
and U19149 (N_19149,N_18963,N_18822);
nor U19150 (N_19150,N_18963,N_18939);
and U19151 (N_19151,N_18866,N_18981);
nor U19152 (N_19152,N_18857,N_18941);
or U19153 (N_19153,N_18872,N_18804);
or U19154 (N_19154,N_18947,N_18789);
xnor U19155 (N_19155,N_18762,N_18887);
nand U19156 (N_19156,N_18862,N_18770);
and U19157 (N_19157,N_18949,N_18771);
nand U19158 (N_19158,N_18815,N_18970);
xor U19159 (N_19159,N_18891,N_18957);
nor U19160 (N_19160,N_18766,N_18865);
nand U19161 (N_19161,N_18958,N_18970);
xnor U19162 (N_19162,N_18838,N_18937);
xor U19163 (N_19163,N_18772,N_18935);
xor U19164 (N_19164,N_18990,N_18847);
or U19165 (N_19165,N_18830,N_18940);
and U19166 (N_19166,N_18806,N_18946);
nor U19167 (N_19167,N_18993,N_18933);
nand U19168 (N_19168,N_18932,N_18918);
and U19169 (N_19169,N_18890,N_18953);
nor U19170 (N_19170,N_18760,N_18918);
nor U19171 (N_19171,N_18812,N_18926);
xor U19172 (N_19172,N_18833,N_18843);
nand U19173 (N_19173,N_18980,N_18760);
xnor U19174 (N_19174,N_18807,N_18823);
and U19175 (N_19175,N_18805,N_18844);
nor U19176 (N_19176,N_18874,N_18808);
xnor U19177 (N_19177,N_18842,N_18855);
nand U19178 (N_19178,N_18890,N_18829);
and U19179 (N_19179,N_18927,N_18827);
and U19180 (N_19180,N_18841,N_18907);
nor U19181 (N_19181,N_18946,N_18900);
xnor U19182 (N_19182,N_18775,N_18964);
and U19183 (N_19183,N_18836,N_18852);
xnor U19184 (N_19184,N_18883,N_18969);
or U19185 (N_19185,N_18825,N_18886);
or U19186 (N_19186,N_18947,N_18965);
nand U19187 (N_19187,N_18883,N_18801);
nand U19188 (N_19188,N_18817,N_18859);
and U19189 (N_19189,N_18794,N_18948);
and U19190 (N_19190,N_18964,N_18776);
or U19191 (N_19191,N_18814,N_18837);
nand U19192 (N_19192,N_18906,N_18854);
nor U19193 (N_19193,N_18882,N_18842);
and U19194 (N_19194,N_18976,N_18947);
and U19195 (N_19195,N_18890,N_18892);
nor U19196 (N_19196,N_18816,N_18826);
or U19197 (N_19197,N_18788,N_18815);
and U19198 (N_19198,N_18806,N_18850);
and U19199 (N_19199,N_18969,N_18790);
and U19200 (N_19200,N_18956,N_18826);
or U19201 (N_19201,N_18808,N_18915);
nor U19202 (N_19202,N_18999,N_18882);
and U19203 (N_19203,N_18912,N_18956);
or U19204 (N_19204,N_18936,N_18993);
and U19205 (N_19205,N_18886,N_18873);
and U19206 (N_19206,N_18929,N_18841);
xor U19207 (N_19207,N_18820,N_18893);
and U19208 (N_19208,N_18954,N_18938);
or U19209 (N_19209,N_18934,N_18755);
nand U19210 (N_19210,N_18997,N_18808);
xnor U19211 (N_19211,N_18849,N_18825);
and U19212 (N_19212,N_18997,N_18835);
xor U19213 (N_19213,N_18814,N_18809);
nor U19214 (N_19214,N_18754,N_18761);
nand U19215 (N_19215,N_18982,N_18863);
and U19216 (N_19216,N_18913,N_18898);
and U19217 (N_19217,N_18860,N_18795);
nor U19218 (N_19218,N_18902,N_18789);
xnor U19219 (N_19219,N_18915,N_18895);
and U19220 (N_19220,N_18891,N_18852);
or U19221 (N_19221,N_18849,N_18856);
and U19222 (N_19222,N_18901,N_18795);
and U19223 (N_19223,N_18999,N_18913);
xor U19224 (N_19224,N_18814,N_18845);
and U19225 (N_19225,N_18932,N_18877);
or U19226 (N_19226,N_18785,N_18963);
nand U19227 (N_19227,N_18915,N_18771);
nand U19228 (N_19228,N_18939,N_18787);
nand U19229 (N_19229,N_18765,N_18831);
nor U19230 (N_19230,N_18775,N_18761);
nand U19231 (N_19231,N_18768,N_18902);
and U19232 (N_19232,N_18792,N_18856);
and U19233 (N_19233,N_18971,N_18952);
xor U19234 (N_19234,N_18814,N_18938);
xnor U19235 (N_19235,N_18809,N_18928);
nand U19236 (N_19236,N_18935,N_18917);
or U19237 (N_19237,N_18904,N_18752);
and U19238 (N_19238,N_18870,N_18958);
xor U19239 (N_19239,N_18805,N_18969);
or U19240 (N_19240,N_18880,N_18847);
or U19241 (N_19241,N_18966,N_18772);
xnor U19242 (N_19242,N_18760,N_18762);
nand U19243 (N_19243,N_18907,N_18953);
and U19244 (N_19244,N_18807,N_18819);
nor U19245 (N_19245,N_18936,N_18797);
and U19246 (N_19246,N_18943,N_18917);
or U19247 (N_19247,N_18794,N_18912);
or U19248 (N_19248,N_18809,N_18825);
or U19249 (N_19249,N_18828,N_18819);
and U19250 (N_19250,N_19061,N_19190);
xnor U19251 (N_19251,N_19134,N_19112);
or U19252 (N_19252,N_19045,N_19060);
or U19253 (N_19253,N_19221,N_19063);
nand U19254 (N_19254,N_19176,N_19021);
or U19255 (N_19255,N_19120,N_19095);
xnor U19256 (N_19256,N_19144,N_19121);
nor U19257 (N_19257,N_19042,N_19213);
nand U19258 (N_19258,N_19037,N_19018);
or U19259 (N_19259,N_19089,N_19030);
nand U19260 (N_19260,N_19065,N_19180);
xnor U19261 (N_19261,N_19109,N_19117);
nand U19262 (N_19262,N_19192,N_19249);
and U19263 (N_19263,N_19047,N_19188);
or U19264 (N_19264,N_19223,N_19187);
nand U19265 (N_19265,N_19158,N_19022);
nor U19266 (N_19266,N_19220,N_19104);
or U19267 (N_19267,N_19165,N_19012);
xor U19268 (N_19268,N_19010,N_19092);
and U19269 (N_19269,N_19205,N_19241);
nor U19270 (N_19270,N_19210,N_19247);
nor U19271 (N_19271,N_19074,N_19027);
and U19272 (N_19272,N_19067,N_19206);
nand U19273 (N_19273,N_19224,N_19195);
or U19274 (N_19274,N_19020,N_19240);
nor U19275 (N_19275,N_19024,N_19154);
nor U19276 (N_19276,N_19172,N_19142);
or U19277 (N_19277,N_19098,N_19203);
nand U19278 (N_19278,N_19183,N_19186);
xor U19279 (N_19279,N_19185,N_19100);
nor U19280 (N_19280,N_19141,N_19001);
nor U19281 (N_19281,N_19118,N_19152);
or U19282 (N_19282,N_19034,N_19028);
and U19283 (N_19283,N_19171,N_19078);
nand U19284 (N_19284,N_19058,N_19036);
nor U19285 (N_19285,N_19127,N_19248);
nand U19286 (N_19286,N_19115,N_19227);
or U19287 (N_19287,N_19218,N_19236);
nand U19288 (N_19288,N_19135,N_19105);
xor U19289 (N_19289,N_19107,N_19108);
and U19290 (N_19290,N_19164,N_19099);
or U19291 (N_19291,N_19040,N_19149);
and U19292 (N_19292,N_19069,N_19169);
and U19293 (N_19293,N_19184,N_19177);
xor U19294 (N_19294,N_19246,N_19151);
and U19295 (N_19295,N_19200,N_19070);
or U19296 (N_19296,N_19032,N_19029);
or U19297 (N_19297,N_19160,N_19179);
nor U19298 (N_19298,N_19055,N_19011);
or U19299 (N_19299,N_19243,N_19101);
or U19300 (N_19300,N_19096,N_19130);
xnor U19301 (N_19301,N_19191,N_19103);
xor U19302 (N_19302,N_19041,N_19097);
xnor U19303 (N_19303,N_19052,N_19202);
or U19304 (N_19304,N_19170,N_19138);
nor U19305 (N_19305,N_19093,N_19082);
xor U19306 (N_19306,N_19166,N_19150);
nand U19307 (N_19307,N_19016,N_19133);
nand U19308 (N_19308,N_19219,N_19031);
xnor U19309 (N_19309,N_19145,N_19194);
and U19310 (N_19310,N_19015,N_19126);
xnor U19311 (N_19311,N_19214,N_19173);
and U19312 (N_19312,N_19242,N_19085);
nor U19313 (N_19313,N_19043,N_19196);
or U19314 (N_19314,N_19232,N_19147);
and U19315 (N_19315,N_19075,N_19000);
xor U19316 (N_19316,N_19209,N_19178);
nand U19317 (N_19317,N_19228,N_19233);
or U19318 (N_19318,N_19086,N_19009);
nor U19319 (N_19319,N_19129,N_19122);
and U19320 (N_19320,N_19159,N_19123);
or U19321 (N_19321,N_19182,N_19056);
and U19322 (N_19322,N_19080,N_19163);
nand U19323 (N_19323,N_19051,N_19136);
and U19324 (N_19324,N_19155,N_19013);
nand U19325 (N_19325,N_19064,N_19161);
or U19326 (N_19326,N_19002,N_19119);
nand U19327 (N_19327,N_19077,N_19019);
or U19328 (N_19328,N_19057,N_19201);
nand U19329 (N_19329,N_19197,N_19167);
and U19330 (N_19330,N_19072,N_19068);
nor U19331 (N_19331,N_19017,N_19153);
nor U19332 (N_19332,N_19083,N_19076);
nor U19333 (N_19333,N_19087,N_19157);
nand U19334 (N_19334,N_19073,N_19198);
nand U19335 (N_19335,N_19225,N_19212);
or U19336 (N_19336,N_19050,N_19181);
nor U19337 (N_19337,N_19162,N_19059);
nor U19338 (N_19338,N_19023,N_19237);
nor U19339 (N_19339,N_19189,N_19007);
nand U19340 (N_19340,N_19046,N_19084);
nor U19341 (N_19341,N_19208,N_19156);
or U19342 (N_19342,N_19140,N_19091);
or U19343 (N_19343,N_19204,N_19038);
and U19344 (N_19344,N_19148,N_19199);
nand U19345 (N_19345,N_19005,N_19207);
nand U19346 (N_19346,N_19143,N_19244);
xor U19347 (N_19347,N_19215,N_19131);
or U19348 (N_19348,N_19216,N_19039);
nor U19349 (N_19349,N_19239,N_19044);
nor U19350 (N_19350,N_19125,N_19245);
or U19351 (N_19351,N_19222,N_19193);
nand U19352 (N_19352,N_19175,N_19231);
or U19353 (N_19353,N_19116,N_19106);
nor U19354 (N_19354,N_19229,N_19111);
and U19355 (N_19355,N_19062,N_19234);
and U19356 (N_19356,N_19025,N_19014);
and U19357 (N_19357,N_19008,N_19071);
nand U19358 (N_19358,N_19128,N_19139);
xnor U19359 (N_19359,N_19217,N_19003);
nand U19360 (N_19360,N_19110,N_19235);
xor U19361 (N_19361,N_19035,N_19090);
or U19362 (N_19362,N_19174,N_19168);
nor U19363 (N_19363,N_19088,N_19114);
or U19364 (N_19364,N_19102,N_19054);
and U19365 (N_19365,N_19048,N_19079);
and U19366 (N_19366,N_19004,N_19124);
or U19367 (N_19367,N_19137,N_19066);
xor U19368 (N_19368,N_19026,N_19049);
xnor U19369 (N_19369,N_19113,N_19132);
xor U19370 (N_19370,N_19033,N_19094);
nand U19371 (N_19371,N_19006,N_19211);
xnor U19372 (N_19372,N_19053,N_19230);
nor U19373 (N_19373,N_19081,N_19146);
and U19374 (N_19374,N_19238,N_19226);
nor U19375 (N_19375,N_19075,N_19241);
nand U19376 (N_19376,N_19144,N_19201);
or U19377 (N_19377,N_19244,N_19196);
nand U19378 (N_19378,N_19032,N_19098);
nor U19379 (N_19379,N_19101,N_19018);
and U19380 (N_19380,N_19178,N_19154);
nor U19381 (N_19381,N_19044,N_19113);
nor U19382 (N_19382,N_19220,N_19208);
xor U19383 (N_19383,N_19234,N_19219);
nand U19384 (N_19384,N_19052,N_19024);
nor U19385 (N_19385,N_19006,N_19029);
nand U19386 (N_19386,N_19007,N_19160);
xor U19387 (N_19387,N_19205,N_19101);
or U19388 (N_19388,N_19126,N_19241);
nor U19389 (N_19389,N_19011,N_19014);
or U19390 (N_19390,N_19068,N_19157);
xor U19391 (N_19391,N_19203,N_19015);
and U19392 (N_19392,N_19249,N_19048);
nor U19393 (N_19393,N_19116,N_19136);
or U19394 (N_19394,N_19215,N_19160);
nor U19395 (N_19395,N_19206,N_19216);
or U19396 (N_19396,N_19230,N_19249);
nor U19397 (N_19397,N_19111,N_19191);
and U19398 (N_19398,N_19175,N_19123);
nor U19399 (N_19399,N_19032,N_19223);
nand U19400 (N_19400,N_19068,N_19159);
nor U19401 (N_19401,N_19196,N_19079);
or U19402 (N_19402,N_19243,N_19064);
and U19403 (N_19403,N_19007,N_19135);
nand U19404 (N_19404,N_19214,N_19107);
or U19405 (N_19405,N_19098,N_19061);
nand U19406 (N_19406,N_19188,N_19143);
xnor U19407 (N_19407,N_19142,N_19162);
and U19408 (N_19408,N_19191,N_19199);
xnor U19409 (N_19409,N_19014,N_19195);
nor U19410 (N_19410,N_19231,N_19068);
xnor U19411 (N_19411,N_19209,N_19131);
and U19412 (N_19412,N_19016,N_19242);
xor U19413 (N_19413,N_19072,N_19125);
xnor U19414 (N_19414,N_19161,N_19200);
nand U19415 (N_19415,N_19100,N_19196);
nor U19416 (N_19416,N_19056,N_19174);
nand U19417 (N_19417,N_19219,N_19067);
xnor U19418 (N_19418,N_19082,N_19008);
or U19419 (N_19419,N_19212,N_19104);
or U19420 (N_19420,N_19083,N_19242);
or U19421 (N_19421,N_19202,N_19175);
or U19422 (N_19422,N_19067,N_19193);
nand U19423 (N_19423,N_19161,N_19193);
nand U19424 (N_19424,N_19164,N_19016);
or U19425 (N_19425,N_19197,N_19004);
and U19426 (N_19426,N_19094,N_19072);
nand U19427 (N_19427,N_19222,N_19051);
and U19428 (N_19428,N_19039,N_19104);
nor U19429 (N_19429,N_19236,N_19009);
or U19430 (N_19430,N_19171,N_19155);
xor U19431 (N_19431,N_19231,N_19097);
xor U19432 (N_19432,N_19238,N_19063);
and U19433 (N_19433,N_19083,N_19072);
and U19434 (N_19434,N_19225,N_19050);
xnor U19435 (N_19435,N_19139,N_19201);
or U19436 (N_19436,N_19031,N_19059);
nand U19437 (N_19437,N_19247,N_19083);
xor U19438 (N_19438,N_19109,N_19018);
or U19439 (N_19439,N_19172,N_19156);
or U19440 (N_19440,N_19075,N_19247);
or U19441 (N_19441,N_19023,N_19026);
xnor U19442 (N_19442,N_19208,N_19036);
xnor U19443 (N_19443,N_19175,N_19154);
nor U19444 (N_19444,N_19066,N_19016);
and U19445 (N_19445,N_19024,N_19192);
and U19446 (N_19446,N_19210,N_19057);
and U19447 (N_19447,N_19020,N_19201);
nor U19448 (N_19448,N_19122,N_19225);
nand U19449 (N_19449,N_19067,N_19209);
xnor U19450 (N_19450,N_19123,N_19125);
nor U19451 (N_19451,N_19217,N_19093);
nand U19452 (N_19452,N_19114,N_19148);
xnor U19453 (N_19453,N_19194,N_19173);
nand U19454 (N_19454,N_19193,N_19170);
xnor U19455 (N_19455,N_19037,N_19104);
nor U19456 (N_19456,N_19113,N_19243);
nor U19457 (N_19457,N_19028,N_19087);
nand U19458 (N_19458,N_19139,N_19229);
xnor U19459 (N_19459,N_19123,N_19191);
nand U19460 (N_19460,N_19168,N_19160);
nand U19461 (N_19461,N_19220,N_19235);
and U19462 (N_19462,N_19158,N_19036);
xnor U19463 (N_19463,N_19182,N_19193);
and U19464 (N_19464,N_19037,N_19186);
xor U19465 (N_19465,N_19053,N_19096);
nor U19466 (N_19466,N_19008,N_19040);
or U19467 (N_19467,N_19079,N_19237);
nand U19468 (N_19468,N_19181,N_19124);
or U19469 (N_19469,N_19221,N_19163);
and U19470 (N_19470,N_19193,N_19052);
and U19471 (N_19471,N_19140,N_19038);
xnor U19472 (N_19472,N_19068,N_19062);
or U19473 (N_19473,N_19217,N_19086);
nor U19474 (N_19474,N_19148,N_19038);
nor U19475 (N_19475,N_19201,N_19060);
or U19476 (N_19476,N_19037,N_19039);
and U19477 (N_19477,N_19221,N_19238);
xor U19478 (N_19478,N_19194,N_19066);
nor U19479 (N_19479,N_19007,N_19228);
nand U19480 (N_19480,N_19200,N_19189);
and U19481 (N_19481,N_19016,N_19214);
and U19482 (N_19482,N_19037,N_19068);
and U19483 (N_19483,N_19202,N_19130);
nor U19484 (N_19484,N_19144,N_19073);
xnor U19485 (N_19485,N_19167,N_19119);
or U19486 (N_19486,N_19200,N_19172);
xnor U19487 (N_19487,N_19160,N_19082);
xnor U19488 (N_19488,N_19066,N_19139);
nand U19489 (N_19489,N_19015,N_19248);
nand U19490 (N_19490,N_19120,N_19180);
nand U19491 (N_19491,N_19126,N_19176);
or U19492 (N_19492,N_19089,N_19110);
nor U19493 (N_19493,N_19044,N_19227);
nand U19494 (N_19494,N_19083,N_19170);
nor U19495 (N_19495,N_19046,N_19228);
and U19496 (N_19496,N_19037,N_19093);
or U19497 (N_19497,N_19044,N_19006);
nor U19498 (N_19498,N_19049,N_19240);
nand U19499 (N_19499,N_19168,N_19246);
and U19500 (N_19500,N_19419,N_19470);
nand U19501 (N_19501,N_19463,N_19365);
xnor U19502 (N_19502,N_19412,N_19439);
xor U19503 (N_19503,N_19332,N_19388);
nor U19504 (N_19504,N_19459,N_19280);
xor U19505 (N_19505,N_19417,N_19333);
and U19506 (N_19506,N_19448,N_19485);
nor U19507 (N_19507,N_19473,N_19305);
nor U19508 (N_19508,N_19454,N_19442);
nor U19509 (N_19509,N_19284,N_19398);
xor U19510 (N_19510,N_19287,N_19447);
nor U19511 (N_19511,N_19471,N_19432);
and U19512 (N_19512,N_19299,N_19352);
xnor U19513 (N_19513,N_19272,N_19358);
or U19514 (N_19514,N_19295,N_19413);
or U19515 (N_19515,N_19257,N_19356);
nand U19516 (N_19516,N_19343,N_19478);
nand U19517 (N_19517,N_19393,N_19495);
xnor U19518 (N_19518,N_19452,N_19251);
nor U19519 (N_19519,N_19335,N_19405);
nand U19520 (N_19520,N_19488,N_19306);
nand U19521 (N_19521,N_19318,N_19274);
xor U19522 (N_19522,N_19347,N_19465);
or U19523 (N_19523,N_19386,N_19469);
or U19524 (N_19524,N_19291,N_19409);
or U19525 (N_19525,N_19346,N_19453);
or U19526 (N_19526,N_19309,N_19256);
nand U19527 (N_19527,N_19373,N_19403);
xor U19528 (N_19528,N_19354,N_19360);
and U19529 (N_19529,N_19314,N_19323);
xnor U19530 (N_19530,N_19428,N_19285);
and U19531 (N_19531,N_19408,N_19477);
xor U19532 (N_19532,N_19279,N_19391);
nand U19533 (N_19533,N_19493,N_19292);
nand U19534 (N_19534,N_19445,N_19311);
or U19535 (N_19535,N_19400,N_19407);
xnor U19536 (N_19536,N_19380,N_19293);
and U19537 (N_19537,N_19484,N_19384);
nor U19538 (N_19538,N_19476,N_19336);
nor U19539 (N_19539,N_19344,N_19423);
or U19540 (N_19540,N_19374,N_19298);
xor U19541 (N_19541,N_19422,N_19331);
xor U19542 (N_19542,N_19414,N_19369);
xor U19543 (N_19543,N_19371,N_19322);
or U19544 (N_19544,N_19366,N_19316);
nand U19545 (N_19545,N_19479,N_19313);
nand U19546 (N_19546,N_19330,N_19431);
xor U19547 (N_19547,N_19328,N_19253);
nand U19548 (N_19548,N_19261,N_19361);
xor U19549 (N_19549,N_19351,N_19434);
and U19550 (N_19550,N_19399,N_19321);
xnor U19551 (N_19551,N_19466,N_19348);
xor U19552 (N_19552,N_19427,N_19483);
nand U19553 (N_19553,N_19278,N_19326);
nand U19554 (N_19554,N_19372,N_19353);
xor U19555 (N_19555,N_19269,N_19387);
nand U19556 (N_19556,N_19468,N_19266);
xor U19557 (N_19557,N_19276,N_19464);
or U19558 (N_19558,N_19416,N_19490);
or U19559 (N_19559,N_19449,N_19341);
nor U19560 (N_19560,N_19397,N_19320);
and U19561 (N_19561,N_19492,N_19268);
nor U19562 (N_19562,N_19482,N_19264);
and U19563 (N_19563,N_19345,N_19496);
nor U19564 (N_19564,N_19433,N_19286);
xnor U19565 (N_19565,N_19392,N_19355);
nor U19566 (N_19566,N_19282,N_19429);
and U19567 (N_19567,N_19404,N_19455);
or U19568 (N_19568,N_19467,N_19340);
nor U19569 (N_19569,N_19270,N_19451);
nor U19570 (N_19570,N_19390,N_19273);
or U19571 (N_19571,N_19440,N_19494);
nand U19572 (N_19572,N_19489,N_19394);
xor U19573 (N_19573,N_19438,N_19277);
xnor U19574 (N_19574,N_19255,N_19363);
nand U19575 (N_19575,N_19370,N_19375);
or U19576 (N_19576,N_19420,N_19324);
and U19577 (N_19577,N_19315,N_19379);
nor U19578 (N_19578,N_19342,N_19406);
nand U19579 (N_19579,N_19436,N_19462);
nand U19580 (N_19580,N_19319,N_19294);
or U19581 (N_19581,N_19385,N_19258);
nand U19582 (N_19582,N_19444,N_19259);
nor U19583 (N_19583,N_19317,N_19446);
and U19584 (N_19584,N_19304,N_19443);
and U19585 (N_19585,N_19300,N_19497);
and U19586 (N_19586,N_19437,N_19458);
or U19587 (N_19587,N_19302,N_19418);
xor U19588 (N_19588,N_19325,N_19396);
or U19589 (N_19589,N_19275,N_19262);
nand U19590 (N_19590,N_19383,N_19450);
nor U19591 (N_19591,N_19389,N_19308);
or U19592 (N_19592,N_19424,N_19378);
xor U19593 (N_19593,N_19368,N_19426);
xnor U19594 (N_19594,N_19441,N_19338);
and U19595 (N_19595,N_19339,N_19395);
nand U19596 (N_19596,N_19312,N_19349);
nor U19597 (N_19597,N_19254,N_19410);
nand U19598 (N_19598,N_19472,N_19475);
or U19599 (N_19599,N_19480,N_19283);
or U19600 (N_19600,N_19435,N_19487);
xor U19601 (N_19601,N_19260,N_19461);
or U19602 (N_19602,N_19290,N_19364);
nand U19603 (N_19603,N_19271,N_19252);
nor U19604 (N_19604,N_19281,N_19474);
nor U19605 (N_19605,N_19498,N_19288);
nor U19606 (N_19606,N_19289,N_19421);
nor U19607 (N_19607,N_19402,N_19296);
nand U19608 (N_19608,N_19297,N_19415);
nor U19609 (N_19609,N_19382,N_19357);
xnor U19610 (N_19610,N_19303,N_19430);
and U19611 (N_19611,N_19381,N_19499);
nand U19612 (N_19612,N_19367,N_19359);
xor U19613 (N_19613,N_19362,N_19265);
and U19614 (N_19614,N_19486,N_19460);
nand U19615 (N_19615,N_19411,N_19337);
xor U19616 (N_19616,N_19334,N_19377);
and U19617 (N_19617,N_19481,N_19456);
and U19618 (N_19618,N_19327,N_19376);
nand U19619 (N_19619,N_19491,N_19263);
nor U19620 (N_19620,N_19267,N_19307);
xor U19621 (N_19621,N_19401,N_19425);
or U19622 (N_19622,N_19350,N_19457);
xor U19623 (N_19623,N_19250,N_19310);
nor U19624 (N_19624,N_19329,N_19301);
or U19625 (N_19625,N_19259,N_19337);
and U19626 (N_19626,N_19472,N_19326);
and U19627 (N_19627,N_19263,N_19325);
nor U19628 (N_19628,N_19466,N_19477);
and U19629 (N_19629,N_19345,N_19309);
or U19630 (N_19630,N_19350,N_19451);
and U19631 (N_19631,N_19404,N_19255);
and U19632 (N_19632,N_19392,N_19431);
and U19633 (N_19633,N_19265,N_19278);
and U19634 (N_19634,N_19454,N_19382);
or U19635 (N_19635,N_19294,N_19329);
xor U19636 (N_19636,N_19460,N_19334);
and U19637 (N_19637,N_19310,N_19257);
xnor U19638 (N_19638,N_19393,N_19397);
or U19639 (N_19639,N_19488,N_19256);
nand U19640 (N_19640,N_19331,N_19343);
xnor U19641 (N_19641,N_19437,N_19314);
nand U19642 (N_19642,N_19431,N_19398);
or U19643 (N_19643,N_19271,N_19436);
and U19644 (N_19644,N_19470,N_19445);
or U19645 (N_19645,N_19449,N_19279);
and U19646 (N_19646,N_19379,N_19341);
xor U19647 (N_19647,N_19333,N_19419);
nand U19648 (N_19648,N_19292,N_19384);
xnor U19649 (N_19649,N_19432,N_19416);
xnor U19650 (N_19650,N_19495,N_19259);
nand U19651 (N_19651,N_19387,N_19303);
xnor U19652 (N_19652,N_19493,N_19485);
xnor U19653 (N_19653,N_19472,N_19272);
xor U19654 (N_19654,N_19320,N_19290);
xnor U19655 (N_19655,N_19386,N_19485);
xnor U19656 (N_19656,N_19319,N_19419);
xor U19657 (N_19657,N_19266,N_19285);
nor U19658 (N_19658,N_19367,N_19408);
or U19659 (N_19659,N_19444,N_19446);
xnor U19660 (N_19660,N_19259,N_19334);
and U19661 (N_19661,N_19319,N_19395);
and U19662 (N_19662,N_19346,N_19471);
and U19663 (N_19663,N_19325,N_19333);
nand U19664 (N_19664,N_19369,N_19264);
nand U19665 (N_19665,N_19284,N_19300);
xor U19666 (N_19666,N_19261,N_19350);
and U19667 (N_19667,N_19364,N_19347);
nand U19668 (N_19668,N_19476,N_19333);
nand U19669 (N_19669,N_19487,N_19460);
nand U19670 (N_19670,N_19313,N_19391);
or U19671 (N_19671,N_19458,N_19255);
nor U19672 (N_19672,N_19327,N_19488);
and U19673 (N_19673,N_19282,N_19411);
nand U19674 (N_19674,N_19391,N_19303);
or U19675 (N_19675,N_19326,N_19443);
xor U19676 (N_19676,N_19411,N_19343);
xor U19677 (N_19677,N_19401,N_19342);
xor U19678 (N_19678,N_19381,N_19352);
nor U19679 (N_19679,N_19440,N_19258);
and U19680 (N_19680,N_19317,N_19403);
nor U19681 (N_19681,N_19489,N_19429);
and U19682 (N_19682,N_19285,N_19299);
nor U19683 (N_19683,N_19406,N_19295);
nor U19684 (N_19684,N_19281,N_19268);
or U19685 (N_19685,N_19319,N_19329);
or U19686 (N_19686,N_19457,N_19376);
xor U19687 (N_19687,N_19462,N_19258);
or U19688 (N_19688,N_19298,N_19430);
or U19689 (N_19689,N_19287,N_19252);
and U19690 (N_19690,N_19298,N_19378);
xor U19691 (N_19691,N_19394,N_19330);
nor U19692 (N_19692,N_19423,N_19363);
or U19693 (N_19693,N_19337,N_19348);
and U19694 (N_19694,N_19378,N_19490);
and U19695 (N_19695,N_19292,N_19272);
and U19696 (N_19696,N_19341,N_19490);
and U19697 (N_19697,N_19282,N_19345);
nor U19698 (N_19698,N_19304,N_19486);
and U19699 (N_19699,N_19301,N_19462);
and U19700 (N_19700,N_19368,N_19457);
nor U19701 (N_19701,N_19390,N_19361);
or U19702 (N_19702,N_19325,N_19264);
and U19703 (N_19703,N_19453,N_19339);
nand U19704 (N_19704,N_19350,N_19293);
and U19705 (N_19705,N_19312,N_19481);
or U19706 (N_19706,N_19429,N_19338);
nor U19707 (N_19707,N_19476,N_19261);
or U19708 (N_19708,N_19285,N_19350);
nand U19709 (N_19709,N_19277,N_19356);
nand U19710 (N_19710,N_19426,N_19408);
xnor U19711 (N_19711,N_19360,N_19303);
xnor U19712 (N_19712,N_19250,N_19491);
nor U19713 (N_19713,N_19271,N_19317);
or U19714 (N_19714,N_19394,N_19387);
nand U19715 (N_19715,N_19297,N_19354);
and U19716 (N_19716,N_19492,N_19434);
and U19717 (N_19717,N_19272,N_19465);
and U19718 (N_19718,N_19428,N_19348);
xor U19719 (N_19719,N_19413,N_19278);
nand U19720 (N_19720,N_19360,N_19446);
or U19721 (N_19721,N_19391,N_19381);
nand U19722 (N_19722,N_19422,N_19477);
nand U19723 (N_19723,N_19257,N_19474);
or U19724 (N_19724,N_19488,N_19487);
and U19725 (N_19725,N_19400,N_19314);
nor U19726 (N_19726,N_19413,N_19484);
nand U19727 (N_19727,N_19335,N_19364);
xor U19728 (N_19728,N_19480,N_19468);
nor U19729 (N_19729,N_19455,N_19342);
xor U19730 (N_19730,N_19464,N_19318);
nor U19731 (N_19731,N_19388,N_19429);
or U19732 (N_19732,N_19355,N_19301);
xnor U19733 (N_19733,N_19307,N_19470);
nor U19734 (N_19734,N_19322,N_19495);
xnor U19735 (N_19735,N_19461,N_19426);
or U19736 (N_19736,N_19383,N_19346);
nor U19737 (N_19737,N_19269,N_19380);
nor U19738 (N_19738,N_19287,N_19250);
nand U19739 (N_19739,N_19282,N_19432);
nand U19740 (N_19740,N_19472,N_19484);
xnor U19741 (N_19741,N_19314,N_19353);
or U19742 (N_19742,N_19433,N_19492);
nor U19743 (N_19743,N_19422,N_19256);
nor U19744 (N_19744,N_19343,N_19424);
xnor U19745 (N_19745,N_19346,N_19460);
nand U19746 (N_19746,N_19286,N_19493);
nand U19747 (N_19747,N_19457,N_19355);
or U19748 (N_19748,N_19345,N_19420);
xor U19749 (N_19749,N_19317,N_19430);
nor U19750 (N_19750,N_19530,N_19680);
xor U19751 (N_19751,N_19699,N_19591);
nor U19752 (N_19752,N_19713,N_19595);
or U19753 (N_19753,N_19665,N_19717);
or U19754 (N_19754,N_19513,N_19674);
nand U19755 (N_19755,N_19536,N_19597);
and U19756 (N_19756,N_19650,N_19686);
or U19757 (N_19757,N_19669,N_19567);
nor U19758 (N_19758,N_19635,N_19577);
or U19759 (N_19759,N_19640,N_19537);
or U19760 (N_19760,N_19731,N_19552);
nor U19761 (N_19761,N_19644,N_19582);
nor U19762 (N_19762,N_19570,N_19627);
and U19763 (N_19763,N_19676,N_19526);
nand U19764 (N_19764,N_19589,N_19726);
nor U19765 (N_19765,N_19578,N_19512);
or U19766 (N_19766,N_19656,N_19572);
xnor U19767 (N_19767,N_19535,N_19606);
nand U19768 (N_19768,N_19617,N_19651);
or U19769 (N_19769,N_19706,N_19690);
xor U19770 (N_19770,N_19695,N_19707);
or U19771 (N_19771,N_19613,N_19603);
and U19772 (N_19772,N_19648,N_19594);
nor U19773 (N_19773,N_19500,N_19637);
nor U19774 (N_19774,N_19716,N_19510);
and U19775 (N_19775,N_19704,N_19660);
xor U19776 (N_19776,N_19691,N_19612);
nand U19777 (N_19777,N_19569,N_19505);
and U19778 (N_19778,N_19715,N_19621);
and U19779 (N_19779,N_19508,N_19700);
nor U19780 (N_19780,N_19598,N_19571);
and U19781 (N_19781,N_19659,N_19681);
xnor U19782 (N_19782,N_19502,N_19693);
nand U19783 (N_19783,N_19729,N_19639);
nor U19784 (N_19784,N_19596,N_19657);
xnor U19785 (N_19785,N_19531,N_19679);
or U19786 (N_19786,N_19645,N_19517);
nand U19787 (N_19787,N_19583,N_19702);
or U19788 (N_19788,N_19661,N_19554);
and U19789 (N_19789,N_19566,N_19641);
or U19790 (N_19790,N_19728,N_19633);
xor U19791 (N_19791,N_19742,N_19559);
nor U19792 (N_19792,N_19576,N_19564);
and U19793 (N_19793,N_19671,N_19685);
nand U19794 (N_19794,N_19615,N_19556);
nor U19795 (N_19795,N_19545,N_19522);
xor U19796 (N_19796,N_19732,N_19561);
nor U19797 (N_19797,N_19701,N_19562);
xor U19798 (N_19798,N_19719,N_19548);
nor U19799 (N_19799,N_19740,N_19737);
and U19800 (N_19800,N_19553,N_19692);
xnor U19801 (N_19801,N_19672,N_19609);
nor U19802 (N_19802,N_19724,N_19518);
nor U19803 (N_19803,N_19698,N_19551);
or U19804 (N_19804,N_19525,N_19743);
nand U19805 (N_19805,N_19563,N_19668);
nand U19806 (N_19806,N_19654,N_19614);
nand U19807 (N_19807,N_19574,N_19542);
or U19808 (N_19808,N_19629,N_19540);
or U19809 (N_19809,N_19619,N_19565);
and U19810 (N_19810,N_19528,N_19543);
xor U19811 (N_19811,N_19722,N_19585);
and U19812 (N_19812,N_19688,N_19532);
nand U19813 (N_19813,N_19558,N_19733);
nor U19814 (N_19814,N_19515,N_19611);
nor U19815 (N_19815,N_19549,N_19705);
xnor U19816 (N_19816,N_19523,N_19599);
xnor U19817 (N_19817,N_19642,N_19587);
xor U19818 (N_19818,N_19581,N_19664);
xor U19819 (N_19819,N_19696,N_19634);
xor U19820 (N_19820,N_19623,N_19678);
or U19821 (N_19821,N_19573,N_19745);
xor U19822 (N_19822,N_19618,N_19747);
or U19823 (N_19823,N_19625,N_19703);
or U19824 (N_19824,N_19655,N_19721);
xnor U19825 (N_19825,N_19605,N_19521);
and U19826 (N_19826,N_19519,N_19520);
and U19827 (N_19827,N_19632,N_19744);
nor U19828 (N_19828,N_19602,N_19670);
or U19829 (N_19829,N_19514,N_19636);
nor U19830 (N_19830,N_19620,N_19630);
or U19831 (N_19831,N_19550,N_19601);
or U19832 (N_19832,N_19653,N_19673);
nand U19833 (N_19833,N_19723,N_19643);
and U19834 (N_19834,N_19511,N_19580);
and U19835 (N_19835,N_19711,N_19604);
or U19836 (N_19836,N_19626,N_19662);
nor U19837 (N_19837,N_19516,N_19682);
or U19838 (N_19838,N_19547,N_19507);
or U19839 (N_19839,N_19610,N_19712);
xnor U19840 (N_19840,N_19622,N_19709);
nand U19841 (N_19841,N_19631,N_19718);
or U19842 (N_19842,N_19608,N_19503);
nand U19843 (N_19843,N_19689,N_19663);
nand U19844 (N_19844,N_19730,N_19541);
nand U19845 (N_19845,N_19735,N_19579);
xnor U19846 (N_19846,N_19546,N_19647);
and U19847 (N_19847,N_19720,N_19588);
or U19848 (N_19848,N_19557,N_19533);
xnor U19849 (N_19849,N_19638,N_19593);
nor U19850 (N_19850,N_19649,N_19509);
xor U19851 (N_19851,N_19646,N_19727);
nor U19852 (N_19852,N_19738,N_19616);
xnor U19853 (N_19853,N_19555,N_19584);
xor U19854 (N_19854,N_19624,N_19684);
nor U19855 (N_19855,N_19710,N_19628);
nor U19856 (N_19856,N_19675,N_19734);
nand U19857 (N_19857,N_19600,N_19749);
or U19858 (N_19858,N_19501,N_19736);
and U19859 (N_19859,N_19568,N_19741);
and U19860 (N_19860,N_19607,N_19504);
nor U19861 (N_19861,N_19534,N_19586);
or U19862 (N_19862,N_19506,N_19697);
or U19863 (N_19863,N_19544,N_19590);
nand U19864 (N_19864,N_19539,N_19725);
and U19865 (N_19865,N_19746,N_19748);
nand U19866 (N_19866,N_19667,N_19560);
and U19867 (N_19867,N_19658,N_19575);
nand U19868 (N_19868,N_19666,N_19694);
nand U19869 (N_19869,N_19677,N_19529);
and U19870 (N_19870,N_19527,N_19652);
xnor U19871 (N_19871,N_19714,N_19739);
nand U19872 (N_19872,N_19592,N_19687);
nor U19873 (N_19873,N_19524,N_19683);
nor U19874 (N_19874,N_19538,N_19708);
xnor U19875 (N_19875,N_19535,N_19615);
nor U19876 (N_19876,N_19746,N_19671);
and U19877 (N_19877,N_19502,N_19745);
nand U19878 (N_19878,N_19569,N_19525);
or U19879 (N_19879,N_19563,N_19619);
xnor U19880 (N_19880,N_19700,N_19513);
and U19881 (N_19881,N_19604,N_19578);
and U19882 (N_19882,N_19535,N_19685);
and U19883 (N_19883,N_19570,N_19642);
or U19884 (N_19884,N_19556,N_19594);
xor U19885 (N_19885,N_19640,N_19729);
nor U19886 (N_19886,N_19572,N_19637);
nor U19887 (N_19887,N_19558,N_19608);
nor U19888 (N_19888,N_19671,N_19580);
xor U19889 (N_19889,N_19503,N_19722);
nor U19890 (N_19890,N_19503,N_19716);
nor U19891 (N_19891,N_19589,N_19535);
or U19892 (N_19892,N_19650,N_19511);
nor U19893 (N_19893,N_19719,N_19742);
xor U19894 (N_19894,N_19738,N_19671);
nor U19895 (N_19895,N_19688,N_19704);
xnor U19896 (N_19896,N_19638,N_19689);
or U19897 (N_19897,N_19686,N_19611);
nor U19898 (N_19898,N_19539,N_19573);
or U19899 (N_19899,N_19699,N_19726);
and U19900 (N_19900,N_19711,N_19617);
nand U19901 (N_19901,N_19506,N_19627);
nand U19902 (N_19902,N_19626,N_19681);
or U19903 (N_19903,N_19675,N_19660);
nand U19904 (N_19904,N_19552,N_19532);
nor U19905 (N_19905,N_19605,N_19539);
nand U19906 (N_19906,N_19692,N_19600);
nor U19907 (N_19907,N_19550,N_19638);
and U19908 (N_19908,N_19514,N_19709);
or U19909 (N_19909,N_19717,N_19625);
and U19910 (N_19910,N_19658,N_19661);
nand U19911 (N_19911,N_19698,N_19612);
or U19912 (N_19912,N_19673,N_19666);
and U19913 (N_19913,N_19692,N_19706);
and U19914 (N_19914,N_19502,N_19555);
or U19915 (N_19915,N_19571,N_19696);
or U19916 (N_19916,N_19664,N_19537);
or U19917 (N_19917,N_19532,N_19698);
xor U19918 (N_19918,N_19502,N_19579);
or U19919 (N_19919,N_19634,N_19597);
xor U19920 (N_19920,N_19602,N_19654);
or U19921 (N_19921,N_19748,N_19637);
nand U19922 (N_19922,N_19509,N_19629);
nand U19923 (N_19923,N_19666,N_19728);
nor U19924 (N_19924,N_19572,N_19743);
nor U19925 (N_19925,N_19528,N_19639);
xnor U19926 (N_19926,N_19547,N_19650);
or U19927 (N_19927,N_19651,N_19632);
nor U19928 (N_19928,N_19610,N_19717);
and U19929 (N_19929,N_19660,N_19537);
xnor U19930 (N_19930,N_19742,N_19606);
and U19931 (N_19931,N_19559,N_19675);
nand U19932 (N_19932,N_19680,N_19596);
and U19933 (N_19933,N_19714,N_19518);
nand U19934 (N_19934,N_19520,N_19569);
and U19935 (N_19935,N_19624,N_19645);
or U19936 (N_19936,N_19711,N_19565);
xnor U19937 (N_19937,N_19545,N_19547);
or U19938 (N_19938,N_19574,N_19584);
and U19939 (N_19939,N_19538,N_19711);
or U19940 (N_19940,N_19659,N_19633);
xnor U19941 (N_19941,N_19524,N_19576);
xnor U19942 (N_19942,N_19557,N_19749);
and U19943 (N_19943,N_19533,N_19712);
nor U19944 (N_19944,N_19623,N_19657);
or U19945 (N_19945,N_19629,N_19581);
nand U19946 (N_19946,N_19573,N_19741);
nand U19947 (N_19947,N_19708,N_19533);
nor U19948 (N_19948,N_19578,N_19633);
nand U19949 (N_19949,N_19614,N_19631);
nand U19950 (N_19950,N_19515,N_19740);
and U19951 (N_19951,N_19637,N_19593);
and U19952 (N_19952,N_19738,N_19502);
and U19953 (N_19953,N_19697,N_19715);
nand U19954 (N_19954,N_19564,N_19527);
xor U19955 (N_19955,N_19563,N_19702);
nand U19956 (N_19956,N_19605,N_19739);
xor U19957 (N_19957,N_19545,N_19738);
nor U19958 (N_19958,N_19500,N_19663);
and U19959 (N_19959,N_19678,N_19714);
nor U19960 (N_19960,N_19703,N_19614);
xor U19961 (N_19961,N_19690,N_19632);
nand U19962 (N_19962,N_19692,N_19624);
and U19963 (N_19963,N_19533,N_19580);
xnor U19964 (N_19964,N_19508,N_19704);
xnor U19965 (N_19965,N_19614,N_19638);
nor U19966 (N_19966,N_19727,N_19728);
or U19967 (N_19967,N_19529,N_19613);
nand U19968 (N_19968,N_19625,N_19691);
or U19969 (N_19969,N_19566,N_19634);
or U19970 (N_19970,N_19655,N_19668);
nor U19971 (N_19971,N_19568,N_19575);
and U19972 (N_19972,N_19691,N_19662);
and U19973 (N_19973,N_19664,N_19682);
nand U19974 (N_19974,N_19629,N_19514);
nand U19975 (N_19975,N_19705,N_19529);
or U19976 (N_19976,N_19532,N_19562);
nand U19977 (N_19977,N_19686,N_19541);
or U19978 (N_19978,N_19507,N_19597);
and U19979 (N_19979,N_19578,N_19652);
xnor U19980 (N_19980,N_19692,N_19646);
xor U19981 (N_19981,N_19585,N_19747);
or U19982 (N_19982,N_19744,N_19523);
nand U19983 (N_19983,N_19679,N_19528);
or U19984 (N_19984,N_19684,N_19669);
and U19985 (N_19985,N_19737,N_19612);
nor U19986 (N_19986,N_19611,N_19669);
nand U19987 (N_19987,N_19622,N_19743);
or U19988 (N_19988,N_19623,N_19591);
and U19989 (N_19989,N_19591,N_19596);
nand U19990 (N_19990,N_19725,N_19693);
nand U19991 (N_19991,N_19681,N_19724);
nand U19992 (N_19992,N_19557,N_19689);
xor U19993 (N_19993,N_19553,N_19523);
nand U19994 (N_19994,N_19579,N_19519);
nand U19995 (N_19995,N_19704,N_19687);
and U19996 (N_19996,N_19655,N_19660);
xnor U19997 (N_19997,N_19628,N_19656);
or U19998 (N_19998,N_19580,N_19512);
nor U19999 (N_19999,N_19520,N_19711);
and U20000 (N_20000,N_19848,N_19780);
xnor U20001 (N_20001,N_19979,N_19940);
xnor U20002 (N_20002,N_19958,N_19866);
nor U20003 (N_20003,N_19825,N_19903);
or U20004 (N_20004,N_19778,N_19872);
or U20005 (N_20005,N_19907,N_19967);
nor U20006 (N_20006,N_19857,N_19884);
nand U20007 (N_20007,N_19793,N_19776);
and U20008 (N_20008,N_19901,N_19752);
nand U20009 (N_20009,N_19831,N_19797);
or U20010 (N_20010,N_19948,N_19845);
and U20011 (N_20011,N_19881,N_19791);
or U20012 (N_20012,N_19863,N_19916);
nand U20013 (N_20013,N_19926,N_19993);
nand U20014 (N_20014,N_19782,N_19919);
and U20015 (N_20015,N_19750,N_19813);
or U20016 (N_20016,N_19763,N_19897);
nand U20017 (N_20017,N_19783,N_19998);
nor U20018 (N_20018,N_19837,N_19839);
nor U20019 (N_20019,N_19808,N_19868);
or U20020 (N_20020,N_19854,N_19867);
xor U20021 (N_20021,N_19798,N_19805);
or U20022 (N_20022,N_19879,N_19771);
nand U20023 (N_20023,N_19833,N_19895);
nor U20024 (N_20024,N_19943,N_19761);
nand U20025 (N_20025,N_19883,N_19772);
or U20026 (N_20026,N_19947,N_19836);
and U20027 (N_20027,N_19924,N_19822);
or U20028 (N_20028,N_19835,N_19991);
xor U20029 (N_20029,N_19774,N_19806);
and U20030 (N_20030,N_19978,N_19892);
or U20031 (N_20031,N_19904,N_19952);
or U20032 (N_20032,N_19853,N_19850);
nor U20033 (N_20033,N_19796,N_19869);
xor U20034 (N_20034,N_19803,N_19814);
xnor U20035 (N_20035,N_19859,N_19936);
and U20036 (N_20036,N_19959,N_19939);
and U20037 (N_20037,N_19942,N_19807);
nor U20038 (N_20038,N_19874,N_19912);
or U20039 (N_20039,N_19975,N_19759);
and U20040 (N_20040,N_19760,N_19921);
nand U20041 (N_20041,N_19865,N_19784);
nor U20042 (N_20042,N_19905,N_19891);
nand U20043 (N_20043,N_19846,N_19777);
nor U20044 (N_20044,N_19894,N_19847);
or U20045 (N_20045,N_19974,N_19862);
nor U20046 (N_20046,N_19900,N_19787);
nor U20047 (N_20047,N_19955,N_19932);
or U20048 (N_20048,N_19913,N_19844);
and U20049 (N_20049,N_19789,N_19908);
nor U20050 (N_20050,N_19909,N_19842);
and U20051 (N_20051,N_19937,N_19786);
nor U20052 (N_20052,N_19792,N_19785);
or U20053 (N_20053,N_19911,N_19969);
nand U20054 (N_20054,N_19801,N_19946);
or U20055 (N_20055,N_19804,N_19928);
and U20056 (N_20056,N_19992,N_19963);
and U20057 (N_20057,N_19961,N_19964);
or U20058 (N_20058,N_19826,N_19795);
or U20059 (N_20059,N_19794,N_19945);
xnor U20060 (N_20060,N_19769,N_19953);
or U20061 (N_20061,N_19843,N_19893);
nand U20062 (N_20062,N_19925,N_19820);
and U20063 (N_20063,N_19989,N_19767);
nor U20064 (N_20064,N_19941,N_19968);
nor U20065 (N_20065,N_19887,N_19775);
nand U20066 (N_20066,N_19827,N_19756);
nor U20067 (N_20067,N_19965,N_19758);
nand U20068 (N_20068,N_19849,N_19990);
xnor U20069 (N_20069,N_19930,N_19976);
xnor U20070 (N_20070,N_19927,N_19768);
nand U20071 (N_20071,N_19973,N_19882);
and U20072 (N_20072,N_19950,N_19999);
nor U20073 (N_20073,N_19951,N_19935);
and U20074 (N_20074,N_19815,N_19988);
or U20075 (N_20075,N_19832,N_19773);
and U20076 (N_20076,N_19922,N_19762);
or U20077 (N_20077,N_19915,N_19956);
or U20078 (N_20078,N_19878,N_19987);
nand U20079 (N_20079,N_19982,N_19949);
nand U20080 (N_20080,N_19755,N_19985);
or U20081 (N_20081,N_19817,N_19934);
or U20082 (N_20082,N_19821,N_19823);
nand U20083 (N_20083,N_19754,N_19962);
or U20084 (N_20084,N_19858,N_19864);
and U20085 (N_20085,N_19981,N_19886);
nand U20086 (N_20086,N_19779,N_19944);
xor U20087 (N_20087,N_19824,N_19770);
nor U20088 (N_20088,N_19781,N_19929);
nand U20089 (N_20089,N_19995,N_19880);
xnor U20090 (N_20090,N_19970,N_19855);
and U20091 (N_20091,N_19753,N_19829);
xor U20092 (N_20092,N_19885,N_19828);
nand U20093 (N_20093,N_19876,N_19918);
xnor U20094 (N_20094,N_19984,N_19766);
or U20095 (N_20095,N_19800,N_19898);
and U20096 (N_20096,N_19816,N_19888);
and U20097 (N_20097,N_19861,N_19811);
xor U20098 (N_20098,N_19819,N_19966);
or U20099 (N_20099,N_19852,N_19830);
and U20100 (N_20100,N_19870,N_19960);
xnor U20101 (N_20101,N_19997,N_19764);
nor U20102 (N_20102,N_19931,N_19954);
and U20103 (N_20103,N_19980,N_19938);
and U20104 (N_20104,N_19957,N_19910);
xnor U20105 (N_20105,N_19994,N_19751);
nand U20106 (N_20106,N_19790,N_19838);
nand U20107 (N_20107,N_19877,N_19841);
nor U20108 (N_20108,N_19906,N_19890);
xor U20109 (N_20109,N_19757,N_19986);
nand U20110 (N_20110,N_19902,N_19834);
xnor U20111 (N_20111,N_19809,N_19860);
nand U20112 (N_20112,N_19914,N_19818);
nand U20113 (N_20113,N_19810,N_19873);
and U20114 (N_20114,N_19875,N_19977);
xnor U20115 (N_20115,N_19788,N_19802);
xor U20116 (N_20116,N_19896,N_19851);
nand U20117 (N_20117,N_19917,N_19856);
xnor U20118 (N_20118,N_19972,N_19923);
xnor U20119 (N_20119,N_19871,N_19765);
nor U20120 (N_20120,N_19996,N_19920);
or U20121 (N_20121,N_19983,N_19971);
xnor U20122 (N_20122,N_19812,N_19840);
xnor U20123 (N_20123,N_19899,N_19889);
or U20124 (N_20124,N_19799,N_19933);
or U20125 (N_20125,N_19881,N_19888);
nand U20126 (N_20126,N_19936,N_19860);
and U20127 (N_20127,N_19887,N_19873);
or U20128 (N_20128,N_19924,N_19857);
xor U20129 (N_20129,N_19786,N_19988);
or U20130 (N_20130,N_19769,N_19813);
xnor U20131 (N_20131,N_19776,N_19939);
and U20132 (N_20132,N_19925,N_19833);
and U20133 (N_20133,N_19848,N_19837);
nand U20134 (N_20134,N_19855,N_19937);
xnor U20135 (N_20135,N_19984,N_19755);
and U20136 (N_20136,N_19892,N_19783);
nand U20137 (N_20137,N_19961,N_19902);
or U20138 (N_20138,N_19945,N_19946);
and U20139 (N_20139,N_19875,N_19851);
or U20140 (N_20140,N_19861,N_19792);
or U20141 (N_20141,N_19990,N_19767);
or U20142 (N_20142,N_19944,N_19871);
or U20143 (N_20143,N_19965,N_19775);
or U20144 (N_20144,N_19807,N_19783);
nor U20145 (N_20145,N_19923,N_19784);
nor U20146 (N_20146,N_19776,N_19870);
xnor U20147 (N_20147,N_19816,N_19895);
xor U20148 (N_20148,N_19954,N_19929);
nand U20149 (N_20149,N_19851,N_19887);
xor U20150 (N_20150,N_19840,N_19976);
nand U20151 (N_20151,N_19827,N_19974);
or U20152 (N_20152,N_19881,N_19802);
or U20153 (N_20153,N_19977,N_19944);
xor U20154 (N_20154,N_19873,N_19993);
nand U20155 (N_20155,N_19814,N_19891);
nand U20156 (N_20156,N_19942,N_19751);
or U20157 (N_20157,N_19789,N_19872);
xnor U20158 (N_20158,N_19884,N_19812);
nor U20159 (N_20159,N_19873,N_19998);
nor U20160 (N_20160,N_19806,N_19920);
and U20161 (N_20161,N_19869,N_19890);
and U20162 (N_20162,N_19791,N_19906);
xnor U20163 (N_20163,N_19972,N_19906);
and U20164 (N_20164,N_19972,N_19775);
nor U20165 (N_20165,N_19958,N_19807);
nor U20166 (N_20166,N_19773,N_19988);
nand U20167 (N_20167,N_19811,N_19923);
and U20168 (N_20168,N_19908,N_19940);
nor U20169 (N_20169,N_19990,N_19906);
xnor U20170 (N_20170,N_19897,N_19869);
nand U20171 (N_20171,N_19759,N_19999);
xor U20172 (N_20172,N_19801,N_19840);
xor U20173 (N_20173,N_19825,N_19865);
nand U20174 (N_20174,N_19810,N_19896);
or U20175 (N_20175,N_19776,N_19962);
nand U20176 (N_20176,N_19988,N_19882);
or U20177 (N_20177,N_19887,N_19876);
or U20178 (N_20178,N_19848,N_19859);
xnor U20179 (N_20179,N_19771,N_19868);
and U20180 (N_20180,N_19817,N_19750);
and U20181 (N_20181,N_19905,N_19963);
or U20182 (N_20182,N_19822,N_19956);
nand U20183 (N_20183,N_19921,N_19893);
xnor U20184 (N_20184,N_19841,N_19932);
and U20185 (N_20185,N_19833,N_19945);
or U20186 (N_20186,N_19948,N_19912);
or U20187 (N_20187,N_19929,N_19848);
and U20188 (N_20188,N_19889,N_19773);
nand U20189 (N_20189,N_19911,N_19800);
and U20190 (N_20190,N_19841,N_19871);
nor U20191 (N_20191,N_19972,N_19990);
nor U20192 (N_20192,N_19940,N_19883);
and U20193 (N_20193,N_19934,N_19873);
xor U20194 (N_20194,N_19929,N_19888);
nand U20195 (N_20195,N_19973,N_19955);
or U20196 (N_20196,N_19759,N_19858);
or U20197 (N_20197,N_19812,N_19876);
nor U20198 (N_20198,N_19953,N_19879);
or U20199 (N_20199,N_19882,N_19757);
xor U20200 (N_20200,N_19895,N_19785);
nor U20201 (N_20201,N_19823,N_19898);
nand U20202 (N_20202,N_19926,N_19789);
or U20203 (N_20203,N_19861,N_19976);
and U20204 (N_20204,N_19954,N_19814);
nand U20205 (N_20205,N_19836,N_19873);
xor U20206 (N_20206,N_19756,N_19906);
xor U20207 (N_20207,N_19753,N_19761);
nand U20208 (N_20208,N_19949,N_19751);
or U20209 (N_20209,N_19937,N_19817);
and U20210 (N_20210,N_19766,N_19916);
nor U20211 (N_20211,N_19874,N_19788);
xor U20212 (N_20212,N_19918,N_19756);
or U20213 (N_20213,N_19931,N_19830);
nand U20214 (N_20214,N_19964,N_19944);
or U20215 (N_20215,N_19809,N_19969);
nor U20216 (N_20216,N_19925,N_19782);
nand U20217 (N_20217,N_19932,N_19781);
nor U20218 (N_20218,N_19767,N_19825);
nand U20219 (N_20219,N_19893,N_19760);
nand U20220 (N_20220,N_19920,N_19969);
nor U20221 (N_20221,N_19979,N_19772);
and U20222 (N_20222,N_19967,N_19856);
and U20223 (N_20223,N_19852,N_19791);
nor U20224 (N_20224,N_19800,N_19760);
nand U20225 (N_20225,N_19793,N_19843);
or U20226 (N_20226,N_19815,N_19952);
xnor U20227 (N_20227,N_19893,N_19755);
nand U20228 (N_20228,N_19840,N_19920);
xnor U20229 (N_20229,N_19938,N_19832);
or U20230 (N_20230,N_19815,N_19905);
xor U20231 (N_20231,N_19823,N_19804);
and U20232 (N_20232,N_19841,N_19844);
nand U20233 (N_20233,N_19895,N_19795);
nand U20234 (N_20234,N_19836,N_19860);
nor U20235 (N_20235,N_19864,N_19925);
nor U20236 (N_20236,N_19767,N_19975);
and U20237 (N_20237,N_19851,N_19759);
nand U20238 (N_20238,N_19941,N_19986);
and U20239 (N_20239,N_19798,N_19864);
or U20240 (N_20240,N_19846,N_19828);
nand U20241 (N_20241,N_19898,N_19891);
and U20242 (N_20242,N_19990,N_19852);
nand U20243 (N_20243,N_19930,N_19783);
xor U20244 (N_20244,N_19911,N_19845);
nor U20245 (N_20245,N_19821,N_19965);
and U20246 (N_20246,N_19904,N_19985);
xor U20247 (N_20247,N_19915,N_19957);
nor U20248 (N_20248,N_19808,N_19977);
xnor U20249 (N_20249,N_19973,N_19874);
xor U20250 (N_20250,N_20108,N_20000);
nand U20251 (N_20251,N_20032,N_20004);
nand U20252 (N_20252,N_20107,N_20012);
nor U20253 (N_20253,N_20139,N_20015);
xor U20254 (N_20254,N_20216,N_20071);
xor U20255 (N_20255,N_20212,N_20144);
or U20256 (N_20256,N_20023,N_20193);
nand U20257 (N_20257,N_20044,N_20030);
xnor U20258 (N_20258,N_20091,N_20122);
nor U20259 (N_20259,N_20117,N_20240);
nor U20260 (N_20260,N_20183,N_20196);
xnor U20261 (N_20261,N_20199,N_20180);
and U20262 (N_20262,N_20060,N_20088);
nor U20263 (N_20263,N_20110,N_20231);
and U20264 (N_20264,N_20152,N_20135);
nor U20265 (N_20265,N_20018,N_20035);
xor U20266 (N_20266,N_20058,N_20086);
xnor U20267 (N_20267,N_20186,N_20082);
xnor U20268 (N_20268,N_20038,N_20208);
nand U20269 (N_20269,N_20169,N_20119);
nor U20270 (N_20270,N_20151,N_20051);
nor U20271 (N_20271,N_20205,N_20085);
nand U20272 (N_20272,N_20120,N_20039);
or U20273 (N_20273,N_20153,N_20201);
and U20274 (N_20274,N_20111,N_20174);
nand U20275 (N_20275,N_20202,N_20198);
xnor U20276 (N_20276,N_20170,N_20024);
xnor U20277 (N_20277,N_20220,N_20211);
xor U20278 (N_20278,N_20072,N_20222);
or U20279 (N_20279,N_20187,N_20184);
xnor U20280 (N_20280,N_20214,N_20241);
or U20281 (N_20281,N_20116,N_20014);
nand U20282 (N_20282,N_20138,N_20195);
or U20283 (N_20283,N_20227,N_20017);
nor U20284 (N_20284,N_20092,N_20133);
nand U20285 (N_20285,N_20011,N_20146);
nand U20286 (N_20286,N_20057,N_20140);
or U20287 (N_20287,N_20073,N_20137);
nor U20288 (N_20288,N_20043,N_20010);
or U20289 (N_20289,N_20191,N_20097);
xnor U20290 (N_20290,N_20221,N_20100);
xor U20291 (N_20291,N_20114,N_20130);
or U20292 (N_20292,N_20026,N_20064);
nand U20293 (N_20293,N_20089,N_20176);
nand U20294 (N_20294,N_20020,N_20008);
and U20295 (N_20295,N_20127,N_20162);
or U20296 (N_20296,N_20123,N_20019);
nand U20297 (N_20297,N_20059,N_20042);
nand U20298 (N_20298,N_20161,N_20063);
nor U20299 (N_20299,N_20056,N_20143);
or U20300 (N_20300,N_20048,N_20192);
nand U20301 (N_20301,N_20109,N_20054);
nand U20302 (N_20302,N_20159,N_20141);
nor U20303 (N_20303,N_20239,N_20155);
xnor U20304 (N_20304,N_20021,N_20207);
and U20305 (N_20305,N_20188,N_20209);
nor U20306 (N_20306,N_20081,N_20182);
nor U20307 (N_20307,N_20052,N_20041);
nand U20308 (N_20308,N_20025,N_20145);
xor U20309 (N_20309,N_20105,N_20165);
or U20310 (N_20310,N_20112,N_20179);
nand U20311 (N_20311,N_20104,N_20232);
or U20312 (N_20312,N_20069,N_20093);
or U20313 (N_20313,N_20234,N_20156);
nor U20314 (N_20314,N_20027,N_20167);
nand U20315 (N_20315,N_20206,N_20094);
or U20316 (N_20316,N_20009,N_20163);
nand U20317 (N_20317,N_20236,N_20247);
nor U20318 (N_20318,N_20077,N_20173);
nor U20319 (N_20319,N_20246,N_20068);
nand U20320 (N_20320,N_20243,N_20045);
or U20321 (N_20321,N_20217,N_20053);
xnor U20322 (N_20322,N_20219,N_20095);
nand U20323 (N_20323,N_20062,N_20194);
or U20324 (N_20324,N_20076,N_20142);
or U20325 (N_20325,N_20128,N_20079);
and U20326 (N_20326,N_20157,N_20099);
nor U20327 (N_20327,N_20022,N_20047);
and U20328 (N_20328,N_20096,N_20102);
nor U20329 (N_20329,N_20037,N_20178);
nor U20330 (N_20330,N_20185,N_20101);
or U20331 (N_20331,N_20040,N_20129);
xnor U20332 (N_20332,N_20166,N_20225);
and U20333 (N_20333,N_20171,N_20131);
or U20334 (N_20334,N_20002,N_20050);
or U20335 (N_20335,N_20106,N_20168);
xnor U20336 (N_20336,N_20033,N_20235);
xor U20337 (N_20337,N_20055,N_20223);
or U20338 (N_20338,N_20150,N_20164);
or U20339 (N_20339,N_20249,N_20248);
or U20340 (N_20340,N_20005,N_20224);
nor U20341 (N_20341,N_20113,N_20134);
nand U20342 (N_20342,N_20080,N_20090);
xor U20343 (N_20343,N_20158,N_20244);
nand U20344 (N_20344,N_20204,N_20226);
and U20345 (N_20345,N_20233,N_20149);
nor U20346 (N_20346,N_20098,N_20125);
or U20347 (N_20347,N_20013,N_20160);
xnor U20348 (N_20348,N_20006,N_20007);
and U20349 (N_20349,N_20049,N_20238);
or U20350 (N_20350,N_20177,N_20083);
or U20351 (N_20351,N_20016,N_20242);
or U20352 (N_20352,N_20003,N_20036);
nand U20353 (N_20353,N_20148,N_20031);
and U20354 (N_20354,N_20126,N_20200);
nor U20355 (N_20355,N_20065,N_20175);
nand U20356 (N_20356,N_20118,N_20190);
nor U20357 (N_20357,N_20132,N_20213);
xnor U20358 (N_20358,N_20203,N_20087);
nand U20359 (N_20359,N_20074,N_20067);
nand U20360 (N_20360,N_20229,N_20215);
nor U20361 (N_20361,N_20136,N_20218);
xnor U20362 (N_20362,N_20189,N_20028);
and U20363 (N_20363,N_20197,N_20181);
xnor U20364 (N_20364,N_20210,N_20115);
and U20365 (N_20365,N_20075,N_20001);
xor U20366 (N_20366,N_20228,N_20084);
nand U20367 (N_20367,N_20121,N_20034);
or U20368 (N_20368,N_20172,N_20103);
xnor U20369 (N_20369,N_20066,N_20245);
nand U20370 (N_20370,N_20124,N_20029);
nor U20371 (N_20371,N_20046,N_20061);
nand U20372 (N_20372,N_20230,N_20237);
xor U20373 (N_20373,N_20078,N_20154);
xnor U20374 (N_20374,N_20147,N_20070);
nor U20375 (N_20375,N_20065,N_20139);
xnor U20376 (N_20376,N_20236,N_20208);
nand U20377 (N_20377,N_20016,N_20135);
nor U20378 (N_20378,N_20149,N_20104);
nand U20379 (N_20379,N_20207,N_20187);
xnor U20380 (N_20380,N_20069,N_20200);
xor U20381 (N_20381,N_20191,N_20052);
xor U20382 (N_20382,N_20094,N_20156);
nand U20383 (N_20383,N_20039,N_20083);
or U20384 (N_20384,N_20155,N_20001);
and U20385 (N_20385,N_20042,N_20248);
or U20386 (N_20386,N_20239,N_20184);
and U20387 (N_20387,N_20004,N_20069);
and U20388 (N_20388,N_20000,N_20219);
and U20389 (N_20389,N_20053,N_20189);
nand U20390 (N_20390,N_20085,N_20229);
or U20391 (N_20391,N_20051,N_20027);
and U20392 (N_20392,N_20114,N_20058);
xnor U20393 (N_20393,N_20013,N_20023);
nand U20394 (N_20394,N_20071,N_20195);
xor U20395 (N_20395,N_20177,N_20211);
nor U20396 (N_20396,N_20094,N_20142);
or U20397 (N_20397,N_20127,N_20041);
xor U20398 (N_20398,N_20202,N_20024);
nor U20399 (N_20399,N_20209,N_20143);
and U20400 (N_20400,N_20050,N_20188);
xnor U20401 (N_20401,N_20107,N_20063);
nor U20402 (N_20402,N_20186,N_20147);
and U20403 (N_20403,N_20125,N_20121);
nand U20404 (N_20404,N_20236,N_20100);
xnor U20405 (N_20405,N_20012,N_20132);
nor U20406 (N_20406,N_20238,N_20075);
nand U20407 (N_20407,N_20063,N_20245);
and U20408 (N_20408,N_20068,N_20041);
xnor U20409 (N_20409,N_20103,N_20226);
nand U20410 (N_20410,N_20039,N_20199);
nand U20411 (N_20411,N_20187,N_20046);
xor U20412 (N_20412,N_20049,N_20244);
nand U20413 (N_20413,N_20032,N_20180);
or U20414 (N_20414,N_20185,N_20140);
xor U20415 (N_20415,N_20008,N_20184);
nand U20416 (N_20416,N_20014,N_20152);
nor U20417 (N_20417,N_20008,N_20246);
nand U20418 (N_20418,N_20125,N_20075);
nand U20419 (N_20419,N_20025,N_20195);
nand U20420 (N_20420,N_20071,N_20120);
nand U20421 (N_20421,N_20014,N_20171);
nor U20422 (N_20422,N_20225,N_20093);
nor U20423 (N_20423,N_20168,N_20071);
nand U20424 (N_20424,N_20124,N_20061);
or U20425 (N_20425,N_20102,N_20175);
or U20426 (N_20426,N_20234,N_20019);
nor U20427 (N_20427,N_20075,N_20192);
nor U20428 (N_20428,N_20028,N_20172);
and U20429 (N_20429,N_20048,N_20071);
or U20430 (N_20430,N_20038,N_20218);
or U20431 (N_20431,N_20041,N_20018);
or U20432 (N_20432,N_20013,N_20028);
and U20433 (N_20433,N_20067,N_20160);
xor U20434 (N_20434,N_20037,N_20242);
xnor U20435 (N_20435,N_20084,N_20051);
nor U20436 (N_20436,N_20199,N_20235);
or U20437 (N_20437,N_20095,N_20237);
nor U20438 (N_20438,N_20176,N_20127);
nor U20439 (N_20439,N_20079,N_20240);
and U20440 (N_20440,N_20039,N_20100);
nor U20441 (N_20441,N_20201,N_20146);
nor U20442 (N_20442,N_20093,N_20116);
nand U20443 (N_20443,N_20153,N_20089);
xnor U20444 (N_20444,N_20210,N_20202);
nor U20445 (N_20445,N_20237,N_20168);
nand U20446 (N_20446,N_20215,N_20089);
nor U20447 (N_20447,N_20180,N_20053);
nand U20448 (N_20448,N_20051,N_20209);
and U20449 (N_20449,N_20081,N_20100);
nor U20450 (N_20450,N_20027,N_20098);
xor U20451 (N_20451,N_20015,N_20092);
or U20452 (N_20452,N_20101,N_20121);
nor U20453 (N_20453,N_20045,N_20127);
nand U20454 (N_20454,N_20198,N_20008);
xnor U20455 (N_20455,N_20052,N_20051);
or U20456 (N_20456,N_20148,N_20240);
nand U20457 (N_20457,N_20138,N_20037);
nand U20458 (N_20458,N_20105,N_20193);
nand U20459 (N_20459,N_20043,N_20049);
nand U20460 (N_20460,N_20017,N_20194);
nand U20461 (N_20461,N_20046,N_20067);
nand U20462 (N_20462,N_20178,N_20222);
or U20463 (N_20463,N_20227,N_20148);
nor U20464 (N_20464,N_20223,N_20190);
or U20465 (N_20465,N_20249,N_20022);
nand U20466 (N_20466,N_20033,N_20223);
nand U20467 (N_20467,N_20107,N_20109);
nand U20468 (N_20468,N_20117,N_20247);
or U20469 (N_20469,N_20093,N_20009);
xor U20470 (N_20470,N_20239,N_20234);
nand U20471 (N_20471,N_20125,N_20208);
nor U20472 (N_20472,N_20207,N_20063);
xnor U20473 (N_20473,N_20143,N_20236);
nand U20474 (N_20474,N_20210,N_20016);
nand U20475 (N_20475,N_20037,N_20003);
xnor U20476 (N_20476,N_20136,N_20134);
or U20477 (N_20477,N_20085,N_20016);
nor U20478 (N_20478,N_20023,N_20101);
xnor U20479 (N_20479,N_20225,N_20167);
nand U20480 (N_20480,N_20239,N_20004);
nor U20481 (N_20481,N_20006,N_20113);
nor U20482 (N_20482,N_20091,N_20186);
nand U20483 (N_20483,N_20068,N_20224);
xor U20484 (N_20484,N_20023,N_20191);
or U20485 (N_20485,N_20092,N_20028);
or U20486 (N_20486,N_20071,N_20020);
or U20487 (N_20487,N_20104,N_20077);
nor U20488 (N_20488,N_20059,N_20246);
and U20489 (N_20489,N_20026,N_20155);
nand U20490 (N_20490,N_20159,N_20231);
or U20491 (N_20491,N_20105,N_20242);
or U20492 (N_20492,N_20141,N_20213);
nor U20493 (N_20493,N_20075,N_20115);
and U20494 (N_20494,N_20230,N_20055);
nor U20495 (N_20495,N_20151,N_20170);
xnor U20496 (N_20496,N_20084,N_20235);
or U20497 (N_20497,N_20184,N_20018);
nand U20498 (N_20498,N_20204,N_20005);
nor U20499 (N_20499,N_20002,N_20146);
or U20500 (N_20500,N_20279,N_20320);
or U20501 (N_20501,N_20444,N_20305);
xnor U20502 (N_20502,N_20371,N_20433);
xnor U20503 (N_20503,N_20403,N_20280);
nand U20504 (N_20504,N_20267,N_20362);
nor U20505 (N_20505,N_20361,N_20263);
nor U20506 (N_20506,N_20349,N_20391);
and U20507 (N_20507,N_20442,N_20368);
and U20508 (N_20508,N_20259,N_20485);
and U20509 (N_20509,N_20375,N_20494);
and U20510 (N_20510,N_20430,N_20443);
xor U20511 (N_20511,N_20340,N_20301);
xnor U20512 (N_20512,N_20473,N_20441);
or U20513 (N_20513,N_20316,N_20299);
and U20514 (N_20514,N_20469,N_20312);
nand U20515 (N_20515,N_20468,N_20434);
nand U20516 (N_20516,N_20405,N_20282);
and U20517 (N_20517,N_20297,N_20483);
xor U20518 (N_20518,N_20358,N_20363);
nand U20519 (N_20519,N_20489,N_20429);
nand U20520 (N_20520,N_20360,N_20264);
nand U20521 (N_20521,N_20343,N_20439);
or U20522 (N_20522,N_20445,N_20428);
nand U20523 (N_20523,N_20265,N_20479);
or U20524 (N_20524,N_20425,N_20426);
nor U20525 (N_20525,N_20411,N_20355);
nor U20526 (N_20526,N_20332,N_20376);
nand U20527 (N_20527,N_20431,N_20386);
and U20528 (N_20528,N_20304,N_20330);
xnor U20529 (N_20529,N_20497,N_20394);
nor U20530 (N_20530,N_20339,N_20390);
nor U20531 (N_20531,N_20453,N_20315);
or U20532 (N_20532,N_20409,N_20486);
and U20533 (N_20533,N_20462,N_20333);
and U20534 (N_20534,N_20463,N_20350);
xor U20535 (N_20535,N_20250,N_20261);
or U20536 (N_20536,N_20374,N_20308);
nor U20537 (N_20537,N_20459,N_20323);
nand U20538 (N_20538,N_20290,N_20392);
nor U20539 (N_20539,N_20289,N_20474);
and U20540 (N_20540,N_20447,N_20311);
and U20541 (N_20541,N_20256,N_20370);
and U20542 (N_20542,N_20336,N_20257);
xnor U20543 (N_20543,N_20295,N_20399);
xor U20544 (N_20544,N_20342,N_20396);
and U20545 (N_20545,N_20417,N_20287);
nor U20546 (N_20546,N_20341,N_20306);
nand U20547 (N_20547,N_20464,N_20266);
and U20548 (N_20548,N_20413,N_20373);
or U20549 (N_20549,N_20388,N_20416);
nor U20550 (N_20550,N_20283,N_20458);
nor U20551 (N_20551,N_20328,N_20379);
nand U20552 (N_20552,N_20356,N_20414);
and U20553 (N_20553,N_20456,N_20288);
nand U20554 (N_20554,N_20346,N_20344);
and U20555 (N_20555,N_20406,N_20377);
xor U20556 (N_20556,N_20271,N_20300);
or U20557 (N_20557,N_20372,N_20412);
xnor U20558 (N_20558,N_20369,N_20382);
nor U20559 (N_20559,N_20421,N_20296);
xnor U20560 (N_20560,N_20407,N_20477);
nor U20561 (N_20561,N_20493,N_20278);
xor U20562 (N_20562,N_20490,N_20269);
or U20563 (N_20563,N_20471,N_20326);
or U20564 (N_20564,N_20423,N_20260);
and U20565 (N_20565,N_20364,N_20270);
or U20566 (N_20566,N_20451,N_20460);
nand U20567 (N_20567,N_20488,N_20310);
or U20568 (N_20568,N_20321,N_20365);
xnor U20569 (N_20569,N_20436,N_20378);
xnor U20570 (N_20570,N_20400,N_20366);
or U20571 (N_20571,N_20495,N_20455);
and U20572 (N_20572,N_20334,N_20251);
xnor U20573 (N_20573,N_20353,N_20415);
nand U20574 (N_20574,N_20401,N_20424);
nand U20575 (N_20575,N_20293,N_20276);
nand U20576 (N_20576,N_20307,N_20285);
and U20577 (N_20577,N_20383,N_20393);
and U20578 (N_20578,N_20291,N_20492);
or U20579 (N_20579,N_20466,N_20454);
and U20580 (N_20580,N_20435,N_20384);
and U20581 (N_20581,N_20452,N_20313);
nand U20582 (N_20582,N_20498,N_20472);
nand U20583 (N_20583,N_20461,N_20327);
nor U20584 (N_20584,N_20319,N_20255);
or U20585 (N_20585,N_20410,N_20337);
nor U20586 (N_20586,N_20418,N_20432);
or U20587 (N_20587,N_20298,N_20357);
and U20588 (N_20588,N_20397,N_20440);
xor U20589 (N_20589,N_20380,N_20385);
nand U20590 (N_20590,N_20481,N_20450);
or U20591 (N_20591,N_20359,N_20348);
or U20592 (N_20592,N_20499,N_20347);
xnor U20593 (N_20593,N_20387,N_20395);
nand U20594 (N_20594,N_20258,N_20389);
nand U20595 (N_20595,N_20273,N_20254);
nand U20596 (N_20596,N_20437,N_20478);
nand U20597 (N_20597,N_20345,N_20335);
nand U20598 (N_20598,N_20480,N_20317);
or U20599 (N_20599,N_20482,N_20272);
or U20600 (N_20600,N_20475,N_20324);
nor U20601 (N_20601,N_20496,N_20284);
nor U20602 (N_20602,N_20470,N_20419);
and U20603 (N_20603,N_20277,N_20398);
and U20604 (N_20604,N_20329,N_20338);
and U20605 (N_20605,N_20253,N_20281);
or U20606 (N_20606,N_20476,N_20438);
xor U20607 (N_20607,N_20292,N_20252);
and U20608 (N_20608,N_20427,N_20351);
nor U20609 (N_20609,N_20467,N_20302);
nor U20610 (N_20610,N_20408,N_20402);
and U20611 (N_20611,N_20325,N_20275);
nor U20612 (N_20612,N_20294,N_20268);
and U20613 (N_20613,N_20465,N_20367);
or U20614 (N_20614,N_20457,N_20354);
or U20615 (N_20615,N_20448,N_20381);
xnor U20616 (N_20616,N_20487,N_20322);
and U20617 (N_20617,N_20446,N_20274);
or U20618 (N_20618,N_20318,N_20309);
and U20619 (N_20619,N_20303,N_20491);
and U20620 (N_20620,N_20422,N_20420);
or U20621 (N_20621,N_20314,N_20484);
or U20622 (N_20622,N_20286,N_20331);
nor U20623 (N_20623,N_20404,N_20262);
nand U20624 (N_20624,N_20352,N_20449);
nor U20625 (N_20625,N_20284,N_20314);
or U20626 (N_20626,N_20468,N_20490);
or U20627 (N_20627,N_20265,N_20402);
xnor U20628 (N_20628,N_20361,N_20332);
and U20629 (N_20629,N_20430,N_20479);
xnor U20630 (N_20630,N_20388,N_20301);
and U20631 (N_20631,N_20449,N_20310);
or U20632 (N_20632,N_20263,N_20481);
nor U20633 (N_20633,N_20361,N_20358);
nor U20634 (N_20634,N_20269,N_20337);
or U20635 (N_20635,N_20354,N_20281);
nand U20636 (N_20636,N_20367,N_20437);
and U20637 (N_20637,N_20454,N_20491);
nand U20638 (N_20638,N_20255,N_20288);
nor U20639 (N_20639,N_20441,N_20364);
and U20640 (N_20640,N_20396,N_20312);
or U20641 (N_20641,N_20275,N_20372);
nor U20642 (N_20642,N_20303,N_20280);
or U20643 (N_20643,N_20252,N_20451);
nor U20644 (N_20644,N_20475,N_20273);
xnor U20645 (N_20645,N_20302,N_20468);
and U20646 (N_20646,N_20325,N_20459);
nor U20647 (N_20647,N_20429,N_20364);
or U20648 (N_20648,N_20317,N_20257);
nand U20649 (N_20649,N_20424,N_20466);
nand U20650 (N_20650,N_20363,N_20499);
nand U20651 (N_20651,N_20405,N_20437);
nand U20652 (N_20652,N_20336,N_20378);
nor U20653 (N_20653,N_20277,N_20358);
xor U20654 (N_20654,N_20477,N_20332);
xnor U20655 (N_20655,N_20453,N_20434);
and U20656 (N_20656,N_20286,N_20385);
nand U20657 (N_20657,N_20432,N_20460);
or U20658 (N_20658,N_20427,N_20396);
nand U20659 (N_20659,N_20423,N_20283);
or U20660 (N_20660,N_20471,N_20293);
and U20661 (N_20661,N_20347,N_20352);
or U20662 (N_20662,N_20495,N_20469);
or U20663 (N_20663,N_20283,N_20269);
and U20664 (N_20664,N_20259,N_20479);
nor U20665 (N_20665,N_20283,N_20293);
xnor U20666 (N_20666,N_20351,N_20316);
and U20667 (N_20667,N_20478,N_20343);
nand U20668 (N_20668,N_20374,N_20402);
or U20669 (N_20669,N_20318,N_20443);
nor U20670 (N_20670,N_20419,N_20496);
xor U20671 (N_20671,N_20260,N_20297);
nor U20672 (N_20672,N_20496,N_20449);
nand U20673 (N_20673,N_20497,N_20339);
nor U20674 (N_20674,N_20284,N_20478);
nor U20675 (N_20675,N_20382,N_20459);
nand U20676 (N_20676,N_20428,N_20492);
and U20677 (N_20677,N_20488,N_20442);
or U20678 (N_20678,N_20477,N_20377);
or U20679 (N_20679,N_20413,N_20348);
and U20680 (N_20680,N_20264,N_20418);
or U20681 (N_20681,N_20388,N_20367);
and U20682 (N_20682,N_20349,N_20355);
nand U20683 (N_20683,N_20422,N_20414);
or U20684 (N_20684,N_20395,N_20291);
xor U20685 (N_20685,N_20329,N_20362);
nor U20686 (N_20686,N_20384,N_20473);
or U20687 (N_20687,N_20443,N_20367);
nor U20688 (N_20688,N_20484,N_20268);
nand U20689 (N_20689,N_20477,N_20333);
nand U20690 (N_20690,N_20254,N_20372);
xor U20691 (N_20691,N_20461,N_20346);
or U20692 (N_20692,N_20427,N_20486);
nor U20693 (N_20693,N_20366,N_20329);
nand U20694 (N_20694,N_20353,N_20356);
nand U20695 (N_20695,N_20282,N_20298);
and U20696 (N_20696,N_20461,N_20336);
xor U20697 (N_20697,N_20455,N_20468);
and U20698 (N_20698,N_20367,N_20341);
and U20699 (N_20699,N_20305,N_20282);
xnor U20700 (N_20700,N_20350,N_20320);
xor U20701 (N_20701,N_20480,N_20324);
xnor U20702 (N_20702,N_20355,N_20306);
nor U20703 (N_20703,N_20287,N_20405);
nor U20704 (N_20704,N_20358,N_20464);
nand U20705 (N_20705,N_20445,N_20426);
nand U20706 (N_20706,N_20266,N_20319);
or U20707 (N_20707,N_20266,N_20493);
or U20708 (N_20708,N_20460,N_20278);
nand U20709 (N_20709,N_20310,N_20439);
and U20710 (N_20710,N_20493,N_20495);
nor U20711 (N_20711,N_20469,N_20289);
xnor U20712 (N_20712,N_20487,N_20358);
nor U20713 (N_20713,N_20462,N_20417);
or U20714 (N_20714,N_20312,N_20262);
xnor U20715 (N_20715,N_20363,N_20488);
nor U20716 (N_20716,N_20435,N_20363);
nand U20717 (N_20717,N_20413,N_20484);
nor U20718 (N_20718,N_20262,N_20396);
xor U20719 (N_20719,N_20356,N_20279);
or U20720 (N_20720,N_20370,N_20353);
and U20721 (N_20721,N_20255,N_20279);
or U20722 (N_20722,N_20351,N_20387);
or U20723 (N_20723,N_20366,N_20469);
xor U20724 (N_20724,N_20401,N_20340);
or U20725 (N_20725,N_20261,N_20477);
xor U20726 (N_20726,N_20399,N_20358);
or U20727 (N_20727,N_20451,N_20388);
or U20728 (N_20728,N_20398,N_20422);
nand U20729 (N_20729,N_20489,N_20456);
xor U20730 (N_20730,N_20297,N_20405);
and U20731 (N_20731,N_20460,N_20406);
xnor U20732 (N_20732,N_20492,N_20493);
and U20733 (N_20733,N_20461,N_20374);
xor U20734 (N_20734,N_20381,N_20410);
xnor U20735 (N_20735,N_20383,N_20273);
nand U20736 (N_20736,N_20438,N_20441);
nor U20737 (N_20737,N_20435,N_20406);
nand U20738 (N_20738,N_20416,N_20473);
nor U20739 (N_20739,N_20444,N_20260);
nand U20740 (N_20740,N_20457,N_20429);
nand U20741 (N_20741,N_20397,N_20277);
nand U20742 (N_20742,N_20383,N_20397);
xor U20743 (N_20743,N_20357,N_20317);
nand U20744 (N_20744,N_20438,N_20383);
nor U20745 (N_20745,N_20268,N_20443);
and U20746 (N_20746,N_20405,N_20399);
nor U20747 (N_20747,N_20266,N_20468);
xor U20748 (N_20748,N_20447,N_20349);
and U20749 (N_20749,N_20469,N_20274);
nand U20750 (N_20750,N_20677,N_20596);
nor U20751 (N_20751,N_20529,N_20632);
or U20752 (N_20752,N_20648,N_20572);
and U20753 (N_20753,N_20744,N_20679);
xor U20754 (N_20754,N_20644,N_20737);
nand U20755 (N_20755,N_20702,N_20608);
and U20756 (N_20756,N_20602,N_20694);
nand U20757 (N_20757,N_20687,N_20613);
nor U20758 (N_20758,N_20740,N_20688);
nor U20759 (N_20759,N_20542,N_20731);
nor U20760 (N_20760,N_20532,N_20664);
and U20761 (N_20761,N_20705,N_20564);
or U20762 (N_20762,N_20696,N_20745);
nor U20763 (N_20763,N_20743,N_20627);
nor U20764 (N_20764,N_20519,N_20631);
nand U20765 (N_20765,N_20601,N_20655);
or U20766 (N_20766,N_20622,N_20734);
nor U20767 (N_20767,N_20517,N_20579);
nor U20768 (N_20768,N_20553,N_20560);
or U20769 (N_20769,N_20660,N_20645);
and U20770 (N_20770,N_20656,N_20510);
nand U20771 (N_20771,N_20653,N_20649);
or U20772 (N_20772,N_20727,N_20605);
nand U20773 (N_20773,N_20685,N_20728);
or U20774 (N_20774,N_20524,N_20698);
xnor U20775 (N_20775,N_20531,N_20668);
and U20776 (N_20776,N_20665,N_20673);
xor U20777 (N_20777,N_20625,N_20508);
nor U20778 (N_20778,N_20573,N_20707);
or U20779 (N_20779,N_20551,N_20538);
nor U20780 (N_20780,N_20738,N_20512);
or U20781 (N_20781,N_20650,N_20616);
nand U20782 (N_20782,N_20599,N_20516);
xnor U20783 (N_20783,N_20507,N_20712);
nor U20784 (N_20784,N_20555,N_20500);
and U20785 (N_20785,N_20518,N_20501);
and U20786 (N_20786,N_20701,N_20629);
or U20787 (N_20787,N_20704,N_20504);
or U20788 (N_20788,N_20611,N_20556);
xor U20789 (N_20789,N_20614,N_20689);
nand U20790 (N_20790,N_20536,N_20624);
nand U20791 (N_20791,N_20747,N_20628);
or U20792 (N_20792,N_20678,N_20659);
or U20793 (N_20793,N_20526,N_20683);
nor U20794 (N_20794,N_20746,N_20580);
xor U20795 (N_20795,N_20515,N_20569);
xnor U20796 (N_20796,N_20640,N_20511);
xnor U20797 (N_20797,N_20597,N_20588);
or U20798 (N_20798,N_20574,N_20533);
or U20799 (N_20799,N_20594,N_20509);
xor U20800 (N_20800,N_20635,N_20722);
xor U20801 (N_20801,N_20530,N_20534);
xnor U20802 (N_20802,N_20612,N_20558);
or U20803 (N_20803,N_20720,N_20584);
and U20804 (N_20804,N_20642,N_20742);
or U20805 (N_20805,N_20716,N_20578);
or U20806 (N_20806,N_20709,N_20541);
nand U20807 (N_20807,N_20523,N_20658);
or U20808 (N_20808,N_20670,N_20549);
nand U20809 (N_20809,N_20714,N_20647);
xnor U20810 (N_20810,N_20711,N_20686);
xnor U20811 (N_20811,N_20563,N_20577);
xnor U20812 (N_20812,N_20733,N_20641);
and U20813 (N_20813,N_20674,N_20719);
nand U20814 (N_20814,N_20672,N_20527);
nand U20815 (N_20815,N_20600,N_20684);
nor U20816 (N_20816,N_20643,N_20646);
nor U20817 (N_20817,N_20732,N_20592);
xnor U20818 (N_20818,N_20706,N_20675);
nand U20819 (N_20819,N_20559,N_20703);
xor U20820 (N_20820,N_20595,N_20514);
and U20821 (N_20821,N_20585,N_20654);
nand U20822 (N_20822,N_20544,N_20561);
and U20823 (N_20823,N_20520,N_20657);
or U20824 (N_20824,N_20617,N_20552);
nand U20825 (N_20825,N_20651,N_20626);
xor U20826 (N_20826,N_20699,N_20591);
and U20827 (N_20827,N_20663,N_20535);
or U20828 (N_20828,N_20662,N_20506);
and U20829 (N_20829,N_20713,N_20726);
nand U20830 (N_20830,N_20708,N_20637);
or U20831 (N_20831,N_20715,N_20598);
nand U20832 (N_20832,N_20607,N_20676);
or U20833 (N_20833,N_20691,N_20741);
or U20834 (N_20834,N_20749,N_20606);
nor U20835 (N_20835,N_20525,N_20521);
nand U20836 (N_20836,N_20697,N_20576);
nand U20837 (N_20837,N_20636,N_20583);
nand U20838 (N_20838,N_20550,N_20575);
xnor U20839 (N_20839,N_20695,N_20603);
or U20840 (N_20840,N_20522,N_20502);
and U20841 (N_20841,N_20610,N_20671);
xnor U20842 (N_20842,N_20639,N_20537);
or U20843 (N_20843,N_20739,N_20593);
nand U20844 (N_20844,N_20634,N_20586);
xnor U20845 (N_20845,N_20729,N_20590);
nand U20846 (N_20846,N_20615,N_20604);
or U20847 (N_20847,N_20736,N_20582);
and U20848 (N_20848,N_20717,N_20540);
nand U20849 (N_20849,N_20547,N_20620);
nand U20850 (N_20850,N_20693,N_20589);
or U20851 (N_20851,N_20546,N_20587);
nor U20852 (N_20852,N_20619,N_20690);
or U20853 (N_20853,N_20667,N_20730);
and U20854 (N_20854,N_20666,N_20638);
nor U20855 (N_20855,N_20570,N_20528);
xnor U20856 (N_20856,N_20721,N_20568);
nor U20857 (N_20857,N_20581,N_20725);
or U20858 (N_20858,N_20681,N_20557);
or U20859 (N_20859,N_20543,N_20669);
and U20860 (N_20860,N_20567,N_20539);
nor U20861 (N_20861,N_20633,N_20554);
nand U20862 (N_20862,N_20723,N_20513);
nor U20863 (N_20863,N_20571,N_20652);
or U20864 (N_20864,N_20710,N_20618);
nand U20865 (N_20865,N_20609,N_20548);
nand U20866 (N_20866,N_20565,N_20623);
nand U20867 (N_20867,N_20724,N_20661);
nand U20868 (N_20868,N_20566,N_20748);
nor U20869 (N_20869,N_20505,N_20545);
nand U20870 (N_20870,N_20692,N_20503);
nand U20871 (N_20871,N_20680,N_20718);
or U20872 (N_20872,N_20735,N_20682);
nand U20873 (N_20873,N_20562,N_20700);
nand U20874 (N_20874,N_20621,N_20630);
and U20875 (N_20875,N_20548,N_20748);
nand U20876 (N_20876,N_20503,N_20509);
nand U20877 (N_20877,N_20603,N_20500);
nor U20878 (N_20878,N_20550,N_20704);
or U20879 (N_20879,N_20746,N_20610);
nor U20880 (N_20880,N_20590,N_20737);
and U20881 (N_20881,N_20710,N_20665);
nand U20882 (N_20882,N_20682,N_20632);
xnor U20883 (N_20883,N_20638,N_20736);
or U20884 (N_20884,N_20563,N_20732);
or U20885 (N_20885,N_20649,N_20689);
xnor U20886 (N_20886,N_20577,N_20593);
nor U20887 (N_20887,N_20650,N_20748);
nor U20888 (N_20888,N_20704,N_20586);
xnor U20889 (N_20889,N_20560,N_20547);
xnor U20890 (N_20890,N_20604,N_20743);
nand U20891 (N_20891,N_20660,N_20507);
or U20892 (N_20892,N_20524,N_20686);
or U20893 (N_20893,N_20710,N_20727);
nor U20894 (N_20894,N_20516,N_20549);
xnor U20895 (N_20895,N_20508,N_20688);
and U20896 (N_20896,N_20749,N_20562);
nand U20897 (N_20897,N_20701,N_20607);
or U20898 (N_20898,N_20557,N_20545);
xor U20899 (N_20899,N_20747,N_20713);
or U20900 (N_20900,N_20510,N_20734);
nor U20901 (N_20901,N_20655,N_20617);
and U20902 (N_20902,N_20685,N_20738);
and U20903 (N_20903,N_20691,N_20645);
and U20904 (N_20904,N_20550,N_20570);
nand U20905 (N_20905,N_20666,N_20532);
or U20906 (N_20906,N_20576,N_20655);
and U20907 (N_20907,N_20571,N_20542);
nor U20908 (N_20908,N_20548,N_20681);
nor U20909 (N_20909,N_20609,N_20607);
nand U20910 (N_20910,N_20620,N_20531);
nand U20911 (N_20911,N_20669,N_20522);
nand U20912 (N_20912,N_20690,N_20593);
and U20913 (N_20913,N_20650,N_20516);
and U20914 (N_20914,N_20520,N_20518);
nand U20915 (N_20915,N_20595,N_20700);
or U20916 (N_20916,N_20646,N_20601);
nor U20917 (N_20917,N_20732,N_20699);
xor U20918 (N_20918,N_20609,N_20584);
and U20919 (N_20919,N_20641,N_20691);
or U20920 (N_20920,N_20700,N_20741);
and U20921 (N_20921,N_20665,N_20661);
xor U20922 (N_20922,N_20576,N_20503);
nand U20923 (N_20923,N_20500,N_20526);
nand U20924 (N_20924,N_20691,N_20528);
or U20925 (N_20925,N_20616,N_20747);
nor U20926 (N_20926,N_20573,N_20678);
nand U20927 (N_20927,N_20639,N_20659);
xor U20928 (N_20928,N_20582,N_20732);
nor U20929 (N_20929,N_20710,N_20713);
nor U20930 (N_20930,N_20620,N_20647);
or U20931 (N_20931,N_20561,N_20501);
nor U20932 (N_20932,N_20685,N_20565);
nor U20933 (N_20933,N_20702,N_20676);
xor U20934 (N_20934,N_20635,N_20718);
xnor U20935 (N_20935,N_20690,N_20696);
nand U20936 (N_20936,N_20693,N_20549);
nor U20937 (N_20937,N_20678,N_20733);
nor U20938 (N_20938,N_20655,N_20709);
nand U20939 (N_20939,N_20622,N_20512);
or U20940 (N_20940,N_20720,N_20580);
or U20941 (N_20941,N_20570,N_20653);
nor U20942 (N_20942,N_20571,N_20712);
nor U20943 (N_20943,N_20545,N_20729);
or U20944 (N_20944,N_20597,N_20560);
and U20945 (N_20945,N_20639,N_20570);
xor U20946 (N_20946,N_20709,N_20678);
or U20947 (N_20947,N_20727,N_20565);
and U20948 (N_20948,N_20653,N_20618);
xor U20949 (N_20949,N_20675,N_20741);
nor U20950 (N_20950,N_20620,N_20566);
xor U20951 (N_20951,N_20683,N_20678);
or U20952 (N_20952,N_20531,N_20579);
nand U20953 (N_20953,N_20722,N_20609);
nand U20954 (N_20954,N_20546,N_20653);
or U20955 (N_20955,N_20624,N_20747);
or U20956 (N_20956,N_20541,N_20560);
nand U20957 (N_20957,N_20608,N_20615);
xor U20958 (N_20958,N_20620,N_20645);
or U20959 (N_20959,N_20662,N_20639);
or U20960 (N_20960,N_20666,N_20693);
or U20961 (N_20961,N_20558,N_20583);
nor U20962 (N_20962,N_20612,N_20743);
nor U20963 (N_20963,N_20666,N_20735);
nand U20964 (N_20964,N_20719,N_20709);
nand U20965 (N_20965,N_20671,N_20637);
nor U20966 (N_20966,N_20624,N_20651);
nand U20967 (N_20967,N_20749,N_20577);
or U20968 (N_20968,N_20715,N_20548);
nor U20969 (N_20969,N_20632,N_20531);
and U20970 (N_20970,N_20639,N_20566);
and U20971 (N_20971,N_20572,N_20638);
or U20972 (N_20972,N_20748,N_20728);
nor U20973 (N_20973,N_20547,N_20696);
xor U20974 (N_20974,N_20689,N_20605);
or U20975 (N_20975,N_20651,N_20568);
or U20976 (N_20976,N_20714,N_20624);
nand U20977 (N_20977,N_20577,N_20568);
xor U20978 (N_20978,N_20747,N_20728);
and U20979 (N_20979,N_20509,N_20522);
and U20980 (N_20980,N_20636,N_20732);
nand U20981 (N_20981,N_20521,N_20663);
nand U20982 (N_20982,N_20725,N_20658);
or U20983 (N_20983,N_20688,N_20511);
or U20984 (N_20984,N_20747,N_20706);
nor U20985 (N_20985,N_20518,N_20623);
and U20986 (N_20986,N_20674,N_20576);
nor U20987 (N_20987,N_20657,N_20621);
nor U20988 (N_20988,N_20733,N_20670);
nand U20989 (N_20989,N_20573,N_20692);
nor U20990 (N_20990,N_20694,N_20615);
or U20991 (N_20991,N_20702,N_20585);
nor U20992 (N_20992,N_20570,N_20650);
and U20993 (N_20993,N_20621,N_20580);
nor U20994 (N_20994,N_20600,N_20645);
nor U20995 (N_20995,N_20700,N_20594);
nor U20996 (N_20996,N_20655,N_20692);
xnor U20997 (N_20997,N_20708,N_20574);
nand U20998 (N_20998,N_20590,N_20669);
nor U20999 (N_20999,N_20551,N_20708);
nor U21000 (N_21000,N_20815,N_20764);
or U21001 (N_21001,N_20950,N_20990);
and U21002 (N_21002,N_20868,N_20839);
nor U21003 (N_21003,N_20967,N_20768);
xnor U21004 (N_21004,N_20958,N_20751);
or U21005 (N_21005,N_20808,N_20770);
xnor U21006 (N_21006,N_20983,N_20830);
nand U21007 (N_21007,N_20991,N_20833);
and U21008 (N_21008,N_20820,N_20921);
or U21009 (N_21009,N_20865,N_20925);
or U21010 (N_21010,N_20875,N_20846);
or U21011 (N_21011,N_20943,N_20787);
xnor U21012 (N_21012,N_20767,N_20858);
or U21013 (N_21013,N_20989,N_20763);
xor U21014 (N_21014,N_20962,N_20776);
xnor U21015 (N_21015,N_20933,N_20963);
nand U21016 (N_21016,N_20999,N_20765);
and U21017 (N_21017,N_20784,N_20826);
xnor U21018 (N_21018,N_20900,N_20936);
xor U21019 (N_21019,N_20806,N_20997);
xnor U21020 (N_21020,N_20812,N_20807);
xnor U21021 (N_21021,N_20759,N_20877);
or U21022 (N_21022,N_20932,N_20895);
xor U21023 (N_21023,N_20831,N_20977);
nor U21024 (N_21024,N_20859,N_20948);
and U21025 (N_21025,N_20988,N_20785);
nand U21026 (N_21026,N_20952,N_20917);
nor U21027 (N_21027,N_20802,N_20824);
and U21028 (N_21028,N_20836,N_20891);
and U21029 (N_21029,N_20881,N_20845);
xor U21030 (N_21030,N_20788,N_20918);
and U21031 (N_21031,N_20772,N_20754);
or U21032 (N_21032,N_20916,N_20973);
nand U21033 (N_21033,N_20811,N_20797);
xor U21034 (N_21034,N_20857,N_20834);
nor U21035 (N_21035,N_20888,N_20984);
or U21036 (N_21036,N_20955,N_20804);
and U21037 (N_21037,N_20796,N_20885);
nor U21038 (N_21038,N_20994,N_20927);
xnor U21039 (N_21039,N_20795,N_20930);
nor U21040 (N_21040,N_20896,N_20957);
xor U21041 (N_21041,N_20819,N_20931);
or U21042 (N_21042,N_20926,N_20904);
and U21043 (N_21043,N_20898,N_20982);
and U21044 (N_21044,N_20774,N_20870);
or U21045 (N_21045,N_20777,N_20861);
and U21046 (N_21046,N_20901,N_20899);
xor U21047 (N_21047,N_20854,N_20908);
nor U21048 (N_21048,N_20869,N_20756);
nor U21049 (N_21049,N_20817,N_20934);
nor U21050 (N_21050,N_20954,N_20947);
nor U21051 (N_21051,N_20938,N_20769);
and U21052 (N_21052,N_20829,N_20970);
or U21053 (N_21053,N_20856,N_20987);
and U21054 (N_21054,N_20922,N_20941);
nand U21055 (N_21055,N_20832,N_20873);
nand U21056 (N_21056,N_20940,N_20883);
xnor U21057 (N_21057,N_20949,N_20993);
nand U21058 (N_21058,N_20907,N_20841);
nand U21059 (N_21059,N_20974,N_20844);
or U21060 (N_21060,N_20814,N_20969);
or U21061 (N_21061,N_20976,N_20848);
xnor U21062 (N_21062,N_20880,N_20799);
and U21063 (N_21063,N_20971,N_20783);
xor U21064 (N_21064,N_20909,N_20851);
and U21065 (N_21065,N_20913,N_20876);
and U21066 (N_21066,N_20850,N_20864);
nor U21067 (N_21067,N_20779,N_20871);
or U21068 (N_21068,N_20985,N_20965);
nand U21069 (N_21069,N_20755,N_20752);
nand U21070 (N_21070,N_20942,N_20920);
or U21071 (N_21071,N_20966,N_20758);
or U21072 (N_21072,N_20929,N_20939);
nand U21073 (N_21073,N_20872,N_20995);
nor U21074 (N_21074,N_20937,N_20975);
nand U21075 (N_21075,N_20910,N_20778);
or U21076 (N_21076,N_20803,N_20894);
xnor U21077 (N_21077,N_20790,N_20761);
nor U21078 (N_21078,N_20810,N_20825);
and U21079 (N_21079,N_20843,N_20786);
nor U21080 (N_21080,N_20842,N_20757);
nand U21081 (N_21081,N_20890,N_20809);
and U21082 (N_21082,N_20914,N_20912);
and U21083 (N_21083,N_20944,N_20775);
nor U21084 (N_21084,N_20813,N_20903);
or U21085 (N_21085,N_20905,N_20882);
and U21086 (N_21086,N_20863,N_20791);
nand U21087 (N_21087,N_20821,N_20853);
and U21088 (N_21088,N_20911,N_20961);
and U21089 (N_21089,N_20782,N_20915);
xor U21090 (N_21090,N_20798,N_20886);
and U21091 (N_21091,N_20823,N_20818);
nand U21092 (N_21092,N_20766,N_20980);
and U21093 (N_21093,N_20945,N_20884);
nand U21094 (N_21094,N_20816,N_20773);
or U21095 (N_21095,N_20847,N_20959);
or U21096 (N_21096,N_20855,N_20960);
and U21097 (N_21097,N_20860,N_20906);
xor U21098 (N_21098,N_20781,N_20878);
nor U21099 (N_21099,N_20835,N_20789);
nand U21100 (N_21100,N_20919,N_20981);
or U21101 (N_21101,N_20794,N_20968);
nand U21102 (N_21102,N_20889,N_20964);
nand U21103 (N_21103,N_20923,N_20771);
nand U21104 (N_21104,N_20998,N_20753);
nor U21105 (N_21105,N_20827,N_20996);
nand U21106 (N_21106,N_20838,N_20992);
and U21107 (N_21107,N_20828,N_20972);
xor U21108 (N_21108,N_20953,N_20951);
nand U21109 (N_21109,N_20840,N_20879);
nand U21110 (N_21110,N_20874,N_20793);
nand U21111 (N_21111,N_20892,N_20792);
nor U21112 (N_21112,N_20979,N_20862);
or U21113 (N_21113,N_20801,N_20897);
xnor U21114 (N_21114,N_20893,N_20978);
nand U21115 (N_21115,N_20946,N_20762);
nor U21116 (N_21116,N_20805,N_20837);
nand U21117 (N_21117,N_20866,N_20928);
or U21118 (N_21118,N_20849,N_20780);
nor U21119 (N_21119,N_20986,N_20800);
or U21120 (N_21120,N_20822,N_20887);
xor U21121 (N_21121,N_20750,N_20867);
xor U21122 (N_21122,N_20852,N_20902);
xor U21123 (N_21123,N_20935,N_20924);
nand U21124 (N_21124,N_20956,N_20760);
xor U21125 (N_21125,N_20793,N_20978);
and U21126 (N_21126,N_20972,N_20947);
nand U21127 (N_21127,N_20912,N_20902);
or U21128 (N_21128,N_20952,N_20915);
nor U21129 (N_21129,N_20920,N_20975);
and U21130 (N_21130,N_20899,N_20960);
xnor U21131 (N_21131,N_20987,N_20818);
xor U21132 (N_21132,N_20792,N_20805);
nand U21133 (N_21133,N_20782,N_20993);
nand U21134 (N_21134,N_20755,N_20799);
xnor U21135 (N_21135,N_20974,N_20902);
xnor U21136 (N_21136,N_20767,N_20954);
nor U21137 (N_21137,N_20992,N_20993);
nand U21138 (N_21138,N_20949,N_20793);
nor U21139 (N_21139,N_20866,N_20910);
or U21140 (N_21140,N_20901,N_20766);
nand U21141 (N_21141,N_20793,N_20794);
xor U21142 (N_21142,N_20906,N_20777);
or U21143 (N_21143,N_20876,N_20812);
or U21144 (N_21144,N_20967,N_20974);
and U21145 (N_21145,N_20976,N_20897);
xor U21146 (N_21146,N_20948,N_20925);
xnor U21147 (N_21147,N_20805,N_20806);
xor U21148 (N_21148,N_20902,N_20853);
nand U21149 (N_21149,N_20766,N_20879);
nand U21150 (N_21150,N_20752,N_20847);
and U21151 (N_21151,N_20996,N_20927);
or U21152 (N_21152,N_20837,N_20924);
and U21153 (N_21153,N_20967,N_20962);
xnor U21154 (N_21154,N_20989,N_20851);
xor U21155 (N_21155,N_20936,N_20916);
and U21156 (N_21156,N_20941,N_20758);
or U21157 (N_21157,N_20915,N_20785);
nand U21158 (N_21158,N_20867,N_20887);
nor U21159 (N_21159,N_20793,N_20931);
xnor U21160 (N_21160,N_20973,N_20897);
or U21161 (N_21161,N_20913,N_20983);
and U21162 (N_21162,N_20975,N_20882);
nor U21163 (N_21163,N_20779,N_20985);
xnor U21164 (N_21164,N_20850,N_20808);
xor U21165 (N_21165,N_20928,N_20820);
nor U21166 (N_21166,N_20875,N_20784);
and U21167 (N_21167,N_20977,N_20958);
nand U21168 (N_21168,N_20857,N_20782);
nor U21169 (N_21169,N_20958,N_20885);
and U21170 (N_21170,N_20763,N_20935);
nor U21171 (N_21171,N_20882,N_20839);
or U21172 (N_21172,N_20803,N_20972);
nor U21173 (N_21173,N_20915,N_20995);
and U21174 (N_21174,N_20966,N_20766);
and U21175 (N_21175,N_20810,N_20881);
xor U21176 (N_21176,N_20825,N_20865);
nor U21177 (N_21177,N_20852,N_20879);
xnor U21178 (N_21178,N_20982,N_20953);
and U21179 (N_21179,N_20788,N_20800);
xor U21180 (N_21180,N_20766,N_20964);
or U21181 (N_21181,N_20961,N_20985);
and U21182 (N_21182,N_20969,N_20984);
xnor U21183 (N_21183,N_20925,N_20964);
xor U21184 (N_21184,N_20828,N_20949);
and U21185 (N_21185,N_20870,N_20799);
or U21186 (N_21186,N_20933,N_20834);
and U21187 (N_21187,N_20898,N_20921);
nand U21188 (N_21188,N_20857,N_20773);
nand U21189 (N_21189,N_20996,N_20830);
nand U21190 (N_21190,N_20874,N_20910);
nand U21191 (N_21191,N_20940,N_20757);
nand U21192 (N_21192,N_20989,N_20999);
nand U21193 (N_21193,N_20771,N_20828);
xor U21194 (N_21194,N_20953,N_20829);
and U21195 (N_21195,N_20972,N_20920);
or U21196 (N_21196,N_20999,N_20858);
nand U21197 (N_21197,N_20854,N_20915);
nor U21198 (N_21198,N_20945,N_20867);
or U21199 (N_21199,N_20801,N_20836);
nor U21200 (N_21200,N_20814,N_20855);
and U21201 (N_21201,N_20789,N_20780);
nor U21202 (N_21202,N_20849,N_20905);
xor U21203 (N_21203,N_20960,N_20998);
nand U21204 (N_21204,N_20891,N_20840);
nand U21205 (N_21205,N_20804,N_20788);
or U21206 (N_21206,N_20985,N_20929);
or U21207 (N_21207,N_20811,N_20997);
or U21208 (N_21208,N_20817,N_20921);
and U21209 (N_21209,N_20999,N_20851);
xor U21210 (N_21210,N_20899,N_20937);
xnor U21211 (N_21211,N_20992,N_20976);
xnor U21212 (N_21212,N_20842,N_20999);
nor U21213 (N_21213,N_20931,N_20943);
or U21214 (N_21214,N_20991,N_20866);
nor U21215 (N_21215,N_20856,N_20921);
nor U21216 (N_21216,N_20778,N_20751);
and U21217 (N_21217,N_20914,N_20808);
and U21218 (N_21218,N_20863,N_20824);
or U21219 (N_21219,N_20881,N_20820);
nor U21220 (N_21220,N_20993,N_20972);
nor U21221 (N_21221,N_20852,N_20886);
or U21222 (N_21222,N_20758,N_20760);
nor U21223 (N_21223,N_20873,N_20821);
nor U21224 (N_21224,N_20951,N_20766);
xnor U21225 (N_21225,N_20847,N_20872);
nand U21226 (N_21226,N_20949,N_20959);
and U21227 (N_21227,N_20812,N_20883);
or U21228 (N_21228,N_20893,N_20919);
nand U21229 (N_21229,N_20985,N_20791);
xor U21230 (N_21230,N_20802,N_20894);
nand U21231 (N_21231,N_20817,N_20945);
xor U21232 (N_21232,N_20999,N_20957);
or U21233 (N_21233,N_20925,N_20847);
nor U21234 (N_21234,N_20924,N_20764);
or U21235 (N_21235,N_20969,N_20878);
xnor U21236 (N_21236,N_20973,N_20909);
nor U21237 (N_21237,N_20944,N_20859);
or U21238 (N_21238,N_20863,N_20843);
and U21239 (N_21239,N_20991,N_20913);
xnor U21240 (N_21240,N_20811,N_20852);
nand U21241 (N_21241,N_20784,N_20752);
nor U21242 (N_21242,N_20854,N_20944);
xor U21243 (N_21243,N_20772,N_20898);
xor U21244 (N_21244,N_20919,N_20977);
and U21245 (N_21245,N_20992,N_20817);
nand U21246 (N_21246,N_20948,N_20906);
nor U21247 (N_21247,N_20882,N_20915);
nand U21248 (N_21248,N_20965,N_20964);
nand U21249 (N_21249,N_20985,N_20787);
and U21250 (N_21250,N_21212,N_21205);
xor U21251 (N_21251,N_21243,N_21005);
or U21252 (N_21252,N_21246,N_21001);
nand U21253 (N_21253,N_21194,N_21007);
nor U21254 (N_21254,N_21126,N_21010);
nand U21255 (N_21255,N_21223,N_21198);
nor U21256 (N_21256,N_21053,N_21081);
and U21257 (N_21257,N_21030,N_21049);
nand U21258 (N_21258,N_21119,N_21201);
xor U21259 (N_21259,N_21233,N_21141);
nor U21260 (N_21260,N_21057,N_21112);
nor U21261 (N_21261,N_21241,N_21036);
and U21262 (N_21262,N_21115,N_21156);
nor U21263 (N_21263,N_21166,N_21035);
nor U21264 (N_21264,N_21144,N_21229);
nor U21265 (N_21265,N_21244,N_21026);
xnor U21266 (N_21266,N_21074,N_21134);
xnor U21267 (N_21267,N_21140,N_21217);
xnor U21268 (N_21268,N_21143,N_21164);
nor U21269 (N_21269,N_21025,N_21228);
and U21270 (N_21270,N_21152,N_21042);
nand U21271 (N_21271,N_21127,N_21031);
nand U21272 (N_21272,N_21017,N_21102);
nand U21273 (N_21273,N_21145,N_21169);
nand U21274 (N_21274,N_21065,N_21050);
and U21275 (N_21275,N_21063,N_21003);
nor U21276 (N_21276,N_21104,N_21182);
and U21277 (N_21277,N_21037,N_21231);
nand U21278 (N_21278,N_21022,N_21162);
nand U21279 (N_21279,N_21148,N_21114);
or U21280 (N_21280,N_21062,N_21086);
nand U21281 (N_21281,N_21069,N_21135);
and U21282 (N_21282,N_21096,N_21172);
nand U21283 (N_21283,N_21206,N_21167);
nor U21284 (N_21284,N_21240,N_21099);
nand U21285 (N_21285,N_21165,N_21097);
or U21286 (N_21286,N_21103,N_21098);
and U21287 (N_21287,N_21041,N_21207);
or U21288 (N_21288,N_21218,N_21208);
xnor U21289 (N_21289,N_21123,N_21046);
and U21290 (N_21290,N_21236,N_21058);
xor U21291 (N_21291,N_21157,N_21109);
xnor U21292 (N_21292,N_21091,N_21138);
xor U21293 (N_21293,N_21133,N_21193);
and U21294 (N_21294,N_21130,N_21178);
xor U21295 (N_21295,N_21021,N_21000);
or U21296 (N_21296,N_21237,N_21158);
xnor U21297 (N_21297,N_21070,N_21071);
xor U21298 (N_21298,N_21048,N_21120);
and U21299 (N_21299,N_21214,N_21171);
xnor U21300 (N_21300,N_21200,N_21234);
and U21301 (N_21301,N_21192,N_21044);
and U21302 (N_21302,N_21202,N_21004);
xor U21303 (N_21303,N_21073,N_21146);
nand U21304 (N_21304,N_21242,N_21018);
and U21305 (N_21305,N_21177,N_21189);
nor U21306 (N_21306,N_21075,N_21006);
or U21307 (N_21307,N_21088,N_21105);
xor U21308 (N_21308,N_21082,N_21161);
nand U21309 (N_21309,N_21084,N_21154);
nand U21310 (N_21310,N_21064,N_21122);
xor U21311 (N_21311,N_21121,N_21222);
nand U21312 (N_21312,N_21078,N_21029);
xor U21313 (N_21313,N_21174,N_21173);
or U21314 (N_21314,N_21137,N_21072);
and U21315 (N_21315,N_21113,N_21068);
xnor U21316 (N_21316,N_21232,N_21219);
nor U21317 (N_21317,N_21187,N_21188);
or U21318 (N_21318,N_21052,N_21209);
xor U21319 (N_21319,N_21083,N_21226);
nor U21320 (N_21320,N_21195,N_21125);
or U21321 (N_21321,N_21080,N_21221);
or U21322 (N_21322,N_21028,N_21110);
and U21323 (N_21323,N_21040,N_21094);
xor U21324 (N_21324,N_21248,N_21227);
nand U21325 (N_21325,N_21225,N_21160);
and U21326 (N_21326,N_21054,N_21067);
nand U21327 (N_21327,N_21090,N_21016);
nand U21328 (N_21328,N_21211,N_21034);
xor U21329 (N_21329,N_21213,N_21131);
xor U21330 (N_21330,N_21111,N_21047);
nor U21331 (N_21331,N_21076,N_21089);
nand U21332 (N_21332,N_21061,N_21051);
nor U21333 (N_21333,N_21224,N_21033);
and U21334 (N_21334,N_21093,N_21181);
nor U21335 (N_21335,N_21011,N_21235);
and U21336 (N_21336,N_21204,N_21203);
nor U21337 (N_21337,N_21185,N_21176);
nand U21338 (N_21338,N_21183,N_21118);
nand U21339 (N_21339,N_21190,N_21077);
nor U21340 (N_21340,N_21085,N_21139);
and U21341 (N_21341,N_21024,N_21002);
or U21342 (N_21342,N_21249,N_21092);
xor U21343 (N_21343,N_21100,N_21039);
and U21344 (N_21344,N_21106,N_21015);
and U21345 (N_21345,N_21136,N_21163);
nor U21346 (N_21346,N_21142,N_21199);
nand U21347 (N_21347,N_21132,N_21032);
or U21348 (N_21348,N_21168,N_21151);
or U21349 (N_21349,N_21055,N_21230);
nand U21350 (N_21350,N_21196,N_21009);
nand U21351 (N_21351,N_21155,N_21095);
nand U21352 (N_21352,N_21056,N_21013);
nor U21353 (N_21353,N_21184,N_21175);
nand U21354 (N_21354,N_21060,N_21128);
xnor U21355 (N_21355,N_21043,N_21186);
or U21356 (N_21356,N_21179,N_21215);
or U21357 (N_21357,N_21238,N_21059);
nand U21358 (N_21358,N_21008,N_21159);
xor U21359 (N_21359,N_21012,N_21023);
and U21360 (N_21360,N_21116,N_21038);
nand U21361 (N_21361,N_21027,N_21108);
or U21362 (N_21362,N_21170,N_21019);
nand U21363 (N_21363,N_21101,N_21247);
or U21364 (N_21364,N_21216,N_21107);
or U21365 (N_21365,N_21220,N_21197);
nor U21366 (N_21366,N_21147,N_21117);
xnor U21367 (N_21367,N_21014,N_21191);
and U21368 (N_21368,N_21079,N_21210);
and U21369 (N_21369,N_21239,N_21045);
nand U21370 (N_21370,N_21066,N_21124);
nand U21371 (N_21371,N_21087,N_21153);
or U21372 (N_21372,N_21245,N_21129);
and U21373 (N_21373,N_21180,N_21149);
nand U21374 (N_21374,N_21150,N_21020);
nor U21375 (N_21375,N_21213,N_21228);
xor U21376 (N_21376,N_21211,N_21122);
xor U21377 (N_21377,N_21032,N_21203);
or U21378 (N_21378,N_21144,N_21091);
and U21379 (N_21379,N_21055,N_21227);
and U21380 (N_21380,N_21224,N_21151);
nand U21381 (N_21381,N_21167,N_21222);
and U21382 (N_21382,N_21233,N_21106);
xnor U21383 (N_21383,N_21120,N_21206);
nand U21384 (N_21384,N_21225,N_21050);
xor U21385 (N_21385,N_21042,N_21121);
xnor U21386 (N_21386,N_21180,N_21160);
xnor U21387 (N_21387,N_21100,N_21049);
nor U21388 (N_21388,N_21208,N_21100);
xor U21389 (N_21389,N_21191,N_21039);
nor U21390 (N_21390,N_21137,N_21044);
nand U21391 (N_21391,N_21076,N_21074);
nand U21392 (N_21392,N_21204,N_21244);
nor U21393 (N_21393,N_21133,N_21137);
nand U21394 (N_21394,N_21008,N_21198);
and U21395 (N_21395,N_21097,N_21096);
and U21396 (N_21396,N_21011,N_21223);
and U21397 (N_21397,N_21003,N_21171);
or U21398 (N_21398,N_21087,N_21233);
and U21399 (N_21399,N_21236,N_21168);
and U21400 (N_21400,N_21200,N_21067);
xor U21401 (N_21401,N_21100,N_21162);
nor U21402 (N_21402,N_21241,N_21086);
nor U21403 (N_21403,N_21231,N_21056);
or U21404 (N_21404,N_21185,N_21103);
nand U21405 (N_21405,N_21150,N_21247);
and U21406 (N_21406,N_21202,N_21137);
nand U21407 (N_21407,N_21068,N_21037);
nor U21408 (N_21408,N_21084,N_21176);
or U21409 (N_21409,N_21241,N_21235);
and U21410 (N_21410,N_21190,N_21242);
xnor U21411 (N_21411,N_21189,N_21241);
and U21412 (N_21412,N_21222,N_21055);
xor U21413 (N_21413,N_21237,N_21057);
or U21414 (N_21414,N_21152,N_21249);
and U21415 (N_21415,N_21061,N_21230);
or U21416 (N_21416,N_21119,N_21240);
nand U21417 (N_21417,N_21017,N_21079);
xnor U21418 (N_21418,N_21107,N_21218);
xor U21419 (N_21419,N_21059,N_21010);
nand U21420 (N_21420,N_21109,N_21053);
and U21421 (N_21421,N_21173,N_21000);
and U21422 (N_21422,N_21068,N_21039);
nand U21423 (N_21423,N_21090,N_21222);
xor U21424 (N_21424,N_21164,N_21087);
or U21425 (N_21425,N_21130,N_21038);
nand U21426 (N_21426,N_21013,N_21095);
and U21427 (N_21427,N_21213,N_21055);
or U21428 (N_21428,N_21185,N_21121);
or U21429 (N_21429,N_21095,N_21087);
nand U21430 (N_21430,N_21135,N_21121);
and U21431 (N_21431,N_21121,N_21084);
and U21432 (N_21432,N_21190,N_21139);
or U21433 (N_21433,N_21062,N_21010);
nor U21434 (N_21434,N_21214,N_21124);
nand U21435 (N_21435,N_21163,N_21047);
nor U21436 (N_21436,N_21137,N_21021);
xnor U21437 (N_21437,N_21096,N_21222);
or U21438 (N_21438,N_21137,N_21050);
xor U21439 (N_21439,N_21218,N_21151);
or U21440 (N_21440,N_21190,N_21194);
xnor U21441 (N_21441,N_21047,N_21125);
nor U21442 (N_21442,N_21077,N_21233);
xnor U21443 (N_21443,N_21201,N_21200);
xor U21444 (N_21444,N_21068,N_21122);
xnor U21445 (N_21445,N_21146,N_21136);
xnor U21446 (N_21446,N_21175,N_21165);
and U21447 (N_21447,N_21084,N_21234);
nand U21448 (N_21448,N_21030,N_21215);
and U21449 (N_21449,N_21003,N_21042);
or U21450 (N_21450,N_21051,N_21105);
nand U21451 (N_21451,N_21152,N_21081);
nor U21452 (N_21452,N_21173,N_21225);
and U21453 (N_21453,N_21084,N_21110);
nor U21454 (N_21454,N_21054,N_21076);
nor U21455 (N_21455,N_21034,N_21204);
nand U21456 (N_21456,N_21234,N_21222);
nand U21457 (N_21457,N_21086,N_21208);
and U21458 (N_21458,N_21229,N_21057);
or U21459 (N_21459,N_21003,N_21038);
nand U21460 (N_21460,N_21041,N_21164);
nor U21461 (N_21461,N_21096,N_21138);
nand U21462 (N_21462,N_21148,N_21010);
or U21463 (N_21463,N_21145,N_21018);
and U21464 (N_21464,N_21232,N_21183);
xnor U21465 (N_21465,N_21248,N_21042);
nor U21466 (N_21466,N_21114,N_21206);
nand U21467 (N_21467,N_21089,N_21099);
nor U21468 (N_21468,N_21107,N_21131);
and U21469 (N_21469,N_21065,N_21230);
xnor U21470 (N_21470,N_21154,N_21015);
and U21471 (N_21471,N_21078,N_21209);
or U21472 (N_21472,N_21210,N_21163);
xor U21473 (N_21473,N_21031,N_21244);
nand U21474 (N_21474,N_21113,N_21128);
and U21475 (N_21475,N_21146,N_21173);
nand U21476 (N_21476,N_21090,N_21033);
xor U21477 (N_21477,N_21152,N_21238);
xnor U21478 (N_21478,N_21231,N_21015);
nor U21479 (N_21479,N_21074,N_21057);
or U21480 (N_21480,N_21034,N_21235);
nand U21481 (N_21481,N_21127,N_21213);
xor U21482 (N_21482,N_21234,N_21053);
nor U21483 (N_21483,N_21215,N_21005);
and U21484 (N_21484,N_21122,N_21153);
and U21485 (N_21485,N_21000,N_21166);
nor U21486 (N_21486,N_21094,N_21139);
xnor U21487 (N_21487,N_21135,N_21134);
or U21488 (N_21488,N_21212,N_21146);
nand U21489 (N_21489,N_21147,N_21240);
nand U21490 (N_21490,N_21219,N_21238);
nand U21491 (N_21491,N_21232,N_21115);
nor U21492 (N_21492,N_21001,N_21115);
nand U21493 (N_21493,N_21136,N_21175);
and U21494 (N_21494,N_21209,N_21244);
nand U21495 (N_21495,N_21239,N_21024);
and U21496 (N_21496,N_21146,N_21000);
xor U21497 (N_21497,N_21024,N_21004);
nor U21498 (N_21498,N_21122,N_21089);
xor U21499 (N_21499,N_21038,N_21089);
nor U21500 (N_21500,N_21365,N_21351);
nand U21501 (N_21501,N_21259,N_21318);
xor U21502 (N_21502,N_21454,N_21373);
nor U21503 (N_21503,N_21412,N_21312);
nand U21504 (N_21504,N_21385,N_21397);
nand U21505 (N_21505,N_21427,N_21350);
xnor U21506 (N_21506,N_21422,N_21374);
and U21507 (N_21507,N_21409,N_21381);
nor U21508 (N_21508,N_21466,N_21478);
xor U21509 (N_21509,N_21430,N_21278);
and U21510 (N_21510,N_21276,N_21489);
nor U21511 (N_21511,N_21487,N_21462);
and U21512 (N_21512,N_21260,N_21436);
and U21513 (N_21513,N_21303,N_21379);
nor U21514 (N_21514,N_21459,N_21299);
xnor U21515 (N_21515,N_21283,N_21419);
xnor U21516 (N_21516,N_21370,N_21393);
and U21517 (N_21517,N_21463,N_21302);
nor U21518 (N_21518,N_21407,N_21333);
or U21519 (N_21519,N_21477,N_21306);
or U21520 (N_21520,N_21414,N_21438);
and U21521 (N_21521,N_21343,N_21496);
or U21522 (N_21522,N_21335,N_21420);
nor U21523 (N_21523,N_21482,N_21354);
nor U21524 (N_21524,N_21458,N_21258);
nor U21525 (N_21525,N_21417,N_21456);
or U21526 (N_21526,N_21392,N_21433);
nor U21527 (N_21527,N_21326,N_21254);
nor U21528 (N_21528,N_21310,N_21411);
and U21529 (N_21529,N_21358,N_21285);
nand U21530 (N_21530,N_21263,N_21428);
xnor U21531 (N_21531,N_21323,N_21348);
and U21532 (N_21532,N_21395,N_21368);
nor U21533 (N_21533,N_21415,N_21396);
nand U21534 (N_21534,N_21342,N_21360);
nor U21535 (N_21535,N_21495,N_21324);
or U21536 (N_21536,N_21284,N_21329);
nand U21537 (N_21537,N_21455,N_21322);
nand U21538 (N_21538,N_21431,N_21451);
or U21539 (N_21539,N_21378,N_21346);
nor U21540 (N_21540,N_21443,N_21340);
or U21541 (N_21541,N_21446,N_21376);
and U21542 (N_21542,N_21253,N_21344);
nand U21543 (N_21543,N_21405,N_21265);
nand U21544 (N_21544,N_21286,N_21304);
nor U21545 (N_21545,N_21311,N_21319);
xor U21546 (N_21546,N_21293,N_21315);
or U21547 (N_21547,N_21426,N_21290);
nor U21548 (N_21548,N_21316,N_21300);
or U21549 (N_21549,N_21400,N_21382);
nor U21550 (N_21550,N_21484,N_21366);
or U21551 (N_21551,N_21398,N_21367);
xnor U21552 (N_21552,N_21251,N_21467);
and U21553 (N_21553,N_21464,N_21475);
or U21554 (N_21554,N_21255,N_21468);
and U21555 (N_21555,N_21364,N_21356);
and U21556 (N_21556,N_21390,N_21491);
or U21557 (N_21557,N_21252,N_21408);
nand U21558 (N_21558,N_21490,N_21410);
xor U21559 (N_21559,N_21272,N_21476);
nor U21560 (N_21560,N_21372,N_21387);
xnor U21561 (N_21561,N_21347,N_21359);
nor U21562 (N_21562,N_21361,N_21352);
xor U21563 (N_21563,N_21314,N_21256);
and U21564 (N_21564,N_21404,N_21271);
and U21565 (N_21565,N_21289,N_21295);
xor U21566 (N_21566,N_21401,N_21309);
nand U21567 (N_21567,N_21472,N_21413);
nand U21568 (N_21568,N_21273,N_21345);
nor U21569 (N_21569,N_21432,N_21429);
and U21570 (N_21570,N_21386,N_21406);
or U21571 (N_21571,N_21341,N_21403);
nor U21572 (N_21572,N_21479,N_21388);
nor U21573 (N_21573,N_21380,N_21357);
xnor U21574 (N_21574,N_21377,N_21457);
nor U21575 (N_21575,N_21317,N_21442);
and U21576 (N_21576,N_21444,N_21434);
or U21577 (N_21577,N_21305,N_21362);
nand U21578 (N_21578,N_21355,N_21371);
nor U21579 (N_21579,N_21450,N_21287);
and U21580 (N_21580,N_21474,N_21307);
nor U21581 (N_21581,N_21391,N_21288);
and U21582 (N_21582,N_21339,N_21369);
nand U21583 (N_21583,N_21470,N_21447);
xnor U21584 (N_21584,N_21337,N_21330);
nand U21585 (N_21585,N_21269,N_21469);
or U21586 (N_21586,N_21353,N_21402);
xor U21587 (N_21587,N_21325,N_21449);
xor U21588 (N_21588,N_21296,N_21279);
nor U21589 (N_21589,N_21461,N_21298);
nor U21590 (N_21590,N_21483,N_21270);
xnor U21591 (N_21591,N_21338,N_21445);
xnor U21592 (N_21592,N_21282,N_21275);
nand U21593 (N_21593,N_21308,N_21257);
nor U21594 (N_21594,N_21332,N_21418);
xnor U21595 (N_21595,N_21320,N_21448);
nand U21596 (N_21596,N_21480,N_21416);
or U21597 (N_21597,N_21264,N_21473);
xor U21598 (N_21598,N_21375,N_21423);
nand U21599 (N_21599,N_21266,N_21331);
or U21600 (N_21600,N_21327,N_21493);
nor U21601 (N_21601,N_21453,N_21349);
or U21602 (N_21602,N_21250,N_21452);
nand U21603 (N_21603,N_21262,N_21313);
nor U21604 (N_21604,N_21280,N_21460);
nand U21605 (N_21605,N_21439,N_21425);
nand U21606 (N_21606,N_21384,N_21297);
or U21607 (N_21607,N_21485,N_21499);
or U21608 (N_21608,N_21494,N_21437);
nor U21609 (N_21609,N_21267,N_21294);
nor U21610 (N_21610,N_21383,N_21301);
nand U21611 (N_21611,N_21328,N_21281);
nand U21612 (N_21612,N_21421,N_21277);
nor U21613 (N_21613,N_21481,N_21488);
or U21614 (N_21614,N_21291,N_21389);
nor U21615 (N_21615,N_21399,N_21492);
nand U21616 (N_21616,N_21336,N_21268);
nand U21617 (N_21617,N_21334,N_21363);
or U21618 (N_21618,N_21440,N_21498);
nand U21619 (N_21619,N_21292,N_21394);
or U21620 (N_21620,N_21486,N_21441);
and U21621 (N_21621,N_21465,N_21424);
and U21622 (N_21622,N_21261,N_21321);
nand U21623 (N_21623,N_21471,N_21435);
and U21624 (N_21624,N_21274,N_21497);
nor U21625 (N_21625,N_21312,N_21337);
and U21626 (N_21626,N_21407,N_21319);
nand U21627 (N_21627,N_21322,N_21466);
nand U21628 (N_21628,N_21292,N_21400);
and U21629 (N_21629,N_21343,N_21401);
and U21630 (N_21630,N_21426,N_21381);
nand U21631 (N_21631,N_21309,N_21268);
or U21632 (N_21632,N_21496,N_21276);
nand U21633 (N_21633,N_21472,N_21494);
nor U21634 (N_21634,N_21320,N_21381);
and U21635 (N_21635,N_21372,N_21356);
or U21636 (N_21636,N_21270,N_21262);
and U21637 (N_21637,N_21321,N_21460);
xnor U21638 (N_21638,N_21396,N_21380);
nand U21639 (N_21639,N_21253,N_21464);
and U21640 (N_21640,N_21388,N_21458);
xor U21641 (N_21641,N_21325,N_21462);
nand U21642 (N_21642,N_21320,N_21327);
and U21643 (N_21643,N_21352,N_21453);
or U21644 (N_21644,N_21425,N_21435);
nand U21645 (N_21645,N_21484,N_21250);
or U21646 (N_21646,N_21338,N_21287);
xor U21647 (N_21647,N_21337,N_21490);
xnor U21648 (N_21648,N_21391,N_21402);
nor U21649 (N_21649,N_21310,N_21407);
nor U21650 (N_21650,N_21473,N_21332);
nand U21651 (N_21651,N_21423,N_21463);
nand U21652 (N_21652,N_21334,N_21319);
nor U21653 (N_21653,N_21281,N_21380);
and U21654 (N_21654,N_21348,N_21306);
xnor U21655 (N_21655,N_21256,N_21366);
or U21656 (N_21656,N_21442,N_21321);
and U21657 (N_21657,N_21266,N_21491);
xor U21658 (N_21658,N_21437,N_21425);
nand U21659 (N_21659,N_21442,N_21362);
xnor U21660 (N_21660,N_21343,N_21452);
xor U21661 (N_21661,N_21265,N_21426);
and U21662 (N_21662,N_21347,N_21330);
or U21663 (N_21663,N_21340,N_21252);
nor U21664 (N_21664,N_21484,N_21352);
nor U21665 (N_21665,N_21475,N_21406);
xnor U21666 (N_21666,N_21472,N_21499);
nor U21667 (N_21667,N_21367,N_21361);
nand U21668 (N_21668,N_21491,N_21476);
nand U21669 (N_21669,N_21466,N_21264);
xor U21670 (N_21670,N_21436,N_21476);
nand U21671 (N_21671,N_21276,N_21338);
and U21672 (N_21672,N_21343,N_21482);
nand U21673 (N_21673,N_21311,N_21378);
nor U21674 (N_21674,N_21285,N_21403);
nand U21675 (N_21675,N_21418,N_21382);
or U21676 (N_21676,N_21468,N_21326);
nand U21677 (N_21677,N_21438,N_21356);
and U21678 (N_21678,N_21408,N_21327);
and U21679 (N_21679,N_21316,N_21322);
nor U21680 (N_21680,N_21495,N_21455);
and U21681 (N_21681,N_21413,N_21420);
nor U21682 (N_21682,N_21387,N_21405);
nor U21683 (N_21683,N_21257,N_21350);
and U21684 (N_21684,N_21432,N_21478);
nand U21685 (N_21685,N_21484,N_21422);
and U21686 (N_21686,N_21490,N_21252);
and U21687 (N_21687,N_21444,N_21277);
xnor U21688 (N_21688,N_21342,N_21277);
and U21689 (N_21689,N_21369,N_21441);
nand U21690 (N_21690,N_21425,N_21273);
nand U21691 (N_21691,N_21315,N_21304);
nor U21692 (N_21692,N_21289,N_21253);
nor U21693 (N_21693,N_21369,N_21415);
xor U21694 (N_21694,N_21270,N_21294);
nor U21695 (N_21695,N_21366,N_21381);
or U21696 (N_21696,N_21252,N_21271);
and U21697 (N_21697,N_21464,N_21366);
and U21698 (N_21698,N_21467,N_21279);
nor U21699 (N_21699,N_21400,N_21414);
nand U21700 (N_21700,N_21398,N_21429);
xnor U21701 (N_21701,N_21449,N_21499);
xnor U21702 (N_21702,N_21339,N_21440);
xnor U21703 (N_21703,N_21375,N_21475);
and U21704 (N_21704,N_21255,N_21497);
nor U21705 (N_21705,N_21480,N_21389);
xor U21706 (N_21706,N_21389,N_21420);
or U21707 (N_21707,N_21402,N_21398);
or U21708 (N_21708,N_21432,N_21343);
nand U21709 (N_21709,N_21460,N_21384);
nor U21710 (N_21710,N_21439,N_21490);
xnor U21711 (N_21711,N_21385,N_21363);
nor U21712 (N_21712,N_21284,N_21297);
or U21713 (N_21713,N_21426,N_21419);
or U21714 (N_21714,N_21445,N_21358);
nor U21715 (N_21715,N_21493,N_21498);
or U21716 (N_21716,N_21325,N_21327);
or U21717 (N_21717,N_21367,N_21334);
xnor U21718 (N_21718,N_21291,N_21360);
xnor U21719 (N_21719,N_21495,N_21463);
nand U21720 (N_21720,N_21334,N_21421);
nand U21721 (N_21721,N_21458,N_21474);
nor U21722 (N_21722,N_21352,N_21364);
nor U21723 (N_21723,N_21267,N_21358);
nor U21724 (N_21724,N_21278,N_21347);
and U21725 (N_21725,N_21290,N_21292);
xnor U21726 (N_21726,N_21369,N_21250);
or U21727 (N_21727,N_21256,N_21499);
or U21728 (N_21728,N_21317,N_21319);
nor U21729 (N_21729,N_21363,N_21476);
nand U21730 (N_21730,N_21293,N_21255);
nand U21731 (N_21731,N_21347,N_21496);
nor U21732 (N_21732,N_21258,N_21289);
and U21733 (N_21733,N_21306,N_21374);
nor U21734 (N_21734,N_21280,N_21419);
and U21735 (N_21735,N_21421,N_21292);
nand U21736 (N_21736,N_21471,N_21269);
or U21737 (N_21737,N_21252,N_21411);
or U21738 (N_21738,N_21415,N_21385);
nor U21739 (N_21739,N_21383,N_21366);
and U21740 (N_21740,N_21303,N_21401);
and U21741 (N_21741,N_21255,N_21432);
nor U21742 (N_21742,N_21267,N_21436);
and U21743 (N_21743,N_21438,N_21433);
nor U21744 (N_21744,N_21289,N_21301);
xnor U21745 (N_21745,N_21268,N_21313);
nand U21746 (N_21746,N_21250,N_21487);
and U21747 (N_21747,N_21276,N_21330);
nand U21748 (N_21748,N_21405,N_21426);
and U21749 (N_21749,N_21266,N_21441);
xnor U21750 (N_21750,N_21653,N_21532);
or U21751 (N_21751,N_21586,N_21625);
nand U21752 (N_21752,N_21642,N_21633);
nor U21753 (N_21753,N_21675,N_21683);
nor U21754 (N_21754,N_21596,N_21672);
xor U21755 (N_21755,N_21583,N_21643);
or U21756 (N_21756,N_21537,N_21598);
and U21757 (N_21757,N_21521,N_21613);
and U21758 (N_21758,N_21562,N_21579);
and U21759 (N_21759,N_21713,N_21748);
xor U21760 (N_21760,N_21727,N_21529);
xor U21761 (N_21761,N_21716,N_21735);
nor U21762 (N_21762,N_21730,N_21592);
nand U21763 (N_21763,N_21684,N_21539);
nor U21764 (N_21764,N_21569,N_21743);
nand U21765 (N_21765,N_21589,N_21605);
and U21766 (N_21766,N_21651,N_21720);
or U21767 (N_21767,N_21600,N_21594);
or U21768 (N_21768,N_21565,N_21658);
xnor U21769 (N_21769,N_21558,N_21506);
or U21770 (N_21770,N_21513,N_21527);
xnor U21771 (N_21771,N_21706,N_21515);
or U21772 (N_21772,N_21645,N_21508);
or U21773 (N_21773,N_21501,N_21610);
and U21774 (N_21774,N_21574,N_21563);
xor U21775 (N_21775,N_21522,N_21674);
xnor U21776 (N_21776,N_21557,N_21657);
and U21777 (N_21777,N_21536,N_21571);
or U21778 (N_21778,N_21622,N_21662);
and U21779 (N_21779,N_21620,N_21719);
or U21780 (N_21780,N_21544,N_21746);
and U21781 (N_21781,N_21612,N_21699);
nor U21782 (N_21782,N_21697,N_21604);
nand U21783 (N_21783,N_21688,N_21677);
nor U21784 (N_21784,N_21577,N_21603);
and U21785 (N_21785,N_21647,N_21680);
nand U21786 (N_21786,N_21654,N_21686);
or U21787 (N_21787,N_21663,N_21567);
or U21788 (N_21788,N_21718,N_21714);
nor U21789 (N_21789,N_21690,N_21619);
xnor U21790 (N_21790,N_21650,N_21512);
and U21791 (N_21791,N_21561,N_21676);
and U21792 (N_21792,N_21599,N_21597);
xor U21793 (N_21793,N_21668,N_21570);
nor U21794 (N_21794,N_21649,N_21543);
nand U21795 (N_21795,N_21670,N_21514);
or U21796 (N_21796,N_21568,N_21664);
xnor U21797 (N_21797,N_21593,N_21656);
and U21798 (N_21798,N_21629,N_21660);
or U21799 (N_21799,N_21530,N_21511);
or U21800 (N_21800,N_21737,N_21505);
or U21801 (N_21801,N_21548,N_21715);
xor U21802 (N_21802,N_21538,N_21559);
or U21803 (N_21803,N_21726,N_21627);
xnor U21804 (N_21804,N_21646,N_21608);
or U21805 (N_21805,N_21736,N_21724);
nor U21806 (N_21806,N_21703,N_21671);
and U21807 (N_21807,N_21673,N_21692);
nand U21808 (N_21808,N_21623,N_21694);
nor U21809 (N_21809,N_21523,N_21580);
or U21810 (N_21810,N_21723,N_21609);
nor U21811 (N_21811,N_21744,N_21507);
nor U21812 (N_21812,N_21742,N_21510);
and U21813 (N_21813,N_21524,N_21528);
xor U21814 (N_21814,N_21549,N_21631);
nor U21815 (N_21815,N_21704,N_21659);
or U21816 (N_21816,N_21552,N_21667);
nand U21817 (N_21817,N_21541,N_21624);
nor U21818 (N_21818,N_21578,N_21740);
and U21819 (N_21819,N_21518,N_21711);
nor U21820 (N_21820,N_21682,N_21734);
nor U21821 (N_21821,N_21534,N_21636);
xnor U21822 (N_21822,N_21635,N_21587);
or U21823 (N_21823,N_21560,N_21601);
xor U21824 (N_21824,N_21526,N_21705);
xor U21825 (N_21825,N_21572,N_21591);
xnor U21826 (N_21826,N_21732,N_21707);
nand U21827 (N_21827,N_21553,N_21621);
xor U21828 (N_21828,N_21687,N_21747);
and U21829 (N_21829,N_21693,N_21729);
or U21830 (N_21830,N_21566,N_21545);
or U21831 (N_21831,N_21733,N_21554);
nand U21832 (N_21832,N_21644,N_21585);
or U21833 (N_21833,N_21722,N_21638);
xnor U21834 (N_21834,N_21519,N_21710);
xnor U21835 (N_21835,N_21655,N_21590);
xnor U21836 (N_21836,N_21738,N_21731);
nor U21837 (N_21837,N_21531,N_21576);
or U21838 (N_21838,N_21588,N_21616);
nand U21839 (N_21839,N_21542,N_21728);
nor U21840 (N_21840,N_21626,N_21678);
xnor U21841 (N_21841,N_21509,N_21634);
or U21842 (N_21842,N_21745,N_21695);
or U21843 (N_21843,N_21637,N_21500);
and U21844 (N_21844,N_21614,N_21661);
nor U21845 (N_21845,N_21652,N_21696);
nand U21846 (N_21846,N_21611,N_21640);
xor U21847 (N_21847,N_21630,N_21556);
nor U21848 (N_21848,N_21739,N_21669);
nand U21849 (N_21849,N_21535,N_21628);
or U21850 (N_21850,N_21717,N_21648);
and U21851 (N_21851,N_21709,N_21641);
or U21852 (N_21852,N_21691,N_21679);
nor U21853 (N_21853,N_21607,N_21584);
or U21854 (N_21854,N_21525,N_21749);
xor U21855 (N_21855,N_21602,N_21581);
nand U21856 (N_21856,N_21547,N_21575);
nor U21857 (N_21857,N_21504,N_21632);
nand U21858 (N_21858,N_21550,N_21551);
xnor U21859 (N_21859,N_21573,N_21639);
nand U21860 (N_21860,N_21618,N_21617);
nand U21861 (N_21861,N_21503,N_21533);
xor U21862 (N_21862,N_21708,N_21689);
or U21863 (N_21863,N_21546,N_21595);
or U21864 (N_21864,N_21681,N_21725);
nand U21865 (N_21865,N_21564,N_21721);
nor U21866 (N_21866,N_21516,N_21555);
and U21867 (N_21867,N_21615,N_21665);
xor U21868 (N_21868,N_21741,N_21582);
xor U21869 (N_21869,N_21502,N_21666);
and U21870 (N_21870,N_21517,N_21702);
xor U21871 (N_21871,N_21712,N_21520);
nand U21872 (N_21872,N_21701,N_21685);
nand U21873 (N_21873,N_21606,N_21700);
nand U21874 (N_21874,N_21698,N_21540);
or U21875 (N_21875,N_21558,N_21612);
and U21876 (N_21876,N_21595,N_21578);
or U21877 (N_21877,N_21689,N_21564);
and U21878 (N_21878,N_21689,N_21733);
nor U21879 (N_21879,N_21615,N_21526);
nor U21880 (N_21880,N_21578,N_21742);
or U21881 (N_21881,N_21610,N_21556);
or U21882 (N_21882,N_21735,N_21580);
xor U21883 (N_21883,N_21517,N_21708);
or U21884 (N_21884,N_21573,N_21512);
nor U21885 (N_21885,N_21652,N_21660);
xor U21886 (N_21886,N_21725,N_21578);
or U21887 (N_21887,N_21510,N_21562);
or U21888 (N_21888,N_21707,N_21529);
or U21889 (N_21889,N_21521,N_21658);
or U21890 (N_21890,N_21538,N_21697);
xor U21891 (N_21891,N_21567,N_21568);
and U21892 (N_21892,N_21608,N_21605);
nor U21893 (N_21893,N_21664,N_21615);
and U21894 (N_21894,N_21573,N_21576);
xnor U21895 (N_21895,N_21704,N_21633);
and U21896 (N_21896,N_21507,N_21541);
xnor U21897 (N_21897,N_21734,N_21614);
nor U21898 (N_21898,N_21550,N_21645);
nand U21899 (N_21899,N_21650,N_21504);
or U21900 (N_21900,N_21556,N_21705);
xor U21901 (N_21901,N_21651,N_21672);
nor U21902 (N_21902,N_21584,N_21523);
and U21903 (N_21903,N_21516,N_21648);
xor U21904 (N_21904,N_21507,N_21527);
nand U21905 (N_21905,N_21548,N_21673);
and U21906 (N_21906,N_21673,N_21572);
xor U21907 (N_21907,N_21595,N_21615);
xnor U21908 (N_21908,N_21682,N_21730);
and U21909 (N_21909,N_21579,N_21667);
and U21910 (N_21910,N_21702,N_21600);
and U21911 (N_21911,N_21560,N_21558);
nand U21912 (N_21912,N_21710,N_21672);
nand U21913 (N_21913,N_21725,N_21645);
and U21914 (N_21914,N_21623,N_21673);
xor U21915 (N_21915,N_21662,N_21691);
or U21916 (N_21916,N_21718,N_21704);
and U21917 (N_21917,N_21545,N_21749);
nand U21918 (N_21918,N_21553,N_21665);
nand U21919 (N_21919,N_21600,N_21744);
xnor U21920 (N_21920,N_21709,N_21582);
nand U21921 (N_21921,N_21574,N_21517);
xor U21922 (N_21922,N_21714,N_21554);
or U21923 (N_21923,N_21693,N_21540);
and U21924 (N_21924,N_21505,N_21671);
or U21925 (N_21925,N_21555,N_21638);
xnor U21926 (N_21926,N_21511,N_21675);
or U21927 (N_21927,N_21735,N_21687);
or U21928 (N_21928,N_21548,N_21546);
xnor U21929 (N_21929,N_21627,N_21538);
and U21930 (N_21930,N_21660,N_21664);
or U21931 (N_21931,N_21653,N_21534);
nor U21932 (N_21932,N_21589,N_21546);
or U21933 (N_21933,N_21730,N_21732);
nor U21934 (N_21934,N_21591,N_21602);
and U21935 (N_21935,N_21643,N_21705);
or U21936 (N_21936,N_21715,N_21620);
xor U21937 (N_21937,N_21515,N_21504);
or U21938 (N_21938,N_21687,N_21688);
nand U21939 (N_21939,N_21553,N_21739);
nand U21940 (N_21940,N_21626,N_21633);
and U21941 (N_21941,N_21601,N_21736);
and U21942 (N_21942,N_21553,N_21692);
or U21943 (N_21943,N_21705,N_21575);
xnor U21944 (N_21944,N_21577,N_21520);
nand U21945 (N_21945,N_21561,N_21721);
xor U21946 (N_21946,N_21566,N_21687);
xor U21947 (N_21947,N_21738,N_21613);
nor U21948 (N_21948,N_21512,N_21738);
nand U21949 (N_21949,N_21740,N_21732);
nand U21950 (N_21950,N_21731,N_21730);
nand U21951 (N_21951,N_21734,N_21727);
xnor U21952 (N_21952,N_21695,N_21615);
xnor U21953 (N_21953,N_21638,N_21515);
and U21954 (N_21954,N_21682,N_21572);
and U21955 (N_21955,N_21646,N_21691);
nand U21956 (N_21956,N_21719,N_21500);
nand U21957 (N_21957,N_21504,N_21688);
xnor U21958 (N_21958,N_21678,N_21589);
and U21959 (N_21959,N_21699,N_21564);
or U21960 (N_21960,N_21737,N_21541);
and U21961 (N_21961,N_21511,N_21630);
and U21962 (N_21962,N_21707,N_21696);
nor U21963 (N_21963,N_21506,N_21614);
xnor U21964 (N_21964,N_21730,N_21515);
nor U21965 (N_21965,N_21560,N_21646);
and U21966 (N_21966,N_21542,N_21581);
and U21967 (N_21967,N_21685,N_21563);
or U21968 (N_21968,N_21575,N_21566);
or U21969 (N_21969,N_21659,N_21718);
and U21970 (N_21970,N_21542,N_21577);
and U21971 (N_21971,N_21668,N_21519);
nand U21972 (N_21972,N_21708,N_21536);
xor U21973 (N_21973,N_21594,N_21740);
nor U21974 (N_21974,N_21526,N_21603);
xor U21975 (N_21975,N_21567,N_21579);
nor U21976 (N_21976,N_21507,N_21740);
or U21977 (N_21977,N_21537,N_21605);
nand U21978 (N_21978,N_21642,N_21632);
and U21979 (N_21979,N_21604,N_21657);
and U21980 (N_21980,N_21635,N_21576);
xor U21981 (N_21981,N_21623,N_21632);
and U21982 (N_21982,N_21675,N_21509);
or U21983 (N_21983,N_21713,N_21703);
nor U21984 (N_21984,N_21509,N_21715);
xor U21985 (N_21985,N_21741,N_21608);
xnor U21986 (N_21986,N_21552,N_21582);
and U21987 (N_21987,N_21620,N_21525);
and U21988 (N_21988,N_21668,N_21649);
nand U21989 (N_21989,N_21582,N_21644);
nand U21990 (N_21990,N_21615,N_21522);
xnor U21991 (N_21991,N_21541,N_21650);
nor U21992 (N_21992,N_21563,N_21570);
and U21993 (N_21993,N_21666,N_21742);
nand U21994 (N_21994,N_21580,N_21617);
nand U21995 (N_21995,N_21669,N_21531);
nand U21996 (N_21996,N_21640,N_21605);
nor U21997 (N_21997,N_21603,N_21702);
xor U21998 (N_21998,N_21695,N_21634);
nand U21999 (N_21999,N_21679,N_21522);
or U22000 (N_22000,N_21935,N_21920);
xnor U22001 (N_22001,N_21969,N_21883);
xnor U22002 (N_22002,N_21786,N_21846);
or U22003 (N_22003,N_21824,N_21823);
nand U22004 (N_22004,N_21832,N_21819);
or U22005 (N_22005,N_21964,N_21976);
nand U22006 (N_22006,N_21947,N_21818);
nor U22007 (N_22007,N_21765,N_21766);
or U22008 (N_22008,N_21862,N_21955);
nor U22009 (N_22009,N_21871,N_21879);
nor U22010 (N_22010,N_21926,N_21813);
xor U22011 (N_22011,N_21796,N_21866);
xnor U22012 (N_22012,N_21779,N_21854);
nor U22013 (N_22013,N_21804,N_21830);
and U22014 (N_22014,N_21960,N_21762);
nand U22015 (N_22015,N_21915,N_21867);
or U22016 (N_22016,N_21812,N_21948);
nor U22017 (N_22017,N_21918,N_21931);
or U22018 (N_22018,N_21774,N_21761);
or U22019 (N_22019,N_21869,N_21886);
xnor U22020 (N_22020,N_21921,N_21954);
xor U22021 (N_22021,N_21777,N_21968);
xor U22022 (N_22022,N_21755,N_21899);
xnor U22023 (N_22023,N_21949,N_21875);
or U22024 (N_22024,N_21999,N_21900);
xor U22025 (N_22025,N_21942,N_21885);
or U22026 (N_22026,N_21923,N_21870);
nor U22027 (N_22027,N_21973,N_21946);
nand U22028 (N_22028,N_21930,N_21961);
and U22029 (N_22029,N_21843,N_21892);
and U22030 (N_22030,N_21877,N_21993);
and U22031 (N_22031,N_21971,N_21790);
or U22032 (N_22032,N_21884,N_21927);
nor U22033 (N_22033,N_21943,N_21811);
or U22034 (N_22034,N_21863,N_21939);
or U22035 (N_22035,N_21836,N_21778);
xnor U22036 (N_22036,N_21963,N_21994);
nor U22037 (N_22037,N_21834,N_21768);
nor U22038 (N_22038,N_21996,N_21895);
or U22039 (N_22039,N_21965,N_21751);
and U22040 (N_22040,N_21983,N_21838);
and U22041 (N_22041,N_21896,N_21882);
and U22042 (N_22042,N_21853,N_21929);
xnor U22043 (N_22043,N_21922,N_21910);
and U22044 (N_22044,N_21905,N_21801);
and U22045 (N_22045,N_21820,N_21924);
or U22046 (N_22046,N_21912,N_21835);
nand U22047 (N_22047,N_21917,N_21855);
and U22048 (N_22048,N_21798,N_21986);
or U22049 (N_22049,N_21980,N_21767);
nand U22050 (N_22050,N_21962,N_21898);
nor U22051 (N_22051,N_21858,N_21860);
or U22052 (N_22052,N_21831,N_21894);
nor U22053 (N_22053,N_21764,N_21967);
or U22054 (N_22054,N_21848,N_21932);
or U22055 (N_22055,N_21906,N_21889);
nand U22056 (N_22056,N_21881,N_21814);
and U22057 (N_22057,N_21776,N_21785);
nand U22058 (N_22058,N_21850,N_21990);
and U22059 (N_22059,N_21979,N_21771);
xor U22060 (N_22060,N_21757,N_21989);
and U22061 (N_22061,N_21933,N_21950);
nand U22062 (N_22062,N_21822,N_21919);
xor U22063 (N_22063,N_21893,N_21878);
nor U22064 (N_22064,N_21940,N_21840);
xor U22065 (N_22065,N_21995,N_21988);
xnor U22066 (N_22066,N_21998,N_21966);
xnor U22067 (N_22067,N_21857,N_21756);
and U22068 (N_22068,N_21972,N_21826);
xnor U22069 (N_22069,N_21752,N_21815);
nand U22070 (N_22070,N_21902,N_21958);
and U22071 (N_22071,N_21991,N_21974);
xnor U22072 (N_22072,N_21849,N_21890);
or U22073 (N_22073,N_21829,N_21852);
nor U22074 (N_22074,N_21783,N_21944);
and U22075 (N_22075,N_21945,N_21951);
nand U22076 (N_22076,N_21975,N_21861);
nor U22077 (N_22077,N_21799,N_21800);
and U22078 (N_22078,N_21833,N_21789);
and U22079 (N_22079,N_21821,N_21903);
and U22080 (N_22080,N_21997,N_21982);
and U22081 (N_22081,N_21876,N_21909);
nand U22082 (N_22082,N_21753,N_21803);
nand U22083 (N_22083,N_21908,N_21773);
or U22084 (N_22084,N_21987,N_21816);
nor U22085 (N_22085,N_21793,N_21763);
xor U22086 (N_22086,N_21788,N_21891);
nand U22087 (N_22087,N_21797,N_21772);
nand U22088 (N_22088,N_21805,N_21952);
and U22089 (N_22089,N_21758,N_21981);
xor U22090 (N_22090,N_21957,N_21978);
and U22091 (N_22091,N_21775,N_21754);
xnor U22092 (N_22092,N_21873,N_21817);
nand U22093 (N_22093,N_21839,N_21934);
xnor U22094 (N_22094,N_21825,N_21888);
nor U22095 (N_22095,N_21916,N_21844);
nor U22096 (N_22096,N_21759,N_21938);
or U22097 (N_22097,N_21913,N_21925);
nand U22098 (N_22098,N_21956,N_21959);
nor U22099 (N_22099,N_21780,N_21806);
or U22100 (N_22100,N_21937,N_21936);
xor U22101 (N_22101,N_21807,N_21911);
and U22102 (N_22102,N_21897,N_21770);
nor U22103 (N_22103,N_21985,N_21901);
xor U22104 (N_22104,N_21795,N_21904);
nand U22105 (N_22105,N_21992,N_21864);
xor U22106 (N_22106,N_21984,N_21970);
or U22107 (N_22107,N_21856,N_21859);
nor U22108 (N_22108,N_21842,N_21809);
or U22109 (N_22109,N_21841,N_21828);
or U22110 (N_22110,N_21847,N_21792);
and U22111 (N_22111,N_21880,N_21914);
nand U22112 (N_22112,N_21941,N_21794);
xnor U22113 (N_22113,N_21887,N_21750);
nor U22114 (N_22114,N_21868,N_21760);
and U22115 (N_22115,N_21872,N_21928);
or U22116 (N_22116,N_21837,N_21977);
and U22117 (N_22117,N_21845,N_21865);
or U22118 (N_22118,N_21874,N_21827);
and U22119 (N_22119,N_21784,N_21810);
xor U22120 (N_22120,N_21808,N_21907);
and U22121 (N_22121,N_21781,N_21782);
nand U22122 (N_22122,N_21769,N_21787);
xnor U22123 (N_22123,N_21791,N_21802);
or U22124 (N_22124,N_21851,N_21953);
or U22125 (N_22125,N_21980,N_21901);
nand U22126 (N_22126,N_21895,N_21807);
nor U22127 (N_22127,N_21781,N_21901);
nand U22128 (N_22128,N_21885,N_21980);
or U22129 (N_22129,N_21818,N_21812);
and U22130 (N_22130,N_21989,N_21928);
and U22131 (N_22131,N_21845,N_21920);
or U22132 (N_22132,N_21887,N_21894);
nor U22133 (N_22133,N_21921,N_21792);
and U22134 (N_22134,N_21811,N_21920);
and U22135 (N_22135,N_21962,N_21904);
and U22136 (N_22136,N_21803,N_21794);
nor U22137 (N_22137,N_21845,N_21760);
or U22138 (N_22138,N_21859,N_21771);
xor U22139 (N_22139,N_21992,N_21840);
and U22140 (N_22140,N_21857,N_21852);
nor U22141 (N_22141,N_21757,N_21933);
or U22142 (N_22142,N_21938,N_21869);
and U22143 (N_22143,N_21966,N_21954);
xor U22144 (N_22144,N_21872,N_21815);
and U22145 (N_22145,N_21912,N_21937);
nand U22146 (N_22146,N_21976,N_21849);
or U22147 (N_22147,N_21941,N_21865);
and U22148 (N_22148,N_21969,N_21852);
or U22149 (N_22149,N_21785,N_21927);
nor U22150 (N_22150,N_21820,N_21916);
and U22151 (N_22151,N_21987,N_21855);
or U22152 (N_22152,N_21970,N_21997);
and U22153 (N_22153,N_21949,N_21982);
nand U22154 (N_22154,N_21764,N_21868);
and U22155 (N_22155,N_21886,N_21887);
nor U22156 (N_22156,N_21936,N_21813);
nand U22157 (N_22157,N_21866,N_21947);
or U22158 (N_22158,N_21920,N_21806);
nand U22159 (N_22159,N_21912,N_21905);
nor U22160 (N_22160,N_21852,N_21752);
and U22161 (N_22161,N_21846,N_21901);
and U22162 (N_22162,N_21993,N_21787);
and U22163 (N_22163,N_21827,N_21994);
nor U22164 (N_22164,N_21779,N_21841);
xnor U22165 (N_22165,N_21817,N_21756);
and U22166 (N_22166,N_21869,N_21902);
and U22167 (N_22167,N_21989,N_21765);
nand U22168 (N_22168,N_21915,N_21777);
or U22169 (N_22169,N_21825,N_21800);
or U22170 (N_22170,N_21884,N_21987);
or U22171 (N_22171,N_21830,N_21773);
nand U22172 (N_22172,N_21994,N_21953);
nor U22173 (N_22173,N_21803,N_21927);
and U22174 (N_22174,N_21915,N_21884);
or U22175 (N_22175,N_21956,N_21827);
xor U22176 (N_22176,N_21902,N_21833);
xnor U22177 (N_22177,N_21868,N_21978);
nand U22178 (N_22178,N_21859,N_21804);
and U22179 (N_22179,N_21762,N_21779);
nor U22180 (N_22180,N_21827,N_21876);
or U22181 (N_22181,N_21835,N_21995);
or U22182 (N_22182,N_21947,N_21901);
or U22183 (N_22183,N_21905,N_21965);
xor U22184 (N_22184,N_21828,N_21774);
nand U22185 (N_22185,N_21757,N_21905);
nor U22186 (N_22186,N_21873,N_21940);
xor U22187 (N_22187,N_21866,N_21790);
nor U22188 (N_22188,N_21993,N_21775);
and U22189 (N_22189,N_21988,N_21777);
or U22190 (N_22190,N_21880,N_21939);
nor U22191 (N_22191,N_21956,N_21800);
and U22192 (N_22192,N_21781,N_21884);
and U22193 (N_22193,N_21973,N_21894);
nand U22194 (N_22194,N_21800,N_21969);
nand U22195 (N_22195,N_21887,N_21939);
xor U22196 (N_22196,N_21934,N_21948);
or U22197 (N_22197,N_21986,N_21897);
or U22198 (N_22198,N_21788,N_21943);
and U22199 (N_22199,N_21791,N_21948);
xnor U22200 (N_22200,N_21947,N_21765);
nor U22201 (N_22201,N_21850,N_21988);
or U22202 (N_22202,N_21919,N_21926);
or U22203 (N_22203,N_21866,N_21906);
or U22204 (N_22204,N_21794,N_21809);
and U22205 (N_22205,N_21860,N_21856);
nand U22206 (N_22206,N_21896,N_21955);
nand U22207 (N_22207,N_21975,N_21954);
nand U22208 (N_22208,N_21935,N_21820);
and U22209 (N_22209,N_21820,N_21889);
and U22210 (N_22210,N_21753,N_21856);
nand U22211 (N_22211,N_21987,N_21813);
and U22212 (N_22212,N_21878,N_21818);
or U22213 (N_22213,N_21906,N_21804);
nand U22214 (N_22214,N_21847,N_21786);
nor U22215 (N_22215,N_21776,N_21930);
and U22216 (N_22216,N_21824,N_21960);
xor U22217 (N_22217,N_21933,N_21984);
nand U22218 (N_22218,N_21922,N_21840);
nor U22219 (N_22219,N_21916,N_21882);
or U22220 (N_22220,N_21775,N_21769);
or U22221 (N_22221,N_21851,N_21933);
nand U22222 (N_22222,N_21918,N_21912);
or U22223 (N_22223,N_21991,N_21891);
or U22224 (N_22224,N_21902,N_21960);
and U22225 (N_22225,N_21974,N_21901);
and U22226 (N_22226,N_21750,N_21923);
and U22227 (N_22227,N_21973,N_21844);
xnor U22228 (N_22228,N_21807,N_21769);
nor U22229 (N_22229,N_21807,N_21812);
and U22230 (N_22230,N_21848,N_21960);
nor U22231 (N_22231,N_21988,N_21820);
nand U22232 (N_22232,N_21810,N_21833);
xor U22233 (N_22233,N_21935,N_21999);
or U22234 (N_22234,N_21926,N_21969);
nand U22235 (N_22235,N_21821,N_21789);
or U22236 (N_22236,N_21957,N_21931);
or U22237 (N_22237,N_21943,N_21956);
nand U22238 (N_22238,N_21892,N_21778);
xnor U22239 (N_22239,N_21957,N_21971);
or U22240 (N_22240,N_21972,N_21966);
nor U22241 (N_22241,N_21924,N_21878);
xnor U22242 (N_22242,N_21894,N_21775);
or U22243 (N_22243,N_21840,N_21800);
or U22244 (N_22244,N_21830,N_21884);
xnor U22245 (N_22245,N_21904,N_21979);
xor U22246 (N_22246,N_21799,N_21984);
or U22247 (N_22247,N_21909,N_21762);
xor U22248 (N_22248,N_21787,N_21945);
or U22249 (N_22249,N_21887,N_21934);
or U22250 (N_22250,N_22031,N_22128);
nand U22251 (N_22251,N_22145,N_22037);
nor U22252 (N_22252,N_22046,N_22183);
nand U22253 (N_22253,N_22131,N_22245);
nand U22254 (N_22254,N_22074,N_22085);
xor U22255 (N_22255,N_22039,N_22162);
xnor U22256 (N_22256,N_22073,N_22076);
nor U22257 (N_22257,N_22099,N_22096);
or U22258 (N_22258,N_22088,N_22040);
nand U22259 (N_22259,N_22198,N_22056);
xnor U22260 (N_22260,N_22014,N_22208);
nand U22261 (N_22261,N_22120,N_22024);
nand U22262 (N_22262,N_22036,N_22100);
or U22263 (N_22263,N_22147,N_22050);
and U22264 (N_22264,N_22227,N_22214);
xnor U22265 (N_22265,N_22166,N_22155);
nand U22266 (N_22266,N_22029,N_22055);
and U22267 (N_22267,N_22243,N_22034);
nand U22268 (N_22268,N_22028,N_22143);
nand U22269 (N_22269,N_22038,N_22080);
nor U22270 (N_22270,N_22215,N_22157);
nor U22271 (N_22271,N_22044,N_22236);
nand U22272 (N_22272,N_22090,N_22079);
nor U22273 (N_22273,N_22216,N_22149);
or U22274 (N_22274,N_22141,N_22247);
xor U22275 (N_22275,N_22191,N_22204);
and U22276 (N_22276,N_22212,N_22209);
nand U22277 (N_22277,N_22144,N_22093);
nor U22278 (N_22278,N_22150,N_22153);
or U22279 (N_22279,N_22118,N_22207);
or U22280 (N_22280,N_22121,N_22152);
xor U22281 (N_22281,N_22222,N_22065);
nor U22282 (N_22282,N_22070,N_22217);
or U22283 (N_22283,N_22159,N_22167);
nor U22284 (N_22284,N_22160,N_22242);
xnor U22285 (N_22285,N_22221,N_22027);
nor U22286 (N_22286,N_22184,N_22091);
nor U22287 (N_22287,N_22061,N_22016);
or U22288 (N_22288,N_22195,N_22101);
nor U22289 (N_22289,N_22219,N_22084);
and U22290 (N_22290,N_22023,N_22108);
nand U22291 (N_22291,N_22220,N_22043);
nand U22292 (N_22292,N_22064,N_22241);
xor U22293 (N_22293,N_22114,N_22103);
nand U22294 (N_22294,N_22051,N_22169);
nand U22295 (N_22295,N_22164,N_22122);
or U22296 (N_22296,N_22098,N_22146);
nor U22297 (N_22297,N_22110,N_22087);
or U22298 (N_22298,N_22201,N_22186);
xor U22299 (N_22299,N_22097,N_22246);
or U22300 (N_22300,N_22053,N_22178);
or U22301 (N_22301,N_22134,N_22190);
xnor U22302 (N_22302,N_22229,N_22199);
or U22303 (N_22303,N_22000,N_22062);
nor U22304 (N_22304,N_22127,N_22094);
nand U22305 (N_22305,N_22136,N_22235);
or U22306 (N_22306,N_22017,N_22116);
and U22307 (N_22307,N_22193,N_22007);
and U22308 (N_22308,N_22197,N_22081);
nand U22309 (N_22309,N_22185,N_22058);
and U22310 (N_22310,N_22225,N_22068);
nand U22311 (N_22311,N_22192,N_22135);
xnor U22312 (N_22312,N_22111,N_22211);
or U22313 (N_22313,N_22172,N_22086);
xor U22314 (N_22314,N_22196,N_22168);
nand U22315 (N_22315,N_22206,N_22106);
nor U22316 (N_22316,N_22181,N_22200);
and U22317 (N_22317,N_22239,N_22138);
nand U22318 (N_22318,N_22018,N_22026);
and U22319 (N_22319,N_22182,N_22148);
nand U22320 (N_22320,N_22011,N_22123);
and U22321 (N_22321,N_22112,N_22170);
nor U22322 (N_22322,N_22226,N_22077);
nor U22323 (N_22323,N_22041,N_22234);
and U22324 (N_22324,N_22004,N_22047);
and U22325 (N_22325,N_22105,N_22066);
or U22326 (N_22326,N_22042,N_22012);
nor U22327 (N_22327,N_22237,N_22248);
nor U22328 (N_22328,N_22161,N_22109);
xor U22329 (N_22329,N_22140,N_22060);
and U22330 (N_22330,N_22132,N_22228);
or U22331 (N_22331,N_22163,N_22231);
or U22332 (N_22332,N_22224,N_22035);
and U22333 (N_22333,N_22057,N_22188);
nand U22334 (N_22334,N_22151,N_22249);
nand U22335 (N_22335,N_22173,N_22069);
nand U22336 (N_22336,N_22001,N_22133);
xor U22337 (N_22337,N_22119,N_22213);
or U22338 (N_22338,N_22015,N_22022);
nand U22339 (N_22339,N_22075,N_22154);
and U22340 (N_22340,N_22071,N_22002);
nand U22341 (N_22341,N_22082,N_22019);
xor U22342 (N_22342,N_22189,N_22020);
or U22343 (N_22343,N_22223,N_22115);
or U22344 (N_22344,N_22139,N_22045);
xnor U22345 (N_22345,N_22092,N_22156);
nand U22346 (N_22346,N_22180,N_22124);
nor U22347 (N_22347,N_22104,N_22063);
or U22348 (N_22348,N_22078,N_22194);
and U22349 (N_22349,N_22003,N_22175);
and U22350 (N_22350,N_22032,N_22025);
nor U22351 (N_22351,N_22126,N_22052);
or U22352 (N_22352,N_22010,N_22205);
xnor U22353 (N_22353,N_22240,N_22171);
xor U22354 (N_22354,N_22059,N_22244);
nor U22355 (N_22355,N_22202,N_22067);
and U22356 (N_22356,N_22083,N_22006);
nand U22357 (N_22357,N_22218,N_22117);
and U22358 (N_22358,N_22177,N_22107);
or U22359 (N_22359,N_22158,N_22009);
and U22360 (N_22360,N_22089,N_22049);
nand U22361 (N_22361,N_22232,N_22233);
xnor U22362 (N_22362,N_22008,N_22179);
or U22363 (N_22363,N_22102,N_22142);
and U22364 (N_22364,N_22203,N_22048);
nor U22365 (N_22365,N_22021,N_22113);
nand U22366 (N_22366,N_22230,N_22165);
nor U22367 (N_22367,N_22210,N_22129);
and U22368 (N_22368,N_22030,N_22187);
xnor U22369 (N_22369,N_22137,N_22130);
xnor U22370 (N_22370,N_22033,N_22238);
and U22371 (N_22371,N_22095,N_22005);
and U22372 (N_22372,N_22013,N_22072);
nand U22373 (N_22373,N_22125,N_22176);
nor U22374 (N_22374,N_22174,N_22054);
xnor U22375 (N_22375,N_22135,N_22196);
and U22376 (N_22376,N_22245,N_22246);
xor U22377 (N_22377,N_22052,N_22067);
and U22378 (N_22378,N_22226,N_22225);
xnor U22379 (N_22379,N_22128,N_22214);
xor U22380 (N_22380,N_22147,N_22141);
and U22381 (N_22381,N_22229,N_22141);
nor U22382 (N_22382,N_22124,N_22184);
nor U22383 (N_22383,N_22019,N_22071);
nor U22384 (N_22384,N_22040,N_22016);
or U22385 (N_22385,N_22241,N_22010);
and U22386 (N_22386,N_22018,N_22191);
or U22387 (N_22387,N_22156,N_22122);
nor U22388 (N_22388,N_22203,N_22236);
xor U22389 (N_22389,N_22107,N_22034);
nor U22390 (N_22390,N_22216,N_22199);
or U22391 (N_22391,N_22126,N_22222);
xnor U22392 (N_22392,N_22086,N_22019);
or U22393 (N_22393,N_22114,N_22198);
nor U22394 (N_22394,N_22045,N_22065);
nor U22395 (N_22395,N_22224,N_22213);
nor U22396 (N_22396,N_22078,N_22177);
and U22397 (N_22397,N_22104,N_22107);
nand U22398 (N_22398,N_22000,N_22143);
or U22399 (N_22399,N_22089,N_22051);
and U22400 (N_22400,N_22026,N_22163);
and U22401 (N_22401,N_22225,N_22054);
and U22402 (N_22402,N_22123,N_22234);
nand U22403 (N_22403,N_22237,N_22022);
or U22404 (N_22404,N_22023,N_22020);
or U22405 (N_22405,N_22228,N_22180);
nand U22406 (N_22406,N_22003,N_22244);
nor U22407 (N_22407,N_22062,N_22089);
or U22408 (N_22408,N_22249,N_22065);
or U22409 (N_22409,N_22051,N_22154);
or U22410 (N_22410,N_22209,N_22126);
xnor U22411 (N_22411,N_22182,N_22013);
xnor U22412 (N_22412,N_22058,N_22182);
and U22413 (N_22413,N_22006,N_22221);
and U22414 (N_22414,N_22226,N_22043);
xnor U22415 (N_22415,N_22233,N_22110);
nand U22416 (N_22416,N_22238,N_22226);
xor U22417 (N_22417,N_22071,N_22091);
nor U22418 (N_22418,N_22018,N_22017);
and U22419 (N_22419,N_22048,N_22010);
nand U22420 (N_22420,N_22246,N_22238);
nand U22421 (N_22421,N_22015,N_22137);
and U22422 (N_22422,N_22084,N_22210);
xnor U22423 (N_22423,N_22060,N_22169);
or U22424 (N_22424,N_22199,N_22065);
and U22425 (N_22425,N_22110,N_22248);
or U22426 (N_22426,N_22142,N_22133);
nand U22427 (N_22427,N_22207,N_22034);
nor U22428 (N_22428,N_22007,N_22036);
and U22429 (N_22429,N_22092,N_22124);
and U22430 (N_22430,N_22119,N_22129);
and U22431 (N_22431,N_22078,N_22233);
and U22432 (N_22432,N_22090,N_22192);
nor U22433 (N_22433,N_22032,N_22197);
nand U22434 (N_22434,N_22101,N_22115);
nand U22435 (N_22435,N_22164,N_22206);
or U22436 (N_22436,N_22091,N_22083);
and U22437 (N_22437,N_22175,N_22207);
xor U22438 (N_22438,N_22114,N_22132);
or U22439 (N_22439,N_22113,N_22119);
or U22440 (N_22440,N_22156,N_22147);
and U22441 (N_22441,N_22056,N_22234);
nor U22442 (N_22442,N_22175,N_22019);
xor U22443 (N_22443,N_22109,N_22103);
nand U22444 (N_22444,N_22041,N_22203);
nor U22445 (N_22445,N_22223,N_22145);
or U22446 (N_22446,N_22140,N_22129);
nand U22447 (N_22447,N_22221,N_22110);
and U22448 (N_22448,N_22119,N_22080);
and U22449 (N_22449,N_22091,N_22057);
xor U22450 (N_22450,N_22108,N_22152);
xnor U22451 (N_22451,N_22041,N_22168);
and U22452 (N_22452,N_22176,N_22097);
xor U22453 (N_22453,N_22007,N_22234);
or U22454 (N_22454,N_22000,N_22006);
xor U22455 (N_22455,N_22105,N_22028);
and U22456 (N_22456,N_22103,N_22118);
or U22457 (N_22457,N_22201,N_22003);
and U22458 (N_22458,N_22228,N_22027);
or U22459 (N_22459,N_22247,N_22013);
or U22460 (N_22460,N_22163,N_22021);
nand U22461 (N_22461,N_22233,N_22021);
or U22462 (N_22462,N_22216,N_22237);
and U22463 (N_22463,N_22209,N_22032);
nand U22464 (N_22464,N_22112,N_22226);
xnor U22465 (N_22465,N_22207,N_22006);
and U22466 (N_22466,N_22000,N_22024);
and U22467 (N_22467,N_22088,N_22164);
nor U22468 (N_22468,N_22203,N_22227);
nand U22469 (N_22469,N_22179,N_22248);
xnor U22470 (N_22470,N_22004,N_22221);
xor U22471 (N_22471,N_22005,N_22108);
xor U22472 (N_22472,N_22164,N_22190);
nand U22473 (N_22473,N_22171,N_22044);
nor U22474 (N_22474,N_22180,N_22201);
or U22475 (N_22475,N_22217,N_22234);
nand U22476 (N_22476,N_22147,N_22051);
or U22477 (N_22477,N_22031,N_22129);
and U22478 (N_22478,N_22182,N_22175);
nor U22479 (N_22479,N_22091,N_22216);
xor U22480 (N_22480,N_22144,N_22194);
xnor U22481 (N_22481,N_22031,N_22107);
or U22482 (N_22482,N_22031,N_22211);
xnor U22483 (N_22483,N_22076,N_22175);
and U22484 (N_22484,N_22054,N_22049);
and U22485 (N_22485,N_22195,N_22077);
and U22486 (N_22486,N_22018,N_22200);
nand U22487 (N_22487,N_22229,N_22066);
xor U22488 (N_22488,N_22188,N_22240);
or U22489 (N_22489,N_22058,N_22008);
and U22490 (N_22490,N_22117,N_22137);
nand U22491 (N_22491,N_22175,N_22068);
nor U22492 (N_22492,N_22111,N_22057);
nor U22493 (N_22493,N_22057,N_22162);
nand U22494 (N_22494,N_22115,N_22249);
and U22495 (N_22495,N_22036,N_22197);
and U22496 (N_22496,N_22060,N_22101);
xor U22497 (N_22497,N_22213,N_22135);
nor U22498 (N_22498,N_22064,N_22117);
nand U22499 (N_22499,N_22144,N_22235);
nor U22500 (N_22500,N_22345,N_22335);
nor U22501 (N_22501,N_22361,N_22250);
nand U22502 (N_22502,N_22397,N_22492);
nor U22503 (N_22503,N_22466,N_22256);
or U22504 (N_22504,N_22385,N_22367);
nand U22505 (N_22505,N_22273,N_22368);
and U22506 (N_22506,N_22482,N_22452);
or U22507 (N_22507,N_22423,N_22262);
nor U22508 (N_22508,N_22371,N_22438);
nor U22509 (N_22509,N_22344,N_22359);
nor U22510 (N_22510,N_22447,N_22319);
and U22511 (N_22511,N_22356,N_22263);
nand U22512 (N_22512,N_22471,N_22360);
nand U22513 (N_22513,N_22404,N_22310);
nand U22514 (N_22514,N_22324,N_22464);
nor U22515 (N_22515,N_22257,N_22472);
or U22516 (N_22516,N_22435,N_22389);
nor U22517 (N_22517,N_22469,N_22354);
xor U22518 (N_22518,N_22275,N_22362);
or U22519 (N_22519,N_22421,N_22496);
nor U22520 (N_22520,N_22462,N_22425);
nand U22521 (N_22521,N_22413,N_22346);
or U22522 (N_22522,N_22475,N_22430);
xor U22523 (N_22523,N_22432,N_22280);
nand U22524 (N_22524,N_22429,N_22331);
or U22525 (N_22525,N_22486,N_22443);
nand U22526 (N_22526,N_22392,N_22308);
xnor U22527 (N_22527,N_22488,N_22405);
xor U22528 (N_22528,N_22293,N_22406);
nand U22529 (N_22529,N_22409,N_22291);
nand U22530 (N_22530,N_22304,N_22382);
or U22531 (N_22531,N_22266,N_22480);
and U22532 (N_22532,N_22441,N_22408);
or U22533 (N_22533,N_22463,N_22440);
or U22534 (N_22534,N_22289,N_22267);
nor U22535 (N_22535,N_22288,N_22305);
nand U22536 (N_22536,N_22399,N_22270);
or U22537 (N_22537,N_22459,N_22387);
nand U22538 (N_22538,N_22370,N_22316);
or U22539 (N_22539,N_22332,N_22450);
or U22540 (N_22540,N_22442,N_22251);
xor U22541 (N_22541,N_22414,N_22325);
nor U22542 (N_22542,N_22272,N_22278);
nor U22543 (N_22543,N_22285,N_22436);
nand U22544 (N_22544,N_22393,N_22449);
nand U22545 (N_22545,N_22254,N_22470);
xor U22546 (N_22546,N_22300,N_22333);
nand U22547 (N_22547,N_22295,N_22372);
and U22548 (N_22548,N_22252,N_22313);
or U22549 (N_22549,N_22473,N_22411);
or U22550 (N_22550,N_22468,N_22255);
nor U22551 (N_22551,N_22365,N_22461);
nand U22552 (N_22552,N_22339,N_22376);
xor U22553 (N_22553,N_22437,N_22302);
nand U22554 (N_22554,N_22327,N_22342);
or U22555 (N_22555,N_22297,N_22259);
xnor U22556 (N_22556,N_22444,N_22315);
or U22557 (N_22557,N_22424,N_22498);
nand U22558 (N_22558,N_22374,N_22484);
and U22559 (N_22559,N_22433,N_22321);
or U22560 (N_22560,N_22326,N_22446);
nand U22561 (N_22561,N_22329,N_22298);
nand U22562 (N_22562,N_22428,N_22373);
nand U22563 (N_22563,N_22350,N_22296);
xnor U22564 (N_22564,N_22363,N_22261);
or U22565 (N_22565,N_22476,N_22290);
and U22566 (N_22566,N_22448,N_22276);
and U22567 (N_22567,N_22301,N_22391);
nand U22568 (N_22568,N_22268,N_22318);
nand U22569 (N_22569,N_22403,N_22400);
or U22570 (N_22570,N_22264,N_22284);
nor U22571 (N_22571,N_22322,N_22456);
nand U22572 (N_22572,N_22282,N_22306);
xnor U22573 (N_22573,N_22422,N_22292);
xor U22574 (N_22574,N_22426,N_22402);
nand U22575 (N_22575,N_22269,N_22351);
nor U22576 (N_22576,N_22481,N_22348);
and U22577 (N_22577,N_22353,N_22383);
nand U22578 (N_22578,N_22401,N_22253);
xnor U22579 (N_22579,N_22380,N_22330);
and U22580 (N_22580,N_22418,N_22491);
nand U22581 (N_22581,N_22467,N_22479);
nor U22582 (N_22582,N_22341,N_22489);
xnor U22583 (N_22583,N_22485,N_22460);
nor U22584 (N_22584,N_22303,N_22309);
xnor U22585 (N_22585,N_22455,N_22317);
nand U22586 (N_22586,N_22271,N_22357);
xor U22587 (N_22587,N_22258,N_22415);
xnor U22588 (N_22588,N_22337,N_22299);
or U22589 (N_22589,N_22390,N_22323);
xnor U22590 (N_22590,N_22427,N_22458);
nand U22591 (N_22591,N_22343,N_22445);
nand U22592 (N_22592,N_22260,N_22494);
xor U22593 (N_22593,N_22474,N_22386);
nor U22594 (N_22594,N_22396,N_22388);
and U22595 (N_22595,N_22294,N_22265);
or U22596 (N_22596,N_22287,N_22487);
nor U22597 (N_22597,N_22434,N_22311);
nor U22598 (N_22598,N_22328,N_22431);
and U22599 (N_22599,N_22477,N_22465);
and U22600 (N_22600,N_22381,N_22274);
and U22601 (N_22601,N_22349,N_22495);
nor U22602 (N_22602,N_22307,N_22394);
nor U22603 (N_22603,N_22395,N_22281);
nand U22604 (N_22604,N_22410,N_22369);
xnor U22605 (N_22605,N_22412,N_22453);
nor U22606 (N_22606,N_22352,N_22417);
xnor U22607 (N_22607,N_22366,N_22375);
xor U22608 (N_22608,N_22419,N_22499);
nor U22609 (N_22609,N_22312,N_22483);
xnor U22610 (N_22610,N_22379,N_22407);
nand U22611 (N_22611,N_22378,N_22355);
nand U22612 (N_22612,N_22358,N_22497);
or U22613 (N_22613,N_22364,N_22286);
nor U22614 (N_22614,N_22454,N_22493);
and U22615 (N_22615,N_22277,N_22377);
nor U22616 (N_22616,N_22416,N_22457);
or U22617 (N_22617,N_22336,N_22398);
and U22618 (N_22618,N_22279,N_22420);
nor U22619 (N_22619,N_22347,N_22334);
and U22620 (N_22620,N_22340,N_22314);
xor U22621 (N_22621,N_22338,N_22451);
xnor U22622 (N_22622,N_22439,N_22490);
and U22623 (N_22623,N_22320,N_22384);
nand U22624 (N_22624,N_22283,N_22478);
xnor U22625 (N_22625,N_22371,N_22318);
nor U22626 (N_22626,N_22429,N_22358);
xor U22627 (N_22627,N_22441,N_22493);
or U22628 (N_22628,N_22295,N_22478);
nand U22629 (N_22629,N_22307,N_22496);
or U22630 (N_22630,N_22272,N_22437);
xor U22631 (N_22631,N_22270,N_22273);
nor U22632 (N_22632,N_22475,N_22303);
nor U22633 (N_22633,N_22369,N_22399);
nor U22634 (N_22634,N_22291,N_22426);
nor U22635 (N_22635,N_22253,N_22438);
and U22636 (N_22636,N_22367,N_22474);
nand U22637 (N_22637,N_22379,N_22499);
or U22638 (N_22638,N_22475,N_22349);
nor U22639 (N_22639,N_22299,N_22261);
nor U22640 (N_22640,N_22336,N_22429);
nor U22641 (N_22641,N_22421,N_22312);
xor U22642 (N_22642,N_22293,N_22350);
and U22643 (N_22643,N_22288,N_22271);
and U22644 (N_22644,N_22374,N_22367);
or U22645 (N_22645,N_22359,N_22435);
and U22646 (N_22646,N_22302,N_22327);
nand U22647 (N_22647,N_22452,N_22342);
or U22648 (N_22648,N_22354,N_22305);
nand U22649 (N_22649,N_22336,N_22459);
nor U22650 (N_22650,N_22404,N_22333);
and U22651 (N_22651,N_22412,N_22488);
and U22652 (N_22652,N_22431,N_22497);
or U22653 (N_22653,N_22334,N_22443);
nor U22654 (N_22654,N_22374,N_22441);
xor U22655 (N_22655,N_22378,N_22312);
and U22656 (N_22656,N_22386,N_22376);
nor U22657 (N_22657,N_22397,N_22267);
nand U22658 (N_22658,N_22386,N_22338);
and U22659 (N_22659,N_22253,N_22373);
and U22660 (N_22660,N_22299,N_22428);
or U22661 (N_22661,N_22321,N_22460);
and U22662 (N_22662,N_22368,N_22412);
or U22663 (N_22663,N_22499,N_22475);
nor U22664 (N_22664,N_22352,N_22438);
nand U22665 (N_22665,N_22470,N_22349);
xnor U22666 (N_22666,N_22433,N_22259);
nor U22667 (N_22667,N_22322,N_22487);
nand U22668 (N_22668,N_22488,N_22348);
or U22669 (N_22669,N_22282,N_22374);
or U22670 (N_22670,N_22385,N_22448);
xnor U22671 (N_22671,N_22329,N_22363);
xor U22672 (N_22672,N_22368,N_22365);
nor U22673 (N_22673,N_22399,N_22420);
xor U22674 (N_22674,N_22473,N_22443);
xor U22675 (N_22675,N_22279,N_22391);
nand U22676 (N_22676,N_22369,N_22474);
nor U22677 (N_22677,N_22474,N_22296);
and U22678 (N_22678,N_22486,N_22290);
nor U22679 (N_22679,N_22462,N_22457);
nor U22680 (N_22680,N_22433,N_22307);
nor U22681 (N_22681,N_22458,N_22251);
nor U22682 (N_22682,N_22404,N_22312);
and U22683 (N_22683,N_22404,N_22309);
xor U22684 (N_22684,N_22405,N_22275);
and U22685 (N_22685,N_22279,N_22340);
nor U22686 (N_22686,N_22344,N_22393);
nor U22687 (N_22687,N_22490,N_22325);
and U22688 (N_22688,N_22285,N_22304);
and U22689 (N_22689,N_22312,N_22376);
nand U22690 (N_22690,N_22372,N_22349);
nor U22691 (N_22691,N_22263,N_22363);
or U22692 (N_22692,N_22416,N_22469);
xnor U22693 (N_22693,N_22458,N_22307);
nor U22694 (N_22694,N_22263,N_22257);
xor U22695 (N_22695,N_22492,N_22405);
nor U22696 (N_22696,N_22376,N_22347);
or U22697 (N_22697,N_22256,N_22373);
and U22698 (N_22698,N_22411,N_22389);
or U22699 (N_22699,N_22449,N_22405);
or U22700 (N_22700,N_22316,N_22265);
xor U22701 (N_22701,N_22315,N_22337);
nand U22702 (N_22702,N_22419,N_22310);
or U22703 (N_22703,N_22281,N_22280);
nand U22704 (N_22704,N_22439,N_22329);
nand U22705 (N_22705,N_22464,N_22407);
and U22706 (N_22706,N_22387,N_22274);
and U22707 (N_22707,N_22361,N_22263);
or U22708 (N_22708,N_22370,N_22339);
or U22709 (N_22709,N_22385,N_22321);
and U22710 (N_22710,N_22375,N_22389);
nor U22711 (N_22711,N_22362,N_22353);
and U22712 (N_22712,N_22339,N_22408);
xnor U22713 (N_22713,N_22317,N_22373);
or U22714 (N_22714,N_22309,N_22386);
and U22715 (N_22715,N_22408,N_22426);
nor U22716 (N_22716,N_22459,N_22494);
or U22717 (N_22717,N_22360,N_22449);
xor U22718 (N_22718,N_22446,N_22313);
or U22719 (N_22719,N_22332,N_22415);
and U22720 (N_22720,N_22286,N_22456);
nor U22721 (N_22721,N_22380,N_22314);
or U22722 (N_22722,N_22357,N_22446);
nand U22723 (N_22723,N_22389,N_22349);
xor U22724 (N_22724,N_22378,N_22352);
nor U22725 (N_22725,N_22350,N_22481);
and U22726 (N_22726,N_22333,N_22481);
or U22727 (N_22727,N_22368,N_22307);
and U22728 (N_22728,N_22371,N_22345);
xor U22729 (N_22729,N_22274,N_22438);
nand U22730 (N_22730,N_22294,N_22368);
nor U22731 (N_22731,N_22457,N_22403);
nand U22732 (N_22732,N_22480,N_22462);
xor U22733 (N_22733,N_22475,N_22272);
or U22734 (N_22734,N_22350,N_22397);
nand U22735 (N_22735,N_22465,N_22310);
xor U22736 (N_22736,N_22494,N_22273);
or U22737 (N_22737,N_22319,N_22409);
xor U22738 (N_22738,N_22436,N_22318);
nand U22739 (N_22739,N_22435,N_22280);
nor U22740 (N_22740,N_22455,N_22440);
nor U22741 (N_22741,N_22406,N_22326);
or U22742 (N_22742,N_22310,N_22374);
nor U22743 (N_22743,N_22297,N_22452);
nor U22744 (N_22744,N_22369,N_22279);
nor U22745 (N_22745,N_22334,N_22261);
xnor U22746 (N_22746,N_22295,N_22269);
and U22747 (N_22747,N_22309,N_22306);
or U22748 (N_22748,N_22423,N_22449);
and U22749 (N_22749,N_22495,N_22303);
or U22750 (N_22750,N_22622,N_22716);
and U22751 (N_22751,N_22693,N_22655);
nor U22752 (N_22752,N_22729,N_22703);
and U22753 (N_22753,N_22651,N_22713);
nor U22754 (N_22754,N_22584,N_22510);
or U22755 (N_22755,N_22726,N_22678);
nor U22756 (N_22756,N_22530,N_22691);
nor U22757 (N_22757,N_22748,N_22677);
or U22758 (N_22758,N_22562,N_22537);
nand U22759 (N_22759,N_22502,N_22709);
xnor U22760 (N_22760,N_22558,N_22632);
nor U22761 (N_22761,N_22590,N_22598);
and U22762 (N_22762,N_22675,N_22565);
and U22763 (N_22763,N_22612,N_22711);
or U22764 (N_22764,N_22659,N_22582);
nor U22765 (N_22765,N_22564,N_22626);
nor U22766 (N_22766,N_22557,N_22734);
and U22767 (N_22767,N_22513,N_22695);
xor U22768 (N_22768,N_22700,N_22618);
and U22769 (N_22769,N_22610,N_22587);
nor U22770 (N_22770,N_22597,N_22721);
xnor U22771 (N_22771,N_22657,N_22527);
or U22772 (N_22772,N_22544,N_22615);
or U22773 (N_22773,N_22560,N_22525);
and U22774 (N_22774,N_22600,N_22681);
nor U22775 (N_22775,N_22717,N_22634);
or U22776 (N_22776,N_22572,N_22629);
and U22777 (N_22777,N_22722,N_22539);
and U22778 (N_22778,N_22742,N_22672);
and U22779 (N_22779,N_22563,N_22633);
nor U22780 (N_22780,N_22535,N_22674);
and U22781 (N_22781,N_22686,N_22676);
or U22782 (N_22782,N_22715,N_22736);
or U22783 (N_22783,N_22723,N_22611);
xor U22784 (N_22784,N_22714,N_22624);
or U22785 (N_22785,N_22708,N_22706);
nor U22786 (N_22786,N_22650,N_22641);
and U22787 (N_22787,N_22712,N_22556);
xor U22788 (N_22788,N_22500,N_22570);
xor U22789 (N_22789,N_22546,N_22662);
nand U22790 (N_22790,N_22550,N_22620);
and U22791 (N_22791,N_22749,N_22621);
xor U22792 (N_22792,N_22566,N_22517);
or U22793 (N_22793,N_22534,N_22707);
and U22794 (N_22794,N_22648,N_22553);
nand U22795 (N_22795,N_22652,N_22705);
nor U22796 (N_22796,N_22595,N_22545);
and U22797 (N_22797,N_22561,N_22653);
xor U22798 (N_22798,N_22719,N_22506);
or U22799 (N_22799,N_22580,N_22586);
nand U22800 (N_22800,N_22540,N_22746);
nor U22801 (N_22801,N_22609,N_22606);
xor U22802 (N_22802,N_22614,N_22669);
nand U22803 (N_22803,N_22528,N_22636);
nand U22804 (N_22804,N_22581,N_22520);
or U22805 (N_22805,N_22745,N_22735);
xor U22806 (N_22806,N_22568,N_22668);
and U22807 (N_22807,N_22623,N_22656);
nand U22808 (N_22808,N_22688,N_22727);
nand U22809 (N_22809,N_22603,N_22596);
and U22810 (N_22810,N_22720,N_22730);
xnor U22811 (N_22811,N_22543,N_22601);
nand U22812 (N_22812,N_22532,N_22683);
and U22813 (N_22813,N_22733,N_22680);
nand U22814 (N_22814,N_22747,N_22725);
and U22815 (N_22815,N_22607,N_22679);
xnor U22816 (N_22816,N_22646,N_22697);
and U22817 (N_22817,N_22744,N_22661);
and U22818 (N_22818,N_22531,N_22739);
and U22819 (N_22819,N_22696,N_22718);
and U22820 (N_22820,N_22567,N_22670);
nor U22821 (N_22821,N_22664,N_22536);
xnor U22822 (N_22822,N_22549,N_22710);
nand U22823 (N_22823,N_22640,N_22645);
or U22824 (N_22824,N_22740,N_22616);
or U22825 (N_22825,N_22699,N_22635);
or U22826 (N_22826,N_22613,N_22591);
or U22827 (N_22827,N_22728,N_22523);
xnor U22828 (N_22828,N_22559,N_22701);
nand U22829 (N_22829,N_22724,N_22663);
or U22830 (N_22830,N_22516,N_22605);
or U22831 (N_22831,N_22522,N_22512);
or U22832 (N_22832,N_22643,N_22619);
xnor U22833 (N_22833,N_22658,N_22524);
or U22834 (N_22834,N_22538,N_22519);
and U22835 (N_22835,N_22630,N_22573);
xnor U22836 (N_22836,N_22576,N_22660);
nor U22837 (N_22837,N_22731,N_22667);
nand U22838 (N_22838,N_22589,N_22687);
xor U22839 (N_22839,N_22503,N_22583);
xor U22840 (N_22840,N_22533,N_22738);
and U22841 (N_22841,N_22666,N_22585);
and U22842 (N_22842,N_22508,N_22594);
xnor U22843 (N_22843,N_22644,N_22698);
nand U22844 (N_22844,N_22637,N_22617);
nor U22845 (N_22845,N_22608,N_22505);
or U22846 (N_22846,N_22593,N_22518);
and U22847 (N_22847,N_22592,N_22665);
or U22848 (N_22848,N_22682,N_22509);
nand U22849 (N_22849,N_22654,N_22599);
or U22850 (N_22850,N_22604,N_22542);
or U22851 (N_22851,N_22689,N_22547);
xor U22852 (N_22852,N_22673,N_22692);
or U22853 (N_22853,N_22526,N_22515);
nor U22854 (N_22854,N_22552,N_22504);
nor U22855 (N_22855,N_22511,N_22529);
nand U22856 (N_22856,N_22602,N_22694);
nor U22857 (N_22857,N_22571,N_22627);
nor U22858 (N_22858,N_22514,N_22541);
or U22859 (N_22859,N_22578,N_22649);
and U22860 (N_22860,N_22684,N_22507);
xor U22861 (N_22861,N_22690,N_22577);
and U22862 (N_22862,N_22741,N_22625);
xor U22863 (N_22863,N_22569,N_22642);
nand U22864 (N_22864,N_22574,N_22638);
nor U22865 (N_22865,N_22647,N_22628);
nand U22866 (N_22866,N_22579,N_22671);
nand U22867 (N_22867,N_22743,N_22555);
and U22868 (N_22868,N_22501,N_22631);
xnor U22869 (N_22869,N_22554,N_22521);
xnor U22870 (N_22870,N_22702,N_22737);
nand U22871 (N_22871,N_22551,N_22639);
nand U22872 (N_22872,N_22704,N_22732);
xnor U22873 (N_22873,N_22588,N_22575);
or U22874 (N_22874,N_22685,N_22548);
and U22875 (N_22875,N_22591,N_22656);
nand U22876 (N_22876,N_22666,N_22641);
and U22877 (N_22877,N_22519,N_22598);
or U22878 (N_22878,N_22660,N_22538);
nand U22879 (N_22879,N_22657,N_22554);
nor U22880 (N_22880,N_22553,N_22685);
nor U22881 (N_22881,N_22717,N_22578);
nand U22882 (N_22882,N_22634,N_22722);
and U22883 (N_22883,N_22569,N_22681);
and U22884 (N_22884,N_22546,N_22718);
nor U22885 (N_22885,N_22646,N_22598);
and U22886 (N_22886,N_22514,N_22605);
nand U22887 (N_22887,N_22685,N_22672);
or U22888 (N_22888,N_22596,N_22694);
xor U22889 (N_22889,N_22639,N_22742);
nor U22890 (N_22890,N_22743,N_22717);
or U22891 (N_22891,N_22730,N_22649);
xnor U22892 (N_22892,N_22659,N_22621);
nor U22893 (N_22893,N_22626,N_22516);
xor U22894 (N_22894,N_22663,N_22744);
and U22895 (N_22895,N_22600,N_22561);
nor U22896 (N_22896,N_22711,N_22638);
and U22897 (N_22897,N_22682,N_22681);
nand U22898 (N_22898,N_22663,N_22691);
xor U22899 (N_22899,N_22516,N_22707);
xor U22900 (N_22900,N_22533,N_22695);
and U22901 (N_22901,N_22616,N_22666);
nand U22902 (N_22902,N_22747,N_22517);
nor U22903 (N_22903,N_22697,N_22530);
and U22904 (N_22904,N_22591,N_22539);
and U22905 (N_22905,N_22592,N_22630);
and U22906 (N_22906,N_22542,N_22728);
nor U22907 (N_22907,N_22507,N_22745);
or U22908 (N_22908,N_22710,N_22558);
or U22909 (N_22909,N_22652,N_22728);
nand U22910 (N_22910,N_22719,N_22501);
nor U22911 (N_22911,N_22505,N_22684);
xnor U22912 (N_22912,N_22546,N_22675);
and U22913 (N_22913,N_22688,N_22574);
xnor U22914 (N_22914,N_22615,N_22682);
nor U22915 (N_22915,N_22600,N_22574);
nor U22916 (N_22916,N_22533,N_22598);
or U22917 (N_22917,N_22631,N_22523);
or U22918 (N_22918,N_22554,N_22673);
and U22919 (N_22919,N_22695,N_22742);
xnor U22920 (N_22920,N_22640,N_22604);
nand U22921 (N_22921,N_22571,N_22691);
nor U22922 (N_22922,N_22527,N_22740);
and U22923 (N_22923,N_22678,N_22539);
xor U22924 (N_22924,N_22535,N_22554);
and U22925 (N_22925,N_22739,N_22702);
and U22926 (N_22926,N_22617,N_22725);
or U22927 (N_22927,N_22586,N_22540);
nand U22928 (N_22928,N_22557,N_22616);
or U22929 (N_22929,N_22625,N_22710);
or U22930 (N_22930,N_22711,N_22581);
xnor U22931 (N_22931,N_22557,N_22662);
xor U22932 (N_22932,N_22614,N_22566);
nor U22933 (N_22933,N_22703,N_22648);
or U22934 (N_22934,N_22728,N_22642);
nand U22935 (N_22935,N_22662,N_22672);
xor U22936 (N_22936,N_22559,N_22537);
or U22937 (N_22937,N_22736,N_22644);
or U22938 (N_22938,N_22571,N_22567);
xor U22939 (N_22939,N_22581,N_22715);
xnor U22940 (N_22940,N_22629,N_22720);
or U22941 (N_22941,N_22595,N_22680);
nand U22942 (N_22942,N_22703,N_22742);
nor U22943 (N_22943,N_22599,N_22583);
nor U22944 (N_22944,N_22611,N_22657);
nor U22945 (N_22945,N_22705,N_22695);
and U22946 (N_22946,N_22504,N_22581);
or U22947 (N_22947,N_22559,N_22515);
nor U22948 (N_22948,N_22557,N_22705);
nor U22949 (N_22949,N_22687,N_22573);
and U22950 (N_22950,N_22741,N_22666);
nor U22951 (N_22951,N_22602,N_22738);
xnor U22952 (N_22952,N_22549,N_22601);
and U22953 (N_22953,N_22640,N_22575);
xnor U22954 (N_22954,N_22626,N_22523);
xor U22955 (N_22955,N_22691,N_22740);
and U22956 (N_22956,N_22717,N_22730);
or U22957 (N_22957,N_22670,N_22519);
and U22958 (N_22958,N_22500,N_22577);
nand U22959 (N_22959,N_22726,N_22545);
nor U22960 (N_22960,N_22567,N_22698);
nor U22961 (N_22961,N_22511,N_22738);
or U22962 (N_22962,N_22665,N_22588);
nor U22963 (N_22963,N_22662,N_22570);
nor U22964 (N_22964,N_22670,N_22735);
or U22965 (N_22965,N_22673,N_22580);
nand U22966 (N_22966,N_22620,N_22680);
nor U22967 (N_22967,N_22681,N_22559);
nand U22968 (N_22968,N_22693,N_22710);
nand U22969 (N_22969,N_22516,N_22748);
nand U22970 (N_22970,N_22602,N_22599);
xnor U22971 (N_22971,N_22695,N_22706);
nor U22972 (N_22972,N_22502,N_22538);
nand U22973 (N_22973,N_22578,N_22727);
xnor U22974 (N_22974,N_22662,N_22538);
nor U22975 (N_22975,N_22583,N_22530);
or U22976 (N_22976,N_22609,N_22531);
nor U22977 (N_22977,N_22685,N_22522);
xor U22978 (N_22978,N_22620,N_22657);
or U22979 (N_22979,N_22736,N_22682);
and U22980 (N_22980,N_22618,N_22662);
and U22981 (N_22981,N_22630,N_22580);
nand U22982 (N_22982,N_22597,N_22740);
xnor U22983 (N_22983,N_22583,N_22686);
or U22984 (N_22984,N_22664,N_22668);
and U22985 (N_22985,N_22505,N_22669);
nor U22986 (N_22986,N_22744,N_22621);
nand U22987 (N_22987,N_22721,N_22690);
and U22988 (N_22988,N_22544,N_22658);
nor U22989 (N_22989,N_22709,N_22556);
nand U22990 (N_22990,N_22728,N_22740);
nand U22991 (N_22991,N_22652,N_22621);
nor U22992 (N_22992,N_22674,N_22693);
xnor U22993 (N_22993,N_22578,N_22540);
or U22994 (N_22994,N_22654,N_22576);
or U22995 (N_22995,N_22548,N_22707);
nand U22996 (N_22996,N_22628,N_22558);
nor U22997 (N_22997,N_22662,N_22511);
nor U22998 (N_22998,N_22618,N_22549);
and U22999 (N_22999,N_22707,N_22668);
nor U23000 (N_23000,N_22761,N_22804);
or U23001 (N_23001,N_22955,N_22951);
and U23002 (N_23002,N_22997,N_22885);
nor U23003 (N_23003,N_22888,N_22891);
or U23004 (N_23004,N_22822,N_22904);
and U23005 (N_23005,N_22855,N_22970);
and U23006 (N_23006,N_22949,N_22856);
or U23007 (N_23007,N_22959,N_22988);
nand U23008 (N_23008,N_22847,N_22807);
and U23009 (N_23009,N_22849,N_22875);
nand U23010 (N_23010,N_22957,N_22775);
nand U23011 (N_23011,N_22884,N_22964);
or U23012 (N_23012,N_22985,N_22950);
nand U23013 (N_23013,N_22859,N_22866);
and U23014 (N_23014,N_22924,N_22889);
nand U23015 (N_23015,N_22994,N_22938);
nand U23016 (N_23016,N_22757,N_22786);
or U23017 (N_23017,N_22784,N_22917);
nand U23018 (N_23018,N_22844,N_22800);
and U23019 (N_23019,N_22863,N_22790);
xor U23020 (N_23020,N_22795,N_22810);
and U23021 (N_23021,N_22901,N_22882);
nand U23022 (N_23022,N_22978,N_22987);
nand U23023 (N_23023,N_22782,N_22835);
nor U23024 (N_23024,N_22868,N_22945);
or U23025 (N_23025,N_22909,N_22990);
nor U23026 (N_23026,N_22817,N_22843);
xor U23027 (N_23027,N_22797,N_22829);
xor U23028 (N_23028,N_22864,N_22971);
xnor U23029 (N_23029,N_22911,N_22975);
and U23030 (N_23030,N_22759,N_22780);
xnor U23031 (N_23031,N_22893,N_22941);
and U23032 (N_23032,N_22871,N_22976);
and U23033 (N_23033,N_22887,N_22922);
nor U23034 (N_23034,N_22979,N_22896);
and U23035 (N_23035,N_22862,N_22956);
or U23036 (N_23036,N_22999,N_22842);
and U23037 (N_23037,N_22894,N_22993);
nor U23038 (N_23038,N_22878,N_22837);
or U23039 (N_23039,N_22865,N_22915);
nor U23040 (N_23040,N_22883,N_22787);
and U23041 (N_23041,N_22921,N_22992);
or U23042 (N_23042,N_22753,N_22813);
or U23043 (N_23043,N_22845,N_22792);
xnor U23044 (N_23044,N_22902,N_22953);
or U23045 (N_23045,N_22919,N_22857);
nand U23046 (N_23046,N_22838,N_22903);
xnor U23047 (N_23047,N_22793,N_22954);
xor U23048 (N_23048,N_22989,N_22886);
and U23049 (N_23049,N_22880,N_22890);
nor U23050 (N_23050,N_22934,N_22834);
and U23051 (N_23051,N_22806,N_22939);
and U23052 (N_23052,N_22769,N_22861);
nand U23053 (N_23053,N_22852,N_22832);
xnor U23054 (N_23054,N_22751,N_22984);
and U23055 (N_23055,N_22819,N_22765);
and U23056 (N_23056,N_22928,N_22848);
nand U23057 (N_23057,N_22969,N_22828);
nor U23058 (N_23058,N_22972,N_22826);
or U23059 (N_23059,N_22820,N_22824);
or U23060 (N_23060,N_22998,N_22799);
nand U23061 (N_23061,N_22967,N_22879);
or U23062 (N_23062,N_22965,N_22815);
nand U23063 (N_23063,N_22977,N_22974);
xnor U23064 (N_23064,N_22756,N_22867);
and U23065 (N_23065,N_22899,N_22986);
xnor U23066 (N_23066,N_22791,N_22860);
xor U23067 (N_23067,N_22913,N_22906);
nand U23068 (N_23068,N_22962,N_22777);
xor U23069 (N_23069,N_22774,N_22910);
nor U23070 (N_23070,N_22771,N_22814);
and U23071 (N_23071,N_22764,N_22783);
nor U23072 (N_23072,N_22948,N_22762);
and U23073 (N_23073,N_22839,N_22981);
nor U23074 (N_23074,N_22973,N_22770);
or U23075 (N_23075,N_22933,N_22869);
or U23076 (N_23076,N_22767,N_22961);
nor U23077 (N_23077,N_22755,N_22779);
and U23078 (N_23078,N_22932,N_22912);
nand U23079 (N_23079,N_22943,N_22827);
nand U23080 (N_23080,N_22929,N_22947);
nor U23081 (N_23081,N_22872,N_22805);
and U23082 (N_23082,N_22966,N_22831);
or U23083 (N_23083,N_22881,N_22931);
nor U23084 (N_23084,N_22823,N_22853);
nor U23085 (N_23085,N_22960,N_22768);
or U23086 (N_23086,N_22916,N_22942);
or U23087 (N_23087,N_22801,N_22796);
nand U23088 (N_23088,N_22940,N_22968);
nand U23089 (N_23089,N_22809,N_22907);
and U23090 (N_23090,N_22811,N_22920);
xor U23091 (N_23091,N_22846,N_22982);
nand U23092 (N_23092,N_22788,N_22850);
nor U23093 (N_23093,N_22803,N_22925);
xor U23094 (N_23094,N_22825,N_22773);
and U23095 (N_23095,N_22918,N_22754);
and U23096 (N_23096,N_22851,N_22840);
nand U23097 (N_23097,N_22766,N_22996);
xor U23098 (N_23098,N_22946,N_22892);
xnor U23099 (N_23099,N_22854,N_22776);
nor U23100 (N_23100,N_22798,N_22991);
and U23101 (N_23101,N_22812,N_22836);
nor U23102 (N_23102,N_22874,N_22895);
xnor U23103 (N_23103,N_22833,N_22778);
xor U23104 (N_23104,N_22952,N_22936);
and U23105 (N_23105,N_22980,N_22926);
xor U23106 (N_23106,N_22935,N_22794);
and U23107 (N_23107,N_22752,N_22914);
and U23108 (N_23108,N_22930,N_22858);
xnor U23109 (N_23109,N_22873,N_22905);
xnor U23110 (N_23110,N_22995,N_22763);
and U23111 (N_23111,N_22958,N_22816);
or U23112 (N_23112,N_22808,N_22785);
xnor U23113 (N_23113,N_22781,N_22821);
or U23114 (N_23114,N_22897,N_22760);
or U23115 (N_23115,N_22963,N_22789);
xnor U23116 (N_23116,N_22877,N_22876);
and U23117 (N_23117,N_22908,N_22983);
nand U23118 (N_23118,N_22818,N_22898);
or U23119 (N_23119,N_22944,N_22841);
nor U23120 (N_23120,N_22927,N_22802);
nand U23121 (N_23121,N_22937,N_22870);
xnor U23122 (N_23122,N_22758,N_22900);
nand U23123 (N_23123,N_22750,N_22830);
xor U23124 (N_23124,N_22772,N_22923);
nor U23125 (N_23125,N_22886,N_22918);
nand U23126 (N_23126,N_22947,N_22844);
nor U23127 (N_23127,N_22914,N_22971);
or U23128 (N_23128,N_22875,N_22900);
nand U23129 (N_23129,N_22786,N_22874);
nor U23130 (N_23130,N_22978,N_22808);
and U23131 (N_23131,N_22959,N_22768);
and U23132 (N_23132,N_22815,N_22910);
nor U23133 (N_23133,N_22919,N_22921);
or U23134 (N_23134,N_22879,N_22841);
nor U23135 (N_23135,N_22947,N_22794);
and U23136 (N_23136,N_22907,N_22833);
or U23137 (N_23137,N_22918,N_22854);
and U23138 (N_23138,N_22932,N_22969);
nand U23139 (N_23139,N_22938,N_22983);
nand U23140 (N_23140,N_22955,N_22911);
xnor U23141 (N_23141,N_22906,N_22847);
nand U23142 (N_23142,N_22908,N_22837);
nor U23143 (N_23143,N_22904,N_22763);
nand U23144 (N_23144,N_22852,N_22900);
xor U23145 (N_23145,N_22776,N_22843);
and U23146 (N_23146,N_22827,N_22833);
nand U23147 (N_23147,N_22794,N_22969);
or U23148 (N_23148,N_22954,N_22852);
nor U23149 (N_23149,N_22903,N_22978);
nor U23150 (N_23150,N_22800,N_22787);
and U23151 (N_23151,N_22846,N_22772);
nand U23152 (N_23152,N_22990,N_22839);
nor U23153 (N_23153,N_22939,N_22876);
nand U23154 (N_23154,N_22958,N_22924);
and U23155 (N_23155,N_22789,N_22865);
nor U23156 (N_23156,N_22968,N_22900);
nand U23157 (N_23157,N_22917,N_22938);
and U23158 (N_23158,N_22857,N_22785);
nand U23159 (N_23159,N_22883,N_22785);
or U23160 (N_23160,N_22778,N_22886);
nor U23161 (N_23161,N_22955,N_22797);
nand U23162 (N_23162,N_22975,N_22944);
nand U23163 (N_23163,N_22960,N_22890);
or U23164 (N_23164,N_22829,N_22961);
or U23165 (N_23165,N_22882,N_22752);
or U23166 (N_23166,N_22951,N_22753);
xnor U23167 (N_23167,N_22973,N_22939);
nand U23168 (N_23168,N_22787,N_22831);
nor U23169 (N_23169,N_22807,N_22964);
nand U23170 (N_23170,N_22875,N_22863);
nand U23171 (N_23171,N_22868,N_22947);
or U23172 (N_23172,N_22797,N_22815);
or U23173 (N_23173,N_22803,N_22909);
and U23174 (N_23174,N_22806,N_22998);
nor U23175 (N_23175,N_22822,N_22815);
xor U23176 (N_23176,N_22984,N_22752);
nor U23177 (N_23177,N_22860,N_22933);
xor U23178 (N_23178,N_22770,N_22935);
nand U23179 (N_23179,N_22934,N_22878);
or U23180 (N_23180,N_22857,N_22776);
xnor U23181 (N_23181,N_22856,N_22929);
or U23182 (N_23182,N_22757,N_22905);
nand U23183 (N_23183,N_22785,N_22753);
nand U23184 (N_23184,N_22895,N_22919);
nor U23185 (N_23185,N_22751,N_22910);
xor U23186 (N_23186,N_22908,N_22874);
nor U23187 (N_23187,N_22806,N_22841);
xnor U23188 (N_23188,N_22804,N_22960);
and U23189 (N_23189,N_22875,N_22785);
nand U23190 (N_23190,N_22909,N_22765);
nor U23191 (N_23191,N_22796,N_22794);
nor U23192 (N_23192,N_22927,N_22934);
xor U23193 (N_23193,N_22926,N_22782);
nand U23194 (N_23194,N_22856,N_22920);
nand U23195 (N_23195,N_22837,N_22758);
nor U23196 (N_23196,N_22796,N_22824);
and U23197 (N_23197,N_22862,N_22889);
nand U23198 (N_23198,N_22916,N_22770);
nand U23199 (N_23199,N_22996,N_22773);
xor U23200 (N_23200,N_22780,N_22853);
or U23201 (N_23201,N_22969,N_22943);
nor U23202 (N_23202,N_22933,N_22956);
nand U23203 (N_23203,N_22848,N_22791);
or U23204 (N_23204,N_22964,N_22887);
xnor U23205 (N_23205,N_22828,N_22813);
or U23206 (N_23206,N_22987,N_22916);
nor U23207 (N_23207,N_22846,N_22992);
or U23208 (N_23208,N_22973,N_22951);
nor U23209 (N_23209,N_22877,N_22928);
xor U23210 (N_23210,N_22954,N_22763);
xnor U23211 (N_23211,N_22811,N_22977);
and U23212 (N_23212,N_22790,N_22934);
and U23213 (N_23213,N_22915,N_22780);
nor U23214 (N_23214,N_22915,N_22973);
nand U23215 (N_23215,N_22939,N_22945);
nand U23216 (N_23216,N_22829,N_22777);
nand U23217 (N_23217,N_22775,N_22780);
nand U23218 (N_23218,N_22767,N_22948);
or U23219 (N_23219,N_22885,N_22825);
and U23220 (N_23220,N_22802,N_22909);
xnor U23221 (N_23221,N_22776,N_22831);
nand U23222 (N_23222,N_22939,N_22855);
nand U23223 (N_23223,N_22867,N_22900);
nor U23224 (N_23224,N_22859,N_22804);
and U23225 (N_23225,N_22998,N_22917);
and U23226 (N_23226,N_22827,N_22881);
and U23227 (N_23227,N_22862,N_22818);
xnor U23228 (N_23228,N_22985,N_22781);
and U23229 (N_23229,N_22973,N_22803);
and U23230 (N_23230,N_22991,N_22879);
and U23231 (N_23231,N_22825,N_22928);
xor U23232 (N_23232,N_22828,N_22946);
xnor U23233 (N_23233,N_22995,N_22909);
and U23234 (N_23234,N_22994,N_22765);
or U23235 (N_23235,N_22848,N_22897);
nor U23236 (N_23236,N_22947,N_22956);
nand U23237 (N_23237,N_22913,N_22821);
nand U23238 (N_23238,N_22911,N_22948);
xnor U23239 (N_23239,N_22939,N_22923);
xnor U23240 (N_23240,N_22988,N_22752);
and U23241 (N_23241,N_22808,N_22898);
nand U23242 (N_23242,N_22906,N_22911);
nand U23243 (N_23243,N_22755,N_22979);
nand U23244 (N_23244,N_22959,N_22933);
and U23245 (N_23245,N_22963,N_22759);
nor U23246 (N_23246,N_22960,N_22879);
nand U23247 (N_23247,N_22836,N_22987);
or U23248 (N_23248,N_22892,N_22939);
or U23249 (N_23249,N_22842,N_22817);
xnor U23250 (N_23250,N_23213,N_23054);
or U23251 (N_23251,N_23006,N_23036);
nand U23252 (N_23252,N_23155,N_23074);
nor U23253 (N_23253,N_23218,N_23138);
nand U23254 (N_23254,N_23078,N_23148);
nor U23255 (N_23255,N_23048,N_23002);
and U23256 (N_23256,N_23115,N_23146);
xnor U23257 (N_23257,N_23189,N_23034);
and U23258 (N_23258,N_23145,N_23119);
nor U23259 (N_23259,N_23045,N_23226);
and U23260 (N_23260,N_23086,N_23195);
xor U23261 (N_23261,N_23039,N_23116);
or U23262 (N_23262,N_23181,N_23170);
and U23263 (N_23263,N_23124,N_23245);
and U23264 (N_23264,N_23171,N_23016);
or U23265 (N_23265,N_23239,N_23033);
nand U23266 (N_23266,N_23214,N_23201);
nand U23267 (N_23267,N_23069,N_23126);
xnor U23268 (N_23268,N_23202,N_23219);
nand U23269 (N_23269,N_23096,N_23169);
and U23270 (N_23270,N_23117,N_23234);
xor U23271 (N_23271,N_23089,N_23157);
and U23272 (N_23272,N_23075,N_23029);
nand U23273 (N_23273,N_23024,N_23136);
and U23274 (N_23274,N_23184,N_23191);
nor U23275 (N_23275,N_23000,N_23076);
nor U23276 (N_23276,N_23166,N_23244);
xor U23277 (N_23277,N_23068,N_23200);
xnor U23278 (N_23278,N_23102,N_23211);
nor U23279 (N_23279,N_23176,N_23122);
nand U23280 (N_23280,N_23204,N_23070);
nand U23281 (N_23281,N_23158,N_23090);
or U23282 (N_23282,N_23099,N_23123);
nand U23283 (N_23283,N_23107,N_23229);
xor U23284 (N_23284,N_23153,N_23167);
or U23285 (N_23285,N_23030,N_23240);
nor U23286 (N_23286,N_23110,N_23025);
nor U23287 (N_23287,N_23179,N_23005);
nor U23288 (N_23288,N_23134,N_23080);
nor U23289 (N_23289,N_23083,N_23185);
or U23290 (N_23290,N_23132,N_23040);
nand U23291 (N_23291,N_23142,N_23101);
or U23292 (N_23292,N_23130,N_23233);
nand U23293 (N_23293,N_23174,N_23066);
and U23294 (N_23294,N_23223,N_23209);
nand U23295 (N_23295,N_23178,N_23015);
nand U23296 (N_23296,N_23088,N_23023);
nor U23297 (N_23297,N_23231,N_23183);
and U23298 (N_23298,N_23073,N_23051);
and U23299 (N_23299,N_23063,N_23053);
nor U23300 (N_23300,N_23220,N_23222);
xnor U23301 (N_23301,N_23084,N_23060);
nand U23302 (N_23302,N_23061,N_23206);
or U23303 (N_23303,N_23182,N_23205);
and U23304 (N_23304,N_23129,N_23236);
or U23305 (N_23305,N_23164,N_23019);
nor U23306 (N_23306,N_23192,N_23010);
and U23307 (N_23307,N_23003,N_23237);
nand U23308 (N_23308,N_23215,N_23028);
xor U23309 (N_23309,N_23022,N_23199);
and U23310 (N_23310,N_23121,N_23049);
or U23311 (N_23311,N_23103,N_23143);
or U23312 (N_23312,N_23091,N_23046);
and U23313 (N_23313,N_23248,N_23020);
nand U23314 (N_23314,N_23112,N_23026);
xor U23315 (N_23315,N_23198,N_23092);
xnor U23316 (N_23316,N_23127,N_23125);
or U23317 (N_23317,N_23071,N_23186);
and U23318 (N_23318,N_23044,N_23150);
nand U23319 (N_23319,N_23141,N_23007);
nand U23320 (N_23320,N_23197,N_23095);
and U23321 (N_23321,N_23012,N_23173);
and U23322 (N_23322,N_23057,N_23052);
xor U23323 (N_23323,N_23149,N_23047);
nand U23324 (N_23324,N_23072,N_23235);
xnor U23325 (N_23325,N_23108,N_23188);
or U23326 (N_23326,N_23177,N_23227);
and U23327 (N_23327,N_23131,N_23113);
nand U23328 (N_23328,N_23135,N_23104);
nand U23329 (N_23329,N_23175,N_23059);
nor U23330 (N_23330,N_23203,N_23137);
and U23331 (N_23331,N_23147,N_23154);
nand U23332 (N_23332,N_23207,N_23249);
and U23333 (N_23333,N_23050,N_23043);
or U23334 (N_23334,N_23065,N_23001);
xor U23335 (N_23335,N_23011,N_23105);
xor U23336 (N_23336,N_23027,N_23087);
nor U23337 (N_23337,N_23225,N_23111);
and U23338 (N_23338,N_23081,N_23221);
nand U23339 (N_23339,N_23187,N_23161);
nand U23340 (N_23340,N_23159,N_23120);
xnor U23341 (N_23341,N_23210,N_23064);
nand U23342 (N_23342,N_23114,N_23038);
xor U23343 (N_23343,N_23241,N_23180);
nor U23344 (N_23344,N_23021,N_23042);
nor U23345 (N_23345,N_23017,N_23208);
and U23346 (N_23346,N_23031,N_23098);
and U23347 (N_23347,N_23242,N_23032);
and U23348 (N_23348,N_23041,N_23156);
nand U23349 (N_23349,N_23014,N_23212);
and U23350 (N_23350,N_23172,N_23009);
and U23351 (N_23351,N_23160,N_23168);
or U23352 (N_23352,N_23085,N_23194);
nor U23353 (N_23353,N_23056,N_23139);
nor U23354 (N_23354,N_23193,N_23109);
xor U23355 (N_23355,N_23037,N_23232);
or U23356 (N_23356,N_23162,N_23118);
nor U23357 (N_23357,N_23062,N_23055);
or U23358 (N_23358,N_23246,N_23018);
nor U23359 (N_23359,N_23077,N_23152);
nor U23360 (N_23360,N_23100,N_23140);
and U23361 (N_23361,N_23196,N_23165);
and U23362 (N_23362,N_23097,N_23228);
xor U23363 (N_23363,N_23238,N_23008);
xor U23364 (N_23364,N_23106,N_23133);
and U23365 (N_23365,N_23013,N_23224);
or U23366 (N_23366,N_23093,N_23004);
and U23367 (N_23367,N_23247,N_23151);
nor U23368 (N_23368,N_23094,N_23216);
nand U23369 (N_23369,N_23144,N_23230);
and U23370 (N_23370,N_23190,N_23163);
and U23371 (N_23371,N_23243,N_23079);
and U23372 (N_23372,N_23067,N_23058);
or U23373 (N_23373,N_23217,N_23128);
nand U23374 (N_23374,N_23035,N_23082);
nand U23375 (N_23375,N_23058,N_23130);
xnor U23376 (N_23376,N_23220,N_23219);
nand U23377 (N_23377,N_23071,N_23156);
and U23378 (N_23378,N_23068,N_23172);
nor U23379 (N_23379,N_23173,N_23081);
nor U23380 (N_23380,N_23160,N_23025);
or U23381 (N_23381,N_23128,N_23127);
xnor U23382 (N_23382,N_23164,N_23101);
and U23383 (N_23383,N_23098,N_23221);
nand U23384 (N_23384,N_23205,N_23024);
and U23385 (N_23385,N_23130,N_23240);
and U23386 (N_23386,N_23110,N_23241);
and U23387 (N_23387,N_23059,N_23082);
nand U23388 (N_23388,N_23160,N_23111);
or U23389 (N_23389,N_23205,N_23146);
or U23390 (N_23390,N_23019,N_23157);
xor U23391 (N_23391,N_23163,N_23139);
or U23392 (N_23392,N_23069,N_23186);
xor U23393 (N_23393,N_23001,N_23045);
or U23394 (N_23394,N_23196,N_23097);
and U23395 (N_23395,N_23199,N_23008);
and U23396 (N_23396,N_23181,N_23202);
xnor U23397 (N_23397,N_23196,N_23016);
nand U23398 (N_23398,N_23112,N_23051);
and U23399 (N_23399,N_23015,N_23154);
xor U23400 (N_23400,N_23193,N_23021);
nor U23401 (N_23401,N_23006,N_23102);
and U23402 (N_23402,N_23128,N_23184);
or U23403 (N_23403,N_23208,N_23118);
or U23404 (N_23404,N_23157,N_23204);
xnor U23405 (N_23405,N_23123,N_23040);
xnor U23406 (N_23406,N_23191,N_23185);
or U23407 (N_23407,N_23059,N_23137);
xor U23408 (N_23408,N_23007,N_23200);
xnor U23409 (N_23409,N_23156,N_23077);
nor U23410 (N_23410,N_23225,N_23050);
xor U23411 (N_23411,N_23048,N_23127);
and U23412 (N_23412,N_23099,N_23104);
or U23413 (N_23413,N_23247,N_23020);
nand U23414 (N_23414,N_23054,N_23134);
and U23415 (N_23415,N_23128,N_23167);
or U23416 (N_23416,N_23082,N_23211);
and U23417 (N_23417,N_23166,N_23107);
and U23418 (N_23418,N_23114,N_23131);
nand U23419 (N_23419,N_23185,N_23212);
nand U23420 (N_23420,N_23188,N_23054);
nor U23421 (N_23421,N_23136,N_23106);
nor U23422 (N_23422,N_23050,N_23241);
nor U23423 (N_23423,N_23058,N_23170);
nand U23424 (N_23424,N_23173,N_23035);
nor U23425 (N_23425,N_23076,N_23037);
or U23426 (N_23426,N_23160,N_23040);
xnor U23427 (N_23427,N_23188,N_23123);
nor U23428 (N_23428,N_23247,N_23106);
or U23429 (N_23429,N_23194,N_23149);
or U23430 (N_23430,N_23117,N_23096);
and U23431 (N_23431,N_23003,N_23245);
xor U23432 (N_23432,N_23034,N_23188);
nand U23433 (N_23433,N_23122,N_23062);
nor U23434 (N_23434,N_23046,N_23014);
xor U23435 (N_23435,N_23249,N_23216);
or U23436 (N_23436,N_23001,N_23174);
nand U23437 (N_23437,N_23139,N_23010);
xnor U23438 (N_23438,N_23212,N_23092);
and U23439 (N_23439,N_23030,N_23006);
xnor U23440 (N_23440,N_23179,N_23206);
xor U23441 (N_23441,N_23099,N_23188);
nor U23442 (N_23442,N_23105,N_23052);
and U23443 (N_23443,N_23084,N_23041);
nand U23444 (N_23444,N_23209,N_23244);
nand U23445 (N_23445,N_23110,N_23090);
nor U23446 (N_23446,N_23089,N_23079);
xor U23447 (N_23447,N_23147,N_23019);
and U23448 (N_23448,N_23145,N_23109);
nor U23449 (N_23449,N_23243,N_23001);
xnor U23450 (N_23450,N_23087,N_23105);
and U23451 (N_23451,N_23006,N_23225);
and U23452 (N_23452,N_23098,N_23047);
nor U23453 (N_23453,N_23178,N_23190);
or U23454 (N_23454,N_23008,N_23101);
nor U23455 (N_23455,N_23184,N_23032);
and U23456 (N_23456,N_23229,N_23150);
xor U23457 (N_23457,N_23185,N_23094);
nand U23458 (N_23458,N_23204,N_23232);
xnor U23459 (N_23459,N_23157,N_23238);
xnor U23460 (N_23460,N_23121,N_23144);
or U23461 (N_23461,N_23163,N_23052);
nor U23462 (N_23462,N_23161,N_23072);
nand U23463 (N_23463,N_23019,N_23025);
nor U23464 (N_23464,N_23095,N_23235);
nand U23465 (N_23465,N_23215,N_23112);
or U23466 (N_23466,N_23048,N_23067);
and U23467 (N_23467,N_23131,N_23175);
nand U23468 (N_23468,N_23236,N_23024);
or U23469 (N_23469,N_23175,N_23219);
nand U23470 (N_23470,N_23107,N_23159);
or U23471 (N_23471,N_23096,N_23140);
xor U23472 (N_23472,N_23034,N_23136);
nor U23473 (N_23473,N_23176,N_23085);
or U23474 (N_23474,N_23170,N_23213);
or U23475 (N_23475,N_23248,N_23140);
xor U23476 (N_23476,N_23083,N_23054);
xor U23477 (N_23477,N_23098,N_23025);
xnor U23478 (N_23478,N_23022,N_23086);
or U23479 (N_23479,N_23161,N_23092);
or U23480 (N_23480,N_23222,N_23076);
or U23481 (N_23481,N_23068,N_23192);
xor U23482 (N_23482,N_23032,N_23112);
or U23483 (N_23483,N_23151,N_23081);
xor U23484 (N_23484,N_23169,N_23094);
xnor U23485 (N_23485,N_23126,N_23197);
and U23486 (N_23486,N_23026,N_23076);
and U23487 (N_23487,N_23173,N_23144);
xnor U23488 (N_23488,N_23089,N_23156);
or U23489 (N_23489,N_23193,N_23087);
xnor U23490 (N_23490,N_23205,N_23143);
or U23491 (N_23491,N_23202,N_23012);
and U23492 (N_23492,N_23206,N_23078);
nand U23493 (N_23493,N_23103,N_23156);
or U23494 (N_23494,N_23076,N_23019);
nor U23495 (N_23495,N_23228,N_23237);
and U23496 (N_23496,N_23051,N_23069);
nor U23497 (N_23497,N_23225,N_23237);
nand U23498 (N_23498,N_23041,N_23164);
nand U23499 (N_23499,N_23136,N_23008);
and U23500 (N_23500,N_23278,N_23439);
and U23501 (N_23501,N_23335,N_23444);
and U23502 (N_23502,N_23391,N_23294);
nor U23503 (N_23503,N_23306,N_23314);
and U23504 (N_23504,N_23480,N_23349);
and U23505 (N_23505,N_23256,N_23326);
or U23506 (N_23506,N_23279,N_23342);
nor U23507 (N_23507,N_23420,N_23348);
xnor U23508 (N_23508,N_23400,N_23453);
or U23509 (N_23509,N_23458,N_23380);
xor U23510 (N_23510,N_23300,N_23396);
xor U23511 (N_23511,N_23383,N_23435);
and U23512 (N_23512,N_23336,N_23486);
nand U23513 (N_23513,N_23432,N_23448);
xor U23514 (N_23514,N_23265,N_23473);
nor U23515 (N_23515,N_23327,N_23301);
nand U23516 (N_23516,N_23333,N_23264);
xnor U23517 (N_23517,N_23476,N_23364);
nand U23518 (N_23518,N_23489,N_23491);
nor U23519 (N_23519,N_23367,N_23496);
and U23520 (N_23520,N_23467,N_23465);
and U23521 (N_23521,N_23460,N_23251);
nand U23522 (N_23522,N_23276,N_23266);
or U23523 (N_23523,N_23449,N_23477);
xor U23524 (N_23524,N_23413,N_23255);
or U23525 (N_23525,N_23484,N_23464);
nor U23526 (N_23526,N_23317,N_23463);
nor U23527 (N_23527,N_23299,N_23378);
nor U23528 (N_23528,N_23381,N_23341);
and U23529 (N_23529,N_23321,N_23398);
and U23530 (N_23530,N_23472,N_23382);
nor U23531 (N_23531,N_23292,N_23431);
and U23532 (N_23532,N_23332,N_23457);
nor U23533 (N_23533,N_23297,N_23483);
and U23534 (N_23534,N_23268,N_23282);
nand U23535 (N_23535,N_23310,N_23356);
or U23536 (N_23536,N_23273,N_23423);
xor U23537 (N_23537,N_23395,N_23416);
nor U23538 (N_23538,N_23343,N_23359);
xor U23539 (N_23539,N_23459,N_23320);
nand U23540 (N_23540,N_23375,N_23281);
nor U23541 (N_23541,N_23291,N_23355);
or U23542 (N_23542,N_23417,N_23414);
and U23543 (N_23543,N_23482,N_23269);
nand U23544 (N_23544,N_23402,N_23346);
xor U23545 (N_23545,N_23328,N_23452);
and U23546 (N_23546,N_23475,N_23271);
xnor U23547 (N_23547,N_23471,N_23370);
xor U23548 (N_23548,N_23428,N_23286);
xnor U23549 (N_23549,N_23311,N_23366);
nand U23550 (N_23550,N_23258,N_23451);
or U23551 (N_23551,N_23426,N_23401);
xnor U23552 (N_23552,N_23325,N_23322);
nand U23553 (N_23553,N_23334,N_23371);
or U23554 (N_23554,N_23280,N_23481);
nand U23555 (N_23555,N_23390,N_23302);
nor U23556 (N_23556,N_23408,N_23354);
nor U23557 (N_23557,N_23450,N_23261);
nand U23558 (N_23558,N_23365,N_23495);
xnor U23559 (N_23559,N_23309,N_23454);
xor U23560 (N_23560,N_23340,N_23368);
or U23561 (N_23561,N_23376,N_23296);
nand U23562 (N_23562,N_23393,N_23468);
or U23563 (N_23563,N_23339,N_23338);
nor U23564 (N_23564,N_23316,N_23474);
and U23565 (N_23565,N_23419,N_23331);
nor U23566 (N_23566,N_23399,N_23403);
and U23567 (N_23567,N_23352,N_23360);
nand U23568 (N_23568,N_23350,N_23290);
nand U23569 (N_23569,N_23440,N_23461);
xnor U23570 (N_23570,N_23319,N_23295);
nand U23571 (N_23571,N_23386,N_23397);
xor U23572 (N_23572,N_23389,N_23384);
nand U23573 (N_23573,N_23410,N_23443);
or U23574 (N_23574,N_23425,N_23323);
nor U23575 (N_23575,N_23363,N_23353);
nand U23576 (N_23576,N_23490,N_23254);
nor U23577 (N_23577,N_23379,N_23313);
and U23578 (N_23578,N_23492,N_23385);
and U23579 (N_23579,N_23424,N_23388);
nand U23580 (N_23580,N_23307,N_23422);
nand U23581 (N_23581,N_23498,N_23442);
or U23582 (N_23582,N_23446,N_23369);
nor U23583 (N_23583,N_23330,N_23287);
nand U23584 (N_23584,N_23257,N_23466);
or U23585 (N_23585,N_23304,N_23298);
xnor U23586 (N_23586,N_23437,N_23411);
or U23587 (N_23587,N_23318,N_23479);
nor U23588 (N_23588,N_23358,N_23303);
and U23589 (N_23589,N_23315,N_23387);
and U23590 (N_23590,N_23493,N_23262);
and U23591 (N_23591,N_23324,N_23374);
or U23592 (N_23592,N_23404,N_23427);
xnor U23593 (N_23593,N_23329,N_23361);
or U23594 (N_23594,N_23259,N_23434);
xnor U23595 (N_23595,N_23308,N_23293);
nor U23596 (N_23596,N_23429,N_23283);
or U23597 (N_23597,N_23288,N_23272);
xor U23598 (N_23598,N_23285,N_23469);
or U23599 (N_23599,N_23415,N_23267);
nand U23600 (N_23600,N_23478,N_23270);
and U23601 (N_23601,N_23305,N_23277);
nor U23602 (N_23602,N_23289,N_23487);
or U23603 (N_23603,N_23497,N_23284);
xor U23604 (N_23604,N_23394,N_23436);
and U23605 (N_23605,N_23412,N_23392);
nand U23606 (N_23606,N_23456,N_23337);
and U23607 (N_23607,N_23351,N_23362);
xnor U23608 (N_23608,N_23263,N_23445);
and U23609 (N_23609,N_23433,N_23409);
and U23610 (N_23610,N_23462,N_23455);
and U23611 (N_23611,N_23250,N_23260);
or U23612 (N_23612,N_23312,N_23344);
nand U23613 (N_23613,N_23438,N_23441);
and U23614 (N_23614,N_23418,N_23275);
and U23615 (N_23615,N_23407,N_23252);
xnor U23616 (N_23616,N_23447,N_23357);
or U23617 (N_23617,N_23405,N_23253);
xnor U23618 (N_23618,N_23274,N_23347);
xnor U23619 (N_23619,N_23406,N_23345);
nand U23620 (N_23620,N_23485,N_23372);
nand U23621 (N_23621,N_23499,N_23488);
xnor U23622 (N_23622,N_23494,N_23430);
nor U23623 (N_23623,N_23377,N_23421);
or U23624 (N_23624,N_23373,N_23470);
nand U23625 (N_23625,N_23411,N_23480);
xor U23626 (N_23626,N_23448,N_23293);
nand U23627 (N_23627,N_23478,N_23312);
nor U23628 (N_23628,N_23315,N_23277);
xnor U23629 (N_23629,N_23491,N_23429);
xnor U23630 (N_23630,N_23266,N_23288);
xor U23631 (N_23631,N_23415,N_23257);
nand U23632 (N_23632,N_23489,N_23322);
nand U23633 (N_23633,N_23362,N_23263);
nand U23634 (N_23634,N_23487,N_23305);
and U23635 (N_23635,N_23427,N_23297);
and U23636 (N_23636,N_23407,N_23402);
or U23637 (N_23637,N_23450,N_23404);
nand U23638 (N_23638,N_23489,N_23393);
or U23639 (N_23639,N_23284,N_23385);
nor U23640 (N_23640,N_23293,N_23315);
nand U23641 (N_23641,N_23373,N_23251);
nor U23642 (N_23642,N_23353,N_23362);
or U23643 (N_23643,N_23283,N_23498);
nand U23644 (N_23644,N_23373,N_23288);
or U23645 (N_23645,N_23456,N_23259);
nand U23646 (N_23646,N_23403,N_23370);
or U23647 (N_23647,N_23442,N_23326);
and U23648 (N_23648,N_23379,N_23329);
nand U23649 (N_23649,N_23298,N_23439);
nand U23650 (N_23650,N_23435,N_23468);
and U23651 (N_23651,N_23285,N_23327);
nor U23652 (N_23652,N_23295,N_23322);
nand U23653 (N_23653,N_23351,N_23419);
xnor U23654 (N_23654,N_23363,N_23425);
and U23655 (N_23655,N_23338,N_23297);
and U23656 (N_23656,N_23270,N_23348);
or U23657 (N_23657,N_23272,N_23257);
or U23658 (N_23658,N_23396,N_23475);
xor U23659 (N_23659,N_23315,N_23337);
xnor U23660 (N_23660,N_23313,N_23475);
nor U23661 (N_23661,N_23257,N_23273);
or U23662 (N_23662,N_23317,N_23268);
nor U23663 (N_23663,N_23250,N_23293);
nand U23664 (N_23664,N_23329,N_23397);
and U23665 (N_23665,N_23422,N_23372);
or U23666 (N_23666,N_23338,N_23315);
xor U23667 (N_23667,N_23431,N_23324);
or U23668 (N_23668,N_23302,N_23277);
xnor U23669 (N_23669,N_23444,N_23403);
nor U23670 (N_23670,N_23402,N_23416);
xnor U23671 (N_23671,N_23320,N_23367);
xor U23672 (N_23672,N_23322,N_23302);
nor U23673 (N_23673,N_23397,N_23361);
xor U23674 (N_23674,N_23473,N_23387);
xor U23675 (N_23675,N_23293,N_23345);
or U23676 (N_23676,N_23491,N_23457);
and U23677 (N_23677,N_23355,N_23430);
and U23678 (N_23678,N_23291,N_23338);
nor U23679 (N_23679,N_23341,N_23411);
nand U23680 (N_23680,N_23493,N_23255);
xnor U23681 (N_23681,N_23343,N_23386);
and U23682 (N_23682,N_23439,N_23319);
xnor U23683 (N_23683,N_23395,N_23422);
and U23684 (N_23684,N_23346,N_23473);
nor U23685 (N_23685,N_23342,N_23327);
nor U23686 (N_23686,N_23342,N_23353);
nand U23687 (N_23687,N_23345,N_23403);
xnor U23688 (N_23688,N_23449,N_23445);
and U23689 (N_23689,N_23338,N_23422);
and U23690 (N_23690,N_23325,N_23482);
or U23691 (N_23691,N_23455,N_23435);
xnor U23692 (N_23692,N_23343,N_23342);
and U23693 (N_23693,N_23252,N_23300);
nand U23694 (N_23694,N_23453,N_23469);
xor U23695 (N_23695,N_23496,N_23262);
nor U23696 (N_23696,N_23297,N_23270);
nor U23697 (N_23697,N_23285,N_23351);
or U23698 (N_23698,N_23489,N_23319);
and U23699 (N_23699,N_23392,N_23337);
nor U23700 (N_23700,N_23344,N_23360);
xor U23701 (N_23701,N_23389,N_23256);
or U23702 (N_23702,N_23430,N_23454);
nor U23703 (N_23703,N_23269,N_23451);
and U23704 (N_23704,N_23252,N_23493);
xor U23705 (N_23705,N_23488,N_23287);
nand U23706 (N_23706,N_23383,N_23388);
and U23707 (N_23707,N_23304,N_23406);
nor U23708 (N_23708,N_23367,N_23255);
xnor U23709 (N_23709,N_23496,N_23470);
or U23710 (N_23710,N_23432,N_23394);
xnor U23711 (N_23711,N_23368,N_23356);
nand U23712 (N_23712,N_23494,N_23383);
and U23713 (N_23713,N_23251,N_23454);
xnor U23714 (N_23714,N_23479,N_23483);
nor U23715 (N_23715,N_23288,N_23305);
and U23716 (N_23716,N_23455,N_23307);
xor U23717 (N_23717,N_23341,N_23283);
nor U23718 (N_23718,N_23386,N_23412);
or U23719 (N_23719,N_23283,N_23270);
nand U23720 (N_23720,N_23397,N_23433);
or U23721 (N_23721,N_23343,N_23363);
xor U23722 (N_23722,N_23328,N_23438);
nand U23723 (N_23723,N_23287,N_23254);
xor U23724 (N_23724,N_23271,N_23477);
nand U23725 (N_23725,N_23482,N_23491);
nor U23726 (N_23726,N_23494,N_23309);
nor U23727 (N_23727,N_23268,N_23406);
nor U23728 (N_23728,N_23469,N_23350);
nor U23729 (N_23729,N_23398,N_23311);
xnor U23730 (N_23730,N_23418,N_23255);
xnor U23731 (N_23731,N_23279,N_23399);
nand U23732 (N_23732,N_23293,N_23400);
nand U23733 (N_23733,N_23484,N_23300);
nand U23734 (N_23734,N_23457,N_23378);
nand U23735 (N_23735,N_23494,N_23344);
nand U23736 (N_23736,N_23354,N_23466);
and U23737 (N_23737,N_23380,N_23256);
nand U23738 (N_23738,N_23303,N_23373);
nor U23739 (N_23739,N_23447,N_23278);
and U23740 (N_23740,N_23350,N_23445);
nand U23741 (N_23741,N_23321,N_23265);
nor U23742 (N_23742,N_23327,N_23347);
nor U23743 (N_23743,N_23381,N_23327);
nand U23744 (N_23744,N_23276,N_23488);
and U23745 (N_23745,N_23420,N_23330);
or U23746 (N_23746,N_23359,N_23465);
and U23747 (N_23747,N_23260,N_23355);
and U23748 (N_23748,N_23348,N_23471);
xnor U23749 (N_23749,N_23261,N_23437);
or U23750 (N_23750,N_23545,N_23560);
nand U23751 (N_23751,N_23578,N_23732);
or U23752 (N_23752,N_23726,N_23556);
nor U23753 (N_23753,N_23729,N_23553);
or U23754 (N_23754,N_23738,N_23586);
nor U23755 (N_23755,N_23503,N_23609);
nand U23756 (N_23756,N_23510,N_23639);
nand U23757 (N_23757,N_23698,N_23680);
or U23758 (N_23758,N_23615,N_23572);
or U23759 (N_23759,N_23633,N_23636);
or U23760 (N_23760,N_23708,N_23713);
xnor U23761 (N_23761,N_23654,N_23623);
nand U23762 (N_23762,N_23538,N_23569);
nand U23763 (N_23763,N_23735,N_23705);
and U23764 (N_23764,N_23638,N_23563);
and U23765 (N_23765,N_23692,N_23576);
xnor U23766 (N_23766,N_23683,N_23663);
and U23767 (N_23767,N_23512,N_23618);
nand U23768 (N_23768,N_23678,N_23703);
nand U23769 (N_23769,N_23540,N_23524);
nand U23770 (N_23770,N_23621,N_23519);
or U23771 (N_23771,N_23627,N_23635);
nand U23772 (N_23772,N_23535,N_23714);
xor U23773 (N_23773,N_23715,N_23597);
nor U23774 (N_23774,N_23724,N_23605);
and U23775 (N_23775,N_23583,N_23555);
nor U23776 (N_23776,N_23607,N_23733);
nand U23777 (N_23777,N_23602,N_23650);
or U23778 (N_23778,N_23568,N_23592);
nand U23779 (N_23779,N_23646,N_23608);
or U23780 (N_23780,N_23667,N_23580);
nor U23781 (N_23781,N_23653,N_23675);
and U23782 (N_23782,N_23644,N_23711);
and U23783 (N_23783,N_23525,N_23591);
xnor U23784 (N_23784,N_23536,N_23679);
nor U23785 (N_23785,N_23722,N_23588);
nand U23786 (N_23786,N_23529,N_23682);
or U23787 (N_23787,N_23651,N_23517);
nand U23788 (N_23788,N_23730,N_23532);
and U23789 (N_23789,N_23515,N_23527);
or U23790 (N_23790,N_23640,N_23725);
and U23791 (N_23791,N_23507,N_23603);
and U23792 (N_23792,N_23659,N_23604);
nand U23793 (N_23793,N_23547,N_23561);
nor U23794 (N_23794,N_23501,N_23672);
nand U23795 (N_23795,N_23551,N_23745);
or U23796 (N_23796,N_23665,N_23528);
nand U23797 (N_23797,N_23731,N_23534);
xor U23798 (N_23798,N_23649,N_23617);
nor U23799 (N_23799,N_23674,N_23614);
and U23800 (N_23800,N_23531,N_23700);
or U23801 (N_23801,N_23626,N_23685);
or U23802 (N_23802,N_23690,N_23641);
nand U23803 (N_23803,N_23704,N_23557);
xor U23804 (N_23804,N_23643,N_23620);
nand U23805 (N_23805,N_23552,N_23579);
xnor U23806 (N_23806,N_23648,N_23743);
xor U23807 (N_23807,N_23634,N_23566);
or U23808 (N_23808,N_23619,N_23622);
xor U23809 (N_23809,N_23598,N_23741);
or U23810 (N_23810,N_23736,N_23574);
nor U23811 (N_23811,N_23642,N_23548);
and U23812 (N_23812,N_23625,N_23696);
nand U23813 (N_23813,N_23554,N_23739);
or U23814 (N_23814,N_23664,N_23508);
nand U23815 (N_23815,N_23697,N_23657);
and U23816 (N_23816,N_23587,N_23514);
xor U23817 (N_23817,N_23710,N_23709);
xnor U23818 (N_23818,N_23595,N_23567);
and U23819 (N_23819,N_23742,N_23593);
nand U23820 (N_23820,N_23689,N_23694);
nor U23821 (N_23821,N_23681,N_23523);
or U23822 (N_23822,N_23656,N_23590);
nand U23823 (N_23823,N_23570,N_23550);
nor U23824 (N_23824,N_23565,N_23575);
or U23825 (N_23825,N_23699,N_23668);
xnor U23826 (N_23826,N_23585,N_23613);
and U23827 (N_23827,N_23533,N_23718);
nor U23828 (N_23828,N_23546,N_23526);
or U23829 (N_23829,N_23695,N_23505);
nand U23830 (N_23830,N_23676,N_23717);
nand U23831 (N_23831,N_23701,N_23748);
and U23832 (N_23832,N_23734,N_23544);
or U23833 (N_23833,N_23584,N_23611);
nand U23834 (N_23834,N_23721,N_23606);
xnor U23835 (N_23835,N_23712,N_23594);
nor U23836 (N_23836,N_23596,N_23647);
xnor U23837 (N_23837,N_23673,N_23543);
nor U23838 (N_23838,N_23599,N_23581);
or U23839 (N_23839,N_23562,N_23662);
nor U23840 (N_23840,N_23702,N_23521);
and U23841 (N_23841,N_23577,N_23506);
or U23842 (N_23842,N_23637,N_23500);
nand U23843 (N_23843,N_23746,N_23658);
and U23844 (N_23844,N_23530,N_23616);
nor U23845 (N_23845,N_23513,N_23559);
nand U23846 (N_23846,N_23686,N_23660);
or U23847 (N_23847,N_23541,N_23693);
nor U23848 (N_23848,N_23688,N_23632);
and U23849 (N_23849,N_23589,N_23744);
nor U23850 (N_23850,N_23707,N_23601);
or U23851 (N_23851,N_23728,N_23537);
xnor U23852 (N_23852,N_23511,N_23539);
nor U23853 (N_23853,N_23504,N_23652);
and U23854 (N_23854,N_23666,N_23723);
nand U23855 (N_23855,N_23737,N_23558);
and U23856 (N_23856,N_23610,N_23684);
or U23857 (N_23857,N_23624,N_23691);
nand U23858 (N_23858,N_23687,N_23655);
xor U23859 (N_23859,N_23600,N_23720);
xnor U23860 (N_23860,N_23740,N_23661);
xnor U23861 (N_23861,N_23612,N_23582);
nor U23862 (N_23862,N_23628,N_23670);
and U23863 (N_23863,N_23677,N_23542);
nand U23864 (N_23864,N_23669,N_23645);
or U23865 (N_23865,N_23571,N_23631);
nand U23866 (N_23866,N_23564,N_23518);
xor U23867 (N_23867,N_23573,N_23522);
and U23868 (N_23868,N_23727,N_23716);
and U23869 (N_23869,N_23719,N_23671);
nand U23870 (N_23870,N_23747,N_23706);
nor U23871 (N_23871,N_23629,N_23549);
xnor U23872 (N_23872,N_23520,N_23749);
and U23873 (N_23873,N_23630,N_23502);
nor U23874 (N_23874,N_23509,N_23516);
and U23875 (N_23875,N_23655,N_23529);
nor U23876 (N_23876,N_23698,N_23564);
xor U23877 (N_23877,N_23679,N_23739);
xnor U23878 (N_23878,N_23503,N_23628);
or U23879 (N_23879,N_23509,N_23689);
nand U23880 (N_23880,N_23579,N_23732);
and U23881 (N_23881,N_23604,N_23672);
or U23882 (N_23882,N_23580,N_23504);
nand U23883 (N_23883,N_23597,N_23645);
or U23884 (N_23884,N_23636,N_23689);
nand U23885 (N_23885,N_23664,N_23715);
nand U23886 (N_23886,N_23582,N_23621);
nand U23887 (N_23887,N_23600,N_23616);
nor U23888 (N_23888,N_23624,N_23607);
nor U23889 (N_23889,N_23628,N_23728);
nor U23890 (N_23890,N_23674,N_23609);
and U23891 (N_23891,N_23550,N_23694);
and U23892 (N_23892,N_23700,N_23729);
nand U23893 (N_23893,N_23684,N_23718);
and U23894 (N_23894,N_23565,N_23692);
nor U23895 (N_23895,N_23616,N_23720);
nor U23896 (N_23896,N_23560,N_23628);
and U23897 (N_23897,N_23648,N_23741);
nor U23898 (N_23898,N_23562,N_23598);
xnor U23899 (N_23899,N_23658,N_23529);
or U23900 (N_23900,N_23537,N_23579);
or U23901 (N_23901,N_23629,N_23611);
or U23902 (N_23902,N_23601,N_23561);
xnor U23903 (N_23903,N_23565,N_23589);
nor U23904 (N_23904,N_23693,N_23578);
and U23905 (N_23905,N_23693,N_23611);
or U23906 (N_23906,N_23738,N_23660);
xnor U23907 (N_23907,N_23517,N_23504);
and U23908 (N_23908,N_23524,N_23621);
xor U23909 (N_23909,N_23521,N_23623);
xnor U23910 (N_23910,N_23617,N_23538);
or U23911 (N_23911,N_23553,N_23582);
and U23912 (N_23912,N_23703,N_23732);
or U23913 (N_23913,N_23533,N_23682);
or U23914 (N_23914,N_23533,N_23637);
and U23915 (N_23915,N_23639,N_23602);
and U23916 (N_23916,N_23577,N_23628);
and U23917 (N_23917,N_23725,N_23611);
nor U23918 (N_23918,N_23747,N_23538);
and U23919 (N_23919,N_23503,N_23647);
or U23920 (N_23920,N_23719,N_23702);
xnor U23921 (N_23921,N_23516,N_23557);
xor U23922 (N_23922,N_23659,N_23588);
or U23923 (N_23923,N_23615,N_23549);
and U23924 (N_23924,N_23546,N_23687);
nor U23925 (N_23925,N_23745,N_23523);
nor U23926 (N_23926,N_23603,N_23595);
nor U23927 (N_23927,N_23580,N_23569);
nand U23928 (N_23928,N_23595,N_23693);
nand U23929 (N_23929,N_23604,N_23715);
or U23930 (N_23930,N_23695,N_23500);
or U23931 (N_23931,N_23673,N_23721);
nand U23932 (N_23932,N_23670,N_23704);
and U23933 (N_23933,N_23528,N_23544);
xor U23934 (N_23934,N_23670,N_23539);
xor U23935 (N_23935,N_23686,N_23584);
and U23936 (N_23936,N_23680,N_23632);
nor U23937 (N_23937,N_23698,N_23645);
and U23938 (N_23938,N_23659,N_23559);
and U23939 (N_23939,N_23593,N_23576);
and U23940 (N_23940,N_23716,N_23563);
or U23941 (N_23941,N_23694,N_23604);
nand U23942 (N_23942,N_23562,N_23700);
xor U23943 (N_23943,N_23643,N_23665);
and U23944 (N_23944,N_23505,N_23582);
xnor U23945 (N_23945,N_23535,N_23644);
nor U23946 (N_23946,N_23741,N_23554);
nand U23947 (N_23947,N_23679,N_23651);
or U23948 (N_23948,N_23578,N_23575);
or U23949 (N_23949,N_23640,N_23647);
or U23950 (N_23950,N_23503,N_23566);
nand U23951 (N_23951,N_23687,N_23562);
and U23952 (N_23952,N_23551,N_23645);
xnor U23953 (N_23953,N_23524,N_23537);
nor U23954 (N_23954,N_23559,N_23594);
xor U23955 (N_23955,N_23548,N_23580);
xnor U23956 (N_23956,N_23601,N_23701);
xor U23957 (N_23957,N_23645,N_23592);
nand U23958 (N_23958,N_23632,N_23696);
nor U23959 (N_23959,N_23626,N_23565);
and U23960 (N_23960,N_23660,N_23652);
nor U23961 (N_23961,N_23540,N_23527);
and U23962 (N_23962,N_23631,N_23617);
and U23963 (N_23963,N_23638,N_23693);
or U23964 (N_23964,N_23657,N_23681);
and U23965 (N_23965,N_23647,N_23675);
xnor U23966 (N_23966,N_23673,N_23656);
xnor U23967 (N_23967,N_23609,N_23736);
nand U23968 (N_23968,N_23634,N_23668);
nor U23969 (N_23969,N_23714,N_23503);
xor U23970 (N_23970,N_23586,N_23672);
xnor U23971 (N_23971,N_23667,N_23701);
nor U23972 (N_23972,N_23658,N_23524);
nand U23973 (N_23973,N_23687,N_23584);
nor U23974 (N_23974,N_23590,N_23586);
nand U23975 (N_23975,N_23703,N_23540);
and U23976 (N_23976,N_23521,N_23745);
xor U23977 (N_23977,N_23617,N_23667);
xor U23978 (N_23978,N_23608,N_23628);
and U23979 (N_23979,N_23712,N_23626);
or U23980 (N_23980,N_23535,N_23518);
and U23981 (N_23981,N_23658,N_23689);
and U23982 (N_23982,N_23576,N_23560);
or U23983 (N_23983,N_23643,N_23534);
nor U23984 (N_23984,N_23566,N_23715);
nand U23985 (N_23985,N_23514,N_23745);
nand U23986 (N_23986,N_23555,N_23655);
xor U23987 (N_23987,N_23616,N_23529);
xnor U23988 (N_23988,N_23736,N_23600);
nor U23989 (N_23989,N_23659,N_23658);
xor U23990 (N_23990,N_23681,N_23640);
or U23991 (N_23991,N_23523,N_23716);
nor U23992 (N_23992,N_23748,N_23644);
or U23993 (N_23993,N_23536,N_23642);
nor U23994 (N_23994,N_23506,N_23744);
nor U23995 (N_23995,N_23654,N_23575);
xor U23996 (N_23996,N_23529,N_23574);
and U23997 (N_23997,N_23684,N_23541);
nor U23998 (N_23998,N_23747,N_23697);
or U23999 (N_23999,N_23693,N_23509);
nand U24000 (N_24000,N_23802,N_23878);
nand U24001 (N_24001,N_23914,N_23796);
and U24002 (N_24002,N_23947,N_23800);
or U24003 (N_24003,N_23877,N_23783);
xor U24004 (N_24004,N_23859,N_23979);
and U24005 (N_24005,N_23756,N_23797);
nor U24006 (N_24006,N_23827,N_23789);
xnor U24007 (N_24007,N_23932,N_23836);
or U24008 (N_24008,N_23821,N_23845);
and U24009 (N_24009,N_23940,N_23955);
and U24010 (N_24010,N_23790,N_23757);
nand U24011 (N_24011,N_23931,N_23772);
and U24012 (N_24012,N_23780,N_23822);
and U24013 (N_24013,N_23785,N_23776);
xor U24014 (N_24014,N_23963,N_23857);
xnor U24015 (N_24015,N_23766,N_23843);
and U24016 (N_24016,N_23812,N_23853);
nor U24017 (N_24017,N_23751,N_23846);
or U24018 (N_24018,N_23787,N_23909);
nand U24019 (N_24019,N_23786,N_23907);
nand U24020 (N_24020,N_23881,N_23788);
or U24021 (N_24021,N_23825,N_23828);
and U24022 (N_24022,N_23818,N_23806);
and U24023 (N_24023,N_23847,N_23960);
or U24024 (N_24024,N_23992,N_23837);
and U24025 (N_24025,N_23781,N_23918);
nor U24026 (N_24026,N_23950,N_23968);
and U24027 (N_24027,N_23880,N_23937);
and U24028 (N_24028,N_23978,N_23830);
or U24029 (N_24029,N_23867,N_23919);
nand U24030 (N_24030,N_23817,N_23905);
nor U24031 (N_24031,N_23993,N_23869);
nand U24032 (N_24032,N_23989,N_23858);
nor U24033 (N_24033,N_23910,N_23750);
xnor U24034 (N_24034,N_23906,N_23936);
and U24035 (N_24035,N_23799,N_23855);
and U24036 (N_24036,N_23754,N_23793);
or U24037 (N_24037,N_23770,N_23888);
nand U24038 (N_24038,N_23804,N_23969);
nand U24039 (N_24039,N_23927,N_23895);
nand U24040 (N_24040,N_23777,N_23798);
xnor U24041 (N_24041,N_23889,N_23985);
nand U24042 (N_24042,N_23928,N_23832);
or U24043 (N_24043,N_23807,N_23874);
and U24044 (N_24044,N_23782,N_23924);
nor U24045 (N_24045,N_23764,N_23856);
xor U24046 (N_24046,N_23941,N_23824);
nand U24047 (N_24047,N_23815,N_23850);
or U24048 (N_24048,N_23879,N_23916);
nand U24049 (N_24049,N_23994,N_23801);
xor U24050 (N_24050,N_23902,N_23819);
and U24051 (N_24051,N_23769,N_23943);
or U24052 (N_24052,N_23980,N_23935);
and U24053 (N_24053,N_23952,N_23860);
and U24054 (N_24054,N_23921,N_23840);
xor U24055 (N_24055,N_23765,N_23894);
or U24056 (N_24056,N_23987,N_23891);
nand U24057 (N_24057,N_23930,N_23873);
or U24058 (N_24058,N_23791,N_23938);
xor U24059 (N_24059,N_23976,N_23904);
nand U24060 (N_24060,N_23886,N_23755);
and U24061 (N_24061,N_23887,N_23792);
nand U24062 (N_24062,N_23851,N_23948);
or U24063 (N_24063,N_23820,N_23923);
nand U24064 (N_24064,N_23875,N_23839);
xnor U24065 (N_24065,N_23778,N_23883);
and U24066 (N_24066,N_23899,N_23865);
nand U24067 (N_24067,N_23920,N_23958);
xor U24068 (N_24068,N_23849,N_23934);
or U24069 (N_24069,N_23823,N_23962);
nand U24070 (N_24070,N_23771,N_23988);
nand U24071 (N_24071,N_23805,N_23926);
or U24072 (N_24072,N_23885,N_23946);
nor U24073 (N_24073,N_23949,N_23871);
or U24074 (N_24074,N_23774,N_23996);
and U24075 (N_24075,N_23997,N_23761);
and U24076 (N_24076,N_23763,N_23870);
and U24077 (N_24077,N_23752,N_23959);
or U24078 (N_24078,N_23898,N_23808);
nand U24079 (N_24079,N_23835,N_23896);
and U24080 (N_24080,N_23917,N_23912);
xnor U24081 (N_24081,N_23933,N_23861);
nor U24082 (N_24082,N_23762,N_23795);
nor U24083 (N_24083,N_23897,N_23901);
nor U24084 (N_24084,N_23779,N_23922);
or U24085 (N_24085,N_23977,N_23981);
and U24086 (N_24086,N_23939,N_23970);
xor U24087 (N_24087,N_23900,N_23951);
or U24088 (N_24088,N_23848,N_23942);
xor U24089 (N_24089,N_23834,N_23929);
nand U24090 (N_24090,N_23915,N_23925);
xnor U24091 (N_24091,N_23998,N_23999);
nand U24092 (N_24092,N_23954,N_23775);
and U24093 (N_24093,N_23967,N_23971);
nand U24094 (N_24094,N_23983,N_23831);
nor U24095 (N_24095,N_23768,N_23953);
and U24096 (N_24096,N_23957,N_23965);
or U24097 (N_24097,N_23813,N_23833);
and U24098 (N_24098,N_23913,N_23872);
nand U24099 (N_24099,N_23826,N_23986);
and U24100 (N_24100,N_23903,N_23829);
or U24101 (N_24101,N_23868,N_23841);
and U24102 (N_24102,N_23984,N_23784);
and U24103 (N_24103,N_23961,N_23884);
nor U24104 (N_24104,N_23966,N_23911);
nand U24105 (N_24105,N_23864,N_23995);
and U24106 (N_24106,N_23956,N_23852);
nor U24107 (N_24107,N_23892,N_23982);
xor U24108 (N_24108,N_23876,N_23973);
nor U24109 (N_24109,N_23866,N_23974);
or U24110 (N_24110,N_23814,N_23758);
or U24111 (N_24111,N_23862,N_23816);
nor U24112 (N_24112,N_23759,N_23972);
xnor U24113 (N_24113,N_23809,N_23991);
or U24114 (N_24114,N_23854,N_23810);
xor U24115 (N_24115,N_23863,N_23975);
or U24116 (N_24116,N_23893,N_23773);
nor U24117 (N_24117,N_23811,N_23753);
nand U24118 (N_24118,N_23944,N_23990);
nor U24119 (N_24119,N_23842,N_23838);
xor U24120 (N_24120,N_23882,N_23890);
nand U24121 (N_24121,N_23908,N_23794);
nand U24122 (N_24122,N_23964,N_23945);
xnor U24123 (N_24123,N_23844,N_23760);
or U24124 (N_24124,N_23767,N_23803);
and U24125 (N_24125,N_23750,N_23868);
nor U24126 (N_24126,N_23887,N_23982);
or U24127 (N_24127,N_23973,N_23824);
and U24128 (N_24128,N_23857,N_23770);
xor U24129 (N_24129,N_23885,N_23876);
xnor U24130 (N_24130,N_23987,N_23931);
xor U24131 (N_24131,N_23876,N_23986);
and U24132 (N_24132,N_23856,N_23775);
nand U24133 (N_24133,N_23775,N_23813);
nand U24134 (N_24134,N_23819,N_23948);
and U24135 (N_24135,N_23980,N_23834);
nor U24136 (N_24136,N_23806,N_23917);
xnor U24137 (N_24137,N_23998,N_23862);
or U24138 (N_24138,N_23821,N_23910);
nor U24139 (N_24139,N_23762,N_23976);
nor U24140 (N_24140,N_23930,N_23943);
nand U24141 (N_24141,N_23929,N_23843);
and U24142 (N_24142,N_23878,N_23947);
nand U24143 (N_24143,N_23939,N_23925);
nand U24144 (N_24144,N_23990,N_23900);
nor U24145 (N_24145,N_23827,N_23901);
and U24146 (N_24146,N_23915,N_23834);
xor U24147 (N_24147,N_23988,N_23763);
xor U24148 (N_24148,N_23930,N_23796);
nand U24149 (N_24149,N_23955,N_23821);
xor U24150 (N_24150,N_23889,N_23851);
nand U24151 (N_24151,N_23985,N_23846);
nand U24152 (N_24152,N_23851,N_23771);
or U24153 (N_24153,N_23930,N_23989);
xor U24154 (N_24154,N_23803,N_23827);
and U24155 (N_24155,N_23987,N_23885);
and U24156 (N_24156,N_23878,N_23774);
xor U24157 (N_24157,N_23986,N_23982);
and U24158 (N_24158,N_23861,N_23894);
nand U24159 (N_24159,N_23811,N_23792);
nand U24160 (N_24160,N_23805,N_23758);
nand U24161 (N_24161,N_23843,N_23948);
or U24162 (N_24162,N_23794,N_23789);
and U24163 (N_24163,N_23966,N_23994);
and U24164 (N_24164,N_23809,N_23889);
nand U24165 (N_24165,N_23855,N_23826);
nor U24166 (N_24166,N_23774,N_23956);
xor U24167 (N_24167,N_23940,N_23763);
or U24168 (N_24168,N_23861,N_23972);
nand U24169 (N_24169,N_23965,N_23906);
nor U24170 (N_24170,N_23800,N_23915);
xnor U24171 (N_24171,N_23824,N_23988);
nand U24172 (N_24172,N_23894,N_23919);
or U24173 (N_24173,N_23846,N_23955);
or U24174 (N_24174,N_23879,N_23824);
or U24175 (N_24175,N_23906,N_23778);
and U24176 (N_24176,N_23870,N_23987);
and U24177 (N_24177,N_23887,N_23779);
or U24178 (N_24178,N_23816,N_23805);
nand U24179 (N_24179,N_23816,N_23832);
and U24180 (N_24180,N_23885,N_23891);
or U24181 (N_24181,N_23867,N_23761);
nand U24182 (N_24182,N_23974,N_23860);
nand U24183 (N_24183,N_23839,N_23792);
or U24184 (N_24184,N_23813,N_23861);
and U24185 (N_24185,N_23862,N_23781);
and U24186 (N_24186,N_23993,N_23992);
or U24187 (N_24187,N_23822,N_23957);
nor U24188 (N_24188,N_23937,N_23906);
xnor U24189 (N_24189,N_23806,N_23864);
nand U24190 (N_24190,N_23755,N_23764);
nand U24191 (N_24191,N_23848,N_23780);
nand U24192 (N_24192,N_23946,N_23905);
or U24193 (N_24193,N_23894,N_23811);
or U24194 (N_24194,N_23828,N_23969);
and U24195 (N_24195,N_23912,N_23859);
nor U24196 (N_24196,N_23783,N_23892);
xnor U24197 (N_24197,N_23839,N_23793);
nand U24198 (N_24198,N_23979,N_23965);
or U24199 (N_24199,N_23953,N_23938);
or U24200 (N_24200,N_23974,N_23939);
and U24201 (N_24201,N_23960,N_23895);
or U24202 (N_24202,N_23928,N_23990);
xor U24203 (N_24203,N_23943,N_23879);
and U24204 (N_24204,N_23904,N_23887);
xor U24205 (N_24205,N_23763,N_23957);
nand U24206 (N_24206,N_23926,N_23960);
nand U24207 (N_24207,N_23979,N_23996);
xnor U24208 (N_24208,N_23786,N_23994);
xnor U24209 (N_24209,N_23910,N_23963);
or U24210 (N_24210,N_23763,N_23922);
or U24211 (N_24211,N_23922,N_23772);
and U24212 (N_24212,N_23868,N_23934);
nand U24213 (N_24213,N_23873,N_23825);
xnor U24214 (N_24214,N_23945,N_23805);
and U24215 (N_24215,N_23756,N_23767);
nor U24216 (N_24216,N_23849,N_23943);
xnor U24217 (N_24217,N_23773,N_23835);
xnor U24218 (N_24218,N_23884,N_23878);
nand U24219 (N_24219,N_23998,N_23958);
and U24220 (N_24220,N_23873,N_23918);
or U24221 (N_24221,N_23959,N_23870);
or U24222 (N_24222,N_23946,N_23928);
or U24223 (N_24223,N_23999,N_23830);
nor U24224 (N_24224,N_23831,N_23920);
and U24225 (N_24225,N_23980,N_23774);
nand U24226 (N_24226,N_23978,N_23828);
nand U24227 (N_24227,N_23939,N_23949);
nand U24228 (N_24228,N_23861,N_23838);
or U24229 (N_24229,N_23777,N_23939);
nand U24230 (N_24230,N_23987,N_23956);
or U24231 (N_24231,N_23890,N_23964);
xor U24232 (N_24232,N_23830,N_23918);
nand U24233 (N_24233,N_23888,N_23994);
nor U24234 (N_24234,N_23931,N_23926);
nor U24235 (N_24235,N_23914,N_23862);
nand U24236 (N_24236,N_23862,N_23853);
or U24237 (N_24237,N_23863,N_23761);
and U24238 (N_24238,N_23758,N_23916);
nand U24239 (N_24239,N_23975,N_23779);
or U24240 (N_24240,N_23857,N_23964);
xor U24241 (N_24241,N_23753,N_23821);
nor U24242 (N_24242,N_23771,N_23874);
nor U24243 (N_24243,N_23832,N_23763);
or U24244 (N_24244,N_23830,N_23814);
and U24245 (N_24245,N_23842,N_23975);
nand U24246 (N_24246,N_23908,N_23837);
nor U24247 (N_24247,N_23813,N_23960);
or U24248 (N_24248,N_23882,N_23798);
or U24249 (N_24249,N_23780,N_23804);
xor U24250 (N_24250,N_24039,N_24185);
or U24251 (N_24251,N_24009,N_24057);
nand U24252 (N_24252,N_24017,N_24180);
or U24253 (N_24253,N_24097,N_24157);
xnor U24254 (N_24254,N_24119,N_24102);
nor U24255 (N_24255,N_24012,N_24082);
xor U24256 (N_24256,N_24192,N_24048);
and U24257 (N_24257,N_24007,N_24058);
nand U24258 (N_24258,N_24055,N_24183);
nor U24259 (N_24259,N_24233,N_24123);
nand U24260 (N_24260,N_24236,N_24044);
and U24261 (N_24261,N_24224,N_24066);
and U24262 (N_24262,N_24244,N_24117);
nand U24263 (N_24263,N_24188,N_24127);
nand U24264 (N_24264,N_24161,N_24156);
xor U24265 (N_24265,N_24143,N_24249);
and U24266 (N_24266,N_24042,N_24096);
nor U24267 (N_24267,N_24028,N_24037);
nand U24268 (N_24268,N_24032,N_24003);
nor U24269 (N_24269,N_24235,N_24201);
nand U24270 (N_24270,N_24002,N_24225);
nor U24271 (N_24271,N_24166,N_24122);
nand U24272 (N_24272,N_24051,N_24172);
xor U24273 (N_24273,N_24021,N_24176);
xor U24274 (N_24274,N_24041,N_24214);
nand U24275 (N_24275,N_24070,N_24206);
nor U24276 (N_24276,N_24043,N_24147);
xnor U24277 (N_24277,N_24124,N_24047);
xor U24278 (N_24278,N_24113,N_24076);
or U24279 (N_24279,N_24030,N_24020);
or U24280 (N_24280,N_24005,N_24100);
or U24281 (N_24281,N_24241,N_24022);
xor U24282 (N_24282,N_24142,N_24075);
or U24283 (N_24283,N_24088,N_24212);
or U24284 (N_24284,N_24062,N_24167);
xor U24285 (N_24285,N_24160,N_24219);
nor U24286 (N_24286,N_24054,N_24046);
xor U24287 (N_24287,N_24171,N_24243);
nand U24288 (N_24288,N_24136,N_24248);
nor U24289 (N_24289,N_24145,N_24099);
or U24290 (N_24290,N_24178,N_24061);
or U24291 (N_24291,N_24036,N_24155);
xnor U24292 (N_24292,N_24013,N_24079);
nand U24293 (N_24293,N_24053,N_24239);
nand U24294 (N_24294,N_24000,N_24189);
nor U24295 (N_24295,N_24015,N_24050);
or U24296 (N_24296,N_24182,N_24121);
xnor U24297 (N_24297,N_24223,N_24218);
or U24298 (N_24298,N_24179,N_24129);
xnor U24299 (N_24299,N_24168,N_24184);
xnor U24300 (N_24300,N_24141,N_24023);
and U24301 (N_24301,N_24217,N_24073);
and U24302 (N_24302,N_24169,N_24133);
nor U24303 (N_24303,N_24247,N_24090);
nand U24304 (N_24304,N_24067,N_24210);
or U24305 (N_24305,N_24089,N_24240);
or U24306 (N_24306,N_24106,N_24229);
and U24307 (N_24307,N_24131,N_24052);
nand U24308 (N_24308,N_24034,N_24150);
nand U24309 (N_24309,N_24071,N_24152);
and U24310 (N_24310,N_24208,N_24220);
or U24311 (N_24311,N_24114,N_24010);
or U24312 (N_24312,N_24008,N_24056);
and U24313 (N_24313,N_24109,N_24033);
nor U24314 (N_24314,N_24011,N_24139);
nand U24315 (N_24315,N_24215,N_24221);
nand U24316 (N_24316,N_24019,N_24228);
and U24317 (N_24317,N_24081,N_24238);
nand U24318 (N_24318,N_24080,N_24181);
nand U24319 (N_24319,N_24092,N_24035);
nand U24320 (N_24320,N_24025,N_24198);
or U24321 (N_24321,N_24173,N_24196);
nand U24322 (N_24322,N_24091,N_24126);
and U24323 (N_24323,N_24191,N_24077);
xnor U24324 (N_24324,N_24083,N_24014);
nor U24325 (N_24325,N_24200,N_24027);
xnor U24326 (N_24326,N_24205,N_24232);
and U24327 (N_24327,N_24230,N_24004);
xnor U24328 (N_24328,N_24163,N_24105);
or U24329 (N_24329,N_24207,N_24153);
and U24330 (N_24330,N_24199,N_24065);
nor U24331 (N_24331,N_24064,N_24060);
or U24332 (N_24332,N_24197,N_24068);
xor U24333 (N_24333,N_24149,N_24135);
xor U24334 (N_24334,N_24137,N_24138);
or U24335 (N_24335,N_24024,N_24162);
or U24336 (N_24336,N_24242,N_24111);
and U24337 (N_24337,N_24087,N_24193);
nor U24338 (N_24338,N_24158,N_24186);
and U24339 (N_24339,N_24174,N_24148);
nor U24340 (N_24340,N_24170,N_24072);
nor U24341 (N_24341,N_24098,N_24226);
nor U24342 (N_24342,N_24222,N_24078);
nor U24343 (N_24343,N_24095,N_24118);
and U24344 (N_24344,N_24016,N_24209);
nand U24345 (N_24345,N_24040,N_24069);
xnor U24346 (N_24346,N_24026,N_24038);
nand U24347 (N_24347,N_24175,N_24063);
xnor U24348 (N_24348,N_24154,N_24108);
or U24349 (N_24349,N_24125,N_24132);
nor U24350 (N_24350,N_24202,N_24134);
or U24351 (N_24351,N_24001,N_24246);
or U24352 (N_24352,N_24049,N_24146);
nor U24353 (N_24353,N_24194,N_24128);
or U24354 (N_24354,N_24045,N_24074);
or U24355 (N_24355,N_24227,N_24187);
nor U24356 (N_24356,N_24140,N_24164);
nor U24357 (N_24357,N_24195,N_24101);
or U24358 (N_24358,N_24085,N_24204);
and U24359 (N_24359,N_24144,N_24177);
xnor U24360 (N_24360,N_24059,N_24165);
nor U24361 (N_24361,N_24213,N_24211);
and U24362 (N_24362,N_24029,N_24086);
nand U24363 (N_24363,N_24031,N_24006);
nand U24364 (N_24364,N_24120,N_24231);
nor U24365 (N_24365,N_24112,N_24159);
nand U24366 (N_24366,N_24190,N_24018);
nor U24367 (N_24367,N_24116,N_24104);
nand U24368 (N_24368,N_24203,N_24115);
and U24369 (N_24369,N_24237,N_24110);
and U24370 (N_24370,N_24103,N_24245);
or U24371 (N_24371,N_24216,N_24130);
or U24372 (N_24372,N_24084,N_24234);
and U24373 (N_24373,N_24093,N_24151);
xor U24374 (N_24374,N_24107,N_24094);
nor U24375 (N_24375,N_24098,N_24033);
or U24376 (N_24376,N_24048,N_24081);
or U24377 (N_24377,N_24034,N_24039);
nand U24378 (N_24378,N_24245,N_24084);
nor U24379 (N_24379,N_24021,N_24028);
and U24380 (N_24380,N_24247,N_24211);
and U24381 (N_24381,N_24146,N_24136);
or U24382 (N_24382,N_24012,N_24182);
or U24383 (N_24383,N_24108,N_24023);
or U24384 (N_24384,N_24100,N_24060);
nand U24385 (N_24385,N_24009,N_24077);
xor U24386 (N_24386,N_24067,N_24069);
nand U24387 (N_24387,N_24145,N_24231);
or U24388 (N_24388,N_24036,N_24171);
or U24389 (N_24389,N_24011,N_24175);
xor U24390 (N_24390,N_24170,N_24178);
or U24391 (N_24391,N_24172,N_24042);
and U24392 (N_24392,N_24225,N_24135);
nor U24393 (N_24393,N_24082,N_24056);
nor U24394 (N_24394,N_24014,N_24091);
xor U24395 (N_24395,N_24122,N_24149);
nand U24396 (N_24396,N_24052,N_24057);
nor U24397 (N_24397,N_24060,N_24184);
xor U24398 (N_24398,N_24064,N_24173);
nand U24399 (N_24399,N_24237,N_24212);
xor U24400 (N_24400,N_24016,N_24085);
or U24401 (N_24401,N_24190,N_24093);
nor U24402 (N_24402,N_24034,N_24226);
nand U24403 (N_24403,N_24247,N_24078);
and U24404 (N_24404,N_24141,N_24170);
xnor U24405 (N_24405,N_24074,N_24008);
and U24406 (N_24406,N_24072,N_24076);
or U24407 (N_24407,N_24243,N_24233);
xnor U24408 (N_24408,N_24187,N_24025);
and U24409 (N_24409,N_24006,N_24212);
or U24410 (N_24410,N_24225,N_24003);
and U24411 (N_24411,N_24197,N_24141);
or U24412 (N_24412,N_24177,N_24097);
xnor U24413 (N_24413,N_24024,N_24084);
and U24414 (N_24414,N_24091,N_24165);
nand U24415 (N_24415,N_24000,N_24206);
and U24416 (N_24416,N_24021,N_24119);
or U24417 (N_24417,N_24054,N_24005);
or U24418 (N_24418,N_24057,N_24243);
xor U24419 (N_24419,N_24037,N_24175);
and U24420 (N_24420,N_24160,N_24214);
and U24421 (N_24421,N_24211,N_24045);
nand U24422 (N_24422,N_24199,N_24114);
nand U24423 (N_24423,N_24190,N_24067);
xnor U24424 (N_24424,N_24065,N_24135);
nor U24425 (N_24425,N_24107,N_24141);
and U24426 (N_24426,N_24067,N_24103);
or U24427 (N_24427,N_24055,N_24175);
or U24428 (N_24428,N_24035,N_24227);
nor U24429 (N_24429,N_24040,N_24166);
nand U24430 (N_24430,N_24173,N_24236);
or U24431 (N_24431,N_24240,N_24058);
nor U24432 (N_24432,N_24008,N_24146);
nand U24433 (N_24433,N_24225,N_24183);
nor U24434 (N_24434,N_24058,N_24232);
xnor U24435 (N_24435,N_24116,N_24208);
and U24436 (N_24436,N_24026,N_24125);
xor U24437 (N_24437,N_24197,N_24092);
nand U24438 (N_24438,N_24011,N_24214);
nor U24439 (N_24439,N_24162,N_24198);
and U24440 (N_24440,N_24074,N_24012);
and U24441 (N_24441,N_24248,N_24114);
nor U24442 (N_24442,N_24133,N_24161);
xor U24443 (N_24443,N_24078,N_24243);
and U24444 (N_24444,N_24069,N_24192);
or U24445 (N_24445,N_24076,N_24186);
and U24446 (N_24446,N_24045,N_24005);
and U24447 (N_24447,N_24120,N_24079);
and U24448 (N_24448,N_24200,N_24129);
nand U24449 (N_24449,N_24071,N_24101);
and U24450 (N_24450,N_24158,N_24137);
xnor U24451 (N_24451,N_24104,N_24087);
nor U24452 (N_24452,N_24012,N_24046);
and U24453 (N_24453,N_24031,N_24093);
and U24454 (N_24454,N_24020,N_24214);
xnor U24455 (N_24455,N_24242,N_24203);
or U24456 (N_24456,N_24093,N_24243);
nand U24457 (N_24457,N_24197,N_24073);
or U24458 (N_24458,N_24031,N_24009);
nand U24459 (N_24459,N_24125,N_24033);
nor U24460 (N_24460,N_24117,N_24068);
nand U24461 (N_24461,N_24040,N_24071);
nand U24462 (N_24462,N_24115,N_24188);
and U24463 (N_24463,N_24034,N_24153);
xnor U24464 (N_24464,N_24249,N_24132);
or U24465 (N_24465,N_24218,N_24063);
xnor U24466 (N_24466,N_24218,N_24109);
or U24467 (N_24467,N_24166,N_24139);
nand U24468 (N_24468,N_24004,N_24231);
and U24469 (N_24469,N_24134,N_24050);
nand U24470 (N_24470,N_24207,N_24055);
nand U24471 (N_24471,N_24188,N_24205);
nand U24472 (N_24472,N_24130,N_24109);
or U24473 (N_24473,N_24017,N_24048);
or U24474 (N_24474,N_24248,N_24165);
nand U24475 (N_24475,N_24123,N_24045);
xor U24476 (N_24476,N_24075,N_24131);
nand U24477 (N_24477,N_24001,N_24096);
xor U24478 (N_24478,N_24085,N_24099);
nor U24479 (N_24479,N_24103,N_24206);
nand U24480 (N_24480,N_24053,N_24179);
nor U24481 (N_24481,N_24116,N_24085);
nor U24482 (N_24482,N_24061,N_24163);
nor U24483 (N_24483,N_24150,N_24148);
nor U24484 (N_24484,N_24018,N_24010);
and U24485 (N_24485,N_24194,N_24021);
xor U24486 (N_24486,N_24155,N_24101);
nor U24487 (N_24487,N_24097,N_24129);
nor U24488 (N_24488,N_24225,N_24078);
or U24489 (N_24489,N_24102,N_24129);
or U24490 (N_24490,N_24003,N_24045);
xnor U24491 (N_24491,N_24130,N_24218);
or U24492 (N_24492,N_24137,N_24103);
nand U24493 (N_24493,N_24249,N_24169);
nand U24494 (N_24494,N_24111,N_24076);
nand U24495 (N_24495,N_24226,N_24024);
xnor U24496 (N_24496,N_24209,N_24131);
nand U24497 (N_24497,N_24192,N_24231);
or U24498 (N_24498,N_24095,N_24244);
nand U24499 (N_24499,N_24143,N_24021);
nor U24500 (N_24500,N_24337,N_24462);
or U24501 (N_24501,N_24445,N_24361);
and U24502 (N_24502,N_24269,N_24342);
nand U24503 (N_24503,N_24378,N_24453);
and U24504 (N_24504,N_24341,N_24356);
nand U24505 (N_24505,N_24321,N_24432);
or U24506 (N_24506,N_24431,N_24355);
or U24507 (N_24507,N_24472,N_24409);
or U24508 (N_24508,N_24314,N_24480);
and U24509 (N_24509,N_24438,N_24497);
xnor U24510 (N_24510,N_24304,N_24452);
xnor U24511 (N_24511,N_24275,N_24411);
xnor U24512 (N_24512,N_24448,N_24490);
xor U24513 (N_24513,N_24426,N_24360);
xor U24514 (N_24514,N_24352,N_24386);
and U24515 (N_24515,N_24493,N_24464);
nor U24516 (N_24516,N_24371,N_24329);
or U24517 (N_24517,N_24330,N_24351);
nor U24518 (N_24518,N_24383,N_24469);
nor U24519 (N_24519,N_24297,N_24403);
and U24520 (N_24520,N_24289,N_24325);
or U24521 (N_24521,N_24447,N_24475);
nand U24522 (N_24522,N_24473,N_24307);
or U24523 (N_24523,N_24394,N_24320);
and U24524 (N_24524,N_24488,N_24486);
or U24525 (N_24525,N_24332,N_24368);
nor U24526 (N_24526,N_24279,N_24293);
and U24527 (N_24527,N_24465,N_24422);
xor U24528 (N_24528,N_24415,N_24471);
nand U24529 (N_24529,N_24366,N_24449);
xnor U24530 (N_24530,N_24463,N_24260);
xnor U24531 (N_24531,N_24272,N_24308);
xnor U24532 (N_24532,N_24306,N_24292);
and U24533 (N_24533,N_24347,N_24285);
xor U24534 (N_24534,N_24435,N_24429);
xor U24535 (N_24535,N_24310,N_24345);
nand U24536 (N_24536,N_24499,N_24282);
nand U24537 (N_24537,N_24414,N_24397);
nor U24538 (N_24538,N_24377,N_24401);
nor U24539 (N_24539,N_24333,N_24494);
nand U24540 (N_24540,N_24468,N_24420);
xnor U24541 (N_24541,N_24461,N_24322);
and U24542 (N_24542,N_24258,N_24387);
nand U24543 (N_24543,N_24391,N_24417);
xnor U24544 (N_24544,N_24287,N_24267);
xnor U24545 (N_24545,N_24425,N_24340);
nand U24546 (N_24546,N_24412,N_24353);
and U24547 (N_24547,N_24479,N_24358);
or U24548 (N_24548,N_24410,N_24354);
nand U24549 (N_24549,N_24393,N_24338);
xnor U24550 (N_24550,N_24441,N_24348);
nor U24551 (N_24551,N_24444,N_24362);
xor U24552 (N_24552,N_24492,N_24263);
nor U24553 (N_24553,N_24323,N_24266);
nor U24554 (N_24554,N_24481,N_24373);
xor U24555 (N_24555,N_24288,N_24419);
nor U24556 (N_24556,N_24390,N_24319);
nand U24557 (N_24557,N_24396,N_24395);
nor U24558 (N_24558,N_24485,N_24498);
or U24559 (N_24559,N_24359,N_24392);
nor U24560 (N_24560,N_24489,N_24376);
and U24561 (N_24561,N_24398,N_24335);
nand U24562 (N_24562,N_24311,N_24271);
xor U24563 (N_24563,N_24291,N_24389);
or U24564 (N_24564,N_24264,N_24384);
and U24565 (N_24565,N_24300,N_24303);
and U24566 (N_24566,N_24428,N_24433);
and U24567 (N_24567,N_24459,N_24456);
or U24568 (N_24568,N_24331,N_24370);
nand U24569 (N_24569,N_24446,N_24413);
and U24570 (N_24570,N_24343,N_24262);
nand U24571 (N_24571,N_24315,N_24408);
nor U24572 (N_24572,N_24457,N_24309);
and U24573 (N_24573,N_24295,N_24455);
and U24574 (N_24574,N_24430,N_24402);
or U24575 (N_24575,N_24277,N_24301);
xnor U24576 (N_24576,N_24252,N_24367);
or U24577 (N_24577,N_24484,N_24339);
or U24578 (N_24578,N_24405,N_24253);
or U24579 (N_24579,N_24369,N_24491);
xnor U24580 (N_24580,N_24372,N_24458);
or U24581 (N_24581,N_24443,N_24364);
nand U24582 (N_24582,N_24278,N_24363);
and U24583 (N_24583,N_24296,N_24427);
xnor U24584 (N_24584,N_24424,N_24406);
and U24585 (N_24585,N_24284,N_24460);
xor U24586 (N_24586,N_24294,N_24254);
or U24587 (N_24587,N_24313,N_24283);
or U24588 (N_24588,N_24299,N_24326);
nand U24589 (N_24589,N_24451,N_24440);
nand U24590 (N_24590,N_24281,N_24434);
and U24591 (N_24591,N_24344,N_24316);
or U24592 (N_24592,N_24379,N_24467);
xnor U24593 (N_24593,N_24381,N_24251);
nor U24594 (N_24594,N_24404,N_24317);
xnor U24595 (N_24595,N_24286,N_24436);
or U24596 (N_24596,N_24375,N_24273);
xor U24597 (N_24597,N_24302,N_24482);
nor U24598 (N_24598,N_24478,N_24385);
nor U24599 (N_24599,N_24407,N_24418);
or U24600 (N_24600,N_24268,N_24399);
xnor U24601 (N_24601,N_24466,N_24265);
and U24602 (N_24602,N_24483,N_24327);
xnor U24603 (N_24603,N_24290,N_24346);
xor U24604 (N_24604,N_24380,N_24350);
and U24605 (N_24605,N_24357,N_24334);
nand U24606 (N_24606,N_24280,N_24476);
xnor U24607 (N_24607,N_24470,N_24274);
nor U24608 (N_24608,N_24442,N_24382);
or U24609 (N_24609,N_24305,N_24324);
nand U24610 (N_24610,N_24450,N_24259);
and U24611 (N_24611,N_24423,N_24250);
nor U24612 (N_24612,N_24276,N_24270);
and U24613 (N_24613,N_24374,N_24454);
and U24614 (N_24614,N_24400,N_24328);
or U24615 (N_24615,N_24477,N_24261);
xor U24616 (N_24616,N_24388,N_24439);
or U24617 (N_24617,N_24349,N_24257);
nand U24618 (N_24618,N_24474,N_24255);
nor U24619 (N_24619,N_24312,N_24487);
and U24620 (N_24620,N_24365,N_24437);
or U24621 (N_24621,N_24421,N_24495);
or U24622 (N_24622,N_24256,N_24416);
nand U24623 (N_24623,N_24336,N_24318);
or U24624 (N_24624,N_24298,N_24496);
xor U24625 (N_24625,N_24284,N_24368);
nand U24626 (N_24626,N_24483,N_24469);
and U24627 (N_24627,N_24410,N_24451);
and U24628 (N_24628,N_24449,N_24308);
and U24629 (N_24629,N_24433,N_24344);
and U24630 (N_24630,N_24323,N_24327);
and U24631 (N_24631,N_24266,N_24343);
xnor U24632 (N_24632,N_24455,N_24277);
xnor U24633 (N_24633,N_24259,N_24301);
nand U24634 (N_24634,N_24331,N_24441);
nand U24635 (N_24635,N_24340,N_24447);
or U24636 (N_24636,N_24450,N_24432);
or U24637 (N_24637,N_24463,N_24437);
and U24638 (N_24638,N_24497,N_24498);
nand U24639 (N_24639,N_24480,N_24404);
nand U24640 (N_24640,N_24280,N_24342);
or U24641 (N_24641,N_24428,N_24358);
nand U24642 (N_24642,N_24404,N_24289);
nor U24643 (N_24643,N_24371,N_24314);
and U24644 (N_24644,N_24443,N_24296);
nand U24645 (N_24645,N_24462,N_24276);
or U24646 (N_24646,N_24378,N_24432);
xnor U24647 (N_24647,N_24310,N_24435);
nand U24648 (N_24648,N_24327,N_24367);
nand U24649 (N_24649,N_24331,N_24276);
nand U24650 (N_24650,N_24410,N_24425);
nor U24651 (N_24651,N_24415,N_24447);
xnor U24652 (N_24652,N_24343,N_24289);
xnor U24653 (N_24653,N_24324,N_24342);
or U24654 (N_24654,N_24384,N_24428);
xnor U24655 (N_24655,N_24378,N_24369);
nand U24656 (N_24656,N_24386,N_24473);
and U24657 (N_24657,N_24486,N_24466);
xor U24658 (N_24658,N_24468,N_24261);
xor U24659 (N_24659,N_24299,N_24305);
xnor U24660 (N_24660,N_24307,N_24271);
xnor U24661 (N_24661,N_24408,N_24328);
or U24662 (N_24662,N_24331,N_24419);
nand U24663 (N_24663,N_24306,N_24372);
xor U24664 (N_24664,N_24488,N_24329);
nor U24665 (N_24665,N_24497,N_24263);
or U24666 (N_24666,N_24479,N_24413);
and U24667 (N_24667,N_24301,N_24408);
nand U24668 (N_24668,N_24294,N_24280);
nand U24669 (N_24669,N_24264,N_24318);
xnor U24670 (N_24670,N_24361,N_24435);
nand U24671 (N_24671,N_24346,N_24328);
nand U24672 (N_24672,N_24480,N_24377);
nor U24673 (N_24673,N_24398,N_24452);
or U24674 (N_24674,N_24252,N_24262);
nor U24675 (N_24675,N_24436,N_24414);
nor U24676 (N_24676,N_24288,N_24287);
nor U24677 (N_24677,N_24424,N_24440);
or U24678 (N_24678,N_24350,N_24383);
nand U24679 (N_24679,N_24297,N_24255);
nor U24680 (N_24680,N_24289,N_24314);
nand U24681 (N_24681,N_24440,N_24386);
or U24682 (N_24682,N_24373,N_24494);
and U24683 (N_24683,N_24372,N_24349);
and U24684 (N_24684,N_24340,N_24444);
nand U24685 (N_24685,N_24442,N_24370);
and U24686 (N_24686,N_24293,N_24262);
and U24687 (N_24687,N_24467,N_24403);
or U24688 (N_24688,N_24327,N_24383);
xnor U24689 (N_24689,N_24251,N_24417);
nand U24690 (N_24690,N_24282,N_24303);
or U24691 (N_24691,N_24317,N_24258);
or U24692 (N_24692,N_24446,N_24345);
nand U24693 (N_24693,N_24274,N_24325);
nor U24694 (N_24694,N_24378,N_24423);
nand U24695 (N_24695,N_24308,N_24269);
xnor U24696 (N_24696,N_24271,N_24492);
or U24697 (N_24697,N_24451,N_24462);
nor U24698 (N_24698,N_24342,N_24374);
and U24699 (N_24699,N_24287,N_24367);
xnor U24700 (N_24700,N_24357,N_24478);
nor U24701 (N_24701,N_24259,N_24390);
and U24702 (N_24702,N_24279,N_24258);
and U24703 (N_24703,N_24370,N_24429);
xor U24704 (N_24704,N_24362,N_24405);
xnor U24705 (N_24705,N_24373,N_24325);
xor U24706 (N_24706,N_24382,N_24287);
or U24707 (N_24707,N_24303,N_24396);
nor U24708 (N_24708,N_24475,N_24409);
nand U24709 (N_24709,N_24357,N_24331);
xnor U24710 (N_24710,N_24340,N_24400);
nor U24711 (N_24711,N_24443,N_24327);
xor U24712 (N_24712,N_24418,N_24296);
nor U24713 (N_24713,N_24479,N_24320);
nand U24714 (N_24714,N_24365,N_24291);
and U24715 (N_24715,N_24291,N_24362);
nand U24716 (N_24716,N_24468,N_24301);
xnor U24717 (N_24717,N_24385,N_24329);
and U24718 (N_24718,N_24342,N_24276);
nand U24719 (N_24719,N_24476,N_24263);
and U24720 (N_24720,N_24465,N_24262);
xnor U24721 (N_24721,N_24457,N_24275);
nand U24722 (N_24722,N_24423,N_24293);
nor U24723 (N_24723,N_24388,N_24413);
or U24724 (N_24724,N_24365,N_24419);
or U24725 (N_24725,N_24265,N_24261);
and U24726 (N_24726,N_24405,N_24415);
or U24727 (N_24727,N_24311,N_24270);
nand U24728 (N_24728,N_24346,N_24261);
and U24729 (N_24729,N_24352,N_24419);
or U24730 (N_24730,N_24288,N_24396);
xnor U24731 (N_24731,N_24410,N_24465);
xor U24732 (N_24732,N_24466,N_24464);
or U24733 (N_24733,N_24329,N_24261);
and U24734 (N_24734,N_24299,N_24321);
xor U24735 (N_24735,N_24488,N_24322);
and U24736 (N_24736,N_24367,N_24402);
nor U24737 (N_24737,N_24367,N_24405);
and U24738 (N_24738,N_24310,N_24401);
nor U24739 (N_24739,N_24250,N_24348);
nor U24740 (N_24740,N_24408,N_24387);
nor U24741 (N_24741,N_24253,N_24275);
xor U24742 (N_24742,N_24283,N_24476);
nor U24743 (N_24743,N_24275,N_24339);
nor U24744 (N_24744,N_24444,N_24369);
or U24745 (N_24745,N_24475,N_24305);
nor U24746 (N_24746,N_24298,N_24479);
xor U24747 (N_24747,N_24342,N_24464);
xnor U24748 (N_24748,N_24339,N_24362);
xor U24749 (N_24749,N_24361,N_24437);
nor U24750 (N_24750,N_24621,N_24518);
or U24751 (N_24751,N_24735,N_24656);
xnor U24752 (N_24752,N_24536,N_24626);
or U24753 (N_24753,N_24602,N_24614);
nand U24754 (N_24754,N_24516,N_24574);
nor U24755 (N_24755,N_24661,N_24500);
and U24756 (N_24756,N_24540,N_24640);
nor U24757 (N_24757,N_24731,N_24634);
nor U24758 (N_24758,N_24583,N_24562);
nand U24759 (N_24759,N_24742,N_24556);
and U24760 (N_24760,N_24607,N_24718);
or U24761 (N_24761,N_24561,N_24748);
xnor U24762 (N_24762,N_24557,N_24563);
nand U24763 (N_24763,N_24542,N_24527);
nand U24764 (N_24764,N_24631,N_24613);
or U24765 (N_24765,N_24593,N_24615);
xor U24766 (N_24766,N_24658,N_24676);
nor U24767 (N_24767,N_24598,N_24530);
and U24768 (N_24768,N_24618,N_24700);
and U24769 (N_24769,N_24665,N_24649);
and U24770 (N_24770,N_24708,N_24739);
nor U24771 (N_24771,N_24571,N_24539);
and U24772 (N_24772,N_24732,N_24682);
or U24773 (N_24773,N_24501,N_24701);
and U24774 (N_24774,N_24715,N_24720);
nor U24775 (N_24775,N_24669,N_24528);
nand U24776 (N_24776,N_24508,N_24589);
and U24777 (N_24777,N_24622,N_24605);
xnor U24778 (N_24778,N_24723,N_24675);
nand U24779 (N_24779,N_24670,N_24729);
xnor U24780 (N_24780,N_24570,N_24654);
or U24781 (N_24781,N_24509,N_24623);
and U24782 (N_24782,N_24599,N_24687);
and U24783 (N_24783,N_24513,N_24688);
nand U24784 (N_24784,N_24624,N_24514);
nor U24785 (N_24785,N_24625,N_24657);
nor U24786 (N_24786,N_24600,N_24722);
nand U24787 (N_24787,N_24512,N_24653);
nor U24788 (N_24788,N_24719,N_24597);
nand U24789 (N_24789,N_24726,N_24585);
xor U24790 (N_24790,N_24525,N_24523);
and U24791 (N_24791,N_24677,N_24587);
nand U24792 (N_24792,N_24660,N_24672);
nor U24793 (N_24793,N_24590,N_24695);
or U24794 (N_24794,N_24546,N_24667);
xor U24795 (N_24795,N_24572,N_24681);
nand U24796 (N_24796,N_24633,N_24703);
and U24797 (N_24797,N_24646,N_24713);
or U24798 (N_24798,N_24537,N_24548);
nor U24799 (N_24799,N_24588,N_24610);
xnor U24800 (N_24800,N_24573,N_24521);
nor U24801 (N_24801,N_24679,N_24690);
nor U24802 (N_24802,N_24745,N_24650);
or U24803 (N_24803,N_24747,N_24707);
or U24804 (N_24804,N_24741,N_24705);
xnor U24805 (N_24805,N_24533,N_24566);
or U24806 (N_24806,N_24706,N_24689);
and U24807 (N_24807,N_24738,N_24697);
xnor U24808 (N_24808,N_24730,N_24692);
nand U24809 (N_24809,N_24520,N_24505);
xnor U24810 (N_24810,N_24596,N_24532);
or U24811 (N_24811,N_24642,N_24616);
xnor U24812 (N_24812,N_24611,N_24538);
or U24813 (N_24813,N_24645,N_24734);
nand U24814 (N_24814,N_24647,N_24552);
and U24815 (N_24815,N_24641,N_24567);
nor U24816 (N_24816,N_24511,N_24629);
xnor U24817 (N_24817,N_24673,N_24635);
nand U24818 (N_24818,N_24560,N_24603);
xnor U24819 (N_24819,N_24709,N_24643);
xor U24820 (N_24820,N_24666,N_24724);
or U24821 (N_24821,N_24699,N_24693);
and U24822 (N_24822,N_24659,N_24502);
or U24823 (N_24823,N_24584,N_24606);
or U24824 (N_24824,N_24721,N_24619);
and U24825 (N_24825,N_24569,N_24651);
nand U24826 (N_24826,N_24579,N_24627);
nor U24827 (N_24827,N_24683,N_24694);
nor U24828 (N_24828,N_24522,N_24652);
nand U24829 (N_24829,N_24506,N_24737);
nand U24830 (N_24830,N_24534,N_24524);
nand U24831 (N_24831,N_24507,N_24517);
and U24832 (N_24832,N_24743,N_24663);
xnor U24833 (N_24833,N_24549,N_24685);
nor U24834 (N_24834,N_24580,N_24620);
or U24835 (N_24835,N_24578,N_24725);
nand U24836 (N_24836,N_24728,N_24577);
nand U24837 (N_24837,N_24655,N_24740);
xor U24838 (N_24838,N_24591,N_24541);
nand U24839 (N_24839,N_24559,N_24550);
nand U24840 (N_24840,N_24733,N_24581);
xnor U24841 (N_24841,N_24630,N_24531);
xnor U24842 (N_24842,N_24608,N_24671);
and U24843 (N_24843,N_24717,N_24503);
nand U24844 (N_24844,N_24637,N_24736);
and U24845 (N_24845,N_24547,N_24594);
nor U24846 (N_24846,N_24696,N_24568);
xnor U24847 (N_24847,N_24555,N_24691);
or U24848 (N_24848,N_24698,N_24526);
and U24849 (N_24849,N_24680,N_24586);
nand U24850 (N_24850,N_24544,N_24749);
nand U24851 (N_24851,N_24716,N_24575);
xnor U24852 (N_24852,N_24515,N_24553);
nor U24853 (N_24853,N_24564,N_24648);
or U24854 (N_24854,N_24558,N_24636);
and U24855 (N_24855,N_24639,N_24710);
nand U24856 (N_24856,N_24576,N_24628);
nor U24857 (N_24857,N_24711,N_24668);
xor U24858 (N_24858,N_24545,N_24612);
nand U24859 (N_24859,N_24529,N_24674);
nor U24860 (N_24860,N_24678,N_24592);
nor U24861 (N_24861,N_24686,N_24543);
or U24862 (N_24862,N_24644,N_24714);
nor U24863 (N_24863,N_24504,N_24609);
nor U24864 (N_24864,N_24535,N_24604);
nand U24865 (N_24865,N_24664,N_24601);
or U24866 (N_24866,N_24510,N_24617);
and U24867 (N_24867,N_24554,N_24519);
xor U24868 (N_24868,N_24551,N_24632);
and U24869 (N_24869,N_24727,N_24595);
or U24870 (N_24870,N_24582,N_24744);
or U24871 (N_24871,N_24638,N_24662);
and U24872 (N_24872,N_24684,N_24712);
and U24873 (N_24873,N_24704,N_24565);
or U24874 (N_24874,N_24746,N_24702);
xor U24875 (N_24875,N_24639,N_24550);
and U24876 (N_24876,N_24619,N_24507);
and U24877 (N_24877,N_24691,N_24536);
and U24878 (N_24878,N_24516,N_24538);
nand U24879 (N_24879,N_24594,N_24526);
and U24880 (N_24880,N_24569,N_24719);
nand U24881 (N_24881,N_24503,N_24683);
xor U24882 (N_24882,N_24719,N_24506);
and U24883 (N_24883,N_24649,N_24630);
nor U24884 (N_24884,N_24555,N_24605);
xnor U24885 (N_24885,N_24597,N_24582);
nand U24886 (N_24886,N_24628,N_24655);
nor U24887 (N_24887,N_24558,N_24601);
xor U24888 (N_24888,N_24744,N_24567);
nand U24889 (N_24889,N_24661,N_24606);
or U24890 (N_24890,N_24735,N_24593);
nor U24891 (N_24891,N_24690,N_24718);
or U24892 (N_24892,N_24727,N_24725);
nor U24893 (N_24893,N_24678,N_24508);
xnor U24894 (N_24894,N_24749,N_24733);
xor U24895 (N_24895,N_24558,N_24603);
and U24896 (N_24896,N_24581,N_24720);
xnor U24897 (N_24897,N_24650,N_24679);
nand U24898 (N_24898,N_24536,N_24528);
and U24899 (N_24899,N_24506,N_24749);
xor U24900 (N_24900,N_24617,N_24597);
nand U24901 (N_24901,N_24701,N_24708);
nand U24902 (N_24902,N_24694,N_24657);
xnor U24903 (N_24903,N_24628,N_24724);
or U24904 (N_24904,N_24658,N_24574);
nor U24905 (N_24905,N_24675,N_24557);
xor U24906 (N_24906,N_24568,N_24594);
or U24907 (N_24907,N_24645,N_24658);
or U24908 (N_24908,N_24667,N_24561);
and U24909 (N_24909,N_24572,N_24590);
nand U24910 (N_24910,N_24625,N_24565);
and U24911 (N_24911,N_24616,N_24620);
nor U24912 (N_24912,N_24661,N_24634);
xnor U24913 (N_24913,N_24560,N_24632);
or U24914 (N_24914,N_24574,N_24663);
nand U24915 (N_24915,N_24694,N_24700);
or U24916 (N_24916,N_24500,N_24713);
and U24917 (N_24917,N_24573,N_24591);
nor U24918 (N_24918,N_24640,N_24618);
nand U24919 (N_24919,N_24699,N_24521);
nand U24920 (N_24920,N_24580,N_24734);
nand U24921 (N_24921,N_24572,N_24741);
nand U24922 (N_24922,N_24656,N_24605);
nor U24923 (N_24923,N_24599,N_24526);
xnor U24924 (N_24924,N_24619,N_24644);
and U24925 (N_24925,N_24678,N_24645);
nor U24926 (N_24926,N_24572,N_24674);
nor U24927 (N_24927,N_24708,N_24538);
and U24928 (N_24928,N_24688,N_24594);
nor U24929 (N_24929,N_24715,N_24650);
nor U24930 (N_24930,N_24652,N_24540);
or U24931 (N_24931,N_24575,N_24502);
nand U24932 (N_24932,N_24688,N_24716);
and U24933 (N_24933,N_24745,N_24698);
xnor U24934 (N_24934,N_24550,N_24553);
nor U24935 (N_24935,N_24630,N_24600);
nand U24936 (N_24936,N_24748,N_24588);
or U24937 (N_24937,N_24724,N_24567);
nand U24938 (N_24938,N_24711,N_24612);
or U24939 (N_24939,N_24696,N_24741);
and U24940 (N_24940,N_24502,N_24525);
nand U24941 (N_24941,N_24648,N_24700);
and U24942 (N_24942,N_24711,N_24707);
and U24943 (N_24943,N_24683,N_24543);
and U24944 (N_24944,N_24724,N_24526);
or U24945 (N_24945,N_24685,N_24529);
nand U24946 (N_24946,N_24727,N_24569);
xor U24947 (N_24947,N_24665,N_24599);
nor U24948 (N_24948,N_24632,N_24625);
nor U24949 (N_24949,N_24664,N_24570);
nand U24950 (N_24950,N_24668,N_24699);
or U24951 (N_24951,N_24574,N_24520);
and U24952 (N_24952,N_24722,N_24581);
or U24953 (N_24953,N_24573,N_24715);
xor U24954 (N_24954,N_24586,N_24605);
or U24955 (N_24955,N_24667,N_24645);
and U24956 (N_24956,N_24521,N_24700);
or U24957 (N_24957,N_24668,N_24683);
nand U24958 (N_24958,N_24548,N_24574);
nand U24959 (N_24959,N_24558,N_24698);
xor U24960 (N_24960,N_24553,N_24704);
or U24961 (N_24961,N_24674,N_24532);
nand U24962 (N_24962,N_24687,N_24544);
or U24963 (N_24963,N_24586,N_24669);
or U24964 (N_24964,N_24609,N_24596);
or U24965 (N_24965,N_24644,N_24566);
nor U24966 (N_24966,N_24738,N_24668);
or U24967 (N_24967,N_24518,N_24738);
nand U24968 (N_24968,N_24565,N_24746);
nor U24969 (N_24969,N_24626,N_24605);
xnor U24970 (N_24970,N_24635,N_24584);
and U24971 (N_24971,N_24573,N_24719);
and U24972 (N_24972,N_24584,N_24669);
and U24973 (N_24973,N_24528,N_24663);
nor U24974 (N_24974,N_24579,N_24501);
or U24975 (N_24975,N_24513,N_24601);
and U24976 (N_24976,N_24704,N_24688);
and U24977 (N_24977,N_24508,N_24500);
nand U24978 (N_24978,N_24622,N_24554);
nand U24979 (N_24979,N_24748,N_24574);
or U24980 (N_24980,N_24635,N_24505);
and U24981 (N_24981,N_24558,N_24749);
xnor U24982 (N_24982,N_24714,N_24749);
xnor U24983 (N_24983,N_24732,N_24706);
nor U24984 (N_24984,N_24719,N_24636);
nor U24985 (N_24985,N_24528,N_24629);
and U24986 (N_24986,N_24568,N_24573);
nand U24987 (N_24987,N_24616,N_24670);
or U24988 (N_24988,N_24651,N_24696);
or U24989 (N_24989,N_24508,N_24599);
and U24990 (N_24990,N_24533,N_24687);
and U24991 (N_24991,N_24722,N_24679);
nor U24992 (N_24992,N_24666,N_24554);
and U24993 (N_24993,N_24736,N_24567);
nand U24994 (N_24994,N_24749,N_24634);
xor U24995 (N_24995,N_24515,N_24637);
and U24996 (N_24996,N_24671,N_24719);
and U24997 (N_24997,N_24665,N_24715);
or U24998 (N_24998,N_24522,N_24690);
nor U24999 (N_24999,N_24591,N_24618);
or UO_0 (O_0,N_24961,N_24875);
xor UO_1 (O_1,N_24886,N_24768);
and UO_2 (O_2,N_24869,N_24891);
nand UO_3 (O_3,N_24926,N_24933);
and UO_4 (O_4,N_24750,N_24937);
nor UO_5 (O_5,N_24919,N_24994);
xnor UO_6 (O_6,N_24997,N_24798);
nor UO_7 (O_7,N_24806,N_24953);
and UO_8 (O_8,N_24861,N_24955);
and UO_9 (O_9,N_24868,N_24895);
and UO_10 (O_10,N_24931,N_24837);
xnor UO_11 (O_11,N_24782,N_24870);
and UO_12 (O_12,N_24901,N_24962);
nand UO_13 (O_13,N_24871,N_24847);
xor UO_14 (O_14,N_24756,N_24893);
nand UO_15 (O_15,N_24945,N_24940);
nor UO_16 (O_16,N_24779,N_24909);
or UO_17 (O_17,N_24758,N_24885);
or UO_18 (O_18,N_24966,N_24946);
nand UO_19 (O_19,N_24924,N_24925);
and UO_20 (O_20,N_24797,N_24920);
nor UO_21 (O_21,N_24970,N_24786);
and UO_22 (O_22,N_24984,N_24843);
xor UO_23 (O_23,N_24880,N_24856);
and UO_24 (O_24,N_24833,N_24838);
nand UO_25 (O_25,N_24910,N_24899);
nor UO_26 (O_26,N_24840,N_24948);
xnor UO_27 (O_27,N_24975,N_24776);
nor UO_28 (O_28,N_24904,N_24855);
or UO_29 (O_29,N_24845,N_24809);
or UO_30 (O_30,N_24803,N_24889);
nand UO_31 (O_31,N_24853,N_24978);
xnor UO_32 (O_32,N_24791,N_24848);
or UO_33 (O_33,N_24993,N_24888);
and UO_34 (O_34,N_24942,N_24813);
or UO_35 (O_35,N_24958,N_24752);
nand UO_36 (O_36,N_24763,N_24824);
and UO_37 (O_37,N_24842,N_24898);
nand UO_38 (O_38,N_24804,N_24916);
nand UO_39 (O_39,N_24979,N_24815);
xnor UO_40 (O_40,N_24836,N_24960);
nand UO_41 (O_41,N_24774,N_24821);
or UO_42 (O_42,N_24773,N_24943);
xor UO_43 (O_43,N_24911,N_24989);
and UO_44 (O_44,N_24969,N_24915);
nor UO_45 (O_45,N_24762,N_24789);
or UO_46 (O_46,N_24985,N_24936);
or UO_47 (O_47,N_24929,N_24822);
or UO_48 (O_48,N_24995,N_24968);
and UO_49 (O_49,N_24864,N_24878);
nand UO_50 (O_50,N_24785,N_24783);
nor UO_51 (O_51,N_24757,N_24980);
nor UO_52 (O_52,N_24883,N_24765);
nand UO_53 (O_53,N_24780,N_24932);
or UO_54 (O_54,N_24902,N_24884);
and UO_55 (O_55,N_24811,N_24754);
xor UO_56 (O_56,N_24907,N_24852);
nand UO_57 (O_57,N_24810,N_24977);
nor UO_58 (O_58,N_24830,N_24944);
nand UO_59 (O_59,N_24956,N_24874);
nand UO_60 (O_60,N_24796,N_24867);
and UO_61 (O_61,N_24918,N_24828);
nor UO_62 (O_62,N_24787,N_24777);
and UO_63 (O_63,N_24831,N_24832);
nor UO_64 (O_64,N_24794,N_24860);
nor UO_65 (O_65,N_24849,N_24835);
xor UO_66 (O_66,N_24972,N_24974);
or UO_67 (O_67,N_24921,N_24983);
nor UO_68 (O_68,N_24927,N_24971);
nand UO_69 (O_69,N_24854,N_24872);
nand UO_70 (O_70,N_24807,N_24817);
and UO_71 (O_71,N_24959,N_24954);
or UO_72 (O_72,N_24819,N_24957);
xor UO_73 (O_73,N_24890,N_24930);
nand UO_74 (O_74,N_24952,N_24894);
and UO_75 (O_75,N_24814,N_24963);
xnor UO_76 (O_76,N_24912,N_24887);
nor UO_77 (O_77,N_24771,N_24986);
nand UO_78 (O_78,N_24976,N_24761);
and UO_79 (O_79,N_24947,N_24795);
xor UO_80 (O_80,N_24876,N_24766);
xor UO_81 (O_81,N_24850,N_24873);
or UO_82 (O_82,N_24862,N_24964);
nor UO_83 (O_83,N_24981,N_24865);
nor UO_84 (O_84,N_24764,N_24775);
nand UO_85 (O_85,N_24825,N_24839);
nand UO_86 (O_86,N_24950,N_24951);
xor UO_87 (O_87,N_24914,N_24917);
nand UO_88 (O_88,N_24903,N_24882);
xor UO_89 (O_89,N_24772,N_24896);
nand UO_90 (O_90,N_24973,N_24879);
and UO_91 (O_91,N_24799,N_24788);
and UO_92 (O_92,N_24857,N_24858);
nor UO_93 (O_93,N_24991,N_24769);
nand UO_94 (O_94,N_24866,N_24965);
xnor UO_95 (O_95,N_24990,N_24941);
and UO_96 (O_96,N_24826,N_24881);
xor UO_97 (O_97,N_24928,N_24851);
or UO_98 (O_98,N_24751,N_24923);
and UO_99 (O_99,N_24987,N_24805);
or UO_100 (O_100,N_24897,N_24988);
xor UO_101 (O_101,N_24820,N_24992);
and UO_102 (O_102,N_24800,N_24801);
and UO_103 (O_103,N_24998,N_24753);
or UO_104 (O_104,N_24900,N_24759);
nand UO_105 (O_105,N_24938,N_24934);
and UO_106 (O_106,N_24834,N_24808);
and UO_107 (O_107,N_24859,N_24760);
xnor UO_108 (O_108,N_24846,N_24767);
or UO_109 (O_109,N_24841,N_24863);
nor UO_110 (O_110,N_24877,N_24829);
xor UO_111 (O_111,N_24982,N_24935);
and UO_112 (O_112,N_24906,N_24793);
nor UO_113 (O_113,N_24778,N_24770);
nor UO_114 (O_114,N_24792,N_24781);
xnor UO_115 (O_115,N_24844,N_24967);
and UO_116 (O_116,N_24949,N_24818);
and UO_117 (O_117,N_24755,N_24939);
and UO_118 (O_118,N_24999,N_24790);
or UO_119 (O_119,N_24827,N_24996);
and UO_120 (O_120,N_24892,N_24812);
or UO_121 (O_121,N_24913,N_24784);
nor UO_122 (O_122,N_24816,N_24823);
xnor UO_123 (O_123,N_24908,N_24905);
nor UO_124 (O_124,N_24922,N_24802);
xnor UO_125 (O_125,N_24758,N_24823);
or UO_126 (O_126,N_24812,N_24899);
or UO_127 (O_127,N_24902,N_24881);
xnor UO_128 (O_128,N_24891,N_24759);
and UO_129 (O_129,N_24840,N_24936);
and UO_130 (O_130,N_24930,N_24962);
nor UO_131 (O_131,N_24826,N_24783);
xor UO_132 (O_132,N_24876,N_24967);
or UO_133 (O_133,N_24866,N_24751);
and UO_134 (O_134,N_24996,N_24971);
and UO_135 (O_135,N_24820,N_24936);
or UO_136 (O_136,N_24848,N_24944);
nand UO_137 (O_137,N_24791,N_24892);
xnor UO_138 (O_138,N_24951,N_24895);
xor UO_139 (O_139,N_24805,N_24884);
nand UO_140 (O_140,N_24802,N_24844);
nor UO_141 (O_141,N_24945,N_24886);
nand UO_142 (O_142,N_24886,N_24872);
or UO_143 (O_143,N_24765,N_24879);
nor UO_144 (O_144,N_24816,N_24800);
or UO_145 (O_145,N_24921,N_24968);
or UO_146 (O_146,N_24898,N_24869);
nand UO_147 (O_147,N_24859,N_24834);
nand UO_148 (O_148,N_24770,N_24853);
nor UO_149 (O_149,N_24818,N_24861);
xor UO_150 (O_150,N_24896,N_24826);
xor UO_151 (O_151,N_24890,N_24797);
nor UO_152 (O_152,N_24993,N_24828);
nand UO_153 (O_153,N_24916,N_24852);
and UO_154 (O_154,N_24948,N_24816);
nor UO_155 (O_155,N_24858,N_24750);
and UO_156 (O_156,N_24878,N_24939);
nor UO_157 (O_157,N_24934,N_24889);
nor UO_158 (O_158,N_24843,N_24854);
xnor UO_159 (O_159,N_24794,N_24770);
nand UO_160 (O_160,N_24905,N_24782);
or UO_161 (O_161,N_24855,N_24829);
xnor UO_162 (O_162,N_24943,N_24953);
or UO_163 (O_163,N_24755,N_24968);
or UO_164 (O_164,N_24803,N_24940);
nor UO_165 (O_165,N_24807,N_24838);
nor UO_166 (O_166,N_24832,N_24761);
xor UO_167 (O_167,N_24803,N_24863);
and UO_168 (O_168,N_24920,N_24940);
nand UO_169 (O_169,N_24914,N_24910);
xor UO_170 (O_170,N_24939,N_24872);
xor UO_171 (O_171,N_24966,N_24810);
or UO_172 (O_172,N_24848,N_24920);
and UO_173 (O_173,N_24871,N_24794);
nand UO_174 (O_174,N_24777,N_24866);
nor UO_175 (O_175,N_24800,N_24932);
nand UO_176 (O_176,N_24917,N_24962);
and UO_177 (O_177,N_24979,N_24886);
xnor UO_178 (O_178,N_24820,N_24796);
or UO_179 (O_179,N_24966,N_24993);
xor UO_180 (O_180,N_24913,N_24810);
and UO_181 (O_181,N_24980,N_24759);
or UO_182 (O_182,N_24775,N_24839);
nor UO_183 (O_183,N_24986,N_24962);
and UO_184 (O_184,N_24821,N_24777);
xnor UO_185 (O_185,N_24854,N_24947);
nand UO_186 (O_186,N_24904,N_24949);
nor UO_187 (O_187,N_24925,N_24892);
and UO_188 (O_188,N_24910,N_24953);
and UO_189 (O_189,N_24824,N_24857);
xor UO_190 (O_190,N_24975,N_24873);
nor UO_191 (O_191,N_24923,N_24816);
nand UO_192 (O_192,N_24928,N_24766);
xnor UO_193 (O_193,N_24960,N_24773);
and UO_194 (O_194,N_24947,N_24952);
or UO_195 (O_195,N_24891,N_24806);
nand UO_196 (O_196,N_24962,N_24826);
or UO_197 (O_197,N_24970,N_24802);
and UO_198 (O_198,N_24989,N_24926);
and UO_199 (O_199,N_24867,N_24834);
xor UO_200 (O_200,N_24826,N_24973);
and UO_201 (O_201,N_24970,N_24939);
nor UO_202 (O_202,N_24848,N_24830);
xor UO_203 (O_203,N_24989,N_24859);
and UO_204 (O_204,N_24905,N_24785);
nor UO_205 (O_205,N_24928,N_24787);
and UO_206 (O_206,N_24759,N_24991);
and UO_207 (O_207,N_24781,N_24772);
xnor UO_208 (O_208,N_24921,N_24885);
xnor UO_209 (O_209,N_24835,N_24775);
nor UO_210 (O_210,N_24945,N_24795);
nor UO_211 (O_211,N_24990,N_24931);
xor UO_212 (O_212,N_24963,N_24797);
or UO_213 (O_213,N_24755,N_24853);
nor UO_214 (O_214,N_24770,N_24776);
nor UO_215 (O_215,N_24905,N_24765);
xnor UO_216 (O_216,N_24998,N_24821);
or UO_217 (O_217,N_24958,N_24780);
xor UO_218 (O_218,N_24951,N_24856);
or UO_219 (O_219,N_24967,N_24768);
nor UO_220 (O_220,N_24955,N_24959);
and UO_221 (O_221,N_24821,N_24950);
or UO_222 (O_222,N_24947,N_24891);
or UO_223 (O_223,N_24780,N_24793);
and UO_224 (O_224,N_24751,N_24950);
xnor UO_225 (O_225,N_24772,N_24756);
nand UO_226 (O_226,N_24826,N_24909);
and UO_227 (O_227,N_24767,N_24782);
and UO_228 (O_228,N_24921,N_24966);
nand UO_229 (O_229,N_24805,N_24844);
or UO_230 (O_230,N_24876,N_24937);
and UO_231 (O_231,N_24780,N_24837);
nor UO_232 (O_232,N_24889,N_24918);
nor UO_233 (O_233,N_24961,N_24976);
nand UO_234 (O_234,N_24931,N_24796);
nand UO_235 (O_235,N_24845,N_24836);
xor UO_236 (O_236,N_24850,N_24773);
or UO_237 (O_237,N_24957,N_24884);
or UO_238 (O_238,N_24751,N_24806);
nand UO_239 (O_239,N_24929,N_24829);
xor UO_240 (O_240,N_24911,N_24897);
xnor UO_241 (O_241,N_24752,N_24813);
xor UO_242 (O_242,N_24920,N_24822);
nand UO_243 (O_243,N_24817,N_24798);
or UO_244 (O_244,N_24992,N_24915);
nand UO_245 (O_245,N_24779,N_24987);
xor UO_246 (O_246,N_24910,N_24966);
or UO_247 (O_247,N_24943,N_24930);
and UO_248 (O_248,N_24987,N_24975);
xnor UO_249 (O_249,N_24989,N_24930);
nand UO_250 (O_250,N_24843,N_24807);
xor UO_251 (O_251,N_24842,N_24992);
xor UO_252 (O_252,N_24970,N_24858);
and UO_253 (O_253,N_24812,N_24863);
and UO_254 (O_254,N_24812,N_24866);
nor UO_255 (O_255,N_24929,N_24767);
nand UO_256 (O_256,N_24822,N_24983);
and UO_257 (O_257,N_24801,N_24768);
or UO_258 (O_258,N_24922,N_24755);
and UO_259 (O_259,N_24909,N_24889);
or UO_260 (O_260,N_24923,N_24995);
xor UO_261 (O_261,N_24804,N_24901);
and UO_262 (O_262,N_24956,N_24997);
nand UO_263 (O_263,N_24993,N_24813);
and UO_264 (O_264,N_24790,N_24868);
and UO_265 (O_265,N_24854,N_24814);
xnor UO_266 (O_266,N_24784,N_24887);
and UO_267 (O_267,N_24844,N_24989);
and UO_268 (O_268,N_24776,N_24981);
nor UO_269 (O_269,N_24994,N_24892);
and UO_270 (O_270,N_24845,N_24883);
nor UO_271 (O_271,N_24775,N_24921);
xor UO_272 (O_272,N_24910,N_24809);
xnor UO_273 (O_273,N_24856,N_24884);
and UO_274 (O_274,N_24876,N_24931);
xnor UO_275 (O_275,N_24773,N_24825);
nor UO_276 (O_276,N_24905,N_24973);
and UO_277 (O_277,N_24951,N_24917);
or UO_278 (O_278,N_24972,N_24811);
xor UO_279 (O_279,N_24925,N_24820);
xor UO_280 (O_280,N_24761,N_24783);
and UO_281 (O_281,N_24995,N_24799);
or UO_282 (O_282,N_24854,N_24896);
nand UO_283 (O_283,N_24883,N_24840);
and UO_284 (O_284,N_24952,N_24954);
nor UO_285 (O_285,N_24823,N_24933);
xnor UO_286 (O_286,N_24830,N_24828);
and UO_287 (O_287,N_24931,N_24830);
or UO_288 (O_288,N_24902,N_24911);
and UO_289 (O_289,N_24937,N_24863);
and UO_290 (O_290,N_24885,N_24965);
nor UO_291 (O_291,N_24917,N_24767);
nand UO_292 (O_292,N_24786,N_24778);
nor UO_293 (O_293,N_24910,N_24925);
or UO_294 (O_294,N_24824,N_24978);
nor UO_295 (O_295,N_24932,N_24848);
and UO_296 (O_296,N_24782,N_24964);
or UO_297 (O_297,N_24845,N_24808);
nand UO_298 (O_298,N_24952,N_24845);
nor UO_299 (O_299,N_24891,N_24926);
nand UO_300 (O_300,N_24836,N_24801);
nand UO_301 (O_301,N_24905,N_24899);
nor UO_302 (O_302,N_24958,N_24761);
and UO_303 (O_303,N_24791,N_24766);
xnor UO_304 (O_304,N_24765,N_24846);
and UO_305 (O_305,N_24873,N_24891);
or UO_306 (O_306,N_24888,N_24906);
nor UO_307 (O_307,N_24803,N_24781);
and UO_308 (O_308,N_24853,N_24868);
or UO_309 (O_309,N_24845,N_24840);
nor UO_310 (O_310,N_24786,N_24787);
nand UO_311 (O_311,N_24815,N_24952);
xor UO_312 (O_312,N_24857,N_24937);
or UO_313 (O_313,N_24795,N_24904);
xnor UO_314 (O_314,N_24957,N_24851);
nor UO_315 (O_315,N_24913,N_24896);
nand UO_316 (O_316,N_24762,N_24872);
nor UO_317 (O_317,N_24867,N_24843);
xor UO_318 (O_318,N_24987,N_24888);
nor UO_319 (O_319,N_24883,N_24802);
nand UO_320 (O_320,N_24987,N_24877);
or UO_321 (O_321,N_24813,N_24933);
xnor UO_322 (O_322,N_24800,N_24770);
or UO_323 (O_323,N_24824,N_24781);
nor UO_324 (O_324,N_24979,N_24834);
nand UO_325 (O_325,N_24906,N_24982);
nor UO_326 (O_326,N_24975,N_24828);
xnor UO_327 (O_327,N_24857,N_24865);
nor UO_328 (O_328,N_24968,N_24809);
nand UO_329 (O_329,N_24999,N_24955);
xor UO_330 (O_330,N_24836,N_24934);
xor UO_331 (O_331,N_24968,N_24906);
nor UO_332 (O_332,N_24855,N_24808);
xor UO_333 (O_333,N_24800,N_24997);
nor UO_334 (O_334,N_24878,N_24813);
nand UO_335 (O_335,N_24917,N_24758);
nand UO_336 (O_336,N_24865,N_24805);
xor UO_337 (O_337,N_24841,N_24781);
xor UO_338 (O_338,N_24949,N_24777);
or UO_339 (O_339,N_24935,N_24821);
nand UO_340 (O_340,N_24889,N_24845);
nor UO_341 (O_341,N_24840,N_24968);
nor UO_342 (O_342,N_24807,N_24874);
or UO_343 (O_343,N_24836,N_24850);
xor UO_344 (O_344,N_24762,N_24962);
and UO_345 (O_345,N_24926,N_24765);
or UO_346 (O_346,N_24871,N_24756);
nand UO_347 (O_347,N_24805,N_24836);
nand UO_348 (O_348,N_24752,N_24822);
or UO_349 (O_349,N_24874,N_24899);
xnor UO_350 (O_350,N_24772,N_24811);
and UO_351 (O_351,N_24832,N_24849);
xnor UO_352 (O_352,N_24816,N_24811);
or UO_353 (O_353,N_24932,N_24818);
nor UO_354 (O_354,N_24981,N_24781);
or UO_355 (O_355,N_24867,N_24872);
xor UO_356 (O_356,N_24827,N_24997);
and UO_357 (O_357,N_24894,N_24900);
nor UO_358 (O_358,N_24812,N_24805);
nor UO_359 (O_359,N_24912,N_24961);
or UO_360 (O_360,N_24966,N_24973);
nor UO_361 (O_361,N_24984,N_24763);
nor UO_362 (O_362,N_24755,N_24770);
and UO_363 (O_363,N_24977,N_24990);
and UO_364 (O_364,N_24850,N_24871);
nor UO_365 (O_365,N_24801,N_24901);
or UO_366 (O_366,N_24990,N_24993);
and UO_367 (O_367,N_24939,N_24772);
nor UO_368 (O_368,N_24999,N_24859);
nand UO_369 (O_369,N_24909,N_24812);
nor UO_370 (O_370,N_24900,N_24899);
or UO_371 (O_371,N_24803,N_24947);
and UO_372 (O_372,N_24778,N_24897);
nor UO_373 (O_373,N_24996,N_24933);
or UO_374 (O_374,N_24969,N_24794);
nor UO_375 (O_375,N_24911,N_24769);
nand UO_376 (O_376,N_24752,N_24815);
or UO_377 (O_377,N_24999,N_24755);
and UO_378 (O_378,N_24819,N_24899);
xor UO_379 (O_379,N_24946,N_24846);
nand UO_380 (O_380,N_24939,N_24765);
nor UO_381 (O_381,N_24924,N_24960);
and UO_382 (O_382,N_24750,N_24992);
nand UO_383 (O_383,N_24859,N_24826);
nor UO_384 (O_384,N_24905,N_24836);
or UO_385 (O_385,N_24988,N_24946);
and UO_386 (O_386,N_24870,N_24983);
or UO_387 (O_387,N_24834,N_24909);
nor UO_388 (O_388,N_24780,N_24993);
nand UO_389 (O_389,N_24999,N_24783);
and UO_390 (O_390,N_24984,N_24977);
xnor UO_391 (O_391,N_24757,N_24894);
nor UO_392 (O_392,N_24775,N_24993);
nor UO_393 (O_393,N_24919,N_24795);
or UO_394 (O_394,N_24813,N_24907);
xnor UO_395 (O_395,N_24768,N_24988);
and UO_396 (O_396,N_24927,N_24972);
xnor UO_397 (O_397,N_24968,N_24940);
nor UO_398 (O_398,N_24783,N_24777);
nor UO_399 (O_399,N_24870,N_24963);
nand UO_400 (O_400,N_24901,N_24913);
nand UO_401 (O_401,N_24751,N_24773);
xnor UO_402 (O_402,N_24965,N_24971);
nor UO_403 (O_403,N_24751,N_24871);
nand UO_404 (O_404,N_24821,N_24948);
xnor UO_405 (O_405,N_24974,N_24805);
or UO_406 (O_406,N_24851,N_24978);
nand UO_407 (O_407,N_24820,N_24918);
and UO_408 (O_408,N_24865,N_24838);
nor UO_409 (O_409,N_24984,N_24870);
and UO_410 (O_410,N_24787,N_24766);
xnor UO_411 (O_411,N_24955,N_24931);
or UO_412 (O_412,N_24950,N_24958);
xor UO_413 (O_413,N_24782,N_24779);
and UO_414 (O_414,N_24892,N_24887);
nor UO_415 (O_415,N_24803,N_24951);
and UO_416 (O_416,N_24799,N_24836);
nor UO_417 (O_417,N_24992,N_24891);
nand UO_418 (O_418,N_24807,N_24998);
xnor UO_419 (O_419,N_24998,N_24872);
and UO_420 (O_420,N_24954,N_24976);
xor UO_421 (O_421,N_24932,N_24792);
nor UO_422 (O_422,N_24970,N_24846);
or UO_423 (O_423,N_24894,N_24826);
or UO_424 (O_424,N_24753,N_24910);
xnor UO_425 (O_425,N_24754,N_24900);
or UO_426 (O_426,N_24757,N_24860);
or UO_427 (O_427,N_24821,N_24884);
xor UO_428 (O_428,N_24996,N_24912);
nand UO_429 (O_429,N_24951,N_24942);
or UO_430 (O_430,N_24916,N_24873);
nand UO_431 (O_431,N_24907,N_24893);
nand UO_432 (O_432,N_24911,N_24788);
xor UO_433 (O_433,N_24997,N_24869);
and UO_434 (O_434,N_24838,N_24858);
and UO_435 (O_435,N_24760,N_24852);
or UO_436 (O_436,N_24990,N_24955);
xnor UO_437 (O_437,N_24791,N_24862);
nand UO_438 (O_438,N_24892,N_24854);
or UO_439 (O_439,N_24779,N_24953);
nor UO_440 (O_440,N_24825,N_24774);
nor UO_441 (O_441,N_24794,N_24820);
or UO_442 (O_442,N_24946,N_24831);
xor UO_443 (O_443,N_24823,N_24984);
nor UO_444 (O_444,N_24906,N_24779);
and UO_445 (O_445,N_24762,N_24782);
xor UO_446 (O_446,N_24773,N_24783);
or UO_447 (O_447,N_24888,N_24985);
nand UO_448 (O_448,N_24885,N_24828);
or UO_449 (O_449,N_24831,N_24822);
or UO_450 (O_450,N_24941,N_24853);
nand UO_451 (O_451,N_24933,N_24851);
xor UO_452 (O_452,N_24809,N_24917);
nand UO_453 (O_453,N_24888,N_24996);
and UO_454 (O_454,N_24778,N_24854);
nand UO_455 (O_455,N_24796,N_24769);
nand UO_456 (O_456,N_24782,N_24859);
or UO_457 (O_457,N_24817,N_24905);
nor UO_458 (O_458,N_24807,N_24884);
nand UO_459 (O_459,N_24798,N_24964);
and UO_460 (O_460,N_24921,N_24816);
nor UO_461 (O_461,N_24920,N_24956);
and UO_462 (O_462,N_24852,N_24904);
and UO_463 (O_463,N_24808,N_24910);
nor UO_464 (O_464,N_24880,N_24831);
or UO_465 (O_465,N_24907,N_24971);
nand UO_466 (O_466,N_24907,N_24987);
or UO_467 (O_467,N_24847,N_24979);
or UO_468 (O_468,N_24886,N_24894);
or UO_469 (O_469,N_24895,N_24865);
nor UO_470 (O_470,N_24834,N_24886);
and UO_471 (O_471,N_24855,N_24867);
or UO_472 (O_472,N_24878,N_24861);
and UO_473 (O_473,N_24830,N_24762);
nor UO_474 (O_474,N_24768,N_24804);
and UO_475 (O_475,N_24898,N_24915);
nand UO_476 (O_476,N_24803,N_24868);
and UO_477 (O_477,N_24910,N_24759);
nand UO_478 (O_478,N_24764,N_24798);
xnor UO_479 (O_479,N_24807,N_24961);
xor UO_480 (O_480,N_24789,N_24836);
or UO_481 (O_481,N_24751,N_24859);
and UO_482 (O_482,N_24926,N_24966);
xnor UO_483 (O_483,N_24947,N_24750);
xnor UO_484 (O_484,N_24947,N_24876);
xnor UO_485 (O_485,N_24983,N_24836);
xor UO_486 (O_486,N_24972,N_24884);
or UO_487 (O_487,N_24963,N_24839);
and UO_488 (O_488,N_24903,N_24984);
nand UO_489 (O_489,N_24949,N_24835);
and UO_490 (O_490,N_24762,N_24796);
or UO_491 (O_491,N_24853,N_24969);
nor UO_492 (O_492,N_24863,N_24982);
xor UO_493 (O_493,N_24808,N_24778);
xnor UO_494 (O_494,N_24978,N_24910);
nand UO_495 (O_495,N_24980,N_24941);
and UO_496 (O_496,N_24835,N_24756);
and UO_497 (O_497,N_24768,N_24906);
nand UO_498 (O_498,N_24803,N_24857);
or UO_499 (O_499,N_24992,N_24875);
xor UO_500 (O_500,N_24755,N_24769);
nor UO_501 (O_501,N_24962,N_24919);
xor UO_502 (O_502,N_24961,N_24880);
or UO_503 (O_503,N_24966,N_24798);
nand UO_504 (O_504,N_24878,N_24841);
or UO_505 (O_505,N_24881,N_24851);
nand UO_506 (O_506,N_24818,N_24881);
nand UO_507 (O_507,N_24872,N_24801);
nand UO_508 (O_508,N_24981,N_24916);
or UO_509 (O_509,N_24974,N_24960);
and UO_510 (O_510,N_24902,N_24870);
xnor UO_511 (O_511,N_24816,N_24848);
or UO_512 (O_512,N_24846,N_24914);
xnor UO_513 (O_513,N_24922,N_24862);
nor UO_514 (O_514,N_24970,N_24945);
xor UO_515 (O_515,N_24782,N_24823);
or UO_516 (O_516,N_24852,N_24812);
or UO_517 (O_517,N_24975,N_24992);
or UO_518 (O_518,N_24833,N_24901);
or UO_519 (O_519,N_24833,N_24770);
and UO_520 (O_520,N_24939,N_24810);
and UO_521 (O_521,N_24838,N_24864);
nor UO_522 (O_522,N_24887,N_24803);
nand UO_523 (O_523,N_24885,N_24878);
and UO_524 (O_524,N_24882,N_24890);
and UO_525 (O_525,N_24987,N_24827);
nor UO_526 (O_526,N_24814,N_24975);
xor UO_527 (O_527,N_24761,N_24883);
xor UO_528 (O_528,N_24953,N_24977);
and UO_529 (O_529,N_24929,N_24864);
and UO_530 (O_530,N_24957,N_24972);
or UO_531 (O_531,N_24847,N_24905);
and UO_532 (O_532,N_24767,N_24908);
xor UO_533 (O_533,N_24949,N_24805);
nand UO_534 (O_534,N_24958,N_24976);
nor UO_535 (O_535,N_24985,N_24794);
or UO_536 (O_536,N_24885,N_24879);
nor UO_537 (O_537,N_24779,N_24955);
and UO_538 (O_538,N_24841,N_24816);
nor UO_539 (O_539,N_24985,N_24991);
xor UO_540 (O_540,N_24995,N_24800);
or UO_541 (O_541,N_24768,N_24798);
nor UO_542 (O_542,N_24914,N_24918);
or UO_543 (O_543,N_24837,N_24978);
and UO_544 (O_544,N_24752,N_24976);
nor UO_545 (O_545,N_24967,N_24860);
nor UO_546 (O_546,N_24917,N_24864);
nand UO_547 (O_547,N_24910,N_24845);
and UO_548 (O_548,N_24884,N_24825);
nor UO_549 (O_549,N_24955,N_24780);
nor UO_550 (O_550,N_24866,N_24937);
nand UO_551 (O_551,N_24774,N_24811);
nor UO_552 (O_552,N_24989,N_24985);
nand UO_553 (O_553,N_24917,N_24755);
xor UO_554 (O_554,N_24839,N_24992);
and UO_555 (O_555,N_24797,N_24817);
nand UO_556 (O_556,N_24869,N_24811);
or UO_557 (O_557,N_24988,N_24823);
nand UO_558 (O_558,N_24939,N_24927);
nor UO_559 (O_559,N_24893,N_24883);
and UO_560 (O_560,N_24841,N_24902);
or UO_561 (O_561,N_24770,N_24837);
nor UO_562 (O_562,N_24760,N_24980);
nand UO_563 (O_563,N_24940,N_24933);
xnor UO_564 (O_564,N_24815,N_24826);
and UO_565 (O_565,N_24860,N_24930);
and UO_566 (O_566,N_24880,N_24784);
nor UO_567 (O_567,N_24785,N_24800);
nor UO_568 (O_568,N_24784,N_24957);
xor UO_569 (O_569,N_24963,N_24951);
xnor UO_570 (O_570,N_24905,N_24934);
xor UO_571 (O_571,N_24859,N_24993);
nor UO_572 (O_572,N_24765,N_24855);
and UO_573 (O_573,N_24778,N_24872);
and UO_574 (O_574,N_24878,N_24905);
nand UO_575 (O_575,N_24792,N_24988);
xnor UO_576 (O_576,N_24915,N_24820);
xor UO_577 (O_577,N_24874,N_24849);
or UO_578 (O_578,N_24818,N_24987);
nand UO_579 (O_579,N_24874,N_24770);
nor UO_580 (O_580,N_24869,N_24767);
nor UO_581 (O_581,N_24954,N_24864);
xor UO_582 (O_582,N_24972,N_24877);
or UO_583 (O_583,N_24993,N_24820);
and UO_584 (O_584,N_24775,N_24904);
and UO_585 (O_585,N_24879,N_24842);
xnor UO_586 (O_586,N_24759,N_24777);
and UO_587 (O_587,N_24888,N_24882);
and UO_588 (O_588,N_24993,N_24972);
nor UO_589 (O_589,N_24889,N_24990);
xor UO_590 (O_590,N_24764,N_24950);
nor UO_591 (O_591,N_24899,N_24766);
xnor UO_592 (O_592,N_24786,N_24935);
xnor UO_593 (O_593,N_24908,N_24815);
xnor UO_594 (O_594,N_24992,N_24753);
xnor UO_595 (O_595,N_24964,N_24787);
xor UO_596 (O_596,N_24858,N_24854);
nor UO_597 (O_597,N_24803,N_24829);
nand UO_598 (O_598,N_24872,N_24879);
or UO_599 (O_599,N_24820,N_24768);
and UO_600 (O_600,N_24796,N_24865);
nor UO_601 (O_601,N_24828,N_24876);
nand UO_602 (O_602,N_24956,N_24880);
or UO_603 (O_603,N_24879,N_24892);
nand UO_604 (O_604,N_24930,N_24769);
or UO_605 (O_605,N_24830,N_24876);
and UO_606 (O_606,N_24946,N_24906);
nand UO_607 (O_607,N_24842,N_24774);
nor UO_608 (O_608,N_24895,N_24763);
and UO_609 (O_609,N_24906,N_24964);
nor UO_610 (O_610,N_24997,N_24909);
nand UO_611 (O_611,N_24869,N_24937);
nor UO_612 (O_612,N_24928,N_24903);
xnor UO_613 (O_613,N_24820,N_24972);
and UO_614 (O_614,N_24880,N_24753);
and UO_615 (O_615,N_24800,N_24908);
and UO_616 (O_616,N_24988,N_24948);
or UO_617 (O_617,N_24794,N_24795);
and UO_618 (O_618,N_24764,N_24959);
nor UO_619 (O_619,N_24785,N_24851);
nand UO_620 (O_620,N_24942,N_24956);
and UO_621 (O_621,N_24789,N_24808);
nor UO_622 (O_622,N_24975,N_24870);
nor UO_623 (O_623,N_24908,N_24948);
xnor UO_624 (O_624,N_24903,N_24827);
or UO_625 (O_625,N_24824,N_24992);
or UO_626 (O_626,N_24936,N_24873);
or UO_627 (O_627,N_24990,N_24750);
nand UO_628 (O_628,N_24792,N_24859);
and UO_629 (O_629,N_24822,N_24819);
nor UO_630 (O_630,N_24855,N_24892);
nor UO_631 (O_631,N_24766,N_24941);
xor UO_632 (O_632,N_24917,N_24760);
nor UO_633 (O_633,N_24935,N_24983);
or UO_634 (O_634,N_24888,N_24938);
xnor UO_635 (O_635,N_24875,N_24989);
or UO_636 (O_636,N_24785,N_24914);
and UO_637 (O_637,N_24918,N_24788);
and UO_638 (O_638,N_24830,N_24797);
nor UO_639 (O_639,N_24863,N_24839);
nor UO_640 (O_640,N_24869,N_24797);
or UO_641 (O_641,N_24920,N_24991);
xnor UO_642 (O_642,N_24750,N_24932);
nor UO_643 (O_643,N_24881,N_24997);
xnor UO_644 (O_644,N_24835,N_24763);
or UO_645 (O_645,N_24933,N_24966);
and UO_646 (O_646,N_24940,N_24821);
or UO_647 (O_647,N_24874,N_24982);
or UO_648 (O_648,N_24757,N_24938);
xnor UO_649 (O_649,N_24759,N_24808);
nor UO_650 (O_650,N_24852,N_24966);
xnor UO_651 (O_651,N_24852,N_24778);
nor UO_652 (O_652,N_24848,N_24959);
and UO_653 (O_653,N_24975,N_24941);
nor UO_654 (O_654,N_24855,N_24901);
nand UO_655 (O_655,N_24805,N_24975);
nand UO_656 (O_656,N_24761,N_24766);
xnor UO_657 (O_657,N_24974,N_24844);
and UO_658 (O_658,N_24914,N_24964);
nor UO_659 (O_659,N_24927,N_24877);
nor UO_660 (O_660,N_24849,N_24978);
xor UO_661 (O_661,N_24846,N_24838);
nand UO_662 (O_662,N_24974,N_24785);
nand UO_663 (O_663,N_24926,N_24903);
nor UO_664 (O_664,N_24936,N_24980);
nand UO_665 (O_665,N_24880,N_24836);
nor UO_666 (O_666,N_24754,N_24784);
and UO_667 (O_667,N_24950,N_24887);
and UO_668 (O_668,N_24987,N_24810);
nand UO_669 (O_669,N_24856,N_24849);
nor UO_670 (O_670,N_24953,N_24898);
xor UO_671 (O_671,N_24765,N_24955);
nor UO_672 (O_672,N_24784,N_24899);
xor UO_673 (O_673,N_24788,N_24931);
nor UO_674 (O_674,N_24978,N_24895);
or UO_675 (O_675,N_24996,N_24817);
xor UO_676 (O_676,N_24990,N_24754);
nand UO_677 (O_677,N_24776,N_24936);
nor UO_678 (O_678,N_24822,N_24991);
or UO_679 (O_679,N_24774,N_24991);
xnor UO_680 (O_680,N_24987,N_24880);
xor UO_681 (O_681,N_24912,N_24764);
and UO_682 (O_682,N_24980,N_24893);
and UO_683 (O_683,N_24920,N_24770);
xor UO_684 (O_684,N_24924,N_24983);
or UO_685 (O_685,N_24840,N_24945);
or UO_686 (O_686,N_24791,N_24750);
or UO_687 (O_687,N_24906,N_24777);
xnor UO_688 (O_688,N_24960,N_24978);
and UO_689 (O_689,N_24823,N_24989);
and UO_690 (O_690,N_24976,N_24950);
and UO_691 (O_691,N_24762,N_24973);
or UO_692 (O_692,N_24897,N_24819);
xnor UO_693 (O_693,N_24790,N_24919);
nor UO_694 (O_694,N_24878,N_24776);
xnor UO_695 (O_695,N_24793,N_24879);
nor UO_696 (O_696,N_24875,N_24784);
nand UO_697 (O_697,N_24845,N_24829);
xnor UO_698 (O_698,N_24921,N_24828);
and UO_699 (O_699,N_24943,N_24908);
nor UO_700 (O_700,N_24778,N_24954);
nand UO_701 (O_701,N_24761,N_24996);
or UO_702 (O_702,N_24810,N_24927);
nor UO_703 (O_703,N_24902,N_24913);
xor UO_704 (O_704,N_24799,N_24903);
or UO_705 (O_705,N_24853,N_24917);
nor UO_706 (O_706,N_24835,N_24961);
and UO_707 (O_707,N_24795,N_24857);
nand UO_708 (O_708,N_24819,N_24930);
or UO_709 (O_709,N_24811,N_24888);
and UO_710 (O_710,N_24964,N_24874);
xnor UO_711 (O_711,N_24958,N_24963);
or UO_712 (O_712,N_24915,N_24801);
xnor UO_713 (O_713,N_24975,N_24905);
nand UO_714 (O_714,N_24924,N_24840);
nand UO_715 (O_715,N_24999,N_24851);
xnor UO_716 (O_716,N_24804,N_24890);
or UO_717 (O_717,N_24830,N_24900);
or UO_718 (O_718,N_24865,N_24933);
and UO_719 (O_719,N_24961,N_24842);
nor UO_720 (O_720,N_24874,N_24866);
xnor UO_721 (O_721,N_24885,N_24948);
nand UO_722 (O_722,N_24991,N_24873);
xor UO_723 (O_723,N_24791,N_24836);
xnor UO_724 (O_724,N_24870,N_24939);
or UO_725 (O_725,N_24858,N_24784);
xnor UO_726 (O_726,N_24967,N_24915);
or UO_727 (O_727,N_24967,N_24946);
and UO_728 (O_728,N_24891,N_24904);
xor UO_729 (O_729,N_24789,N_24769);
nor UO_730 (O_730,N_24824,N_24817);
and UO_731 (O_731,N_24799,N_24969);
nand UO_732 (O_732,N_24925,N_24848);
xnor UO_733 (O_733,N_24780,N_24987);
nor UO_734 (O_734,N_24880,N_24776);
nor UO_735 (O_735,N_24853,N_24935);
nor UO_736 (O_736,N_24917,N_24990);
xnor UO_737 (O_737,N_24834,N_24902);
nand UO_738 (O_738,N_24931,N_24776);
or UO_739 (O_739,N_24940,N_24910);
and UO_740 (O_740,N_24930,N_24911);
xor UO_741 (O_741,N_24806,N_24846);
and UO_742 (O_742,N_24884,N_24951);
nor UO_743 (O_743,N_24949,N_24900);
and UO_744 (O_744,N_24817,N_24793);
nor UO_745 (O_745,N_24930,N_24754);
nand UO_746 (O_746,N_24875,N_24887);
nand UO_747 (O_747,N_24941,N_24781);
and UO_748 (O_748,N_24845,N_24855);
and UO_749 (O_749,N_24890,N_24896);
and UO_750 (O_750,N_24995,N_24789);
nor UO_751 (O_751,N_24822,N_24933);
or UO_752 (O_752,N_24996,N_24839);
and UO_753 (O_753,N_24928,N_24864);
nand UO_754 (O_754,N_24926,N_24917);
and UO_755 (O_755,N_24978,N_24948);
nand UO_756 (O_756,N_24764,N_24915);
or UO_757 (O_757,N_24893,N_24848);
nand UO_758 (O_758,N_24933,N_24893);
nor UO_759 (O_759,N_24798,N_24854);
xnor UO_760 (O_760,N_24986,N_24872);
nor UO_761 (O_761,N_24843,N_24759);
xor UO_762 (O_762,N_24859,N_24809);
or UO_763 (O_763,N_24769,N_24910);
nand UO_764 (O_764,N_24939,N_24907);
or UO_765 (O_765,N_24828,N_24787);
nor UO_766 (O_766,N_24760,N_24797);
nand UO_767 (O_767,N_24937,N_24858);
or UO_768 (O_768,N_24971,N_24999);
nor UO_769 (O_769,N_24817,N_24787);
and UO_770 (O_770,N_24798,N_24836);
or UO_771 (O_771,N_24953,N_24902);
or UO_772 (O_772,N_24974,N_24765);
nor UO_773 (O_773,N_24828,N_24793);
nor UO_774 (O_774,N_24972,N_24858);
and UO_775 (O_775,N_24819,N_24797);
nand UO_776 (O_776,N_24874,N_24934);
nand UO_777 (O_777,N_24779,N_24833);
nand UO_778 (O_778,N_24794,N_24841);
nor UO_779 (O_779,N_24834,N_24758);
nor UO_780 (O_780,N_24951,N_24935);
xor UO_781 (O_781,N_24894,N_24954);
nand UO_782 (O_782,N_24822,N_24811);
xor UO_783 (O_783,N_24964,N_24984);
nor UO_784 (O_784,N_24920,N_24766);
xor UO_785 (O_785,N_24920,N_24843);
nand UO_786 (O_786,N_24846,N_24909);
or UO_787 (O_787,N_24841,N_24827);
xor UO_788 (O_788,N_24808,N_24763);
or UO_789 (O_789,N_24797,N_24850);
nor UO_790 (O_790,N_24852,N_24837);
xnor UO_791 (O_791,N_24935,N_24799);
or UO_792 (O_792,N_24946,N_24981);
xnor UO_793 (O_793,N_24882,N_24962);
and UO_794 (O_794,N_24945,N_24891);
and UO_795 (O_795,N_24801,N_24896);
and UO_796 (O_796,N_24823,N_24880);
and UO_797 (O_797,N_24915,N_24905);
or UO_798 (O_798,N_24862,N_24769);
nor UO_799 (O_799,N_24763,N_24879);
and UO_800 (O_800,N_24760,N_24788);
xnor UO_801 (O_801,N_24937,N_24903);
nand UO_802 (O_802,N_24885,N_24990);
xnor UO_803 (O_803,N_24935,N_24973);
xor UO_804 (O_804,N_24780,N_24970);
nor UO_805 (O_805,N_24821,N_24836);
nor UO_806 (O_806,N_24849,N_24830);
or UO_807 (O_807,N_24977,N_24839);
and UO_808 (O_808,N_24906,N_24884);
nor UO_809 (O_809,N_24773,N_24780);
xor UO_810 (O_810,N_24896,N_24918);
and UO_811 (O_811,N_24819,N_24882);
xnor UO_812 (O_812,N_24792,N_24801);
nor UO_813 (O_813,N_24816,N_24803);
and UO_814 (O_814,N_24862,N_24849);
nor UO_815 (O_815,N_24891,N_24833);
nand UO_816 (O_816,N_24835,N_24948);
and UO_817 (O_817,N_24835,N_24807);
nand UO_818 (O_818,N_24970,N_24831);
nand UO_819 (O_819,N_24955,N_24946);
or UO_820 (O_820,N_24928,N_24880);
and UO_821 (O_821,N_24994,N_24950);
xor UO_822 (O_822,N_24934,N_24854);
and UO_823 (O_823,N_24916,N_24862);
xnor UO_824 (O_824,N_24985,N_24892);
and UO_825 (O_825,N_24985,N_24823);
xor UO_826 (O_826,N_24753,N_24818);
or UO_827 (O_827,N_24906,N_24822);
and UO_828 (O_828,N_24753,N_24760);
and UO_829 (O_829,N_24862,N_24970);
nor UO_830 (O_830,N_24950,N_24819);
nand UO_831 (O_831,N_24986,N_24896);
nand UO_832 (O_832,N_24975,N_24848);
nor UO_833 (O_833,N_24994,N_24887);
nor UO_834 (O_834,N_24838,N_24755);
nor UO_835 (O_835,N_24905,N_24983);
nand UO_836 (O_836,N_24864,N_24767);
or UO_837 (O_837,N_24975,N_24923);
nor UO_838 (O_838,N_24900,N_24806);
or UO_839 (O_839,N_24893,N_24998);
xnor UO_840 (O_840,N_24789,N_24916);
nand UO_841 (O_841,N_24782,N_24914);
nor UO_842 (O_842,N_24865,N_24826);
xnor UO_843 (O_843,N_24900,N_24911);
nand UO_844 (O_844,N_24811,N_24929);
xnor UO_845 (O_845,N_24938,N_24971);
and UO_846 (O_846,N_24962,N_24972);
nor UO_847 (O_847,N_24897,N_24838);
xor UO_848 (O_848,N_24834,N_24848);
nor UO_849 (O_849,N_24779,N_24971);
nand UO_850 (O_850,N_24775,N_24754);
xor UO_851 (O_851,N_24972,N_24928);
or UO_852 (O_852,N_24915,N_24978);
and UO_853 (O_853,N_24949,N_24966);
and UO_854 (O_854,N_24861,N_24961);
nor UO_855 (O_855,N_24937,N_24968);
or UO_856 (O_856,N_24999,N_24989);
or UO_857 (O_857,N_24827,N_24865);
and UO_858 (O_858,N_24889,N_24818);
or UO_859 (O_859,N_24801,N_24851);
xor UO_860 (O_860,N_24900,N_24943);
or UO_861 (O_861,N_24951,N_24932);
and UO_862 (O_862,N_24925,N_24781);
nand UO_863 (O_863,N_24880,N_24995);
nand UO_864 (O_864,N_24795,N_24899);
nand UO_865 (O_865,N_24839,N_24990);
nor UO_866 (O_866,N_24971,N_24945);
and UO_867 (O_867,N_24885,N_24992);
nor UO_868 (O_868,N_24954,N_24831);
nand UO_869 (O_869,N_24869,N_24775);
or UO_870 (O_870,N_24924,N_24966);
nor UO_871 (O_871,N_24943,N_24989);
nand UO_872 (O_872,N_24797,N_24941);
or UO_873 (O_873,N_24771,N_24875);
nor UO_874 (O_874,N_24926,N_24974);
xor UO_875 (O_875,N_24973,N_24779);
and UO_876 (O_876,N_24966,N_24935);
nand UO_877 (O_877,N_24776,N_24780);
or UO_878 (O_878,N_24863,N_24761);
xor UO_879 (O_879,N_24788,N_24840);
xnor UO_880 (O_880,N_24977,N_24845);
nor UO_881 (O_881,N_24775,N_24759);
xnor UO_882 (O_882,N_24973,N_24956);
and UO_883 (O_883,N_24756,N_24842);
nand UO_884 (O_884,N_24955,N_24800);
nand UO_885 (O_885,N_24933,N_24930);
and UO_886 (O_886,N_24843,N_24754);
and UO_887 (O_887,N_24831,N_24824);
xnor UO_888 (O_888,N_24903,N_24756);
or UO_889 (O_889,N_24857,N_24859);
or UO_890 (O_890,N_24987,N_24847);
nor UO_891 (O_891,N_24857,N_24802);
or UO_892 (O_892,N_24793,N_24845);
nand UO_893 (O_893,N_24977,N_24823);
nand UO_894 (O_894,N_24951,N_24781);
nor UO_895 (O_895,N_24871,N_24778);
and UO_896 (O_896,N_24797,N_24849);
or UO_897 (O_897,N_24817,N_24771);
nor UO_898 (O_898,N_24968,N_24793);
nand UO_899 (O_899,N_24846,N_24963);
nand UO_900 (O_900,N_24922,N_24813);
nand UO_901 (O_901,N_24843,N_24770);
nand UO_902 (O_902,N_24853,N_24987);
xnor UO_903 (O_903,N_24998,N_24846);
xor UO_904 (O_904,N_24846,N_24857);
nand UO_905 (O_905,N_24930,N_24827);
nor UO_906 (O_906,N_24926,N_24920);
or UO_907 (O_907,N_24867,N_24884);
xnor UO_908 (O_908,N_24781,N_24840);
xor UO_909 (O_909,N_24908,N_24830);
or UO_910 (O_910,N_24807,N_24764);
nor UO_911 (O_911,N_24922,N_24792);
and UO_912 (O_912,N_24955,N_24996);
or UO_913 (O_913,N_24926,N_24754);
nor UO_914 (O_914,N_24962,N_24939);
xnor UO_915 (O_915,N_24826,N_24851);
nand UO_916 (O_916,N_24843,N_24814);
xor UO_917 (O_917,N_24898,N_24767);
and UO_918 (O_918,N_24764,N_24894);
and UO_919 (O_919,N_24823,N_24751);
xor UO_920 (O_920,N_24832,N_24857);
nand UO_921 (O_921,N_24968,N_24986);
xor UO_922 (O_922,N_24807,N_24827);
nand UO_923 (O_923,N_24807,N_24893);
nand UO_924 (O_924,N_24980,N_24822);
xnor UO_925 (O_925,N_24896,N_24939);
nor UO_926 (O_926,N_24859,N_24974);
and UO_927 (O_927,N_24859,N_24822);
nand UO_928 (O_928,N_24917,N_24834);
nand UO_929 (O_929,N_24845,N_24858);
and UO_930 (O_930,N_24977,N_24786);
and UO_931 (O_931,N_24840,N_24933);
and UO_932 (O_932,N_24797,N_24756);
and UO_933 (O_933,N_24842,N_24903);
nor UO_934 (O_934,N_24750,N_24873);
xor UO_935 (O_935,N_24994,N_24796);
nand UO_936 (O_936,N_24995,N_24945);
nor UO_937 (O_937,N_24820,N_24910);
xor UO_938 (O_938,N_24904,N_24758);
or UO_939 (O_939,N_24767,N_24832);
nand UO_940 (O_940,N_24960,N_24950);
nand UO_941 (O_941,N_24968,N_24956);
and UO_942 (O_942,N_24824,N_24956);
and UO_943 (O_943,N_24906,N_24921);
xnor UO_944 (O_944,N_24870,N_24820);
nor UO_945 (O_945,N_24827,N_24963);
or UO_946 (O_946,N_24953,N_24986);
nor UO_947 (O_947,N_24937,N_24951);
and UO_948 (O_948,N_24767,N_24761);
nor UO_949 (O_949,N_24831,N_24876);
nand UO_950 (O_950,N_24996,N_24846);
and UO_951 (O_951,N_24869,N_24765);
nor UO_952 (O_952,N_24943,N_24846);
or UO_953 (O_953,N_24956,N_24881);
nand UO_954 (O_954,N_24948,N_24827);
nor UO_955 (O_955,N_24801,N_24893);
or UO_956 (O_956,N_24799,N_24961);
nand UO_957 (O_957,N_24899,N_24793);
and UO_958 (O_958,N_24999,N_24766);
or UO_959 (O_959,N_24974,N_24893);
or UO_960 (O_960,N_24782,N_24775);
nand UO_961 (O_961,N_24857,N_24876);
or UO_962 (O_962,N_24931,N_24826);
nand UO_963 (O_963,N_24943,N_24996);
xnor UO_964 (O_964,N_24819,N_24848);
xnor UO_965 (O_965,N_24956,N_24980);
nor UO_966 (O_966,N_24907,N_24801);
xnor UO_967 (O_967,N_24835,N_24957);
or UO_968 (O_968,N_24810,N_24863);
xnor UO_969 (O_969,N_24850,N_24840);
nor UO_970 (O_970,N_24797,N_24781);
and UO_971 (O_971,N_24837,N_24853);
nand UO_972 (O_972,N_24751,N_24896);
nor UO_973 (O_973,N_24855,N_24760);
xor UO_974 (O_974,N_24884,N_24817);
xnor UO_975 (O_975,N_24813,N_24792);
xor UO_976 (O_976,N_24856,N_24925);
or UO_977 (O_977,N_24854,N_24884);
or UO_978 (O_978,N_24832,N_24847);
nor UO_979 (O_979,N_24880,N_24861);
or UO_980 (O_980,N_24912,N_24955);
or UO_981 (O_981,N_24931,N_24806);
xor UO_982 (O_982,N_24964,N_24764);
nand UO_983 (O_983,N_24917,N_24983);
or UO_984 (O_984,N_24770,N_24958);
and UO_985 (O_985,N_24871,N_24962);
and UO_986 (O_986,N_24880,N_24806);
nor UO_987 (O_987,N_24776,N_24874);
xor UO_988 (O_988,N_24789,N_24797);
nand UO_989 (O_989,N_24772,N_24949);
nor UO_990 (O_990,N_24965,N_24991);
or UO_991 (O_991,N_24874,N_24833);
and UO_992 (O_992,N_24916,N_24818);
xor UO_993 (O_993,N_24854,N_24838);
nor UO_994 (O_994,N_24852,N_24764);
nor UO_995 (O_995,N_24933,N_24920);
xnor UO_996 (O_996,N_24918,N_24829);
or UO_997 (O_997,N_24919,N_24811);
xor UO_998 (O_998,N_24908,N_24959);
and UO_999 (O_999,N_24796,N_24766);
xnor UO_1000 (O_1000,N_24897,N_24960);
nand UO_1001 (O_1001,N_24861,N_24858);
xnor UO_1002 (O_1002,N_24843,N_24864);
and UO_1003 (O_1003,N_24787,N_24757);
nor UO_1004 (O_1004,N_24754,N_24790);
nand UO_1005 (O_1005,N_24804,N_24884);
or UO_1006 (O_1006,N_24818,N_24967);
nor UO_1007 (O_1007,N_24990,N_24986);
xnor UO_1008 (O_1008,N_24798,N_24897);
nand UO_1009 (O_1009,N_24797,N_24821);
xnor UO_1010 (O_1010,N_24973,N_24754);
xnor UO_1011 (O_1011,N_24917,N_24795);
and UO_1012 (O_1012,N_24940,N_24999);
and UO_1013 (O_1013,N_24761,N_24808);
nor UO_1014 (O_1014,N_24838,N_24750);
nand UO_1015 (O_1015,N_24922,N_24971);
and UO_1016 (O_1016,N_24805,N_24885);
nor UO_1017 (O_1017,N_24792,N_24921);
nor UO_1018 (O_1018,N_24942,N_24975);
xnor UO_1019 (O_1019,N_24782,N_24904);
xor UO_1020 (O_1020,N_24799,N_24890);
xor UO_1021 (O_1021,N_24963,N_24952);
nor UO_1022 (O_1022,N_24875,N_24873);
xor UO_1023 (O_1023,N_24917,N_24782);
xnor UO_1024 (O_1024,N_24914,N_24754);
xor UO_1025 (O_1025,N_24797,N_24906);
nor UO_1026 (O_1026,N_24955,N_24934);
nor UO_1027 (O_1027,N_24780,N_24911);
xnor UO_1028 (O_1028,N_24974,N_24981);
nand UO_1029 (O_1029,N_24960,N_24865);
xnor UO_1030 (O_1030,N_24833,N_24974);
nand UO_1031 (O_1031,N_24960,N_24903);
nor UO_1032 (O_1032,N_24783,N_24965);
and UO_1033 (O_1033,N_24892,N_24858);
or UO_1034 (O_1034,N_24816,N_24867);
xnor UO_1035 (O_1035,N_24943,N_24866);
xor UO_1036 (O_1036,N_24847,N_24775);
or UO_1037 (O_1037,N_24771,N_24992);
nand UO_1038 (O_1038,N_24898,N_24773);
nor UO_1039 (O_1039,N_24846,N_24794);
nand UO_1040 (O_1040,N_24983,N_24813);
nor UO_1041 (O_1041,N_24878,N_24799);
or UO_1042 (O_1042,N_24818,N_24896);
nand UO_1043 (O_1043,N_24769,N_24842);
or UO_1044 (O_1044,N_24949,N_24933);
xnor UO_1045 (O_1045,N_24803,N_24930);
and UO_1046 (O_1046,N_24764,N_24838);
or UO_1047 (O_1047,N_24910,N_24770);
nand UO_1048 (O_1048,N_24811,N_24862);
or UO_1049 (O_1049,N_24891,N_24815);
xor UO_1050 (O_1050,N_24806,N_24978);
nor UO_1051 (O_1051,N_24922,N_24968);
or UO_1052 (O_1052,N_24979,N_24981);
or UO_1053 (O_1053,N_24848,N_24859);
nor UO_1054 (O_1054,N_24790,N_24824);
xor UO_1055 (O_1055,N_24919,N_24946);
or UO_1056 (O_1056,N_24813,N_24963);
or UO_1057 (O_1057,N_24772,N_24958);
xor UO_1058 (O_1058,N_24969,N_24808);
and UO_1059 (O_1059,N_24894,N_24824);
or UO_1060 (O_1060,N_24990,N_24860);
xnor UO_1061 (O_1061,N_24900,N_24963);
or UO_1062 (O_1062,N_24956,N_24969);
nor UO_1063 (O_1063,N_24967,N_24878);
nand UO_1064 (O_1064,N_24838,N_24785);
or UO_1065 (O_1065,N_24902,N_24766);
and UO_1066 (O_1066,N_24818,N_24763);
xnor UO_1067 (O_1067,N_24843,N_24769);
nor UO_1068 (O_1068,N_24941,N_24943);
xnor UO_1069 (O_1069,N_24755,N_24831);
and UO_1070 (O_1070,N_24896,N_24819);
nand UO_1071 (O_1071,N_24813,N_24793);
nor UO_1072 (O_1072,N_24963,N_24811);
nor UO_1073 (O_1073,N_24784,N_24945);
and UO_1074 (O_1074,N_24945,N_24939);
or UO_1075 (O_1075,N_24863,N_24941);
xor UO_1076 (O_1076,N_24905,N_24952);
or UO_1077 (O_1077,N_24937,N_24842);
or UO_1078 (O_1078,N_24761,N_24776);
and UO_1079 (O_1079,N_24949,N_24927);
xor UO_1080 (O_1080,N_24795,N_24885);
nand UO_1081 (O_1081,N_24935,N_24922);
nor UO_1082 (O_1082,N_24966,N_24795);
nor UO_1083 (O_1083,N_24862,N_24948);
xnor UO_1084 (O_1084,N_24915,N_24867);
nand UO_1085 (O_1085,N_24808,N_24891);
and UO_1086 (O_1086,N_24951,N_24905);
xor UO_1087 (O_1087,N_24770,N_24842);
xor UO_1088 (O_1088,N_24830,N_24778);
and UO_1089 (O_1089,N_24790,N_24781);
nand UO_1090 (O_1090,N_24775,N_24758);
nand UO_1091 (O_1091,N_24940,N_24806);
xnor UO_1092 (O_1092,N_24780,N_24810);
or UO_1093 (O_1093,N_24791,N_24986);
and UO_1094 (O_1094,N_24823,N_24908);
or UO_1095 (O_1095,N_24871,N_24780);
nor UO_1096 (O_1096,N_24993,N_24902);
xnor UO_1097 (O_1097,N_24770,N_24997);
or UO_1098 (O_1098,N_24896,N_24861);
and UO_1099 (O_1099,N_24901,N_24915);
or UO_1100 (O_1100,N_24755,N_24813);
nand UO_1101 (O_1101,N_24817,N_24975);
or UO_1102 (O_1102,N_24965,N_24834);
and UO_1103 (O_1103,N_24852,N_24978);
nand UO_1104 (O_1104,N_24750,N_24928);
or UO_1105 (O_1105,N_24937,N_24848);
and UO_1106 (O_1106,N_24839,N_24860);
nand UO_1107 (O_1107,N_24782,N_24906);
nor UO_1108 (O_1108,N_24843,N_24962);
nor UO_1109 (O_1109,N_24824,N_24867);
nand UO_1110 (O_1110,N_24770,N_24909);
nor UO_1111 (O_1111,N_24815,N_24851);
nor UO_1112 (O_1112,N_24850,N_24959);
nor UO_1113 (O_1113,N_24973,N_24877);
xor UO_1114 (O_1114,N_24787,N_24886);
and UO_1115 (O_1115,N_24980,N_24850);
nand UO_1116 (O_1116,N_24824,N_24862);
or UO_1117 (O_1117,N_24981,N_24802);
or UO_1118 (O_1118,N_24846,N_24860);
nand UO_1119 (O_1119,N_24992,N_24832);
and UO_1120 (O_1120,N_24928,N_24788);
nor UO_1121 (O_1121,N_24852,N_24761);
nand UO_1122 (O_1122,N_24764,N_24756);
xnor UO_1123 (O_1123,N_24985,N_24955);
and UO_1124 (O_1124,N_24818,N_24995);
and UO_1125 (O_1125,N_24827,N_24843);
or UO_1126 (O_1126,N_24781,N_24959);
and UO_1127 (O_1127,N_24923,N_24804);
or UO_1128 (O_1128,N_24827,N_24856);
and UO_1129 (O_1129,N_24798,N_24930);
and UO_1130 (O_1130,N_24836,N_24922);
and UO_1131 (O_1131,N_24927,N_24868);
nor UO_1132 (O_1132,N_24784,N_24965);
and UO_1133 (O_1133,N_24924,N_24814);
xor UO_1134 (O_1134,N_24787,N_24997);
and UO_1135 (O_1135,N_24765,N_24849);
and UO_1136 (O_1136,N_24954,N_24944);
nor UO_1137 (O_1137,N_24951,N_24808);
xor UO_1138 (O_1138,N_24896,N_24906);
and UO_1139 (O_1139,N_24866,N_24872);
xnor UO_1140 (O_1140,N_24826,N_24969);
and UO_1141 (O_1141,N_24791,N_24955);
or UO_1142 (O_1142,N_24882,N_24823);
xnor UO_1143 (O_1143,N_24935,N_24768);
xor UO_1144 (O_1144,N_24753,N_24826);
nor UO_1145 (O_1145,N_24880,N_24898);
or UO_1146 (O_1146,N_24790,N_24922);
nand UO_1147 (O_1147,N_24832,N_24793);
and UO_1148 (O_1148,N_24832,N_24958);
nor UO_1149 (O_1149,N_24808,N_24879);
and UO_1150 (O_1150,N_24776,N_24793);
nand UO_1151 (O_1151,N_24980,N_24952);
xor UO_1152 (O_1152,N_24934,N_24864);
nand UO_1153 (O_1153,N_24840,N_24905);
nand UO_1154 (O_1154,N_24776,N_24983);
xnor UO_1155 (O_1155,N_24763,N_24961);
or UO_1156 (O_1156,N_24937,N_24943);
nor UO_1157 (O_1157,N_24985,N_24943);
nor UO_1158 (O_1158,N_24967,N_24901);
or UO_1159 (O_1159,N_24802,N_24903);
nor UO_1160 (O_1160,N_24773,N_24811);
and UO_1161 (O_1161,N_24929,N_24906);
or UO_1162 (O_1162,N_24904,N_24995);
or UO_1163 (O_1163,N_24894,N_24976);
and UO_1164 (O_1164,N_24839,N_24848);
nand UO_1165 (O_1165,N_24955,N_24816);
nor UO_1166 (O_1166,N_24821,N_24862);
or UO_1167 (O_1167,N_24781,N_24970);
xnor UO_1168 (O_1168,N_24862,N_24760);
and UO_1169 (O_1169,N_24855,N_24921);
xor UO_1170 (O_1170,N_24871,N_24997);
xnor UO_1171 (O_1171,N_24809,N_24894);
or UO_1172 (O_1172,N_24908,N_24894);
nor UO_1173 (O_1173,N_24994,N_24927);
or UO_1174 (O_1174,N_24788,N_24916);
or UO_1175 (O_1175,N_24939,N_24839);
and UO_1176 (O_1176,N_24938,N_24896);
nand UO_1177 (O_1177,N_24797,N_24885);
xnor UO_1178 (O_1178,N_24792,N_24894);
and UO_1179 (O_1179,N_24839,N_24960);
and UO_1180 (O_1180,N_24792,N_24805);
and UO_1181 (O_1181,N_24965,N_24922);
or UO_1182 (O_1182,N_24874,N_24929);
nor UO_1183 (O_1183,N_24877,N_24789);
and UO_1184 (O_1184,N_24936,N_24960);
xor UO_1185 (O_1185,N_24921,N_24802);
xnor UO_1186 (O_1186,N_24817,N_24973);
xor UO_1187 (O_1187,N_24925,N_24812);
nor UO_1188 (O_1188,N_24818,N_24864);
nor UO_1189 (O_1189,N_24875,N_24967);
nand UO_1190 (O_1190,N_24946,N_24896);
nor UO_1191 (O_1191,N_24798,N_24868);
and UO_1192 (O_1192,N_24963,N_24988);
xor UO_1193 (O_1193,N_24825,N_24865);
and UO_1194 (O_1194,N_24757,N_24865);
and UO_1195 (O_1195,N_24973,N_24831);
nor UO_1196 (O_1196,N_24771,N_24786);
xor UO_1197 (O_1197,N_24929,N_24789);
nand UO_1198 (O_1198,N_24829,N_24886);
nand UO_1199 (O_1199,N_24928,N_24857);
or UO_1200 (O_1200,N_24774,N_24911);
and UO_1201 (O_1201,N_24883,N_24958);
nand UO_1202 (O_1202,N_24820,N_24874);
and UO_1203 (O_1203,N_24819,N_24902);
nor UO_1204 (O_1204,N_24933,N_24801);
xor UO_1205 (O_1205,N_24873,N_24838);
nand UO_1206 (O_1206,N_24914,N_24815);
nor UO_1207 (O_1207,N_24985,N_24806);
or UO_1208 (O_1208,N_24774,N_24922);
nand UO_1209 (O_1209,N_24801,N_24953);
and UO_1210 (O_1210,N_24866,N_24831);
nor UO_1211 (O_1211,N_24888,N_24813);
xnor UO_1212 (O_1212,N_24939,N_24912);
nand UO_1213 (O_1213,N_24848,N_24908);
and UO_1214 (O_1214,N_24889,N_24915);
nand UO_1215 (O_1215,N_24998,N_24859);
and UO_1216 (O_1216,N_24801,N_24770);
or UO_1217 (O_1217,N_24828,N_24813);
and UO_1218 (O_1218,N_24986,N_24899);
xnor UO_1219 (O_1219,N_24815,N_24860);
and UO_1220 (O_1220,N_24913,N_24908);
or UO_1221 (O_1221,N_24889,N_24910);
nand UO_1222 (O_1222,N_24791,N_24833);
xor UO_1223 (O_1223,N_24820,N_24986);
nor UO_1224 (O_1224,N_24820,N_24804);
or UO_1225 (O_1225,N_24815,N_24863);
nand UO_1226 (O_1226,N_24901,N_24998);
nor UO_1227 (O_1227,N_24932,N_24967);
or UO_1228 (O_1228,N_24785,N_24752);
and UO_1229 (O_1229,N_24902,N_24970);
nor UO_1230 (O_1230,N_24811,N_24768);
nand UO_1231 (O_1231,N_24868,N_24960);
nor UO_1232 (O_1232,N_24861,N_24766);
or UO_1233 (O_1233,N_24906,N_24819);
and UO_1234 (O_1234,N_24900,N_24841);
nor UO_1235 (O_1235,N_24990,N_24927);
and UO_1236 (O_1236,N_24759,N_24830);
and UO_1237 (O_1237,N_24978,N_24989);
nor UO_1238 (O_1238,N_24949,N_24855);
and UO_1239 (O_1239,N_24832,N_24798);
xor UO_1240 (O_1240,N_24820,N_24962);
and UO_1241 (O_1241,N_24958,N_24917);
and UO_1242 (O_1242,N_24996,N_24818);
nand UO_1243 (O_1243,N_24942,N_24963);
or UO_1244 (O_1244,N_24845,N_24902);
xor UO_1245 (O_1245,N_24980,N_24972);
and UO_1246 (O_1246,N_24912,N_24956);
xor UO_1247 (O_1247,N_24925,N_24841);
or UO_1248 (O_1248,N_24763,N_24967);
nor UO_1249 (O_1249,N_24995,N_24928);
or UO_1250 (O_1250,N_24795,N_24897);
and UO_1251 (O_1251,N_24785,N_24799);
or UO_1252 (O_1252,N_24814,N_24888);
xnor UO_1253 (O_1253,N_24847,N_24858);
or UO_1254 (O_1254,N_24753,N_24996);
and UO_1255 (O_1255,N_24752,N_24790);
nor UO_1256 (O_1256,N_24917,N_24784);
nand UO_1257 (O_1257,N_24816,N_24895);
nand UO_1258 (O_1258,N_24908,N_24757);
or UO_1259 (O_1259,N_24983,N_24790);
xor UO_1260 (O_1260,N_24810,N_24971);
or UO_1261 (O_1261,N_24822,N_24898);
or UO_1262 (O_1262,N_24887,N_24843);
xor UO_1263 (O_1263,N_24913,N_24914);
and UO_1264 (O_1264,N_24866,N_24811);
nor UO_1265 (O_1265,N_24814,N_24916);
xnor UO_1266 (O_1266,N_24897,N_24888);
nor UO_1267 (O_1267,N_24811,N_24851);
or UO_1268 (O_1268,N_24963,N_24770);
and UO_1269 (O_1269,N_24869,N_24851);
xor UO_1270 (O_1270,N_24892,N_24783);
nand UO_1271 (O_1271,N_24992,N_24800);
nand UO_1272 (O_1272,N_24865,N_24913);
nand UO_1273 (O_1273,N_24952,N_24906);
xnor UO_1274 (O_1274,N_24787,N_24870);
and UO_1275 (O_1275,N_24778,N_24887);
and UO_1276 (O_1276,N_24839,N_24994);
and UO_1277 (O_1277,N_24879,N_24913);
and UO_1278 (O_1278,N_24769,N_24761);
and UO_1279 (O_1279,N_24981,N_24852);
nand UO_1280 (O_1280,N_24934,N_24923);
or UO_1281 (O_1281,N_24958,N_24764);
or UO_1282 (O_1282,N_24807,N_24812);
and UO_1283 (O_1283,N_24866,N_24881);
nor UO_1284 (O_1284,N_24794,N_24953);
nand UO_1285 (O_1285,N_24954,N_24815);
xor UO_1286 (O_1286,N_24851,N_24906);
nand UO_1287 (O_1287,N_24998,N_24902);
nand UO_1288 (O_1288,N_24932,N_24885);
or UO_1289 (O_1289,N_24766,N_24996);
and UO_1290 (O_1290,N_24980,N_24777);
nor UO_1291 (O_1291,N_24903,N_24958);
nand UO_1292 (O_1292,N_24989,N_24755);
nor UO_1293 (O_1293,N_24895,N_24964);
or UO_1294 (O_1294,N_24924,N_24879);
nand UO_1295 (O_1295,N_24960,N_24825);
xnor UO_1296 (O_1296,N_24838,N_24811);
xor UO_1297 (O_1297,N_24982,N_24976);
or UO_1298 (O_1298,N_24750,N_24817);
nand UO_1299 (O_1299,N_24969,N_24763);
and UO_1300 (O_1300,N_24922,N_24859);
nand UO_1301 (O_1301,N_24912,N_24884);
nand UO_1302 (O_1302,N_24846,N_24915);
nor UO_1303 (O_1303,N_24843,N_24916);
xor UO_1304 (O_1304,N_24773,N_24819);
nand UO_1305 (O_1305,N_24833,N_24836);
or UO_1306 (O_1306,N_24993,N_24821);
and UO_1307 (O_1307,N_24791,N_24757);
nand UO_1308 (O_1308,N_24794,N_24785);
xor UO_1309 (O_1309,N_24960,N_24798);
and UO_1310 (O_1310,N_24969,N_24824);
nor UO_1311 (O_1311,N_24816,N_24825);
and UO_1312 (O_1312,N_24835,N_24923);
nor UO_1313 (O_1313,N_24969,N_24971);
or UO_1314 (O_1314,N_24922,N_24924);
or UO_1315 (O_1315,N_24958,N_24806);
xnor UO_1316 (O_1316,N_24957,N_24966);
nor UO_1317 (O_1317,N_24978,N_24879);
nor UO_1318 (O_1318,N_24995,N_24939);
or UO_1319 (O_1319,N_24774,N_24940);
or UO_1320 (O_1320,N_24860,N_24780);
nand UO_1321 (O_1321,N_24929,N_24830);
xnor UO_1322 (O_1322,N_24961,N_24832);
nand UO_1323 (O_1323,N_24982,N_24909);
nor UO_1324 (O_1324,N_24765,N_24763);
and UO_1325 (O_1325,N_24908,N_24869);
and UO_1326 (O_1326,N_24968,N_24862);
xnor UO_1327 (O_1327,N_24932,N_24845);
xor UO_1328 (O_1328,N_24779,N_24917);
or UO_1329 (O_1329,N_24753,N_24927);
nand UO_1330 (O_1330,N_24909,N_24820);
or UO_1331 (O_1331,N_24863,N_24772);
xor UO_1332 (O_1332,N_24752,N_24915);
nand UO_1333 (O_1333,N_24816,N_24960);
and UO_1334 (O_1334,N_24965,N_24917);
and UO_1335 (O_1335,N_24988,N_24997);
or UO_1336 (O_1336,N_24765,N_24963);
and UO_1337 (O_1337,N_24790,N_24890);
nand UO_1338 (O_1338,N_24753,N_24854);
or UO_1339 (O_1339,N_24959,N_24887);
nor UO_1340 (O_1340,N_24995,N_24916);
nand UO_1341 (O_1341,N_24930,N_24910);
xnor UO_1342 (O_1342,N_24813,N_24913);
and UO_1343 (O_1343,N_24878,N_24855);
nor UO_1344 (O_1344,N_24950,N_24867);
xor UO_1345 (O_1345,N_24945,N_24942);
or UO_1346 (O_1346,N_24825,N_24925);
nand UO_1347 (O_1347,N_24888,N_24988);
nor UO_1348 (O_1348,N_24859,N_24883);
xor UO_1349 (O_1349,N_24879,N_24846);
nor UO_1350 (O_1350,N_24779,N_24975);
and UO_1351 (O_1351,N_24841,N_24800);
and UO_1352 (O_1352,N_24871,N_24952);
nor UO_1353 (O_1353,N_24942,N_24929);
or UO_1354 (O_1354,N_24805,N_24826);
or UO_1355 (O_1355,N_24907,N_24763);
nor UO_1356 (O_1356,N_24823,N_24762);
nand UO_1357 (O_1357,N_24971,N_24882);
nor UO_1358 (O_1358,N_24781,N_24863);
xnor UO_1359 (O_1359,N_24779,N_24841);
and UO_1360 (O_1360,N_24940,N_24819);
nor UO_1361 (O_1361,N_24889,N_24876);
nand UO_1362 (O_1362,N_24799,N_24847);
or UO_1363 (O_1363,N_24994,N_24968);
xor UO_1364 (O_1364,N_24920,N_24908);
or UO_1365 (O_1365,N_24857,N_24943);
xnor UO_1366 (O_1366,N_24760,N_24971);
nor UO_1367 (O_1367,N_24770,N_24795);
nand UO_1368 (O_1368,N_24973,N_24924);
nor UO_1369 (O_1369,N_24820,N_24861);
nand UO_1370 (O_1370,N_24764,N_24840);
or UO_1371 (O_1371,N_24958,N_24881);
and UO_1372 (O_1372,N_24969,N_24920);
xor UO_1373 (O_1373,N_24767,N_24862);
xor UO_1374 (O_1374,N_24899,N_24847);
nor UO_1375 (O_1375,N_24982,N_24768);
and UO_1376 (O_1376,N_24967,N_24830);
and UO_1377 (O_1377,N_24908,N_24837);
xor UO_1378 (O_1378,N_24983,N_24920);
nand UO_1379 (O_1379,N_24873,N_24830);
or UO_1380 (O_1380,N_24878,N_24825);
and UO_1381 (O_1381,N_24976,N_24909);
xor UO_1382 (O_1382,N_24903,N_24854);
or UO_1383 (O_1383,N_24936,N_24887);
or UO_1384 (O_1384,N_24842,N_24812);
and UO_1385 (O_1385,N_24788,N_24953);
nor UO_1386 (O_1386,N_24937,N_24875);
nand UO_1387 (O_1387,N_24999,N_24857);
nor UO_1388 (O_1388,N_24810,N_24850);
nor UO_1389 (O_1389,N_24895,N_24928);
and UO_1390 (O_1390,N_24846,N_24952);
nor UO_1391 (O_1391,N_24942,N_24763);
nor UO_1392 (O_1392,N_24958,N_24956);
nand UO_1393 (O_1393,N_24838,N_24912);
nor UO_1394 (O_1394,N_24999,N_24855);
or UO_1395 (O_1395,N_24942,N_24910);
xnor UO_1396 (O_1396,N_24797,N_24861);
and UO_1397 (O_1397,N_24885,N_24902);
xor UO_1398 (O_1398,N_24982,N_24794);
xor UO_1399 (O_1399,N_24818,N_24782);
nor UO_1400 (O_1400,N_24965,N_24853);
nor UO_1401 (O_1401,N_24777,N_24853);
and UO_1402 (O_1402,N_24872,N_24894);
or UO_1403 (O_1403,N_24801,N_24936);
nand UO_1404 (O_1404,N_24805,N_24839);
xnor UO_1405 (O_1405,N_24782,N_24755);
and UO_1406 (O_1406,N_24964,N_24769);
or UO_1407 (O_1407,N_24757,N_24988);
nor UO_1408 (O_1408,N_24758,N_24817);
nand UO_1409 (O_1409,N_24870,N_24953);
or UO_1410 (O_1410,N_24886,N_24846);
or UO_1411 (O_1411,N_24844,N_24790);
nand UO_1412 (O_1412,N_24897,N_24927);
nor UO_1413 (O_1413,N_24781,N_24782);
xor UO_1414 (O_1414,N_24792,N_24836);
nor UO_1415 (O_1415,N_24869,N_24847);
nor UO_1416 (O_1416,N_24781,N_24881);
or UO_1417 (O_1417,N_24792,N_24780);
and UO_1418 (O_1418,N_24887,N_24800);
or UO_1419 (O_1419,N_24781,N_24846);
and UO_1420 (O_1420,N_24942,N_24750);
and UO_1421 (O_1421,N_24838,N_24797);
or UO_1422 (O_1422,N_24969,N_24833);
nand UO_1423 (O_1423,N_24899,N_24791);
xnor UO_1424 (O_1424,N_24910,N_24992);
nor UO_1425 (O_1425,N_24829,N_24799);
or UO_1426 (O_1426,N_24902,N_24945);
nand UO_1427 (O_1427,N_24866,N_24758);
nand UO_1428 (O_1428,N_24980,N_24801);
xnor UO_1429 (O_1429,N_24971,N_24859);
nand UO_1430 (O_1430,N_24879,N_24985);
nor UO_1431 (O_1431,N_24812,N_24755);
and UO_1432 (O_1432,N_24985,N_24793);
nand UO_1433 (O_1433,N_24776,N_24887);
or UO_1434 (O_1434,N_24914,N_24844);
and UO_1435 (O_1435,N_24798,N_24982);
nor UO_1436 (O_1436,N_24886,N_24990);
and UO_1437 (O_1437,N_24772,N_24758);
nand UO_1438 (O_1438,N_24836,N_24912);
or UO_1439 (O_1439,N_24838,N_24828);
or UO_1440 (O_1440,N_24940,N_24841);
nor UO_1441 (O_1441,N_24920,N_24915);
and UO_1442 (O_1442,N_24993,N_24895);
xor UO_1443 (O_1443,N_24805,N_24753);
xor UO_1444 (O_1444,N_24985,N_24829);
nor UO_1445 (O_1445,N_24924,N_24844);
nor UO_1446 (O_1446,N_24872,N_24870);
and UO_1447 (O_1447,N_24993,N_24963);
nor UO_1448 (O_1448,N_24929,N_24902);
xnor UO_1449 (O_1449,N_24953,N_24888);
nor UO_1450 (O_1450,N_24883,N_24975);
nor UO_1451 (O_1451,N_24889,N_24988);
xor UO_1452 (O_1452,N_24881,N_24917);
xnor UO_1453 (O_1453,N_24790,N_24766);
nand UO_1454 (O_1454,N_24919,N_24786);
nor UO_1455 (O_1455,N_24903,N_24765);
and UO_1456 (O_1456,N_24766,N_24776);
and UO_1457 (O_1457,N_24867,N_24753);
nand UO_1458 (O_1458,N_24913,N_24926);
xnor UO_1459 (O_1459,N_24981,N_24824);
xor UO_1460 (O_1460,N_24776,N_24965);
nand UO_1461 (O_1461,N_24851,N_24898);
or UO_1462 (O_1462,N_24981,N_24854);
or UO_1463 (O_1463,N_24865,N_24771);
nor UO_1464 (O_1464,N_24949,N_24769);
and UO_1465 (O_1465,N_24976,N_24937);
and UO_1466 (O_1466,N_24948,N_24854);
and UO_1467 (O_1467,N_24797,N_24999);
or UO_1468 (O_1468,N_24926,N_24888);
or UO_1469 (O_1469,N_24834,N_24809);
nor UO_1470 (O_1470,N_24777,N_24927);
or UO_1471 (O_1471,N_24890,N_24942);
nand UO_1472 (O_1472,N_24864,N_24800);
and UO_1473 (O_1473,N_24873,N_24899);
nand UO_1474 (O_1474,N_24874,N_24915);
or UO_1475 (O_1475,N_24900,N_24977);
nor UO_1476 (O_1476,N_24839,N_24954);
xnor UO_1477 (O_1477,N_24750,N_24811);
or UO_1478 (O_1478,N_24967,N_24855);
or UO_1479 (O_1479,N_24860,N_24821);
nor UO_1480 (O_1480,N_24900,N_24776);
nor UO_1481 (O_1481,N_24764,N_24792);
xor UO_1482 (O_1482,N_24843,N_24822);
and UO_1483 (O_1483,N_24915,N_24825);
and UO_1484 (O_1484,N_24865,N_24929);
xor UO_1485 (O_1485,N_24853,N_24926);
xnor UO_1486 (O_1486,N_24756,N_24993);
nor UO_1487 (O_1487,N_24813,N_24779);
or UO_1488 (O_1488,N_24982,N_24908);
xor UO_1489 (O_1489,N_24919,N_24767);
xor UO_1490 (O_1490,N_24801,N_24766);
nor UO_1491 (O_1491,N_24878,N_24800);
nand UO_1492 (O_1492,N_24863,N_24756);
and UO_1493 (O_1493,N_24867,N_24764);
or UO_1494 (O_1494,N_24960,N_24993);
xor UO_1495 (O_1495,N_24862,N_24905);
and UO_1496 (O_1496,N_24781,N_24805);
nand UO_1497 (O_1497,N_24927,N_24987);
nand UO_1498 (O_1498,N_24936,N_24988);
nor UO_1499 (O_1499,N_24893,N_24798);
or UO_1500 (O_1500,N_24775,N_24762);
xor UO_1501 (O_1501,N_24931,N_24818);
and UO_1502 (O_1502,N_24774,N_24858);
or UO_1503 (O_1503,N_24791,N_24877);
nor UO_1504 (O_1504,N_24985,N_24890);
or UO_1505 (O_1505,N_24932,N_24760);
and UO_1506 (O_1506,N_24998,N_24914);
xor UO_1507 (O_1507,N_24755,N_24760);
nand UO_1508 (O_1508,N_24929,N_24954);
and UO_1509 (O_1509,N_24859,N_24982);
nand UO_1510 (O_1510,N_24799,N_24905);
or UO_1511 (O_1511,N_24966,N_24787);
or UO_1512 (O_1512,N_24768,N_24788);
or UO_1513 (O_1513,N_24860,N_24994);
nor UO_1514 (O_1514,N_24767,N_24902);
or UO_1515 (O_1515,N_24816,N_24962);
nor UO_1516 (O_1516,N_24779,N_24929);
and UO_1517 (O_1517,N_24754,N_24982);
xnor UO_1518 (O_1518,N_24821,N_24890);
and UO_1519 (O_1519,N_24968,N_24890);
xnor UO_1520 (O_1520,N_24998,N_24899);
nor UO_1521 (O_1521,N_24982,N_24752);
or UO_1522 (O_1522,N_24897,N_24861);
nor UO_1523 (O_1523,N_24754,N_24941);
nand UO_1524 (O_1524,N_24957,N_24933);
or UO_1525 (O_1525,N_24859,N_24755);
and UO_1526 (O_1526,N_24974,N_24976);
nand UO_1527 (O_1527,N_24947,N_24828);
nor UO_1528 (O_1528,N_24765,N_24865);
xnor UO_1529 (O_1529,N_24773,N_24844);
xor UO_1530 (O_1530,N_24936,N_24789);
and UO_1531 (O_1531,N_24890,N_24805);
or UO_1532 (O_1532,N_24883,N_24941);
xor UO_1533 (O_1533,N_24878,N_24846);
xor UO_1534 (O_1534,N_24758,N_24909);
and UO_1535 (O_1535,N_24942,N_24918);
nor UO_1536 (O_1536,N_24910,N_24893);
nand UO_1537 (O_1537,N_24989,N_24863);
or UO_1538 (O_1538,N_24901,N_24920);
xnor UO_1539 (O_1539,N_24973,N_24810);
nor UO_1540 (O_1540,N_24910,N_24752);
or UO_1541 (O_1541,N_24906,N_24922);
or UO_1542 (O_1542,N_24797,N_24974);
and UO_1543 (O_1543,N_24834,N_24849);
xnor UO_1544 (O_1544,N_24986,N_24915);
xor UO_1545 (O_1545,N_24935,N_24910);
nor UO_1546 (O_1546,N_24822,N_24856);
or UO_1547 (O_1547,N_24917,N_24895);
nor UO_1548 (O_1548,N_24961,N_24841);
xor UO_1549 (O_1549,N_24772,N_24911);
nor UO_1550 (O_1550,N_24801,N_24765);
and UO_1551 (O_1551,N_24761,N_24847);
or UO_1552 (O_1552,N_24774,N_24865);
xor UO_1553 (O_1553,N_24941,N_24757);
xnor UO_1554 (O_1554,N_24797,N_24995);
and UO_1555 (O_1555,N_24901,N_24861);
nand UO_1556 (O_1556,N_24797,N_24944);
xnor UO_1557 (O_1557,N_24988,N_24810);
and UO_1558 (O_1558,N_24758,N_24818);
nor UO_1559 (O_1559,N_24981,N_24866);
nand UO_1560 (O_1560,N_24781,N_24935);
nor UO_1561 (O_1561,N_24764,N_24896);
nand UO_1562 (O_1562,N_24910,N_24972);
nand UO_1563 (O_1563,N_24903,N_24862);
nor UO_1564 (O_1564,N_24825,N_24822);
or UO_1565 (O_1565,N_24800,N_24803);
or UO_1566 (O_1566,N_24814,N_24927);
nand UO_1567 (O_1567,N_24890,N_24885);
nand UO_1568 (O_1568,N_24974,N_24774);
nor UO_1569 (O_1569,N_24895,N_24806);
nor UO_1570 (O_1570,N_24913,N_24957);
nand UO_1571 (O_1571,N_24865,N_24925);
xnor UO_1572 (O_1572,N_24760,N_24857);
xor UO_1573 (O_1573,N_24798,N_24804);
or UO_1574 (O_1574,N_24809,N_24947);
and UO_1575 (O_1575,N_24904,N_24886);
or UO_1576 (O_1576,N_24973,N_24890);
nand UO_1577 (O_1577,N_24973,N_24903);
and UO_1578 (O_1578,N_24772,N_24918);
nand UO_1579 (O_1579,N_24960,N_24922);
or UO_1580 (O_1580,N_24859,N_24917);
and UO_1581 (O_1581,N_24945,N_24958);
or UO_1582 (O_1582,N_24803,N_24944);
xor UO_1583 (O_1583,N_24958,N_24866);
nor UO_1584 (O_1584,N_24848,N_24775);
nand UO_1585 (O_1585,N_24963,N_24877);
nand UO_1586 (O_1586,N_24792,N_24891);
xnor UO_1587 (O_1587,N_24839,N_24762);
xor UO_1588 (O_1588,N_24958,N_24851);
xor UO_1589 (O_1589,N_24889,N_24777);
and UO_1590 (O_1590,N_24891,N_24966);
xor UO_1591 (O_1591,N_24955,N_24871);
and UO_1592 (O_1592,N_24890,N_24855);
xor UO_1593 (O_1593,N_24778,N_24926);
or UO_1594 (O_1594,N_24978,N_24873);
nand UO_1595 (O_1595,N_24763,N_24917);
or UO_1596 (O_1596,N_24942,N_24860);
or UO_1597 (O_1597,N_24799,N_24941);
or UO_1598 (O_1598,N_24944,N_24971);
and UO_1599 (O_1599,N_24855,N_24771);
nand UO_1600 (O_1600,N_24944,N_24903);
nand UO_1601 (O_1601,N_24847,N_24843);
and UO_1602 (O_1602,N_24872,N_24767);
or UO_1603 (O_1603,N_24776,N_24861);
or UO_1604 (O_1604,N_24847,N_24915);
or UO_1605 (O_1605,N_24769,N_24786);
nand UO_1606 (O_1606,N_24862,N_24859);
xnor UO_1607 (O_1607,N_24842,N_24790);
or UO_1608 (O_1608,N_24773,N_24981);
or UO_1609 (O_1609,N_24944,N_24926);
nor UO_1610 (O_1610,N_24845,N_24776);
nor UO_1611 (O_1611,N_24999,N_24781);
or UO_1612 (O_1612,N_24896,N_24836);
or UO_1613 (O_1613,N_24831,N_24895);
and UO_1614 (O_1614,N_24760,N_24782);
nor UO_1615 (O_1615,N_24790,N_24946);
xor UO_1616 (O_1616,N_24967,N_24981);
nor UO_1617 (O_1617,N_24782,N_24751);
or UO_1618 (O_1618,N_24964,N_24986);
nand UO_1619 (O_1619,N_24963,N_24978);
nand UO_1620 (O_1620,N_24940,N_24839);
and UO_1621 (O_1621,N_24796,N_24823);
and UO_1622 (O_1622,N_24847,N_24971);
nor UO_1623 (O_1623,N_24831,N_24821);
nor UO_1624 (O_1624,N_24813,N_24898);
nor UO_1625 (O_1625,N_24986,N_24981);
nor UO_1626 (O_1626,N_24783,N_24996);
nor UO_1627 (O_1627,N_24751,N_24852);
nor UO_1628 (O_1628,N_24784,N_24950);
nand UO_1629 (O_1629,N_24890,N_24843);
or UO_1630 (O_1630,N_24844,N_24850);
and UO_1631 (O_1631,N_24765,N_24959);
nor UO_1632 (O_1632,N_24962,N_24848);
and UO_1633 (O_1633,N_24876,N_24922);
nand UO_1634 (O_1634,N_24908,N_24842);
nor UO_1635 (O_1635,N_24813,N_24860);
and UO_1636 (O_1636,N_24944,N_24889);
nand UO_1637 (O_1637,N_24970,N_24927);
nor UO_1638 (O_1638,N_24814,N_24884);
or UO_1639 (O_1639,N_24865,N_24939);
nor UO_1640 (O_1640,N_24778,N_24961);
xor UO_1641 (O_1641,N_24893,N_24795);
xor UO_1642 (O_1642,N_24855,N_24796);
nand UO_1643 (O_1643,N_24857,N_24766);
and UO_1644 (O_1644,N_24932,N_24995);
xor UO_1645 (O_1645,N_24816,N_24838);
nand UO_1646 (O_1646,N_24878,N_24751);
and UO_1647 (O_1647,N_24977,N_24856);
xnor UO_1648 (O_1648,N_24805,N_24756);
nand UO_1649 (O_1649,N_24799,N_24911);
nor UO_1650 (O_1650,N_24984,N_24990);
nor UO_1651 (O_1651,N_24751,N_24789);
nor UO_1652 (O_1652,N_24901,N_24881);
nand UO_1653 (O_1653,N_24857,N_24855);
or UO_1654 (O_1654,N_24763,N_24918);
xnor UO_1655 (O_1655,N_24817,N_24845);
and UO_1656 (O_1656,N_24961,N_24948);
and UO_1657 (O_1657,N_24838,N_24904);
xor UO_1658 (O_1658,N_24780,N_24770);
or UO_1659 (O_1659,N_24840,N_24844);
or UO_1660 (O_1660,N_24885,N_24918);
and UO_1661 (O_1661,N_24868,N_24782);
or UO_1662 (O_1662,N_24759,N_24985);
xor UO_1663 (O_1663,N_24968,N_24824);
or UO_1664 (O_1664,N_24936,N_24807);
nor UO_1665 (O_1665,N_24814,N_24784);
and UO_1666 (O_1666,N_24948,N_24986);
nand UO_1667 (O_1667,N_24992,N_24765);
and UO_1668 (O_1668,N_24835,N_24997);
nor UO_1669 (O_1669,N_24898,N_24826);
or UO_1670 (O_1670,N_24750,N_24813);
nor UO_1671 (O_1671,N_24879,N_24903);
nand UO_1672 (O_1672,N_24912,N_24778);
xnor UO_1673 (O_1673,N_24946,N_24835);
or UO_1674 (O_1674,N_24835,N_24975);
and UO_1675 (O_1675,N_24916,N_24965);
or UO_1676 (O_1676,N_24986,N_24900);
nor UO_1677 (O_1677,N_24890,N_24809);
nor UO_1678 (O_1678,N_24945,N_24863);
and UO_1679 (O_1679,N_24917,N_24787);
xor UO_1680 (O_1680,N_24879,N_24811);
xor UO_1681 (O_1681,N_24877,N_24755);
nor UO_1682 (O_1682,N_24821,N_24982);
and UO_1683 (O_1683,N_24929,N_24886);
and UO_1684 (O_1684,N_24860,N_24971);
nand UO_1685 (O_1685,N_24790,N_24848);
nand UO_1686 (O_1686,N_24841,N_24913);
nand UO_1687 (O_1687,N_24940,N_24870);
and UO_1688 (O_1688,N_24790,N_24840);
or UO_1689 (O_1689,N_24980,N_24853);
or UO_1690 (O_1690,N_24921,N_24990);
nand UO_1691 (O_1691,N_24846,N_24896);
and UO_1692 (O_1692,N_24800,N_24946);
nand UO_1693 (O_1693,N_24823,N_24895);
or UO_1694 (O_1694,N_24964,N_24856);
and UO_1695 (O_1695,N_24839,N_24856);
and UO_1696 (O_1696,N_24934,N_24890);
or UO_1697 (O_1697,N_24834,N_24803);
or UO_1698 (O_1698,N_24870,N_24971);
nand UO_1699 (O_1699,N_24815,N_24970);
nor UO_1700 (O_1700,N_24986,N_24993);
nor UO_1701 (O_1701,N_24945,N_24969);
or UO_1702 (O_1702,N_24799,N_24767);
or UO_1703 (O_1703,N_24949,N_24962);
nand UO_1704 (O_1704,N_24952,N_24884);
nor UO_1705 (O_1705,N_24846,N_24810);
xor UO_1706 (O_1706,N_24754,N_24820);
and UO_1707 (O_1707,N_24821,N_24791);
or UO_1708 (O_1708,N_24806,N_24876);
or UO_1709 (O_1709,N_24843,N_24756);
nor UO_1710 (O_1710,N_24894,N_24852);
and UO_1711 (O_1711,N_24938,N_24999);
or UO_1712 (O_1712,N_24760,N_24806);
nand UO_1713 (O_1713,N_24869,N_24781);
nand UO_1714 (O_1714,N_24935,N_24838);
nor UO_1715 (O_1715,N_24828,N_24986);
and UO_1716 (O_1716,N_24865,N_24983);
and UO_1717 (O_1717,N_24941,N_24928);
nor UO_1718 (O_1718,N_24924,N_24911);
nor UO_1719 (O_1719,N_24986,N_24865);
and UO_1720 (O_1720,N_24915,N_24932);
and UO_1721 (O_1721,N_24998,N_24814);
and UO_1722 (O_1722,N_24814,N_24925);
xor UO_1723 (O_1723,N_24906,N_24876);
nor UO_1724 (O_1724,N_24863,N_24845);
and UO_1725 (O_1725,N_24893,N_24830);
and UO_1726 (O_1726,N_24899,N_24859);
nor UO_1727 (O_1727,N_24845,N_24890);
xnor UO_1728 (O_1728,N_24796,N_24954);
or UO_1729 (O_1729,N_24823,N_24986);
or UO_1730 (O_1730,N_24865,N_24772);
and UO_1731 (O_1731,N_24928,N_24997);
xnor UO_1732 (O_1732,N_24805,N_24965);
xor UO_1733 (O_1733,N_24777,N_24899);
nor UO_1734 (O_1734,N_24784,N_24825);
nor UO_1735 (O_1735,N_24818,N_24778);
and UO_1736 (O_1736,N_24766,N_24842);
and UO_1737 (O_1737,N_24891,N_24995);
or UO_1738 (O_1738,N_24834,N_24995);
or UO_1739 (O_1739,N_24824,N_24924);
xnor UO_1740 (O_1740,N_24769,N_24859);
nor UO_1741 (O_1741,N_24995,N_24922);
and UO_1742 (O_1742,N_24756,N_24931);
or UO_1743 (O_1743,N_24847,N_24803);
or UO_1744 (O_1744,N_24855,N_24886);
nor UO_1745 (O_1745,N_24936,N_24890);
xor UO_1746 (O_1746,N_24780,N_24927);
or UO_1747 (O_1747,N_24887,N_24965);
nand UO_1748 (O_1748,N_24957,N_24959);
nor UO_1749 (O_1749,N_24993,N_24950);
or UO_1750 (O_1750,N_24923,N_24856);
or UO_1751 (O_1751,N_24872,N_24938);
or UO_1752 (O_1752,N_24846,N_24928);
or UO_1753 (O_1753,N_24868,N_24936);
and UO_1754 (O_1754,N_24889,N_24814);
nand UO_1755 (O_1755,N_24893,N_24796);
nor UO_1756 (O_1756,N_24866,N_24755);
nor UO_1757 (O_1757,N_24850,N_24903);
nand UO_1758 (O_1758,N_24880,N_24867);
nor UO_1759 (O_1759,N_24871,N_24813);
nor UO_1760 (O_1760,N_24888,N_24963);
xor UO_1761 (O_1761,N_24958,N_24776);
nand UO_1762 (O_1762,N_24903,N_24995);
or UO_1763 (O_1763,N_24966,N_24978);
nor UO_1764 (O_1764,N_24892,N_24978);
nor UO_1765 (O_1765,N_24870,N_24948);
xnor UO_1766 (O_1766,N_24933,N_24855);
xor UO_1767 (O_1767,N_24982,N_24930);
or UO_1768 (O_1768,N_24937,N_24957);
and UO_1769 (O_1769,N_24967,N_24794);
or UO_1770 (O_1770,N_24832,N_24923);
nor UO_1771 (O_1771,N_24817,N_24852);
nand UO_1772 (O_1772,N_24976,N_24938);
xor UO_1773 (O_1773,N_24870,N_24769);
nor UO_1774 (O_1774,N_24884,N_24898);
xnor UO_1775 (O_1775,N_24825,N_24948);
or UO_1776 (O_1776,N_24913,N_24767);
or UO_1777 (O_1777,N_24761,N_24912);
xnor UO_1778 (O_1778,N_24762,N_24939);
xor UO_1779 (O_1779,N_24870,N_24796);
xor UO_1780 (O_1780,N_24992,N_24911);
and UO_1781 (O_1781,N_24975,N_24876);
or UO_1782 (O_1782,N_24862,N_24965);
nor UO_1783 (O_1783,N_24989,N_24855);
or UO_1784 (O_1784,N_24916,N_24999);
or UO_1785 (O_1785,N_24771,N_24887);
nor UO_1786 (O_1786,N_24757,N_24982);
nor UO_1787 (O_1787,N_24978,N_24843);
xnor UO_1788 (O_1788,N_24789,N_24794);
or UO_1789 (O_1789,N_24775,N_24978);
nor UO_1790 (O_1790,N_24986,N_24874);
and UO_1791 (O_1791,N_24899,N_24932);
xor UO_1792 (O_1792,N_24753,N_24981);
xor UO_1793 (O_1793,N_24952,N_24872);
xor UO_1794 (O_1794,N_24787,N_24855);
xor UO_1795 (O_1795,N_24910,N_24912);
nand UO_1796 (O_1796,N_24904,N_24936);
and UO_1797 (O_1797,N_24974,N_24861);
and UO_1798 (O_1798,N_24928,N_24977);
nor UO_1799 (O_1799,N_24954,N_24755);
or UO_1800 (O_1800,N_24956,N_24902);
and UO_1801 (O_1801,N_24849,N_24851);
nand UO_1802 (O_1802,N_24860,N_24752);
xor UO_1803 (O_1803,N_24994,N_24859);
and UO_1804 (O_1804,N_24918,N_24960);
xnor UO_1805 (O_1805,N_24878,N_24758);
xor UO_1806 (O_1806,N_24853,N_24858);
nor UO_1807 (O_1807,N_24842,N_24954);
nor UO_1808 (O_1808,N_24815,N_24934);
xor UO_1809 (O_1809,N_24842,N_24927);
or UO_1810 (O_1810,N_24891,N_24958);
and UO_1811 (O_1811,N_24923,N_24932);
xor UO_1812 (O_1812,N_24862,N_24932);
nand UO_1813 (O_1813,N_24977,N_24898);
xnor UO_1814 (O_1814,N_24849,N_24925);
nor UO_1815 (O_1815,N_24920,N_24996);
or UO_1816 (O_1816,N_24996,N_24806);
or UO_1817 (O_1817,N_24866,N_24780);
xor UO_1818 (O_1818,N_24766,N_24844);
nand UO_1819 (O_1819,N_24790,N_24992);
nand UO_1820 (O_1820,N_24932,N_24901);
xnor UO_1821 (O_1821,N_24763,N_24937);
nand UO_1822 (O_1822,N_24998,N_24999);
and UO_1823 (O_1823,N_24781,N_24991);
nor UO_1824 (O_1824,N_24893,N_24924);
nor UO_1825 (O_1825,N_24848,N_24872);
nor UO_1826 (O_1826,N_24770,N_24774);
or UO_1827 (O_1827,N_24818,N_24823);
and UO_1828 (O_1828,N_24945,N_24775);
and UO_1829 (O_1829,N_24883,N_24795);
or UO_1830 (O_1830,N_24751,N_24921);
xor UO_1831 (O_1831,N_24823,N_24854);
and UO_1832 (O_1832,N_24979,N_24794);
nor UO_1833 (O_1833,N_24963,N_24867);
or UO_1834 (O_1834,N_24780,N_24898);
nand UO_1835 (O_1835,N_24889,N_24887);
nand UO_1836 (O_1836,N_24856,N_24956);
and UO_1837 (O_1837,N_24784,N_24982);
or UO_1838 (O_1838,N_24999,N_24791);
or UO_1839 (O_1839,N_24945,N_24989);
or UO_1840 (O_1840,N_24835,N_24798);
nor UO_1841 (O_1841,N_24759,N_24880);
nand UO_1842 (O_1842,N_24971,N_24798);
and UO_1843 (O_1843,N_24864,N_24805);
xor UO_1844 (O_1844,N_24933,N_24974);
nand UO_1845 (O_1845,N_24969,N_24825);
xnor UO_1846 (O_1846,N_24904,N_24764);
and UO_1847 (O_1847,N_24962,N_24964);
and UO_1848 (O_1848,N_24798,N_24867);
xor UO_1849 (O_1849,N_24959,N_24785);
and UO_1850 (O_1850,N_24937,N_24801);
and UO_1851 (O_1851,N_24964,N_24817);
and UO_1852 (O_1852,N_24989,N_24851);
xor UO_1853 (O_1853,N_24842,N_24882);
xnor UO_1854 (O_1854,N_24824,N_24997);
nand UO_1855 (O_1855,N_24827,N_24797);
nor UO_1856 (O_1856,N_24969,N_24858);
and UO_1857 (O_1857,N_24797,N_24864);
or UO_1858 (O_1858,N_24887,N_24891);
and UO_1859 (O_1859,N_24925,N_24873);
xnor UO_1860 (O_1860,N_24847,N_24956);
xor UO_1861 (O_1861,N_24949,N_24839);
nor UO_1862 (O_1862,N_24874,N_24863);
xnor UO_1863 (O_1863,N_24966,N_24959);
xor UO_1864 (O_1864,N_24876,N_24814);
nand UO_1865 (O_1865,N_24913,N_24948);
nand UO_1866 (O_1866,N_24893,N_24972);
or UO_1867 (O_1867,N_24871,N_24999);
nand UO_1868 (O_1868,N_24983,N_24990);
or UO_1869 (O_1869,N_24969,N_24883);
nor UO_1870 (O_1870,N_24911,N_24855);
nor UO_1871 (O_1871,N_24835,N_24750);
nor UO_1872 (O_1872,N_24931,N_24794);
nor UO_1873 (O_1873,N_24887,N_24760);
and UO_1874 (O_1874,N_24934,N_24900);
nand UO_1875 (O_1875,N_24903,N_24880);
or UO_1876 (O_1876,N_24900,N_24952);
xor UO_1877 (O_1877,N_24845,N_24991);
xnor UO_1878 (O_1878,N_24958,N_24842);
nand UO_1879 (O_1879,N_24804,N_24896);
or UO_1880 (O_1880,N_24882,N_24998);
xnor UO_1881 (O_1881,N_24869,N_24938);
nor UO_1882 (O_1882,N_24991,N_24869);
and UO_1883 (O_1883,N_24870,N_24808);
or UO_1884 (O_1884,N_24755,N_24993);
nand UO_1885 (O_1885,N_24834,N_24756);
xnor UO_1886 (O_1886,N_24862,N_24958);
nor UO_1887 (O_1887,N_24771,N_24881);
and UO_1888 (O_1888,N_24859,N_24853);
or UO_1889 (O_1889,N_24773,N_24948);
and UO_1890 (O_1890,N_24965,N_24973);
or UO_1891 (O_1891,N_24983,N_24863);
nand UO_1892 (O_1892,N_24889,N_24770);
or UO_1893 (O_1893,N_24750,N_24876);
nand UO_1894 (O_1894,N_24929,N_24760);
and UO_1895 (O_1895,N_24782,N_24854);
nand UO_1896 (O_1896,N_24954,N_24909);
xnor UO_1897 (O_1897,N_24785,N_24759);
nor UO_1898 (O_1898,N_24754,N_24822);
or UO_1899 (O_1899,N_24980,N_24776);
xor UO_1900 (O_1900,N_24820,N_24781);
xnor UO_1901 (O_1901,N_24952,N_24989);
or UO_1902 (O_1902,N_24831,N_24924);
or UO_1903 (O_1903,N_24992,N_24829);
nand UO_1904 (O_1904,N_24935,N_24892);
or UO_1905 (O_1905,N_24916,N_24929);
and UO_1906 (O_1906,N_24946,N_24939);
and UO_1907 (O_1907,N_24840,N_24886);
nand UO_1908 (O_1908,N_24870,N_24907);
xnor UO_1909 (O_1909,N_24803,N_24907);
xnor UO_1910 (O_1910,N_24784,N_24844);
nand UO_1911 (O_1911,N_24962,N_24877);
xnor UO_1912 (O_1912,N_24824,N_24869);
xor UO_1913 (O_1913,N_24766,N_24762);
nand UO_1914 (O_1914,N_24790,N_24939);
or UO_1915 (O_1915,N_24885,N_24973);
nor UO_1916 (O_1916,N_24839,N_24770);
or UO_1917 (O_1917,N_24978,N_24893);
or UO_1918 (O_1918,N_24931,N_24971);
and UO_1919 (O_1919,N_24895,N_24753);
xnor UO_1920 (O_1920,N_24771,N_24898);
nor UO_1921 (O_1921,N_24780,N_24953);
xnor UO_1922 (O_1922,N_24924,N_24881);
xnor UO_1923 (O_1923,N_24999,N_24978);
nor UO_1924 (O_1924,N_24799,N_24946);
and UO_1925 (O_1925,N_24879,N_24925);
and UO_1926 (O_1926,N_24838,N_24979);
or UO_1927 (O_1927,N_24793,N_24926);
nor UO_1928 (O_1928,N_24997,N_24836);
xnor UO_1929 (O_1929,N_24844,N_24943);
or UO_1930 (O_1930,N_24891,N_24836);
and UO_1931 (O_1931,N_24860,N_24958);
or UO_1932 (O_1932,N_24944,N_24943);
or UO_1933 (O_1933,N_24828,N_24936);
or UO_1934 (O_1934,N_24887,N_24866);
nor UO_1935 (O_1935,N_24770,N_24791);
or UO_1936 (O_1936,N_24779,N_24866);
nand UO_1937 (O_1937,N_24931,N_24836);
nand UO_1938 (O_1938,N_24902,N_24782);
or UO_1939 (O_1939,N_24954,N_24797);
nor UO_1940 (O_1940,N_24794,N_24784);
nand UO_1941 (O_1941,N_24934,N_24915);
nor UO_1942 (O_1942,N_24783,N_24937);
or UO_1943 (O_1943,N_24823,N_24959);
or UO_1944 (O_1944,N_24770,N_24931);
nor UO_1945 (O_1945,N_24801,N_24767);
and UO_1946 (O_1946,N_24944,N_24913);
xnor UO_1947 (O_1947,N_24938,N_24909);
xor UO_1948 (O_1948,N_24863,N_24968);
and UO_1949 (O_1949,N_24934,N_24841);
xor UO_1950 (O_1950,N_24804,N_24774);
nand UO_1951 (O_1951,N_24871,N_24924);
xnor UO_1952 (O_1952,N_24927,N_24885);
and UO_1953 (O_1953,N_24854,N_24984);
nor UO_1954 (O_1954,N_24956,N_24864);
nand UO_1955 (O_1955,N_24807,N_24789);
xnor UO_1956 (O_1956,N_24896,N_24914);
or UO_1957 (O_1957,N_24866,N_24843);
nand UO_1958 (O_1958,N_24953,N_24798);
and UO_1959 (O_1959,N_24997,N_24880);
nor UO_1960 (O_1960,N_24851,N_24981);
and UO_1961 (O_1961,N_24993,N_24982);
nor UO_1962 (O_1962,N_24863,N_24778);
xnor UO_1963 (O_1963,N_24933,N_24835);
xor UO_1964 (O_1964,N_24757,N_24810);
and UO_1965 (O_1965,N_24926,N_24907);
or UO_1966 (O_1966,N_24950,N_24754);
xor UO_1967 (O_1967,N_24837,N_24877);
or UO_1968 (O_1968,N_24860,N_24922);
nor UO_1969 (O_1969,N_24809,N_24895);
nand UO_1970 (O_1970,N_24911,N_24952);
or UO_1971 (O_1971,N_24993,N_24792);
xnor UO_1972 (O_1972,N_24955,N_24764);
or UO_1973 (O_1973,N_24817,N_24976);
xnor UO_1974 (O_1974,N_24832,N_24768);
nor UO_1975 (O_1975,N_24821,N_24880);
and UO_1976 (O_1976,N_24902,N_24869);
and UO_1977 (O_1977,N_24882,N_24846);
nor UO_1978 (O_1978,N_24799,N_24994);
nand UO_1979 (O_1979,N_24924,N_24815);
or UO_1980 (O_1980,N_24977,N_24982);
and UO_1981 (O_1981,N_24794,N_24936);
xnor UO_1982 (O_1982,N_24776,N_24917);
or UO_1983 (O_1983,N_24822,N_24862);
xor UO_1984 (O_1984,N_24799,N_24775);
xor UO_1985 (O_1985,N_24998,N_24978);
xor UO_1986 (O_1986,N_24751,N_24845);
nor UO_1987 (O_1987,N_24980,N_24929);
nor UO_1988 (O_1988,N_24768,N_24921);
or UO_1989 (O_1989,N_24758,N_24809);
xnor UO_1990 (O_1990,N_24980,N_24927);
xnor UO_1991 (O_1991,N_24940,N_24987);
xor UO_1992 (O_1992,N_24770,N_24786);
and UO_1993 (O_1993,N_24768,N_24864);
and UO_1994 (O_1994,N_24964,N_24975);
xnor UO_1995 (O_1995,N_24762,N_24819);
xor UO_1996 (O_1996,N_24941,N_24963);
and UO_1997 (O_1997,N_24934,N_24958);
nand UO_1998 (O_1998,N_24792,N_24991);
and UO_1999 (O_1999,N_24984,N_24872);
or UO_2000 (O_2000,N_24990,N_24762);
nand UO_2001 (O_2001,N_24940,N_24890);
nor UO_2002 (O_2002,N_24839,N_24777);
or UO_2003 (O_2003,N_24926,N_24860);
nor UO_2004 (O_2004,N_24952,N_24754);
xnor UO_2005 (O_2005,N_24868,N_24841);
xor UO_2006 (O_2006,N_24946,N_24817);
nand UO_2007 (O_2007,N_24766,N_24924);
nor UO_2008 (O_2008,N_24787,N_24903);
nor UO_2009 (O_2009,N_24985,N_24819);
nor UO_2010 (O_2010,N_24949,N_24964);
nand UO_2011 (O_2011,N_24998,N_24982);
or UO_2012 (O_2012,N_24979,N_24836);
and UO_2013 (O_2013,N_24910,N_24868);
nor UO_2014 (O_2014,N_24873,N_24863);
or UO_2015 (O_2015,N_24803,N_24810);
and UO_2016 (O_2016,N_24870,N_24804);
nor UO_2017 (O_2017,N_24846,N_24832);
nand UO_2018 (O_2018,N_24820,N_24872);
and UO_2019 (O_2019,N_24954,N_24922);
nand UO_2020 (O_2020,N_24761,N_24805);
nand UO_2021 (O_2021,N_24810,N_24836);
nor UO_2022 (O_2022,N_24912,N_24874);
nand UO_2023 (O_2023,N_24779,N_24977);
xnor UO_2024 (O_2024,N_24994,N_24981);
and UO_2025 (O_2025,N_24825,N_24967);
nor UO_2026 (O_2026,N_24750,N_24859);
nor UO_2027 (O_2027,N_24991,N_24844);
or UO_2028 (O_2028,N_24860,N_24876);
and UO_2029 (O_2029,N_24761,N_24870);
and UO_2030 (O_2030,N_24755,N_24896);
and UO_2031 (O_2031,N_24762,N_24861);
xor UO_2032 (O_2032,N_24991,N_24959);
and UO_2033 (O_2033,N_24805,N_24908);
xor UO_2034 (O_2034,N_24823,N_24814);
nand UO_2035 (O_2035,N_24885,N_24841);
xnor UO_2036 (O_2036,N_24900,N_24801);
nand UO_2037 (O_2037,N_24961,N_24787);
nor UO_2038 (O_2038,N_24777,N_24816);
nor UO_2039 (O_2039,N_24801,N_24847);
xor UO_2040 (O_2040,N_24816,N_24881);
xor UO_2041 (O_2041,N_24990,N_24877);
and UO_2042 (O_2042,N_24990,N_24878);
nor UO_2043 (O_2043,N_24891,N_24905);
xnor UO_2044 (O_2044,N_24973,N_24952);
and UO_2045 (O_2045,N_24970,N_24992);
xnor UO_2046 (O_2046,N_24927,N_24904);
nand UO_2047 (O_2047,N_24878,N_24943);
nor UO_2048 (O_2048,N_24810,N_24815);
and UO_2049 (O_2049,N_24795,N_24870);
nand UO_2050 (O_2050,N_24967,N_24767);
or UO_2051 (O_2051,N_24873,N_24752);
nor UO_2052 (O_2052,N_24925,N_24963);
xor UO_2053 (O_2053,N_24968,N_24869);
xor UO_2054 (O_2054,N_24835,N_24890);
nor UO_2055 (O_2055,N_24783,N_24757);
xor UO_2056 (O_2056,N_24967,N_24822);
or UO_2057 (O_2057,N_24781,N_24756);
and UO_2058 (O_2058,N_24762,N_24802);
nor UO_2059 (O_2059,N_24987,N_24786);
nand UO_2060 (O_2060,N_24760,N_24849);
nor UO_2061 (O_2061,N_24803,N_24850);
and UO_2062 (O_2062,N_24784,N_24765);
nor UO_2063 (O_2063,N_24788,N_24792);
xor UO_2064 (O_2064,N_24845,N_24906);
xor UO_2065 (O_2065,N_24798,N_24839);
and UO_2066 (O_2066,N_24917,N_24878);
nor UO_2067 (O_2067,N_24751,N_24872);
nand UO_2068 (O_2068,N_24778,N_24842);
and UO_2069 (O_2069,N_24937,N_24897);
or UO_2070 (O_2070,N_24839,N_24917);
or UO_2071 (O_2071,N_24757,N_24803);
nand UO_2072 (O_2072,N_24783,N_24936);
xor UO_2073 (O_2073,N_24964,N_24942);
or UO_2074 (O_2074,N_24947,N_24859);
or UO_2075 (O_2075,N_24778,N_24777);
nand UO_2076 (O_2076,N_24880,N_24850);
xor UO_2077 (O_2077,N_24805,N_24979);
xnor UO_2078 (O_2078,N_24885,N_24982);
and UO_2079 (O_2079,N_24976,N_24819);
or UO_2080 (O_2080,N_24757,N_24767);
or UO_2081 (O_2081,N_24990,N_24908);
and UO_2082 (O_2082,N_24897,N_24984);
and UO_2083 (O_2083,N_24952,N_24876);
or UO_2084 (O_2084,N_24803,N_24939);
and UO_2085 (O_2085,N_24763,N_24995);
or UO_2086 (O_2086,N_24836,N_24855);
xor UO_2087 (O_2087,N_24981,N_24871);
or UO_2088 (O_2088,N_24778,N_24948);
xnor UO_2089 (O_2089,N_24994,N_24757);
nor UO_2090 (O_2090,N_24943,N_24769);
nor UO_2091 (O_2091,N_24845,N_24908);
xor UO_2092 (O_2092,N_24995,N_24898);
nor UO_2093 (O_2093,N_24926,N_24959);
and UO_2094 (O_2094,N_24923,N_24895);
nor UO_2095 (O_2095,N_24836,N_24814);
nor UO_2096 (O_2096,N_24756,N_24892);
or UO_2097 (O_2097,N_24971,N_24855);
nand UO_2098 (O_2098,N_24802,N_24958);
or UO_2099 (O_2099,N_24941,N_24905);
nor UO_2100 (O_2100,N_24869,N_24856);
xnor UO_2101 (O_2101,N_24896,N_24998);
nand UO_2102 (O_2102,N_24945,N_24815);
or UO_2103 (O_2103,N_24823,N_24833);
or UO_2104 (O_2104,N_24887,N_24876);
nand UO_2105 (O_2105,N_24752,N_24782);
and UO_2106 (O_2106,N_24948,N_24810);
nand UO_2107 (O_2107,N_24770,N_24960);
and UO_2108 (O_2108,N_24951,N_24823);
and UO_2109 (O_2109,N_24806,N_24888);
or UO_2110 (O_2110,N_24917,N_24959);
xnor UO_2111 (O_2111,N_24926,N_24916);
and UO_2112 (O_2112,N_24955,N_24798);
xor UO_2113 (O_2113,N_24840,N_24779);
nand UO_2114 (O_2114,N_24828,N_24854);
and UO_2115 (O_2115,N_24955,N_24759);
and UO_2116 (O_2116,N_24880,N_24984);
or UO_2117 (O_2117,N_24932,N_24758);
and UO_2118 (O_2118,N_24859,N_24987);
nand UO_2119 (O_2119,N_24979,N_24964);
nand UO_2120 (O_2120,N_24974,N_24863);
nor UO_2121 (O_2121,N_24822,N_24766);
nor UO_2122 (O_2122,N_24995,N_24954);
nand UO_2123 (O_2123,N_24835,N_24916);
and UO_2124 (O_2124,N_24990,N_24973);
xnor UO_2125 (O_2125,N_24908,N_24942);
xor UO_2126 (O_2126,N_24828,N_24934);
nand UO_2127 (O_2127,N_24765,N_24968);
nor UO_2128 (O_2128,N_24792,N_24943);
or UO_2129 (O_2129,N_24984,N_24983);
and UO_2130 (O_2130,N_24854,N_24966);
and UO_2131 (O_2131,N_24856,N_24832);
nor UO_2132 (O_2132,N_24802,N_24852);
nor UO_2133 (O_2133,N_24842,N_24779);
xnor UO_2134 (O_2134,N_24853,N_24819);
and UO_2135 (O_2135,N_24960,N_24757);
xnor UO_2136 (O_2136,N_24813,N_24862);
xor UO_2137 (O_2137,N_24751,N_24999);
nand UO_2138 (O_2138,N_24782,N_24918);
and UO_2139 (O_2139,N_24964,N_24852);
and UO_2140 (O_2140,N_24822,N_24790);
or UO_2141 (O_2141,N_24806,N_24957);
or UO_2142 (O_2142,N_24933,N_24871);
and UO_2143 (O_2143,N_24856,N_24965);
xnor UO_2144 (O_2144,N_24876,N_24904);
or UO_2145 (O_2145,N_24950,N_24903);
or UO_2146 (O_2146,N_24838,N_24758);
nand UO_2147 (O_2147,N_24979,N_24753);
nand UO_2148 (O_2148,N_24838,N_24917);
nor UO_2149 (O_2149,N_24910,N_24862);
nand UO_2150 (O_2150,N_24988,N_24962);
nor UO_2151 (O_2151,N_24755,N_24885);
nor UO_2152 (O_2152,N_24767,N_24798);
nand UO_2153 (O_2153,N_24875,N_24996);
and UO_2154 (O_2154,N_24753,N_24962);
and UO_2155 (O_2155,N_24876,N_24954);
or UO_2156 (O_2156,N_24856,N_24795);
nor UO_2157 (O_2157,N_24854,N_24907);
or UO_2158 (O_2158,N_24941,N_24791);
xnor UO_2159 (O_2159,N_24917,N_24826);
or UO_2160 (O_2160,N_24864,N_24755);
nor UO_2161 (O_2161,N_24926,N_24968);
nor UO_2162 (O_2162,N_24772,N_24981);
or UO_2163 (O_2163,N_24978,N_24795);
nor UO_2164 (O_2164,N_24936,N_24805);
xnor UO_2165 (O_2165,N_24942,N_24833);
nor UO_2166 (O_2166,N_24789,N_24942);
or UO_2167 (O_2167,N_24843,N_24889);
nand UO_2168 (O_2168,N_24871,N_24967);
nand UO_2169 (O_2169,N_24905,N_24837);
nor UO_2170 (O_2170,N_24820,N_24955);
nand UO_2171 (O_2171,N_24815,N_24781);
and UO_2172 (O_2172,N_24856,N_24840);
nand UO_2173 (O_2173,N_24869,N_24782);
nand UO_2174 (O_2174,N_24930,N_24845);
nor UO_2175 (O_2175,N_24825,N_24943);
nor UO_2176 (O_2176,N_24806,N_24919);
nand UO_2177 (O_2177,N_24855,N_24977);
or UO_2178 (O_2178,N_24786,N_24937);
xnor UO_2179 (O_2179,N_24780,N_24834);
or UO_2180 (O_2180,N_24890,N_24924);
xor UO_2181 (O_2181,N_24801,N_24759);
or UO_2182 (O_2182,N_24936,N_24798);
or UO_2183 (O_2183,N_24806,N_24763);
nand UO_2184 (O_2184,N_24958,N_24965);
nor UO_2185 (O_2185,N_24888,N_24973);
and UO_2186 (O_2186,N_24759,N_24810);
nor UO_2187 (O_2187,N_24877,N_24883);
or UO_2188 (O_2188,N_24801,N_24779);
nor UO_2189 (O_2189,N_24980,N_24833);
or UO_2190 (O_2190,N_24976,N_24948);
nor UO_2191 (O_2191,N_24871,N_24906);
nor UO_2192 (O_2192,N_24820,N_24911);
or UO_2193 (O_2193,N_24877,N_24795);
or UO_2194 (O_2194,N_24968,N_24874);
xor UO_2195 (O_2195,N_24804,N_24987);
or UO_2196 (O_2196,N_24779,N_24871);
nor UO_2197 (O_2197,N_24907,N_24818);
or UO_2198 (O_2198,N_24765,N_24785);
nor UO_2199 (O_2199,N_24770,N_24964);
and UO_2200 (O_2200,N_24887,N_24789);
xnor UO_2201 (O_2201,N_24984,N_24851);
xnor UO_2202 (O_2202,N_24950,N_24874);
xor UO_2203 (O_2203,N_24897,N_24966);
nand UO_2204 (O_2204,N_24867,N_24961);
nand UO_2205 (O_2205,N_24763,N_24851);
nor UO_2206 (O_2206,N_24824,N_24809);
nor UO_2207 (O_2207,N_24933,N_24946);
or UO_2208 (O_2208,N_24826,N_24761);
nand UO_2209 (O_2209,N_24856,N_24878);
nor UO_2210 (O_2210,N_24899,N_24923);
xor UO_2211 (O_2211,N_24817,N_24939);
or UO_2212 (O_2212,N_24929,N_24766);
and UO_2213 (O_2213,N_24981,N_24985);
and UO_2214 (O_2214,N_24980,N_24858);
xor UO_2215 (O_2215,N_24784,N_24936);
nor UO_2216 (O_2216,N_24787,N_24806);
nor UO_2217 (O_2217,N_24758,N_24800);
xor UO_2218 (O_2218,N_24987,N_24901);
and UO_2219 (O_2219,N_24880,N_24786);
and UO_2220 (O_2220,N_24899,N_24931);
nor UO_2221 (O_2221,N_24933,N_24890);
nand UO_2222 (O_2222,N_24971,N_24883);
nand UO_2223 (O_2223,N_24927,N_24907);
and UO_2224 (O_2224,N_24896,N_24851);
and UO_2225 (O_2225,N_24840,N_24760);
nor UO_2226 (O_2226,N_24882,N_24790);
and UO_2227 (O_2227,N_24849,N_24750);
and UO_2228 (O_2228,N_24837,N_24824);
and UO_2229 (O_2229,N_24768,N_24900);
or UO_2230 (O_2230,N_24769,N_24775);
and UO_2231 (O_2231,N_24776,N_24911);
nor UO_2232 (O_2232,N_24818,N_24913);
and UO_2233 (O_2233,N_24933,N_24842);
nor UO_2234 (O_2234,N_24914,N_24956);
and UO_2235 (O_2235,N_24908,N_24761);
nor UO_2236 (O_2236,N_24906,N_24935);
nor UO_2237 (O_2237,N_24847,N_24951);
nand UO_2238 (O_2238,N_24899,N_24939);
xnor UO_2239 (O_2239,N_24780,N_24821);
and UO_2240 (O_2240,N_24816,N_24904);
nor UO_2241 (O_2241,N_24984,N_24926);
nand UO_2242 (O_2242,N_24890,N_24840);
xor UO_2243 (O_2243,N_24759,N_24861);
nor UO_2244 (O_2244,N_24780,N_24941);
nand UO_2245 (O_2245,N_24962,N_24994);
or UO_2246 (O_2246,N_24962,N_24915);
or UO_2247 (O_2247,N_24835,N_24854);
or UO_2248 (O_2248,N_24763,N_24951);
nor UO_2249 (O_2249,N_24910,N_24861);
nand UO_2250 (O_2250,N_24919,N_24793);
and UO_2251 (O_2251,N_24956,N_24795);
xnor UO_2252 (O_2252,N_24759,N_24979);
xnor UO_2253 (O_2253,N_24905,N_24841);
xor UO_2254 (O_2254,N_24769,N_24890);
nor UO_2255 (O_2255,N_24781,N_24829);
nor UO_2256 (O_2256,N_24877,N_24849);
nand UO_2257 (O_2257,N_24785,N_24892);
or UO_2258 (O_2258,N_24795,N_24819);
xor UO_2259 (O_2259,N_24825,N_24876);
nor UO_2260 (O_2260,N_24871,N_24985);
xnor UO_2261 (O_2261,N_24814,N_24846);
nand UO_2262 (O_2262,N_24821,N_24776);
and UO_2263 (O_2263,N_24883,N_24933);
nand UO_2264 (O_2264,N_24906,N_24802);
nand UO_2265 (O_2265,N_24966,N_24784);
or UO_2266 (O_2266,N_24984,N_24790);
nor UO_2267 (O_2267,N_24823,N_24821);
or UO_2268 (O_2268,N_24957,N_24813);
nor UO_2269 (O_2269,N_24842,N_24759);
nor UO_2270 (O_2270,N_24785,N_24870);
and UO_2271 (O_2271,N_24829,N_24876);
nand UO_2272 (O_2272,N_24837,N_24937);
nand UO_2273 (O_2273,N_24869,N_24970);
nand UO_2274 (O_2274,N_24786,N_24806);
and UO_2275 (O_2275,N_24835,N_24983);
and UO_2276 (O_2276,N_24810,N_24881);
or UO_2277 (O_2277,N_24887,N_24855);
xor UO_2278 (O_2278,N_24908,N_24816);
nor UO_2279 (O_2279,N_24819,N_24863);
or UO_2280 (O_2280,N_24943,N_24882);
nand UO_2281 (O_2281,N_24853,N_24993);
or UO_2282 (O_2282,N_24877,N_24964);
or UO_2283 (O_2283,N_24784,N_24891);
nor UO_2284 (O_2284,N_24889,N_24829);
and UO_2285 (O_2285,N_24860,N_24795);
or UO_2286 (O_2286,N_24926,N_24872);
nand UO_2287 (O_2287,N_24793,N_24892);
or UO_2288 (O_2288,N_24783,N_24811);
and UO_2289 (O_2289,N_24982,N_24801);
xnor UO_2290 (O_2290,N_24909,N_24877);
nor UO_2291 (O_2291,N_24830,N_24866);
xor UO_2292 (O_2292,N_24839,N_24811);
or UO_2293 (O_2293,N_24830,N_24769);
xnor UO_2294 (O_2294,N_24802,N_24817);
and UO_2295 (O_2295,N_24970,N_24847);
or UO_2296 (O_2296,N_24980,N_24978);
and UO_2297 (O_2297,N_24778,N_24924);
nand UO_2298 (O_2298,N_24819,N_24754);
or UO_2299 (O_2299,N_24784,N_24860);
nand UO_2300 (O_2300,N_24851,N_24816);
nor UO_2301 (O_2301,N_24844,N_24882);
and UO_2302 (O_2302,N_24903,N_24851);
or UO_2303 (O_2303,N_24989,N_24769);
nand UO_2304 (O_2304,N_24859,N_24832);
or UO_2305 (O_2305,N_24774,N_24866);
and UO_2306 (O_2306,N_24831,N_24816);
nor UO_2307 (O_2307,N_24911,N_24953);
or UO_2308 (O_2308,N_24966,N_24757);
xor UO_2309 (O_2309,N_24818,N_24751);
and UO_2310 (O_2310,N_24925,N_24821);
nand UO_2311 (O_2311,N_24932,N_24950);
and UO_2312 (O_2312,N_24883,N_24862);
xor UO_2313 (O_2313,N_24816,N_24767);
or UO_2314 (O_2314,N_24778,N_24963);
nand UO_2315 (O_2315,N_24887,N_24882);
nand UO_2316 (O_2316,N_24897,N_24864);
nor UO_2317 (O_2317,N_24867,N_24899);
xnor UO_2318 (O_2318,N_24838,N_24787);
or UO_2319 (O_2319,N_24754,N_24800);
and UO_2320 (O_2320,N_24992,N_24936);
nor UO_2321 (O_2321,N_24887,N_24787);
nand UO_2322 (O_2322,N_24803,N_24763);
nand UO_2323 (O_2323,N_24801,N_24938);
or UO_2324 (O_2324,N_24803,N_24773);
or UO_2325 (O_2325,N_24978,N_24796);
nor UO_2326 (O_2326,N_24817,N_24913);
nand UO_2327 (O_2327,N_24919,N_24769);
and UO_2328 (O_2328,N_24904,N_24755);
and UO_2329 (O_2329,N_24846,N_24804);
and UO_2330 (O_2330,N_24850,N_24878);
and UO_2331 (O_2331,N_24834,N_24845);
nor UO_2332 (O_2332,N_24771,N_24961);
or UO_2333 (O_2333,N_24841,N_24893);
nor UO_2334 (O_2334,N_24799,N_24922);
and UO_2335 (O_2335,N_24766,N_24860);
nand UO_2336 (O_2336,N_24948,N_24937);
or UO_2337 (O_2337,N_24901,N_24793);
and UO_2338 (O_2338,N_24960,N_24977);
xor UO_2339 (O_2339,N_24833,N_24971);
xor UO_2340 (O_2340,N_24937,N_24967);
and UO_2341 (O_2341,N_24927,N_24945);
nand UO_2342 (O_2342,N_24912,N_24883);
xor UO_2343 (O_2343,N_24790,N_24901);
or UO_2344 (O_2344,N_24832,N_24770);
xor UO_2345 (O_2345,N_24956,N_24769);
and UO_2346 (O_2346,N_24912,N_24820);
and UO_2347 (O_2347,N_24939,N_24834);
xor UO_2348 (O_2348,N_24822,N_24915);
and UO_2349 (O_2349,N_24952,N_24773);
or UO_2350 (O_2350,N_24993,N_24830);
or UO_2351 (O_2351,N_24859,N_24920);
or UO_2352 (O_2352,N_24951,N_24830);
or UO_2353 (O_2353,N_24898,N_24943);
xor UO_2354 (O_2354,N_24786,N_24849);
xnor UO_2355 (O_2355,N_24911,N_24966);
or UO_2356 (O_2356,N_24898,N_24970);
or UO_2357 (O_2357,N_24875,N_24860);
nand UO_2358 (O_2358,N_24757,N_24916);
or UO_2359 (O_2359,N_24815,N_24794);
nand UO_2360 (O_2360,N_24768,N_24983);
nand UO_2361 (O_2361,N_24814,N_24852);
nor UO_2362 (O_2362,N_24840,N_24827);
nand UO_2363 (O_2363,N_24883,N_24847);
nor UO_2364 (O_2364,N_24868,N_24941);
nor UO_2365 (O_2365,N_24779,N_24950);
nand UO_2366 (O_2366,N_24889,N_24861);
nand UO_2367 (O_2367,N_24878,N_24956);
nor UO_2368 (O_2368,N_24843,N_24968);
nand UO_2369 (O_2369,N_24818,N_24999);
or UO_2370 (O_2370,N_24808,N_24784);
or UO_2371 (O_2371,N_24972,N_24753);
and UO_2372 (O_2372,N_24996,N_24958);
or UO_2373 (O_2373,N_24836,N_24786);
and UO_2374 (O_2374,N_24750,N_24927);
nor UO_2375 (O_2375,N_24838,N_24775);
or UO_2376 (O_2376,N_24880,N_24942);
nand UO_2377 (O_2377,N_24982,N_24763);
or UO_2378 (O_2378,N_24994,N_24814);
xor UO_2379 (O_2379,N_24899,N_24984);
and UO_2380 (O_2380,N_24792,N_24868);
or UO_2381 (O_2381,N_24969,N_24807);
or UO_2382 (O_2382,N_24759,N_24998);
or UO_2383 (O_2383,N_24793,N_24998);
and UO_2384 (O_2384,N_24819,N_24982);
or UO_2385 (O_2385,N_24981,N_24938);
and UO_2386 (O_2386,N_24851,N_24966);
nand UO_2387 (O_2387,N_24764,N_24944);
or UO_2388 (O_2388,N_24816,N_24847);
xor UO_2389 (O_2389,N_24954,N_24819);
xnor UO_2390 (O_2390,N_24809,N_24804);
nor UO_2391 (O_2391,N_24967,N_24942);
and UO_2392 (O_2392,N_24790,N_24947);
or UO_2393 (O_2393,N_24886,N_24938);
nand UO_2394 (O_2394,N_24904,N_24980);
xnor UO_2395 (O_2395,N_24957,N_24918);
and UO_2396 (O_2396,N_24759,N_24807);
nand UO_2397 (O_2397,N_24836,N_24818);
nand UO_2398 (O_2398,N_24975,N_24928);
and UO_2399 (O_2399,N_24959,N_24805);
nor UO_2400 (O_2400,N_24944,N_24755);
xnor UO_2401 (O_2401,N_24934,N_24859);
nand UO_2402 (O_2402,N_24874,N_24908);
or UO_2403 (O_2403,N_24996,N_24824);
nand UO_2404 (O_2404,N_24883,N_24945);
nor UO_2405 (O_2405,N_24911,N_24991);
and UO_2406 (O_2406,N_24893,N_24909);
nor UO_2407 (O_2407,N_24937,N_24778);
and UO_2408 (O_2408,N_24761,N_24787);
nor UO_2409 (O_2409,N_24814,N_24999);
nand UO_2410 (O_2410,N_24793,N_24812);
and UO_2411 (O_2411,N_24783,N_24782);
and UO_2412 (O_2412,N_24846,N_24987);
and UO_2413 (O_2413,N_24976,N_24858);
xnor UO_2414 (O_2414,N_24786,N_24885);
nand UO_2415 (O_2415,N_24951,N_24931);
xnor UO_2416 (O_2416,N_24905,N_24912);
or UO_2417 (O_2417,N_24867,N_24758);
nor UO_2418 (O_2418,N_24812,N_24893);
and UO_2419 (O_2419,N_24834,N_24795);
and UO_2420 (O_2420,N_24966,N_24774);
and UO_2421 (O_2421,N_24810,N_24918);
and UO_2422 (O_2422,N_24767,N_24773);
or UO_2423 (O_2423,N_24858,N_24989);
and UO_2424 (O_2424,N_24838,N_24756);
xnor UO_2425 (O_2425,N_24968,N_24879);
or UO_2426 (O_2426,N_24861,N_24866);
nor UO_2427 (O_2427,N_24829,N_24809);
and UO_2428 (O_2428,N_24904,N_24765);
xor UO_2429 (O_2429,N_24790,N_24873);
nand UO_2430 (O_2430,N_24799,N_24819);
nor UO_2431 (O_2431,N_24764,N_24765);
nand UO_2432 (O_2432,N_24889,N_24866);
xor UO_2433 (O_2433,N_24787,N_24778);
or UO_2434 (O_2434,N_24827,N_24943);
xor UO_2435 (O_2435,N_24912,N_24915);
or UO_2436 (O_2436,N_24922,N_24838);
and UO_2437 (O_2437,N_24959,N_24818);
xnor UO_2438 (O_2438,N_24972,N_24797);
and UO_2439 (O_2439,N_24877,N_24968);
or UO_2440 (O_2440,N_24776,N_24805);
nand UO_2441 (O_2441,N_24831,N_24926);
or UO_2442 (O_2442,N_24927,N_24840);
nand UO_2443 (O_2443,N_24973,N_24875);
and UO_2444 (O_2444,N_24787,N_24940);
xnor UO_2445 (O_2445,N_24939,N_24935);
nor UO_2446 (O_2446,N_24980,N_24983);
or UO_2447 (O_2447,N_24994,N_24840);
nand UO_2448 (O_2448,N_24820,N_24997);
nand UO_2449 (O_2449,N_24976,N_24892);
xor UO_2450 (O_2450,N_24989,N_24905);
nor UO_2451 (O_2451,N_24952,N_24984);
nand UO_2452 (O_2452,N_24757,N_24773);
xor UO_2453 (O_2453,N_24762,N_24885);
nor UO_2454 (O_2454,N_24755,N_24858);
nor UO_2455 (O_2455,N_24774,N_24798);
nand UO_2456 (O_2456,N_24865,N_24813);
nor UO_2457 (O_2457,N_24816,N_24966);
xor UO_2458 (O_2458,N_24966,N_24981);
nand UO_2459 (O_2459,N_24761,N_24825);
nor UO_2460 (O_2460,N_24817,N_24936);
or UO_2461 (O_2461,N_24820,N_24815);
nand UO_2462 (O_2462,N_24820,N_24876);
or UO_2463 (O_2463,N_24963,N_24975);
nand UO_2464 (O_2464,N_24782,N_24977);
or UO_2465 (O_2465,N_24804,N_24854);
nand UO_2466 (O_2466,N_24843,N_24844);
nand UO_2467 (O_2467,N_24842,N_24923);
nor UO_2468 (O_2468,N_24788,N_24829);
xor UO_2469 (O_2469,N_24934,N_24911);
xnor UO_2470 (O_2470,N_24817,N_24812);
and UO_2471 (O_2471,N_24865,N_24786);
or UO_2472 (O_2472,N_24880,N_24883);
nand UO_2473 (O_2473,N_24834,N_24997);
nor UO_2474 (O_2474,N_24831,N_24977);
nand UO_2475 (O_2475,N_24843,N_24921);
and UO_2476 (O_2476,N_24918,N_24858);
or UO_2477 (O_2477,N_24993,N_24864);
or UO_2478 (O_2478,N_24997,N_24792);
or UO_2479 (O_2479,N_24890,N_24943);
xnor UO_2480 (O_2480,N_24958,N_24919);
nor UO_2481 (O_2481,N_24893,N_24818);
and UO_2482 (O_2482,N_24963,N_24899);
nor UO_2483 (O_2483,N_24800,N_24825);
nor UO_2484 (O_2484,N_24827,N_24767);
nor UO_2485 (O_2485,N_24750,N_24840);
nand UO_2486 (O_2486,N_24960,N_24927);
and UO_2487 (O_2487,N_24757,N_24785);
and UO_2488 (O_2488,N_24983,N_24882);
nand UO_2489 (O_2489,N_24901,N_24863);
xor UO_2490 (O_2490,N_24916,N_24970);
nor UO_2491 (O_2491,N_24878,N_24964);
nor UO_2492 (O_2492,N_24780,N_24979);
xor UO_2493 (O_2493,N_24938,N_24822);
or UO_2494 (O_2494,N_24956,N_24779);
xnor UO_2495 (O_2495,N_24840,N_24919);
nand UO_2496 (O_2496,N_24917,N_24941);
or UO_2497 (O_2497,N_24941,N_24851);
nor UO_2498 (O_2498,N_24804,N_24773);
nor UO_2499 (O_2499,N_24924,N_24755);
xnor UO_2500 (O_2500,N_24897,N_24814);
or UO_2501 (O_2501,N_24800,N_24795);
and UO_2502 (O_2502,N_24918,N_24767);
xor UO_2503 (O_2503,N_24812,N_24958);
or UO_2504 (O_2504,N_24993,N_24874);
nor UO_2505 (O_2505,N_24902,N_24863);
and UO_2506 (O_2506,N_24824,N_24808);
xnor UO_2507 (O_2507,N_24957,N_24889);
and UO_2508 (O_2508,N_24966,N_24975);
or UO_2509 (O_2509,N_24803,N_24998);
and UO_2510 (O_2510,N_24842,N_24860);
or UO_2511 (O_2511,N_24883,N_24863);
nor UO_2512 (O_2512,N_24785,N_24863);
nor UO_2513 (O_2513,N_24777,N_24834);
and UO_2514 (O_2514,N_24883,N_24770);
xnor UO_2515 (O_2515,N_24938,N_24942);
nand UO_2516 (O_2516,N_24764,N_24757);
nor UO_2517 (O_2517,N_24924,N_24781);
nand UO_2518 (O_2518,N_24829,N_24851);
and UO_2519 (O_2519,N_24943,N_24902);
xor UO_2520 (O_2520,N_24927,N_24961);
xnor UO_2521 (O_2521,N_24843,N_24911);
and UO_2522 (O_2522,N_24750,N_24772);
nor UO_2523 (O_2523,N_24957,N_24876);
or UO_2524 (O_2524,N_24958,N_24940);
nor UO_2525 (O_2525,N_24830,N_24982);
nor UO_2526 (O_2526,N_24979,N_24948);
and UO_2527 (O_2527,N_24833,N_24761);
or UO_2528 (O_2528,N_24954,N_24992);
or UO_2529 (O_2529,N_24984,N_24882);
or UO_2530 (O_2530,N_24768,N_24808);
nor UO_2531 (O_2531,N_24949,N_24881);
or UO_2532 (O_2532,N_24827,N_24773);
nor UO_2533 (O_2533,N_24869,N_24918);
or UO_2534 (O_2534,N_24858,N_24962);
and UO_2535 (O_2535,N_24982,N_24887);
xnor UO_2536 (O_2536,N_24869,N_24772);
nand UO_2537 (O_2537,N_24944,N_24762);
or UO_2538 (O_2538,N_24853,N_24968);
or UO_2539 (O_2539,N_24983,N_24900);
and UO_2540 (O_2540,N_24866,N_24801);
nand UO_2541 (O_2541,N_24971,N_24988);
nand UO_2542 (O_2542,N_24754,N_24839);
and UO_2543 (O_2543,N_24793,N_24984);
nand UO_2544 (O_2544,N_24933,N_24786);
nor UO_2545 (O_2545,N_24870,N_24988);
and UO_2546 (O_2546,N_24936,N_24912);
or UO_2547 (O_2547,N_24766,N_24990);
nor UO_2548 (O_2548,N_24793,N_24787);
nor UO_2549 (O_2549,N_24797,N_24909);
nand UO_2550 (O_2550,N_24775,N_24910);
nor UO_2551 (O_2551,N_24962,N_24916);
nand UO_2552 (O_2552,N_24851,N_24814);
or UO_2553 (O_2553,N_24835,N_24768);
nor UO_2554 (O_2554,N_24842,N_24893);
nor UO_2555 (O_2555,N_24907,N_24799);
xor UO_2556 (O_2556,N_24769,N_24782);
nand UO_2557 (O_2557,N_24789,N_24896);
xnor UO_2558 (O_2558,N_24983,N_24894);
nor UO_2559 (O_2559,N_24841,N_24889);
nand UO_2560 (O_2560,N_24833,N_24990);
and UO_2561 (O_2561,N_24873,N_24766);
nor UO_2562 (O_2562,N_24773,N_24838);
nor UO_2563 (O_2563,N_24763,N_24780);
or UO_2564 (O_2564,N_24927,N_24886);
xor UO_2565 (O_2565,N_24848,N_24952);
or UO_2566 (O_2566,N_24886,N_24909);
and UO_2567 (O_2567,N_24845,N_24831);
or UO_2568 (O_2568,N_24825,N_24779);
nor UO_2569 (O_2569,N_24864,N_24851);
or UO_2570 (O_2570,N_24811,N_24775);
and UO_2571 (O_2571,N_24957,N_24922);
nand UO_2572 (O_2572,N_24944,N_24788);
nand UO_2573 (O_2573,N_24960,N_24949);
nand UO_2574 (O_2574,N_24894,N_24779);
nand UO_2575 (O_2575,N_24942,N_24762);
nand UO_2576 (O_2576,N_24784,N_24986);
or UO_2577 (O_2577,N_24816,N_24900);
or UO_2578 (O_2578,N_24893,N_24935);
nand UO_2579 (O_2579,N_24941,N_24776);
xnor UO_2580 (O_2580,N_24755,N_24965);
nand UO_2581 (O_2581,N_24976,N_24845);
and UO_2582 (O_2582,N_24952,N_24966);
nand UO_2583 (O_2583,N_24983,N_24948);
and UO_2584 (O_2584,N_24955,N_24880);
nand UO_2585 (O_2585,N_24973,N_24873);
or UO_2586 (O_2586,N_24933,N_24959);
nand UO_2587 (O_2587,N_24811,N_24986);
and UO_2588 (O_2588,N_24788,N_24776);
nand UO_2589 (O_2589,N_24884,N_24996);
nor UO_2590 (O_2590,N_24835,N_24779);
nor UO_2591 (O_2591,N_24923,N_24937);
nand UO_2592 (O_2592,N_24952,N_24800);
xor UO_2593 (O_2593,N_24811,N_24817);
and UO_2594 (O_2594,N_24778,N_24779);
nand UO_2595 (O_2595,N_24851,N_24965);
or UO_2596 (O_2596,N_24840,N_24848);
xnor UO_2597 (O_2597,N_24882,N_24942);
and UO_2598 (O_2598,N_24959,N_24752);
nand UO_2599 (O_2599,N_24854,N_24881);
or UO_2600 (O_2600,N_24829,N_24848);
nand UO_2601 (O_2601,N_24981,N_24838);
xnor UO_2602 (O_2602,N_24864,N_24812);
xnor UO_2603 (O_2603,N_24787,N_24873);
nand UO_2604 (O_2604,N_24821,N_24995);
xnor UO_2605 (O_2605,N_24997,N_24786);
nor UO_2606 (O_2606,N_24852,N_24793);
nand UO_2607 (O_2607,N_24863,N_24991);
nor UO_2608 (O_2608,N_24788,N_24921);
nand UO_2609 (O_2609,N_24783,N_24871);
or UO_2610 (O_2610,N_24791,N_24932);
or UO_2611 (O_2611,N_24974,N_24966);
or UO_2612 (O_2612,N_24904,N_24806);
and UO_2613 (O_2613,N_24826,N_24905);
xor UO_2614 (O_2614,N_24806,N_24916);
or UO_2615 (O_2615,N_24844,N_24928);
nand UO_2616 (O_2616,N_24968,N_24811);
nand UO_2617 (O_2617,N_24894,N_24980);
and UO_2618 (O_2618,N_24873,N_24820);
xor UO_2619 (O_2619,N_24838,N_24860);
xor UO_2620 (O_2620,N_24765,N_24766);
and UO_2621 (O_2621,N_24930,N_24856);
xnor UO_2622 (O_2622,N_24855,N_24853);
or UO_2623 (O_2623,N_24898,N_24902);
xnor UO_2624 (O_2624,N_24790,N_24783);
nor UO_2625 (O_2625,N_24848,N_24924);
nor UO_2626 (O_2626,N_24924,N_24965);
and UO_2627 (O_2627,N_24916,N_24910);
nor UO_2628 (O_2628,N_24821,N_24878);
nor UO_2629 (O_2629,N_24881,N_24824);
nor UO_2630 (O_2630,N_24789,N_24774);
nand UO_2631 (O_2631,N_24827,N_24985);
and UO_2632 (O_2632,N_24787,N_24956);
nor UO_2633 (O_2633,N_24948,N_24873);
and UO_2634 (O_2634,N_24780,N_24883);
nor UO_2635 (O_2635,N_24762,N_24774);
nor UO_2636 (O_2636,N_24966,N_24884);
nor UO_2637 (O_2637,N_24914,N_24751);
xnor UO_2638 (O_2638,N_24800,N_24925);
nand UO_2639 (O_2639,N_24854,N_24986);
nor UO_2640 (O_2640,N_24886,N_24973);
nand UO_2641 (O_2641,N_24820,N_24805);
nand UO_2642 (O_2642,N_24847,N_24866);
and UO_2643 (O_2643,N_24962,N_24935);
and UO_2644 (O_2644,N_24989,N_24797);
and UO_2645 (O_2645,N_24824,N_24967);
or UO_2646 (O_2646,N_24972,N_24894);
xnor UO_2647 (O_2647,N_24771,N_24978);
nand UO_2648 (O_2648,N_24776,N_24999);
and UO_2649 (O_2649,N_24893,N_24891);
xnor UO_2650 (O_2650,N_24810,N_24914);
nand UO_2651 (O_2651,N_24995,N_24848);
xor UO_2652 (O_2652,N_24973,N_24775);
xor UO_2653 (O_2653,N_24888,N_24796);
xnor UO_2654 (O_2654,N_24814,N_24900);
nand UO_2655 (O_2655,N_24991,N_24934);
or UO_2656 (O_2656,N_24809,N_24852);
nand UO_2657 (O_2657,N_24773,N_24781);
nand UO_2658 (O_2658,N_24769,N_24990);
and UO_2659 (O_2659,N_24886,N_24817);
xnor UO_2660 (O_2660,N_24820,N_24819);
and UO_2661 (O_2661,N_24751,N_24954);
or UO_2662 (O_2662,N_24834,N_24825);
nand UO_2663 (O_2663,N_24862,N_24802);
nand UO_2664 (O_2664,N_24992,N_24934);
and UO_2665 (O_2665,N_24912,N_24952);
or UO_2666 (O_2666,N_24834,N_24900);
xor UO_2667 (O_2667,N_24937,N_24807);
nor UO_2668 (O_2668,N_24933,N_24998);
and UO_2669 (O_2669,N_24936,N_24813);
or UO_2670 (O_2670,N_24897,N_24790);
xnor UO_2671 (O_2671,N_24750,N_24966);
xor UO_2672 (O_2672,N_24837,N_24936);
xnor UO_2673 (O_2673,N_24803,N_24966);
nand UO_2674 (O_2674,N_24992,N_24866);
xnor UO_2675 (O_2675,N_24964,N_24859);
nand UO_2676 (O_2676,N_24907,N_24756);
and UO_2677 (O_2677,N_24831,N_24794);
xnor UO_2678 (O_2678,N_24833,N_24885);
or UO_2679 (O_2679,N_24857,N_24936);
xor UO_2680 (O_2680,N_24789,N_24915);
or UO_2681 (O_2681,N_24861,N_24953);
nand UO_2682 (O_2682,N_24886,N_24751);
xor UO_2683 (O_2683,N_24812,N_24966);
nand UO_2684 (O_2684,N_24850,N_24791);
xor UO_2685 (O_2685,N_24912,N_24763);
nand UO_2686 (O_2686,N_24796,N_24792);
and UO_2687 (O_2687,N_24857,N_24779);
nand UO_2688 (O_2688,N_24865,N_24944);
nand UO_2689 (O_2689,N_24801,N_24920);
nor UO_2690 (O_2690,N_24766,N_24937);
nor UO_2691 (O_2691,N_24819,N_24942);
nor UO_2692 (O_2692,N_24885,N_24825);
or UO_2693 (O_2693,N_24824,N_24900);
xnor UO_2694 (O_2694,N_24794,N_24834);
and UO_2695 (O_2695,N_24807,N_24783);
or UO_2696 (O_2696,N_24860,N_24886);
nor UO_2697 (O_2697,N_24862,N_24783);
nand UO_2698 (O_2698,N_24899,N_24780);
xor UO_2699 (O_2699,N_24882,N_24920);
and UO_2700 (O_2700,N_24761,N_24885);
nand UO_2701 (O_2701,N_24984,N_24795);
nand UO_2702 (O_2702,N_24940,N_24975);
nand UO_2703 (O_2703,N_24911,N_24786);
or UO_2704 (O_2704,N_24976,N_24850);
and UO_2705 (O_2705,N_24966,N_24900);
or UO_2706 (O_2706,N_24921,N_24942);
and UO_2707 (O_2707,N_24934,N_24757);
nor UO_2708 (O_2708,N_24840,N_24987);
xnor UO_2709 (O_2709,N_24877,N_24951);
or UO_2710 (O_2710,N_24806,N_24966);
and UO_2711 (O_2711,N_24810,N_24800);
xor UO_2712 (O_2712,N_24858,N_24812);
xnor UO_2713 (O_2713,N_24915,N_24768);
or UO_2714 (O_2714,N_24982,N_24884);
xnor UO_2715 (O_2715,N_24903,N_24762);
or UO_2716 (O_2716,N_24803,N_24851);
or UO_2717 (O_2717,N_24976,N_24808);
nor UO_2718 (O_2718,N_24785,N_24888);
and UO_2719 (O_2719,N_24876,N_24992);
nor UO_2720 (O_2720,N_24789,N_24856);
and UO_2721 (O_2721,N_24816,N_24889);
or UO_2722 (O_2722,N_24804,N_24956);
xnor UO_2723 (O_2723,N_24841,N_24858);
nand UO_2724 (O_2724,N_24901,N_24912);
nand UO_2725 (O_2725,N_24929,N_24960);
or UO_2726 (O_2726,N_24911,N_24807);
or UO_2727 (O_2727,N_24954,N_24820);
nor UO_2728 (O_2728,N_24796,N_24751);
and UO_2729 (O_2729,N_24863,N_24948);
xnor UO_2730 (O_2730,N_24776,N_24818);
nor UO_2731 (O_2731,N_24803,N_24832);
nor UO_2732 (O_2732,N_24855,N_24995);
or UO_2733 (O_2733,N_24853,N_24960);
or UO_2734 (O_2734,N_24994,N_24899);
xor UO_2735 (O_2735,N_24982,N_24924);
nand UO_2736 (O_2736,N_24980,N_24974);
and UO_2737 (O_2737,N_24806,N_24885);
xnor UO_2738 (O_2738,N_24841,N_24782);
and UO_2739 (O_2739,N_24862,N_24989);
nor UO_2740 (O_2740,N_24944,N_24859);
xor UO_2741 (O_2741,N_24844,N_24762);
xor UO_2742 (O_2742,N_24780,N_24873);
nor UO_2743 (O_2743,N_24805,N_24780);
xor UO_2744 (O_2744,N_24799,N_24930);
and UO_2745 (O_2745,N_24801,N_24992);
nand UO_2746 (O_2746,N_24994,N_24985);
nor UO_2747 (O_2747,N_24780,N_24995);
or UO_2748 (O_2748,N_24906,N_24882);
nand UO_2749 (O_2749,N_24876,N_24849);
nand UO_2750 (O_2750,N_24839,N_24766);
nor UO_2751 (O_2751,N_24846,N_24949);
or UO_2752 (O_2752,N_24754,N_24922);
or UO_2753 (O_2753,N_24821,N_24772);
and UO_2754 (O_2754,N_24861,N_24892);
or UO_2755 (O_2755,N_24821,N_24794);
or UO_2756 (O_2756,N_24834,N_24920);
nand UO_2757 (O_2757,N_24878,N_24934);
nor UO_2758 (O_2758,N_24788,N_24929);
xnor UO_2759 (O_2759,N_24910,N_24764);
nand UO_2760 (O_2760,N_24844,N_24837);
nor UO_2761 (O_2761,N_24928,N_24759);
and UO_2762 (O_2762,N_24824,N_24849);
xor UO_2763 (O_2763,N_24862,N_24826);
xor UO_2764 (O_2764,N_24900,N_24955);
xnor UO_2765 (O_2765,N_24832,N_24946);
nand UO_2766 (O_2766,N_24774,N_24886);
nor UO_2767 (O_2767,N_24931,N_24761);
or UO_2768 (O_2768,N_24782,N_24995);
nand UO_2769 (O_2769,N_24757,N_24903);
or UO_2770 (O_2770,N_24862,N_24998);
or UO_2771 (O_2771,N_24990,N_24760);
nor UO_2772 (O_2772,N_24853,N_24955);
xor UO_2773 (O_2773,N_24887,N_24814);
xor UO_2774 (O_2774,N_24761,N_24778);
nor UO_2775 (O_2775,N_24803,N_24988);
xor UO_2776 (O_2776,N_24979,N_24965);
and UO_2777 (O_2777,N_24865,N_24779);
or UO_2778 (O_2778,N_24891,N_24931);
xor UO_2779 (O_2779,N_24893,N_24928);
nand UO_2780 (O_2780,N_24915,N_24961);
xor UO_2781 (O_2781,N_24773,N_24777);
nor UO_2782 (O_2782,N_24985,N_24785);
and UO_2783 (O_2783,N_24974,N_24786);
nor UO_2784 (O_2784,N_24838,N_24761);
or UO_2785 (O_2785,N_24774,N_24777);
xnor UO_2786 (O_2786,N_24783,N_24994);
and UO_2787 (O_2787,N_24909,N_24996);
nand UO_2788 (O_2788,N_24786,N_24943);
or UO_2789 (O_2789,N_24796,N_24843);
nor UO_2790 (O_2790,N_24937,N_24883);
xnor UO_2791 (O_2791,N_24883,N_24789);
nand UO_2792 (O_2792,N_24900,N_24923);
or UO_2793 (O_2793,N_24823,N_24969);
or UO_2794 (O_2794,N_24951,N_24948);
xnor UO_2795 (O_2795,N_24928,N_24978);
and UO_2796 (O_2796,N_24831,N_24944);
nor UO_2797 (O_2797,N_24987,N_24958);
and UO_2798 (O_2798,N_24918,N_24904);
nand UO_2799 (O_2799,N_24981,N_24770);
or UO_2800 (O_2800,N_24978,N_24988);
nand UO_2801 (O_2801,N_24861,N_24864);
and UO_2802 (O_2802,N_24933,N_24891);
and UO_2803 (O_2803,N_24879,N_24923);
and UO_2804 (O_2804,N_24897,N_24763);
or UO_2805 (O_2805,N_24788,N_24895);
and UO_2806 (O_2806,N_24933,N_24844);
nor UO_2807 (O_2807,N_24914,N_24756);
or UO_2808 (O_2808,N_24960,N_24881);
nand UO_2809 (O_2809,N_24865,N_24778);
or UO_2810 (O_2810,N_24860,N_24909);
nor UO_2811 (O_2811,N_24944,N_24984);
nand UO_2812 (O_2812,N_24751,N_24753);
xnor UO_2813 (O_2813,N_24848,N_24914);
xnor UO_2814 (O_2814,N_24898,N_24888);
nand UO_2815 (O_2815,N_24823,N_24771);
nor UO_2816 (O_2816,N_24896,N_24910);
or UO_2817 (O_2817,N_24773,N_24764);
or UO_2818 (O_2818,N_24956,N_24913);
and UO_2819 (O_2819,N_24955,N_24918);
and UO_2820 (O_2820,N_24979,N_24869);
nor UO_2821 (O_2821,N_24769,N_24865);
nand UO_2822 (O_2822,N_24859,N_24852);
xnor UO_2823 (O_2823,N_24937,N_24755);
or UO_2824 (O_2824,N_24810,N_24994);
and UO_2825 (O_2825,N_24915,N_24774);
nor UO_2826 (O_2826,N_24848,N_24768);
xnor UO_2827 (O_2827,N_24848,N_24954);
nand UO_2828 (O_2828,N_24972,N_24824);
and UO_2829 (O_2829,N_24832,N_24898);
xor UO_2830 (O_2830,N_24982,N_24822);
xnor UO_2831 (O_2831,N_24884,N_24991);
nand UO_2832 (O_2832,N_24811,N_24940);
nand UO_2833 (O_2833,N_24835,N_24934);
and UO_2834 (O_2834,N_24899,N_24935);
and UO_2835 (O_2835,N_24947,N_24868);
or UO_2836 (O_2836,N_24779,N_24797);
and UO_2837 (O_2837,N_24917,N_24947);
and UO_2838 (O_2838,N_24774,N_24822);
nand UO_2839 (O_2839,N_24763,N_24810);
nor UO_2840 (O_2840,N_24857,N_24877);
or UO_2841 (O_2841,N_24894,N_24769);
nand UO_2842 (O_2842,N_24911,N_24888);
or UO_2843 (O_2843,N_24792,N_24771);
and UO_2844 (O_2844,N_24848,N_24851);
or UO_2845 (O_2845,N_24903,N_24977);
nor UO_2846 (O_2846,N_24881,N_24880);
or UO_2847 (O_2847,N_24872,N_24829);
nor UO_2848 (O_2848,N_24831,N_24950);
xor UO_2849 (O_2849,N_24803,N_24870);
nand UO_2850 (O_2850,N_24805,N_24887);
and UO_2851 (O_2851,N_24772,N_24961);
xor UO_2852 (O_2852,N_24770,N_24824);
xnor UO_2853 (O_2853,N_24836,N_24783);
nor UO_2854 (O_2854,N_24856,N_24992);
and UO_2855 (O_2855,N_24782,N_24817);
xnor UO_2856 (O_2856,N_24908,N_24953);
or UO_2857 (O_2857,N_24968,N_24938);
or UO_2858 (O_2858,N_24777,N_24870);
nand UO_2859 (O_2859,N_24961,N_24750);
nor UO_2860 (O_2860,N_24876,N_24891);
nand UO_2861 (O_2861,N_24860,N_24801);
nand UO_2862 (O_2862,N_24951,N_24822);
nand UO_2863 (O_2863,N_24929,N_24996);
nor UO_2864 (O_2864,N_24940,N_24912);
nor UO_2865 (O_2865,N_24791,N_24855);
xnor UO_2866 (O_2866,N_24976,N_24767);
nor UO_2867 (O_2867,N_24851,N_24916);
nand UO_2868 (O_2868,N_24990,N_24775);
or UO_2869 (O_2869,N_24949,N_24967);
xor UO_2870 (O_2870,N_24903,N_24891);
and UO_2871 (O_2871,N_24985,N_24756);
nor UO_2872 (O_2872,N_24952,N_24949);
nor UO_2873 (O_2873,N_24803,N_24935);
nor UO_2874 (O_2874,N_24767,N_24978);
nor UO_2875 (O_2875,N_24841,N_24853);
nor UO_2876 (O_2876,N_24803,N_24842);
nand UO_2877 (O_2877,N_24948,N_24964);
xnor UO_2878 (O_2878,N_24909,N_24837);
nand UO_2879 (O_2879,N_24779,N_24853);
nand UO_2880 (O_2880,N_24845,N_24832);
xor UO_2881 (O_2881,N_24883,N_24871);
nor UO_2882 (O_2882,N_24997,N_24769);
nor UO_2883 (O_2883,N_24885,N_24931);
nor UO_2884 (O_2884,N_24939,N_24882);
and UO_2885 (O_2885,N_24997,N_24859);
xor UO_2886 (O_2886,N_24997,N_24991);
nor UO_2887 (O_2887,N_24835,N_24760);
and UO_2888 (O_2888,N_24884,N_24760);
and UO_2889 (O_2889,N_24988,N_24769);
nand UO_2890 (O_2890,N_24850,N_24875);
xor UO_2891 (O_2891,N_24912,N_24780);
xnor UO_2892 (O_2892,N_24888,N_24875);
nor UO_2893 (O_2893,N_24766,N_24940);
xor UO_2894 (O_2894,N_24817,N_24999);
xnor UO_2895 (O_2895,N_24816,N_24884);
nand UO_2896 (O_2896,N_24766,N_24907);
or UO_2897 (O_2897,N_24857,N_24975);
and UO_2898 (O_2898,N_24812,N_24987);
nor UO_2899 (O_2899,N_24830,N_24946);
nor UO_2900 (O_2900,N_24955,N_24928);
and UO_2901 (O_2901,N_24809,N_24902);
xor UO_2902 (O_2902,N_24760,N_24951);
nand UO_2903 (O_2903,N_24903,N_24985);
xor UO_2904 (O_2904,N_24961,N_24942);
nor UO_2905 (O_2905,N_24984,N_24797);
xor UO_2906 (O_2906,N_24967,N_24879);
nand UO_2907 (O_2907,N_24846,N_24977);
and UO_2908 (O_2908,N_24817,N_24892);
and UO_2909 (O_2909,N_24894,N_24883);
or UO_2910 (O_2910,N_24894,N_24931);
nand UO_2911 (O_2911,N_24931,N_24829);
xnor UO_2912 (O_2912,N_24993,N_24939);
or UO_2913 (O_2913,N_24981,N_24949);
nand UO_2914 (O_2914,N_24968,N_24876);
and UO_2915 (O_2915,N_24974,N_24946);
nand UO_2916 (O_2916,N_24800,N_24950);
nand UO_2917 (O_2917,N_24813,N_24801);
or UO_2918 (O_2918,N_24964,N_24812);
nand UO_2919 (O_2919,N_24857,N_24890);
xor UO_2920 (O_2920,N_24861,N_24921);
nand UO_2921 (O_2921,N_24893,N_24831);
nand UO_2922 (O_2922,N_24944,N_24914);
xnor UO_2923 (O_2923,N_24763,N_24938);
nand UO_2924 (O_2924,N_24781,N_24905);
nand UO_2925 (O_2925,N_24884,N_24865);
xor UO_2926 (O_2926,N_24870,N_24959);
and UO_2927 (O_2927,N_24851,N_24911);
xnor UO_2928 (O_2928,N_24866,N_24798);
and UO_2929 (O_2929,N_24915,N_24916);
nor UO_2930 (O_2930,N_24874,N_24917);
xor UO_2931 (O_2931,N_24857,N_24768);
and UO_2932 (O_2932,N_24859,N_24991);
nor UO_2933 (O_2933,N_24895,N_24879);
xor UO_2934 (O_2934,N_24759,N_24962);
or UO_2935 (O_2935,N_24962,N_24887);
nand UO_2936 (O_2936,N_24797,N_24926);
or UO_2937 (O_2937,N_24778,N_24951);
nand UO_2938 (O_2938,N_24759,N_24929);
xnor UO_2939 (O_2939,N_24923,N_24930);
nor UO_2940 (O_2940,N_24965,N_24867);
nor UO_2941 (O_2941,N_24874,N_24869);
xnor UO_2942 (O_2942,N_24856,N_24799);
xor UO_2943 (O_2943,N_24838,N_24954);
nor UO_2944 (O_2944,N_24979,N_24960);
nand UO_2945 (O_2945,N_24809,N_24985);
or UO_2946 (O_2946,N_24943,N_24938);
nand UO_2947 (O_2947,N_24855,N_24757);
or UO_2948 (O_2948,N_24758,N_24958);
xnor UO_2949 (O_2949,N_24901,N_24902);
nand UO_2950 (O_2950,N_24905,N_24901);
and UO_2951 (O_2951,N_24855,N_24756);
and UO_2952 (O_2952,N_24761,N_24750);
nor UO_2953 (O_2953,N_24945,N_24909);
nor UO_2954 (O_2954,N_24909,N_24760);
and UO_2955 (O_2955,N_24992,N_24762);
and UO_2956 (O_2956,N_24750,N_24915);
and UO_2957 (O_2957,N_24995,N_24859);
nand UO_2958 (O_2958,N_24841,N_24799);
and UO_2959 (O_2959,N_24978,N_24777);
nor UO_2960 (O_2960,N_24772,N_24803);
or UO_2961 (O_2961,N_24804,N_24838);
xor UO_2962 (O_2962,N_24845,N_24760);
or UO_2963 (O_2963,N_24985,N_24768);
or UO_2964 (O_2964,N_24812,N_24857);
nor UO_2965 (O_2965,N_24897,N_24813);
or UO_2966 (O_2966,N_24787,N_24779);
and UO_2967 (O_2967,N_24940,N_24869);
nor UO_2968 (O_2968,N_24978,N_24975);
xnor UO_2969 (O_2969,N_24799,N_24998);
xor UO_2970 (O_2970,N_24836,N_24865);
or UO_2971 (O_2971,N_24923,N_24865);
and UO_2972 (O_2972,N_24766,N_24938);
xnor UO_2973 (O_2973,N_24977,N_24923);
xnor UO_2974 (O_2974,N_24897,N_24969);
xnor UO_2975 (O_2975,N_24866,N_24923);
xor UO_2976 (O_2976,N_24760,N_24834);
and UO_2977 (O_2977,N_24989,N_24839);
xnor UO_2978 (O_2978,N_24936,N_24923);
and UO_2979 (O_2979,N_24989,N_24934);
nor UO_2980 (O_2980,N_24895,N_24884);
nor UO_2981 (O_2981,N_24811,N_24795);
nor UO_2982 (O_2982,N_24856,N_24859);
and UO_2983 (O_2983,N_24797,N_24945);
nand UO_2984 (O_2984,N_24897,N_24890);
nor UO_2985 (O_2985,N_24847,N_24924);
or UO_2986 (O_2986,N_24848,N_24892);
and UO_2987 (O_2987,N_24968,N_24857);
or UO_2988 (O_2988,N_24851,N_24837);
or UO_2989 (O_2989,N_24794,N_24837);
nand UO_2990 (O_2990,N_24756,N_24930);
xnor UO_2991 (O_2991,N_24907,N_24980);
xnor UO_2992 (O_2992,N_24778,N_24754);
and UO_2993 (O_2993,N_24826,N_24940);
xnor UO_2994 (O_2994,N_24808,N_24833);
or UO_2995 (O_2995,N_24763,N_24766);
and UO_2996 (O_2996,N_24763,N_24759);
nand UO_2997 (O_2997,N_24954,N_24860);
nor UO_2998 (O_2998,N_24972,N_24799);
or UO_2999 (O_2999,N_24752,N_24753);
endmodule