module basic_750_5000_1000_25_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_626,In_389);
and U1 (N_1,In_660,In_593);
and U2 (N_2,In_676,In_373);
nand U3 (N_3,In_737,In_192);
xor U4 (N_4,In_422,In_605);
nor U5 (N_5,In_323,In_410);
or U6 (N_6,In_625,In_187);
and U7 (N_7,In_69,In_519);
nand U8 (N_8,In_161,In_189);
and U9 (N_9,In_469,In_491);
nor U10 (N_10,In_585,In_569);
nand U11 (N_11,In_729,In_36);
xor U12 (N_12,In_116,In_450);
nand U13 (N_13,In_72,In_412);
and U14 (N_14,In_398,In_61);
nand U15 (N_15,In_197,In_378);
nand U16 (N_16,In_468,In_427);
xnor U17 (N_17,In_141,In_13);
xor U18 (N_18,In_163,In_102);
nand U19 (N_19,In_228,In_249);
nor U20 (N_20,In_14,In_202);
nand U21 (N_21,In_52,In_279);
and U22 (N_22,In_83,In_308);
nand U23 (N_23,In_91,In_735);
or U24 (N_24,In_289,In_63);
and U25 (N_25,In_413,In_226);
nor U26 (N_26,In_399,In_171);
nor U27 (N_27,In_407,In_602);
nand U28 (N_28,In_423,In_46);
nand U29 (N_29,In_408,In_143);
and U30 (N_30,In_665,In_478);
nor U31 (N_31,In_333,In_681);
and U32 (N_32,In_154,In_653);
and U33 (N_33,In_432,In_292);
or U34 (N_34,In_122,In_674);
nor U35 (N_35,In_41,In_632);
and U36 (N_36,In_586,In_430);
and U37 (N_37,In_730,In_578);
or U38 (N_38,In_240,In_424);
xnor U39 (N_39,In_343,In_652);
nand U40 (N_40,In_379,In_415);
or U41 (N_41,In_58,In_629);
and U42 (N_42,In_482,In_8);
or U43 (N_43,In_10,In_623);
or U44 (N_44,In_721,In_731);
nor U45 (N_45,In_554,In_120);
nor U46 (N_46,In_417,In_749);
or U47 (N_47,In_179,In_640);
or U48 (N_48,In_261,In_541);
and U49 (N_49,In_12,In_612);
nand U50 (N_50,In_638,In_268);
or U51 (N_51,In_217,In_85);
nor U52 (N_52,In_3,In_195);
nand U53 (N_53,In_474,In_354);
xor U54 (N_54,In_448,In_386);
nor U55 (N_55,In_734,In_700);
xor U56 (N_56,In_551,In_212);
nor U57 (N_57,In_374,In_62);
xnor U58 (N_58,In_156,In_64);
and U59 (N_59,In_57,In_565);
or U60 (N_60,In_732,In_304);
nand U61 (N_61,In_377,In_403);
and U62 (N_62,In_113,In_99);
or U63 (N_63,In_515,In_142);
and U64 (N_64,In_24,In_512);
nand U65 (N_65,In_748,In_743);
or U66 (N_66,In_339,In_370);
and U67 (N_67,In_622,In_724);
and U68 (N_68,In_693,In_742);
and U69 (N_69,In_401,In_131);
xnor U70 (N_70,In_15,In_137);
and U71 (N_71,In_96,In_574);
or U72 (N_72,In_263,In_296);
and U73 (N_73,In_90,In_118);
nand U74 (N_74,In_151,In_522);
and U75 (N_75,In_719,In_500);
nor U76 (N_76,In_738,In_95);
nor U77 (N_77,In_4,In_677);
or U78 (N_78,In_68,In_506);
nand U79 (N_79,In_678,In_656);
and U80 (N_80,In_336,In_411);
nor U81 (N_81,In_53,In_646);
xor U82 (N_82,In_624,In_525);
and U83 (N_83,In_453,In_659);
and U84 (N_84,In_250,In_117);
nand U85 (N_85,In_357,In_293);
nor U86 (N_86,In_556,In_526);
nand U87 (N_87,In_6,In_497);
and U88 (N_88,In_21,In_581);
or U89 (N_89,In_572,In_546);
and U90 (N_90,In_347,In_567);
nand U91 (N_91,In_45,In_209);
nand U92 (N_92,In_211,In_668);
nor U93 (N_93,In_695,In_358);
nand U94 (N_94,In_105,In_319);
nand U95 (N_95,In_534,In_488);
nand U96 (N_96,In_229,In_313);
and U97 (N_97,In_445,In_194);
nand U98 (N_98,In_218,In_260);
and U99 (N_99,In_178,In_455);
or U100 (N_100,In_571,In_404);
or U101 (N_101,In_346,In_663);
or U102 (N_102,In_560,In_577);
nand U103 (N_103,In_717,In_591);
and U104 (N_104,In_144,In_636);
and U105 (N_105,In_307,In_690);
or U106 (N_106,In_387,In_709);
nor U107 (N_107,In_93,In_236);
or U108 (N_108,In_42,In_54);
or U109 (N_109,In_564,In_278);
and U110 (N_110,In_238,In_299);
nor U111 (N_111,In_698,In_691);
or U112 (N_112,In_627,In_705);
and U113 (N_113,In_2,In_380);
nand U114 (N_114,In_50,In_675);
and U115 (N_115,In_504,In_106);
and U116 (N_116,In_685,In_28);
nand U117 (N_117,In_366,In_11);
or U118 (N_118,In_470,In_210);
xnor U119 (N_119,In_26,In_138);
nor U120 (N_120,In_266,In_460);
xor U121 (N_121,In_739,In_265);
nor U122 (N_122,In_561,In_56);
nor U123 (N_123,In_542,In_254);
nand U124 (N_124,In_435,In_312);
and U125 (N_125,In_532,In_222);
and U126 (N_126,In_73,In_670);
xnor U127 (N_127,In_207,In_146);
nor U128 (N_128,In_394,In_110);
nand U129 (N_129,In_606,In_177);
xor U130 (N_130,In_544,In_184);
nand U131 (N_131,In_563,In_485);
nor U132 (N_132,In_37,In_174);
nand U133 (N_133,In_420,In_81);
nand U134 (N_134,In_5,In_598);
nor U135 (N_135,In_123,In_188);
and U136 (N_136,In_449,In_508);
or U137 (N_137,In_277,In_60);
nand U138 (N_138,In_475,In_588);
and U139 (N_139,In_267,In_597);
nor U140 (N_140,In_199,In_216);
or U141 (N_141,In_67,In_434);
nor U142 (N_142,In_558,In_74);
and U143 (N_143,In_327,In_348);
and U144 (N_144,In_301,In_716);
nor U145 (N_145,In_396,In_344);
nor U146 (N_146,In_329,In_35);
xor U147 (N_147,In_555,In_440);
nor U148 (N_148,In_306,In_584);
nand U149 (N_149,In_484,In_227);
or U150 (N_150,In_518,In_426);
or U151 (N_151,In_298,In_490);
and U152 (N_152,In_165,In_230);
nor U153 (N_153,In_364,In_487);
nor U154 (N_154,In_44,In_609);
nor U155 (N_155,In_523,In_84);
nor U156 (N_156,In_23,In_65);
and U157 (N_157,In_334,In_367);
nor U158 (N_158,In_704,In_594);
and U159 (N_159,In_191,In_466);
nand U160 (N_160,In_740,In_129);
and U161 (N_161,In_545,In_124);
and U162 (N_162,In_726,In_309);
and U163 (N_163,In_371,In_352);
or U164 (N_164,In_481,In_295);
xnor U165 (N_165,In_528,In_98);
nor U166 (N_166,In_390,In_645);
or U167 (N_167,In_507,In_248);
and U168 (N_168,In_159,In_642);
nand U169 (N_169,In_176,In_692);
and U170 (N_170,In_40,In_509);
nand U171 (N_171,In_425,In_673);
nor U172 (N_172,In_337,In_573);
or U173 (N_173,In_477,In_140);
and U174 (N_174,In_587,In_237);
nand U175 (N_175,In_479,In_157);
or U176 (N_176,In_172,In_49);
nand U177 (N_177,In_182,In_535);
nand U178 (N_178,In_43,In_583);
xnor U179 (N_179,In_436,In_531);
nand U180 (N_180,In_97,In_70);
xnor U181 (N_181,In_242,In_51);
nor U182 (N_182,In_701,In_158);
and U183 (N_183,In_662,In_125);
or U184 (N_184,In_383,In_282);
nand U185 (N_185,In_667,In_232);
and U186 (N_186,In_233,In_275);
and U187 (N_187,In_747,In_421);
nor U188 (N_188,In_527,In_71);
and U189 (N_189,In_335,In_169);
or U190 (N_190,In_471,In_687);
or U191 (N_191,In_688,In_603);
and U192 (N_192,In_369,In_231);
nor U193 (N_193,In_345,In_649);
and U194 (N_194,In_433,In_280);
or U195 (N_195,In_461,In_437);
and U196 (N_196,In_100,In_127);
and U197 (N_197,In_181,In_221);
nand U198 (N_198,In_702,In_499);
nand U199 (N_199,In_316,In_359);
and U200 (N_200,In_326,In_273);
nand U201 (N_201,N_101,In_286);
and U202 (N_202,N_141,In_214);
xnor U203 (N_203,N_45,N_65);
nor U204 (N_204,N_196,In_297);
xor U205 (N_205,In_589,In_294);
nand U206 (N_206,N_12,N_33);
nor U207 (N_207,In_89,In_145);
nor U208 (N_208,In_9,In_384);
nand U209 (N_209,In_175,In_405);
and U210 (N_210,N_32,In_703);
nor U211 (N_211,N_177,N_193);
nor U212 (N_212,In_203,In_397);
nand U213 (N_213,In_454,In_164);
nor U214 (N_214,N_174,N_176);
nor U215 (N_215,N_164,In_338);
or U216 (N_216,N_168,In_224);
nor U217 (N_217,In_314,N_105);
nand U218 (N_218,In_291,N_165);
and U219 (N_219,N_37,In_392);
or U220 (N_220,In_18,N_70);
or U221 (N_221,In_391,In_310);
and U222 (N_222,In_245,In_262);
and U223 (N_223,In_576,In_243);
and U224 (N_224,In_111,In_633);
and U225 (N_225,N_23,N_10);
xor U226 (N_226,N_83,In_457);
nand U227 (N_227,N_92,N_186);
nor U228 (N_228,In_686,In_672);
and U229 (N_229,In_315,In_283);
and U230 (N_230,In_728,In_575);
xor U231 (N_231,In_451,In_600);
nand U232 (N_232,In_637,N_87);
nand U233 (N_233,N_156,In_416);
nor U234 (N_234,In_135,In_543);
and U235 (N_235,In_630,N_154);
and U236 (N_236,In_382,In_270);
or U237 (N_237,In_38,In_502);
xor U238 (N_238,In_167,In_317);
xor U239 (N_239,N_55,N_24);
or U240 (N_240,In_109,In_616);
xnor U241 (N_241,In_160,In_276);
nor U242 (N_242,N_73,N_145);
or U243 (N_243,In_155,In_119);
nor U244 (N_244,In_537,In_467);
and U245 (N_245,In_269,In_419);
and U246 (N_246,N_30,In_208);
and U247 (N_247,In_514,N_98);
nand U248 (N_248,N_116,N_89);
xnor U249 (N_249,N_63,In_720);
nor U250 (N_250,N_64,N_52);
and U251 (N_251,N_80,In_362);
nor U252 (N_252,In_441,In_643);
and U253 (N_253,In_150,In_718);
xor U254 (N_254,In_332,In_568);
xnor U255 (N_255,In_496,N_113);
or U256 (N_256,In_342,In_548);
or U257 (N_257,In_80,N_88);
and U258 (N_258,N_178,In_439);
nor U259 (N_259,In_17,N_48);
and U260 (N_260,In_682,In_444);
nand U261 (N_261,In_552,In_16);
xor U262 (N_262,In_592,In_274);
or U263 (N_263,N_152,In_213);
or U264 (N_264,N_163,In_406);
nand U265 (N_265,In_480,In_644);
xnor U266 (N_266,In_234,In_353);
xor U267 (N_267,In_385,N_190);
xnor U268 (N_268,In_259,In_320);
nand U269 (N_269,In_112,In_579);
nand U270 (N_270,N_199,In_680);
nand U271 (N_271,In_599,N_155);
and U272 (N_272,In_418,N_90);
and U273 (N_273,In_431,N_97);
and U274 (N_274,N_137,In_284);
and U275 (N_275,N_104,N_11);
and U276 (N_276,In_429,In_247);
nand U277 (N_277,In_305,In_549);
nor U278 (N_278,N_69,N_15);
and U279 (N_279,In_86,N_138);
and U280 (N_280,In_654,N_41);
or U281 (N_281,In_473,In_710);
or U282 (N_282,In_550,In_340);
and U283 (N_283,In_132,In_87);
or U284 (N_284,N_71,In_281);
nor U285 (N_285,In_683,In_511);
nand U286 (N_286,N_161,N_44);
and U287 (N_287,In_255,In_501);
nand U288 (N_288,N_151,In_341);
nand U289 (N_289,N_54,In_498);
nand U290 (N_290,N_28,In_648);
nor U291 (N_291,In_31,In_241);
nand U292 (N_292,N_56,N_153);
nor U293 (N_293,N_171,N_5);
or U294 (N_294,N_170,In_325);
and U295 (N_295,In_559,N_128);
nor U296 (N_296,N_46,N_17);
and U297 (N_297,In_104,In_530);
and U298 (N_298,In_495,N_96);
and U299 (N_299,In_539,In_27);
nand U300 (N_300,In_253,N_47);
and U301 (N_301,In_66,In_607);
nand U302 (N_302,N_27,In_614);
nor U303 (N_303,In_88,In_246);
or U304 (N_304,In_723,In_465);
and U305 (N_305,N_93,In_462);
xor U306 (N_306,In_697,N_182);
nor U307 (N_307,In_0,In_349);
nand U308 (N_308,In_368,N_57);
or U309 (N_309,In_139,In_635);
or U310 (N_310,In_570,In_483);
and U311 (N_311,In_20,N_185);
or U312 (N_312,In_664,In_153);
and U313 (N_313,In_47,In_355);
nand U314 (N_314,In_183,In_442);
or U315 (N_315,In_608,In_736);
xnor U316 (N_316,In_540,In_148);
xnor U317 (N_317,N_82,In_34);
and U318 (N_318,In_76,In_185);
nor U319 (N_319,N_144,N_121);
nor U320 (N_320,In_741,N_132);
nor U321 (N_321,N_139,In_595);
or U322 (N_322,N_166,In_712);
nor U323 (N_323,N_78,N_157);
and U324 (N_324,In_324,N_131);
xnor U325 (N_325,In_162,N_142);
and U326 (N_326,In_714,In_30);
and U327 (N_327,In_356,In_447);
or U328 (N_328,In_621,In_493);
and U329 (N_329,N_94,In_513);
and U330 (N_330,In_494,N_86);
or U331 (N_331,N_79,In_503);
nand U332 (N_332,In_330,In_566);
and U333 (N_333,In_562,In_517);
or U334 (N_334,In_205,N_3);
nor U335 (N_335,In_696,In_39);
nand U336 (N_336,In_631,N_39);
and U337 (N_337,In_147,N_22);
and U338 (N_338,N_21,In_101);
or U339 (N_339,In_198,In_393);
nor U340 (N_340,In_264,N_167);
and U341 (N_341,In_725,N_100);
nor U342 (N_342,N_109,N_124);
nand U343 (N_343,In_428,In_19);
nor U344 (N_344,In_360,In_596);
or U345 (N_345,N_173,N_130);
or U346 (N_346,In_33,N_99);
or U347 (N_347,N_112,In_476);
nor U348 (N_348,In_582,In_464);
or U349 (N_349,In_59,In_29);
nor U350 (N_350,N_42,In_557);
and U351 (N_351,In_524,In_708);
and U352 (N_352,N_76,In_235);
nor U353 (N_353,N_103,In_381);
nor U354 (N_354,In_553,N_172);
and U355 (N_355,N_43,In_201);
or U356 (N_356,N_191,In_168);
and U357 (N_357,N_9,In_452);
nand U358 (N_358,N_7,In_617);
nand U359 (N_359,N_61,In_287);
nand U360 (N_360,N_146,N_35);
or U361 (N_361,In_538,N_187);
or U362 (N_362,In_707,N_38);
or U363 (N_363,In_115,N_25);
and U364 (N_364,N_62,N_72);
or U365 (N_365,In_285,N_160);
nand U366 (N_366,In_744,In_618);
nand U367 (N_367,In_661,N_0);
nand U368 (N_368,N_6,In_400);
nor U369 (N_369,N_175,In_611);
and U370 (N_370,In_489,In_215);
nand U371 (N_371,In_290,In_258);
and U372 (N_372,In_650,In_402);
nor U373 (N_373,N_108,N_127);
nand U374 (N_374,In_82,In_22);
or U375 (N_375,In_322,N_189);
and U376 (N_376,In_170,In_492);
xnor U377 (N_377,In_733,In_679);
and U378 (N_378,N_66,In_79);
xnor U379 (N_379,In_529,In_601);
or U380 (N_380,In_318,In_166);
nor U381 (N_381,In_48,In_409);
nor U382 (N_382,N_81,In_658);
nor U383 (N_383,N_125,N_49);
nand U384 (N_384,In_363,N_77);
and U385 (N_385,In_580,In_300);
nor U386 (N_386,In_7,In_77);
or U387 (N_387,In_134,N_14);
nand U388 (N_388,In_533,In_372);
or U389 (N_389,In_126,N_20);
or U390 (N_390,N_129,N_95);
nand U391 (N_391,N_51,N_58);
nor U392 (N_392,In_395,In_244);
nor U393 (N_393,In_114,N_75);
nand U394 (N_394,In_620,In_414);
nor U395 (N_395,In_302,N_68);
nand U396 (N_396,N_162,In_722);
xor U397 (N_397,N_34,N_60);
xor U398 (N_398,N_147,In_365);
nor U399 (N_399,In_303,N_107);
and U400 (N_400,In_149,N_300);
nand U401 (N_401,N_241,N_313);
and U402 (N_402,N_294,N_255);
and U403 (N_403,N_266,N_123);
and U404 (N_404,N_202,N_286);
xor U405 (N_405,N_143,N_227);
nor U406 (N_406,N_267,In_715);
nor U407 (N_407,In_388,N_254);
xnor U408 (N_408,N_296,In_669);
and U409 (N_409,N_263,N_367);
and U410 (N_410,N_354,N_346);
xor U411 (N_411,N_356,N_203);
nor U412 (N_412,In_510,In_520);
xnor U413 (N_413,N_225,In_459);
and U414 (N_414,N_290,N_268);
or U415 (N_415,N_237,N_304);
nand U416 (N_416,N_310,N_119);
xor U417 (N_417,N_396,N_246);
xor U418 (N_418,In_666,In_94);
nand U419 (N_419,In_136,N_309);
nor U420 (N_420,N_218,In_706);
or U421 (N_421,N_261,N_319);
xor U422 (N_422,N_239,N_311);
nor U423 (N_423,N_272,In_456);
or U424 (N_424,N_2,N_377);
xnor U425 (N_425,N_50,N_215);
and U426 (N_426,N_264,In_204);
nand U427 (N_427,N_334,N_231);
nor U428 (N_428,N_360,N_209);
nand U429 (N_429,N_271,N_381);
nand U430 (N_430,In_619,N_397);
nor U431 (N_431,N_207,In_193);
or U432 (N_432,N_328,N_74);
nor U433 (N_433,In_376,N_376);
and U434 (N_434,N_285,N_353);
and U435 (N_435,N_331,N_110);
and U436 (N_436,N_134,In_107);
nand U437 (N_437,In_75,N_238);
nor U438 (N_438,N_369,In_446);
nand U439 (N_439,N_392,N_342);
nand U440 (N_440,N_262,In_634);
nand U441 (N_441,N_180,In_108);
xor U442 (N_442,N_269,N_149);
nor U443 (N_443,N_253,N_361);
or U444 (N_444,N_395,N_248);
and U445 (N_445,In_590,In_694);
nand U446 (N_446,N_213,N_348);
and U447 (N_447,N_305,N_158);
and U448 (N_448,N_250,In_103);
xor U449 (N_449,N_114,In_32);
or U450 (N_450,N_91,N_198);
xnor U451 (N_451,N_233,N_16);
or U452 (N_452,N_194,In_438);
and U453 (N_453,N_273,In_186);
or U454 (N_454,N_111,N_318);
xnor U455 (N_455,N_26,N_355);
or U456 (N_456,N_295,N_365);
or U457 (N_457,N_359,N_299);
xor U458 (N_458,N_120,N_192);
xor U459 (N_459,N_36,N_13);
nor U460 (N_460,N_133,In_628);
or U461 (N_461,N_228,N_223);
or U462 (N_462,N_352,N_384);
and U463 (N_463,In_206,N_67);
nor U464 (N_464,N_53,In_647);
nand U465 (N_465,N_236,N_288);
and U466 (N_466,In_331,N_84);
and U467 (N_467,N_301,N_385);
nand U468 (N_468,In_458,N_260);
xnor U469 (N_469,In_239,N_251);
xnor U470 (N_470,N_350,N_364);
nand U471 (N_471,N_219,N_349);
nor U472 (N_472,In_727,N_181);
and U473 (N_473,In_615,N_217);
or U474 (N_474,N_327,N_389);
nand U475 (N_475,N_338,N_29);
or U476 (N_476,N_362,N_201);
nor U477 (N_477,In_200,In_521);
nand U478 (N_478,In_699,N_224);
and U479 (N_479,In_190,N_297);
and U480 (N_480,N_184,N_230);
and U481 (N_481,N_229,N_183);
nor U482 (N_482,In_1,N_393);
and U483 (N_483,In_257,N_235);
nor U484 (N_484,In_55,In_639);
nand U485 (N_485,In_613,In_78);
xnor U486 (N_486,N_280,N_4);
and U487 (N_487,In_225,N_249);
nand U488 (N_488,N_387,N_368);
and U489 (N_489,N_335,N_337);
nand U490 (N_490,N_122,N_220);
and U491 (N_491,N_19,N_234);
or U492 (N_492,N_345,N_289);
and U493 (N_493,N_344,In_671);
nand U494 (N_494,N_257,N_242);
nor U495 (N_495,N_85,In_128);
or U496 (N_496,N_373,N_140);
xnor U497 (N_497,N_278,N_221);
nor U498 (N_498,N_357,N_1);
or U499 (N_499,N_211,N_214);
nor U500 (N_500,N_341,N_276);
or U501 (N_501,N_366,N_383);
and U502 (N_502,N_394,N_279);
and U503 (N_503,In_472,N_302);
nand U504 (N_504,N_358,N_371);
nor U505 (N_505,N_18,N_31);
nor U506 (N_506,N_148,In_256);
nand U507 (N_507,N_247,N_222);
nand U508 (N_508,In_152,In_641);
nor U509 (N_509,N_205,In_133);
nor U510 (N_510,N_382,N_390);
xor U511 (N_511,N_258,N_117);
nor U512 (N_512,N_306,N_308);
nand U513 (N_513,N_150,In_547);
nand U514 (N_514,N_315,N_284);
nor U515 (N_515,In_173,N_135);
nand U516 (N_516,N_363,N_206);
and U517 (N_517,N_391,N_347);
and U518 (N_518,N_323,N_336);
and U519 (N_519,N_256,In_486);
nand U520 (N_520,In_651,N_339);
or U521 (N_521,In_251,N_226);
nor U522 (N_522,In_219,N_188);
nor U523 (N_523,N_115,N_40);
nor U524 (N_524,N_118,In_196);
nor U525 (N_525,In_745,N_378);
or U526 (N_526,N_333,In_536);
nand U527 (N_527,N_169,N_204);
nand U528 (N_528,N_321,In_220);
nor U529 (N_529,N_277,N_136);
nor U530 (N_530,N_325,N_245);
nor U531 (N_531,N_332,N_386);
or U532 (N_532,N_282,In_443);
nor U533 (N_533,N_293,In_657);
nand U534 (N_534,N_330,N_283);
nand U535 (N_535,N_298,In_180);
nor U536 (N_536,N_244,N_351);
nand U537 (N_537,N_208,N_252);
and U538 (N_538,N_197,In_516);
or U539 (N_539,In_311,In_711);
nand U540 (N_540,N_375,In_272);
nand U541 (N_541,In_505,In_463);
and U542 (N_542,N_126,N_380);
xor U543 (N_543,N_8,In_25);
nor U544 (N_544,N_200,N_270);
and U545 (N_545,N_210,In_328);
nand U546 (N_546,N_216,N_179);
or U547 (N_547,N_388,N_324);
nand U548 (N_548,N_159,In_375);
or U549 (N_549,N_106,In_271);
nor U550 (N_550,In_361,N_343);
and U551 (N_551,N_379,N_195);
nor U552 (N_552,In_655,N_316);
or U553 (N_553,In_350,In_604);
nor U554 (N_554,N_232,N_240);
xnor U555 (N_555,N_326,N_291);
xor U556 (N_556,N_281,N_259);
and U557 (N_557,N_265,In_610);
nand U558 (N_558,N_329,N_398);
nor U559 (N_559,In_252,In_351);
xor U560 (N_560,N_370,In_92);
and U561 (N_561,N_287,In_689);
and U562 (N_562,In_130,N_274);
nor U563 (N_563,In_746,N_374);
and U564 (N_564,N_292,In_713);
and U565 (N_565,N_102,N_275);
xnor U566 (N_566,N_320,In_321);
and U567 (N_567,N_59,N_322);
nor U568 (N_568,N_243,N_212);
and U569 (N_569,N_372,N_399);
or U570 (N_570,N_314,N_340);
nand U571 (N_571,N_312,In_684);
and U572 (N_572,In_121,In_223);
and U573 (N_573,N_307,N_303);
nand U574 (N_574,N_317,In_288);
or U575 (N_575,N_384,In_375);
xor U576 (N_576,N_229,N_396);
or U577 (N_577,N_273,In_634);
xnor U578 (N_578,N_380,N_284);
and U579 (N_579,N_143,In_173);
or U580 (N_580,N_110,N_336);
nand U581 (N_581,N_259,N_318);
nand U582 (N_582,N_324,N_272);
nor U583 (N_583,N_84,N_209);
and U584 (N_584,In_149,N_359);
xnor U585 (N_585,N_283,In_220);
nor U586 (N_586,N_222,N_331);
or U587 (N_587,N_324,N_247);
and U588 (N_588,In_459,N_134);
nor U589 (N_589,In_225,N_288);
nand U590 (N_590,N_261,N_265);
xor U591 (N_591,N_332,N_270);
or U592 (N_592,N_29,N_135);
xor U593 (N_593,N_310,N_179);
nand U594 (N_594,N_26,In_657);
or U595 (N_595,N_245,N_353);
nor U596 (N_596,N_8,In_438);
nand U597 (N_597,N_288,In_55);
or U598 (N_598,N_367,N_286);
and U599 (N_599,N_275,N_221);
and U600 (N_600,N_555,N_562);
or U601 (N_601,N_460,N_465);
nor U602 (N_602,N_581,N_444);
or U603 (N_603,N_407,N_492);
nand U604 (N_604,N_495,N_554);
and U605 (N_605,N_578,N_408);
and U606 (N_606,N_461,N_467);
nor U607 (N_607,N_530,N_450);
or U608 (N_608,N_464,N_511);
or U609 (N_609,N_456,N_587);
nand U610 (N_610,N_412,N_589);
xor U611 (N_611,N_426,N_550);
nor U612 (N_612,N_570,N_519);
nand U613 (N_613,N_590,N_430);
and U614 (N_614,N_505,N_498);
xnor U615 (N_615,N_551,N_537);
nand U616 (N_616,N_538,N_406);
nor U617 (N_617,N_473,N_502);
nor U618 (N_618,N_471,N_575);
xor U619 (N_619,N_453,N_522);
and U620 (N_620,N_496,N_488);
nor U621 (N_621,N_503,N_422);
or U622 (N_622,N_576,N_524);
and U623 (N_623,N_525,N_486);
nor U624 (N_624,N_445,N_415);
and U625 (N_625,N_418,N_501);
or U626 (N_626,N_565,N_588);
or U627 (N_627,N_485,N_404);
nand U628 (N_628,N_535,N_515);
and U629 (N_629,N_596,N_468);
nor U630 (N_630,N_401,N_474);
or U631 (N_631,N_523,N_459);
or U632 (N_632,N_476,N_521);
and U633 (N_633,N_480,N_429);
xnor U634 (N_634,N_574,N_592);
nand U635 (N_635,N_599,N_434);
and U636 (N_636,N_470,N_402);
nor U637 (N_637,N_514,N_543);
nor U638 (N_638,N_403,N_478);
or U639 (N_639,N_499,N_559);
nand U640 (N_640,N_516,N_489);
and U641 (N_641,N_481,N_520);
nand U642 (N_642,N_567,N_506);
nand U643 (N_643,N_424,N_561);
nor U644 (N_644,N_556,N_549);
xnor U645 (N_645,N_457,N_593);
nor U646 (N_646,N_528,N_449);
and U647 (N_647,N_534,N_544);
and U648 (N_648,N_431,N_420);
nand U649 (N_649,N_491,N_440);
nand U650 (N_650,N_583,N_573);
nor U651 (N_651,N_569,N_563);
and U652 (N_652,N_437,N_493);
nor U653 (N_653,N_564,N_597);
nor U654 (N_654,N_446,N_585);
and U655 (N_655,N_423,N_455);
nor U656 (N_656,N_584,N_409);
nand U657 (N_657,N_410,N_405);
and U658 (N_658,N_518,N_414);
nand U659 (N_659,N_508,N_416);
nand U660 (N_660,N_517,N_494);
and U661 (N_661,N_512,N_580);
and U662 (N_662,N_572,N_472);
nand U663 (N_663,N_482,N_432);
and U664 (N_664,N_526,N_500);
or U665 (N_665,N_497,N_463);
and U666 (N_666,N_539,N_490);
nor U667 (N_667,N_504,N_438);
nand U668 (N_668,N_529,N_421);
nand U669 (N_669,N_451,N_542);
or U670 (N_670,N_571,N_413);
nor U671 (N_671,N_479,N_586);
and U672 (N_672,N_532,N_527);
nor U673 (N_673,N_541,N_419);
or U674 (N_674,N_428,N_546);
nand U675 (N_675,N_442,N_487);
nand U676 (N_676,N_441,N_452);
or U677 (N_677,N_568,N_458);
nand U678 (N_678,N_411,N_547);
nand U679 (N_679,N_582,N_531);
and U680 (N_680,N_454,N_469);
nand U681 (N_681,N_536,N_448);
nor U682 (N_682,N_425,N_439);
or U683 (N_683,N_483,N_433);
and U684 (N_684,N_552,N_400);
nand U685 (N_685,N_591,N_466);
nor U686 (N_686,N_477,N_443);
nand U687 (N_687,N_594,N_545);
nor U688 (N_688,N_540,N_553);
nor U689 (N_689,N_595,N_427);
or U690 (N_690,N_447,N_509);
or U691 (N_691,N_507,N_560);
nor U692 (N_692,N_557,N_548);
and U693 (N_693,N_579,N_417);
nand U694 (N_694,N_558,N_598);
and U695 (N_695,N_484,N_513);
or U696 (N_696,N_435,N_577);
or U697 (N_697,N_462,N_475);
nand U698 (N_698,N_510,N_436);
nand U699 (N_699,N_533,N_566);
nor U700 (N_700,N_589,N_485);
nor U701 (N_701,N_584,N_417);
and U702 (N_702,N_550,N_553);
nand U703 (N_703,N_444,N_450);
or U704 (N_704,N_595,N_597);
and U705 (N_705,N_558,N_429);
and U706 (N_706,N_578,N_513);
and U707 (N_707,N_587,N_520);
nand U708 (N_708,N_561,N_566);
nor U709 (N_709,N_478,N_535);
xor U710 (N_710,N_461,N_498);
and U711 (N_711,N_437,N_471);
nand U712 (N_712,N_475,N_448);
nand U713 (N_713,N_428,N_524);
nor U714 (N_714,N_523,N_507);
nand U715 (N_715,N_471,N_482);
or U716 (N_716,N_481,N_418);
and U717 (N_717,N_426,N_598);
nand U718 (N_718,N_537,N_572);
and U719 (N_719,N_441,N_536);
nand U720 (N_720,N_598,N_594);
or U721 (N_721,N_440,N_529);
or U722 (N_722,N_429,N_487);
or U723 (N_723,N_535,N_440);
or U724 (N_724,N_460,N_528);
and U725 (N_725,N_446,N_531);
nand U726 (N_726,N_572,N_569);
nand U727 (N_727,N_594,N_463);
xor U728 (N_728,N_417,N_562);
nand U729 (N_729,N_474,N_420);
nand U730 (N_730,N_559,N_484);
nand U731 (N_731,N_443,N_426);
nand U732 (N_732,N_578,N_495);
nor U733 (N_733,N_431,N_446);
nand U734 (N_734,N_524,N_545);
xor U735 (N_735,N_400,N_446);
xor U736 (N_736,N_427,N_432);
and U737 (N_737,N_459,N_412);
or U738 (N_738,N_520,N_440);
xnor U739 (N_739,N_477,N_524);
nand U740 (N_740,N_517,N_462);
nand U741 (N_741,N_444,N_445);
and U742 (N_742,N_527,N_545);
or U743 (N_743,N_596,N_592);
xnor U744 (N_744,N_521,N_518);
or U745 (N_745,N_545,N_546);
xor U746 (N_746,N_533,N_590);
nand U747 (N_747,N_568,N_539);
nand U748 (N_748,N_461,N_597);
and U749 (N_749,N_549,N_541);
and U750 (N_750,N_553,N_569);
nand U751 (N_751,N_518,N_524);
xor U752 (N_752,N_598,N_565);
or U753 (N_753,N_522,N_466);
nor U754 (N_754,N_441,N_447);
xnor U755 (N_755,N_569,N_593);
or U756 (N_756,N_449,N_582);
nand U757 (N_757,N_534,N_445);
nand U758 (N_758,N_485,N_549);
nor U759 (N_759,N_516,N_460);
and U760 (N_760,N_493,N_411);
nor U761 (N_761,N_563,N_559);
nand U762 (N_762,N_588,N_447);
nand U763 (N_763,N_443,N_576);
or U764 (N_764,N_423,N_542);
or U765 (N_765,N_583,N_562);
or U766 (N_766,N_413,N_453);
nand U767 (N_767,N_599,N_431);
nor U768 (N_768,N_505,N_440);
or U769 (N_769,N_597,N_535);
xnor U770 (N_770,N_444,N_427);
xor U771 (N_771,N_410,N_474);
nor U772 (N_772,N_536,N_412);
or U773 (N_773,N_459,N_507);
and U774 (N_774,N_478,N_524);
and U775 (N_775,N_421,N_560);
nand U776 (N_776,N_535,N_561);
and U777 (N_777,N_561,N_558);
nand U778 (N_778,N_561,N_505);
nor U779 (N_779,N_547,N_457);
nand U780 (N_780,N_406,N_493);
or U781 (N_781,N_467,N_443);
nand U782 (N_782,N_531,N_533);
xnor U783 (N_783,N_468,N_436);
or U784 (N_784,N_566,N_427);
and U785 (N_785,N_422,N_517);
nor U786 (N_786,N_564,N_521);
nand U787 (N_787,N_593,N_475);
or U788 (N_788,N_567,N_469);
xor U789 (N_789,N_404,N_590);
or U790 (N_790,N_569,N_442);
nor U791 (N_791,N_443,N_556);
nor U792 (N_792,N_453,N_428);
nor U793 (N_793,N_467,N_421);
and U794 (N_794,N_570,N_486);
and U795 (N_795,N_428,N_411);
and U796 (N_796,N_431,N_528);
xnor U797 (N_797,N_541,N_410);
xnor U798 (N_798,N_495,N_492);
and U799 (N_799,N_428,N_492);
nor U800 (N_800,N_784,N_764);
or U801 (N_801,N_617,N_611);
and U802 (N_802,N_604,N_769);
and U803 (N_803,N_733,N_762);
nor U804 (N_804,N_686,N_630);
nor U805 (N_805,N_696,N_745);
xor U806 (N_806,N_632,N_777);
nand U807 (N_807,N_736,N_662);
or U808 (N_808,N_609,N_712);
and U809 (N_809,N_602,N_759);
nor U810 (N_810,N_658,N_657);
or U811 (N_811,N_795,N_684);
nor U812 (N_812,N_616,N_688);
and U813 (N_813,N_625,N_739);
xnor U814 (N_814,N_787,N_664);
nand U815 (N_815,N_678,N_797);
and U816 (N_816,N_674,N_750);
and U817 (N_817,N_633,N_610);
nand U818 (N_818,N_744,N_668);
and U819 (N_819,N_785,N_707);
and U820 (N_820,N_786,N_773);
and U821 (N_821,N_730,N_715);
or U822 (N_822,N_644,N_791);
nand U823 (N_823,N_685,N_605);
and U824 (N_824,N_734,N_702);
and U825 (N_825,N_725,N_789);
nand U826 (N_826,N_613,N_695);
nor U827 (N_827,N_722,N_758);
and U828 (N_828,N_755,N_672);
xnor U829 (N_829,N_682,N_631);
or U830 (N_830,N_689,N_681);
or U831 (N_831,N_727,N_746);
nor U832 (N_832,N_623,N_651);
and U833 (N_833,N_723,N_629);
or U834 (N_834,N_737,N_765);
nor U835 (N_835,N_792,N_783);
nor U836 (N_836,N_772,N_661);
nor U837 (N_837,N_635,N_788);
or U838 (N_838,N_781,N_705);
and U839 (N_839,N_692,N_771);
xnor U840 (N_840,N_710,N_694);
or U841 (N_841,N_697,N_753);
or U842 (N_842,N_768,N_763);
nand U843 (N_843,N_646,N_760);
nor U844 (N_844,N_700,N_726);
nand U845 (N_845,N_680,N_667);
or U846 (N_846,N_603,N_738);
and U847 (N_847,N_647,N_756);
nor U848 (N_848,N_641,N_708);
xor U849 (N_849,N_648,N_751);
and U850 (N_850,N_743,N_780);
or U851 (N_851,N_655,N_676);
nand U852 (N_852,N_634,N_652);
nand U853 (N_853,N_754,N_636);
and U854 (N_854,N_615,N_677);
nor U855 (N_855,N_770,N_628);
xnor U856 (N_856,N_683,N_671);
or U857 (N_857,N_794,N_701);
nor U858 (N_858,N_721,N_637);
nor U859 (N_859,N_711,N_600);
and U860 (N_860,N_608,N_698);
or U861 (N_861,N_690,N_741);
and U862 (N_862,N_621,N_638);
nor U863 (N_863,N_618,N_757);
and U864 (N_864,N_656,N_767);
xnor U865 (N_865,N_714,N_706);
nor U866 (N_866,N_673,N_776);
xor U867 (N_867,N_717,N_642);
or U868 (N_868,N_660,N_649);
nor U869 (N_869,N_670,N_793);
xor U870 (N_870,N_622,N_798);
nand U871 (N_871,N_752,N_687);
nand U872 (N_872,N_669,N_747);
nand U873 (N_873,N_650,N_729);
nor U874 (N_874,N_704,N_620);
nand U875 (N_875,N_612,N_774);
nand U876 (N_876,N_748,N_766);
or U877 (N_877,N_679,N_790);
and U878 (N_878,N_693,N_699);
xor U879 (N_879,N_675,N_779);
or U880 (N_880,N_713,N_735);
nand U881 (N_881,N_639,N_716);
nor U882 (N_882,N_659,N_643);
or U883 (N_883,N_719,N_601);
and U884 (N_884,N_645,N_703);
nand U885 (N_885,N_626,N_665);
or U886 (N_886,N_782,N_663);
or U887 (N_887,N_799,N_640);
nand U888 (N_888,N_761,N_606);
or U889 (N_889,N_728,N_742);
or U890 (N_890,N_624,N_666);
or U891 (N_891,N_775,N_718);
nor U892 (N_892,N_607,N_720);
and U893 (N_893,N_731,N_627);
nand U894 (N_894,N_619,N_614);
and U895 (N_895,N_732,N_709);
nor U896 (N_896,N_796,N_691);
or U897 (N_897,N_724,N_749);
or U898 (N_898,N_653,N_654);
or U899 (N_899,N_778,N_740);
and U900 (N_900,N_718,N_660);
or U901 (N_901,N_606,N_645);
nor U902 (N_902,N_652,N_657);
or U903 (N_903,N_796,N_620);
nor U904 (N_904,N_690,N_712);
and U905 (N_905,N_645,N_789);
and U906 (N_906,N_771,N_734);
or U907 (N_907,N_799,N_673);
or U908 (N_908,N_674,N_616);
nor U909 (N_909,N_693,N_687);
xnor U910 (N_910,N_633,N_753);
or U911 (N_911,N_632,N_700);
nor U912 (N_912,N_652,N_731);
and U913 (N_913,N_752,N_753);
or U914 (N_914,N_741,N_719);
nor U915 (N_915,N_744,N_636);
nor U916 (N_916,N_705,N_772);
nor U917 (N_917,N_604,N_723);
xor U918 (N_918,N_797,N_732);
and U919 (N_919,N_655,N_648);
nor U920 (N_920,N_614,N_637);
or U921 (N_921,N_765,N_607);
nor U922 (N_922,N_761,N_603);
nand U923 (N_923,N_789,N_717);
or U924 (N_924,N_761,N_727);
and U925 (N_925,N_726,N_732);
or U926 (N_926,N_730,N_774);
and U927 (N_927,N_613,N_629);
nor U928 (N_928,N_604,N_797);
xnor U929 (N_929,N_741,N_632);
nand U930 (N_930,N_791,N_731);
or U931 (N_931,N_623,N_721);
nand U932 (N_932,N_787,N_645);
nor U933 (N_933,N_776,N_785);
and U934 (N_934,N_669,N_640);
nor U935 (N_935,N_751,N_649);
and U936 (N_936,N_655,N_769);
nand U937 (N_937,N_785,N_770);
xor U938 (N_938,N_657,N_777);
nor U939 (N_939,N_688,N_767);
nand U940 (N_940,N_609,N_734);
nor U941 (N_941,N_633,N_671);
nor U942 (N_942,N_618,N_669);
nand U943 (N_943,N_784,N_773);
nand U944 (N_944,N_799,N_657);
or U945 (N_945,N_732,N_628);
nand U946 (N_946,N_651,N_693);
nand U947 (N_947,N_637,N_655);
xnor U948 (N_948,N_699,N_666);
or U949 (N_949,N_711,N_731);
and U950 (N_950,N_667,N_677);
nor U951 (N_951,N_633,N_687);
and U952 (N_952,N_636,N_705);
xnor U953 (N_953,N_687,N_759);
or U954 (N_954,N_715,N_635);
and U955 (N_955,N_767,N_787);
nor U956 (N_956,N_610,N_635);
nor U957 (N_957,N_649,N_617);
xor U958 (N_958,N_776,N_638);
and U959 (N_959,N_674,N_665);
xnor U960 (N_960,N_650,N_631);
and U961 (N_961,N_775,N_725);
or U962 (N_962,N_713,N_646);
nand U963 (N_963,N_689,N_685);
and U964 (N_964,N_708,N_784);
nand U965 (N_965,N_729,N_752);
xnor U966 (N_966,N_604,N_607);
or U967 (N_967,N_759,N_751);
or U968 (N_968,N_649,N_671);
nor U969 (N_969,N_632,N_780);
nand U970 (N_970,N_625,N_708);
nand U971 (N_971,N_669,N_628);
or U972 (N_972,N_609,N_702);
nand U973 (N_973,N_625,N_628);
nor U974 (N_974,N_726,N_743);
and U975 (N_975,N_670,N_786);
nor U976 (N_976,N_798,N_643);
or U977 (N_977,N_627,N_680);
and U978 (N_978,N_642,N_613);
nor U979 (N_979,N_788,N_638);
and U980 (N_980,N_673,N_782);
or U981 (N_981,N_708,N_622);
nor U982 (N_982,N_644,N_637);
or U983 (N_983,N_797,N_708);
nor U984 (N_984,N_607,N_778);
nand U985 (N_985,N_758,N_738);
nor U986 (N_986,N_601,N_706);
and U987 (N_987,N_770,N_711);
xor U988 (N_988,N_736,N_786);
and U989 (N_989,N_725,N_776);
nor U990 (N_990,N_762,N_739);
and U991 (N_991,N_725,N_631);
nand U992 (N_992,N_751,N_796);
nor U993 (N_993,N_712,N_608);
nor U994 (N_994,N_762,N_763);
nor U995 (N_995,N_646,N_687);
nor U996 (N_996,N_702,N_684);
nand U997 (N_997,N_766,N_749);
nor U998 (N_998,N_610,N_636);
and U999 (N_999,N_782,N_622);
nand U1000 (N_1000,N_820,N_870);
nand U1001 (N_1001,N_919,N_909);
and U1002 (N_1002,N_997,N_889);
and U1003 (N_1003,N_935,N_969);
or U1004 (N_1004,N_973,N_960);
nand U1005 (N_1005,N_983,N_926);
nand U1006 (N_1006,N_892,N_873);
and U1007 (N_1007,N_976,N_970);
xnor U1008 (N_1008,N_962,N_925);
nor U1009 (N_1009,N_989,N_972);
and U1010 (N_1010,N_884,N_936);
xor U1011 (N_1011,N_805,N_860);
xor U1012 (N_1012,N_918,N_880);
nor U1013 (N_1013,N_982,N_941);
or U1014 (N_1014,N_816,N_928);
nand U1015 (N_1015,N_888,N_874);
or U1016 (N_1016,N_806,N_859);
and U1017 (N_1017,N_900,N_869);
or U1018 (N_1018,N_971,N_887);
nand U1019 (N_1019,N_848,N_836);
and U1020 (N_1020,N_804,N_975);
nand U1021 (N_1021,N_824,N_908);
nand U1022 (N_1022,N_837,N_871);
nand U1023 (N_1023,N_966,N_951);
nor U1024 (N_1024,N_904,N_952);
and U1025 (N_1025,N_930,N_977);
nand U1026 (N_1026,N_854,N_886);
or U1027 (N_1027,N_921,N_986);
nand U1028 (N_1028,N_979,N_839);
and U1029 (N_1029,N_939,N_841);
and U1030 (N_1030,N_835,N_963);
nand U1031 (N_1031,N_993,N_846);
or U1032 (N_1032,N_883,N_980);
and U1033 (N_1033,N_810,N_920);
nor U1034 (N_1034,N_948,N_853);
and U1035 (N_1035,N_834,N_898);
nor U1036 (N_1036,N_857,N_821);
and U1037 (N_1037,N_876,N_801);
and U1038 (N_1038,N_855,N_851);
nand U1039 (N_1039,N_897,N_800);
nand U1040 (N_1040,N_812,N_863);
nand U1041 (N_1041,N_831,N_894);
nor U1042 (N_1042,N_856,N_917);
nor U1043 (N_1043,N_866,N_809);
nor U1044 (N_1044,N_845,N_872);
and U1045 (N_1045,N_890,N_944);
nand U1046 (N_1046,N_956,N_912);
nand U1047 (N_1047,N_877,N_838);
nor U1048 (N_1048,N_961,N_907);
nor U1049 (N_1049,N_814,N_885);
or U1050 (N_1050,N_847,N_955);
or U1051 (N_1051,N_942,N_929);
nand U1052 (N_1052,N_899,N_865);
nor U1053 (N_1053,N_861,N_945);
nor U1054 (N_1054,N_832,N_818);
nand U1055 (N_1055,N_896,N_862);
xnor U1056 (N_1056,N_867,N_826);
nand U1057 (N_1057,N_957,N_813);
nor U1058 (N_1058,N_910,N_881);
nand U1059 (N_1059,N_913,N_827);
nor U1060 (N_1060,N_879,N_927);
nor U1061 (N_1061,N_998,N_947);
nand U1062 (N_1062,N_934,N_891);
nand U1063 (N_1063,N_996,N_985);
nand U1064 (N_1064,N_931,N_893);
nand U1065 (N_1065,N_829,N_882);
and U1066 (N_1066,N_840,N_923);
xnor U1067 (N_1067,N_906,N_938);
and U1068 (N_1068,N_808,N_833);
nor U1069 (N_1069,N_995,N_825);
nand U1070 (N_1070,N_822,N_950);
and U1071 (N_1071,N_815,N_850);
xor U1072 (N_1072,N_864,N_987);
nor U1073 (N_1073,N_940,N_954);
xnor U1074 (N_1074,N_878,N_968);
and U1075 (N_1075,N_807,N_965);
xor U1076 (N_1076,N_858,N_914);
or U1077 (N_1077,N_828,N_984);
and U1078 (N_1078,N_990,N_903);
and U1079 (N_1079,N_974,N_922);
and U1080 (N_1080,N_978,N_844);
and U1081 (N_1081,N_819,N_823);
and U1082 (N_1082,N_946,N_959);
xor U1083 (N_1083,N_994,N_915);
or U1084 (N_1084,N_988,N_811);
and U1085 (N_1085,N_902,N_911);
nor U1086 (N_1086,N_933,N_964);
and U1087 (N_1087,N_895,N_916);
xor U1088 (N_1088,N_981,N_852);
nor U1089 (N_1089,N_958,N_843);
nand U1090 (N_1090,N_949,N_924);
nor U1091 (N_1091,N_932,N_817);
and U1092 (N_1092,N_999,N_901);
or U1093 (N_1093,N_849,N_992);
xnor U1094 (N_1094,N_937,N_868);
nand U1095 (N_1095,N_943,N_842);
or U1096 (N_1096,N_953,N_803);
nand U1097 (N_1097,N_905,N_830);
nand U1098 (N_1098,N_802,N_875);
or U1099 (N_1099,N_991,N_967);
and U1100 (N_1100,N_949,N_844);
and U1101 (N_1101,N_945,N_839);
xnor U1102 (N_1102,N_830,N_933);
nor U1103 (N_1103,N_876,N_807);
or U1104 (N_1104,N_928,N_901);
xnor U1105 (N_1105,N_832,N_976);
nor U1106 (N_1106,N_927,N_942);
and U1107 (N_1107,N_910,N_899);
xor U1108 (N_1108,N_805,N_972);
nand U1109 (N_1109,N_982,N_811);
nand U1110 (N_1110,N_847,N_822);
or U1111 (N_1111,N_870,N_906);
nand U1112 (N_1112,N_919,N_869);
and U1113 (N_1113,N_872,N_971);
xor U1114 (N_1114,N_983,N_921);
nor U1115 (N_1115,N_964,N_829);
xnor U1116 (N_1116,N_859,N_861);
nor U1117 (N_1117,N_856,N_833);
nor U1118 (N_1118,N_824,N_910);
or U1119 (N_1119,N_969,N_857);
nand U1120 (N_1120,N_959,N_928);
or U1121 (N_1121,N_855,N_846);
nand U1122 (N_1122,N_982,N_990);
or U1123 (N_1123,N_823,N_896);
xnor U1124 (N_1124,N_989,N_980);
and U1125 (N_1125,N_926,N_957);
nand U1126 (N_1126,N_997,N_948);
xnor U1127 (N_1127,N_979,N_971);
nor U1128 (N_1128,N_873,N_953);
and U1129 (N_1129,N_938,N_814);
xnor U1130 (N_1130,N_902,N_984);
nand U1131 (N_1131,N_969,N_915);
nor U1132 (N_1132,N_930,N_861);
xor U1133 (N_1133,N_874,N_895);
and U1134 (N_1134,N_806,N_842);
xor U1135 (N_1135,N_971,N_869);
nor U1136 (N_1136,N_921,N_932);
or U1137 (N_1137,N_884,N_972);
nor U1138 (N_1138,N_942,N_985);
nor U1139 (N_1139,N_976,N_900);
or U1140 (N_1140,N_966,N_866);
nor U1141 (N_1141,N_932,N_977);
and U1142 (N_1142,N_935,N_905);
and U1143 (N_1143,N_915,N_931);
nor U1144 (N_1144,N_961,N_994);
nor U1145 (N_1145,N_829,N_904);
nand U1146 (N_1146,N_964,N_969);
nand U1147 (N_1147,N_823,N_831);
nor U1148 (N_1148,N_965,N_804);
nor U1149 (N_1149,N_986,N_895);
nor U1150 (N_1150,N_807,N_822);
nand U1151 (N_1151,N_892,N_910);
nor U1152 (N_1152,N_991,N_810);
nor U1153 (N_1153,N_957,N_903);
and U1154 (N_1154,N_997,N_960);
nor U1155 (N_1155,N_927,N_933);
xor U1156 (N_1156,N_924,N_972);
nand U1157 (N_1157,N_875,N_822);
and U1158 (N_1158,N_812,N_967);
xor U1159 (N_1159,N_907,N_821);
nor U1160 (N_1160,N_965,N_819);
nand U1161 (N_1161,N_924,N_879);
or U1162 (N_1162,N_921,N_950);
xor U1163 (N_1163,N_976,N_991);
and U1164 (N_1164,N_997,N_800);
nand U1165 (N_1165,N_819,N_891);
and U1166 (N_1166,N_997,N_963);
and U1167 (N_1167,N_952,N_941);
and U1168 (N_1168,N_825,N_866);
or U1169 (N_1169,N_834,N_800);
and U1170 (N_1170,N_998,N_912);
xor U1171 (N_1171,N_964,N_851);
nor U1172 (N_1172,N_894,N_912);
or U1173 (N_1173,N_838,N_806);
nand U1174 (N_1174,N_877,N_889);
xnor U1175 (N_1175,N_988,N_986);
nor U1176 (N_1176,N_901,N_937);
and U1177 (N_1177,N_886,N_835);
or U1178 (N_1178,N_983,N_933);
nand U1179 (N_1179,N_874,N_991);
xnor U1180 (N_1180,N_869,N_991);
nand U1181 (N_1181,N_847,N_989);
or U1182 (N_1182,N_838,N_978);
and U1183 (N_1183,N_845,N_828);
nor U1184 (N_1184,N_837,N_987);
nor U1185 (N_1185,N_823,N_984);
nor U1186 (N_1186,N_850,N_830);
or U1187 (N_1187,N_951,N_897);
or U1188 (N_1188,N_886,N_814);
or U1189 (N_1189,N_942,N_988);
nor U1190 (N_1190,N_874,N_814);
nor U1191 (N_1191,N_892,N_961);
and U1192 (N_1192,N_979,N_939);
and U1193 (N_1193,N_826,N_856);
or U1194 (N_1194,N_804,N_973);
nor U1195 (N_1195,N_974,N_835);
or U1196 (N_1196,N_956,N_812);
nor U1197 (N_1197,N_906,N_847);
or U1198 (N_1198,N_944,N_989);
xor U1199 (N_1199,N_825,N_877);
nand U1200 (N_1200,N_1176,N_1166);
nand U1201 (N_1201,N_1184,N_1119);
xor U1202 (N_1202,N_1060,N_1015);
or U1203 (N_1203,N_1181,N_1000);
and U1204 (N_1204,N_1037,N_1138);
or U1205 (N_1205,N_1073,N_1081);
and U1206 (N_1206,N_1038,N_1159);
and U1207 (N_1207,N_1121,N_1017);
nand U1208 (N_1208,N_1160,N_1144);
and U1209 (N_1209,N_1141,N_1100);
or U1210 (N_1210,N_1168,N_1045);
nor U1211 (N_1211,N_1173,N_1088);
nor U1212 (N_1212,N_1078,N_1114);
nand U1213 (N_1213,N_1182,N_1116);
and U1214 (N_1214,N_1006,N_1190);
nand U1215 (N_1215,N_1009,N_1199);
nand U1216 (N_1216,N_1158,N_1193);
nand U1217 (N_1217,N_1064,N_1062);
nor U1218 (N_1218,N_1174,N_1059);
or U1219 (N_1219,N_1150,N_1093);
and U1220 (N_1220,N_1031,N_1192);
and U1221 (N_1221,N_1113,N_1186);
nand U1222 (N_1222,N_1033,N_1044);
nor U1223 (N_1223,N_1165,N_1147);
nand U1224 (N_1224,N_1110,N_1101);
or U1225 (N_1225,N_1012,N_1066);
and U1226 (N_1226,N_1051,N_1154);
xor U1227 (N_1227,N_1097,N_1122);
nand U1228 (N_1228,N_1002,N_1030);
nand U1229 (N_1229,N_1067,N_1068);
nand U1230 (N_1230,N_1195,N_1071);
nand U1231 (N_1231,N_1089,N_1130);
xnor U1232 (N_1232,N_1055,N_1126);
nand U1233 (N_1233,N_1198,N_1143);
or U1234 (N_1234,N_1058,N_1180);
or U1235 (N_1235,N_1028,N_1145);
nand U1236 (N_1236,N_1169,N_1133);
nand U1237 (N_1237,N_1061,N_1164);
nor U1238 (N_1238,N_1065,N_1079);
nor U1239 (N_1239,N_1083,N_1135);
and U1240 (N_1240,N_1170,N_1098);
nand U1241 (N_1241,N_1011,N_1027);
nand U1242 (N_1242,N_1085,N_1106);
xnor U1243 (N_1243,N_1082,N_1148);
or U1244 (N_1244,N_1023,N_1105);
or U1245 (N_1245,N_1022,N_1157);
and U1246 (N_1246,N_1032,N_1125);
xnor U1247 (N_1247,N_1139,N_1131);
and U1248 (N_1248,N_1096,N_1043);
nor U1249 (N_1249,N_1189,N_1053);
nand U1250 (N_1250,N_1137,N_1172);
and U1251 (N_1251,N_1003,N_1124);
or U1252 (N_1252,N_1140,N_1013);
or U1253 (N_1253,N_1099,N_1036);
or U1254 (N_1254,N_1161,N_1018);
or U1255 (N_1255,N_1049,N_1054);
nand U1256 (N_1256,N_1103,N_1149);
nand U1257 (N_1257,N_1109,N_1048);
or U1258 (N_1258,N_1152,N_1151);
nor U1259 (N_1259,N_1041,N_1118);
or U1260 (N_1260,N_1040,N_1026);
nor U1261 (N_1261,N_1084,N_1004);
or U1262 (N_1262,N_1178,N_1086);
nor U1263 (N_1263,N_1175,N_1029);
nor U1264 (N_1264,N_1162,N_1142);
nor U1265 (N_1265,N_1123,N_1102);
or U1266 (N_1266,N_1008,N_1171);
nand U1267 (N_1267,N_1196,N_1034);
nand U1268 (N_1268,N_1127,N_1024);
nor U1269 (N_1269,N_1146,N_1197);
nand U1270 (N_1270,N_1128,N_1115);
nor U1271 (N_1271,N_1194,N_1187);
and U1272 (N_1272,N_1108,N_1156);
nand U1273 (N_1273,N_1179,N_1076);
nand U1274 (N_1274,N_1177,N_1001);
nor U1275 (N_1275,N_1090,N_1070);
nand U1276 (N_1276,N_1075,N_1163);
nand U1277 (N_1277,N_1072,N_1167);
and U1278 (N_1278,N_1183,N_1050);
nand U1279 (N_1279,N_1052,N_1107);
xor U1280 (N_1280,N_1134,N_1111);
or U1281 (N_1281,N_1132,N_1025);
or U1282 (N_1282,N_1091,N_1035);
or U1283 (N_1283,N_1010,N_1063);
or U1284 (N_1284,N_1019,N_1005);
xnor U1285 (N_1285,N_1112,N_1042);
nor U1286 (N_1286,N_1020,N_1117);
or U1287 (N_1287,N_1007,N_1074);
or U1288 (N_1288,N_1057,N_1136);
or U1289 (N_1289,N_1080,N_1021);
or U1290 (N_1290,N_1092,N_1016);
and U1291 (N_1291,N_1155,N_1094);
or U1292 (N_1292,N_1047,N_1191);
or U1293 (N_1293,N_1014,N_1046);
and U1294 (N_1294,N_1120,N_1087);
and U1295 (N_1295,N_1188,N_1095);
and U1296 (N_1296,N_1185,N_1077);
and U1297 (N_1297,N_1039,N_1153);
nor U1298 (N_1298,N_1129,N_1104);
and U1299 (N_1299,N_1069,N_1056);
nand U1300 (N_1300,N_1138,N_1083);
nor U1301 (N_1301,N_1011,N_1048);
or U1302 (N_1302,N_1134,N_1178);
nand U1303 (N_1303,N_1113,N_1037);
or U1304 (N_1304,N_1086,N_1032);
and U1305 (N_1305,N_1033,N_1092);
or U1306 (N_1306,N_1069,N_1125);
and U1307 (N_1307,N_1080,N_1017);
nand U1308 (N_1308,N_1188,N_1156);
or U1309 (N_1309,N_1101,N_1043);
nor U1310 (N_1310,N_1151,N_1159);
xnor U1311 (N_1311,N_1039,N_1187);
nor U1312 (N_1312,N_1192,N_1052);
nand U1313 (N_1313,N_1036,N_1110);
nand U1314 (N_1314,N_1086,N_1016);
nand U1315 (N_1315,N_1196,N_1073);
nor U1316 (N_1316,N_1074,N_1122);
and U1317 (N_1317,N_1053,N_1124);
nand U1318 (N_1318,N_1016,N_1104);
and U1319 (N_1319,N_1123,N_1146);
nand U1320 (N_1320,N_1118,N_1028);
or U1321 (N_1321,N_1119,N_1140);
or U1322 (N_1322,N_1124,N_1102);
and U1323 (N_1323,N_1077,N_1067);
and U1324 (N_1324,N_1157,N_1152);
xnor U1325 (N_1325,N_1077,N_1156);
and U1326 (N_1326,N_1026,N_1162);
nand U1327 (N_1327,N_1044,N_1103);
nand U1328 (N_1328,N_1179,N_1023);
nand U1329 (N_1329,N_1180,N_1051);
nor U1330 (N_1330,N_1028,N_1033);
xor U1331 (N_1331,N_1182,N_1090);
and U1332 (N_1332,N_1192,N_1168);
or U1333 (N_1333,N_1008,N_1007);
or U1334 (N_1334,N_1082,N_1008);
nor U1335 (N_1335,N_1131,N_1140);
nor U1336 (N_1336,N_1193,N_1119);
and U1337 (N_1337,N_1062,N_1038);
and U1338 (N_1338,N_1068,N_1069);
and U1339 (N_1339,N_1000,N_1166);
nand U1340 (N_1340,N_1042,N_1181);
and U1341 (N_1341,N_1003,N_1062);
and U1342 (N_1342,N_1122,N_1102);
and U1343 (N_1343,N_1161,N_1033);
or U1344 (N_1344,N_1126,N_1175);
nand U1345 (N_1345,N_1063,N_1021);
and U1346 (N_1346,N_1022,N_1146);
or U1347 (N_1347,N_1156,N_1074);
xor U1348 (N_1348,N_1084,N_1134);
or U1349 (N_1349,N_1191,N_1006);
and U1350 (N_1350,N_1056,N_1086);
nor U1351 (N_1351,N_1058,N_1028);
xnor U1352 (N_1352,N_1047,N_1166);
nand U1353 (N_1353,N_1179,N_1084);
nand U1354 (N_1354,N_1020,N_1127);
nand U1355 (N_1355,N_1148,N_1111);
or U1356 (N_1356,N_1087,N_1000);
or U1357 (N_1357,N_1057,N_1159);
and U1358 (N_1358,N_1110,N_1015);
xnor U1359 (N_1359,N_1021,N_1082);
nand U1360 (N_1360,N_1126,N_1084);
xnor U1361 (N_1361,N_1060,N_1148);
and U1362 (N_1362,N_1175,N_1006);
nor U1363 (N_1363,N_1082,N_1101);
or U1364 (N_1364,N_1124,N_1031);
nand U1365 (N_1365,N_1062,N_1155);
and U1366 (N_1366,N_1079,N_1078);
nor U1367 (N_1367,N_1185,N_1000);
and U1368 (N_1368,N_1131,N_1009);
and U1369 (N_1369,N_1135,N_1122);
nand U1370 (N_1370,N_1191,N_1090);
or U1371 (N_1371,N_1195,N_1110);
nand U1372 (N_1372,N_1038,N_1168);
or U1373 (N_1373,N_1092,N_1005);
nand U1374 (N_1374,N_1032,N_1043);
or U1375 (N_1375,N_1146,N_1158);
and U1376 (N_1376,N_1085,N_1071);
xor U1377 (N_1377,N_1137,N_1099);
or U1378 (N_1378,N_1182,N_1098);
or U1379 (N_1379,N_1048,N_1045);
or U1380 (N_1380,N_1067,N_1132);
nor U1381 (N_1381,N_1121,N_1061);
or U1382 (N_1382,N_1131,N_1095);
or U1383 (N_1383,N_1112,N_1051);
and U1384 (N_1384,N_1059,N_1000);
or U1385 (N_1385,N_1116,N_1102);
and U1386 (N_1386,N_1115,N_1168);
nor U1387 (N_1387,N_1076,N_1159);
and U1388 (N_1388,N_1072,N_1052);
and U1389 (N_1389,N_1189,N_1175);
or U1390 (N_1390,N_1037,N_1137);
nor U1391 (N_1391,N_1079,N_1034);
or U1392 (N_1392,N_1038,N_1198);
or U1393 (N_1393,N_1120,N_1191);
and U1394 (N_1394,N_1021,N_1015);
and U1395 (N_1395,N_1025,N_1018);
or U1396 (N_1396,N_1024,N_1025);
nor U1397 (N_1397,N_1072,N_1068);
nor U1398 (N_1398,N_1035,N_1044);
nor U1399 (N_1399,N_1153,N_1058);
nand U1400 (N_1400,N_1262,N_1306);
and U1401 (N_1401,N_1378,N_1261);
or U1402 (N_1402,N_1204,N_1309);
nand U1403 (N_1403,N_1252,N_1342);
and U1404 (N_1404,N_1275,N_1379);
nor U1405 (N_1405,N_1200,N_1277);
xnor U1406 (N_1406,N_1303,N_1373);
nor U1407 (N_1407,N_1238,N_1335);
or U1408 (N_1408,N_1233,N_1307);
and U1409 (N_1409,N_1302,N_1214);
and U1410 (N_1410,N_1241,N_1232);
nor U1411 (N_1411,N_1208,N_1237);
and U1412 (N_1412,N_1380,N_1301);
nand U1413 (N_1413,N_1210,N_1231);
and U1414 (N_1414,N_1257,N_1329);
or U1415 (N_1415,N_1256,N_1315);
or U1416 (N_1416,N_1202,N_1247);
or U1417 (N_1417,N_1212,N_1345);
xor U1418 (N_1418,N_1254,N_1226);
nand U1419 (N_1419,N_1331,N_1205);
and U1420 (N_1420,N_1300,N_1398);
nor U1421 (N_1421,N_1221,N_1328);
and U1422 (N_1422,N_1295,N_1340);
and U1423 (N_1423,N_1381,N_1370);
and U1424 (N_1424,N_1230,N_1351);
or U1425 (N_1425,N_1339,N_1293);
or U1426 (N_1426,N_1269,N_1222);
and U1427 (N_1427,N_1282,N_1228);
nand U1428 (N_1428,N_1227,N_1397);
nor U1429 (N_1429,N_1350,N_1244);
or U1430 (N_1430,N_1362,N_1366);
and U1431 (N_1431,N_1292,N_1368);
and U1432 (N_1432,N_1258,N_1286);
or U1433 (N_1433,N_1201,N_1251);
nor U1434 (N_1434,N_1217,N_1296);
and U1435 (N_1435,N_1326,N_1384);
xnor U1436 (N_1436,N_1325,N_1203);
or U1437 (N_1437,N_1278,N_1213);
nor U1438 (N_1438,N_1284,N_1280);
nand U1439 (N_1439,N_1347,N_1312);
nand U1440 (N_1440,N_1291,N_1388);
nor U1441 (N_1441,N_1255,N_1240);
and U1442 (N_1442,N_1394,N_1246);
nor U1443 (N_1443,N_1338,N_1389);
xor U1444 (N_1444,N_1316,N_1356);
nor U1445 (N_1445,N_1390,N_1290);
nand U1446 (N_1446,N_1317,N_1359);
nand U1447 (N_1447,N_1371,N_1383);
nor U1448 (N_1448,N_1206,N_1245);
or U1449 (N_1449,N_1321,N_1341);
nand U1450 (N_1450,N_1313,N_1288);
and U1451 (N_1451,N_1330,N_1357);
nand U1452 (N_1452,N_1333,N_1376);
xnor U1453 (N_1453,N_1248,N_1259);
nand U1454 (N_1454,N_1395,N_1386);
nand U1455 (N_1455,N_1216,N_1385);
xnor U1456 (N_1456,N_1391,N_1322);
nor U1457 (N_1457,N_1314,N_1294);
nor U1458 (N_1458,N_1365,N_1318);
nand U1459 (N_1459,N_1234,N_1229);
and U1460 (N_1460,N_1285,N_1355);
and U1461 (N_1461,N_1207,N_1346);
and U1462 (N_1462,N_1297,N_1353);
nor U1463 (N_1463,N_1396,N_1249);
nor U1464 (N_1464,N_1224,N_1264);
xor U1465 (N_1465,N_1393,N_1250);
or U1466 (N_1466,N_1283,N_1289);
or U1467 (N_1467,N_1253,N_1361);
xor U1468 (N_1468,N_1265,N_1358);
nor U1469 (N_1469,N_1235,N_1375);
nand U1470 (N_1470,N_1334,N_1219);
nor U1471 (N_1471,N_1272,N_1374);
and U1472 (N_1472,N_1363,N_1319);
and U1473 (N_1473,N_1281,N_1268);
xor U1474 (N_1474,N_1364,N_1360);
or U1475 (N_1475,N_1276,N_1260);
and U1476 (N_1476,N_1299,N_1266);
or U1477 (N_1477,N_1223,N_1323);
nor U1478 (N_1478,N_1337,N_1336);
or U1479 (N_1479,N_1311,N_1399);
nand U1480 (N_1480,N_1369,N_1287);
and U1481 (N_1481,N_1382,N_1270);
xor U1482 (N_1482,N_1377,N_1305);
and U1483 (N_1483,N_1344,N_1242);
or U1484 (N_1484,N_1218,N_1343);
and U1485 (N_1485,N_1239,N_1387);
nand U1486 (N_1486,N_1324,N_1367);
nand U1487 (N_1487,N_1279,N_1215);
xor U1488 (N_1488,N_1392,N_1354);
and U1489 (N_1489,N_1220,N_1352);
nand U1490 (N_1490,N_1372,N_1327);
and U1491 (N_1491,N_1349,N_1209);
and U1492 (N_1492,N_1267,N_1211);
xor U1493 (N_1493,N_1274,N_1320);
or U1494 (N_1494,N_1308,N_1273);
nand U1495 (N_1495,N_1332,N_1298);
and U1496 (N_1496,N_1225,N_1243);
nor U1497 (N_1497,N_1310,N_1236);
nand U1498 (N_1498,N_1348,N_1304);
nor U1499 (N_1499,N_1263,N_1271);
or U1500 (N_1500,N_1310,N_1203);
xnor U1501 (N_1501,N_1297,N_1336);
nand U1502 (N_1502,N_1316,N_1311);
nand U1503 (N_1503,N_1365,N_1391);
or U1504 (N_1504,N_1232,N_1207);
nor U1505 (N_1505,N_1225,N_1233);
or U1506 (N_1506,N_1288,N_1221);
nor U1507 (N_1507,N_1218,N_1217);
or U1508 (N_1508,N_1206,N_1235);
or U1509 (N_1509,N_1330,N_1261);
nand U1510 (N_1510,N_1245,N_1305);
nor U1511 (N_1511,N_1315,N_1354);
nand U1512 (N_1512,N_1344,N_1313);
or U1513 (N_1513,N_1323,N_1237);
nand U1514 (N_1514,N_1266,N_1307);
and U1515 (N_1515,N_1354,N_1321);
nand U1516 (N_1516,N_1253,N_1236);
nor U1517 (N_1517,N_1394,N_1281);
and U1518 (N_1518,N_1220,N_1328);
xnor U1519 (N_1519,N_1313,N_1307);
or U1520 (N_1520,N_1304,N_1202);
nor U1521 (N_1521,N_1307,N_1249);
and U1522 (N_1522,N_1292,N_1356);
nand U1523 (N_1523,N_1247,N_1302);
nand U1524 (N_1524,N_1289,N_1276);
or U1525 (N_1525,N_1217,N_1365);
nor U1526 (N_1526,N_1306,N_1282);
xor U1527 (N_1527,N_1322,N_1336);
or U1528 (N_1528,N_1232,N_1344);
nor U1529 (N_1529,N_1204,N_1349);
and U1530 (N_1530,N_1233,N_1392);
or U1531 (N_1531,N_1215,N_1330);
nand U1532 (N_1532,N_1323,N_1381);
xor U1533 (N_1533,N_1208,N_1248);
nor U1534 (N_1534,N_1217,N_1275);
xnor U1535 (N_1535,N_1207,N_1353);
or U1536 (N_1536,N_1353,N_1318);
nand U1537 (N_1537,N_1213,N_1341);
nor U1538 (N_1538,N_1328,N_1374);
and U1539 (N_1539,N_1238,N_1310);
and U1540 (N_1540,N_1379,N_1316);
xnor U1541 (N_1541,N_1268,N_1295);
or U1542 (N_1542,N_1333,N_1332);
nand U1543 (N_1543,N_1238,N_1303);
and U1544 (N_1544,N_1323,N_1336);
nor U1545 (N_1545,N_1283,N_1334);
nor U1546 (N_1546,N_1226,N_1358);
xnor U1547 (N_1547,N_1227,N_1311);
nor U1548 (N_1548,N_1261,N_1245);
nand U1549 (N_1549,N_1367,N_1343);
xnor U1550 (N_1550,N_1238,N_1234);
nand U1551 (N_1551,N_1246,N_1264);
and U1552 (N_1552,N_1314,N_1268);
nor U1553 (N_1553,N_1306,N_1331);
nand U1554 (N_1554,N_1328,N_1268);
and U1555 (N_1555,N_1293,N_1252);
xor U1556 (N_1556,N_1369,N_1333);
and U1557 (N_1557,N_1385,N_1301);
or U1558 (N_1558,N_1334,N_1281);
nand U1559 (N_1559,N_1275,N_1262);
nand U1560 (N_1560,N_1257,N_1282);
or U1561 (N_1561,N_1367,N_1326);
or U1562 (N_1562,N_1363,N_1324);
or U1563 (N_1563,N_1267,N_1310);
or U1564 (N_1564,N_1211,N_1325);
and U1565 (N_1565,N_1295,N_1229);
and U1566 (N_1566,N_1229,N_1252);
or U1567 (N_1567,N_1305,N_1391);
xor U1568 (N_1568,N_1252,N_1207);
nand U1569 (N_1569,N_1227,N_1319);
nor U1570 (N_1570,N_1397,N_1297);
and U1571 (N_1571,N_1335,N_1290);
and U1572 (N_1572,N_1384,N_1237);
nand U1573 (N_1573,N_1284,N_1203);
or U1574 (N_1574,N_1229,N_1277);
or U1575 (N_1575,N_1393,N_1351);
nor U1576 (N_1576,N_1227,N_1252);
or U1577 (N_1577,N_1223,N_1258);
nand U1578 (N_1578,N_1358,N_1294);
xor U1579 (N_1579,N_1201,N_1345);
nor U1580 (N_1580,N_1308,N_1399);
or U1581 (N_1581,N_1294,N_1228);
xnor U1582 (N_1582,N_1323,N_1253);
or U1583 (N_1583,N_1294,N_1335);
or U1584 (N_1584,N_1336,N_1330);
nand U1585 (N_1585,N_1241,N_1303);
nand U1586 (N_1586,N_1363,N_1329);
and U1587 (N_1587,N_1244,N_1373);
xor U1588 (N_1588,N_1356,N_1385);
nand U1589 (N_1589,N_1261,N_1295);
or U1590 (N_1590,N_1243,N_1258);
nor U1591 (N_1591,N_1264,N_1327);
or U1592 (N_1592,N_1262,N_1299);
and U1593 (N_1593,N_1337,N_1270);
nand U1594 (N_1594,N_1358,N_1295);
and U1595 (N_1595,N_1390,N_1280);
or U1596 (N_1596,N_1210,N_1354);
and U1597 (N_1597,N_1316,N_1229);
nand U1598 (N_1598,N_1243,N_1306);
or U1599 (N_1599,N_1369,N_1367);
and U1600 (N_1600,N_1507,N_1479);
or U1601 (N_1601,N_1508,N_1489);
or U1602 (N_1602,N_1592,N_1586);
nand U1603 (N_1603,N_1568,N_1525);
xnor U1604 (N_1604,N_1572,N_1443);
and U1605 (N_1605,N_1450,N_1478);
nand U1606 (N_1606,N_1584,N_1449);
nor U1607 (N_1607,N_1545,N_1515);
nand U1608 (N_1608,N_1430,N_1427);
or U1609 (N_1609,N_1419,N_1464);
nand U1610 (N_1610,N_1569,N_1583);
and U1611 (N_1611,N_1537,N_1485);
nand U1612 (N_1612,N_1514,N_1410);
or U1613 (N_1613,N_1442,N_1552);
nand U1614 (N_1614,N_1576,N_1589);
or U1615 (N_1615,N_1454,N_1403);
or U1616 (N_1616,N_1566,N_1599);
nand U1617 (N_1617,N_1404,N_1541);
nand U1618 (N_1618,N_1509,N_1482);
and U1619 (N_1619,N_1455,N_1435);
and U1620 (N_1620,N_1577,N_1581);
nand U1621 (N_1621,N_1495,N_1534);
nor U1622 (N_1622,N_1439,N_1516);
or U1623 (N_1623,N_1470,N_1555);
nor U1624 (N_1624,N_1557,N_1413);
nor U1625 (N_1625,N_1423,N_1594);
or U1626 (N_1626,N_1483,N_1571);
or U1627 (N_1627,N_1521,N_1529);
nand U1628 (N_1628,N_1472,N_1444);
nand U1629 (N_1629,N_1548,N_1400);
or U1630 (N_1630,N_1500,N_1432);
nor U1631 (N_1631,N_1501,N_1585);
and U1632 (N_1632,N_1575,N_1551);
and U1633 (N_1633,N_1418,N_1486);
or U1634 (N_1634,N_1567,N_1590);
nand U1635 (N_1635,N_1417,N_1463);
or U1636 (N_1636,N_1414,N_1491);
and U1637 (N_1637,N_1573,N_1456);
nor U1638 (N_1638,N_1416,N_1492);
or U1639 (N_1639,N_1591,N_1517);
nor U1640 (N_1640,N_1596,N_1593);
nand U1641 (N_1641,N_1532,N_1412);
or U1642 (N_1642,N_1510,N_1461);
xor U1643 (N_1643,N_1502,N_1422);
nand U1644 (N_1644,N_1563,N_1477);
and U1645 (N_1645,N_1465,N_1531);
and U1646 (N_1646,N_1578,N_1448);
and U1647 (N_1647,N_1429,N_1480);
and U1648 (N_1648,N_1499,N_1431);
or U1649 (N_1649,N_1528,N_1428);
nor U1650 (N_1650,N_1504,N_1474);
nand U1651 (N_1651,N_1595,N_1401);
nand U1652 (N_1652,N_1518,N_1560);
or U1653 (N_1653,N_1538,N_1459);
nor U1654 (N_1654,N_1408,N_1524);
nand U1655 (N_1655,N_1445,N_1526);
and U1656 (N_1656,N_1588,N_1497);
and U1657 (N_1657,N_1544,N_1542);
nand U1658 (N_1658,N_1471,N_1457);
or U1659 (N_1659,N_1536,N_1451);
nor U1660 (N_1660,N_1453,N_1582);
nor U1661 (N_1661,N_1433,N_1406);
nor U1662 (N_1662,N_1436,N_1550);
or U1663 (N_1663,N_1540,N_1460);
nand U1664 (N_1664,N_1475,N_1519);
nor U1665 (N_1665,N_1527,N_1434);
or U1666 (N_1666,N_1535,N_1498);
nor U1667 (N_1667,N_1447,N_1547);
or U1668 (N_1668,N_1466,N_1556);
nand U1669 (N_1669,N_1512,N_1462);
and U1670 (N_1670,N_1533,N_1481);
nand U1671 (N_1671,N_1562,N_1409);
or U1672 (N_1672,N_1437,N_1549);
xor U1673 (N_1673,N_1469,N_1496);
nand U1674 (N_1674,N_1598,N_1543);
nor U1675 (N_1675,N_1468,N_1503);
or U1676 (N_1676,N_1452,N_1476);
or U1677 (N_1677,N_1467,N_1438);
nand U1678 (N_1678,N_1415,N_1553);
and U1679 (N_1679,N_1446,N_1411);
nor U1680 (N_1680,N_1574,N_1546);
or U1681 (N_1681,N_1405,N_1579);
and U1682 (N_1682,N_1421,N_1511);
and U1683 (N_1683,N_1554,N_1522);
nor U1684 (N_1684,N_1458,N_1407);
nand U1685 (N_1685,N_1425,N_1490);
nand U1686 (N_1686,N_1565,N_1580);
and U1687 (N_1687,N_1424,N_1505);
nand U1688 (N_1688,N_1484,N_1506);
nor U1689 (N_1689,N_1523,N_1564);
nor U1690 (N_1690,N_1558,N_1487);
or U1691 (N_1691,N_1520,N_1493);
nor U1692 (N_1692,N_1402,N_1530);
nand U1693 (N_1693,N_1559,N_1513);
and U1694 (N_1694,N_1539,N_1597);
or U1695 (N_1695,N_1488,N_1570);
xor U1696 (N_1696,N_1420,N_1587);
nor U1697 (N_1697,N_1441,N_1561);
nand U1698 (N_1698,N_1440,N_1473);
or U1699 (N_1699,N_1494,N_1426);
or U1700 (N_1700,N_1524,N_1406);
nor U1701 (N_1701,N_1485,N_1541);
and U1702 (N_1702,N_1510,N_1569);
and U1703 (N_1703,N_1467,N_1500);
nand U1704 (N_1704,N_1473,N_1402);
nor U1705 (N_1705,N_1473,N_1501);
and U1706 (N_1706,N_1447,N_1576);
or U1707 (N_1707,N_1533,N_1462);
nor U1708 (N_1708,N_1422,N_1494);
or U1709 (N_1709,N_1547,N_1480);
or U1710 (N_1710,N_1508,N_1555);
and U1711 (N_1711,N_1469,N_1409);
nor U1712 (N_1712,N_1411,N_1477);
and U1713 (N_1713,N_1498,N_1425);
and U1714 (N_1714,N_1599,N_1590);
and U1715 (N_1715,N_1420,N_1593);
or U1716 (N_1716,N_1539,N_1501);
nand U1717 (N_1717,N_1452,N_1584);
nand U1718 (N_1718,N_1466,N_1469);
and U1719 (N_1719,N_1501,N_1548);
and U1720 (N_1720,N_1466,N_1486);
or U1721 (N_1721,N_1474,N_1517);
and U1722 (N_1722,N_1422,N_1460);
nand U1723 (N_1723,N_1553,N_1450);
or U1724 (N_1724,N_1414,N_1560);
and U1725 (N_1725,N_1535,N_1501);
and U1726 (N_1726,N_1579,N_1441);
nand U1727 (N_1727,N_1456,N_1417);
nor U1728 (N_1728,N_1429,N_1512);
xnor U1729 (N_1729,N_1464,N_1510);
or U1730 (N_1730,N_1423,N_1433);
and U1731 (N_1731,N_1497,N_1424);
nand U1732 (N_1732,N_1528,N_1550);
nand U1733 (N_1733,N_1405,N_1517);
and U1734 (N_1734,N_1552,N_1450);
nand U1735 (N_1735,N_1512,N_1591);
and U1736 (N_1736,N_1459,N_1574);
nor U1737 (N_1737,N_1507,N_1503);
xor U1738 (N_1738,N_1443,N_1541);
nand U1739 (N_1739,N_1599,N_1489);
and U1740 (N_1740,N_1535,N_1500);
xnor U1741 (N_1741,N_1550,N_1472);
nand U1742 (N_1742,N_1409,N_1533);
nor U1743 (N_1743,N_1570,N_1464);
and U1744 (N_1744,N_1419,N_1444);
and U1745 (N_1745,N_1597,N_1543);
nor U1746 (N_1746,N_1539,N_1596);
nor U1747 (N_1747,N_1507,N_1535);
and U1748 (N_1748,N_1573,N_1594);
nand U1749 (N_1749,N_1439,N_1402);
or U1750 (N_1750,N_1589,N_1475);
xor U1751 (N_1751,N_1560,N_1578);
or U1752 (N_1752,N_1523,N_1432);
or U1753 (N_1753,N_1537,N_1434);
or U1754 (N_1754,N_1410,N_1569);
xnor U1755 (N_1755,N_1543,N_1473);
and U1756 (N_1756,N_1449,N_1554);
or U1757 (N_1757,N_1538,N_1468);
nand U1758 (N_1758,N_1492,N_1581);
and U1759 (N_1759,N_1551,N_1449);
and U1760 (N_1760,N_1556,N_1496);
and U1761 (N_1761,N_1584,N_1480);
nand U1762 (N_1762,N_1462,N_1587);
xnor U1763 (N_1763,N_1560,N_1479);
xnor U1764 (N_1764,N_1461,N_1567);
or U1765 (N_1765,N_1587,N_1431);
nor U1766 (N_1766,N_1545,N_1409);
nor U1767 (N_1767,N_1534,N_1411);
and U1768 (N_1768,N_1491,N_1559);
and U1769 (N_1769,N_1493,N_1497);
nand U1770 (N_1770,N_1450,N_1501);
or U1771 (N_1771,N_1432,N_1572);
nor U1772 (N_1772,N_1511,N_1573);
nor U1773 (N_1773,N_1462,N_1500);
nor U1774 (N_1774,N_1467,N_1510);
and U1775 (N_1775,N_1490,N_1511);
nor U1776 (N_1776,N_1421,N_1547);
nor U1777 (N_1777,N_1420,N_1564);
or U1778 (N_1778,N_1577,N_1408);
nand U1779 (N_1779,N_1579,N_1570);
nor U1780 (N_1780,N_1449,N_1499);
xnor U1781 (N_1781,N_1403,N_1428);
or U1782 (N_1782,N_1577,N_1536);
nor U1783 (N_1783,N_1558,N_1421);
and U1784 (N_1784,N_1536,N_1457);
nor U1785 (N_1785,N_1535,N_1533);
and U1786 (N_1786,N_1570,N_1405);
or U1787 (N_1787,N_1486,N_1461);
or U1788 (N_1788,N_1423,N_1415);
and U1789 (N_1789,N_1581,N_1469);
nand U1790 (N_1790,N_1449,N_1460);
or U1791 (N_1791,N_1497,N_1518);
and U1792 (N_1792,N_1465,N_1427);
nand U1793 (N_1793,N_1415,N_1505);
nor U1794 (N_1794,N_1462,N_1598);
nand U1795 (N_1795,N_1487,N_1474);
nand U1796 (N_1796,N_1541,N_1458);
or U1797 (N_1797,N_1542,N_1553);
xnor U1798 (N_1798,N_1456,N_1497);
or U1799 (N_1799,N_1591,N_1513);
nand U1800 (N_1800,N_1674,N_1604);
nand U1801 (N_1801,N_1698,N_1760);
or U1802 (N_1802,N_1665,N_1720);
or U1803 (N_1803,N_1789,N_1769);
and U1804 (N_1804,N_1645,N_1702);
nand U1805 (N_1805,N_1711,N_1700);
or U1806 (N_1806,N_1642,N_1668);
nand U1807 (N_1807,N_1613,N_1740);
and U1808 (N_1808,N_1751,N_1755);
and U1809 (N_1809,N_1761,N_1683);
and U1810 (N_1810,N_1773,N_1716);
and U1811 (N_1811,N_1731,N_1710);
nor U1812 (N_1812,N_1794,N_1707);
and U1813 (N_1813,N_1697,N_1629);
nand U1814 (N_1814,N_1609,N_1682);
or U1815 (N_1815,N_1603,N_1633);
nor U1816 (N_1816,N_1623,N_1708);
nor U1817 (N_1817,N_1651,N_1791);
or U1818 (N_1818,N_1757,N_1727);
xor U1819 (N_1819,N_1639,N_1601);
and U1820 (N_1820,N_1656,N_1775);
nor U1821 (N_1821,N_1673,N_1774);
xor U1822 (N_1822,N_1787,N_1772);
or U1823 (N_1823,N_1684,N_1738);
or U1824 (N_1824,N_1641,N_1671);
nor U1825 (N_1825,N_1615,N_1765);
or U1826 (N_1826,N_1652,N_1699);
xor U1827 (N_1827,N_1703,N_1725);
and U1828 (N_1828,N_1767,N_1600);
or U1829 (N_1829,N_1732,N_1696);
nor U1830 (N_1830,N_1795,N_1786);
nor U1831 (N_1831,N_1621,N_1632);
or U1832 (N_1832,N_1602,N_1617);
nand U1833 (N_1833,N_1637,N_1655);
nor U1834 (N_1834,N_1677,N_1614);
or U1835 (N_1835,N_1743,N_1759);
nor U1836 (N_1836,N_1692,N_1663);
nor U1837 (N_1837,N_1709,N_1729);
and U1838 (N_1838,N_1622,N_1780);
and U1839 (N_1839,N_1689,N_1610);
or U1840 (N_1840,N_1741,N_1690);
and U1841 (N_1841,N_1763,N_1612);
nand U1842 (N_1842,N_1638,N_1721);
nand U1843 (N_1843,N_1744,N_1753);
xor U1844 (N_1844,N_1664,N_1784);
nand U1845 (N_1845,N_1693,N_1640);
and U1846 (N_1846,N_1799,N_1620);
nor U1847 (N_1847,N_1719,N_1606);
and U1848 (N_1848,N_1653,N_1736);
and U1849 (N_1849,N_1788,N_1717);
nand U1850 (N_1850,N_1666,N_1748);
and U1851 (N_1851,N_1752,N_1734);
nand U1852 (N_1852,N_1718,N_1662);
nor U1853 (N_1853,N_1605,N_1676);
nand U1854 (N_1854,N_1790,N_1627);
nor U1855 (N_1855,N_1750,N_1686);
and U1856 (N_1856,N_1783,N_1675);
nor U1857 (N_1857,N_1715,N_1607);
and U1858 (N_1858,N_1661,N_1793);
nand U1859 (N_1859,N_1694,N_1723);
nor U1860 (N_1860,N_1730,N_1636);
and U1861 (N_1861,N_1728,N_1658);
xnor U1862 (N_1862,N_1619,N_1798);
nand U1863 (N_1863,N_1669,N_1785);
or U1864 (N_1864,N_1737,N_1667);
or U1865 (N_1865,N_1688,N_1680);
nand U1866 (N_1866,N_1792,N_1722);
nor U1867 (N_1867,N_1781,N_1649);
xor U1868 (N_1868,N_1678,N_1749);
xnor U1869 (N_1869,N_1764,N_1779);
nand U1870 (N_1870,N_1766,N_1796);
or U1871 (N_1871,N_1681,N_1644);
or U1872 (N_1872,N_1778,N_1625);
nor U1873 (N_1873,N_1768,N_1782);
nor U1874 (N_1874,N_1776,N_1758);
nand U1875 (N_1875,N_1771,N_1714);
xor U1876 (N_1876,N_1691,N_1630);
nor U1877 (N_1877,N_1626,N_1631);
nor U1878 (N_1878,N_1654,N_1611);
nand U1879 (N_1879,N_1670,N_1745);
and U1880 (N_1880,N_1754,N_1643);
and U1881 (N_1881,N_1635,N_1695);
or U1882 (N_1882,N_1797,N_1616);
or U1883 (N_1883,N_1705,N_1726);
nand U1884 (N_1884,N_1624,N_1735);
nor U1885 (N_1885,N_1706,N_1742);
xnor U1886 (N_1886,N_1660,N_1608);
or U1887 (N_1887,N_1756,N_1646);
nor U1888 (N_1888,N_1704,N_1618);
and U1889 (N_1889,N_1770,N_1672);
xor U1890 (N_1890,N_1747,N_1657);
nor U1891 (N_1891,N_1650,N_1628);
nor U1892 (N_1892,N_1762,N_1724);
and U1893 (N_1893,N_1739,N_1746);
nand U1894 (N_1894,N_1712,N_1634);
or U1895 (N_1895,N_1659,N_1777);
nand U1896 (N_1896,N_1679,N_1648);
xnor U1897 (N_1897,N_1647,N_1687);
and U1898 (N_1898,N_1733,N_1685);
nor U1899 (N_1899,N_1701,N_1713);
xnor U1900 (N_1900,N_1743,N_1742);
or U1901 (N_1901,N_1639,N_1675);
nand U1902 (N_1902,N_1752,N_1621);
nand U1903 (N_1903,N_1649,N_1690);
and U1904 (N_1904,N_1686,N_1652);
nor U1905 (N_1905,N_1725,N_1652);
or U1906 (N_1906,N_1751,N_1690);
nor U1907 (N_1907,N_1698,N_1736);
or U1908 (N_1908,N_1691,N_1760);
or U1909 (N_1909,N_1689,N_1714);
and U1910 (N_1910,N_1777,N_1740);
and U1911 (N_1911,N_1721,N_1780);
and U1912 (N_1912,N_1676,N_1783);
and U1913 (N_1913,N_1664,N_1659);
nand U1914 (N_1914,N_1705,N_1778);
or U1915 (N_1915,N_1690,N_1707);
and U1916 (N_1916,N_1665,N_1706);
and U1917 (N_1917,N_1662,N_1666);
xor U1918 (N_1918,N_1722,N_1602);
nand U1919 (N_1919,N_1799,N_1776);
and U1920 (N_1920,N_1759,N_1670);
and U1921 (N_1921,N_1704,N_1791);
nand U1922 (N_1922,N_1795,N_1749);
nor U1923 (N_1923,N_1611,N_1645);
and U1924 (N_1924,N_1695,N_1676);
nor U1925 (N_1925,N_1621,N_1733);
or U1926 (N_1926,N_1680,N_1756);
nand U1927 (N_1927,N_1734,N_1697);
xor U1928 (N_1928,N_1750,N_1781);
nand U1929 (N_1929,N_1766,N_1630);
nor U1930 (N_1930,N_1682,N_1715);
nand U1931 (N_1931,N_1703,N_1623);
or U1932 (N_1932,N_1650,N_1664);
nand U1933 (N_1933,N_1689,N_1626);
and U1934 (N_1934,N_1794,N_1765);
nor U1935 (N_1935,N_1623,N_1723);
or U1936 (N_1936,N_1652,N_1759);
nor U1937 (N_1937,N_1741,N_1637);
nand U1938 (N_1938,N_1794,N_1611);
nor U1939 (N_1939,N_1763,N_1741);
nor U1940 (N_1940,N_1676,N_1608);
nor U1941 (N_1941,N_1717,N_1641);
or U1942 (N_1942,N_1672,N_1709);
nand U1943 (N_1943,N_1636,N_1691);
xnor U1944 (N_1944,N_1708,N_1781);
or U1945 (N_1945,N_1648,N_1744);
nand U1946 (N_1946,N_1600,N_1765);
and U1947 (N_1947,N_1617,N_1627);
nand U1948 (N_1948,N_1644,N_1634);
and U1949 (N_1949,N_1792,N_1736);
xnor U1950 (N_1950,N_1650,N_1775);
nand U1951 (N_1951,N_1684,N_1628);
nor U1952 (N_1952,N_1681,N_1753);
and U1953 (N_1953,N_1725,N_1645);
nor U1954 (N_1954,N_1612,N_1681);
nand U1955 (N_1955,N_1699,N_1638);
nor U1956 (N_1956,N_1715,N_1665);
nand U1957 (N_1957,N_1647,N_1790);
nand U1958 (N_1958,N_1750,N_1641);
nor U1959 (N_1959,N_1606,N_1782);
and U1960 (N_1960,N_1725,N_1650);
nand U1961 (N_1961,N_1700,N_1606);
and U1962 (N_1962,N_1744,N_1741);
nand U1963 (N_1963,N_1723,N_1731);
nand U1964 (N_1964,N_1794,N_1640);
xor U1965 (N_1965,N_1708,N_1772);
nor U1966 (N_1966,N_1704,N_1746);
nand U1967 (N_1967,N_1723,N_1650);
nand U1968 (N_1968,N_1708,N_1642);
or U1969 (N_1969,N_1757,N_1674);
and U1970 (N_1970,N_1746,N_1611);
and U1971 (N_1971,N_1795,N_1626);
and U1972 (N_1972,N_1731,N_1788);
or U1973 (N_1973,N_1722,N_1668);
nor U1974 (N_1974,N_1738,N_1765);
nor U1975 (N_1975,N_1765,N_1653);
and U1976 (N_1976,N_1742,N_1702);
nand U1977 (N_1977,N_1661,N_1621);
and U1978 (N_1978,N_1744,N_1762);
nand U1979 (N_1979,N_1679,N_1660);
nor U1980 (N_1980,N_1748,N_1774);
nand U1981 (N_1981,N_1793,N_1709);
or U1982 (N_1982,N_1734,N_1725);
or U1983 (N_1983,N_1751,N_1795);
and U1984 (N_1984,N_1789,N_1652);
nor U1985 (N_1985,N_1705,N_1789);
or U1986 (N_1986,N_1786,N_1623);
nor U1987 (N_1987,N_1743,N_1653);
nor U1988 (N_1988,N_1774,N_1724);
or U1989 (N_1989,N_1707,N_1703);
nor U1990 (N_1990,N_1621,N_1738);
and U1991 (N_1991,N_1654,N_1725);
nand U1992 (N_1992,N_1786,N_1642);
nor U1993 (N_1993,N_1775,N_1704);
nand U1994 (N_1994,N_1678,N_1723);
or U1995 (N_1995,N_1783,N_1712);
or U1996 (N_1996,N_1633,N_1714);
nand U1997 (N_1997,N_1790,N_1621);
nand U1998 (N_1998,N_1686,N_1732);
nand U1999 (N_1999,N_1742,N_1650);
nand U2000 (N_2000,N_1819,N_1844);
nand U2001 (N_2001,N_1925,N_1923);
and U2002 (N_2002,N_1857,N_1895);
nor U2003 (N_2003,N_1948,N_1805);
or U2004 (N_2004,N_1973,N_1914);
nand U2005 (N_2005,N_1909,N_1821);
xnor U2006 (N_2006,N_1818,N_1963);
xor U2007 (N_2007,N_1955,N_1950);
nand U2008 (N_2008,N_1831,N_1996);
xor U2009 (N_2009,N_1904,N_1985);
nor U2010 (N_2010,N_1897,N_1867);
nor U2011 (N_2011,N_1824,N_1829);
or U2012 (N_2012,N_1958,N_1969);
nand U2013 (N_2013,N_1920,N_1881);
or U2014 (N_2014,N_1850,N_1999);
xor U2015 (N_2015,N_1970,N_1924);
or U2016 (N_2016,N_1836,N_1875);
or U2017 (N_2017,N_1892,N_1838);
or U2018 (N_2018,N_1942,N_1975);
and U2019 (N_2019,N_1802,N_1801);
xnor U2020 (N_2020,N_1935,N_1862);
or U2021 (N_2021,N_1817,N_1915);
or U2022 (N_2022,N_1858,N_1957);
nor U2023 (N_2023,N_1986,N_1926);
nor U2024 (N_2024,N_1808,N_1843);
xnor U2025 (N_2025,N_1908,N_1855);
nor U2026 (N_2026,N_1882,N_1894);
nand U2027 (N_2027,N_1968,N_1974);
xor U2028 (N_2028,N_1834,N_1859);
and U2029 (N_2029,N_1931,N_1994);
nand U2030 (N_2030,N_1956,N_1848);
xor U2031 (N_2031,N_1959,N_1933);
and U2032 (N_2032,N_1903,N_1871);
nand U2033 (N_2033,N_1938,N_1823);
nor U2034 (N_2034,N_1912,N_1928);
nand U2035 (N_2035,N_1816,N_1980);
nor U2036 (N_2036,N_1868,N_1947);
xnor U2037 (N_2037,N_1847,N_1840);
nor U2038 (N_2038,N_1946,N_1837);
nor U2039 (N_2039,N_1813,N_1981);
nand U2040 (N_2040,N_1993,N_1934);
nor U2041 (N_2041,N_1917,N_1971);
and U2042 (N_2042,N_1893,N_1865);
nor U2043 (N_2043,N_1902,N_1954);
nand U2044 (N_2044,N_1916,N_1879);
or U2045 (N_2045,N_1812,N_1940);
xor U2046 (N_2046,N_1937,N_1827);
nor U2047 (N_2047,N_1851,N_1870);
and U2048 (N_2048,N_1866,N_1886);
nand U2049 (N_2049,N_1890,N_1896);
and U2050 (N_2050,N_1936,N_1811);
nand U2051 (N_2051,N_1911,N_1815);
nand U2052 (N_2052,N_1899,N_1861);
and U2053 (N_2053,N_1863,N_1845);
nor U2054 (N_2054,N_1921,N_1891);
or U2055 (N_2055,N_1989,N_1976);
nand U2056 (N_2056,N_1898,N_1939);
nand U2057 (N_2057,N_1951,N_1807);
and U2058 (N_2058,N_1992,N_1820);
nand U2059 (N_2059,N_1888,N_1952);
and U2060 (N_2060,N_1932,N_1982);
nand U2061 (N_2061,N_1849,N_1835);
nand U2062 (N_2062,N_1967,N_1919);
nor U2063 (N_2063,N_1822,N_1842);
xor U2064 (N_2064,N_1885,N_1826);
nor U2065 (N_2065,N_1809,N_1941);
nand U2066 (N_2066,N_1803,N_1901);
or U2067 (N_2067,N_1828,N_1841);
and U2068 (N_2068,N_1856,N_1918);
and U2069 (N_2069,N_1990,N_1987);
nor U2070 (N_2070,N_1943,N_1874);
nor U2071 (N_2071,N_1966,N_1961);
or U2072 (N_2072,N_1991,N_1988);
or U2073 (N_2073,N_1846,N_1979);
xor U2074 (N_2074,N_1825,N_1944);
nand U2075 (N_2075,N_1929,N_1839);
nand U2076 (N_2076,N_1983,N_1905);
and U2077 (N_2077,N_1814,N_1949);
xor U2078 (N_2078,N_1884,N_1800);
or U2079 (N_2079,N_1804,N_1876);
xnor U2080 (N_2080,N_1972,N_1878);
nor U2081 (N_2081,N_1880,N_1900);
or U2082 (N_2082,N_1910,N_1984);
or U2083 (N_2083,N_1860,N_1830);
nand U2084 (N_2084,N_1964,N_1806);
or U2085 (N_2085,N_1887,N_1853);
nand U2086 (N_2086,N_1883,N_1965);
and U2087 (N_2087,N_1945,N_1997);
xnor U2088 (N_2088,N_1833,N_1922);
or U2089 (N_2089,N_1889,N_1873);
nor U2090 (N_2090,N_1877,N_1913);
nor U2091 (N_2091,N_1995,N_1978);
xor U2092 (N_2092,N_1953,N_1864);
nor U2093 (N_2093,N_1960,N_1962);
or U2094 (N_2094,N_1854,N_1906);
or U2095 (N_2095,N_1998,N_1872);
nor U2096 (N_2096,N_1832,N_1930);
nor U2097 (N_2097,N_1907,N_1852);
and U2098 (N_2098,N_1810,N_1869);
and U2099 (N_2099,N_1977,N_1927);
nor U2100 (N_2100,N_1983,N_1981);
nor U2101 (N_2101,N_1973,N_1879);
or U2102 (N_2102,N_1889,N_1874);
or U2103 (N_2103,N_1811,N_1827);
and U2104 (N_2104,N_1863,N_1997);
and U2105 (N_2105,N_1824,N_1807);
nor U2106 (N_2106,N_1841,N_1981);
and U2107 (N_2107,N_1929,N_1962);
and U2108 (N_2108,N_1944,N_1914);
or U2109 (N_2109,N_1871,N_1938);
and U2110 (N_2110,N_1926,N_1841);
xnor U2111 (N_2111,N_1836,N_1867);
or U2112 (N_2112,N_1972,N_1906);
nand U2113 (N_2113,N_1907,N_1859);
or U2114 (N_2114,N_1937,N_1809);
nand U2115 (N_2115,N_1835,N_1820);
nor U2116 (N_2116,N_1947,N_1909);
nor U2117 (N_2117,N_1998,N_1941);
nand U2118 (N_2118,N_1964,N_1847);
or U2119 (N_2119,N_1938,N_1822);
nand U2120 (N_2120,N_1993,N_1896);
or U2121 (N_2121,N_1897,N_1999);
nand U2122 (N_2122,N_1819,N_1988);
or U2123 (N_2123,N_1843,N_1894);
or U2124 (N_2124,N_1917,N_1821);
or U2125 (N_2125,N_1905,N_1927);
nor U2126 (N_2126,N_1817,N_1976);
nor U2127 (N_2127,N_1871,N_1803);
nor U2128 (N_2128,N_1982,N_1922);
or U2129 (N_2129,N_1989,N_1943);
xnor U2130 (N_2130,N_1839,N_1834);
nor U2131 (N_2131,N_1924,N_1903);
nand U2132 (N_2132,N_1991,N_1811);
and U2133 (N_2133,N_1922,N_1841);
and U2134 (N_2134,N_1815,N_1984);
nand U2135 (N_2135,N_1870,N_1972);
or U2136 (N_2136,N_1993,N_1956);
or U2137 (N_2137,N_1817,N_1899);
or U2138 (N_2138,N_1968,N_1914);
and U2139 (N_2139,N_1876,N_1985);
xor U2140 (N_2140,N_1810,N_1849);
nand U2141 (N_2141,N_1975,N_1897);
nand U2142 (N_2142,N_1916,N_1957);
and U2143 (N_2143,N_1941,N_1992);
xor U2144 (N_2144,N_1883,N_1813);
and U2145 (N_2145,N_1988,N_1950);
nor U2146 (N_2146,N_1921,N_1843);
or U2147 (N_2147,N_1954,N_1907);
nand U2148 (N_2148,N_1881,N_1963);
nor U2149 (N_2149,N_1966,N_1818);
or U2150 (N_2150,N_1876,N_1806);
nor U2151 (N_2151,N_1926,N_1889);
nand U2152 (N_2152,N_1831,N_1976);
nand U2153 (N_2153,N_1878,N_1896);
nor U2154 (N_2154,N_1907,N_1958);
nand U2155 (N_2155,N_1912,N_1895);
or U2156 (N_2156,N_1877,N_1985);
or U2157 (N_2157,N_1898,N_1875);
nor U2158 (N_2158,N_1982,N_1949);
and U2159 (N_2159,N_1955,N_1975);
nor U2160 (N_2160,N_1862,N_1957);
and U2161 (N_2161,N_1843,N_1823);
and U2162 (N_2162,N_1978,N_1903);
nor U2163 (N_2163,N_1947,N_1991);
and U2164 (N_2164,N_1939,N_1855);
nor U2165 (N_2165,N_1873,N_1876);
nand U2166 (N_2166,N_1839,N_1816);
nor U2167 (N_2167,N_1968,N_1947);
xor U2168 (N_2168,N_1890,N_1946);
nor U2169 (N_2169,N_1937,N_1844);
and U2170 (N_2170,N_1937,N_1919);
and U2171 (N_2171,N_1824,N_1958);
or U2172 (N_2172,N_1900,N_1981);
nand U2173 (N_2173,N_1962,N_1976);
nor U2174 (N_2174,N_1812,N_1832);
or U2175 (N_2175,N_1952,N_1987);
and U2176 (N_2176,N_1949,N_1878);
nand U2177 (N_2177,N_1959,N_1882);
nand U2178 (N_2178,N_1878,N_1987);
and U2179 (N_2179,N_1832,N_1950);
nor U2180 (N_2180,N_1800,N_1855);
nor U2181 (N_2181,N_1875,N_1816);
xnor U2182 (N_2182,N_1957,N_1899);
nand U2183 (N_2183,N_1996,N_1900);
or U2184 (N_2184,N_1949,N_1919);
nand U2185 (N_2185,N_1965,N_1838);
and U2186 (N_2186,N_1944,N_1833);
nand U2187 (N_2187,N_1975,N_1927);
xor U2188 (N_2188,N_1994,N_1821);
and U2189 (N_2189,N_1881,N_1962);
nor U2190 (N_2190,N_1886,N_1991);
nor U2191 (N_2191,N_1830,N_1884);
or U2192 (N_2192,N_1898,N_1921);
nand U2193 (N_2193,N_1976,N_1921);
nand U2194 (N_2194,N_1934,N_1925);
or U2195 (N_2195,N_1867,N_1898);
nand U2196 (N_2196,N_1959,N_1938);
nor U2197 (N_2197,N_1994,N_1924);
xor U2198 (N_2198,N_1975,N_1920);
xnor U2199 (N_2199,N_1905,N_1959);
nor U2200 (N_2200,N_2027,N_2078);
or U2201 (N_2201,N_2017,N_2142);
or U2202 (N_2202,N_2186,N_2055);
nor U2203 (N_2203,N_2061,N_2146);
or U2204 (N_2204,N_2115,N_2183);
and U2205 (N_2205,N_2174,N_2148);
or U2206 (N_2206,N_2021,N_2164);
xor U2207 (N_2207,N_2188,N_2050);
nand U2208 (N_2208,N_2119,N_2054);
and U2209 (N_2209,N_2067,N_2172);
nand U2210 (N_2210,N_2006,N_2175);
xnor U2211 (N_2211,N_2039,N_2192);
or U2212 (N_2212,N_2150,N_2170);
nor U2213 (N_2213,N_2058,N_2092);
nand U2214 (N_2214,N_2152,N_2044);
nand U2215 (N_2215,N_2084,N_2029);
nor U2216 (N_2216,N_2035,N_2127);
nor U2217 (N_2217,N_2037,N_2162);
nor U2218 (N_2218,N_2168,N_2060);
or U2219 (N_2219,N_2022,N_2033);
and U2220 (N_2220,N_2081,N_2141);
nand U2221 (N_2221,N_2049,N_2112);
or U2222 (N_2222,N_2056,N_2167);
or U2223 (N_2223,N_2125,N_2197);
or U2224 (N_2224,N_2155,N_2179);
nand U2225 (N_2225,N_2087,N_2064);
or U2226 (N_2226,N_2026,N_2107);
nand U2227 (N_2227,N_2137,N_2117);
xnor U2228 (N_2228,N_2019,N_2130);
or U2229 (N_2229,N_2180,N_2088);
nor U2230 (N_2230,N_2030,N_2189);
nor U2231 (N_2231,N_2118,N_2114);
and U2232 (N_2232,N_2153,N_2063);
nor U2233 (N_2233,N_2124,N_2013);
xnor U2234 (N_2234,N_2139,N_2104);
or U2235 (N_2235,N_2121,N_2096);
nand U2236 (N_2236,N_2102,N_2090);
or U2237 (N_2237,N_2129,N_2069);
and U2238 (N_2238,N_2193,N_2163);
nand U2239 (N_2239,N_2178,N_2089);
nand U2240 (N_2240,N_2065,N_2110);
or U2241 (N_2241,N_2158,N_2147);
xnor U2242 (N_2242,N_2074,N_2181);
and U2243 (N_2243,N_2166,N_2126);
nand U2244 (N_2244,N_2062,N_2028);
nor U2245 (N_2245,N_2161,N_2135);
and U2246 (N_2246,N_2133,N_2196);
and U2247 (N_2247,N_2145,N_2076);
xor U2248 (N_2248,N_2190,N_2177);
or U2249 (N_2249,N_2036,N_2077);
nor U2250 (N_2250,N_2091,N_2016);
or U2251 (N_2251,N_2156,N_2000);
or U2252 (N_2252,N_2199,N_2014);
nand U2253 (N_2253,N_2048,N_2008);
nand U2254 (N_2254,N_2053,N_2111);
or U2255 (N_2255,N_2041,N_2025);
and U2256 (N_2256,N_2009,N_2079);
nor U2257 (N_2257,N_2151,N_2195);
nor U2258 (N_2258,N_2165,N_2080);
nor U2259 (N_2259,N_2085,N_2047);
nor U2260 (N_2260,N_2034,N_2106);
nor U2261 (N_2261,N_2004,N_2038);
nand U2262 (N_2262,N_2105,N_2007);
and U2263 (N_2263,N_2109,N_2154);
and U2264 (N_2264,N_2157,N_2131);
or U2265 (N_2265,N_2171,N_2012);
nand U2266 (N_2266,N_2045,N_2023);
xor U2267 (N_2267,N_2108,N_2099);
and U2268 (N_2268,N_2001,N_2100);
nand U2269 (N_2269,N_2120,N_2169);
or U2270 (N_2270,N_2182,N_2042);
nand U2271 (N_2271,N_2020,N_2176);
xor U2272 (N_2272,N_2015,N_2138);
nand U2273 (N_2273,N_2086,N_2082);
nor U2274 (N_2274,N_2103,N_2185);
xnor U2275 (N_2275,N_2046,N_2194);
and U2276 (N_2276,N_2043,N_2093);
xnor U2277 (N_2277,N_2032,N_2116);
xor U2278 (N_2278,N_2123,N_2052);
and U2279 (N_2279,N_2134,N_2132);
or U2280 (N_2280,N_2005,N_2002);
and U2281 (N_2281,N_2160,N_2136);
or U2282 (N_2282,N_2149,N_2191);
and U2283 (N_2283,N_2057,N_2075);
or U2284 (N_2284,N_2072,N_2128);
or U2285 (N_2285,N_2051,N_2059);
nand U2286 (N_2286,N_2066,N_2010);
or U2287 (N_2287,N_2097,N_2098);
and U2288 (N_2288,N_2122,N_2094);
xnor U2289 (N_2289,N_2073,N_2173);
and U2290 (N_2290,N_2071,N_2040);
and U2291 (N_2291,N_2031,N_2068);
nor U2292 (N_2292,N_2159,N_2140);
or U2293 (N_2293,N_2184,N_2024);
or U2294 (N_2294,N_2198,N_2070);
or U2295 (N_2295,N_2143,N_2018);
or U2296 (N_2296,N_2101,N_2011);
or U2297 (N_2297,N_2095,N_2003);
or U2298 (N_2298,N_2187,N_2083);
nor U2299 (N_2299,N_2113,N_2144);
or U2300 (N_2300,N_2027,N_2195);
or U2301 (N_2301,N_2167,N_2108);
or U2302 (N_2302,N_2118,N_2186);
or U2303 (N_2303,N_2096,N_2002);
nand U2304 (N_2304,N_2003,N_2025);
nor U2305 (N_2305,N_2161,N_2027);
nor U2306 (N_2306,N_2029,N_2197);
nor U2307 (N_2307,N_2005,N_2029);
or U2308 (N_2308,N_2111,N_2114);
xnor U2309 (N_2309,N_2053,N_2156);
and U2310 (N_2310,N_2057,N_2144);
nor U2311 (N_2311,N_2029,N_2054);
nand U2312 (N_2312,N_2033,N_2008);
and U2313 (N_2313,N_2151,N_2060);
nor U2314 (N_2314,N_2112,N_2163);
nand U2315 (N_2315,N_2071,N_2172);
nor U2316 (N_2316,N_2095,N_2150);
or U2317 (N_2317,N_2161,N_2133);
nand U2318 (N_2318,N_2078,N_2163);
or U2319 (N_2319,N_2193,N_2152);
nand U2320 (N_2320,N_2194,N_2093);
nand U2321 (N_2321,N_2020,N_2034);
or U2322 (N_2322,N_2067,N_2154);
nand U2323 (N_2323,N_2143,N_2091);
nand U2324 (N_2324,N_2173,N_2143);
nor U2325 (N_2325,N_2004,N_2159);
or U2326 (N_2326,N_2078,N_2028);
nand U2327 (N_2327,N_2015,N_2004);
or U2328 (N_2328,N_2058,N_2160);
and U2329 (N_2329,N_2123,N_2145);
or U2330 (N_2330,N_2158,N_2082);
and U2331 (N_2331,N_2060,N_2147);
and U2332 (N_2332,N_2022,N_2081);
and U2333 (N_2333,N_2050,N_2045);
and U2334 (N_2334,N_2164,N_2064);
nand U2335 (N_2335,N_2026,N_2142);
or U2336 (N_2336,N_2073,N_2049);
nand U2337 (N_2337,N_2121,N_2186);
xnor U2338 (N_2338,N_2078,N_2095);
nor U2339 (N_2339,N_2084,N_2125);
nor U2340 (N_2340,N_2102,N_2152);
or U2341 (N_2341,N_2128,N_2154);
or U2342 (N_2342,N_2020,N_2194);
nand U2343 (N_2343,N_2117,N_2131);
or U2344 (N_2344,N_2028,N_2012);
nand U2345 (N_2345,N_2047,N_2162);
nor U2346 (N_2346,N_2001,N_2013);
and U2347 (N_2347,N_2042,N_2070);
and U2348 (N_2348,N_2189,N_2083);
nand U2349 (N_2349,N_2147,N_2028);
nand U2350 (N_2350,N_2053,N_2022);
xnor U2351 (N_2351,N_2022,N_2166);
nand U2352 (N_2352,N_2083,N_2004);
xor U2353 (N_2353,N_2046,N_2058);
nand U2354 (N_2354,N_2171,N_2069);
nor U2355 (N_2355,N_2091,N_2000);
and U2356 (N_2356,N_2175,N_2091);
nand U2357 (N_2357,N_2030,N_2043);
and U2358 (N_2358,N_2171,N_2021);
or U2359 (N_2359,N_2032,N_2077);
or U2360 (N_2360,N_2162,N_2004);
nand U2361 (N_2361,N_2192,N_2072);
and U2362 (N_2362,N_2110,N_2150);
nor U2363 (N_2363,N_2008,N_2075);
nand U2364 (N_2364,N_2019,N_2127);
nand U2365 (N_2365,N_2137,N_2114);
nand U2366 (N_2366,N_2035,N_2137);
nor U2367 (N_2367,N_2162,N_2056);
or U2368 (N_2368,N_2017,N_2040);
and U2369 (N_2369,N_2113,N_2017);
xor U2370 (N_2370,N_2121,N_2151);
xor U2371 (N_2371,N_2107,N_2110);
nand U2372 (N_2372,N_2001,N_2041);
nor U2373 (N_2373,N_2032,N_2110);
xnor U2374 (N_2374,N_2075,N_2064);
or U2375 (N_2375,N_2017,N_2084);
nand U2376 (N_2376,N_2054,N_2067);
nand U2377 (N_2377,N_2117,N_2051);
and U2378 (N_2378,N_2090,N_2053);
nand U2379 (N_2379,N_2112,N_2109);
nand U2380 (N_2380,N_2163,N_2114);
nand U2381 (N_2381,N_2121,N_2048);
and U2382 (N_2382,N_2161,N_2141);
or U2383 (N_2383,N_2044,N_2130);
xor U2384 (N_2384,N_2037,N_2108);
and U2385 (N_2385,N_2027,N_2168);
xnor U2386 (N_2386,N_2084,N_2015);
or U2387 (N_2387,N_2167,N_2124);
and U2388 (N_2388,N_2032,N_2001);
and U2389 (N_2389,N_2134,N_2010);
nor U2390 (N_2390,N_2020,N_2187);
and U2391 (N_2391,N_2032,N_2061);
nor U2392 (N_2392,N_2064,N_2137);
and U2393 (N_2393,N_2122,N_2113);
nor U2394 (N_2394,N_2190,N_2199);
and U2395 (N_2395,N_2045,N_2059);
nor U2396 (N_2396,N_2026,N_2030);
or U2397 (N_2397,N_2172,N_2036);
and U2398 (N_2398,N_2020,N_2179);
or U2399 (N_2399,N_2195,N_2144);
nand U2400 (N_2400,N_2205,N_2289);
and U2401 (N_2401,N_2206,N_2285);
or U2402 (N_2402,N_2287,N_2308);
nor U2403 (N_2403,N_2213,N_2257);
nor U2404 (N_2404,N_2275,N_2380);
nand U2405 (N_2405,N_2227,N_2358);
nor U2406 (N_2406,N_2220,N_2346);
nand U2407 (N_2407,N_2207,N_2210);
xnor U2408 (N_2408,N_2381,N_2383);
or U2409 (N_2409,N_2351,N_2232);
nand U2410 (N_2410,N_2284,N_2339);
nand U2411 (N_2411,N_2378,N_2222);
xnor U2412 (N_2412,N_2369,N_2244);
and U2413 (N_2413,N_2215,N_2349);
nor U2414 (N_2414,N_2263,N_2370);
nor U2415 (N_2415,N_2353,N_2367);
xnor U2416 (N_2416,N_2274,N_2325);
nand U2417 (N_2417,N_2262,N_2318);
xor U2418 (N_2418,N_2338,N_2267);
and U2419 (N_2419,N_2343,N_2323);
and U2420 (N_2420,N_2331,N_2359);
xor U2421 (N_2421,N_2390,N_2217);
and U2422 (N_2422,N_2297,N_2395);
nor U2423 (N_2423,N_2397,N_2283);
nand U2424 (N_2424,N_2268,N_2312);
or U2425 (N_2425,N_2240,N_2347);
xnor U2426 (N_2426,N_2354,N_2337);
nand U2427 (N_2427,N_2335,N_2201);
nand U2428 (N_2428,N_2379,N_2326);
and U2429 (N_2429,N_2277,N_2256);
xnor U2430 (N_2430,N_2305,N_2269);
nor U2431 (N_2431,N_2355,N_2365);
xor U2432 (N_2432,N_2307,N_2228);
nand U2433 (N_2433,N_2317,N_2350);
nor U2434 (N_2434,N_2388,N_2316);
or U2435 (N_2435,N_2229,N_2321);
xor U2436 (N_2436,N_2238,N_2341);
nand U2437 (N_2437,N_2310,N_2278);
xnor U2438 (N_2438,N_2234,N_2292);
nand U2439 (N_2439,N_2348,N_2299);
nor U2440 (N_2440,N_2286,N_2243);
or U2441 (N_2441,N_2270,N_2253);
nor U2442 (N_2442,N_2265,N_2280);
nor U2443 (N_2443,N_2264,N_2300);
nand U2444 (N_2444,N_2294,N_2252);
or U2445 (N_2445,N_2324,N_2340);
nand U2446 (N_2446,N_2203,N_2313);
or U2447 (N_2447,N_2342,N_2301);
nor U2448 (N_2448,N_2245,N_2216);
and U2449 (N_2449,N_2291,N_2247);
or U2450 (N_2450,N_2271,N_2363);
and U2451 (N_2451,N_2306,N_2226);
or U2452 (N_2452,N_2385,N_2362);
nand U2453 (N_2453,N_2272,N_2230);
nand U2454 (N_2454,N_2315,N_2394);
nor U2455 (N_2455,N_2237,N_2327);
nor U2456 (N_2456,N_2309,N_2273);
or U2457 (N_2457,N_2218,N_2372);
nand U2458 (N_2458,N_2258,N_2235);
nor U2459 (N_2459,N_2333,N_2223);
or U2460 (N_2460,N_2202,N_2319);
nor U2461 (N_2461,N_2345,N_2224);
nand U2462 (N_2462,N_2281,N_2376);
nor U2463 (N_2463,N_2344,N_2371);
and U2464 (N_2464,N_2374,N_2311);
and U2465 (N_2465,N_2254,N_2304);
and U2466 (N_2466,N_2332,N_2320);
or U2467 (N_2467,N_2361,N_2352);
nand U2468 (N_2468,N_2399,N_2219);
or U2469 (N_2469,N_2255,N_2330);
nor U2470 (N_2470,N_2221,N_2328);
and U2471 (N_2471,N_2360,N_2329);
nand U2472 (N_2472,N_2368,N_2209);
and U2473 (N_2473,N_2248,N_2356);
or U2474 (N_2474,N_2276,N_2242);
xnor U2475 (N_2475,N_2246,N_2251);
xnor U2476 (N_2476,N_2392,N_2233);
xor U2477 (N_2477,N_2398,N_2282);
and U2478 (N_2478,N_2382,N_2236);
nor U2479 (N_2479,N_2239,N_2375);
nor U2480 (N_2480,N_2259,N_2391);
and U2481 (N_2481,N_2231,N_2266);
nor U2482 (N_2482,N_2373,N_2357);
nor U2483 (N_2483,N_2334,N_2288);
and U2484 (N_2484,N_2212,N_2250);
or U2485 (N_2485,N_2208,N_2204);
nand U2486 (N_2486,N_2377,N_2241);
and U2487 (N_2487,N_2303,N_2384);
nor U2488 (N_2488,N_2260,N_2200);
nand U2489 (N_2489,N_2261,N_2389);
and U2490 (N_2490,N_2396,N_2214);
nand U2491 (N_2491,N_2364,N_2298);
nand U2492 (N_2492,N_2366,N_2225);
nor U2493 (N_2493,N_2322,N_2211);
and U2494 (N_2494,N_2295,N_2386);
and U2495 (N_2495,N_2314,N_2302);
nor U2496 (N_2496,N_2393,N_2336);
or U2497 (N_2497,N_2296,N_2290);
or U2498 (N_2498,N_2279,N_2293);
or U2499 (N_2499,N_2387,N_2249);
and U2500 (N_2500,N_2339,N_2281);
and U2501 (N_2501,N_2362,N_2212);
nor U2502 (N_2502,N_2389,N_2202);
and U2503 (N_2503,N_2256,N_2358);
nand U2504 (N_2504,N_2216,N_2394);
nor U2505 (N_2505,N_2308,N_2277);
or U2506 (N_2506,N_2365,N_2256);
nand U2507 (N_2507,N_2329,N_2271);
and U2508 (N_2508,N_2227,N_2278);
or U2509 (N_2509,N_2222,N_2224);
or U2510 (N_2510,N_2306,N_2271);
nand U2511 (N_2511,N_2384,N_2200);
nand U2512 (N_2512,N_2341,N_2355);
and U2513 (N_2513,N_2261,N_2262);
xor U2514 (N_2514,N_2215,N_2368);
xor U2515 (N_2515,N_2291,N_2301);
xnor U2516 (N_2516,N_2213,N_2351);
xor U2517 (N_2517,N_2389,N_2230);
nand U2518 (N_2518,N_2256,N_2254);
and U2519 (N_2519,N_2371,N_2343);
and U2520 (N_2520,N_2370,N_2282);
or U2521 (N_2521,N_2231,N_2312);
and U2522 (N_2522,N_2249,N_2277);
nand U2523 (N_2523,N_2288,N_2251);
xnor U2524 (N_2524,N_2271,N_2370);
nand U2525 (N_2525,N_2247,N_2250);
or U2526 (N_2526,N_2356,N_2274);
nor U2527 (N_2527,N_2334,N_2314);
or U2528 (N_2528,N_2330,N_2253);
nand U2529 (N_2529,N_2393,N_2233);
xnor U2530 (N_2530,N_2359,N_2204);
nor U2531 (N_2531,N_2367,N_2336);
nor U2532 (N_2532,N_2369,N_2379);
or U2533 (N_2533,N_2323,N_2367);
nand U2534 (N_2534,N_2248,N_2200);
or U2535 (N_2535,N_2266,N_2209);
and U2536 (N_2536,N_2354,N_2273);
or U2537 (N_2537,N_2335,N_2353);
nor U2538 (N_2538,N_2286,N_2321);
and U2539 (N_2539,N_2241,N_2254);
and U2540 (N_2540,N_2280,N_2368);
or U2541 (N_2541,N_2210,N_2246);
nor U2542 (N_2542,N_2316,N_2363);
nand U2543 (N_2543,N_2307,N_2264);
or U2544 (N_2544,N_2214,N_2227);
or U2545 (N_2545,N_2259,N_2218);
nor U2546 (N_2546,N_2229,N_2220);
nor U2547 (N_2547,N_2311,N_2289);
or U2548 (N_2548,N_2249,N_2220);
or U2549 (N_2549,N_2366,N_2313);
nor U2550 (N_2550,N_2331,N_2394);
or U2551 (N_2551,N_2255,N_2230);
nand U2552 (N_2552,N_2369,N_2319);
and U2553 (N_2553,N_2203,N_2332);
nand U2554 (N_2554,N_2239,N_2398);
nand U2555 (N_2555,N_2353,N_2380);
nand U2556 (N_2556,N_2257,N_2362);
nor U2557 (N_2557,N_2357,N_2243);
nor U2558 (N_2558,N_2268,N_2290);
nand U2559 (N_2559,N_2261,N_2312);
nand U2560 (N_2560,N_2279,N_2268);
nor U2561 (N_2561,N_2287,N_2257);
nand U2562 (N_2562,N_2214,N_2380);
nor U2563 (N_2563,N_2360,N_2357);
nand U2564 (N_2564,N_2210,N_2358);
nand U2565 (N_2565,N_2299,N_2259);
xor U2566 (N_2566,N_2360,N_2387);
or U2567 (N_2567,N_2339,N_2226);
nand U2568 (N_2568,N_2359,N_2257);
or U2569 (N_2569,N_2276,N_2392);
or U2570 (N_2570,N_2325,N_2284);
nor U2571 (N_2571,N_2289,N_2211);
and U2572 (N_2572,N_2339,N_2224);
xor U2573 (N_2573,N_2295,N_2306);
nor U2574 (N_2574,N_2230,N_2258);
nor U2575 (N_2575,N_2300,N_2392);
nor U2576 (N_2576,N_2388,N_2318);
xor U2577 (N_2577,N_2291,N_2234);
or U2578 (N_2578,N_2273,N_2282);
and U2579 (N_2579,N_2273,N_2307);
or U2580 (N_2580,N_2301,N_2238);
and U2581 (N_2581,N_2270,N_2366);
or U2582 (N_2582,N_2399,N_2215);
nand U2583 (N_2583,N_2345,N_2213);
nor U2584 (N_2584,N_2262,N_2306);
nor U2585 (N_2585,N_2385,N_2223);
xor U2586 (N_2586,N_2241,N_2213);
or U2587 (N_2587,N_2301,N_2399);
or U2588 (N_2588,N_2281,N_2354);
nor U2589 (N_2589,N_2342,N_2241);
nand U2590 (N_2590,N_2277,N_2255);
nand U2591 (N_2591,N_2321,N_2217);
or U2592 (N_2592,N_2257,N_2211);
nand U2593 (N_2593,N_2207,N_2211);
nand U2594 (N_2594,N_2243,N_2215);
nor U2595 (N_2595,N_2289,N_2273);
nand U2596 (N_2596,N_2344,N_2259);
nor U2597 (N_2597,N_2370,N_2227);
nand U2598 (N_2598,N_2360,N_2365);
nor U2599 (N_2599,N_2259,N_2255);
nand U2600 (N_2600,N_2523,N_2486);
nor U2601 (N_2601,N_2442,N_2489);
xor U2602 (N_2602,N_2585,N_2406);
nand U2603 (N_2603,N_2452,N_2465);
nand U2604 (N_2604,N_2451,N_2410);
or U2605 (N_2605,N_2584,N_2598);
or U2606 (N_2606,N_2447,N_2586);
nand U2607 (N_2607,N_2545,N_2468);
nand U2608 (N_2608,N_2548,N_2524);
nand U2609 (N_2609,N_2423,N_2459);
and U2610 (N_2610,N_2466,N_2544);
xnor U2611 (N_2611,N_2424,N_2530);
and U2612 (N_2612,N_2538,N_2507);
nand U2613 (N_2613,N_2470,N_2564);
xnor U2614 (N_2614,N_2418,N_2573);
or U2615 (N_2615,N_2593,N_2482);
or U2616 (N_2616,N_2481,N_2493);
and U2617 (N_2617,N_2582,N_2492);
nor U2618 (N_2618,N_2588,N_2551);
nand U2619 (N_2619,N_2566,N_2401);
or U2620 (N_2620,N_2460,N_2562);
and U2621 (N_2621,N_2549,N_2514);
nand U2622 (N_2622,N_2463,N_2577);
or U2623 (N_2623,N_2509,N_2536);
xnor U2624 (N_2624,N_2483,N_2532);
nand U2625 (N_2625,N_2431,N_2501);
and U2626 (N_2626,N_2429,N_2477);
nand U2627 (N_2627,N_2533,N_2517);
nand U2628 (N_2628,N_2529,N_2455);
nand U2629 (N_2629,N_2415,N_2405);
or U2630 (N_2630,N_2578,N_2449);
or U2631 (N_2631,N_2510,N_2525);
or U2632 (N_2632,N_2400,N_2464);
nand U2633 (N_2633,N_2432,N_2520);
and U2634 (N_2634,N_2554,N_2560);
nor U2635 (N_2635,N_2416,N_2467);
or U2636 (N_2636,N_2445,N_2474);
nand U2637 (N_2637,N_2535,N_2433);
nand U2638 (N_2638,N_2568,N_2462);
and U2639 (N_2639,N_2439,N_2557);
and U2640 (N_2640,N_2440,N_2526);
nand U2641 (N_2641,N_2475,N_2472);
nor U2642 (N_2642,N_2450,N_2441);
nand U2643 (N_2643,N_2414,N_2417);
xnor U2644 (N_2644,N_2518,N_2583);
or U2645 (N_2645,N_2569,N_2487);
or U2646 (N_2646,N_2402,N_2555);
nor U2647 (N_2647,N_2541,N_2500);
and U2648 (N_2648,N_2543,N_2425);
nand U2649 (N_2649,N_2456,N_2575);
or U2650 (N_2650,N_2419,N_2488);
nor U2651 (N_2651,N_2437,N_2559);
or U2652 (N_2652,N_2594,N_2521);
and U2653 (N_2653,N_2494,N_2595);
or U2654 (N_2654,N_2552,N_2576);
nand U2655 (N_2655,N_2561,N_2589);
nor U2656 (N_2656,N_2491,N_2502);
and U2657 (N_2657,N_2574,N_2531);
nand U2658 (N_2658,N_2430,N_2422);
or U2659 (N_2659,N_2565,N_2454);
and U2660 (N_2660,N_2498,N_2408);
xnor U2661 (N_2661,N_2527,N_2484);
or U2662 (N_2662,N_2404,N_2409);
and U2663 (N_2663,N_2499,N_2540);
or U2664 (N_2664,N_2426,N_2438);
and U2665 (N_2665,N_2444,N_2542);
or U2666 (N_2666,N_2485,N_2413);
nor U2667 (N_2667,N_2539,N_2537);
and U2668 (N_2668,N_2547,N_2443);
xnor U2669 (N_2669,N_2495,N_2587);
xnor U2670 (N_2670,N_2504,N_2556);
xor U2671 (N_2671,N_2469,N_2599);
nor U2672 (N_2672,N_2512,N_2479);
nand U2673 (N_2673,N_2420,N_2503);
nand U2674 (N_2674,N_2558,N_2403);
nand U2675 (N_2675,N_2446,N_2546);
and U2676 (N_2676,N_2436,N_2473);
nand U2677 (N_2677,N_2428,N_2579);
xor U2678 (N_2678,N_2434,N_2563);
or U2679 (N_2679,N_2496,N_2421);
nor U2680 (N_2680,N_2457,N_2407);
nor U2681 (N_2681,N_2596,N_2480);
and U2682 (N_2682,N_2592,N_2597);
nand U2683 (N_2683,N_2411,N_2412);
and U2684 (N_2684,N_2553,N_2448);
and U2685 (N_2685,N_2461,N_2435);
or U2686 (N_2686,N_2476,N_2458);
and U2687 (N_2687,N_2513,N_2511);
and U2688 (N_2688,N_2550,N_2471);
nor U2689 (N_2689,N_2591,N_2505);
nand U2690 (N_2690,N_2581,N_2478);
or U2691 (N_2691,N_2572,N_2427);
and U2692 (N_2692,N_2519,N_2590);
and U2693 (N_2693,N_2570,N_2516);
and U2694 (N_2694,N_2508,N_2580);
or U2695 (N_2695,N_2506,N_2453);
nor U2696 (N_2696,N_2522,N_2497);
or U2697 (N_2697,N_2567,N_2571);
xnor U2698 (N_2698,N_2528,N_2515);
and U2699 (N_2699,N_2534,N_2490);
nand U2700 (N_2700,N_2509,N_2520);
nand U2701 (N_2701,N_2445,N_2542);
or U2702 (N_2702,N_2510,N_2595);
and U2703 (N_2703,N_2556,N_2572);
xor U2704 (N_2704,N_2464,N_2559);
or U2705 (N_2705,N_2536,N_2511);
and U2706 (N_2706,N_2420,N_2465);
nor U2707 (N_2707,N_2476,N_2560);
nor U2708 (N_2708,N_2530,N_2460);
nor U2709 (N_2709,N_2438,N_2423);
nand U2710 (N_2710,N_2466,N_2454);
or U2711 (N_2711,N_2548,N_2429);
or U2712 (N_2712,N_2490,N_2565);
nor U2713 (N_2713,N_2446,N_2571);
or U2714 (N_2714,N_2443,N_2405);
and U2715 (N_2715,N_2504,N_2413);
and U2716 (N_2716,N_2507,N_2515);
or U2717 (N_2717,N_2522,N_2548);
and U2718 (N_2718,N_2451,N_2486);
nand U2719 (N_2719,N_2465,N_2538);
or U2720 (N_2720,N_2599,N_2420);
nor U2721 (N_2721,N_2430,N_2566);
nor U2722 (N_2722,N_2543,N_2504);
or U2723 (N_2723,N_2579,N_2430);
xor U2724 (N_2724,N_2428,N_2415);
or U2725 (N_2725,N_2426,N_2528);
xnor U2726 (N_2726,N_2432,N_2457);
nor U2727 (N_2727,N_2537,N_2511);
nor U2728 (N_2728,N_2563,N_2473);
or U2729 (N_2729,N_2474,N_2587);
or U2730 (N_2730,N_2573,N_2434);
nor U2731 (N_2731,N_2455,N_2536);
or U2732 (N_2732,N_2520,N_2478);
xnor U2733 (N_2733,N_2547,N_2553);
xnor U2734 (N_2734,N_2595,N_2402);
or U2735 (N_2735,N_2579,N_2596);
nor U2736 (N_2736,N_2443,N_2595);
and U2737 (N_2737,N_2509,N_2575);
nor U2738 (N_2738,N_2416,N_2457);
nor U2739 (N_2739,N_2553,N_2539);
or U2740 (N_2740,N_2567,N_2557);
nor U2741 (N_2741,N_2545,N_2586);
nor U2742 (N_2742,N_2540,N_2553);
nand U2743 (N_2743,N_2445,N_2468);
xnor U2744 (N_2744,N_2593,N_2430);
and U2745 (N_2745,N_2598,N_2518);
xnor U2746 (N_2746,N_2496,N_2422);
and U2747 (N_2747,N_2487,N_2594);
and U2748 (N_2748,N_2577,N_2530);
and U2749 (N_2749,N_2418,N_2403);
nand U2750 (N_2750,N_2450,N_2403);
or U2751 (N_2751,N_2518,N_2564);
xnor U2752 (N_2752,N_2583,N_2441);
nor U2753 (N_2753,N_2459,N_2442);
nand U2754 (N_2754,N_2431,N_2450);
or U2755 (N_2755,N_2489,N_2485);
xor U2756 (N_2756,N_2510,N_2581);
xnor U2757 (N_2757,N_2419,N_2460);
xor U2758 (N_2758,N_2428,N_2478);
xor U2759 (N_2759,N_2545,N_2481);
nand U2760 (N_2760,N_2407,N_2490);
nand U2761 (N_2761,N_2568,N_2429);
or U2762 (N_2762,N_2516,N_2568);
nor U2763 (N_2763,N_2578,N_2465);
or U2764 (N_2764,N_2418,N_2484);
nor U2765 (N_2765,N_2599,N_2508);
nor U2766 (N_2766,N_2483,N_2499);
nand U2767 (N_2767,N_2513,N_2522);
nand U2768 (N_2768,N_2468,N_2522);
or U2769 (N_2769,N_2515,N_2585);
or U2770 (N_2770,N_2580,N_2463);
and U2771 (N_2771,N_2427,N_2492);
nand U2772 (N_2772,N_2463,N_2456);
nor U2773 (N_2773,N_2478,N_2546);
and U2774 (N_2774,N_2439,N_2567);
nand U2775 (N_2775,N_2531,N_2590);
or U2776 (N_2776,N_2441,N_2400);
nand U2777 (N_2777,N_2530,N_2547);
nand U2778 (N_2778,N_2599,N_2552);
nor U2779 (N_2779,N_2512,N_2400);
nor U2780 (N_2780,N_2455,N_2463);
nand U2781 (N_2781,N_2474,N_2513);
or U2782 (N_2782,N_2416,N_2521);
or U2783 (N_2783,N_2500,N_2426);
nor U2784 (N_2784,N_2460,N_2504);
and U2785 (N_2785,N_2408,N_2462);
nor U2786 (N_2786,N_2466,N_2414);
or U2787 (N_2787,N_2535,N_2519);
and U2788 (N_2788,N_2551,N_2475);
nand U2789 (N_2789,N_2504,N_2526);
or U2790 (N_2790,N_2521,N_2485);
nand U2791 (N_2791,N_2541,N_2495);
or U2792 (N_2792,N_2537,N_2433);
or U2793 (N_2793,N_2513,N_2401);
or U2794 (N_2794,N_2442,N_2586);
and U2795 (N_2795,N_2589,N_2431);
and U2796 (N_2796,N_2449,N_2400);
nand U2797 (N_2797,N_2455,N_2406);
nand U2798 (N_2798,N_2478,N_2589);
nor U2799 (N_2799,N_2552,N_2407);
xnor U2800 (N_2800,N_2639,N_2746);
nor U2801 (N_2801,N_2645,N_2672);
nand U2802 (N_2802,N_2754,N_2619);
nor U2803 (N_2803,N_2647,N_2708);
nand U2804 (N_2804,N_2684,N_2679);
nand U2805 (N_2805,N_2756,N_2603);
or U2806 (N_2806,N_2730,N_2698);
nand U2807 (N_2807,N_2699,N_2649);
and U2808 (N_2808,N_2697,N_2627);
nand U2809 (N_2809,N_2765,N_2626);
xor U2810 (N_2810,N_2682,N_2776);
nand U2811 (N_2811,N_2790,N_2613);
and U2812 (N_2812,N_2767,N_2691);
or U2813 (N_2813,N_2702,N_2662);
or U2814 (N_2814,N_2611,N_2719);
nor U2815 (N_2815,N_2720,N_2782);
nor U2816 (N_2816,N_2640,N_2723);
nor U2817 (N_2817,N_2605,N_2636);
and U2818 (N_2818,N_2617,N_2637);
and U2819 (N_2819,N_2629,N_2631);
and U2820 (N_2820,N_2665,N_2681);
nor U2821 (N_2821,N_2709,N_2722);
nor U2822 (N_2822,N_2721,N_2784);
xnor U2823 (N_2823,N_2751,N_2728);
and U2824 (N_2824,N_2610,N_2628);
or U2825 (N_2825,N_2655,N_2602);
and U2826 (N_2826,N_2692,N_2703);
or U2827 (N_2827,N_2715,N_2607);
or U2828 (N_2828,N_2774,N_2620);
nand U2829 (N_2829,N_2623,N_2695);
or U2830 (N_2830,N_2742,N_2734);
nor U2831 (N_2831,N_2789,N_2771);
or U2832 (N_2832,N_2759,N_2676);
and U2833 (N_2833,N_2741,N_2726);
xnor U2834 (N_2834,N_2614,N_2712);
and U2835 (N_2835,N_2704,N_2764);
nor U2836 (N_2836,N_2729,N_2653);
nor U2837 (N_2837,N_2668,N_2615);
or U2838 (N_2838,N_2641,N_2609);
nor U2839 (N_2839,N_2600,N_2671);
nand U2840 (N_2840,N_2735,N_2747);
and U2841 (N_2841,N_2783,N_2638);
and U2842 (N_2842,N_2750,N_2731);
nor U2843 (N_2843,N_2624,N_2630);
xnor U2844 (N_2844,N_2644,N_2714);
nor U2845 (N_2845,N_2689,N_2744);
nor U2846 (N_2846,N_2710,N_2643);
nand U2847 (N_2847,N_2660,N_2652);
nand U2848 (N_2848,N_2727,N_2748);
nor U2849 (N_2849,N_2778,N_2670);
and U2850 (N_2850,N_2718,N_2745);
or U2851 (N_2851,N_2666,N_2766);
xor U2852 (N_2852,N_2758,N_2687);
and U2853 (N_2853,N_2632,N_2622);
and U2854 (N_2854,N_2799,N_2752);
xnor U2855 (N_2855,N_2673,N_2791);
and U2856 (N_2856,N_2664,N_2635);
nand U2857 (N_2857,N_2794,N_2616);
or U2858 (N_2858,N_2667,N_2795);
and U2859 (N_2859,N_2793,N_2701);
or U2860 (N_2860,N_2733,N_2693);
or U2861 (N_2861,N_2642,N_2680);
nor U2862 (N_2862,N_2705,N_2654);
nor U2863 (N_2863,N_2753,N_2677);
nand U2864 (N_2864,N_2707,N_2732);
or U2865 (N_2865,N_2740,N_2760);
or U2866 (N_2866,N_2775,N_2787);
nor U2867 (N_2867,N_2674,N_2792);
xor U2868 (N_2868,N_2651,N_2621);
and U2869 (N_2869,N_2669,N_2683);
or U2870 (N_2870,N_2763,N_2656);
and U2871 (N_2871,N_2601,N_2755);
and U2872 (N_2872,N_2772,N_2663);
nand U2873 (N_2873,N_2738,N_2657);
and U2874 (N_2874,N_2659,N_2625);
and U2875 (N_2875,N_2604,N_2780);
nor U2876 (N_2876,N_2777,N_2646);
and U2877 (N_2877,N_2608,N_2675);
nor U2878 (N_2878,N_2686,N_2713);
nand U2879 (N_2879,N_2779,N_2706);
xor U2880 (N_2880,N_2737,N_2762);
nor U2881 (N_2881,N_2606,N_2658);
nor U2882 (N_2882,N_2736,N_2757);
nand U2883 (N_2883,N_2612,N_2650);
xor U2884 (N_2884,N_2690,N_2717);
nand U2885 (N_2885,N_2724,N_2785);
nand U2886 (N_2886,N_2769,N_2786);
and U2887 (N_2887,N_2788,N_2739);
nor U2888 (N_2888,N_2781,N_2743);
and U2889 (N_2889,N_2685,N_2798);
nand U2890 (N_2890,N_2749,N_2725);
xnor U2891 (N_2891,N_2694,N_2678);
and U2892 (N_2892,N_2711,N_2796);
nand U2893 (N_2893,N_2661,N_2688);
or U2894 (N_2894,N_2770,N_2648);
nor U2895 (N_2895,N_2700,N_2696);
nor U2896 (N_2896,N_2633,N_2797);
or U2897 (N_2897,N_2634,N_2761);
or U2898 (N_2898,N_2768,N_2773);
nor U2899 (N_2899,N_2716,N_2618);
nand U2900 (N_2900,N_2648,N_2702);
and U2901 (N_2901,N_2719,N_2687);
or U2902 (N_2902,N_2705,N_2605);
or U2903 (N_2903,N_2685,N_2638);
xor U2904 (N_2904,N_2718,N_2601);
nand U2905 (N_2905,N_2658,N_2676);
nand U2906 (N_2906,N_2669,N_2704);
and U2907 (N_2907,N_2744,N_2732);
nand U2908 (N_2908,N_2626,N_2676);
nor U2909 (N_2909,N_2683,N_2661);
and U2910 (N_2910,N_2686,N_2780);
and U2911 (N_2911,N_2722,N_2629);
and U2912 (N_2912,N_2648,N_2707);
and U2913 (N_2913,N_2627,N_2717);
or U2914 (N_2914,N_2778,N_2739);
xnor U2915 (N_2915,N_2655,N_2787);
nand U2916 (N_2916,N_2696,N_2682);
or U2917 (N_2917,N_2679,N_2693);
or U2918 (N_2918,N_2750,N_2726);
or U2919 (N_2919,N_2679,N_2724);
nor U2920 (N_2920,N_2785,N_2757);
nor U2921 (N_2921,N_2754,N_2666);
nor U2922 (N_2922,N_2690,N_2685);
or U2923 (N_2923,N_2673,N_2699);
nand U2924 (N_2924,N_2621,N_2695);
xor U2925 (N_2925,N_2764,N_2760);
nor U2926 (N_2926,N_2715,N_2648);
or U2927 (N_2927,N_2743,N_2698);
nor U2928 (N_2928,N_2703,N_2779);
nor U2929 (N_2929,N_2783,N_2751);
and U2930 (N_2930,N_2605,N_2615);
xnor U2931 (N_2931,N_2674,N_2677);
nor U2932 (N_2932,N_2754,N_2746);
nor U2933 (N_2933,N_2798,N_2624);
nor U2934 (N_2934,N_2713,N_2641);
or U2935 (N_2935,N_2677,N_2602);
or U2936 (N_2936,N_2610,N_2722);
nand U2937 (N_2937,N_2708,N_2650);
nand U2938 (N_2938,N_2675,N_2694);
nand U2939 (N_2939,N_2624,N_2736);
and U2940 (N_2940,N_2752,N_2716);
nor U2941 (N_2941,N_2695,N_2636);
nor U2942 (N_2942,N_2616,N_2610);
and U2943 (N_2943,N_2642,N_2671);
nor U2944 (N_2944,N_2791,N_2782);
nand U2945 (N_2945,N_2738,N_2691);
or U2946 (N_2946,N_2691,N_2616);
nor U2947 (N_2947,N_2715,N_2661);
or U2948 (N_2948,N_2768,N_2619);
and U2949 (N_2949,N_2617,N_2773);
nor U2950 (N_2950,N_2707,N_2701);
nand U2951 (N_2951,N_2686,N_2712);
and U2952 (N_2952,N_2665,N_2660);
or U2953 (N_2953,N_2638,N_2751);
and U2954 (N_2954,N_2773,N_2642);
and U2955 (N_2955,N_2743,N_2751);
and U2956 (N_2956,N_2684,N_2613);
nor U2957 (N_2957,N_2795,N_2698);
or U2958 (N_2958,N_2674,N_2762);
and U2959 (N_2959,N_2653,N_2738);
nor U2960 (N_2960,N_2707,N_2620);
and U2961 (N_2961,N_2699,N_2768);
xor U2962 (N_2962,N_2748,N_2600);
nand U2963 (N_2963,N_2624,N_2699);
xnor U2964 (N_2964,N_2643,N_2639);
xor U2965 (N_2965,N_2676,N_2723);
nand U2966 (N_2966,N_2665,N_2663);
or U2967 (N_2967,N_2679,N_2681);
or U2968 (N_2968,N_2791,N_2620);
or U2969 (N_2969,N_2699,N_2702);
nand U2970 (N_2970,N_2650,N_2631);
and U2971 (N_2971,N_2757,N_2765);
nor U2972 (N_2972,N_2747,N_2731);
and U2973 (N_2973,N_2726,N_2774);
xor U2974 (N_2974,N_2628,N_2793);
and U2975 (N_2975,N_2703,N_2634);
nand U2976 (N_2976,N_2612,N_2641);
nor U2977 (N_2977,N_2736,N_2601);
nand U2978 (N_2978,N_2701,N_2698);
and U2979 (N_2979,N_2721,N_2750);
or U2980 (N_2980,N_2648,N_2631);
and U2981 (N_2981,N_2745,N_2726);
nand U2982 (N_2982,N_2653,N_2632);
xnor U2983 (N_2983,N_2703,N_2711);
or U2984 (N_2984,N_2785,N_2726);
nand U2985 (N_2985,N_2670,N_2650);
nand U2986 (N_2986,N_2659,N_2605);
nor U2987 (N_2987,N_2756,N_2611);
nand U2988 (N_2988,N_2786,N_2678);
nor U2989 (N_2989,N_2787,N_2612);
nand U2990 (N_2990,N_2667,N_2642);
nand U2991 (N_2991,N_2660,N_2680);
nand U2992 (N_2992,N_2723,N_2654);
and U2993 (N_2993,N_2604,N_2758);
or U2994 (N_2994,N_2659,N_2676);
nor U2995 (N_2995,N_2662,N_2691);
or U2996 (N_2996,N_2767,N_2692);
and U2997 (N_2997,N_2606,N_2718);
and U2998 (N_2998,N_2658,N_2783);
nor U2999 (N_2999,N_2761,N_2759);
nand U3000 (N_3000,N_2970,N_2978);
nand U3001 (N_3001,N_2989,N_2945);
or U3002 (N_3002,N_2943,N_2843);
nor U3003 (N_3003,N_2916,N_2999);
nor U3004 (N_3004,N_2832,N_2966);
nor U3005 (N_3005,N_2904,N_2952);
nor U3006 (N_3006,N_2809,N_2925);
and U3007 (N_3007,N_2860,N_2913);
nand U3008 (N_3008,N_2889,N_2825);
or U3009 (N_3009,N_2956,N_2930);
and U3010 (N_3010,N_2907,N_2990);
nand U3011 (N_3011,N_2880,N_2806);
or U3012 (N_3012,N_2802,N_2982);
xnor U3013 (N_3013,N_2828,N_2941);
and U3014 (N_3014,N_2817,N_2834);
and U3015 (N_3015,N_2897,N_2920);
nand U3016 (N_3016,N_2858,N_2938);
nand U3017 (N_3017,N_2900,N_2993);
nor U3018 (N_3018,N_2912,N_2881);
and U3019 (N_3019,N_2926,N_2879);
and U3020 (N_3020,N_2927,N_2827);
or U3021 (N_3021,N_2837,N_2933);
xnor U3022 (N_3022,N_2923,N_2886);
nand U3023 (N_3023,N_2964,N_2901);
nor U3024 (N_3024,N_2885,N_2844);
and U3025 (N_3025,N_2981,N_2968);
nand U3026 (N_3026,N_2995,N_2852);
nand U3027 (N_3027,N_2895,N_2829);
or U3028 (N_3028,N_2842,N_2838);
and U3029 (N_3029,N_2836,N_2915);
and U3030 (N_3030,N_2877,N_2961);
nand U3031 (N_3031,N_2887,N_2973);
and U3032 (N_3032,N_2822,N_2921);
nor U3033 (N_3033,N_2918,N_2908);
nor U3034 (N_3034,N_2902,N_2816);
or U3035 (N_3035,N_2823,N_2818);
or U3036 (N_3036,N_2849,N_2801);
nor U3037 (N_3037,N_2878,N_2946);
or U3038 (N_3038,N_2924,N_2864);
nand U3039 (N_3039,N_2944,N_2977);
and U3040 (N_3040,N_2991,N_2899);
xnor U3041 (N_3041,N_2866,N_2971);
or U3042 (N_3042,N_2965,N_2988);
nor U3043 (N_3043,N_2875,N_2936);
and U3044 (N_3044,N_2958,N_2969);
nand U3045 (N_3045,N_2857,N_2851);
and U3046 (N_3046,N_2985,N_2975);
and U3047 (N_3047,N_2909,N_2810);
nand U3048 (N_3048,N_2984,N_2986);
nand U3049 (N_3049,N_2859,N_2953);
xor U3050 (N_3050,N_2994,N_2876);
and U3051 (N_3051,N_2951,N_2845);
nand U3052 (N_3052,N_2854,N_2869);
xnor U3053 (N_3053,N_2963,N_2939);
xnor U3054 (N_3054,N_2803,N_2955);
or U3055 (N_3055,N_2932,N_2861);
and U3056 (N_3056,N_2931,N_2959);
nor U3057 (N_3057,N_2898,N_2894);
xor U3058 (N_3058,N_2929,N_2826);
and U3059 (N_3059,N_2811,N_2957);
and U3060 (N_3060,N_2824,N_2884);
nand U3061 (N_3061,N_2808,N_2807);
nor U3062 (N_3062,N_2831,N_2893);
nand U3063 (N_3063,N_2888,N_2983);
or U3064 (N_3064,N_2910,N_2865);
nor U3065 (N_3065,N_2855,N_2804);
nand U3066 (N_3066,N_2867,N_2896);
nor U3067 (N_3067,N_2948,N_2972);
xor U3068 (N_3068,N_2928,N_2976);
nor U3069 (N_3069,N_2820,N_2830);
and U3070 (N_3070,N_2962,N_2868);
nor U3071 (N_3071,N_2814,N_2846);
nor U3072 (N_3072,N_2979,N_2949);
and U3073 (N_3073,N_2874,N_2987);
and U3074 (N_3074,N_2997,N_2891);
or U3075 (N_3075,N_2813,N_2819);
and U3076 (N_3076,N_2892,N_2919);
nor U3077 (N_3077,N_2873,N_2821);
and U3078 (N_3078,N_2940,N_2914);
nand U3079 (N_3079,N_2871,N_2911);
or U3080 (N_3080,N_2870,N_2856);
and U3081 (N_3081,N_2992,N_2950);
xor U3082 (N_3082,N_2998,N_2942);
and U3083 (N_3083,N_2863,N_2922);
xor U3084 (N_3084,N_2996,N_2906);
or U3085 (N_3085,N_2815,N_2890);
nand U3086 (N_3086,N_2882,N_2980);
nor U3087 (N_3087,N_2917,N_2974);
nor U3088 (N_3088,N_2805,N_2903);
nand U3089 (N_3089,N_2883,N_2905);
and U3090 (N_3090,N_2947,N_2833);
and U3091 (N_3091,N_2954,N_2960);
nand U3092 (N_3092,N_2937,N_2853);
nor U3093 (N_3093,N_2935,N_2967);
and U3094 (N_3094,N_2839,N_2862);
xnor U3095 (N_3095,N_2847,N_2850);
xnor U3096 (N_3096,N_2934,N_2840);
or U3097 (N_3097,N_2872,N_2800);
and U3098 (N_3098,N_2841,N_2812);
or U3099 (N_3099,N_2848,N_2835);
and U3100 (N_3100,N_2872,N_2835);
nand U3101 (N_3101,N_2843,N_2859);
nor U3102 (N_3102,N_2954,N_2964);
or U3103 (N_3103,N_2812,N_2871);
or U3104 (N_3104,N_2925,N_2888);
nand U3105 (N_3105,N_2902,N_2805);
and U3106 (N_3106,N_2998,N_2922);
or U3107 (N_3107,N_2983,N_2906);
nand U3108 (N_3108,N_2894,N_2818);
nand U3109 (N_3109,N_2908,N_2956);
and U3110 (N_3110,N_2839,N_2945);
and U3111 (N_3111,N_2921,N_2978);
and U3112 (N_3112,N_2970,N_2902);
and U3113 (N_3113,N_2823,N_2994);
nor U3114 (N_3114,N_2900,N_2809);
and U3115 (N_3115,N_2908,N_2878);
and U3116 (N_3116,N_2812,N_2837);
xnor U3117 (N_3117,N_2950,N_2980);
nor U3118 (N_3118,N_2834,N_2879);
or U3119 (N_3119,N_2898,N_2941);
nand U3120 (N_3120,N_2887,N_2863);
xnor U3121 (N_3121,N_2907,N_2956);
nand U3122 (N_3122,N_2868,N_2872);
or U3123 (N_3123,N_2972,N_2916);
nor U3124 (N_3124,N_2913,N_2800);
nand U3125 (N_3125,N_2825,N_2865);
and U3126 (N_3126,N_2983,N_2901);
nor U3127 (N_3127,N_2893,N_2931);
and U3128 (N_3128,N_2890,N_2995);
and U3129 (N_3129,N_2900,N_2927);
nand U3130 (N_3130,N_2858,N_2968);
nor U3131 (N_3131,N_2805,N_2998);
and U3132 (N_3132,N_2885,N_2888);
nor U3133 (N_3133,N_2975,N_2998);
nor U3134 (N_3134,N_2824,N_2817);
xor U3135 (N_3135,N_2846,N_2852);
or U3136 (N_3136,N_2905,N_2889);
or U3137 (N_3137,N_2812,N_2976);
nor U3138 (N_3138,N_2863,N_2810);
nor U3139 (N_3139,N_2851,N_2883);
xnor U3140 (N_3140,N_2928,N_2815);
and U3141 (N_3141,N_2841,N_2947);
or U3142 (N_3142,N_2965,N_2849);
nand U3143 (N_3143,N_2949,N_2977);
nor U3144 (N_3144,N_2821,N_2870);
and U3145 (N_3145,N_2916,N_2877);
nand U3146 (N_3146,N_2838,N_2853);
nor U3147 (N_3147,N_2846,N_2935);
nor U3148 (N_3148,N_2884,N_2832);
nor U3149 (N_3149,N_2946,N_2882);
nand U3150 (N_3150,N_2927,N_2952);
nor U3151 (N_3151,N_2995,N_2984);
nor U3152 (N_3152,N_2827,N_2904);
or U3153 (N_3153,N_2947,N_2931);
and U3154 (N_3154,N_2800,N_2847);
nor U3155 (N_3155,N_2854,N_2839);
or U3156 (N_3156,N_2886,N_2967);
or U3157 (N_3157,N_2971,N_2943);
nand U3158 (N_3158,N_2941,N_2948);
and U3159 (N_3159,N_2880,N_2918);
nand U3160 (N_3160,N_2970,N_2962);
xor U3161 (N_3161,N_2893,N_2994);
nor U3162 (N_3162,N_2892,N_2890);
nand U3163 (N_3163,N_2838,N_2891);
and U3164 (N_3164,N_2960,N_2963);
or U3165 (N_3165,N_2934,N_2904);
xnor U3166 (N_3166,N_2926,N_2824);
nand U3167 (N_3167,N_2908,N_2945);
and U3168 (N_3168,N_2936,N_2905);
nand U3169 (N_3169,N_2886,N_2862);
nand U3170 (N_3170,N_2871,N_2895);
xnor U3171 (N_3171,N_2855,N_2805);
and U3172 (N_3172,N_2809,N_2898);
xnor U3173 (N_3173,N_2828,N_2933);
nand U3174 (N_3174,N_2846,N_2908);
xor U3175 (N_3175,N_2830,N_2916);
and U3176 (N_3176,N_2811,N_2847);
nor U3177 (N_3177,N_2973,N_2838);
nor U3178 (N_3178,N_2800,N_2946);
nand U3179 (N_3179,N_2874,N_2832);
or U3180 (N_3180,N_2935,N_2958);
or U3181 (N_3181,N_2952,N_2868);
nand U3182 (N_3182,N_2954,N_2945);
and U3183 (N_3183,N_2999,N_2834);
xor U3184 (N_3184,N_2861,N_2940);
nor U3185 (N_3185,N_2831,N_2817);
and U3186 (N_3186,N_2967,N_2960);
nand U3187 (N_3187,N_2878,N_2889);
nand U3188 (N_3188,N_2803,N_2902);
nor U3189 (N_3189,N_2882,N_2862);
or U3190 (N_3190,N_2930,N_2898);
nor U3191 (N_3191,N_2944,N_2824);
nand U3192 (N_3192,N_2942,N_2809);
nor U3193 (N_3193,N_2931,N_2845);
nor U3194 (N_3194,N_2876,N_2816);
or U3195 (N_3195,N_2906,N_2995);
or U3196 (N_3196,N_2966,N_2909);
xnor U3197 (N_3197,N_2928,N_2871);
or U3198 (N_3198,N_2837,N_2921);
xnor U3199 (N_3199,N_2990,N_2846);
nand U3200 (N_3200,N_3054,N_3160);
nand U3201 (N_3201,N_3119,N_3131);
nor U3202 (N_3202,N_3064,N_3129);
nor U3203 (N_3203,N_3145,N_3199);
and U3204 (N_3204,N_3061,N_3031);
nor U3205 (N_3205,N_3185,N_3098);
nand U3206 (N_3206,N_3027,N_3159);
and U3207 (N_3207,N_3150,N_3048);
nand U3208 (N_3208,N_3130,N_3147);
nor U3209 (N_3209,N_3001,N_3075);
nand U3210 (N_3210,N_3095,N_3035);
nand U3211 (N_3211,N_3099,N_3026);
nand U3212 (N_3212,N_3074,N_3132);
nor U3213 (N_3213,N_3154,N_3094);
nand U3214 (N_3214,N_3135,N_3003);
nor U3215 (N_3215,N_3085,N_3175);
and U3216 (N_3216,N_3176,N_3124);
nand U3217 (N_3217,N_3022,N_3179);
nor U3218 (N_3218,N_3170,N_3123);
and U3219 (N_3219,N_3146,N_3080);
and U3220 (N_3220,N_3018,N_3172);
and U3221 (N_3221,N_3013,N_3197);
nand U3222 (N_3222,N_3173,N_3009);
nor U3223 (N_3223,N_3072,N_3189);
and U3224 (N_3224,N_3063,N_3113);
nand U3225 (N_3225,N_3196,N_3036);
nor U3226 (N_3226,N_3010,N_3133);
xnor U3227 (N_3227,N_3115,N_3106);
and U3228 (N_3228,N_3125,N_3062);
xor U3229 (N_3229,N_3069,N_3092);
nand U3230 (N_3230,N_3116,N_3066);
nor U3231 (N_3231,N_3162,N_3177);
and U3232 (N_3232,N_3086,N_3141);
nor U3233 (N_3233,N_3166,N_3011);
and U3234 (N_3234,N_3101,N_3093);
or U3235 (N_3235,N_3077,N_3005);
nand U3236 (N_3236,N_3056,N_3060);
nor U3237 (N_3237,N_3041,N_3078);
and U3238 (N_3238,N_3068,N_3088);
nor U3239 (N_3239,N_3050,N_3030);
nor U3240 (N_3240,N_3169,N_3117);
and U3241 (N_3241,N_3014,N_3070);
and U3242 (N_3242,N_3165,N_3112);
or U3243 (N_3243,N_3023,N_3188);
and U3244 (N_3244,N_3087,N_3126);
nor U3245 (N_3245,N_3082,N_3104);
or U3246 (N_3246,N_3045,N_3178);
nand U3247 (N_3247,N_3127,N_3015);
nor U3248 (N_3248,N_3079,N_3144);
or U3249 (N_3249,N_3037,N_3114);
xor U3250 (N_3250,N_3057,N_3052);
nand U3251 (N_3251,N_3183,N_3090);
or U3252 (N_3252,N_3191,N_3025);
and U3253 (N_3253,N_3134,N_3140);
nand U3254 (N_3254,N_3122,N_3091);
or U3255 (N_3255,N_3164,N_3040);
xor U3256 (N_3256,N_3187,N_3019);
or U3257 (N_3257,N_3065,N_3008);
xnor U3258 (N_3258,N_3024,N_3017);
nand U3259 (N_3259,N_3012,N_3121);
nand U3260 (N_3260,N_3152,N_3136);
or U3261 (N_3261,N_3168,N_3006);
and U3262 (N_3262,N_3181,N_3120);
nand U3263 (N_3263,N_3118,N_3186);
nor U3264 (N_3264,N_3021,N_3097);
nor U3265 (N_3265,N_3167,N_3148);
or U3266 (N_3266,N_3139,N_3156);
and U3267 (N_3267,N_3102,N_3076);
or U3268 (N_3268,N_3034,N_3043);
and U3269 (N_3269,N_3110,N_3157);
nor U3270 (N_3270,N_3096,N_3180);
nor U3271 (N_3271,N_3089,N_3049);
or U3272 (N_3272,N_3109,N_3038);
nor U3273 (N_3273,N_3107,N_3171);
nand U3274 (N_3274,N_3016,N_3149);
nor U3275 (N_3275,N_3111,N_3051);
nand U3276 (N_3276,N_3000,N_3004);
nand U3277 (N_3277,N_3163,N_3184);
nand U3278 (N_3278,N_3059,N_3084);
nand U3279 (N_3279,N_3103,N_3194);
nand U3280 (N_3280,N_3073,N_3046);
xor U3281 (N_3281,N_3020,N_3053);
nand U3282 (N_3282,N_3029,N_3044);
nor U3283 (N_3283,N_3083,N_3193);
nor U3284 (N_3284,N_3100,N_3028);
nor U3285 (N_3285,N_3105,N_3174);
and U3286 (N_3286,N_3081,N_3108);
or U3287 (N_3287,N_3192,N_3190);
nor U3288 (N_3288,N_3067,N_3182);
nor U3289 (N_3289,N_3142,N_3055);
nor U3290 (N_3290,N_3198,N_3161);
xnor U3291 (N_3291,N_3158,N_3195);
or U3292 (N_3292,N_3155,N_3032);
or U3293 (N_3293,N_3002,N_3047);
and U3294 (N_3294,N_3143,N_3151);
xor U3295 (N_3295,N_3153,N_3128);
or U3296 (N_3296,N_3058,N_3033);
and U3297 (N_3297,N_3007,N_3042);
or U3298 (N_3298,N_3071,N_3039);
or U3299 (N_3299,N_3137,N_3138);
or U3300 (N_3300,N_3109,N_3111);
and U3301 (N_3301,N_3068,N_3167);
and U3302 (N_3302,N_3164,N_3194);
nor U3303 (N_3303,N_3196,N_3000);
nand U3304 (N_3304,N_3054,N_3186);
nor U3305 (N_3305,N_3007,N_3006);
nor U3306 (N_3306,N_3111,N_3186);
nand U3307 (N_3307,N_3077,N_3050);
or U3308 (N_3308,N_3030,N_3116);
nor U3309 (N_3309,N_3195,N_3183);
nand U3310 (N_3310,N_3022,N_3003);
nand U3311 (N_3311,N_3083,N_3102);
and U3312 (N_3312,N_3176,N_3000);
and U3313 (N_3313,N_3131,N_3040);
xnor U3314 (N_3314,N_3184,N_3148);
nor U3315 (N_3315,N_3152,N_3046);
or U3316 (N_3316,N_3048,N_3166);
nor U3317 (N_3317,N_3171,N_3074);
nand U3318 (N_3318,N_3139,N_3081);
nand U3319 (N_3319,N_3086,N_3037);
nand U3320 (N_3320,N_3189,N_3105);
nor U3321 (N_3321,N_3139,N_3133);
or U3322 (N_3322,N_3072,N_3095);
nor U3323 (N_3323,N_3172,N_3068);
nand U3324 (N_3324,N_3198,N_3047);
nand U3325 (N_3325,N_3173,N_3016);
and U3326 (N_3326,N_3180,N_3129);
nand U3327 (N_3327,N_3028,N_3157);
or U3328 (N_3328,N_3118,N_3142);
nand U3329 (N_3329,N_3103,N_3046);
nor U3330 (N_3330,N_3089,N_3115);
nor U3331 (N_3331,N_3107,N_3086);
nand U3332 (N_3332,N_3082,N_3101);
nand U3333 (N_3333,N_3055,N_3079);
nand U3334 (N_3334,N_3075,N_3163);
and U3335 (N_3335,N_3025,N_3122);
and U3336 (N_3336,N_3056,N_3087);
xnor U3337 (N_3337,N_3152,N_3145);
xnor U3338 (N_3338,N_3145,N_3178);
nand U3339 (N_3339,N_3156,N_3055);
or U3340 (N_3340,N_3143,N_3127);
and U3341 (N_3341,N_3101,N_3135);
nor U3342 (N_3342,N_3103,N_3085);
or U3343 (N_3343,N_3009,N_3124);
nor U3344 (N_3344,N_3019,N_3106);
and U3345 (N_3345,N_3057,N_3070);
and U3346 (N_3346,N_3177,N_3046);
nand U3347 (N_3347,N_3022,N_3164);
or U3348 (N_3348,N_3118,N_3165);
nor U3349 (N_3349,N_3155,N_3028);
nor U3350 (N_3350,N_3170,N_3060);
and U3351 (N_3351,N_3013,N_3014);
nand U3352 (N_3352,N_3075,N_3005);
and U3353 (N_3353,N_3019,N_3052);
nor U3354 (N_3354,N_3118,N_3062);
nor U3355 (N_3355,N_3084,N_3100);
xnor U3356 (N_3356,N_3015,N_3089);
or U3357 (N_3357,N_3059,N_3035);
or U3358 (N_3358,N_3048,N_3121);
nor U3359 (N_3359,N_3105,N_3155);
nand U3360 (N_3360,N_3084,N_3033);
or U3361 (N_3361,N_3072,N_3129);
and U3362 (N_3362,N_3178,N_3165);
nor U3363 (N_3363,N_3083,N_3144);
nor U3364 (N_3364,N_3179,N_3041);
nor U3365 (N_3365,N_3166,N_3031);
nand U3366 (N_3366,N_3063,N_3029);
nor U3367 (N_3367,N_3056,N_3169);
nor U3368 (N_3368,N_3106,N_3026);
nor U3369 (N_3369,N_3018,N_3184);
nand U3370 (N_3370,N_3034,N_3124);
nor U3371 (N_3371,N_3018,N_3088);
nor U3372 (N_3372,N_3160,N_3109);
or U3373 (N_3373,N_3053,N_3056);
nor U3374 (N_3374,N_3019,N_3058);
xnor U3375 (N_3375,N_3170,N_3198);
or U3376 (N_3376,N_3095,N_3081);
or U3377 (N_3377,N_3042,N_3012);
nor U3378 (N_3378,N_3024,N_3101);
nand U3379 (N_3379,N_3083,N_3015);
or U3380 (N_3380,N_3067,N_3148);
nor U3381 (N_3381,N_3179,N_3029);
nor U3382 (N_3382,N_3006,N_3023);
and U3383 (N_3383,N_3061,N_3058);
or U3384 (N_3384,N_3170,N_3161);
or U3385 (N_3385,N_3068,N_3164);
nor U3386 (N_3386,N_3143,N_3188);
and U3387 (N_3387,N_3032,N_3103);
or U3388 (N_3388,N_3184,N_3174);
nor U3389 (N_3389,N_3177,N_3107);
xnor U3390 (N_3390,N_3180,N_3146);
and U3391 (N_3391,N_3076,N_3161);
or U3392 (N_3392,N_3146,N_3015);
and U3393 (N_3393,N_3053,N_3188);
nor U3394 (N_3394,N_3001,N_3027);
nor U3395 (N_3395,N_3085,N_3094);
nand U3396 (N_3396,N_3189,N_3199);
nor U3397 (N_3397,N_3139,N_3105);
nor U3398 (N_3398,N_3163,N_3097);
xnor U3399 (N_3399,N_3175,N_3109);
and U3400 (N_3400,N_3244,N_3222);
and U3401 (N_3401,N_3344,N_3290);
and U3402 (N_3402,N_3300,N_3355);
nand U3403 (N_3403,N_3346,N_3238);
nor U3404 (N_3404,N_3339,N_3280);
nand U3405 (N_3405,N_3377,N_3310);
nor U3406 (N_3406,N_3374,N_3365);
or U3407 (N_3407,N_3240,N_3252);
nor U3408 (N_3408,N_3215,N_3242);
nand U3409 (N_3409,N_3376,N_3316);
nand U3410 (N_3410,N_3314,N_3375);
and U3411 (N_3411,N_3286,N_3273);
nor U3412 (N_3412,N_3358,N_3330);
or U3413 (N_3413,N_3337,N_3216);
or U3414 (N_3414,N_3380,N_3379);
and U3415 (N_3415,N_3317,N_3345);
xor U3416 (N_3416,N_3236,N_3213);
nand U3417 (N_3417,N_3299,N_3385);
xor U3418 (N_3418,N_3292,N_3205);
or U3419 (N_3419,N_3207,N_3361);
and U3420 (N_3420,N_3201,N_3264);
or U3421 (N_3421,N_3396,N_3382);
nor U3422 (N_3422,N_3306,N_3234);
and U3423 (N_3423,N_3217,N_3383);
and U3424 (N_3424,N_3232,N_3325);
nor U3425 (N_3425,N_3359,N_3363);
nand U3426 (N_3426,N_3334,N_3392);
nand U3427 (N_3427,N_3348,N_3308);
nor U3428 (N_3428,N_3356,N_3397);
nor U3429 (N_3429,N_3351,N_3303);
or U3430 (N_3430,N_3386,N_3218);
nor U3431 (N_3431,N_3388,N_3338);
and U3432 (N_3432,N_3319,N_3241);
xor U3433 (N_3433,N_3393,N_3258);
nand U3434 (N_3434,N_3212,N_3221);
and U3435 (N_3435,N_3279,N_3272);
xnor U3436 (N_3436,N_3209,N_3343);
nand U3437 (N_3437,N_3259,N_3384);
xnor U3438 (N_3438,N_3387,N_3277);
nand U3439 (N_3439,N_3247,N_3210);
xor U3440 (N_3440,N_3285,N_3246);
and U3441 (N_3441,N_3267,N_3233);
or U3442 (N_3442,N_3239,N_3318);
nand U3443 (N_3443,N_3371,N_3260);
and U3444 (N_3444,N_3200,N_3288);
nor U3445 (N_3445,N_3326,N_3224);
or U3446 (N_3446,N_3274,N_3322);
and U3447 (N_3447,N_3296,N_3328);
nor U3448 (N_3448,N_3219,N_3204);
or U3449 (N_3449,N_3263,N_3255);
and U3450 (N_3450,N_3270,N_3243);
and U3451 (N_3451,N_3305,N_3271);
and U3452 (N_3452,N_3366,N_3336);
and U3453 (N_3453,N_3323,N_3320);
nor U3454 (N_3454,N_3342,N_3329);
and U3455 (N_3455,N_3381,N_3294);
xor U3456 (N_3456,N_3235,N_3269);
or U3457 (N_3457,N_3226,N_3291);
or U3458 (N_3458,N_3354,N_3253);
nand U3459 (N_3459,N_3257,N_3298);
or U3460 (N_3460,N_3256,N_3262);
nand U3461 (N_3461,N_3208,N_3333);
or U3462 (N_3462,N_3254,N_3399);
xnor U3463 (N_3463,N_3282,N_3357);
or U3464 (N_3464,N_3349,N_3370);
nand U3465 (N_3465,N_3227,N_3304);
and U3466 (N_3466,N_3225,N_3341);
nand U3467 (N_3467,N_3367,N_3289);
nand U3468 (N_3468,N_3315,N_3228);
nor U3469 (N_3469,N_3331,N_3332);
nand U3470 (N_3470,N_3364,N_3245);
or U3471 (N_3471,N_3395,N_3261);
nor U3472 (N_3472,N_3220,N_3312);
nand U3473 (N_3473,N_3327,N_3266);
or U3474 (N_3474,N_3284,N_3302);
nor U3475 (N_3475,N_3350,N_3206);
or U3476 (N_3476,N_3311,N_3237);
nor U3477 (N_3477,N_3268,N_3251);
or U3478 (N_3478,N_3307,N_3276);
or U3479 (N_3479,N_3394,N_3214);
and U3480 (N_3480,N_3278,N_3369);
and U3481 (N_3481,N_3301,N_3373);
or U3482 (N_3482,N_3229,N_3353);
nand U3483 (N_3483,N_3295,N_3321);
or U3484 (N_3484,N_3230,N_3390);
nor U3485 (N_3485,N_3293,N_3203);
nor U3486 (N_3486,N_3249,N_3340);
nand U3487 (N_3487,N_3324,N_3211);
xor U3488 (N_3488,N_3283,N_3309);
and U3489 (N_3489,N_3378,N_3313);
nand U3490 (N_3490,N_3202,N_3297);
or U3491 (N_3491,N_3281,N_3287);
xor U3492 (N_3492,N_3389,N_3362);
nand U3493 (N_3493,N_3391,N_3275);
or U3494 (N_3494,N_3231,N_3223);
nor U3495 (N_3495,N_3360,N_3335);
and U3496 (N_3496,N_3398,N_3347);
nor U3497 (N_3497,N_3250,N_3352);
nor U3498 (N_3498,N_3372,N_3265);
xnor U3499 (N_3499,N_3248,N_3368);
nor U3500 (N_3500,N_3376,N_3309);
nor U3501 (N_3501,N_3369,N_3275);
or U3502 (N_3502,N_3305,N_3328);
nor U3503 (N_3503,N_3339,N_3287);
nor U3504 (N_3504,N_3237,N_3352);
nor U3505 (N_3505,N_3343,N_3321);
or U3506 (N_3506,N_3353,N_3271);
nor U3507 (N_3507,N_3223,N_3349);
or U3508 (N_3508,N_3377,N_3206);
nand U3509 (N_3509,N_3343,N_3274);
and U3510 (N_3510,N_3287,N_3302);
nand U3511 (N_3511,N_3280,N_3216);
or U3512 (N_3512,N_3310,N_3347);
and U3513 (N_3513,N_3327,N_3382);
or U3514 (N_3514,N_3211,N_3248);
or U3515 (N_3515,N_3383,N_3340);
nand U3516 (N_3516,N_3363,N_3330);
nand U3517 (N_3517,N_3321,N_3210);
nor U3518 (N_3518,N_3399,N_3332);
or U3519 (N_3519,N_3279,N_3335);
xnor U3520 (N_3520,N_3252,N_3385);
and U3521 (N_3521,N_3270,N_3373);
nor U3522 (N_3522,N_3200,N_3315);
or U3523 (N_3523,N_3250,N_3312);
nand U3524 (N_3524,N_3227,N_3263);
nand U3525 (N_3525,N_3211,N_3381);
nor U3526 (N_3526,N_3377,N_3254);
nand U3527 (N_3527,N_3217,N_3291);
and U3528 (N_3528,N_3208,N_3311);
nor U3529 (N_3529,N_3390,N_3355);
and U3530 (N_3530,N_3212,N_3279);
xor U3531 (N_3531,N_3351,N_3382);
and U3532 (N_3532,N_3282,N_3204);
and U3533 (N_3533,N_3249,N_3338);
nand U3534 (N_3534,N_3343,N_3386);
and U3535 (N_3535,N_3396,N_3298);
nor U3536 (N_3536,N_3389,N_3297);
nor U3537 (N_3537,N_3284,N_3351);
and U3538 (N_3538,N_3359,N_3261);
xnor U3539 (N_3539,N_3303,N_3252);
nand U3540 (N_3540,N_3269,N_3307);
and U3541 (N_3541,N_3288,N_3372);
and U3542 (N_3542,N_3289,N_3248);
nor U3543 (N_3543,N_3240,N_3272);
xor U3544 (N_3544,N_3394,N_3285);
nor U3545 (N_3545,N_3289,N_3388);
or U3546 (N_3546,N_3320,N_3387);
nor U3547 (N_3547,N_3365,N_3345);
nand U3548 (N_3548,N_3247,N_3369);
nor U3549 (N_3549,N_3256,N_3320);
or U3550 (N_3550,N_3372,N_3246);
nand U3551 (N_3551,N_3245,N_3246);
xnor U3552 (N_3552,N_3318,N_3313);
or U3553 (N_3553,N_3273,N_3284);
nor U3554 (N_3554,N_3361,N_3315);
nor U3555 (N_3555,N_3238,N_3200);
nand U3556 (N_3556,N_3239,N_3326);
xor U3557 (N_3557,N_3260,N_3390);
or U3558 (N_3558,N_3270,N_3290);
nor U3559 (N_3559,N_3348,N_3350);
nor U3560 (N_3560,N_3235,N_3229);
nand U3561 (N_3561,N_3329,N_3321);
and U3562 (N_3562,N_3357,N_3216);
nor U3563 (N_3563,N_3279,N_3259);
nor U3564 (N_3564,N_3316,N_3261);
or U3565 (N_3565,N_3260,N_3388);
xnor U3566 (N_3566,N_3323,N_3314);
and U3567 (N_3567,N_3271,N_3262);
nand U3568 (N_3568,N_3360,N_3225);
nor U3569 (N_3569,N_3254,N_3350);
and U3570 (N_3570,N_3331,N_3205);
or U3571 (N_3571,N_3236,N_3357);
and U3572 (N_3572,N_3246,N_3391);
nand U3573 (N_3573,N_3349,N_3282);
nand U3574 (N_3574,N_3200,N_3383);
nand U3575 (N_3575,N_3284,N_3357);
nand U3576 (N_3576,N_3378,N_3206);
nor U3577 (N_3577,N_3300,N_3361);
xnor U3578 (N_3578,N_3233,N_3220);
nor U3579 (N_3579,N_3287,N_3249);
or U3580 (N_3580,N_3359,N_3243);
and U3581 (N_3581,N_3281,N_3384);
xor U3582 (N_3582,N_3399,N_3347);
nand U3583 (N_3583,N_3263,N_3341);
xnor U3584 (N_3584,N_3214,N_3393);
nor U3585 (N_3585,N_3379,N_3225);
or U3586 (N_3586,N_3339,N_3201);
and U3587 (N_3587,N_3308,N_3313);
nand U3588 (N_3588,N_3346,N_3378);
nand U3589 (N_3589,N_3215,N_3356);
and U3590 (N_3590,N_3210,N_3350);
nand U3591 (N_3591,N_3289,N_3233);
nand U3592 (N_3592,N_3209,N_3332);
or U3593 (N_3593,N_3324,N_3303);
and U3594 (N_3594,N_3230,N_3207);
or U3595 (N_3595,N_3203,N_3261);
nand U3596 (N_3596,N_3299,N_3312);
or U3597 (N_3597,N_3289,N_3288);
xnor U3598 (N_3598,N_3380,N_3230);
or U3599 (N_3599,N_3279,N_3246);
and U3600 (N_3600,N_3592,N_3532);
nor U3601 (N_3601,N_3490,N_3403);
and U3602 (N_3602,N_3414,N_3440);
nand U3603 (N_3603,N_3436,N_3428);
or U3604 (N_3604,N_3559,N_3424);
or U3605 (N_3605,N_3519,N_3509);
and U3606 (N_3606,N_3420,N_3516);
and U3607 (N_3607,N_3419,N_3580);
nand U3608 (N_3608,N_3571,N_3520);
and U3609 (N_3609,N_3437,N_3574);
nand U3610 (N_3610,N_3470,N_3487);
and U3611 (N_3611,N_3449,N_3493);
nand U3612 (N_3612,N_3471,N_3538);
or U3613 (N_3613,N_3466,N_3503);
or U3614 (N_3614,N_3542,N_3517);
or U3615 (N_3615,N_3569,N_3443);
xnor U3616 (N_3616,N_3429,N_3441);
or U3617 (N_3617,N_3557,N_3410);
xor U3618 (N_3618,N_3453,N_3474);
and U3619 (N_3619,N_3537,N_3423);
or U3620 (N_3620,N_3550,N_3467);
nor U3621 (N_3621,N_3568,N_3552);
or U3622 (N_3622,N_3581,N_3402);
or U3623 (N_3623,N_3450,N_3457);
nor U3624 (N_3624,N_3444,N_3448);
and U3625 (N_3625,N_3535,N_3515);
or U3626 (N_3626,N_3475,N_3540);
or U3627 (N_3627,N_3502,N_3521);
xnor U3628 (N_3628,N_3417,N_3587);
nand U3629 (N_3629,N_3489,N_3539);
or U3630 (N_3630,N_3590,N_3563);
and U3631 (N_3631,N_3480,N_3597);
nand U3632 (N_3632,N_3485,N_3473);
nand U3633 (N_3633,N_3551,N_3585);
and U3634 (N_3634,N_3459,N_3479);
nor U3635 (N_3635,N_3577,N_3579);
or U3636 (N_3636,N_3456,N_3598);
or U3637 (N_3637,N_3591,N_3483);
and U3638 (N_3638,N_3566,N_3472);
xor U3639 (N_3639,N_3536,N_3560);
nor U3640 (N_3640,N_3511,N_3492);
nand U3641 (N_3641,N_3561,N_3405);
and U3642 (N_3642,N_3596,N_3458);
nor U3643 (N_3643,N_3496,N_3506);
nand U3644 (N_3644,N_3501,N_3488);
nand U3645 (N_3645,N_3484,N_3546);
nor U3646 (N_3646,N_3527,N_3504);
and U3647 (N_3647,N_3460,N_3524);
or U3648 (N_3648,N_3500,N_3469);
nand U3649 (N_3649,N_3461,N_3576);
or U3650 (N_3650,N_3434,N_3442);
and U3651 (N_3651,N_3553,N_3478);
or U3652 (N_3652,N_3599,N_3523);
and U3653 (N_3653,N_3486,N_3530);
nor U3654 (N_3654,N_3400,N_3505);
or U3655 (N_3655,N_3401,N_3541);
xnor U3656 (N_3656,N_3575,N_3452);
or U3657 (N_3657,N_3499,N_3558);
or U3658 (N_3658,N_3513,N_3462);
and U3659 (N_3659,N_3578,N_3431);
and U3660 (N_3660,N_3545,N_3404);
nand U3661 (N_3661,N_3407,N_3421);
nand U3662 (N_3662,N_3565,N_3432);
and U3663 (N_3663,N_3481,N_3588);
and U3664 (N_3664,N_3507,N_3548);
nor U3665 (N_3665,N_3512,N_3495);
or U3666 (N_3666,N_3584,N_3439);
nand U3667 (N_3667,N_3547,N_3451);
or U3668 (N_3668,N_3593,N_3589);
nand U3669 (N_3669,N_3531,N_3427);
and U3670 (N_3670,N_3433,N_3562);
and U3671 (N_3671,N_3465,N_3556);
nand U3672 (N_3672,N_3518,N_3415);
nand U3673 (N_3673,N_3544,N_3594);
or U3674 (N_3674,N_3426,N_3416);
and U3675 (N_3675,N_3543,N_3438);
nor U3676 (N_3676,N_3406,N_3570);
and U3677 (N_3677,N_3583,N_3464);
and U3678 (N_3678,N_3555,N_3476);
xor U3679 (N_3679,N_3573,N_3510);
and U3680 (N_3680,N_3554,N_3408);
nand U3681 (N_3681,N_3447,N_3411);
xor U3682 (N_3682,N_3413,N_3497);
nand U3683 (N_3683,N_3491,N_3468);
xnor U3684 (N_3684,N_3477,N_3430);
and U3685 (N_3685,N_3567,N_3522);
and U3686 (N_3686,N_3463,N_3435);
nand U3687 (N_3687,N_3454,N_3528);
or U3688 (N_3688,N_3482,N_3525);
and U3689 (N_3689,N_3494,N_3526);
nor U3690 (N_3690,N_3508,N_3564);
and U3691 (N_3691,N_3425,N_3412);
or U3692 (N_3692,N_3533,N_3409);
nand U3693 (N_3693,N_3498,N_3529);
nor U3694 (N_3694,N_3549,N_3586);
or U3695 (N_3695,N_3514,N_3418);
and U3696 (N_3696,N_3534,N_3582);
and U3697 (N_3697,N_3455,N_3422);
or U3698 (N_3698,N_3572,N_3445);
xor U3699 (N_3699,N_3595,N_3446);
nor U3700 (N_3700,N_3408,N_3421);
and U3701 (N_3701,N_3449,N_3434);
nand U3702 (N_3702,N_3583,N_3404);
or U3703 (N_3703,N_3557,N_3409);
or U3704 (N_3704,N_3425,N_3518);
and U3705 (N_3705,N_3581,N_3432);
and U3706 (N_3706,N_3418,N_3599);
nand U3707 (N_3707,N_3416,N_3585);
or U3708 (N_3708,N_3503,N_3432);
nand U3709 (N_3709,N_3525,N_3424);
nand U3710 (N_3710,N_3402,N_3575);
nor U3711 (N_3711,N_3412,N_3487);
nor U3712 (N_3712,N_3518,N_3483);
and U3713 (N_3713,N_3435,N_3508);
or U3714 (N_3714,N_3555,N_3425);
or U3715 (N_3715,N_3519,N_3401);
nand U3716 (N_3716,N_3493,N_3404);
nand U3717 (N_3717,N_3587,N_3566);
and U3718 (N_3718,N_3532,N_3599);
and U3719 (N_3719,N_3428,N_3588);
nor U3720 (N_3720,N_3561,N_3558);
nand U3721 (N_3721,N_3457,N_3493);
and U3722 (N_3722,N_3471,N_3559);
nor U3723 (N_3723,N_3516,N_3422);
xnor U3724 (N_3724,N_3495,N_3541);
and U3725 (N_3725,N_3498,N_3516);
and U3726 (N_3726,N_3513,N_3508);
xnor U3727 (N_3727,N_3455,N_3549);
and U3728 (N_3728,N_3477,N_3537);
xor U3729 (N_3729,N_3453,N_3446);
and U3730 (N_3730,N_3591,N_3571);
and U3731 (N_3731,N_3569,N_3565);
or U3732 (N_3732,N_3405,N_3514);
or U3733 (N_3733,N_3463,N_3456);
or U3734 (N_3734,N_3559,N_3423);
nand U3735 (N_3735,N_3552,N_3510);
and U3736 (N_3736,N_3426,N_3597);
nor U3737 (N_3737,N_3504,N_3595);
and U3738 (N_3738,N_3580,N_3539);
and U3739 (N_3739,N_3596,N_3549);
nor U3740 (N_3740,N_3428,N_3557);
xor U3741 (N_3741,N_3598,N_3532);
nor U3742 (N_3742,N_3434,N_3560);
and U3743 (N_3743,N_3569,N_3429);
nand U3744 (N_3744,N_3490,N_3488);
nand U3745 (N_3745,N_3439,N_3476);
or U3746 (N_3746,N_3598,N_3594);
or U3747 (N_3747,N_3580,N_3404);
nor U3748 (N_3748,N_3496,N_3409);
and U3749 (N_3749,N_3504,N_3513);
and U3750 (N_3750,N_3438,N_3465);
nor U3751 (N_3751,N_3563,N_3427);
nand U3752 (N_3752,N_3458,N_3515);
and U3753 (N_3753,N_3445,N_3543);
nand U3754 (N_3754,N_3402,N_3522);
nand U3755 (N_3755,N_3467,N_3477);
nor U3756 (N_3756,N_3547,N_3430);
and U3757 (N_3757,N_3586,N_3433);
nand U3758 (N_3758,N_3588,N_3545);
or U3759 (N_3759,N_3517,N_3432);
nand U3760 (N_3760,N_3557,N_3443);
and U3761 (N_3761,N_3449,N_3571);
nand U3762 (N_3762,N_3506,N_3578);
nor U3763 (N_3763,N_3551,N_3577);
nor U3764 (N_3764,N_3582,N_3570);
nor U3765 (N_3765,N_3402,N_3513);
and U3766 (N_3766,N_3424,N_3539);
nand U3767 (N_3767,N_3470,N_3555);
nor U3768 (N_3768,N_3580,N_3413);
or U3769 (N_3769,N_3529,N_3421);
xnor U3770 (N_3770,N_3440,N_3538);
and U3771 (N_3771,N_3590,N_3425);
xnor U3772 (N_3772,N_3520,N_3409);
nand U3773 (N_3773,N_3562,N_3592);
or U3774 (N_3774,N_3432,N_3567);
and U3775 (N_3775,N_3560,N_3523);
nor U3776 (N_3776,N_3429,N_3424);
nand U3777 (N_3777,N_3469,N_3418);
xor U3778 (N_3778,N_3539,N_3493);
nand U3779 (N_3779,N_3429,N_3457);
nor U3780 (N_3780,N_3544,N_3470);
nand U3781 (N_3781,N_3421,N_3478);
nand U3782 (N_3782,N_3582,N_3590);
and U3783 (N_3783,N_3579,N_3546);
nor U3784 (N_3784,N_3420,N_3592);
and U3785 (N_3785,N_3499,N_3495);
nor U3786 (N_3786,N_3406,N_3474);
nor U3787 (N_3787,N_3513,N_3490);
xor U3788 (N_3788,N_3566,N_3572);
xor U3789 (N_3789,N_3453,N_3471);
xor U3790 (N_3790,N_3540,N_3410);
nand U3791 (N_3791,N_3560,N_3597);
nor U3792 (N_3792,N_3522,N_3452);
nor U3793 (N_3793,N_3539,N_3497);
nand U3794 (N_3794,N_3432,N_3544);
and U3795 (N_3795,N_3416,N_3436);
xnor U3796 (N_3796,N_3580,N_3432);
nand U3797 (N_3797,N_3405,N_3559);
or U3798 (N_3798,N_3488,N_3527);
and U3799 (N_3799,N_3466,N_3401);
nand U3800 (N_3800,N_3615,N_3665);
and U3801 (N_3801,N_3625,N_3607);
xnor U3802 (N_3802,N_3727,N_3749);
and U3803 (N_3803,N_3734,N_3648);
and U3804 (N_3804,N_3650,N_3758);
nand U3805 (N_3805,N_3671,N_3610);
nand U3806 (N_3806,N_3673,N_3604);
nand U3807 (N_3807,N_3757,N_3747);
xor U3808 (N_3808,N_3643,N_3627);
nand U3809 (N_3809,N_3759,N_3651);
nand U3810 (N_3810,N_3737,N_3623);
nor U3811 (N_3811,N_3751,N_3755);
nor U3812 (N_3812,N_3660,N_3675);
nand U3813 (N_3813,N_3775,N_3646);
nor U3814 (N_3814,N_3666,N_3799);
or U3815 (N_3815,N_3794,N_3601);
nor U3816 (N_3816,N_3782,N_3700);
or U3817 (N_3817,N_3765,N_3622);
nor U3818 (N_3818,N_3715,N_3752);
or U3819 (N_3819,N_3743,N_3729);
and U3820 (N_3820,N_3707,N_3712);
and U3821 (N_3821,N_3656,N_3770);
nand U3822 (N_3822,N_3611,N_3753);
and U3823 (N_3823,N_3696,N_3710);
nand U3824 (N_3824,N_3781,N_3699);
nand U3825 (N_3825,N_3687,N_3620);
and U3826 (N_3826,N_3686,N_3603);
nand U3827 (N_3827,N_3606,N_3621);
nand U3828 (N_3828,N_3684,N_3702);
nor U3829 (N_3829,N_3719,N_3787);
xor U3830 (N_3830,N_3750,N_3632);
nor U3831 (N_3831,N_3798,N_3640);
nor U3832 (N_3832,N_3780,N_3733);
and U3833 (N_3833,N_3630,N_3756);
or U3834 (N_3834,N_3754,N_3681);
nor U3835 (N_3835,N_3642,N_3677);
or U3836 (N_3836,N_3792,N_3772);
nor U3837 (N_3837,N_3773,N_3645);
nor U3838 (N_3838,N_3689,N_3626);
or U3839 (N_3839,N_3631,N_3669);
nand U3840 (N_3840,N_3616,N_3716);
nor U3841 (N_3841,N_3768,N_3653);
or U3842 (N_3842,N_3634,N_3786);
and U3843 (N_3843,N_3670,N_3676);
and U3844 (N_3844,N_3738,N_3682);
and U3845 (N_3845,N_3614,N_3746);
nor U3846 (N_3846,N_3736,N_3748);
xor U3847 (N_3847,N_3629,N_3641);
xor U3848 (N_3848,N_3723,N_3718);
nand U3849 (N_3849,N_3732,N_3709);
nand U3850 (N_3850,N_3674,N_3722);
nor U3851 (N_3851,N_3694,N_3761);
nand U3852 (N_3852,N_3658,N_3654);
or U3853 (N_3853,N_3708,N_3667);
and U3854 (N_3854,N_3778,N_3793);
and U3855 (N_3855,N_3662,N_3672);
nor U3856 (N_3856,N_3647,N_3698);
nand U3857 (N_3857,N_3659,N_3697);
nand U3858 (N_3858,N_3764,N_3766);
or U3859 (N_3859,N_3638,N_3726);
nor U3860 (N_3860,N_3609,N_3649);
or U3861 (N_3861,N_3714,N_3791);
nand U3862 (N_3862,N_3763,N_3668);
and U3863 (N_3863,N_3652,N_3717);
and U3864 (N_3864,N_3613,N_3636);
xor U3865 (N_3865,N_3600,N_3612);
nand U3866 (N_3866,N_3692,N_3602);
nand U3867 (N_3867,N_3691,N_3628);
nor U3868 (N_3868,N_3661,N_3678);
nor U3869 (N_3869,N_3739,N_3774);
nor U3870 (N_3870,N_3725,N_3742);
or U3871 (N_3871,N_3769,N_3663);
nor U3872 (N_3872,N_3728,N_3619);
nand U3873 (N_3873,N_3796,N_3703);
or U3874 (N_3874,N_3771,N_3635);
nand U3875 (N_3875,N_3701,N_3741);
xor U3876 (N_3876,N_3711,N_3618);
or U3877 (N_3877,N_3784,N_3724);
and U3878 (N_3878,N_3767,N_3680);
or U3879 (N_3879,N_3788,N_3633);
or U3880 (N_3880,N_3617,N_3720);
and U3881 (N_3881,N_3608,N_3605);
xor U3882 (N_3882,N_3679,N_3657);
or U3883 (N_3883,N_3745,N_3644);
nand U3884 (N_3884,N_3695,N_3683);
or U3885 (N_3885,N_3779,N_3705);
or U3886 (N_3886,N_3713,N_3740);
nor U3887 (N_3887,N_3730,N_3797);
or U3888 (N_3888,N_3688,N_3685);
nand U3889 (N_3889,N_3690,N_3637);
or U3890 (N_3890,N_3789,N_3731);
and U3891 (N_3891,N_3655,N_3783);
nor U3892 (N_3892,N_3664,N_3777);
or U3893 (N_3893,N_3785,N_3776);
xnor U3894 (N_3894,N_3762,N_3624);
or U3895 (N_3895,N_3735,N_3790);
and U3896 (N_3896,N_3704,N_3721);
xor U3897 (N_3897,N_3760,N_3795);
nor U3898 (N_3898,N_3744,N_3639);
nand U3899 (N_3899,N_3693,N_3706);
nand U3900 (N_3900,N_3662,N_3600);
nor U3901 (N_3901,N_3685,N_3752);
xnor U3902 (N_3902,N_3771,N_3673);
and U3903 (N_3903,N_3662,N_3799);
and U3904 (N_3904,N_3730,N_3690);
or U3905 (N_3905,N_3761,N_3632);
nand U3906 (N_3906,N_3706,N_3602);
or U3907 (N_3907,N_3615,N_3799);
nand U3908 (N_3908,N_3729,N_3740);
nor U3909 (N_3909,N_3633,N_3678);
or U3910 (N_3910,N_3680,N_3783);
and U3911 (N_3911,N_3617,N_3717);
xnor U3912 (N_3912,N_3700,N_3653);
nor U3913 (N_3913,N_3623,N_3618);
and U3914 (N_3914,N_3605,N_3733);
and U3915 (N_3915,N_3637,N_3614);
or U3916 (N_3916,N_3723,N_3740);
nand U3917 (N_3917,N_3617,N_3619);
nand U3918 (N_3918,N_3603,N_3724);
nor U3919 (N_3919,N_3738,N_3679);
xnor U3920 (N_3920,N_3680,N_3768);
and U3921 (N_3921,N_3722,N_3610);
or U3922 (N_3922,N_3718,N_3681);
or U3923 (N_3923,N_3757,N_3701);
nand U3924 (N_3924,N_3689,N_3607);
and U3925 (N_3925,N_3655,N_3761);
and U3926 (N_3926,N_3675,N_3679);
or U3927 (N_3927,N_3730,N_3705);
and U3928 (N_3928,N_3725,N_3681);
nor U3929 (N_3929,N_3670,N_3797);
xnor U3930 (N_3930,N_3644,N_3617);
nor U3931 (N_3931,N_3779,N_3668);
nand U3932 (N_3932,N_3759,N_3641);
nand U3933 (N_3933,N_3605,N_3678);
nand U3934 (N_3934,N_3611,N_3738);
and U3935 (N_3935,N_3638,N_3797);
or U3936 (N_3936,N_3762,N_3640);
or U3937 (N_3937,N_3681,N_3624);
and U3938 (N_3938,N_3695,N_3756);
nand U3939 (N_3939,N_3768,N_3708);
and U3940 (N_3940,N_3676,N_3733);
nand U3941 (N_3941,N_3600,N_3717);
nand U3942 (N_3942,N_3746,N_3747);
nand U3943 (N_3943,N_3707,N_3769);
or U3944 (N_3944,N_3708,N_3674);
nand U3945 (N_3945,N_3611,N_3706);
nor U3946 (N_3946,N_3661,N_3675);
nor U3947 (N_3947,N_3630,N_3682);
nand U3948 (N_3948,N_3699,N_3790);
nand U3949 (N_3949,N_3702,N_3606);
nor U3950 (N_3950,N_3727,N_3710);
xnor U3951 (N_3951,N_3621,N_3752);
and U3952 (N_3952,N_3664,N_3610);
nand U3953 (N_3953,N_3782,N_3655);
nor U3954 (N_3954,N_3779,N_3790);
and U3955 (N_3955,N_3635,N_3668);
and U3956 (N_3956,N_3604,N_3716);
nand U3957 (N_3957,N_3680,N_3762);
nand U3958 (N_3958,N_3697,N_3647);
nand U3959 (N_3959,N_3637,N_3600);
or U3960 (N_3960,N_3606,N_3624);
nor U3961 (N_3961,N_3647,N_3754);
and U3962 (N_3962,N_3629,N_3645);
nand U3963 (N_3963,N_3687,N_3759);
and U3964 (N_3964,N_3734,N_3752);
nor U3965 (N_3965,N_3771,N_3703);
and U3966 (N_3966,N_3764,N_3757);
nand U3967 (N_3967,N_3742,N_3697);
and U3968 (N_3968,N_3625,N_3777);
xor U3969 (N_3969,N_3766,N_3735);
nor U3970 (N_3970,N_3756,N_3768);
or U3971 (N_3971,N_3769,N_3633);
xnor U3972 (N_3972,N_3631,N_3612);
and U3973 (N_3973,N_3778,N_3690);
or U3974 (N_3974,N_3673,N_3723);
nand U3975 (N_3975,N_3626,N_3601);
and U3976 (N_3976,N_3712,N_3602);
nand U3977 (N_3977,N_3740,N_3773);
xnor U3978 (N_3978,N_3600,N_3755);
and U3979 (N_3979,N_3729,N_3783);
nor U3980 (N_3980,N_3730,N_3694);
xor U3981 (N_3981,N_3783,N_3728);
nor U3982 (N_3982,N_3708,N_3704);
nand U3983 (N_3983,N_3649,N_3617);
nor U3984 (N_3984,N_3674,N_3698);
and U3985 (N_3985,N_3628,N_3721);
nor U3986 (N_3986,N_3614,N_3710);
nand U3987 (N_3987,N_3775,N_3774);
or U3988 (N_3988,N_3693,N_3722);
and U3989 (N_3989,N_3615,N_3621);
nor U3990 (N_3990,N_3776,N_3778);
nand U3991 (N_3991,N_3693,N_3716);
or U3992 (N_3992,N_3635,N_3678);
and U3993 (N_3993,N_3713,N_3785);
nand U3994 (N_3994,N_3788,N_3664);
nor U3995 (N_3995,N_3713,N_3647);
and U3996 (N_3996,N_3724,N_3699);
nand U3997 (N_3997,N_3770,N_3732);
nand U3998 (N_3998,N_3782,N_3759);
and U3999 (N_3999,N_3617,N_3636);
and U4000 (N_4000,N_3842,N_3962);
nor U4001 (N_4001,N_3990,N_3883);
nand U4002 (N_4002,N_3820,N_3843);
and U4003 (N_4003,N_3948,N_3933);
nor U4004 (N_4004,N_3874,N_3804);
and U4005 (N_4005,N_3973,N_3960);
and U4006 (N_4006,N_3997,N_3868);
or U4007 (N_4007,N_3993,N_3958);
nand U4008 (N_4008,N_3979,N_3952);
nand U4009 (N_4009,N_3827,N_3940);
or U4010 (N_4010,N_3896,N_3935);
nand U4011 (N_4011,N_3850,N_3999);
and U4012 (N_4012,N_3967,N_3964);
nor U4013 (N_4013,N_3877,N_3888);
xnor U4014 (N_4014,N_3972,N_3801);
xor U4015 (N_4015,N_3969,N_3884);
nand U4016 (N_4016,N_3938,N_3898);
or U4017 (N_4017,N_3899,N_3986);
nand U4018 (N_4018,N_3936,N_3988);
and U4019 (N_4019,N_3816,N_3907);
and U4020 (N_4020,N_3808,N_3859);
nor U4021 (N_4021,N_3949,N_3920);
nand U4022 (N_4022,N_3814,N_3873);
and U4023 (N_4023,N_3974,N_3856);
or U4024 (N_4024,N_3844,N_3824);
and U4025 (N_4025,N_3869,N_3942);
nor U4026 (N_4026,N_3803,N_3832);
or U4027 (N_4027,N_3980,N_3911);
and U4028 (N_4028,N_3914,N_3845);
and U4029 (N_4029,N_3866,N_3813);
nor U4030 (N_4030,N_3860,N_3865);
and U4031 (N_4031,N_3950,N_3821);
nand U4032 (N_4032,N_3887,N_3930);
nor U4033 (N_4033,N_3978,N_3806);
nor U4034 (N_4034,N_3957,N_3959);
and U4035 (N_4035,N_3929,N_3818);
and U4036 (N_4036,N_3852,N_3987);
nor U4037 (N_4037,N_3900,N_3847);
or U4038 (N_4038,N_3965,N_3984);
or U4039 (N_4039,N_3875,N_3829);
or U4040 (N_4040,N_3937,N_3981);
nand U4041 (N_4041,N_3934,N_3886);
nand U4042 (N_4042,N_3846,N_3923);
xor U4043 (N_4043,N_3893,N_3826);
nand U4044 (N_4044,N_3996,N_3837);
nor U4045 (N_4045,N_3840,N_3890);
nand U4046 (N_4046,N_3919,N_3807);
or U4047 (N_4047,N_3944,N_3905);
nand U4048 (N_4048,N_3932,N_3802);
nand U4049 (N_4049,N_3891,N_3915);
nor U4050 (N_4050,N_3882,N_3956);
xor U4051 (N_4051,N_3908,N_3872);
nor U4052 (N_4052,N_3867,N_3941);
or U4053 (N_4053,N_3848,N_3985);
nor U4054 (N_4054,N_3849,N_3946);
and U4055 (N_4055,N_3927,N_3831);
nand U4056 (N_4056,N_3903,N_3862);
xor U4057 (N_4057,N_3830,N_3855);
nand U4058 (N_4058,N_3975,N_3870);
or U4059 (N_4059,N_3971,N_3976);
and U4060 (N_4060,N_3994,N_3857);
nand U4061 (N_4061,N_3894,N_3922);
nand U4062 (N_4062,N_3910,N_3902);
nand U4063 (N_4063,N_3961,N_3851);
or U4064 (N_4064,N_3885,N_3970);
nor U4065 (N_4065,N_3871,N_3881);
or U4066 (N_4066,N_3945,N_3819);
nand U4067 (N_4067,N_3825,N_3853);
nor U4068 (N_4068,N_3982,N_3977);
nand U4069 (N_4069,N_3822,N_3928);
and U4070 (N_4070,N_3805,N_3876);
and U4071 (N_4071,N_3863,N_3963);
and U4072 (N_4072,N_3955,N_3916);
or U4073 (N_4073,N_3906,N_3992);
and U4074 (N_4074,N_3864,N_3858);
and U4075 (N_4075,N_3889,N_3926);
nor U4076 (N_4076,N_3800,N_3815);
nor U4077 (N_4077,N_3823,N_3841);
nor U4078 (N_4078,N_3836,N_3968);
nand U4079 (N_4079,N_3921,N_3861);
and U4080 (N_4080,N_3925,N_3811);
xor U4081 (N_4081,N_3839,N_3880);
or U4082 (N_4082,N_3991,N_3897);
and U4083 (N_4083,N_3901,N_3812);
or U4084 (N_4084,N_3909,N_3892);
and U4085 (N_4085,N_3943,N_3966);
or U4086 (N_4086,N_3828,N_3954);
nor U4087 (N_4087,N_3913,N_3912);
nor U4088 (N_4088,N_3835,N_3917);
xnor U4089 (N_4089,N_3878,N_3953);
or U4090 (N_4090,N_3947,N_3810);
or U4091 (N_4091,N_3951,N_3838);
nand U4092 (N_4092,N_3809,N_3904);
xor U4093 (N_4093,N_3817,N_3931);
and U4094 (N_4094,N_3939,N_3924);
nand U4095 (N_4095,N_3983,N_3995);
and U4096 (N_4096,N_3918,N_3854);
or U4097 (N_4097,N_3879,N_3833);
nand U4098 (N_4098,N_3895,N_3998);
and U4099 (N_4099,N_3834,N_3989);
nand U4100 (N_4100,N_3953,N_3927);
or U4101 (N_4101,N_3928,N_3901);
or U4102 (N_4102,N_3805,N_3926);
and U4103 (N_4103,N_3978,N_3950);
xor U4104 (N_4104,N_3960,N_3840);
nand U4105 (N_4105,N_3887,N_3820);
xnor U4106 (N_4106,N_3871,N_3813);
nand U4107 (N_4107,N_3963,N_3899);
or U4108 (N_4108,N_3830,N_3833);
and U4109 (N_4109,N_3979,N_3953);
xor U4110 (N_4110,N_3908,N_3976);
xnor U4111 (N_4111,N_3929,N_3991);
and U4112 (N_4112,N_3827,N_3887);
xnor U4113 (N_4113,N_3842,N_3936);
nor U4114 (N_4114,N_3831,N_3952);
and U4115 (N_4115,N_3968,N_3933);
nand U4116 (N_4116,N_3972,N_3982);
nor U4117 (N_4117,N_3848,N_3879);
or U4118 (N_4118,N_3842,N_3809);
xor U4119 (N_4119,N_3954,N_3980);
nand U4120 (N_4120,N_3956,N_3896);
nand U4121 (N_4121,N_3874,N_3926);
nor U4122 (N_4122,N_3891,N_3926);
or U4123 (N_4123,N_3949,N_3884);
or U4124 (N_4124,N_3914,N_3862);
and U4125 (N_4125,N_3811,N_3888);
and U4126 (N_4126,N_3886,N_3856);
nand U4127 (N_4127,N_3845,N_3851);
nor U4128 (N_4128,N_3947,N_3848);
xnor U4129 (N_4129,N_3966,N_3821);
nand U4130 (N_4130,N_3861,N_3833);
nand U4131 (N_4131,N_3807,N_3812);
nand U4132 (N_4132,N_3922,N_3854);
and U4133 (N_4133,N_3894,N_3858);
or U4134 (N_4134,N_3814,N_3826);
nand U4135 (N_4135,N_3879,N_3983);
xnor U4136 (N_4136,N_3917,N_3850);
and U4137 (N_4137,N_3999,N_3909);
nor U4138 (N_4138,N_3873,N_3801);
and U4139 (N_4139,N_3923,N_3864);
nor U4140 (N_4140,N_3956,N_3999);
nor U4141 (N_4141,N_3948,N_3847);
nor U4142 (N_4142,N_3999,N_3805);
and U4143 (N_4143,N_3952,N_3911);
nor U4144 (N_4144,N_3989,N_3911);
nor U4145 (N_4145,N_3968,N_3907);
and U4146 (N_4146,N_3949,N_3864);
or U4147 (N_4147,N_3997,N_3805);
and U4148 (N_4148,N_3935,N_3991);
and U4149 (N_4149,N_3997,N_3942);
xnor U4150 (N_4150,N_3885,N_3822);
nor U4151 (N_4151,N_3929,N_3943);
nand U4152 (N_4152,N_3858,N_3866);
nand U4153 (N_4153,N_3972,N_3989);
nand U4154 (N_4154,N_3805,N_3824);
or U4155 (N_4155,N_3851,N_3951);
and U4156 (N_4156,N_3857,N_3833);
nand U4157 (N_4157,N_3826,N_3969);
or U4158 (N_4158,N_3807,N_3986);
and U4159 (N_4159,N_3814,N_3980);
or U4160 (N_4160,N_3981,N_3946);
xnor U4161 (N_4161,N_3933,N_3929);
nor U4162 (N_4162,N_3981,N_3958);
and U4163 (N_4163,N_3862,N_3904);
nor U4164 (N_4164,N_3898,N_3977);
nand U4165 (N_4165,N_3846,N_3871);
or U4166 (N_4166,N_3807,N_3956);
and U4167 (N_4167,N_3900,N_3970);
nand U4168 (N_4168,N_3959,N_3913);
xor U4169 (N_4169,N_3968,N_3848);
nand U4170 (N_4170,N_3989,N_3967);
and U4171 (N_4171,N_3970,N_3867);
nor U4172 (N_4172,N_3955,N_3963);
nor U4173 (N_4173,N_3957,N_3912);
and U4174 (N_4174,N_3966,N_3814);
xor U4175 (N_4175,N_3889,N_3957);
nor U4176 (N_4176,N_3897,N_3852);
nand U4177 (N_4177,N_3959,N_3879);
nor U4178 (N_4178,N_3844,N_3890);
and U4179 (N_4179,N_3832,N_3802);
nor U4180 (N_4180,N_3952,N_3907);
and U4181 (N_4181,N_3861,N_3807);
nor U4182 (N_4182,N_3982,N_3826);
nor U4183 (N_4183,N_3937,N_3814);
xor U4184 (N_4184,N_3964,N_3863);
and U4185 (N_4185,N_3849,N_3817);
nor U4186 (N_4186,N_3819,N_3807);
xor U4187 (N_4187,N_3960,N_3861);
nand U4188 (N_4188,N_3840,N_3891);
nor U4189 (N_4189,N_3865,N_3873);
nor U4190 (N_4190,N_3823,N_3897);
nor U4191 (N_4191,N_3934,N_3835);
nor U4192 (N_4192,N_3890,N_3984);
nand U4193 (N_4193,N_3909,N_3837);
xnor U4194 (N_4194,N_3915,N_3918);
and U4195 (N_4195,N_3934,N_3906);
nand U4196 (N_4196,N_3882,N_3821);
nor U4197 (N_4197,N_3818,N_3826);
or U4198 (N_4198,N_3888,N_3823);
or U4199 (N_4199,N_3976,N_3831);
nand U4200 (N_4200,N_4042,N_4054);
and U4201 (N_4201,N_4085,N_4153);
nor U4202 (N_4202,N_4155,N_4121);
or U4203 (N_4203,N_4120,N_4142);
and U4204 (N_4204,N_4196,N_4029);
and U4205 (N_4205,N_4049,N_4079);
nand U4206 (N_4206,N_4187,N_4081);
and U4207 (N_4207,N_4044,N_4098);
or U4208 (N_4208,N_4119,N_4144);
nand U4209 (N_4209,N_4037,N_4138);
nor U4210 (N_4210,N_4050,N_4104);
or U4211 (N_4211,N_4078,N_4161);
nor U4212 (N_4212,N_4043,N_4130);
nand U4213 (N_4213,N_4176,N_4168);
nor U4214 (N_4214,N_4139,N_4034);
nor U4215 (N_4215,N_4084,N_4177);
xnor U4216 (N_4216,N_4183,N_4158);
xor U4217 (N_4217,N_4106,N_4072);
or U4218 (N_4218,N_4184,N_4173);
nand U4219 (N_4219,N_4093,N_4113);
nor U4220 (N_4220,N_4094,N_4015);
or U4221 (N_4221,N_4148,N_4008);
or U4222 (N_4222,N_4194,N_4033);
nor U4223 (N_4223,N_4115,N_4165);
and U4224 (N_4224,N_4135,N_4164);
and U4225 (N_4225,N_4040,N_4007);
or U4226 (N_4226,N_4112,N_4102);
nand U4227 (N_4227,N_4059,N_4020);
nor U4228 (N_4228,N_4140,N_4082);
nor U4229 (N_4229,N_4002,N_4065);
nand U4230 (N_4230,N_4109,N_4103);
and U4231 (N_4231,N_4068,N_4038);
nand U4232 (N_4232,N_4096,N_4005);
nand U4233 (N_4233,N_4089,N_4001);
xnor U4234 (N_4234,N_4060,N_4167);
and U4235 (N_4235,N_4157,N_4048);
and U4236 (N_4236,N_4051,N_4107);
nand U4237 (N_4237,N_4190,N_4191);
and U4238 (N_4238,N_4199,N_4136);
nor U4239 (N_4239,N_4198,N_4179);
or U4240 (N_4240,N_4129,N_4035);
nor U4241 (N_4241,N_4133,N_4118);
nor U4242 (N_4242,N_4122,N_4087);
and U4243 (N_4243,N_4083,N_4003);
nor U4244 (N_4244,N_4021,N_4066);
nand U4245 (N_4245,N_4032,N_4117);
or U4246 (N_4246,N_4195,N_4058);
and U4247 (N_4247,N_4057,N_4132);
or U4248 (N_4248,N_4010,N_4025);
and U4249 (N_4249,N_4017,N_4143);
nand U4250 (N_4250,N_4101,N_4030);
and U4251 (N_4251,N_4116,N_4163);
or U4252 (N_4252,N_4067,N_4174);
and U4253 (N_4253,N_4039,N_4162);
xor U4254 (N_4254,N_4110,N_4075);
and U4255 (N_4255,N_4031,N_4080);
and U4256 (N_4256,N_4124,N_4172);
and U4257 (N_4257,N_4063,N_4146);
or U4258 (N_4258,N_4105,N_4011);
nor U4259 (N_4259,N_4097,N_4013);
or U4260 (N_4260,N_4006,N_4024);
nand U4261 (N_4261,N_4070,N_4071);
and U4262 (N_4262,N_4149,N_4123);
nand U4263 (N_4263,N_4047,N_4018);
and U4264 (N_4264,N_4086,N_4150);
xnor U4265 (N_4265,N_4088,N_4036);
or U4266 (N_4266,N_4053,N_4188);
xnor U4267 (N_4267,N_4182,N_4052);
nor U4268 (N_4268,N_4197,N_4016);
nor U4269 (N_4269,N_4009,N_4091);
xor U4270 (N_4270,N_4026,N_4126);
and U4271 (N_4271,N_4077,N_4152);
and U4272 (N_4272,N_4064,N_4014);
nor U4273 (N_4273,N_4099,N_4108);
and U4274 (N_4274,N_4074,N_4095);
nand U4275 (N_4275,N_4137,N_4181);
or U4276 (N_4276,N_4169,N_4022);
nand U4277 (N_4277,N_4127,N_4073);
nor U4278 (N_4278,N_4004,N_4125);
nor U4279 (N_4279,N_4178,N_4069);
and U4280 (N_4280,N_4090,N_4154);
xor U4281 (N_4281,N_4000,N_4111);
nor U4282 (N_4282,N_4185,N_4056);
or U4283 (N_4283,N_4145,N_4027);
xnor U4284 (N_4284,N_4147,N_4046);
or U4285 (N_4285,N_4114,N_4166);
and U4286 (N_4286,N_4160,N_4141);
or U4287 (N_4287,N_4159,N_4041);
xnor U4288 (N_4288,N_4156,N_4076);
xnor U4289 (N_4289,N_4175,N_4012);
xnor U4290 (N_4290,N_4100,N_4092);
and U4291 (N_4291,N_4131,N_4180);
nor U4292 (N_4292,N_4055,N_4019);
and U4293 (N_4293,N_4128,N_4186);
nand U4294 (N_4294,N_4193,N_4170);
and U4295 (N_4295,N_4061,N_4171);
nand U4296 (N_4296,N_4192,N_4151);
or U4297 (N_4297,N_4189,N_4028);
nor U4298 (N_4298,N_4062,N_4045);
nor U4299 (N_4299,N_4023,N_4134);
nand U4300 (N_4300,N_4030,N_4173);
xor U4301 (N_4301,N_4188,N_4158);
and U4302 (N_4302,N_4110,N_4109);
or U4303 (N_4303,N_4174,N_4068);
nand U4304 (N_4304,N_4091,N_4130);
nor U4305 (N_4305,N_4074,N_4005);
nand U4306 (N_4306,N_4133,N_4181);
and U4307 (N_4307,N_4145,N_4085);
and U4308 (N_4308,N_4055,N_4013);
and U4309 (N_4309,N_4003,N_4182);
nor U4310 (N_4310,N_4159,N_4162);
and U4311 (N_4311,N_4178,N_4129);
nand U4312 (N_4312,N_4067,N_4173);
nand U4313 (N_4313,N_4191,N_4133);
and U4314 (N_4314,N_4048,N_4103);
and U4315 (N_4315,N_4028,N_4029);
and U4316 (N_4316,N_4142,N_4007);
xnor U4317 (N_4317,N_4002,N_4032);
nand U4318 (N_4318,N_4013,N_4028);
xor U4319 (N_4319,N_4165,N_4011);
nand U4320 (N_4320,N_4081,N_4152);
or U4321 (N_4321,N_4004,N_4182);
nand U4322 (N_4322,N_4012,N_4095);
and U4323 (N_4323,N_4177,N_4137);
nor U4324 (N_4324,N_4095,N_4130);
or U4325 (N_4325,N_4155,N_4165);
xor U4326 (N_4326,N_4158,N_4190);
nand U4327 (N_4327,N_4125,N_4183);
xor U4328 (N_4328,N_4165,N_4150);
or U4329 (N_4329,N_4146,N_4118);
nand U4330 (N_4330,N_4176,N_4117);
nor U4331 (N_4331,N_4041,N_4088);
or U4332 (N_4332,N_4059,N_4084);
and U4333 (N_4333,N_4193,N_4052);
or U4334 (N_4334,N_4090,N_4006);
or U4335 (N_4335,N_4163,N_4082);
and U4336 (N_4336,N_4165,N_4013);
and U4337 (N_4337,N_4083,N_4098);
and U4338 (N_4338,N_4025,N_4106);
nor U4339 (N_4339,N_4152,N_4160);
nor U4340 (N_4340,N_4169,N_4013);
or U4341 (N_4341,N_4074,N_4097);
and U4342 (N_4342,N_4153,N_4011);
nor U4343 (N_4343,N_4168,N_4082);
xnor U4344 (N_4344,N_4066,N_4109);
nor U4345 (N_4345,N_4070,N_4042);
xor U4346 (N_4346,N_4170,N_4144);
and U4347 (N_4347,N_4108,N_4195);
and U4348 (N_4348,N_4082,N_4109);
nor U4349 (N_4349,N_4187,N_4154);
and U4350 (N_4350,N_4097,N_4179);
nor U4351 (N_4351,N_4138,N_4041);
nor U4352 (N_4352,N_4141,N_4185);
nand U4353 (N_4353,N_4115,N_4136);
nand U4354 (N_4354,N_4098,N_4139);
and U4355 (N_4355,N_4189,N_4094);
and U4356 (N_4356,N_4133,N_4079);
nand U4357 (N_4357,N_4036,N_4102);
nand U4358 (N_4358,N_4131,N_4030);
or U4359 (N_4359,N_4084,N_4186);
nand U4360 (N_4360,N_4003,N_4032);
and U4361 (N_4361,N_4091,N_4065);
nand U4362 (N_4362,N_4144,N_4084);
nor U4363 (N_4363,N_4075,N_4037);
and U4364 (N_4364,N_4100,N_4071);
or U4365 (N_4365,N_4023,N_4053);
nor U4366 (N_4366,N_4027,N_4160);
nor U4367 (N_4367,N_4053,N_4132);
and U4368 (N_4368,N_4100,N_4020);
or U4369 (N_4369,N_4034,N_4197);
nor U4370 (N_4370,N_4117,N_4072);
or U4371 (N_4371,N_4040,N_4016);
nand U4372 (N_4372,N_4199,N_4077);
and U4373 (N_4373,N_4102,N_4107);
nor U4374 (N_4374,N_4145,N_4047);
or U4375 (N_4375,N_4154,N_4069);
or U4376 (N_4376,N_4028,N_4081);
nor U4377 (N_4377,N_4167,N_4156);
and U4378 (N_4378,N_4113,N_4108);
xor U4379 (N_4379,N_4124,N_4199);
and U4380 (N_4380,N_4123,N_4168);
nand U4381 (N_4381,N_4069,N_4169);
nand U4382 (N_4382,N_4087,N_4018);
nand U4383 (N_4383,N_4044,N_4108);
nor U4384 (N_4384,N_4047,N_4127);
and U4385 (N_4385,N_4133,N_4051);
and U4386 (N_4386,N_4029,N_4156);
or U4387 (N_4387,N_4130,N_4070);
nor U4388 (N_4388,N_4162,N_4030);
nand U4389 (N_4389,N_4028,N_4057);
xor U4390 (N_4390,N_4140,N_4056);
nand U4391 (N_4391,N_4123,N_4050);
nor U4392 (N_4392,N_4145,N_4174);
nor U4393 (N_4393,N_4031,N_4166);
or U4394 (N_4394,N_4178,N_4158);
nor U4395 (N_4395,N_4162,N_4190);
and U4396 (N_4396,N_4113,N_4132);
or U4397 (N_4397,N_4187,N_4160);
nand U4398 (N_4398,N_4117,N_4115);
nor U4399 (N_4399,N_4081,N_4109);
and U4400 (N_4400,N_4332,N_4319);
or U4401 (N_4401,N_4300,N_4366);
or U4402 (N_4402,N_4227,N_4271);
or U4403 (N_4403,N_4243,N_4387);
or U4404 (N_4404,N_4369,N_4344);
nand U4405 (N_4405,N_4209,N_4298);
and U4406 (N_4406,N_4303,N_4235);
xnor U4407 (N_4407,N_4275,N_4311);
nand U4408 (N_4408,N_4281,N_4256);
xor U4409 (N_4409,N_4381,N_4232);
or U4410 (N_4410,N_4318,N_4384);
nand U4411 (N_4411,N_4399,N_4390);
nand U4412 (N_4412,N_4345,N_4295);
nor U4413 (N_4413,N_4324,N_4376);
and U4414 (N_4414,N_4291,N_4219);
nor U4415 (N_4415,N_4252,N_4350);
nor U4416 (N_4416,N_4353,N_4362);
and U4417 (N_4417,N_4225,N_4296);
xor U4418 (N_4418,N_4357,N_4211);
nor U4419 (N_4419,N_4320,N_4321);
nand U4420 (N_4420,N_4356,N_4282);
xnor U4421 (N_4421,N_4379,N_4327);
nor U4422 (N_4422,N_4386,N_4280);
and U4423 (N_4423,N_4268,N_4391);
xor U4424 (N_4424,N_4279,N_4367);
nand U4425 (N_4425,N_4349,N_4338);
and U4426 (N_4426,N_4316,N_4218);
nand U4427 (N_4427,N_4383,N_4337);
nor U4428 (N_4428,N_4330,N_4237);
and U4429 (N_4429,N_4221,N_4329);
nand U4430 (N_4430,N_4299,N_4297);
or U4431 (N_4431,N_4359,N_4393);
nor U4432 (N_4432,N_4361,N_4250);
and U4433 (N_4433,N_4322,N_4308);
nand U4434 (N_4434,N_4200,N_4233);
and U4435 (N_4435,N_4348,N_4231);
nor U4436 (N_4436,N_4377,N_4292);
and U4437 (N_4437,N_4201,N_4333);
nor U4438 (N_4438,N_4389,N_4278);
or U4439 (N_4439,N_4210,N_4396);
nand U4440 (N_4440,N_4395,N_4392);
or U4441 (N_4441,N_4334,N_4304);
nor U4442 (N_4442,N_4241,N_4336);
or U4443 (N_4443,N_4205,N_4286);
xor U4444 (N_4444,N_4302,N_4240);
xor U4445 (N_4445,N_4347,N_4251);
and U4446 (N_4446,N_4289,N_4223);
nand U4447 (N_4447,N_4394,N_4364);
nand U4448 (N_4448,N_4264,N_4380);
or U4449 (N_4449,N_4236,N_4203);
and U4450 (N_4450,N_4288,N_4375);
or U4451 (N_4451,N_4239,N_4371);
and U4452 (N_4452,N_4212,N_4208);
xor U4453 (N_4453,N_4254,N_4242);
or U4454 (N_4454,N_4217,N_4317);
and U4455 (N_4455,N_4257,N_4307);
nand U4456 (N_4456,N_4397,N_4269);
nor U4457 (N_4457,N_4249,N_4352);
and U4458 (N_4458,N_4226,N_4368);
or U4459 (N_4459,N_4312,N_4259);
and U4460 (N_4460,N_4293,N_4373);
and U4461 (N_4461,N_4370,N_4234);
and U4462 (N_4462,N_4363,N_4262);
nor U4463 (N_4463,N_4255,N_4283);
nand U4464 (N_4464,N_4342,N_4216);
nand U4465 (N_4465,N_4305,N_4314);
nand U4466 (N_4466,N_4253,N_4340);
nand U4467 (N_4467,N_4374,N_4244);
and U4468 (N_4468,N_4267,N_4224);
or U4469 (N_4469,N_4382,N_4310);
xnor U4470 (N_4470,N_4220,N_4246);
nor U4471 (N_4471,N_4358,N_4346);
nor U4472 (N_4472,N_4277,N_4365);
nand U4473 (N_4473,N_4360,N_4229);
nor U4474 (N_4474,N_4215,N_4372);
nand U4475 (N_4475,N_4323,N_4294);
nand U4476 (N_4476,N_4287,N_4385);
nor U4477 (N_4477,N_4228,N_4284);
nor U4478 (N_4478,N_4309,N_4331);
or U4479 (N_4479,N_4315,N_4258);
nor U4480 (N_4480,N_4325,N_4354);
or U4481 (N_4481,N_4339,N_4214);
and U4482 (N_4482,N_4274,N_4230);
nand U4483 (N_4483,N_4355,N_4273);
or U4484 (N_4484,N_4335,N_4328);
nor U4485 (N_4485,N_4266,N_4341);
or U4486 (N_4486,N_4261,N_4247);
nor U4487 (N_4487,N_4301,N_4204);
and U4488 (N_4488,N_4206,N_4388);
nand U4489 (N_4489,N_4222,N_4285);
or U4490 (N_4490,N_4245,N_4248);
nand U4491 (N_4491,N_4313,N_4306);
nor U4492 (N_4492,N_4270,N_4213);
nor U4493 (N_4493,N_4238,N_4378);
and U4494 (N_4494,N_4263,N_4265);
xor U4495 (N_4495,N_4272,N_4398);
nand U4496 (N_4496,N_4260,N_4351);
nand U4497 (N_4497,N_4276,N_4290);
xnor U4498 (N_4498,N_4326,N_4202);
or U4499 (N_4499,N_4343,N_4207);
nor U4500 (N_4500,N_4236,N_4256);
nor U4501 (N_4501,N_4394,N_4322);
nor U4502 (N_4502,N_4233,N_4314);
and U4503 (N_4503,N_4326,N_4329);
nand U4504 (N_4504,N_4360,N_4252);
or U4505 (N_4505,N_4376,N_4237);
and U4506 (N_4506,N_4377,N_4290);
and U4507 (N_4507,N_4216,N_4238);
and U4508 (N_4508,N_4288,N_4294);
nor U4509 (N_4509,N_4237,N_4245);
or U4510 (N_4510,N_4309,N_4249);
nand U4511 (N_4511,N_4283,N_4226);
nand U4512 (N_4512,N_4211,N_4261);
and U4513 (N_4513,N_4276,N_4231);
nand U4514 (N_4514,N_4347,N_4260);
or U4515 (N_4515,N_4249,N_4363);
and U4516 (N_4516,N_4236,N_4356);
and U4517 (N_4517,N_4388,N_4263);
xor U4518 (N_4518,N_4364,N_4363);
nor U4519 (N_4519,N_4353,N_4231);
or U4520 (N_4520,N_4239,N_4222);
nor U4521 (N_4521,N_4332,N_4267);
or U4522 (N_4522,N_4393,N_4306);
nand U4523 (N_4523,N_4334,N_4344);
or U4524 (N_4524,N_4250,N_4233);
nor U4525 (N_4525,N_4368,N_4374);
nor U4526 (N_4526,N_4367,N_4221);
or U4527 (N_4527,N_4269,N_4380);
or U4528 (N_4528,N_4209,N_4315);
and U4529 (N_4529,N_4336,N_4389);
nor U4530 (N_4530,N_4295,N_4341);
nor U4531 (N_4531,N_4329,N_4365);
or U4532 (N_4532,N_4248,N_4380);
nand U4533 (N_4533,N_4305,N_4306);
and U4534 (N_4534,N_4364,N_4358);
or U4535 (N_4535,N_4279,N_4253);
nor U4536 (N_4536,N_4211,N_4244);
nor U4537 (N_4537,N_4293,N_4290);
nor U4538 (N_4538,N_4358,N_4202);
xor U4539 (N_4539,N_4269,N_4317);
nand U4540 (N_4540,N_4246,N_4224);
and U4541 (N_4541,N_4226,N_4250);
nor U4542 (N_4542,N_4334,N_4325);
or U4543 (N_4543,N_4391,N_4205);
nor U4544 (N_4544,N_4398,N_4362);
or U4545 (N_4545,N_4201,N_4216);
or U4546 (N_4546,N_4304,N_4347);
nor U4547 (N_4547,N_4286,N_4375);
nor U4548 (N_4548,N_4200,N_4293);
nand U4549 (N_4549,N_4372,N_4290);
nor U4550 (N_4550,N_4206,N_4274);
and U4551 (N_4551,N_4305,N_4276);
xnor U4552 (N_4552,N_4331,N_4203);
and U4553 (N_4553,N_4209,N_4226);
and U4554 (N_4554,N_4308,N_4247);
xor U4555 (N_4555,N_4245,N_4299);
and U4556 (N_4556,N_4391,N_4349);
nor U4557 (N_4557,N_4228,N_4267);
nand U4558 (N_4558,N_4218,N_4265);
nor U4559 (N_4559,N_4256,N_4289);
xnor U4560 (N_4560,N_4283,N_4281);
nor U4561 (N_4561,N_4292,N_4254);
and U4562 (N_4562,N_4203,N_4287);
and U4563 (N_4563,N_4358,N_4333);
xor U4564 (N_4564,N_4204,N_4395);
xor U4565 (N_4565,N_4316,N_4389);
and U4566 (N_4566,N_4387,N_4246);
and U4567 (N_4567,N_4371,N_4225);
or U4568 (N_4568,N_4393,N_4380);
nor U4569 (N_4569,N_4383,N_4288);
nand U4570 (N_4570,N_4311,N_4323);
and U4571 (N_4571,N_4258,N_4314);
and U4572 (N_4572,N_4398,N_4379);
nand U4573 (N_4573,N_4287,N_4217);
or U4574 (N_4574,N_4375,N_4210);
and U4575 (N_4575,N_4206,N_4336);
and U4576 (N_4576,N_4235,N_4286);
and U4577 (N_4577,N_4251,N_4241);
and U4578 (N_4578,N_4225,N_4367);
or U4579 (N_4579,N_4288,N_4317);
nor U4580 (N_4580,N_4304,N_4278);
nand U4581 (N_4581,N_4277,N_4220);
nand U4582 (N_4582,N_4391,N_4329);
xnor U4583 (N_4583,N_4283,N_4227);
nand U4584 (N_4584,N_4202,N_4255);
or U4585 (N_4585,N_4311,N_4308);
nor U4586 (N_4586,N_4314,N_4241);
nand U4587 (N_4587,N_4295,N_4386);
nor U4588 (N_4588,N_4218,N_4345);
or U4589 (N_4589,N_4343,N_4275);
or U4590 (N_4590,N_4211,N_4225);
or U4591 (N_4591,N_4206,N_4282);
or U4592 (N_4592,N_4302,N_4270);
or U4593 (N_4593,N_4328,N_4387);
or U4594 (N_4594,N_4352,N_4393);
xor U4595 (N_4595,N_4333,N_4310);
nor U4596 (N_4596,N_4231,N_4385);
nand U4597 (N_4597,N_4243,N_4283);
nand U4598 (N_4598,N_4343,N_4293);
and U4599 (N_4599,N_4343,N_4344);
or U4600 (N_4600,N_4456,N_4445);
or U4601 (N_4601,N_4435,N_4590);
nand U4602 (N_4602,N_4457,N_4436);
nand U4603 (N_4603,N_4474,N_4587);
nor U4604 (N_4604,N_4454,N_4552);
and U4605 (N_4605,N_4538,N_4579);
xor U4606 (N_4606,N_4488,N_4517);
and U4607 (N_4607,N_4532,N_4508);
or U4608 (N_4608,N_4547,N_4401);
xnor U4609 (N_4609,N_4495,N_4582);
nor U4610 (N_4610,N_4470,N_4430);
and U4611 (N_4611,N_4599,N_4505);
and U4612 (N_4612,N_4402,N_4419);
or U4613 (N_4613,N_4493,N_4576);
xnor U4614 (N_4614,N_4574,N_4528);
nor U4615 (N_4615,N_4417,N_4506);
or U4616 (N_4616,N_4423,N_4524);
or U4617 (N_4617,N_4521,N_4404);
xnor U4618 (N_4618,N_4561,N_4461);
nor U4619 (N_4619,N_4565,N_4463);
or U4620 (N_4620,N_4472,N_4554);
nand U4621 (N_4621,N_4406,N_4441);
nor U4622 (N_4622,N_4422,N_4555);
and U4623 (N_4623,N_4514,N_4492);
nand U4624 (N_4624,N_4400,N_4433);
or U4625 (N_4625,N_4567,N_4455);
nand U4626 (N_4626,N_4462,N_4497);
nor U4627 (N_4627,N_4546,N_4413);
and U4628 (N_4628,N_4491,N_4450);
nor U4629 (N_4629,N_4515,N_4519);
nor U4630 (N_4630,N_4551,N_4414);
or U4631 (N_4631,N_4584,N_4504);
and U4632 (N_4632,N_4586,N_4486);
xor U4633 (N_4633,N_4481,N_4478);
nor U4634 (N_4634,N_4544,N_4484);
xnor U4635 (N_4635,N_4416,N_4578);
nand U4636 (N_4636,N_4442,N_4467);
xnor U4637 (N_4637,N_4466,N_4432);
xnor U4638 (N_4638,N_4437,N_4499);
nand U4639 (N_4639,N_4440,N_4564);
or U4640 (N_4640,N_4523,N_4500);
and U4641 (N_4641,N_4409,N_4421);
or U4642 (N_4642,N_4558,N_4447);
xnor U4643 (N_4643,N_4560,N_4411);
or U4644 (N_4644,N_4420,N_4591);
nor U4645 (N_4645,N_4516,N_4460);
nand U4646 (N_4646,N_4526,N_4498);
and U4647 (N_4647,N_4448,N_4476);
and U4648 (N_4648,N_4425,N_4465);
xnor U4649 (N_4649,N_4477,N_4464);
nor U4650 (N_4650,N_4503,N_4525);
nand U4651 (N_4651,N_4535,N_4443);
xnor U4652 (N_4652,N_4533,N_4496);
nor U4653 (N_4653,N_4571,N_4512);
and U4654 (N_4654,N_4483,N_4548);
or U4655 (N_4655,N_4407,N_4408);
nor U4656 (N_4656,N_4568,N_4588);
nor U4657 (N_4657,N_4502,N_4410);
and U4658 (N_4658,N_4543,N_4540);
nand U4659 (N_4659,N_4458,N_4471);
or U4660 (N_4660,N_4592,N_4509);
and U4661 (N_4661,N_4549,N_4563);
nor U4662 (N_4662,N_4469,N_4431);
and U4663 (N_4663,N_4415,N_4513);
nor U4664 (N_4664,N_4545,N_4570);
and U4665 (N_4665,N_4553,N_4537);
or U4666 (N_4666,N_4487,N_4480);
xor U4667 (N_4667,N_4459,N_4468);
nand U4668 (N_4668,N_4427,N_4593);
or U4669 (N_4669,N_4580,N_4428);
xnor U4670 (N_4670,N_4403,N_4424);
or U4671 (N_4671,N_4583,N_4518);
and U4672 (N_4672,N_4581,N_4522);
nand U4673 (N_4673,N_4473,N_4438);
and U4674 (N_4674,N_4485,N_4482);
nand U4675 (N_4675,N_4444,N_4595);
or U4676 (N_4676,N_4534,N_4594);
nand U4677 (N_4677,N_4562,N_4575);
and U4678 (N_4678,N_4494,N_4507);
or U4679 (N_4679,N_4520,N_4446);
or U4680 (N_4680,N_4479,N_4529);
and U4681 (N_4681,N_4557,N_4434);
or U4682 (N_4682,N_4589,N_4531);
nand U4683 (N_4683,N_4451,N_4511);
and U4684 (N_4684,N_4550,N_4536);
nand U4685 (N_4685,N_4541,N_4539);
and U4686 (N_4686,N_4405,N_4542);
or U4687 (N_4687,N_4573,N_4489);
nand U4688 (N_4688,N_4596,N_4572);
nor U4689 (N_4689,N_4569,N_4585);
or U4690 (N_4690,N_4475,N_4598);
and U4691 (N_4691,N_4527,N_4577);
xnor U4692 (N_4692,N_4530,N_4418);
or U4693 (N_4693,N_4449,N_4426);
and U4694 (N_4694,N_4597,N_4453);
and U4695 (N_4695,N_4412,N_4452);
nor U4696 (N_4696,N_4501,N_4490);
and U4697 (N_4697,N_4556,N_4429);
nor U4698 (N_4698,N_4510,N_4559);
nand U4699 (N_4699,N_4566,N_4439);
xor U4700 (N_4700,N_4553,N_4428);
or U4701 (N_4701,N_4503,N_4556);
xor U4702 (N_4702,N_4558,N_4566);
nor U4703 (N_4703,N_4569,N_4494);
nand U4704 (N_4704,N_4405,N_4425);
nor U4705 (N_4705,N_4553,N_4434);
nand U4706 (N_4706,N_4412,N_4577);
nand U4707 (N_4707,N_4582,N_4517);
xnor U4708 (N_4708,N_4565,N_4525);
and U4709 (N_4709,N_4538,N_4578);
or U4710 (N_4710,N_4412,N_4474);
nor U4711 (N_4711,N_4584,N_4565);
nor U4712 (N_4712,N_4536,N_4441);
and U4713 (N_4713,N_4582,N_4425);
and U4714 (N_4714,N_4427,N_4571);
or U4715 (N_4715,N_4417,N_4503);
nand U4716 (N_4716,N_4458,N_4465);
and U4717 (N_4717,N_4461,N_4437);
nand U4718 (N_4718,N_4482,N_4447);
nand U4719 (N_4719,N_4530,N_4537);
and U4720 (N_4720,N_4562,N_4514);
nor U4721 (N_4721,N_4538,N_4505);
nand U4722 (N_4722,N_4458,N_4469);
nor U4723 (N_4723,N_4466,N_4421);
nor U4724 (N_4724,N_4414,N_4435);
nand U4725 (N_4725,N_4465,N_4405);
nand U4726 (N_4726,N_4404,N_4569);
nand U4727 (N_4727,N_4406,N_4588);
nor U4728 (N_4728,N_4592,N_4434);
nor U4729 (N_4729,N_4553,N_4477);
nand U4730 (N_4730,N_4463,N_4521);
and U4731 (N_4731,N_4514,N_4571);
or U4732 (N_4732,N_4473,N_4536);
nor U4733 (N_4733,N_4504,N_4552);
or U4734 (N_4734,N_4522,N_4525);
xnor U4735 (N_4735,N_4588,N_4473);
or U4736 (N_4736,N_4472,N_4492);
and U4737 (N_4737,N_4546,N_4447);
nor U4738 (N_4738,N_4449,N_4500);
nor U4739 (N_4739,N_4578,N_4521);
nand U4740 (N_4740,N_4421,N_4547);
nor U4741 (N_4741,N_4533,N_4562);
nand U4742 (N_4742,N_4536,N_4563);
and U4743 (N_4743,N_4519,N_4416);
nor U4744 (N_4744,N_4517,N_4424);
nor U4745 (N_4745,N_4510,N_4509);
nand U4746 (N_4746,N_4571,N_4506);
nand U4747 (N_4747,N_4564,N_4565);
nand U4748 (N_4748,N_4481,N_4592);
nand U4749 (N_4749,N_4457,N_4427);
nand U4750 (N_4750,N_4488,N_4486);
and U4751 (N_4751,N_4554,N_4569);
nand U4752 (N_4752,N_4417,N_4574);
or U4753 (N_4753,N_4575,N_4594);
nor U4754 (N_4754,N_4468,N_4587);
nand U4755 (N_4755,N_4516,N_4511);
xnor U4756 (N_4756,N_4517,N_4435);
and U4757 (N_4757,N_4468,N_4467);
nand U4758 (N_4758,N_4496,N_4418);
nor U4759 (N_4759,N_4431,N_4493);
or U4760 (N_4760,N_4448,N_4420);
nor U4761 (N_4761,N_4499,N_4529);
or U4762 (N_4762,N_4452,N_4533);
or U4763 (N_4763,N_4585,N_4546);
nand U4764 (N_4764,N_4405,N_4592);
or U4765 (N_4765,N_4534,N_4406);
nand U4766 (N_4766,N_4453,N_4445);
and U4767 (N_4767,N_4588,N_4426);
nor U4768 (N_4768,N_4456,N_4517);
nand U4769 (N_4769,N_4521,N_4568);
or U4770 (N_4770,N_4574,N_4551);
nor U4771 (N_4771,N_4558,N_4572);
nand U4772 (N_4772,N_4512,N_4477);
or U4773 (N_4773,N_4490,N_4480);
nor U4774 (N_4774,N_4510,N_4408);
nand U4775 (N_4775,N_4465,N_4550);
nor U4776 (N_4776,N_4466,N_4506);
and U4777 (N_4777,N_4438,N_4546);
nor U4778 (N_4778,N_4518,N_4532);
and U4779 (N_4779,N_4540,N_4510);
xnor U4780 (N_4780,N_4419,N_4416);
or U4781 (N_4781,N_4405,N_4561);
or U4782 (N_4782,N_4425,N_4406);
and U4783 (N_4783,N_4498,N_4445);
or U4784 (N_4784,N_4504,N_4446);
xor U4785 (N_4785,N_4433,N_4593);
xnor U4786 (N_4786,N_4441,N_4554);
nand U4787 (N_4787,N_4520,N_4539);
nand U4788 (N_4788,N_4461,N_4502);
nor U4789 (N_4789,N_4474,N_4588);
nor U4790 (N_4790,N_4471,N_4582);
and U4791 (N_4791,N_4547,N_4414);
nor U4792 (N_4792,N_4530,N_4519);
nand U4793 (N_4793,N_4453,N_4499);
and U4794 (N_4794,N_4463,N_4580);
or U4795 (N_4795,N_4467,N_4482);
and U4796 (N_4796,N_4402,N_4552);
or U4797 (N_4797,N_4407,N_4564);
xnor U4798 (N_4798,N_4564,N_4457);
nor U4799 (N_4799,N_4558,N_4481);
nand U4800 (N_4800,N_4752,N_4749);
or U4801 (N_4801,N_4706,N_4753);
nand U4802 (N_4802,N_4790,N_4628);
or U4803 (N_4803,N_4642,N_4604);
and U4804 (N_4804,N_4646,N_4781);
nor U4805 (N_4805,N_4797,N_4673);
nor U4806 (N_4806,N_4782,N_4788);
nand U4807 (N_4807,N_4674,N_4689);
nand U4808 (N_4808,N_4666,N_4671);
nand U4809 (N_4809,N_4763,N_4651);
or U4810 (N_4810,N_4791,N_4668);
xnor U4811 (N_4811,N_4669,N_4698);
or U4812 (N_4812,N_4631,N_4718);
nand U4813 (N_4813,N_4794,N_4638);
and U4814 (N_4814,N_4769,N_4758);
nand U4815 (N_4815,N_4768,N_4739);
or U4816 (N_4816,N_4741,N_4732);
nor U4817 (N_4817,N_4636,N_4771);
nand U4818 (N_4818,N_4784,N_4606);
nand U4819 (N_4819,N_4662,N_4657);
or U4820 (N_4820,N_4745,N_4640);
or U4821 (N_4821,N_4600,N_4616);
nor U4822 (N_4822,N_4792,N_4759);
and U4823 (N_4823,N_4711,N_4775);
nor U4824 (N_4824,N_4730,N_4619);
and U4825 (N_4825,N_4729,N_4766);
or U4826 (N_4826,N_4654,N_4650);
nor U4827 (N_4827,N_4658,N_4716);
or U4828 (N_4828,N_4723,N_4786);
and U4829 (N_4829,N_4678,N_4704);
nand U4830 (N_4830,N_4693,N_4760);
nor U4831 (N_4831,N_4612,N_4725);
nand U4832 (N_4832,N_4655,N_4762);
nand U4833 (N_4833,N_4682,N_4634);
nor U4834 (N_4834,N_4765,N_4726);
or U4835 (N_4835,N_4694,N_4737);
nor U4836 (N_4836,N_4691,N_4705);
nand U4837 (N_4837,N_4780,N_4796);
nand U4838 (N_4838,N_4617,N_4773);
and U4839 (N_4839,N_4690,N_4747);
nand U4840 (N_4840,N_4667,N_4736);
or U4841 (N_4841,N_4607,N_4755);
nand U4842 (N_4842,N_4707,N_4754);
or U4843 (N_4843,N_4779,N_4645);
nand U4844 (N_4844,N_4630,N_4605);
nand U4845 (N_4845,N_4717,N_4675);
nor U4846 (N_4846,N_4710,N_4601);
and U4847 (N_4847,N_4770,N_4602);
nor U4848 (N_4848,N_4728,N_4799);
xnor U4849 (N_4849,N_4621,N_4798);
or U4850 (N_4850,N_4660,N_4714);
nand U4851 (N_4851,N_4701,N_4618);
and U4852 (N_4852,N_4664,N_4695);
and U4853 (N_4853,N_4686,N_4738);
and U4854 (N_4854,N_4778,N_4708);
nand U4855 (N_4855,N_4720,N_4697);
nand U4856 (N_4856,N_4641,N_4683);
nor U4857 (N_4857,N_4614,N_4672);
or U4858 (N_4858,N_4623,N_4685);
nor U4859 (N_4859,N_4647,N_4665);
or U4860 (N_4860,N_4699,N_4610);
nand U4861 (N_4861,N_4632,N_4635);
or U4862 (N_4862,N_4746,N_4743);
xor U4863 (N_4863,N_4777,N_4783);
and U4864 (N_4864,N_4733,N_4721);
nor U4865 (N_4865,N_4715,N_4757);
and U4866 (N_4866,N_4653,N_4724);
and U4867 (N_4867,N_4620,N_4712);
xnor U4868 (N_4868,N_4793,N_4661);
nor U4869 (N_4869,N_4625,N_4611);
or U4870 (N_4870,N_4663,N_4764);
xnor U4871 (N_4871,N_4677,N_4727);
and U4872 (N_4872,N_4615,N_4659);
xnor U4873 (N_4873,N_4622,N_4643);
nor U4874 (N_4874,N_4649,N_4751);
xnor U4875 (N_4875,N_4734,N_4735);
xor U4876 (N_4876,N_4652,N_4609);
or U4877 (N_4877,N_4722,N_4676);
nor U4878 (N_4878,N_4785,N_4772);
nor U4879 (N_4879,N_4633,N_4703);
nor U4880 (N_4880,N_4639,N_4787);
or U4881 (N_4881,N_4684,N_4627);
and U4882 (N_4882,N_4731,N_4679);
or U4883 (N_4883,N_4709,N_4608);
and U4884 (N_4884,N_4688,N_4761);
nor U4885 (N_4885,N_4648,N_4748);
or U4886 (N_4886,N_4626,N_4700);
nand U4887 (N_4887,N_4670,N_4776);
nand U4888 (N_4888,N_4702,N_4795);
and U4889 (N_4889,N_4603,N_4750);
and U4890 (N_4890,N_4692,N_4624);
nor U4891 (N_4891,N_4744,N_4644);
nand U4892 (N_4892,N_4687,N_4629);
xor U4893 (N_4893,N_4613,N_4713);
or U4894 (N_4894,N_4742,N_4740);
nand U4895 (N_4895,N_4789,N_4696);
nand U4896 (N_4896,N_4680,N_4681);
nand U4897 (N_4897,N_4719,N_4637);
nor U4898 (N_4898,N_4756,N_4656);
nor U4899 (N_4899,N_4767,N_4774);
and U4900 (N_4900,N_4789,N_4706);
nand U4901 (N_4901,N_4741,N_4641);
nor U4902 (N_4902,N_4774,N_4696);
nor U4903 (N_4903,N_4679,N_4780);
nand U4904 (N_4904,N_4673,N_4726);
nor U4905 (N_4905,N_4779,N_4675);
nor U4906 (N_4906,N_4797,N_4790);
and U4907 (N_4907,N_4798,N_4670);
or U4908 (N_4908,N_4668,N_4608);
and U4909 (N_4909,N_4763,N_4788);
nor U4910 (N_4910,N_4675,N_4615);
or U4911 (N_4911,N_4783,N_4602);
nand U4912 (N_4912,N_4722,N_4657);
or U4913 (N_4913,N_4766,N_4769);
nand U4914 (N_4914,N_4713,N_4785);
nor U4915 (N_4915,N_4686,N_4737);
nand U4916 (N_4916,N_4647,N_4609);
or U4917 (N_4917,N_4639,N_4752);
nor U4918 (N_4918,N_4715,N_4675);
nor U4919 (N_4919,N_4763,N_4690);
and U4920 (N_4920,N_4792,N_4637);
nor U4921 (N_4921,N_4678,N_4759);
nand U4922 (N_4922,N_4683,N_4781);
nand U4923 (N_4923,N_4695,N_4606);
nor U4924 (N_4924,N_4735,N_4657);
nor U4925 (N_4925,N_4656,N_4645);
or U4926 (N_4926,N_4678,N_4772);
or U4927 (N_4927,N_4652,N_4658);
nand U4928 (N_4928,N_4749,N_4720);
and U4929 (N_4929,N_4720,N_4677);
nor U4930 (N_4930,N_4774,N_4669);
nand U4931 (N_4931,N_4649,N_4605);
or U4932 (N_4932,N_4725,N_4639);
nor U4933 (N_4933,N_4632,N_4616);
or U4934 (N_4934,N_4652,N_4630);
and U4935 (N_4935,N_4755,N_4700);
or U4936 (N_4936,N_4785,N_4712);
or U4937 (N_4937,N_4667,N_4681);
nor U4938 (N_4938,N_4768,N_4656);
or U4939 (N_4939,N_4746,N_4722);
and U4940 (N_4940,N_4799,N_4761);
nor U4941 (N_4941,N_4675,N_4730);
or U4942 (N_4942,N_4786,N_4622);
xor U4943 (N_4943,N_4615,N_4782);
nand U4944 (N_4944,N_4761,N_4607);
or U4945 (N_4945,N_4664,N_4784);
nand U4946 (N_4946,N_4664,N_4612);
nor U4947 (N_4947,N_4640,N_4694);
nand U4948 (N_4948,N_4786,N_4770);
and U4949 (N_4949,N_4628,N_4604);
and U4950 (N_4950,N_4714,N_4616);
and U4951 (N_4951,N_4655,N_4766);
nor U4952 (N_4952,N_4677,N_4780);
or U4953 (N_4953,N_4673,N_4642);
nand U4954 (N_4954,N_4664,N_4613);
or U4955 (N_4955,N_4625,N_4774);
nand U4956 (N_4956,N_4633,N_4686);
or U4957 (N_4957,N_4748,N_4668);
xnor U4958 (N_4958,N_4682,N_4695);
nor U4959 (N_4959,N_4675,N_4696);
nor U4960 (N_4960,N_4747,N_4624);
and U4961 (N_4961,N_4674,N_4603);
or U4962 (N_4962,N_4718,N_4762);
nand U4963 (N_4963,N_4632,N_4700);
nor U4964 (N_4964,N_4777,N_4784);
xor U4965 (N_4965,N_4663,N_4690);
nand U4966 (N_4966,N_4736,N_4605);
nand U4967 (N_4967,N_4707,N_4623);
and U4968 (N_4968,N_4738,N_4754);
and U4969 (N_4969,N_4654,N_4759);
xor U4970 (N_4970,N_4695,N_4616);
and U4971 (N_4971,N_4628,N_4662);
and U4972 (N_4972,N_4651,N_4753);
nor U4973 (N_4973,N_4786,N_4654);
nor U4974 (N_4974,N_4706,N_4770);
and U4975 (N_4975,N_4733,N_4710);
and U4976 (N_4976,N_4736,N_4730);
or U4977 (N_4977,N_4673,N_4757);
nand U4978 (N_4978,N_4684,N_4672);
or U4979 (N_4979,N_4729,N_4670);
nor U4980 (N_4980,N_4636,N_4696);
or U4981 (N_4981,N_4796,N_4746);
or U4982 (N_4982,N_4796,N_4707);
and U4983 (N_4983,N_4744,N_4714);
nand U4984 (N_4984,N_4675,N_4661);
nand U4985 (N_4985,N_4615,N_4656);
nand U4986 (N_4986,N_4667,N_4795);
nor U4987 (N_4987,N_4607,N_4675);
and U4988 (N_4988,N_4666,N_4770);
nand U4989 (N_4989,N_4747,N_4799);
nor U4990 (N_4990,N_4682,N_4775);
and U4991 (N_4991,N_4695,N_4716);
nand U4992 (N_4992,N_4643,N_4665);
or U4993 (N_4993,N_4762,N_4773);
nand U4994 (N_4994,N_4669,N_4626);
nor U4995 (N_4995,N_4770,N_4782);
nand U4996 (N_4996,N_4731,N_4753);
nand U4997 (N_4997,N_4714,N_4717);
and U4998 (N_4998,N_4651,N_4767);
nand U4999 (N_4999,N_4676,N_4717);
nor UO_0 (O_0,N_4884,N_4925);
xnor UO_1 (O_1,N_4874,N_4941);
xor UO_2 (O_2,N_4830,N_4958);
and UO_3 (O_3,N_4858,N_4851);
nor UO_4 (O_4,N_4934,N_4987);
nor UO_5 (O_5,N_4881,N_4855);
or UO_6 (O_6,N_4914,N_4826);
nor UO_7 (O_7,N_4857,N_4953);
xnor UO_8 (O_8,N_4901,N_4813);
nand UO_9 (O_9,N_4908,N_4880);
xnor UO_10 (O_10,N_4899,N_4823);
nor UO_11 (O_11,N_4814,N_4907);
and UO_12 (O_12,N_4973,N_4936);
and UO_13 (O_13,N_4837,N_4913);
or UO_14 (O_14,N_4897,N_4910);
and UO_15 (O_15,N_4853,N_4892);
nand UO_16 (O_16,N_4954,N_4985);
nor UO_17 (O_17,N_4803,N_4850);
nor UO_18 (O_18,N_4902,N_4950);
and UO_19 (O_19,N_4979,N_4903);
xor UO_20 (O_20,N_4854,N_4801);
or UO_21 (O_21,N_4877,N_4905);
or UO_22 (O_22,N_4827,N_4939);
and UO_23 (O_23,N_4832,N_4983);
or UO_24 (O_24,N_4923,N_4878);
xor UO_25 (O_25,N_4821,N_4900);
and UO_26 (O_26,N_4932,N_4862);
nor UO_27 (O_27,N_4944,N_4842);
nor UO_28 (O_28,N_4981,N_4834);
nand UO_29 (O_29,N_4852,N_4964);
nor UO_30 (O_30,N_4848,N_4949);
or UO_31 (O_31,N_4894,N_4816);
or UO_32 (O_32,N_4806,N_4928);
nor UO_33 (O_33,N_4864,N_4911);
or UO_34 (O_34,N_4906,N_4835);
nor UO_35 (O_35,N_4969,N_4976);
nor UO_36 (O_36,N_4838,N_4990);
nand UO_37 (O_37,N_4868,N_4999);
and UO_38 (O_38,N_4996,N_4933);
nand UO_39 (O_39,N_4943,N_4922);
and UO_40 (O_40,N_4840,N_4822);
xor UO_41 (O_41,N_4886,N_4945);
nor UO_42 (O_42,N_4815,N_4805);
and UO_43 (O_43,N_4918,N_4810);
and UO_44 (O_44,N_4970,N_4982);
nor UO_45 (O_45,N_4825,N_4819);
and UO_46 (O_46,N_4817,N_4802);
or UO_47 (O_47,N_4887,N_4808);
xnor UO_48 (O_48,N_4938,N_4807);
and UO_49 (O_49,N_4866,N_4980);
or UO_50 (O_50,N_4927,N_4948);
or UO_51 (O_51,N_4869,N_4812);
nor UO_52 (O_52,N_4972,N_4820);
or UO_53 (O_53,N_4867,N_4829);
or UO_54 (O_54,N_4861,N_4818);
and UO_55 (O_55,N_4860,N_4916);
nor UO_56 (O_56,N_4912,N_4849);
or UO_57 (O_57,N_4919,N_4891);
or UO_58 (O_58,N_4856,N_4844);
or UO_59 (O_59,N_4909,N_4859);
nor UO_60 (O_60,N_4841,N_4847);
and UO_61 (O_61,N_4800,N_4872);
nand UO_62 (O_62,N_4957,N_4968);
or UO_63 (O_63,N_4967,N_4839);
and UO_64 (O_64,N_4893,N_4896);
or UO_65 (O_65,N_4951,N_4870);
nand UO_66 (O_66,N_4929,N_4947);
and UO_67 (O_67,N_4963,N_4921);
nor UO_68 (O_68,N_4809,N_4833);
and UO_69 (O_69,N_4875,N_4966);
and UO_70 (O_70,N_4811,N_4955);
and UO_71 (O_71,N_4879,N_4975);
nand UO_72 (O_72,N_4882,N_4930);
xor UO_73 (O_73,N_4865,N_4991);
nand UO_74 (O_74,N_4846,N_4989);
or UO_75 (O_75,N_4959,N_4942);
and UO_76 (O_76,N_4920,N_4876);
xor UO_77 (O_77,N_4995,N_4831);
nand UO_78 (O_78,N_4828,N_4997);
nand UO_79 (O_79,N_4915,N_4940);
and UO_80 (O_80,N_4984,N_4935);
nor UO_81 (O_81,N_4836,N_4931);
nor UO_82 (O_82,N_4883,N_4890);
xnor UO_83 (O_83,N_4824,N_4889);
nor UO_84 (O_84,N_4962,N_4895);
or UO_85 (O_85,N_4960,N_4845);
nor UO_86 (O_86,N_4885,N_4994);
and UO_87 (O_87,N_4946,N_4904);
nand UO_88 (O_88,N_4986,N_4998);
nor UO_89 (O_89,N_4926,N_4993);
and UO_90 (O_90,N_4977,N_4988);
nor UO_91 (O_91,N_4924,N_4804);
nand UO_92 (O_92,N_4888,N_4971);
nor UO_93 (O_93,N_4961,N_4992);
xnor UO_94 (O_94,N_4843,N_4871);
nand UO_95 (O_95,N_4952,N_4873);
or UO_96 (O_96,N_4978,N_4956);
nor UO_97 (O_97,N_4863,N_4965);
or UO_98 (O_98,N_4917,N_4974);
and UO_99 (O_99,N_4937,N_4898);
and UO_100 (O_100,N_4923,N_4896);
or UO_101 (O_101,N_4834,N_4984);
or UO_102 (O_102,N_4926,N_4898);
nand UO_103 (O_103,N_4897,N_4929);
nand UO_104 (O_104,N_4910,N_4871);
and UO_105 (O_105,N_4900,N_4933);
nand UO_106 (O_106,N_4882,N_4843);
and UO_107 (O_107,N_4863,N_4963);
nor UO_108 (O_108,N_4956,N_4866);
or UO_109 (O_109,N_4823,N_4951);
nor UO_110 (O_110,N_4818,N_4815);
and UO_111 (O_111,N_4995,N_4869);
nand UO_112 (O_112,N_4841,N_4911);
or UO_113 (O_113,N_4826,N_4833);
or UO_114 (O_114,N_4882,N_4896);
or UO_115 (O_115,N_4922,N_4948);
or UO_116 (O_116,N_4955,N_4870);
and UO_117 (O_117,N_4817,N_4985);
xnor UO_118 (O_118,N_4853,N_4820);
or UO_119 (O_119,N_4935,N_4864);
nand UO_120 (O_120,N_4890,N_4912);
or UO_121 (O_121,N_4990,N_4868);
and UO_122 (O_122,N_4850,N_4897);
nand UO_123 (O_123,N_4869,N_4881);
or UO_124 (O_124,N_4869,N_4873);
xnor UO_125 (O_125,N_4928,N_4869);
or UO_126 (O_126,N_4936,N_4947);
nor UO_127 (O_127,N_4807,N_4942);
or UO_128 (O_128,N_4906,N_4913);
xnor UO_129 (O_129,N_4811,N_4933);
or UO_130 (O_130,N_4910,N_4808);
or UO_131 (O_131,N_4893,N_4885);
or UO_132 (O_132,N_4996,N_4873);
and UO_133 (O_133,N_4927,N_4959);
or UO_134 (O_134,N_4959,N_4912);
and UO_135 (O_135,N_4801,N_4934);
or UO_136 (O_136,N_4977,N_4924);
and UO_137 (O_137,N_4806,N_4860);
nor UO_138 (O_138,N_4934,N_4813);
nand UO_139 (O_139,N_4833,N_4945);
or UO_140 (O_140,N_4876,N_4957);
nand UO_141 (O_141,N_4963,N_4848);
or UO_142 (O_142,N_4812,N_4905);
and UO_143 (O_143,N_4832,N_4872);
or UO_144 (O_144,N_4911,N_4948);
nand UO_145 (O_145,N_4805,N_4848);
nand UO_146 (O_146,N_4841,N_4983);
nand UO_147 (O_147,N_4861,N_4834);
or UO_148 (O_148,N_4876,N_4911);
and UO_149 (O_149,N_4810,N_4973);
xnor UO_150 (O_150,N_4882,N_4983);
or UO_151 (O_151,N_4946,N_4816);
nand UO_152 (O_152,N_4962,N_4896);
and UO_153 (O_153,N_4866,N_4849);
or UO_154 (O_154,N_4861,N_4801);
xnor UO_155 (O_155,N_4939,N_4941);
nor UO_156 (O_156,N_4805,N_4934);
nand UO_157 (O_157,N_4981,N_4959);
nor UO_158 (O_158,N_4954,N_4864);
and UO_159 (O_159,N_4847,N_4925);
xor UO_160 (O_160,N_4848,N_4859);
and UO_161 (O_161,N_4931,N_4866);
nor UO_162 (O_162,N_4950,N_4975);
and UO_163 (O_163,N_4892,N_4834);
or UO_164 (O_164,N_4998,N_4997);
nand UO_165 (O_165,N_4926,N_4911);
nor UO_166 (O_166,N_4828,N_4999);
and UO_167 (O_167,N_4963,N_4877);
nor UO_168 (O_168,N_4863,N_4956);
and UO_169 (O_169,N_4847,N_4938);
or UO_170 (O_170,N_4997,N_4980);
nand UO_171 (O_171,N_4898,N_4837);
nor UO_172 (O_172,N_4974,N_4983);
and UO_173 (O_173,N_4928,N_4823);
nand UO_174 (O_174,N_4898,N_4872);
and UO_175 (O_175,N_4992,N_4902);
nand UO_176 (O_176,N_4931,N_4835);
or UO_177 (O_177,N_4953,N_4962);
nor UO_178 (O_178,N_4880,N_4982);
nor UO_179 (O_179,N_4825,N_4810);
or UO_180 (O_180,N_4848,N_4962);
nand UO_181 (O_181,N_4877,N_4993);
or UO_182 (O_182,N_4957,N_4836);
and UO_183 (O_183,N_4840,N_4839);
nor UO_184 (O_184,N_4971,N_4814);
xnor UO_185 (O_185,N_4833,N_4804);
and UO_186 (O_186,N_4835,N_4970);
nand UO_187 (O_187,N_4969,N_4925);
or UO_188 (O_188,N_4882,N_4927);
and UO_189 (O_189,N_4930,N_4891);
nor UO_190 (O_190,N_4815,N_4933);
nor UO_191 (O_191,N_4880,N_4947);
and UO_192 (O_192,N_4858,N_4859);
and UO_193 (O_193,N_4974,N_4839);
nor UO_194 (O_194,N_4970,N_4935);
and UO_195 (O_195,N_4880,N_4914);
and UO_196 (O_196,N_4890,N_4862);
or UO_197 (O_197,N_4929,N_4996);
xnor UO_198 (O_198,N_4904,N_4894);
xnor UO_199 (O_199,N_4893,N_4940);
and UO_200 (O_200,N_4970,N_4859);
or UO_201 (O_201,N_4914,N_4861);
nand UO_202 (O_202,N_4886,N_4923);
nor UO_203 (O_203,N_4917,N_4877);
and UO_204 (O_204,N_4885,N_4869);
and UO_205 (O_205,N_4844,N_4981);
nor UO_206 (O_206,N_4801,N_4943);
nor UO_207 (O_207,N_4849,N_4900);
nand UO_208 (O_208,N_4819,N_4856);
and UO_209 (O_209,N_4896,N_4876);
nor UO_210 (O_210,N_4847,N_4832);
nand UO_211 (O_211,N_4893,N_4984);
or UO_212 (O_212,N_4868,N_4901);
and UO_213 (O_213,N_4829,N_4931);
and UO_214 (O_214,N_4823,N_4969);
nor UO_215 (O_215,N_4983,N_4858);
or UO_216 (O_216,N_4861,N_4879);
or UO_217 (O_217,N_4910,N_4965);
nand UO_218 (O_218,N_4830,N_4901);
and UO_219 (O_219,N_4920,N_4899);
or UO_220 (O_220,N_4900,N_4880);
nand UO_221 (O_221,N_4823,N_4839);
or UO_222 (O_222,N_4959,N_4825);
or UO_223 (O_223,N_4824,N_4980);
nand UO_224 (O_224,N_4927,N_4986);
xnor UO_225 (O_225,N_4901,N_4933);
or UO_226 (O_226,N_4992,N_4896);
nor UO_227 (O_227,N_4972,N_4834);
nor UO_228 (O_228,N_4975,N_4918);
or UO_229 (O_229,N_4835,N_4822);
nor UO_230 (O_230,N_4907,N_4825);
or UO_231 (O_231,N_4956,N_4920);
or UO_232 (O_232,N_4820,N_4892);
nand UO_233 (O_233,N_4837,N_4892);
nand UO_234 (O_234,N_4822,N_4859);
or UO_235 (O_235,N_4868,N_4933);
nand UO_236 (O_236,N_4995,N_4964);
nor UO_237 (O_237,N_4967,N_4904);
or UO_238 (O_238,N_4917,N_4973);
nand UO_239 (O_239,N_4858,N_4861);
and UO_240 (O_240,N_4861,N_4868);
nor UO_241 (O_241,N_4875,N_4984);
nand UO_242 (O_242,N_4939,N_4859);
nand UO_243 (O_243,N_4980,N_4894);
nand UO_244 (O_244,N_4852,N_4868);
nor UO_245 (O_245,N_4993,N_4837);
nor UO_246 (O_246,N_4876,N_4904);
nor UO_247 (O_247,N_4841,N_4998);
and UO_248 (O_248,N_4983,N_4818);
nor UO_249 (O_249,N_4898,N_4905);
and UO_250 (O_250,N_4986,N_4934);
and UO_251 (O_251,N_4894,N_4930);
nor UO_252 (O_252,N_4850,N_4992);
nand UO_253 (O_253,N_4879,N_4993);
nor UO_254 (O_254,N_4810,N_4951);
nor UO_255 (O_255,N_4952,N_4951);
nand UO_256 (O_256,N_4960,N_4929);
and UO_257 (O_257,N_4931,N_4939);
nor UO_258 (O_258,N_4816,N_4966);
nor UO_259 (O_259,N_4846,N_4844);
and UO_260 (O_260,N_4975,N_4985);
xor UO_261 (O_261,N_4830,N_4915);
nor UO_262 (O_262,N_4943,N_4960);
and UO_263 (O_263,N_4813,N_4816);
nor UO_264 (O_264,N_4957,N_4984);
nor UO_265 (O_265,N_4817,N_4867);
xnor UO_266 (O_266,N_4858,N_4831);
and UO_267 (O_267,N_4891,N_4994);
xor UO_268 (O_268,N_4859,N_4988);
nor UO_269 (O_269,N_4913,N_4857);
xnor UO_270 (O_270,N_4838,N_4897);
nand UO_271 (O_271,N_4968,N_4812);
nand UO_272 (O_272,N_4854,N_4842);
or UO_273 (O_273,N_4947,N_4939);
or UO_274 (O_274,N_4994,N_4863);
nor UO_275 (O_275,N_4932,N_4908);
and UO_276 (O_276,N_4973,N_4870);
or UO_277 (O_277,N_4801,N_4963);
xnor UO_278 (O_278,N_4828,N_4990);
and UO_279 (O_279,N_4971,N_4965);
nor UO_280 (O_280,N_4915,N_4843);
or UO_281 (O_281,N_4896,N_4979);
nor UO_282 (O_282,N_4916,N_4991);
or UO_283 (O_283,N_4957,N_4977);
nor UO_284 (O_284,N_4940,N_4952);
or UO_285 (O_285,N_4938,N_4924);
nand UO_286 (O_286,N_4912,N_4873);
nor UO_287 (O_287,N_4864,N_4801);
nand UO_288 (O_288,N_4950,N_4876);
and UO_289 (O_289,N_4955,N_4932);
nand UO_290 (O_290,N_4896,N_4978);
xnor UO_291 (O_291,N_4935,N_4990);
or UO_292 (O_292,N_4867,N_4888);
nand UO_293 (O_293,N_4934,N_4833);
or UO_294 (O_294,N_4826,N_4932);
or UO_295 (O_295,N_4858,N_4838);
nor UO_296 (O_296,N_4949,N_4872);
xnor UO_297 (O_297,N_4954,N_4925);
or UO_298 (O_298,N_4809,N_4914);
nor UO_299 (O_299,N_4843,N_4976);
xor UO_300 (O_300,N_4878,N_4921);
xor UO_301 (O_301,N_4955,N_4961);
nand UO_302 (O_302,N_4851,N_4857);
xnor UO_303 (O_303,N_4802,N_4835);
and UO_304 (O_304,N_4865,N_4802);
and UO_305 (O_305,N_4876,N_4875);
nand UO_306 (O_306,N_4914,N_4802);
and UO_307 (O_307,N_4872,N_4867);
and UO_308 (O_308,N_4833,N_4978);
xor UO_309 (O_309,N_4891,N_4903);
nand UO_310 (O_310,N_4883,N_4813);
or UO_311 (O_311,N_4901,N_4932);
or UO_312 (O_312,N_4892,N_4868);
nand UO_313 (O_313,N_4960,N_4991);
nor UO_314 (O_314,N_4845,N_4982);
nor UO_315 (O_315,N_4875,N_4985);
or UO_316 (O_316,N_4907,N_4868);
or UO_317 (O_317,N_4912,N_4940);
or UO_318 (O_318,N_4929,N_4999);
nand UO_319 (O_319,N_4983,N_4851);
or UO_320 (O_320,N_4807,N_4929);
and UO_321 (O_321,N_4920,N_4874);
and UO_322 (O_322,N_4867,N_4975);
or UO_323 (O_323,N_4903,N_4911);
and UO_324 (O_324,N_4961,N_4972);
nand UO_325 (O_325,N_4955,N_4904);
nor UO_326 (O_326,N_4927,N_4968);
nor UO_327 (O_327,N_4817,N_4943);
nand UO_328 (O_328,N_4974,N_4884);
and UO_329 (O_329,N_4983,N_4973);
nor UO_330 (O_330,N_4834,N_4894);
nand UO_331 (O_331,N_4885,N_4946);
or UO_332 (O_332,N_4994,N_4912);
or UO_333 (O_333,N_4981,N_4847);
or UO_334 (O_334,N_4950,N_4833);
nand UO_335 (O_335,N_4812,N_4998);
and UO_336 (O_336,N_4873,N_4985);
nand UO_337 (O_337,N_4978,N_4820);
and UO_338 (O_338,N_4876,N_4987);
and UO_339 (O_339,N_4892,N_4897);
nor UO_340 (O_340,N_4841,N_4910);
nor UO_341 (O_341,N_4891,N_4825);
or UO_342 (O_342,N_4863,N_4930);
nor UO_343 (O_343,N_4905,N_4961);
and UO_344 (O_344,N_4836,N_4923);
and UO_345 (O_345,N_4812,N_4868);
nand UO_346 (O_346,N_4985,N_4951);
and UO_347 (O_347,N_4811,N_4975);
and UO_348 (O_348,N_4944,N_4905);
and UO_349 (O_349,N_4951,N_4844);
xor UO_350 (O_350,N_4900,N_4878);
or UO_351 (O_351,N_4976,N_4917);
xor UO_352 (O_352,N_4911,N_4979);
xor UO_353 (O_353,N_4856,N_4867);
xor UO_354 (O_354,N_4854,N_4823);
nor UO_355 (O_355,N_4879,N_4941);
nand UO_356 (O_356,N_4902,N_4895);
nor UO_357 (O_357,N_4855,N_4884);
nor UO_358 (O_358,N_4941,N_4866);
and UO_359 (O_359,N_4880,N_4967);
and UO_360 (O_360,N_4974,N_4830);
or UO_361 (O_361,N_4959,N_4882);
or UO_362 (O_362,N_4937,N_4825);
or UO_363 (O_363,N_4968,N_4956);
nand UO_364 (O_364,N_4855,N_4826);
or UO_365 (O_365,N_4857,N_4842);
or UO_366 (O_366,N_4891,N_4944);
nand UO_367 (O_367,N_4965,N_4990);
nand UO_368 (O_368,N_4939,N_4810);
or UO_369 (O_369,N_4915,N_4985);
and UO_370 (O_370,N_4991,N_4893);
or UO_371 (O_371,N_4888,N_4970);
xor UO_372 (O_372,N_4879,N_4869);
and UO_373 (O_373,N_4810,N_4949);
and UO_374 (O_374,N_4924,N_4909);
xnor UO_375 (O_375,N_4975,N_4932);
and UO_376 (O_376,N_4966,N_4919);
nand UO_377 (O_377,N_4869,N_4950);
or UO_378 (O_378,N_4911,N_4986);
nor UO_379 (O_379,N_4854,N_4973);
or UO_380 (O_380,N_4935,N_4996);
nand UO_381 (O_381,N_4971,N_4948);
nor UO_382 (O_382,N_4882,N_4895);
and UO_383 (O_383,N_4814,N_4961);
nand UO_384 (O_384,N_4870,N_4804);
and UO_385 (O_385,N_4989,N_4974);
xor UO_386 (O_386,N_4987,N_4948);
nor UO_387 (O_387,N_4987,N_4885);
and UO_388 (O_388,N_4830,N_4816);
xor UO_389 (O_389,N_4982,N_4841);
xnor UO_390 (O_390,N_4961,N_4838);
nor UO_391 (O_391,N_4994,N_4978);
nor UO_392 (O_392,N_4987,N_4852);
and UO_393 (O_393,N_4918,N_4998);
nor UO_394 (O_394,N_4863,N_4903);
nand UO_395 (O_395,N_4998,N_4955);
nand UO_396 (O_396,N_4881,N_4906);
or UO_397 (O_397,N_4887,N_4997);
nor UO_398 (O_398,N_4862,N_4888);
nand UO_399 (O_399,N_4937,N_4971);
or UO_400 (O_400,N_4996,N_4815);
or UO_401 (O_401,N_4839,N_4936);
and UO_402 (O_402,N_4849,N_4854);
xor UO_403 (O_403,N_4926,N_4869);
nor UO_404 (O_404,N_4939,N_4934);
xor UO_405 (O_405,N_4906,N_4804);
nand UO_406 (O_406,N_4820,N_4986);
or UO_407 (O_407,N_4903,N_4982);
nor UO_408 (O_408,N_4971,N_4847);
xnor UO_409 (O_409,N_4972,N_4836);
nand UO_410 (O_410,N_4848,N_4925);
nand UO_411 (O_411,N_4845,N_4989);
nor UO_412 (O_412,N_4933,N_4899);
or UO_413 (O_413,N_4828,N_4850);
and UO_414 (O_414,N_4905,N_4923);
nor UO_415 (O_415,N_4808,N_4953);
and UO_416 (O_416,N_4948,N_4864);
nand UO_417 (O_417,N_4877,N_4817);
nor UO_418 (O_418,N_4836,N_4937);
or UO_419 (O_419,N_4944,N_4836);
and UO_420 (O_420,N_4913,N_4935);
or UO_421 (O_421,N_4935,N_4917);
and UO_422 (O_422,N_4868,N_4960);
nand UO_423 (O_423,N_4977,N_4981);
or UO_424 (O_424,N_4882,N_4965);
nor UO_425 (O_425,N_4801,N_4953);
or UO_426 (O_426,N_4824,N_4838);
or UO_427 (O_427,N_4858,N_4870);
nand UO_428 (O_428,N_4905,N_4952);
and UO_429 (O_429,N_4912,N_4988);
or UO_430 (O_430,N_4823,N_4985);
xor UO_431 (O_431,N_4967,N_4884);
xnor UO_432 (O_432,N_4901,N_4879);
nor UO_433 (O_433,N_4926,N_4870);
xnor UO_434 (O_434,N_4822,N_4999);
nor UO_435 (O_435,N_4895,N_4829);
nor UO_436 (O_436,N_4808,N_4922);
or UO_437 (O_437,N_4857,N_4924);
xnor UO_438 (O_438,N_4948,N_4818);
and UO_439 (O_439,N_4871,N_4872);
nand UO_440 (O_440,N_4974,N_4857);
nor UO_441 (O_441,N_4824,N_4832);
nor UO_442 (O_442,N_4846,N_4856);
nand UO_443 (O_443,N_4826,N_4894);
and UO_444 (O_444,N_4953,N_4819);
nor UO_445 (O_445,N_4949,N_4973);
nor UO_446 (O_446,N_4980,N_4821);
xnor UO_447 (O_447,N_4886,N_4904);
nand UO_448 (O_448,N_4968,N_4899);
or UO_449 (O_449,N_4879,N_4899);
or UO_450 (O_450,N_4841,N_4957);
or UO_451 (O_451,N_4812,N_4896);
nor UO_452 (O_452,N_4972,N_4911);
and UO_453 (O_453,N_4870,N_4902);
nor UO_454 (O_454,N_4879,N_4994);
nand UO_455 (O_455,N_4975,N_4904);
or UO_456 (O_456,N_4945,N_4972);
or UO_457 (O_457,N_4997,N_4944);
nor UO_458 (O_458,N_4919,N_4807);
nand UO_459 (O_459,N_4800,N_4846);
nand UO_460 (O_460,N_4949,N_4894);
and UO_461 (O_461,N_4859,N_4806);
and UO_462 (O_462,N_4995,N_4809);
and UO_463 (O_463,N_4931,N_4874);
nor UO_464 (O_464,N_4909,N_4914);
nand UO_465 (O_465,N_4816,N_4989);
and UO_466 (O_466,N_4958,N_4980);
nand UO_467 (O_467,N_4930,N_4995);
nand UO_468 (O_468,N_4824,N_4978);
and UO_469 (O_469,N_4901,N_4917);
or UO_470 (O_470,N_4892,N_4970);
nor UO_471 (O_471,N_4874,N_4817);
or UO_472 (O_472,N_4999,N_4887);
nand UO_473 (O_473,N_4861,N_4803);
nor UO_474 (O_474,N_4830,N_4841);
nor UO_475 (O_475,N_4859,N_4953);
or UO_476 (O_476,N_4833,N_4997);
nor UO_477 (O_477,N_4893,N_4907);
nor UO_478 (O_478,N_4907,N_4842);
nor UO_479 (O_479,N_4969,N_4875);
nand UO_480 (O_480,N_4945,N_4936);
or UO_481 (O_481,N_4930,N_4862);
or UO_482 (O_482,N_4916,N_4840);
or UO_483 (O_483,N_4897,N_4816);
or UO_484 (O_484,N_4814,N_4987);
nand UO_485 (O_485,N_4923,N_4907);
nand UO_486 (O_486,N_4827,N_4805);
or UO_487 (O_487,N_4990,N_4947);
nand UO_488 (O_488,N_4901,N_4989);
nor UO_489 (O_489,N_4941,N_4947);
or UO_490 (O_490,N_4843,N_4963);
and UO_491 (O_491,N_4937,N_4876);
nand UO_492 (O_492,N_4814,N_4922);
nand UO_493 (O_493,N_4805,N_4943);
or UO_494 (O_494,N_4874,N_4953);
or UO_495 (O_495,N_4962,N_4847);
xnor UO_496 (O_496,N_4923,N_4852);
or UO_497 (O_497,N_4966,N_4868);
nor UO_498 (O_498,N_4843,N_4904);
nor UO_499 (O_499,N_4831,N_4972);
nor UO_500 (O_500,N_4992,N_4801);
nor UO_501 (O_501,N_4856,N_4886);
or UO_502 (O_502,N_4828,N_4994);
nor UO_503 (O_503,N_4948,N_4930);
or UO_504 (O_504,N_4830,N_4835);
and UO_505 (O_505,N_4960,N_4827);
and UO_506 (O_506,N_4961,N_4853);
and UO_507 (O_507,N_4991,N_4857);
nor UO_508 (O_508,N_4993,N_4937);
nor UO_509 (O_509,N_4946,N_4992);
or UO_510 (O_510,N_4911,N_4900);
and UO_511 (O_511,N_4987,N_4967);
or UO_512 (O_512,N_4981,N_4934);
nor UO_513 (O_513,N_4882,N_4801);
xor UO_514 (O_514,N_4948,N_4991);
nand UO_515 (O_515,N_4944,N_4949);
nand UO_516 (O_516,N_4946,N_4921);
nand UO_517 (O_517,N_4940,N_4854);
or UO_518 (O_518,N_4985,N_4966);
nand UO_519 (O_519,N_4850,N_4823);
nand UO_520 (O_520,N_4875,N_4943);
xnor UO_521 (O_521,N_4896,N_4941);
or UO_522 (O_522,N_4824,N_4844);
nand UO_523 (O_523,N_4899,N_4984);
and UO_524 (O_524,N_4979,N_4946);
nand UO_525 (O_525,N_4981,N_4816);
nor UO_526 (O_526,N_4957,N_4802);
and UO_527 (O_527,N_4884,N_4913);
and UO_528 (O_528,N_4897,N_4805);
or UO_529 (O_529,N_4842,N_4819);
nor UO_530 (O_530,N_4986,N_4946);
or UO_531 (O_531,N_4862,N_4962);
nor UO_532 (O_532,N_4852,N_4861);
nor UO_533 (O_533,N_4949,N_4868);
and UO_534 (O_534,N_4963,N_4870);
nand UO_535 (O_535,N_4881,N_4816);
nand UO_536 (O_536,N_4971,N_4918);
nor UO_537 (O_537,N_4850,N_4976);
nor UO_538 (O_538,N_4993,N_4941);
nand UO_539 (O_539,N_4802,N_4888);
and UO_540 (O_540,N_4979,N_4961);
nand UO_541 (O_541,N_4853,N_4955);
and UO_542 (O_542,N_4997,N_4810);
and UO_543 (O_543,N_4978,N_4892);
xor UO_544 (O_544,N_4812,N_4891);
and UO_545 (O_545,N_4900,N_4893);
nand UO_546 (O_546,N_4967,N_4837);
nor UO_547 (O_547,N_4941,N_4886);
nand UO_548 (O_548,N_4815,N_4968);
nand UO_549 (O_549,N_4991,N_4996);
or UO_550 (O_550,N_4943,N_4833);
nor UO_551 (O_551,N_4917,N_4912);
xnor UO_552 (O_552,N_4863,N_4923);
and UO_553 (O_553,N_4865,N_4939);
and UO_554 (O_554,N_4866,N_4822);
nand UO_555 (O_555,N_4894,N_4987);
nor UO_556 (O_556,N_4841,N_4896);
xnor UO_557 (O_557,N_4899,N_4889);
and UO_558 (O_558,N_4979,N_4854);
nand UO_559 (O_559,N_4912,N_4905);
nand UO_560 (O_560,N_4819,N_4875);
or UO_561 (O_561,N_4963,N_4827);
nor UO_562 (O_562,N_4852,N_4983);
or UO_563 (O_563,N_4832,N_4931);
or UO_564 (O_564,N_4987,N_4961);
nand UO_565 (O_565,N_4865,N_4993);
xnor UO_566 (O_566,N_4962,N_4832);
nand UO_567 (O_567,N_4993,N_4990);
and UO_568 (O_568,N_4913,N_4871);
and UO_569 (O_569,N_4923,N_4999);
nand UO_570 (O_570,N_4808,N_4959);
nand UO_571 (O_571,N_4960,N_4927);
nand UO_572 (O_572,N_4902,N_4991);
or UO_573 (O_573,N_4966,N_4811);
and UO_574 (O_574,N_4804,N_4823);
nor UO_575 (O_575,N_4882,N_4909);
or UO_576 (O_576,N_4958,N_4884);
or UO_577 (O_577,N_4827,N_4974);
nor UO_578 (O_578,N_4808,N_4884);
or UO_579 (O_579,N_4919,N_4878);
nand UO_580 (O_580,N_4924,N_4846);
nand UO_581 (O_581,N_4823,N_4939);
xnor UO_582 (O_582,N_4975,N_4900);
and UO_583 (O_583,N_4884,N_4987);
xnor UO_584 (O_584,N_4899,N_4979);
nor UO_585 (O_585,N_4864,N_4958);
or UO_586 (O_586,N_4953,N_4891);
and UO_587 (O_587,N_4938,N_4906);
xnor UO_588 (O_588,N_4962,N_4914);
and UO_589 (O_589,N_4880,N_4812);
or UO_590 (O_590,N_4905,N_4886);
xor UO_591 (O_591,N_4891,N_4963);
or UO_592 (O_592,N_4850,N_4847);
nor UO_593 (O_593,N_4902,N_4822);
and UO_594 (O_594,N_4856,N_4919);
xor UO_595 (O_595,N_4887,N_4906);
and UO_596 (O_596,N_4910,N_4805);
or UO_597 (O_597,N_4951,N_4804);
or UO_598 (O_598,N_4979,N_4934);
xor UO_599 (O_599,N_4893,N_4983);
and UO_600 (O_600,N_4983,N_4992);
and UO_601 (O_601,N_4874,N_4814);
or UO_602 (O_602,N_4993,N_4810);
xor UO_603 (O_603,N_4856,N_4939);
or UO_604 (O_604,N_4866,N_4969);
nor UO_605 (O_605,N_4992,N_4962);
xnor UO_606 (O_606,N_4954,N_4823);
and UO_607 (O_607,N_4900,N_4948);
nor UO_608 (O_608,N_4977,N_4810);
and UO_609 (O_609,N_4899,N_4883);
xor UO_610 (O_610,N_4954,N_4858);
nand UO_611 (O_611,N_4930,N_4957);
nor UO_612 (O_612,N_4867,N_4989);
nor UO_613 (O_613,N_4912,N_4834);
and UO_614 (O_614,N_4846,N_4892);
xor UO_615 (O_615,N_4855,N_4871);
xor UO_616 (O_616,N_4859,N_4839);
and UO_617 (O_617,N_4926,N_4979);
and UO_618 (O_618,N_4802,N_4845);
or UO_619 (O_619,N_4947,N_4968);
or UO_620 (O_620,N_4958,N_4806);
and UO_621 (O_621,N_4816,N_4851);
nand UO_622 (O_622,N_4834,N_4868);
and UO_623 (O_623,N_4839,N_4880);
or UO_624 (O_624,N_4910,N_4814);
xnor UO_625 (O_625,N_4934,N_4810);
and UO_626 (O_626,N_4912,N_4869);
or UO_627 (O_627,N_4991,N_4866);
and UO_628 (O_628,N_4972,N_4973);
nand UO_629 (O_629,N_4943,N_4840);
nand UO_630 (O_630,N_4867,N_4923);
nor UO_631 (O_631,N_4843,N_4831);
nand UO_632 (O_632,N_4873,N_4825);
and UO_633 (O_633,N_4940,N_4943);
nor UO_634 (O_634,N_4957,N_4898);
and UO_635 (O_635,N_4944,N_4979);
nor UO_636 (O_636,N_4877,N_4938);
nor UO_637 (O_637,N_4863,N_4833);
nand UO_638 (O_638,N_4890,N_4980);
or UO_639 (O_639,N_4906,N_4929);
nand UO_640 (O_640,N_4933,N_4943);
xor UO_641 (O_641,N_4950,N_4968);
nand UO_642 (O_642,N_4952,N_4919);
or UO_643 (O_643,N_4923,N_4948);
xor UO_644 (O_644,N_4861,N_4977);
nand UO_645 (O_645,N_4871,N_4862);
nand UO_646 (O_646,N_4804,N_4917);
and UO_647 (O_647,N_4921,N_4864);
nand UO_648 (O_648,N_4949,N_4900);
xnor UO_649 (O_649,N_4968,N_4817);
or UO_650 (O_650,N_4965,N_4845);
nor UO_651 (O_651,N_4817,N_4927);
and UO_652 (O_652,N_4988,N_4835);
or UO_653 (O_653,N_4944,N_4845);
nor UO_654 (O_654,N_4950,N_4859);
xnor UO_655 (O_655,N_4896,N_4996);
or UO_656 (O_656,N_4986,N_4992);
or UO_657 (O_657,N_4928,N_4990);
or UO_658 (O_658,N_4905,N_4873);
nand UO_659 (O_659,N_4937,N_4908);
nor UO_660 (O_660,N_4959,N_4972);
or UO_661 (O_661,N_4844,N_4850);
nand UO_662 (O_662,N_4857,N_4900);
nor UO_663 (O_663,N_4900,N_4866);
and UO_664 (O_664,N_4871,N_4880);
nor UO_665 (O_665,N_4853,N_4931);
nor UO_666 (O_666,N_4830,N_4821);
nand UO_667 (O_667,N_4996,N_4813);
nor UO_668 (O_668,N_4859,N_4898);
or UO_669 (O_669,N_4893,N_4986);
or UO_670 (O_670,N_4837,N_4924);
or UO_671 (O_671,N_4909,N_4913);
and UO_672 (O_672,N_4926,N_4904);
nand UO_673 (O_673,N_4964,N_4801);
xor UO_674 (O_674,N_4991,N_4921);
nor UO_675 (O_675,N_4956,N_4928);
nand UO_676 (O_676,N_4866,N_4995);
nor UO_677 (O_677,N_4809,N_4888);
nor UO_678 (O_678,N_4855,N_4859);
and UO_679 (O_679,N_4972,N_4859);
nand UO_680 (O_680,N_4890,N_4908);
or UO_681 (O_681,N_4921,N_4821);
nand UO_682 (O_682,N_4865,N_4887);
nand UO_683 (O_683,N_4987,N_4920);
or UO_684 (O_684,N_4951,N_4982);
nor UO_685 (O_685,N_4848,N_4952);
or UO_686 (O_686,N_4883,N_4848);
or UO_687 (O_687,N_4949,N_4911);
and UO_688 (O_688,N_4930,N_4887);
and UO_689 (O_689,N_4830,N_4914);
nand UO_690 (O_690,N_4919,N_4951);
or UO_691 (O_691,N_4835,N_4860);
or UO_692 (O_692,N_4983,N_4960);
or UO_693 (O_693,N_4902,N_4937);
nand UO_694 (O_694,N_4882,N_4952);
nor UO_695 (O_695,N_4877,N_4821);
nor UO_696 (O_696,N_4957,N_4807);
nor UO_697 (O_697,N_4921,N_4980);
and UO_698 (O_698,N_4957,N_4940);
nor UO_699 (O_699,N_4982,N_4921);
nand UO_700 (O_700,N_4944,N_4811);
nor UO_701 (O_701,N_4867,N_4947);
nand UO_702 (O_702,N_4997,N_4963);
xor UO_703 (O_703,N_4876,N_4932);
nor UO_704 (O_704,N_4995,N_4906);
and UO_705 (O_705,N_4928,N_4829);
xor UO_706 (O_706,N_4818,N_4876);
and UO_707 (O_707,N_4866,N_4824);
or UO_708 (O_708,N_4829,N_4847);
nand UO_709 (O_709,N_4895,N_4886);
or UO_710 (O_710,N_4874,N_4909);
nand UO_711 (O_711,N_4949,N_4828);
nor UO_712 (O_712,N_4966,N_4881);
xor UO_713 (O_713,N_4866,N_4949);
nor UO_714 (O_714,N_4822,N_4813);
nand UO_715 (O_715,N_4872,N_4937);
nand UO_716 (O_716,N_4967,N_4849);
and UO_717 (O_717,N_4954,N_4927);
xor UO_718 (O_718,N_4955,N_4898);
and UO_719 (O_719,N_4835,N_4987);
or UO_720 (O_720,N_4879,N_4961);
xor UO_721 (O_721,N_4974,N_4954);
or UO_722 (O_722,N_4875,N_4913);
nand UO_723 (O_723,N_4863,N_4928);
or UO_724 (O_724,N_4950,N_4835);
nand UO_725 (O_725,N_4843,N_4920);
nand UO_726 (O_726,N_4814,N_4811);
nor UO_727 (O_727,N_4916,N_4843);
nor UO_728 (O_728,N_4853,N_4905);
or UO_729 (O_729,N_4843,N_4983);
nand UO_730 (O_730,N_4928,N_4925);
or UO_731 (O_731,N_4970,N_4864);
xor UO_732 (O_732,N_4917,N_4969);
nand UO_733 (O_733,N_4863,N_4849);
and UO_734 (O_734,N_4867,N_4988);
or UO_735 (O_735,N_4885,N_4887);
or UO_736 (O_736,N_4930,N_4950);
nand UO_737 (O_737,N_4980,N_4823);
nand UO_738 (O_738,N_4951,N_4854);
or UO_739 (O_739,N_4902,N_4883);
and UO_740 (O_740,N_4982,N_4875);
or UO_741 (O_741,N_4851,N_4836);
or UO_742 (O_742,N_4872,N_4989);
or UO_743 (O_743,N_4890,N_4810);
nor UO_744 (O_744,N_4875,N_4926);
nor UO_745 (O_745,N_4964,N_4838);
nand UO_746 (O_746,N_4933,N_4835);
xnor UO_747 (O_747,N_4905,N_4965);
or UO_748 (O_748,N_4850,N_4832);
or UO_749 (O_749,N_4911,N_4874);
or UO_750 (O_750,N_4934,N_4988);
or UO_751 (O_751,N_4935,N_4932);
and UO_752 (O_752,N_4963,N_4973);
nand UO_753 (O_753,N_4896,N_4937);
xnor UO_754 (O_754,N_4935,N_4873);
nor UO_755 (O_755,N_4870,N_4841);
nand UO_756 (O_756,N_4976,N_4955);
or UO_757 (O_757,N_4879,N_4895);
nand UO_758 (O_758,N_4944,N_4858);
nor UO_759 (O_759,N_4960,N_4969);
nand UO_760 (O_760,N_4886,N_4983);
nor UO_761 (O_761,N_4805,N_4803);
nor UO_762 (O_762,N_4807,N_4923);
or UO_763 (O_763,N_4885,N_4881);
nor UO_764 (O_764,N_4976,N_4840);
nor UO_765 (O_765,N_4967,N_4901);
and UO_766 (O_766,N_4924,N_4999);
nand UO_767 (O_767,N_4839,N_4802);
or UO_768 (O_768,N_4816,N_4971);
nor UO_769 (O_769,N_4951,N_4993);
or UO_770 (O_770,N_4962,N_4877);
or UO_771 (O_771,N_4978,N_4893);
xor UO_772 (O_772,N_4921,N_4892);
nor UO_773 (O_773,N_4812,N_4987);
and UO_774 (O_774,N_4920,N_4930);
and UO_775 (O_775,N_4866,N_4993);
xor UO_776 (O_776,N_4923,N_4921);
nor UO_777 (O_777,N_4854,N_4815);
xnor UO_778 (O_778,N_4957,N_4816);
nor UO_779 (O_779,N_4843,N_4928);
nor UO_780 (O_780,N_4971,N_4983);
or UO_781 (O_781,N_4856,N_4911);
nand UO_782 (O_782,N_4827,N_4865);
or UO_783 (O_783,N_4938,N_4921);
nor UO_784 (O_784,N_4963,N_4935);
xnor UO_785 (O_785,N_4849,N_4958);
and UO_786 (O_786,N_4853,N_4863);
nor UO_787 (O_787,N_4814,N_4901);
or UO_788 (O_788,N_4966,N_4900);
nor UO_789 (O_789,N_4993,N_4994);
and UO_790 (O_790,N_4923,N_4861);
or UO_791 (O_791,N_4908,N_4877);
nand UO_792 (O_792,N_4866,N_4951);
xor UO_793 (O_793,N_4928,N_4878);
nand UO_794 (O_794,N_4815,N_4993);
nor UO_795 (O_795,N_4839,N_4992);
nand UO_796 (O_796,N_4905,N_4841);
and UO_797 (O_797,N_4877,N_4957);
nand UO_798 (O_798,N_4811,N_4868);
nand UO_799 (O_799,N_4842,N_4943);
or UO_800 (O_800,N_4898,N_4803);
nand UO_801 (O_801,N_4944,N_4913);
and UO_802 (O_802,N_4963,N_4917);
nor UO_803 (O_803,N_4830,N_4878);
and UO_804 (O_804,N_4931,N_4977);
nand UO_805 (O_805,N_4972,N_4931);
nand UO_806 (O_806,N_4807,N_4911);
or UO_807 (O_807,N_4998,N_4851);
nand UO_808 (O_808,N_4838,N_4962);
or UO_809 (O_809,N_4894,N_4864);
nand UO_810 (O_810,N_4926,N_4931);
xnor UO_811 (O_811,N_4933,N_4957);
nor UO_812 (O_812,N_4809,N_4944);
nand UO_813 (O_813,N_4831,N_4894);
nor UO_814 (O_814,N_4851,N_4877);
xnor UO_815 (O_815,N_4899,N_4848);
and UO_816 (O_816,N_4972,N_4824);
nand UO_817 (O_817,N_4819,N_4944);
xnor UO_818 (O_818,N_4915,N_4824);
or UO_819 (O_819,N_4966,N_4969);
or UO_820 (O_820,N_4820,N_4809);
or UO_821 (O_821,N_4975,N_4841);
or UO_822 (O_822,N_4852,N_4913);
and UO_823 (O_823,N_4989,N_4976);
and UO_824 (O_824,N_4910,N_4962);
and UO_825 (O_825,N_4928,N_4840);
nand UO_826 (O_826,N_4937,N_4890);
or UO_827 (O_827,N_4821,N_4939);
or UO_828 (O_828,N_4975,N_4887);
and UO_829 (O_829,N_4822,N_4838);
or UO_830 (O_830,N_4975,N_4837);
nand UO_831 (O_831,N_4901,N_4942);
xor UO_832 (O_832,N_4913,N_4985);
xor UO_833 (O_833,N_4910,N_4880);
nand UO_834 (O_834,N_4811,N_4863);
nand UO_835 (O_835,N_4953,N_4937);
or UO_836 (O_836,N_4863,N_4950);
or UO_837 (O_837,N_4817,N_4976);
or UO_838 (O_838,N_4913,N_4811);
nand UO_839 (O_839,N_4897,N_4815);
nor UO_840 (O_840,N_4882,N_4976);
nand UO_841 (O_841,N_4970,N_4810);
and UO_842 (O_842,N_4867,N_4836);
xor UO_843 (O_843,N_4966,N_4944);
and UO_844 (O_844,N_4995,N_4853);
nor UO_845 (O_845,N_4988,N_4864);
nand UO_846 (O_846,N_4909,N_4805);
or UO_847 (O_847,N_4956,N_4830);
or UO_848 (O_848,N_4801,N_4978);
or UO_849 (O_849,N_4933,N_4941);
nor UO_850 (O_850,N_4831,N_4973);
nand UO_851 (O_851,N_4860,N_4801);
nor UO_852 (O_852,N_4829,N_4887);
nand UO_853 (O_853,N_4937,N_4918);
nor UO_854 (O_854,N_4890,N_4832);
nor UO_855 (O_855,N_4948,N_4978);
or UO_856 (O_856,N_4939,N_4933);
xnor UO_857 (O_857,N_4917,N_4991);
nor UO_858 (O_858,N_4890,N_4979);
and UO_859 (O_859,N_4809,N_4815);
and UO_860 (O_860,N_4877,N_4859);
or UO_861 (O_861,N_4853,N_4910);
or UO_862 (O_862,N_4921,N_4828);
nor UO_863 (O_863,N_4971,N_4857);
xnor UO_864 (O_864,N_4800,N_4913);
and UO_865 (O_865,N_4821,N_4816);
nor UO_866 (O_866,N_4805,N_4913);
nand UO_867 (O_867,N_4878,N_4826);
xnor UO_868 (O_868,N_4954,N_4973);
nor UO_869 (O_869,N_4855,N_4993);
nor UO_870 (O_870,N_4921,N_4809);
or UO_871 (O_871,N_4864,N_4852);
nand UO_872 (O_872,N_4887,N_4952);
and UO_873 (O_873,N_4874,N_4939);
nor UO_874 (O_874,N_4832,N_4961);
or UO_875 (O_875,N_4954,N_4945);
nand UO_876 (O_876,N_4980,N_4905);
nor UO_877 (O_877,N_4812,N_4847);
or UO_878 (O_878,N_4882,N_4867);
and UO_879 (O_879,N_4883,N_4842);
nand UO_880 (O_880,N_4920,N_4806);
nand UO_881 (O_881,N_4931,N_4917);
or UO_882 (O_882,N_4976,N_4906);
nor UO_883 (O_883,N_4923,N_4822);
or UO_884 (O_884,N_4973,N_4855);
or UO_885 (O_885,N_4991,N_4907);
or UO_886 (O_886,N_4946,N_4819);
xor UO_887 (O_887,N_4895,N_4969);
or UO_888 (O_888,N_4832,N_4841);
and UO_889 (O_889,N_4955,N_4996);
and UO_890 (O_890,N_4935,N_4975);
and UO_891 (O_891,N_4853,N_4984);
and UO_892 (O_892,N_4999,N_4955);
nand UO_893 (O_893,N_4997,N_4884);
nor UO_894 (O_894,N_4827,N_4920);
nand UO_895 (O_895,N_4819,N_4884);
nor UO_896 (O_896,N_4939,N_4841);
nand UO_897 (O_897,N_4974,N_4966);
and UO_898 (O_898,N_4955,N_4839);
nand UO_899 (O_899,N_4831,N_4826);
and UO_900 (O_900,N_4902,N_4952);
nor UO_901 (O_901,N_4849,N_4896);
nand UO_902 (O_902,N_4974,N_4996);
nand UO_903 (O_903,N_4881,N_4848);
nand UO_904 (O_904,N_4916,N_4918);
nand UO_905 (O_905,N_4979,N_4970);
nor UO_906 (O_906,N_4872,N_4954);
or UO_907 (O_907,N_4933,N_4823);
nand UO_908 (O_908,N_4917,N_4989);
nor UO_909 (O_909,N_4934,N_4899);
or UO_910 (O_910,N_4895,N_4815);
xnor UO_911 (O_911,N_4990,N_4863);
nand UO_912 (O_912,N_4932,N_4870);
xor UO_913 (O_913,N_4861,N_4983);
or UO_914 (O_914,N_4844,N_4862);
and UO_915 (O_915,N_4826,N_4884);
or UO_916 (O_916,N_4832,N_4812);
nor UO_917 (O_917,N_4857,N_4828);
nand UO_918 (O_918,N_4897,N_4807);
or UO_919 (O_919,N_4846,N_4963);
and UO_920 (O_920,N_4890,N_4996);
nand UO_921 (O_921,N_4972,N_4987);
or UO_922 (O_922,N_4925,N_4942);
nor UO_923 (O_923,N_4916,N_4803);
or UO_924 (O_924,N_4873,N_4877);
or UO_925 (O_925,N_4900,N_4980);
nor UO_926 (O_926,N_4834,N_4951);
nor UO_927 (O_927,N_4988,N_4898);
nor UO_928 (O_928,N_4991,N_4837);
and UO_929 (O_929,N_4953,N_4951);
nand UO_930 (O_930,N_4864,N_4976);
or UO_931 (O_931,N_4848,N_4892);
nand UO_932 (O_932,N_4992,N_4954);
and UO_933 (O_933,N_4993,N_4919);
or UO_934 (O_934,N_4944,N_4876);
or UO_935 (O_935,N_4907,N_4963);
xnor UO_936 (O_936,N_4979,N_4941);
xnor UO_937 (O_937,N_4827,N_4918);
nor UO_938 (O_938,N_4934,N_4860);
nand UO_939 (O_939,N_4946,N_4959);
nand UO_940 (O_940,N_4947,N_4997);
and UO_941 (O_941,N_4898,N_4820);
xor UO_942 (O_942,N_4854,N_4885);
nor UO_943 (O_943,N_4803,N_4937);
and UO_944 (O_944,N_4810,N_4828);
xnor UO_945 (O_945,N_4938,N_4934);
nand UO_946 (O_946,N_4809,N_4826);
and UO_947 (O_947,N_4983,N_4890);
or UO_948 (O_948,N_4995,N_4870);
xor UO_949 (O_949,N_4818,N_4906);
nand UO_950 (O_950,N_4999,N_4831);
nand UO_951 (O_951,N_4963,N_4912);
and UO_952 (O_952,N_4915,N_4867);
nand UO_953 (O_953,N_4843,N_4872);
xor UO_954 (O_954,N_4879,N_4916);
nor UO_955 (O_955,N_4889,N_4816);
nand UO_956 (O_956,N_4980,N_4964);
or UO_957 (O_957,N_4982,N_4847);
and UO_958 (O_958,N_4850,N_4928);
nor UO_959 (O_959,N_4920,N_4966);
nor UO_960 (O_960,N_4923,N_4845);
or UO_961 (O_961,N_4980,N_4910);
nor UO_962 (O_962,N_4913,N_4915);
and UO_963 (O_963,N_4875,N_4990);
nand UO_964 (O_964,N_4880,N_4943);
nand UO_965 (O_965,N_4943,N_4925);
and UO_966 (O_966,N_4897,N_4935);
nand UO_967 (O_967,N_4907,N_4815);
nand UO_968 (O_968,N_4890,N_4848);
or UO_969 (O_969,N_4843,N_4965);
and UO_970 (O_970,N_4978,N_4816);
and UO_971 (O_971,N_4910,N_4992);
or UO_972 (O_972,N_4831,N_4837);
and UO_973 (O_973,N_4913,N_4844);
nor UO_974 (O_974,N_4948,N_4957);
nor UO_975 (O_975,N_4841,N_4913);
nand UO_976 (O_976,N_4846,N_4811);
nand UO_977 (O_977,N_4822,N_4967);
nand UO_978 (O_978,N_4809,N_4996);
nor UO_979 (O_979,N_4857,N_4840);
nand UO_980 (O_980,N_4984,N_4994);
nand UO_981 (O_981,N_4892,N_4957);
nand UO_982 (O_982,N_4894,N_4947);
or UO_983 (O_983,N_4874,N_4838);
and UO_984 (O_984,N_4859,N_4801);
nor UO_985 (O_985,N_4994,N_4862);
or UO_986 (O_986,N_4802,N_4992);
and UO_987 (O_987,N_4884,N_4954);
and UO_988 (O_988,N_4865,N_4872);
nand UO_989 (O_989,N_4871,N_4984);
or UO_990 (O_990,N_4868,N_4877);
or UO_991 (O_991,N_4844,N_4938);
or UO_992 (O_992,N_4822,N_4895);
nor UO_993 (O_993,N_4849,N_4860);
nor UO_994 (O_994,N_4833,N_4846);
and UO_995 (O_995,N_4807,N_4956);
nor UO_996 (O_996,N_4802,N_4842);
xor UO_997 (O_997,N_4811,N_4845);
xnor UO_998 (O_998,N_4930,N_4923);
nand UO_999 (O_999,N_4875,N_4987);
endmodule