module basic_500_3000_500_50_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_477,In_331);
nand U1 (N_1,In_495,In_37);
and U2 (N_2,In_211,In_459);
or U3 (N_3,In_195,In_475);
or U4 (N_4,In_77,In_476);
and U5 (N_5,In_171,In_167);
nand U6 (N_6,In_122,In_346);
nand U7 (N_7,In_349,In_302);
and U8 (N_8,In_372,In_447);
nor U9 (N_9,In_489,In_401);
nor U10 (N_10,In_449,In_266);
nor U11 (N_11,In_223,In_162);
nor U12 (N_12,In_244,In_370);
nand U13 (N_13,In_281,In_80);
and U14 (N_14,In_61,In_6);
and U15 (N_15,In_201,In_112);
nor U16 (N_16,In_399,In_36);
or U17 (N_17,In_342,In_49);
or U18 (N_18,In_430,In_354);
nand U19 (N_19,In_54,In_200);
and U20 (N_20,In_374,In_91);
or U21 (N_21,In_137,In_294);
and U22 (N_22,In_221,In_395);
and U23 (N_23,In_219,In_472);
and U24 (N_24,In_180,In_404);
or U25 (N_25,In_357,In_499);
nor U26 (N_26,In_166,In_213);
or U27 (N_27,In_460,In_248);
or U28 (N_28,In_194,In_462);
nor U29 (N_29,In_368,In_164);
nor U30 (N_30,In_243,In_156);
nand U31 (N_31,In_301,In_140);
and U32 (N_32,In_13,In_38);
nand U33 (N_33,In_317,In_319);
and U34 (N_34,In_416,In_406);
nor U35 (N_35,In_147,In_226);
or U36 (N_36,In_215,In_242);
nand U37 (N_37,In_239,In_465);
nor U38 (N_38,In_41,In_424);
nand U39 (N_39,In_230,In_407);
nand U40 (N_40,In_310,In_386);
nand U41 (N_41,In_7,In_125);
nor U42 (N_42,In_249,In_102);
or U43 (N_43,In_42,In_139);
or U44 (N_44,In_55,In_116);
and U45 (N_45,In_45,In_29);
or U46 (N_46,In_131,In_78);
or U47 (N_47,In_394,In_245);
and U48 (N_48,In_287,In_9);
nand U49 (N_49,In_99,In_113);
or U50 (N_50,In_56,In_163);
or U51 (N_51,In_385,In_359);
or U52 (N_52,In_47,In_185);
and U53 (N_53,In_121,In_308);
or U54 (N_54,In_8,In_233);
nand U55 (N_55,In_272,In_267);
and U56 (N_56,In_328,In_59);
or U57 (N_57,In_103,In_365);
or U58 (N_58,In_67,In_71);
nor U59 (N_59,In_148,In_280);
nor U60 (N_60,In_182,In_369);
or U61 (N_61,In_312,N_11);
nand U62 (N_62,In_86,In_126);
or U63 (N_63,N_30,In_83);
and U64 (N_64,In_247,In_384);
nor U65 (N_65,In_63,In_145);
nor U66 (N_66,N_5,In_255);
nand U67 (N_67,In_292,In_432);
nand U68 (N_68,In_160,In_389);
nand U69 (N_69,N_48,In_396);
nor U70 (N_70,In_427,In_258);
nor U71 (N_71,In_17,In_332);
or U72 (N_72,N_8,In_144);
nor U73 (N_73,In_20,In_222);
nor U74 (N_74,In_31,In_107);
nor U75 (N_75,In_297,In_471);
nand U76 (N_76,In_498,N_59);
nand U77 (N_77,In_446,In_232);
nand U78 (N_78,In_177,In_345);
and U79 (N_79,In_30,In_228);
or U80 (N_80,In_473,In_106);
and U81 (N_81,In_11,In_174);
nand U82 (N_82,N_26,In_169);
nor U83 (N_83,In_286,In_73);
nand U84 (N_84,In_260,In_313);
and U85 (N_85,N_19,In_5);
nand U86 (N_86,In_420,In_274);
nor U87 (N_87,In_150,In_360);
nor U88 (N_88,In_51,In_358);
or U89 (N_89,N_14,In_277);
and U90 (N_90,In_262,In_237);
xor U91 (N_91,In_75,In_373);
or U92 (N_92,In_143,In_65);
xnor U93 (N_93,N_38,In_190);
and U94 (N_94,In_283,In_253);
nor U95 (N_95,In_241,In_48);
nand U96 (N_96,In_191,In_492);
or U97 (N_97,In_338,In_46);
or U98 (N_98,In_304,In_134);
nand U99 (N_99,In_361,In_377);
nand U100 (N_100,In_28,In_196);
or U101 (N_101,In_161,In_314);
nand U102 (N_102,In_410,In_183);
nor U103 (N_103,In_123,N_23);
nand U104 (N_104,In_326,In_269);
nand U105 (N_105,In_397,In_254);
and U106 (N_106,In_322,In_132);
and U107 (N_107,In_203,In_341);
and U108 (N_108,N_6,In_82);
nor U109 (N_109,N_18,In_275);
nand U110 (N_110,In_484,In_64);
or U111 (N_111,In_480,In_378);
nand U112 (N_112,In_497,In_380);
or U113 (N_113,In_351,In_282);
or U114 (N_114,In_265,In_21);
nor U115 (N_115,In_291,N_22);
and U116 (N_116,In_261,In_97);
or U117 (N_117,In_316,In_325);
nor U118 (N_118,In_375,In_376);
or U119 (N_119,In_426,In_26);
nor U120 (N_120,In_53,In_119);
nand U121 (N_121,In_197,N_41);
nor U122 (N_122,In_273,In_40);
and U123 (N_123,In_408,In_198);
nand U124 (N_124,In_214,In_250);
or U125 (N_125,In_108,In_493);
nor U126 (N_126,N_25,In_165);
nor U127 (N_127,In_300,In_335);
or U128 (N_128,In_176,In_329);
nand U129 (N_129,In_153,In_433);
or U130 (N_130,In_409,In_487);
and U131 (N_131,In_101,In_142);
and U132 (N_132,In_288,In_179);
nor U133 (N_133,In_411,N_103);
and U134 (N_134,N_47,In_189);
nor U135 (N_135,In_16,In_81);
and U136 (N_136,In_417,In_32);
nand U137 (N_137,In_414,In_178);
and U138 (N_138,In_415,N_71);
and U139 (N_139,In_438,In_348);
nor U140 (N_140,In_318,N_13);
or U141 (N_141,In_402,N_106);
nor U142 (N_142,In_138,In_467);
nand U143 (N_143,In_334,N_4);
or U144 (N_144,N_113,N_21);
nor U145 (N_145,N_100,In_405);
nor U146 (N_146,In_23,In_79);
nand U147 (N_147,In_74,In_295);
nor U148 (N_148,In_175,In_238);
nand U149 (N_149,In_251,In_343);
and U150 (N_150,In_57,In_383);
nor U151 (N_151,N_89,In_252);
nand U152 (N_152,N_105,In_96);
or U153 (N_153,N_101,N_58);
nor U154 (N_154,In_478,N_87);
nor U155 (N_155,N_96,N_98);
and U156 (N_156,In_363,In_72);
and U157 (N_157,In_130,In_127);
or U158 (N_158,N_37,In_458);
nor U159 (N_159,In_336,In_434);
nand U160 (N_160,N_78,In_284);
nor U161 (N_161,N_63,In_207);
nand U162 (N_162,N_27,N_82);
nand U163 (N_163,N_75,In_133);
or U164 (N_164,In_118,N_43);
nor U165 (N_165,N_116,In_494);
and U166 (N_166,In_488,In_482);
nor U167 (N_167,N_24,In_146);
or U168 (N_168,N_88,In_84);
nor U169 (N_169,N_56,In_234);
nor U170 (N_170,In_347,N_65);
or U171 (N_171,In_387,In_50);
nand U172 (N_172,In_431,N_119);
nor U173 (N_173,In_403,In_323);
and U174 (N_174,In_44,In_418);
or U175 (N_175,In_470,In_490);
nand U176 (N_176,In_483,In_69);
nor U177 (N_177,In_85,In_263);
and U178 (N_178,In_193,In_285);
nor U179 (N_179,In_324,In_205);
nand U180 (N_180,N_52,N_168);
nand U181 (N_181,N_69,N_42);
and U182 (N_182,In_70,In_173);
nand U183 (N_183,In_330,N_173);
nor U184 (N_184,N_80,In_352);
and U185 (N_185,In_93,In_35);
or U186 (N_186,In_388,In_412);
xnor U187 (N_187,N_133,In_141);
nand U188 (N_188,N_154,In_14);
nor U189 (N_189,N_54,In_413);
nor U190 (N_190,N_45,N_51);
nand U191 (N_191,In_425,In_293);
and U192 (N_192,In_120,N_0);
nand U193 (N_193,In_149,In_27);
and U194 (N_194,In_2,In_202);
and U195 (N_195,In_24,In_464);
or U196 (N_196,In_393,N_143);
nand U197 (N_197,In_43,N_131);
nor U198 (N_198,N_70,N_159);
and U199 (N_199,In_109,N_9);
and U200 (N_200,In_217,In_206);
nand U201 (N_201,N_83,N_31);
nand U202 (N_202,N_111,N_155);
nand U203 (N_203,In_428,N_91);
and U204 (N_204,In_381,N_108);
nor U205 (N_205,N_134,In_136);
nand U206 (N_206,In_439,In_259);
nor U207 (N_207,In_445,In_486);
nand U208 (N_208,In_115,In_364);
nor U209 (N_209,N_68,In_110);
nand U210 (N_210,In_208,N_126);
nor U211 (N_211,N_72,N_64);
or U212 (N_212,N_95,In_469);
nand U213 (N_213,N_171,In_92);
and U214 (N_214,N_12,In_94);
and U215 (N_215,N_147,In_19);
nor U216 (N_216,In_159,In_170);
or U217 (N_217,In_320,In_315);
and U218 (N_218,In_344,In_88);
nor U219 (N_219,N_76,In_276);
nor U220 (N_220,N_29,In_135);
nor U221 (N_221,In_441,In_186);
and U222 (N_222,N_49,In_199);
and U223 (N_223,N_34,N_74);
nor U224 (N_224,In_212,In_184);
nor U225 (N_225,N_85,In_496);
and U226 (N_226,N_114,N_156);
nor U227 (N_227,In_39,In_461);
and U228 (N_228,In_355,In_466);
nand U229 (N_229,In_299,N_117);
and U230 (N_230,In_124,In_298);
or U231 (N_231,N_67,In_390);
nor U232 (N_232,N_92,In_309);
nand U233 (N_233,N_135,N_138);
nand U234 (N_234,N_136,N_127);
or U235 (N_235,In_451,In_296);
and U236 (N_236,In_89,In_400);
or U237 (N_237,N_77,In_419);
nor U238 (N_238,N_36,In_117);
nand U239 (N_239,In_333,N_161);
nor U240 (N_240,N_129,N_112);
or U241 (N_241,N_97,In_481);
nor U242 (N_242,In_33,In_264);
nor U243 (N_243,In_327,N_190);
and U244 (N_244,In_455,N_1);
or U245 (N_245,N_186,In_422);
and U246 (N_246,In_353,N_194);
and U247 (N_247,N_232,In_306);
nor U248 (N_248,N_229,N_191);
and U249 (N_249,N_107,In_52);
nand U250 (N_250,N_104,In_231);
nor U251 (N_251,In_339,N_123);
or U252 (N_252,N_239,N_238);
nand U253 (N_253,In_456,In_435);
and U254 (N_254,N_233,N_66);
and U255 (N_255,N_142,In_491);
and U256 (N_256,N_163,N_124);
nor U257 (N_257,In_268,N_166);
xor U258 (N_258,In_371,N_188);
nand U259 (N_259,In_68,N_211);
nor U260 (N_260,N_17,N_61);
nor U261 (N_261,In_181,In_227);
and U262 (N_262,N_181,N_140);
nand U263 (N_263,In_225,In_421);
and U264 (N_264,N_153,N_174);
nand U265 (N_265,In_321,In_100);
nand U266 (N_266,N_208,In_279);
and U267 (N_267,N_20,In_129);
and U268 (N_268,In_485,N_120);
or U269 (N_269,N_53,In_90);
nand U270 (N_270,N_35,In_155);
and U271 (N_271,In_444,N_196);
and U272 (N_272,In_246,N_152);
nor U273 (N_273,N_224,N_73);
and U274 (N_274,In_10,In_60);
nor U275 (N_275,N_182,N_218);
nor U276 (N_276,In_463,In_0);
and U277 (N_277,N_50,N_183);
or U278 (N_278,N_118,In_188);
or U279 (N_279,N_209,N_160);
nor U280 (N_280,N_10,N_179);
nand U281 (N_281,In_4,N_125);
nand U282 (N_282,N_164,N_214);
or U283 (N_283,N_150,In_218);
nand U284 (N_284,In_209,N_99);
and U285 (N_285,In_3,N_187);
and U286 (N_286,In_362,N_81);
and U287 (N_287,N_172,In_366);
nor U288 (N_288,In_157,In_256);
nand U289 (N_289,N_121,In_436);
or U290 (N_290,N_16,N_115);
and U291 (N_291,In_25,N_234);
and U292 (N_292,N_151,N_46);
nor U293 (N_293,N_165,N_177);
or U294 (N_294,N_205,N_216);
or U295 (N_295,N_149,N_32);
and U296 (N_296,In_423,In_111);
or U297 (N_297,N_228,N_2);
or U298 (N_298,In_128,N_169);
nor U299 (N_299,N_55,In_448);
xor U300 (N_300,N_3,In_216);
or U301 (N_301,N_268,In_452);
and U302 (N_302,N_202,N_180);
nand U303 (N_303,In_66,N_285);
and U304 (N_304,N_245,N_237);
nand U305 (N_305,In_229,N_15);
nor U306 (N_306,In_457,N_261);
or U307 (N_307,N_130,N_265);
nor U308 (N_308,In_450,In_158);
nand U309 (N_309,In_340,N_215);
or U310 (N_310,N_289,In_257);
nand U311 (N_311,N_246,N_297);
and U312 (N_312,N_201,N_219);
nor U313 (N_313,N_137,N_276);
and U314 (N_314,In_114,N_270);
or U315 (N_315,N_220,N_242);
and U316 (N_316,N_84,N_93);
and U317 (N_317,In_204,N_110);
nand U318 (N_318,N_287,In_105);
nand U319 (N_319,N_221,N_263);
or U320 (N_320,N_212,N_189);
nor U321 (N_321,In_311,N_243);
nor U322 (N_322,N_248,N_195);
nand U323 (N_323,N_146,In_454);
and U324 (N_324,In_443,N_185);
or U325 (N_325,N_200,N_39);
and U326 (N_326,In_350,N_199);
or U327 (N_327,N_176,N_278);
and U328 (N_328,In_95,N_178);
and U329 (N_329,N_167,N_250);
nand U330 (N_330,N_252,N_257);
nand U331 (N_331,N_282,In_192);
nand U332 (N_332,N_44,N_292);
or U333 (N_333,N_266,In_87);
and U334 (N_334,N_264,N_296);
or U335 (N_335,In_15,N_192);
and U336 (N_336,N_277,N_184);
nand U337 (N_337,In_104,N_213);
nor U338 (N_338,In_58,In_382);
or U339 (N_339,In_468,In_236);
nor U340 (N_340,In_398,N_197);
and U341 (N_341,N_122,N_79);
nand U342 (N_342,N_60,In_1);
nand U343 (N_343,N_298,N_90);
nor U344 (N_344,N_62,In_22);
nand U345 (N_345,In_220,N_144);
nand U346 (N_346,N_175,N_256);
and U347 (N_347,N_40,N_269);
or U348 (N_348,N_226,In_62);
nand U349 (N_349,In_367,N_193);
nand U350 (N_350,In_18,N_249);
or U351 (N_351,N_94,In_270);
nor U352 (N_352,N_294,In_379);
and U353 (N_353,In_356,N_253);
nor U354 (N_354,N_128,N_262);
or U355 (N_355,In_34,N_141);
or U356 (N_356,In_303,N_299);
nand U357 (N_357,N_28,In_440);
nand U358 (N_358,N_223,In_210);
nand U359 (N_359,N_288,In_437);
and U360 (N_360,N_206,N_258);
nor U361 (N_361,N_251,In_392);
nand U362 (N_362,N_328,N_309);
and U363 (N_363,N_260,In_240);
and U364 (N_364,N_313,N_350);
or U365 (N_365,N_332,In_429);
and U366 (N_366,In_442,N_322);
or U367 (N_367,N_356,N_302);
nand U368 (N_368,N_300,N_343);
and U369 (N_369,In_98,N_7);
or U370 (N_370,N_305,N_325);
or U371 (N_371,N_345,N_279);
nor U372 (N_372,N_217,N_316);
nor U373 (N_373,N_33,N_329);
and U374 (N_374,N_306,N_311);
and U375 (N_375,N_308,N_330);
nand U376 (N_376,In_172,N_272);
or U377 (N_377,N_335,N_319);
and U378 (N_378,N_315,N_327);
or U379 (N_379,In_152,N_240);
nand U380 (N_380,N_337,N_326);
nor U381 (N_381,N_303,N_244);
and U382 (N_382,N_210,In_391);
and U383 (N_383,In_187,N_230);
nand U384 (N_384,N_162,In_76);
and U385 (N_385,N_102,N_352);
and U386 (N_386,N_247,N_357);
or U387 (N_387,N_342,In_168);
nor U388 (N_388,In_479,In_289);
and U389 (N_389,N_286,N_222);
or U390 (N_390,N_290,N_139);
and U391 (N_391,N_336,N_148);
nand U392 (N_392,N_273,N_301);
and U393 (N_393,N_231,N_359);
or U394 (N_394,N_338,N_320);
and U395 (N_395,N_307,N_132);
or U396 (N_396,N_254,N_281);
or U397 (N_397,N_198,N_358);
nor U398 (N_398,N_293,In_12);
and U399 (N_399,N_236,N_347);
or U400 (N_400,N_324,N_318);
nor U401 (N_401,In_235,N_348);
nand U402 (N_402,N_334,N_321);
nor U403 (N_403,N_158,In_307);
nand U404 (N_404,N_341,In_271);
and U405 (N_405,N_351,N_170);
and U406 (N_406,N_227,N_204);
and U407 (N_407,N_314,N_304);
xor U408 (N_408,N_340,In_154);
nor U409 (N_409,In_278,N_312);
nor U410 (N_410,N_295,N_267);
or U411 (N_411,N_57,N_333);
or U412 (N_412,N_274,In_337);
or U413 (N_413,N_344,N_109);
nand U414 (N_414,In_290,N_225);
or U415 (N_415,N_310,In_151);
and U416 (N_416,N_317,N_353);
nor U417 (N_417,In_453,N_157);
or U418 (N_418,N_207,N_259);
nand U419 (N_419,N_145,N_323);
nor U420 (N_420,N_389,N_235);
or U421 (N_421,N_376,N_386);
or U422 (N_422,N_393,N_416);
nor U423 (N_423,N_417,N_384);
and U424 (N_424,N_404,N_283);
nor U425 (N_425,N_394,N_365);
nand U426 (N_426,N_391,N_379);
or U427 (N_427,N_371,N_407);
nand U428 (N_428,N_370,N_410);
or U429 (N_429,N_374,N_398);
and U430 (N_430,N_361,N_399);
or U431 (N_431,N_395,N_400);
nand U432 (N_432,N_280,N_381);
nand U433 (N_433,N_364,N_405);
or U434 (N_434,N_382,N_406);
and U435 (N_435,N_255,N_402);
nand U436 (N_436,N_414,N_373);
nor U437 (N_437,N_367,N_203);
nor U438 (N_438,N_380,N_354);
or U439 (N_439,N_378,N_363);
and U440 (N_440,N_418,N_86);
and U441 (N_441,N_360,N_409);
nor U442 (N_442,N_366,N_291);
nor U443 (N_443,N_419,N_396);
nand U444 (N_444,N_349,N_401);
or U445 (N_445,N_403,N_397);
or U446 (N_446,In_305,N_346);
or U447 (N_447,N_383,In_474);
nand U448 (N_448,N_415,N_375);
nand U449 (N_449,N_275,N_411);
or U450 (N_450,N_377,N_413);
or U451 (N_451,N_369,N_284);
nor U452 (N_452,N_408,N_388);
nor U453 (N_453,N_387,In_224);
nand U454 (N_454,N_368,N_331);
and U455 (N_455,N_390,N_372);
and U456 (N_456,N_412,N_362);
nor U457 (N_457,N_385,N_355);
or U458 (N_458,N_339,N_241);
or U459 (N_459,N_392,N_271);
and U460 (N_460,N_86,N_393);
nand U461 (N_461,N_403,N_346);
and U462 (N_462,N_271,N_407);
nor U463 (N_463,N_375,N_275);
and U464 (N_464,N_241,N_392);
nor U465 (N_465,N_373,N_388);
and U466 (N_466,N_400,N_361);
and U467 (N_467,N_397,N_354);
nor U468 (N_468,N_413,N_418);
nor U469 (N_469,N_381,N_390);
or U470 (N_470,N_331,N_406);
xnor U471 (N_471,N_383,N_403);
and U472 (N_472,N_387,N_275);
nand U473 (N_473,N_404,N_410);
nand U474 (N_474,N_381,N_283);
and U475 (N_475,N_406,N_413);
nand U476 (N_476,N_367,N_366);
or U477 (N_477,N_380,N_402);
and U478 (N_478,N_284,N_372);
nand U479 (N_479,N_414,N_366);
or U480 (N_480,N_463,N_432);
or U481 (N_481,N_428,N_451);
or U482 (N_482,N_476,N_475);
or U483 (N_483,N_450,N_420);
nor U484 (N_484,N_453,N_436);
nand U485 (N_485,N_431,N_429);
and U486 (N_486,N_470,N_460);
and U487 (N_487,N_433,N_430);
nor U488 (N_488,N_454,N_438);
and U489 (N_489,N_465,N_469);
nand U490 (N_490,N_448,N_427);
nor U491 (N_491,N_447,N_442);
and U492 (N_492,N_461,N_449);
or U493 (N_493,N_435,N_473);
nand U494 (N_494,N_467,N_439);
and U495 (N_495,N_437,N_452);
and U496 (N_496,N_423,N_446);
or U497 (N_497,N_458,N_472);
or U498 (N_498,N_424,N_459);
nand U499 (N_499,N_462,N_464);
and U500 (N_500,N_440,N_444);
and U501 (N_501,N_425,N_445);
and U502 (N_502,N_457,N_422);
nand U503 (N_503,N_455,N_441);
nand U504 (N_504,N_477,N_471);
nand U505 (N_505,N_456,N_421);
or U506 (N_506,N_443,N_474);
or U507 (N_507,N_426,N_466);
nand U508 (N_508,N_479,N_478);
xnor U509 (N_509,N_468,N_434);
nor U510 (N_510,N_478,N_462);
or U511 (N_511,N_427,N_456);
nand U512 (N_512,N_430,N_450);
or U513 (N_513,N_434,N_432);
or U514 (N_514,N_444,N_468);
or U515 (N_515,N_435,N_447);
and U516 (N_516,N_478,N_476);
nand U517 (N_517,N_458,N_439);
or U518 (N_518,N_473,N_470);
and U519 (N_519,N_449,N_474);
and U520 (N_520,N_437,N_476);
nand U521 (N_521,N_448,N_422);
nor U522 (N_522,N_448,N_438);
or U523 (N_523,N_472,N_427);
and U524 (N_524,N_462,N_430);
or U525 (N_525,N_443,N_423);
nor U526 (N_526,N_450,N_461);
and U527 (N_527,N_461,N_437);
nand U528 (N_528,N_461,N_475);
nor U529 (N_529,N_464,N_447);
or U530 (N_530,N_459,N_478);
or U531 (N_531,N_476,N_435);
and U532 (N_532,N_423,N_477);
nand U533 (N_533,N_464,N_424);
nand U534 (N_534,N_431,N_423);
or U535 (N_535,N_452,N_438);
and U536 (N_536,N_430,N_424);
nand U537 (N_537,N_467,N_442);
nor U538 (N_538,N_467,N_475);
nand U539 (N_539,N_453,N_435);
or U540 (N_540,N_491,N_537);
nor U541 (N_541,N_517,N_502);
nor U542 (N_542,N_527,N_531);
or U543 (N_543,N_503,N_481);
and U544 (N_544,N_499,N_498);
nor U545 (N_545,N_497,N_492);
nand U546 (N_546,N_509,N_538);
nand U547 (N_547,N_489,N_501);
or U548 (N_548,N_528,N_512);
nand U549 (N_549,N_513,N_530);
or U550 (N_550,N_533,N_496);
nor U551 (N_551,N_488,N_526);
or U552 (N_552,N_523,N_508);
or U553 (N_553,N_516,N_511);
or U554 (N_554,N_505,N_520);
nand U555 (N_555,N_486,N_506);
nand U556 (N_556,N_487,N_500);
nor U557 (N_557,N_518,N_494);
nor U558 (N_558,N_532,N_535);
nand U559 (N_559,N_519,N_521);
nor U560 (N_560,N_515,N_490);
nor U561 (N_561,N_493,N_525);
nor U562 (N_562,N_539,N_522);
or U563 (N_563,N_480,N_507);
and U564 (N_564,N_482,N_504);
or U565 (N_565,N_485,N_514);
nand U566 (N_566,N_495,N_536);
nor U567 (N_567,N_529,N_484);
and U568 (N_568,N_483,N_524);
and U569 (N_569,N_534,N_510);
nand U570 (N_570,N_504,N_512);
and U571 (N_571,N_511,N_505);
nor U572 (N_572,N_534,N_524);
and U573 (N_573,N_518,N_527);
nor U574 (N_574,N_510,N_526);
nor U575 (N_575,N_484,N_524);
or U576 (N_576,N_482,N_488);
xor U577 (N_577,N_519,N_492);
and U578 (N_578,N_511,N_484);
nand U579 (N_579,N_527,N_492);
nand U580 (N_580,N_536,N_493);
or U581 (N_581,N_500,N_538);
nand U582 (N_582,N_533,N_503);
or U583 (N_583,N_528,N_503);
nor U584 (N_584,N_510,N_523);
nand U585 (N_585,N_484,N_521);
nor U586 (N_586,N_499,N_508);
nor U587 (N_587,N_498,N_507);
and U588 (N_588,N_498,N_529);
nor U589 (N_589,N_524,N_533);
and U590 (N_590,N_526,N_507);
nand U591 (N_591,N_519,N_493);
or U592 (N_592,N_504,N_527);
or U593 (N_593,N_513,N_518);
and U594 (N_594,N_509,N_488);
nor U595 (N_595,N_518,N_490);
and U596 (N_596,N_533,N_525);
nor U597 (N_597,N_512,N_518);
nand U598 (N_598,N_515,N_536);
and U599 (N_599,N_512,N_486);
nand U600 (N_600,N_556,N_593);
nor U601 (N_601,N_589,N_576);
nor U602 (N_602,N_586,N_561);
or U603 (N_603,N_559,N_545);
nand U604 (N_604,N_553,N_579);
nand U605 (N_605,N_568,N_547);
or U606 (N_606,N_558,N_570);
nor U607 (N_607,N_582,N_573);
xor U608 (N_608,N_581,N_584);
nand U609 (N_609,N_599,N_566);
nand U610 (N_610,N_563,N_587);
or U611 (N_611,N_574,N_596);
nand U612 (N_612,N_544,N_564);
nand U613 (N_613,N_549,N_540);
nor U614 (N_614,N_548,N_571);
xor U615 (N_615,N_552,N_591);
nor U616 (N_616,N_578,N_575);
and U617 (N_617,N_557,N_551);
nand U618 (N_618,N_543,N_542);
nand U619 (N_619,N_594,N_595);
nand U620 (N_620,N_580,N_541);
or U621 (N_621,N_590,N_569);
and U622 (N_622,N_577,N_588);
xnor U623 (N_623,N_572,N_560);
or U624 (N_624,N_585,N_592);
and U625 (N_625,N_554,N_565);
nand U626 (N_626,N_555,N_562);
nand U627 (N_627,N_598,N_597);
nand U628 (N_628,N_567,N_550);
nor U629 (N_629,N_546,N_583);
nand U630 (N_630,N_577,N_573);
nor U631 (N_631,N_560,N_566);
or U632 (N_632,N_561,N_570);
and U633 (N_633,N_542,N_555);
or U634 (N_634,N_559,N_554);
and U635 (N_635,N_563,N_547);
and U636 (N_636,N_544,N_540);
nand U637 (N_637,N_571,N_594);
and U638 (N_638,N_547,N_589);
or U639 (N_639,N_562,N_546);
xnor U640 (N_640,N_541,N_550);
and U641 (N_641,N_597,N_565);
nor U642 (N_642,N_561,N_559);
nor U643 (N_643,N_548,N_546);
or U644 (N_644,N_596,N_570);
nand U645 (N_645,N_586,N_599);
or U646 (N_646,N_544,N_585);
and U647 (N_647,N_540,N_562);
or U648 (N_648,N_581,N_577);
or U649 (N_649,N_553,N_581);
or U650 (N_650,N_564,N_594);
nand U651 (N_651,N_595,N_566);
and U652 (N_652,N_595,N_584);
nand U653 (N_653,N_563,N_596);
and U654 (N_654,N_595,N_571);
nor U655 (N_655,N_572,N_593);
nand U656 (N_656,N_559,N_593);
nand U657 (N_657,N_543,N_598);
nor U658 (N_658,N_541,N_540);
xor U659 (N_659,N_598,N_592);
or U660 (N_660,N_651,N_603);
and U661 (N_661,N_647,N_655);
nand U662 (N_662,N_640,N_626);
or U663 (N_663,N_659,N_622);
and U664 (N_664,N_652,N_625);
and U665 (N_665,N_648,N_620);
nor U666 (N_666,N_631,N_657);
and U667 (N_667,N_614,N_646);
nand U668 (N_668,N_656,N_612);
or U669 (N_669,N_632,N_600);
nand U670 (N_670,N_630,N_639);
nor U671 (N_671,N_615,N_607);
or U672 (N_672,N_619,N_623);
nand U673 (N_673,N_610,N_650);
nand U674 (N_674,N_605,N_621);
or U675 (N_675,N_604,N_636);
nand U676 (N_676,N_653,N_654);
nand U677 (N_677,N_609,N_645);
or U678 (N_678,N_627,N_633);
nor U679 (N_679,N_618,N_616);
or U680 (N_680,N_617,N_635);
nor U681 (N_681,N_601,N_643);
and U682 (N_682,N_637,N_642);
or U683 (N_683,N_634,N_649);
and U684 (N_684,N_629,N_611);
or U685 (N_685,N_613,N_602);
nor U686 (N_686,N_641,N_624);
nand U687 (N_687,N_608,N_658);
nand U688 (N_688,N_644,N_638);
nor U689 (N_689,N_606,N_628);
or U690 (N_690,N_600,N_650);
and U691 (N_691,N_643,N_630);
and U692 (N_692,N_655,N_600);
and U693 (N_693,N_644,N_645);
nand U694 (N_694,N_655,N_653);
nand U695 (N_695,N_643,N_602);
nor U696 (N_696,N_605,N_600);
nand U697 (N_697,N_640,N_651);
and U698 (N_698,N_644,N_602);
nor U699 (N_699,N_627,N_617);
and U700 (N_700,N_652,N_642);
nand U701 (N_701,N_627,N_650);
xor U702 (N_702,N_615,N_630);
nor U703 (N_703,N_612,N_623);
or U704 (N_704,N_657,N_609);
nor U705 (N_705,N_620,N_655);
or U706 (N_706,N_635,N_629);
and U707 (N_707,N_638,N_613);
nand U708 (N_708,N_638,N_653);
nor U709 (N_709,N_611,N_658);
nand U710 (N_710,N_623,N_631);
and U711 (N_711,N_617,N_620);
nand U712 (N_712,N_650,N_656);
nor U713 (N_713,N_626,N_655);
nand U714 (N_714,N_648,N_607);
and U715 (N_715,N_638,N_609);
nand U716 (N_716,N_607,N_632);
and U717 (N_717,N_613,N_610);
nand U718 (N_718,N_659,N_655);
nor U719 (N_719,N_635,N_639);
nand U720 (N_720,N_688,N_694);
nand U721 (N_721,N_681,N_698);
and U722 (N_722,N_670,N_713);
nand U723 (N_723,N_679,N_705);
and U724 (N_724,N_704,N_707);
or U725 (N_725,N_682,N_697);
or U726 (N_726,N_717,N_684);
nand U727 (N_727,N_677,N_667);
or U728 (N_728,N_689,N_716);
or U729 (N_729,N_701,N_691);
nor U730 (N_730,N_685,N_663);
and U731 (N_731,N_683,N_674);
nor U732 (N_732,N_675,N_666);
nand U733 (N_733,N_664,N_695);
or U734 (N_734,N_706,N_661);
nor U735 (N_735,N_668,N_709);
and U736 (N_736,N_718,N_714);
and U737 (N_737,N_665,N_687);
nor U738 (N_738,N_662,N_690);
nor U739 (N_739,N_715,N_711);
nor U740 (N_740,N_686,N_660);
or U741 (N_741,N_702,N_693);
and U742 (N_742,N_680,N_700);
or U743 (N_743,N_672,N_671);
nand U744 (N_744,N_673,N_699);
and U745 (N_745,N_719,N_676);
or U746 (N_746,N_696,N_708);
or U747 (N_747,N_692,N_678);
or U748 (N_748,N_712,N_710);
nor U749 (N_749,N_669,N_703);
xor U750 (N_750,N_696,N_669);
or U751 (N_751,N_673,N_678);
nor U752 (N_752,N_705,N_660);
or U753 (N_753,N_701,N_677);
nor U754 (N_754,N_685,N_678);
and U755 (N_755,N_691,N_674);
nand U756 (N_756,N_677,N_717);
nor U757 (N_757,N_698,N_690);
or U758 (N_758,N_666,N_682);
and U759 (N_759,N_689,N_710);
nand U760 (N_760,N_686,N_661);
or U761 (N_761,N_712,N_717);
nor U762 (N_762,N_671,N_689);
and U763 (N_763,N_700,N_675);
nor U764 (N_764,N_713,N_705);
nor U765 (N_765,N_713,N_679);
nand U766 (N_766,N_671,N_682);
nor U767 (N_767,N_676,N_672);
or U768 (N_768,N_670,N_673);
nor U769 (N_769,N_690,N_696);
and U770 (N_770,N_716,N_700);
and U771 (N_771,N_674,N_676);
nor U772 (N_772,N_693,N_719);
or U773 (N_773,N_676,N_693);
and U774 (N_774,N_719,N_667);
and U775 (N_775,N_677,N_719);
nor U776 (N_776,N_703,N_718);
or U777 (N_777,N_662,N_702);
nand U778 (N_778,N_671,N_690);
or U779 (N_779,N_666,N_673);
nand U780 (N_780,N_736,N_721);
or U781 (N_781,N_737,N_777);
and U782 (N_782,N_768,N_742);
nand U783 (N_783,N_740,N_741);
nor U784 (N_784,N_772,N_756);
nand U785 (N_785,N_774,N_751);
nand U786 (N_786,N_750,N_730);
or U787 (N_787,N_763,N_753);
nand U788 (N_788,N_727,N_738);
or U789 (N_789,N_765,N_720);
nor U790 (N_790,N_739,N_749);
nand U791 (N_791,N_747,N_755);
and U792 (N_792,N_752,N_758);
nand U793 (N_793,N_762,N_748);
or U794 (N_794,N_776,N_732);
nor U795 (N_795,N_729,N_743);
and U796 (N_796,N_754,N_767);
nand U797 (N_797,N_779,N_746);
and U798 (N_798,N_775,N_735);
xnor U799 (N_799,N_759,N_766);
nand U800 (N_800,N_723,N_760);
nor U801 (N_801,N_734,N_761);
or U802 (N_802,N_770,N_773);
or U803 (N_803,N_722,N_764);
nand U804 (N_804,N_771,N_726);
or U805 (N_805,N_744,N_745);
or U806 (N_806,N_733,N_728);
or U807 (N_807,N_757,N_724);
and U808 (N_808,N_725,N_778);
or U809 (N_809,N_769,N_731);
nor U810 (N_810,N_731,N_746);
or U811 (N_811,N_770,N_777);
and U812 (N_812,N_759,N_731);
nand U813 (N_813,N_729,N_766);
and U814 (N_814,N_731,N_776);
nand U815 (N_815,N_748,N_775);
or U816 (N_816,N_739,N_745);
or U817 (N_817,N_728,N_754);
and U818 (N_818,N_726,N_739);
and U819 (N_819,N_751,N_740);
nand U820 (N_820,N_771,N_762);
nand U821 (N_821,N_743,N_755);
or U822 (N_822,N_724,N_763);
nand U823 (N_823,N_724,N_734);
and U824 (N_824,N_739,N_757);
nand U825 (N_825,N_745,N_761);
or U826 (N_826,N_751,N_725);
and U827 (N_827,N_767,N_771);
nor U828 (N_828,N_730,N_777);
or U829 (N_829,N_732,N_762);
or U830 (N_830,N_724,N_762);
nand U831 (N_831,N_745,N_763);
nor U832 (N_832,N_776,N_756);
nand U833 (N_833,N_774,N_720);
nor U834 (N_834,N_757,N_765);
nand U835 (N_835,N_750,N_726);
and U836 (N_836,N_748,N_758);
nor U837 (N_837,N_740,N_752);
and U838 (N_838,N_761,N_748);
nand U839 (N_839,N_754,N_755);
nor U840 (N_840,N_809,N_808);
nor U841 (N_841,N_805,N_788);
nor U842 (N_842,N_833,N_829);
nand U843 (N_843,N_795,N_837);
or U844 (N_844,N_781,N_835);
nor U845 (N_845,N_815,N_785);
nand U846 (N_846,N_819,N_783);
xnor U847 (N_847,N_828,N_780);
or U848 (N_848,N_798,N_822);
and U849 (N_849,N_791,N_816);
or U850 (N_850,N_824,N_839);
and U851 (N_851,N_813,N_789);
or U852 (N_852,N_818,N_817);
or U853 (N_853,N_793,N_811);
and U854 (N_854,N_801,N_830);
nor U855 (N_855,N_836,N_806);
and U856 (N_856,N_832,N_810);
nand U857 (N_857,N_807,N_787);
and U858 (N_858,N_814,N_786);
nor U859 (N_859,N_796,N_804);
and U860 (N_860,N_797,N_799);
nand U861 (N_861,N_838,N_812);
and U862 (N_862,N_825,N_826);
nand U863 (N_863,N_827,N_800);
nor U864 (N_864,N_790,N_823);
or U865 (N_865,N_782,N_821);
or U866 (N_866,N_803,N_831);
nand U867 (N_867,N_820,N_784);
nand U868 (N_868,N_794,N_802);
nand U869 (N_869,N_834,N_792);
or U870 (N_870,N_800,N_789);
and U871 (N_871,N_821,N_803);
or U872 (N_872,N_827,N_820);
or U873 (N_873,N_829,N_810);
or U874 (N_874,N_790,N_819);
or U875 (N_875,N_813,N_802);
or U876 (N_876,N_799,N_805);
nor U877 (N_877,N_793,N_819);
and U878 (N_878,N_827,N_804);
nand U879 (N_879,N_785,N_790);
nor U880 (N_880,N_785,N_793);
or U881 (N_881,N_808,N_826);
and U882 (N_882,N_826,N_783);
and U883 (N_883,N_809,N_797);
or U884 (N_884,N_826,N_819);
nand U885 (N_885,N_822,N_825);
nor U886 (N_886,N_823,N_802);
and U887 (N_887,N_784,N_838);
and U888 (N_888,N_788,N_792);
and U889 (N_889,N_827,N_793);
nor U890 (N_890,N_788,N_804);
nand U891 (N_891,N_800,N_819);
nor U892 (N_892,N_797,N_834);
or U893 (N_893,N_801,N_785);
nand U894 (N_894,N_824,N_831);
or U895 (N_895,N_807,N_825);
or U896 (N_896,N_819,N_787);
nor U897 (N_897,N_809,N_831);
or U898 (N_898,N_794,N_812);
nand U899 (N_899,N_821,N_796);
nor U900 (N_900,N_867,N_863);
nor U901 (N_901,N_895,N_872);
or U902 (N_902,N_880,N_852);
nand U903 (N_903,N_876,N_892);
or U904 (N_904,N_877,N_888);
and U905 (N_905,N_846,N_843);
nand U906 (N_906,N_854,N_859);
nor U907 (N_907,N_844,N_871);
and U908 (N_908,N_890,N_894);
and U909 (N_909,N_885,N_873);
or U910 (N_910,N_879,N_897);
and U911 (N_911,N_891,N_878);
or U912 (N_912,N_841,N_865);
and U913 (N_913,N_881,N_847);
and U914 (N_914,N_862,N_850);
or U915 (N_915,N_855,N_858);
nand U916 (N_916,N_840,N_857);
and U917 (N_917,N_860,N_886);
and U918 (N_918,N_883,N_842);
and U919 (N_919,N_849,N_853);
nand U920 (N_920,N_870,N_864);
and U921 (N_921,N_893,N_889);
or U922 (N_922,N_884,N_882);
nand U923 (N_923,N_845,N_856);
and U924 (N_924,N_874,N_851);
nand U925 (N_925,N_887,N_899);
nand U926 (N_926,N_869,N_868);
or U927 (N_927,N_848,N_875);
or U928 (N_928,N_866,N_898);
or U929 (N_929,N_861,N_896);
nor U930 (N_930,N_849,N_845);
nand U931 (N_931,N_841,N_880);
nor U932 (N_932,N_868,N_867);
or U933 (N_933,N_894,N_867);
and U934 (N_934,N_869,N_853);
and U935 (N_935,N_895,N_847);
and U936 (N_936,N_883,N_895);
nand U937 (N_937,N_863,N_890);
nor U938 (N_938,N_841,N_850);
or U939 (N_939,N_862,N_844);
nor U940 (N_940,N_846,N_881);
or U941 (N_941,N_849,N_884);
and U942 (N_942,N_890,N_851);
or U943 (N_943,N_865,N_862);
or U944 (N_944,N_879,N_885);
or U945 (N_945,N_856,N_862);
and U946 (N_946,N_853,N_893);
and U947 (N_947,N_895,N_888);
and U948 (N_948,N_883,N_855);
nand U949 (N_949,N_874,N_848);
or U950 (N_950,N_880,N_875);
and U951 (N_951,N_854,N_895);
or U952 (N_952,N_894,N_882);
or U953 (N_953,N_851,N_850);
nor U954 (N_954,N_881,N_875);
and U955 (N_955,N_891,N_887);
and U956 (N_956,N_870,N_866);
nand U957 (N_957,N_888,N_884);
nor U958 (N_958,N_882,N_851);
and U959 (N_959,N_867,N_849);
or U960 (N_960,N_950,N_956);
and U961 (N_961,N_902,N_947);
nor U962 (N_962,N_919,N_953);
nand U963 (N_963,N_946,N_909);
and U964 (N_964,N_930,N_901);
nand U965 (N_965,N_914,N_932);
nor U966 (N_966,N_944,N_913);
nand U967 (N_967,N_943,N_942);
or U968 (N_968,N_908,N_905);
nand U969 (N_969,N_955,N_936);
nand U970 (N_970,N_958,N_952);
and U971 (N_971,N_949,N_940);
nor U972 (N_972,N_915,N_918);
or U973 (N_973,N_906,N_923);
or U974 (N_974,N_951,N_928);
nor U975 (N_975,N_938,N_912);
nor U976 (N_976,N_917,N_904);
or U977 (N_977,N_921,N_927);
nand U978 (N_978,N_925,N_924);
nor U979 (N_979,N_945,N_954);
or U980 (N_980,N_939,N_941);
nand U981 (N_981,N_931,N_926);
nor U982 (N_982,N_920,N_959);
or U983 (N_983,N_900,N_934);
and U984 (N_984,N_922,N_911);
and U985 (N_985,N_929,N_903);
and U986 (N_986,N_916,N_957);
nor U987 (N_987,N_910,N_948);
and U988 (N_988,N_937,N_933);
and U989 (N_989,N_935,N_907);
or U990 (N_990,N_953,N_922);
and U991 (N_991,N_904,N_928);
nor U992 (N_992,N_958,N_931);
and U993 (N_993,N_944,N_939);
and U994 (N_994,N_937,N_930);
nand U995 (N_995,N_946,N_921);
nor U996 (N_996,N_940,N_908);
and U997 (N_997,N_925,N_902);
nor U998 (N_998,N_917,N_918);
nor U999 (N_999,N_956,N_906);
nand U1000 (N_1000,N_939,N_910);
nor U1001 (N_1001,N_932,N_921);
nor U1002 (N_1002,N_919,N_927);
or U1003 (N_1003,N_904,N_953);
or U1004 (N_1004,N_920,N_904);
nand U1005 (N_1005,N_942,N_928);
or U1006 (N_1006,N_900,N_937);
nor U1007 (N_1007,N_936,N_911);
or U1008 (N_1008,N_919,N_914);
or U1009 (N_1009,N_915,N_910);
or U1010 (N_1010,N_951,N_943);
or U1011 (N_1011,N_943,N_922);
and U1012 (N_1012,N_907,N_900);
nor U1013 (N_1013,N_946,N_914);
or U1014 (N_1014,N_909,N_950);
and U1015 (N_1015,N_927,N_945);
nor U1016 (N_1016,N_933,N_940);
and U1017 (N_1017,N_951,N_929);
xor U1018 (N_1018,N_941,N_903);
nand U1019 (N_1019,N_958,N_942);
and U1020 (N_1020,N_975,N_980);
or U1021 (N_1021,N_977,N_986);
and U1022 (N_1022,N_981,N_1000);
nor U1023 (N_1023,N_973,N_964);
nand U1024 (N_1024,N_963,N_960);
or U1025 (N_1025,N_1007,N_982);
xor U1026 (N_1026,N_965,N_1018);
nand U1027 (N_1027,N_970,N_1011);
nor U1028 (N_1028,N_961,N_969);
and U1029 (N_1029,N_1014,N_990);
nand U1030 (N_1030,N_974,N_992);
nand U1031 (N_1031,N_1009,N_968);
or U1032 (N_1032,N_998,N_1019);
nand U1033 (N_1033,N_997,N_999);
nor U1034 (N_1034,N_995,N_967);
nor U1035 (N_1035,N_1013,N_1012);
or U1036 (N_1036,N_1017,N_962);
nor U1037 (N_1037,N_989,N_1006);
nor U1038 (N_1038,N_966,N_976);
nand U1039 (N_1039,N_1010,N_1005);
or U1040 (N_1040,N_972,N_988);
nand U1041 (N_1041,N_1004,N_1002);
nor U1042 (N_1042,N_971,N_993);
and U1043 (N_1043,N_1001,N_1003);
nand U1044 (N_1044,N_1015,N_987);
nand U1045 (N_1045,N_991,N_979);
nand U1046 (N_1046,N_996,N_1008);
nand U1047 (N_1047,N_978,N_984);
and U1048 (N_1048,N_994,N_985);
nor U1049 (N_1049,N_1016,N_983);
or U1050 (N_1050,N_1005,N_973);
nand U1051 (N_1051,N_963,N_989);
nor U1052 (N_1052,N_962,N_979);
or U1053 (N_1053,N_1018,N_994);
nand U1054 (N_1054,N_989,N_996);
nor U1055 (N_1055,N_972,N_997);
nor U1056 (N_1056,N_978,N_964);
nand U1057 (N_1057,N_983,N_974);
or U1058 (N_1058,N_993,N_970);
nor U1059 (N_1059,N_1009,N_995);
nand U1060 (N_1060,N_1002,N_1016);
nor U1061 (N_1061,N_994,N_1005);
nand U1062 (N_1062,N_981,N_975);
and U1063 (N_1063,N_981,N_1007);
nor U1064 (N_1064,N_996,N_973);
nor U1065 (N_1065,N_979,N_961);
or U1066 (N_1066,N_969,N_1017);
and U1067 (N_1067,N_989,N_1005);
or U1068 (N_1068,N_980,N_1000);
nor U1069 (N_1069,N_1002,N_1008);
and U1070 (N_1070,N_968,N_1013);
nand U1071 (N_1071,N_994,N_967);
and U1072 (N_1072,N_985,N_997);
nor U1073 (N_1073,N_1007,N_977);
nor U1074 (N_1074,N_999,N_998);
and U1075 (N_1075,N_979,N_1008);
or U1076 (N_1076,N_1014,N_1008);
or U1077 (N_1077,N_968,N_1010);
nand U1078 (N_1078,N_975,N_976);
nand U1079 (N_1079,N_1002,N_968);
and U1080 (N_1080,N_1049,N_1062);
or U1081 (N_1081,N_1051,N_1058);
nand U1082 (N_1082,N_1063,N_1036);
nand U1083 (N_1083,N_1056,N_1050);
nor U1084 (N_1084,N_1034,N_1047);
and U1085 (N_1085,N_1039,N_1038);
and U1086 (N_1086,N_1037,N_1064);
and U1087 (N_1087,N_1067,N_1076);
nor U1088 (N_1088,N_1065,N_1040);
xor U1089 (N_1089,N_1033,N_1055);
and U1090 (N_1090,N_1054,N_1070);
nand U1091 (N_1091,N_1079,N_1043);
nor U1092 (N_1092,N_1060,N_1045);
nand U1093 (N_1093,N_1030,N_1057);
and U1094 (N_1094,N_1072,N_1068);
nand U1095 (N_1095,N_1020,N_1042);
or U1096 (N_1096,N_1078,N_1061);
nand U1097 (N_1097,N_1023,N_1041);
or U1098 (N_1098,N_1071,N_1022);
nor U1099 (N_1099,N_1077,N_1075);
nor U1100 (N_1100,N_1035,N_1046);
nand U1101 (N_1101,N_1066,N_1032);
nor U1102 (N_1102,N_1021,N_1069);
xnor U1103 (N_1103,N_1073,N_1059);
nor U1104 (N_1104,N_1053,N_1074);
or U1105 (N_1105,N_1029,N_1024);
xor U1106 (N_1106,N_1052,N_1025);
and U1107 (N_1107,N_1044,N_1048);
nand U1108 (N_1108,N_1028,N_1027);
nor U1109 (N_1109,N_1026,N_1031);
and U1110 (N_1110,N_1038,N_1060);
nor U1111 (N_1111,N_1067,N_1035);
or U1112 (N_1112,N_1063,N_1046);
or U1113 (N_1113,N_1032,N_1033);
nand U1114 (N_1114,N_1071,N_1028);
and U1115 (N_1115,N_1045,N_1047);
xor U1116 (N_1116,N_1031,N_1064);
nor U1117 (N_1117,N_1073,N_1075);
and U1118 (N_1118,N_1020,N_1024);
nand U1119 (N_1119,N_1058,N_1045);
nand U1120 (N_1120,N_1036,N_1071);
nand U1121 (N_1121,N_1065,N_1070);
and U1122 (N_1122,N_1074,N_1065);
and U1123 (N_1123,N_1077,N_1076);
and U1124 (N_1124,N_1047,N_1060);
nand U1125 (N_1125,N_1066,N_1040);
or U1126 (N_1126,N_1077,N_1025);
or U1127 (N_1127,N_1059,N_1043);
nor U1128 (N_1128,N_1054,N_1040);
or U1129 (N_1129,N_1064,N_1063);
or U1130 (N_1130,N_1029,N_1076);
nand U1131 (N_1131,N_1025,N_1035);
and U1132 (N_1132,N_1072,N_1021);
and U1133 (N_1133,N_1045,N_1051);
nor U1134 (N_1134,N_1029,N_1045);
or U1135 (N_1135,N_1033,N_1063);
and U1136 (N_1136,N_1057,N_1036);
nor U1137 (N_1137,N_1075,N_1078);
and U1138 (N_1138,N_1052,N_1028);
nor U1139 (N_1139,N_1042,N_1038);
and U1140 (N_1140,N_1088,N_1099);
nor U1141 (N_1141,N_1108,N_1125);
nor U1142 (N_1142,N_1104,N_1119);
or U1143 (N_1143,N_1097,N_1084);
nand U1144 (N_1144,N_1138,N_1123);
or U1145 (N_1145,N_1131,N_1090);
or U1146 (N_1146,N_1130,N_1087);
and U1147 (N_1147,N_1118,N_1107);
or U1148 (N_1148,N_1112,N_1135);
nand U1149 (N_1149,N_1114,N_1082);
nor U1150 (N_1150,N_1120,N_1133);
and U1151 (N_1151,N_1106,N_1122);
nand U1152 (N_1152,N_1096,N_1129);
nand U1153 (N_1153,N_1136,N_1093);
nand U1154 (N_1154,N_1081,N_1117);
or U1155 (N_1155,N_1102,N_1086);
and U1156 (N_1156,N_1116,N_1137);
and U1157 (N_1157,N_1101,N_1139);
nor U1158 (N_1158,N_1113,N_1121);
nor U1159 (N_1159,N_1092,N_1105);
nand U1160 (N_1160,N_1132,N_1094);
nor U1161 (N_1161,N_1127,N_1115);
and U1162 (N_1162,N_1128,N_1110);
or U1163 (N_1163,N_1124,N_1080);
nor U1164 (N_1164,N_1100,N_1109);
and U1165 (N_1165,N_1091,N_1098);
and U1166 (N_1166,N_1103,N_1083);
nand U1167 (N_1167,N_1095,N_1111);
and U1168 (N_1168,N_1134,N_1089);
nand U1169 (N_1169,N_1085,N_1126);
nand U1170 (N_1170,N_1100,N_1113);
nor U1171 (N_1171,N_1114,N_1134);
or U1172 (N_1172,N_1130,N_1102);
nor U1173 (N_1173,N_1090,N_1110);
and U1174 (N_1174,N_1127,N_1134);
or U1175 (N_1175,N_1093,N_1122);
or U1176 (N_1176,N_1082,N_1096);
nor U1177 (N_1177,N_1092,N_1114);
or U1178 (N_1178,N_1095,N_1086);
or U1179 (N_1179,N_1081,N_1089);
or U1180 (N_1180,N_1108,N_1129);
and U1181 (N_1181,N_1098,N_1121);
nand U1182 (N_1182,N_1099,N_1118);
and U1183 (N_1183,N_1127,N_1083);
nand U1184 (N_1184,N_1108,N_1132);
and U1185 (N_1185,N_1106,N_1129);
nor U1186 (N_1186,N_1122,N_1118);
and U1187 (N_1187,N_1107,N_1138);
and U1188 (N_1188,N_1083,N_1114);
or U1189 (N_1189,N_1103,N_1107);
nor U1190 (N_1190,N_1087,N_1091);
or U1191 (N_1191,N_1103,N_1087);
nand U1192 (N_1192,N_1127,N_1137);
or U1193 (N_1193,N_1125,N_1119);
nand U1194 (N_1194,N_1133,N_1116);
nand U1195 (N_1195,N_1132,N_1101);
nor U1196 (N_1196,N_1134,N_1125);
nand U1197 (N_1197,N_1116,N_1101);
and U1198 (N_1198,N_1105,N_1087);
and U1199 (N_1199,N_1096,N_1089);
nor U1200 (N_1200,N_1190,N_1192);
or U1201 (N_1201,N_1193,N_1159);
or U1202 (N_1202,N_1189,N_1143);
and U1203 (N_1203,N_1173,N_1194);
xnor U1204 (N_1204,N_1170,N_1157);
or U1205 (N_1205,N_1153,N_1154);
nand U1206 (N_1206,N_1176,N_1184);
or U1207 (N_1207,N_1197,N_1145);
or U1208 (N_1208,N_1169,N_1147);
or U1209 (N_1209,N_1196,N_1186);
nor U1210 (N_1210,N_1140,N_1178);
or U1211 (N_1211,N_1172,N_1183);
and U1212 (N_1212,N_1162,N_1167);
or U1213 (N_1213,N_1151,N_1185);
nor U1214 (N_1214,N_1187,N_1195);
or U1215 (N_1215,N_1144,N_1148);
nor U1216 (N_1216,N_1155,N_1179);
and U1217 (N_1217,N_1171,N_1182);
or U1218 (N_1218,N_1174,N_1156);
and U1219 (N_1219,N_1141,N_1161);
nor U1220 (N_1220,N_1175,N_1166);
nor U1221 (N_1221,N_1177,N_1188);
and U1222 (N_1222,N_1199,N_1149);
nand U1223 (N_1223,N_1181,N_1152);
and U1224 (N_1224,N_1163,N_1146);
and U1225 (N_1225,N_1158,N_1160);
and U1226 (N_1226,N_1150,N_1142);
or U1227 (N_1227,N_1198,N_1165);
nor U1228 (N_1228,N_1180,N_1164);
nand U1229 (N_1229,N_1168,N_1191);
nand U1230 (N_1230,N_1186,N_1164);
or U1231 (N_1231,N_1164,N_1199);
or U1232 (N_1232,N_1194,N_1140);
nor U1233 (N_1233,N_1166,N_1156);
nand U1234 (N_1234,N_1143,N_1188);
nor U1235 (N_1235,N_1182,N_1160);
nand U1236 (N_1236,N_1189,N_1182);
and U1237 (N_1237,N_1196,N_1167);
nor U1238 (N_1238,N_1191,N_1199);
nand U1239 (N_1239,N_1147,N_1175);
nor U1240 (N_1240,N_1151,N_1161);
nor U1241 (N_1241,N_1170,N_1148);
or U1242 (N_1242,N_1166,N_1163);
nand U1243 (N_1243,N_1146,N_1153);
nor U1244 (N_1244,N_1143,N_1167);
and U1245 (N_1245,N_1170,N_1145);
or U1246 (N_1246,N_1177,N_1149);
nand U1247 (N_1247,N_1198,N_1153);
and U1248 (N_1248,N_1141,N_1143);
nor U1249 (N_1249,N_1141,N_1175);
and U1250 (N_1250,N_1182,N_1146);
nor U1251 (N_1251,N_1195,N_1169);
nor U1252 (N_1252,N_1146,N_1141);
or U1253 (N_1253,N_1158,N_1147);
and U1254 (N_1254,N_1172,N_1178);
nor U1255 (N_1255,N_1174,N_1187);
or U1256 (N_1256,N_1165,N_1196);
or U1257 (N_1257,N_1171,N_1173);
or U1258 (N_1258,N_1166,N_1185);
nor U1259 (N_1259,N_1142,N_1157);
nand U1260 (N_1260,N_1241,N_1228);
or U1261 (N_1261,N_1256,N_1224);
and U1262 (N_1262,N_1226,N_1258);
or U1263 (N_1263,N_1221,N_1211);
or U1264 (N_1264,N_1229,N_1208);
nand U1265 (N_1265,N_1203,N_1254);
or U1266 (N_1266,N_1235,N_1234);
nor U1267 (N_1267,N_1217,N_1248);
and U1268 (N_1268,N_1249,N_1257);
and U1269 (N_1269,N_1253,N_1218);
and U1270 (N_1270,N_1242,N_1232);
or U1271 (N_1271,N_1223,N_1246);
nand U1272 (N_1272,N_1205,N_1219);
nand U1273 (N_1273,N_1237,N_1239);
and U1274 (N_1274,N_1245,N_1210);
or U1275 (N_1275,N_1233,N_1230);
or U1276 (N_1276,N_1240,N_1227);
nor U1277 (N_1277,N_1259,N_1244);
and U1278 (N_1278,N_1251,N_1213);
nand U1279 (N_1279,N_1231,N_1250);
nor U1280 (N_1280,N_1236,N_1216);
nand U1281 (N_1281,N_1204,N_1214);
and U1282 (N_1282,N_1201,N_1225);
nand U1283 (N_1283,N_1255,N_1252);
and U1284 (N_1284,N_1215,N_1200);
nor U1285 (N_1285,N_1202,N_1212);
and U1286 (N_1286,N_1247,N_1206);
nand U1287 (N_1287,N_1209,N_1207);
and U1288 (N_1288,N_1243,N_1222);
nand U1289 (N_1289,N_1220,N_1238);
nand U1290 (N_1290,N_1259,N_1250);
or U1291 (N_1291,N_1219,N_1223);
nor U1292 (N_1292,N_1236,N_1218);
and U1293 (N_1293,N_1222,N_1227);
or U1294 (N_1294,N_1233,N_1208);
nor U1295 (N_1295,N_1243,N_1201);
nand U1296 (N_1296,N_1235,N_1253);
nor U1297 (N_1297,N_1251,N_1201);
nand U1298 (N_1298,N_1230,N_1223);
nand U1299 (N_1299,N_1215,N_1244);
and U1300 (N_1300,N_1226,N_1232);
nor U1301 (N_1301,N_1232,N_1250);
or U1302 (N_1302,N_1228,N_1231);
or U1303 (N_1303,N_1209,N_1256);
nor U1304 (N_1304,N_1202,N_1243);
or U1305 (N_1305,N_1217,N_1239);
nor U1306 (N_1306,N_1250,N_1210);
nor U1307 (N_1307,N_1224,N_1227);
or U1308 (N_1308,N_1255,N_1200);
or U1309 (N_1309,N_1208,N_1214);
nor U1310 (N_1310,N_1239,N_1248);
nor U1311 (N_1311,N_1238,N_1235);
and U1312 (N_1312,N_1216,N_1259);
or U1313 (N_1313,N_1252,N_1222);
or U1314 (N_1314,N_1235,N_1211);
or U1315 (N_1315,N_1249,N_1200);
nand U1316 (N_1316,N_1257,N_1209);
or U1317 (N_1317,N_1208,N_1249);
nor U1318 (N_1318,N_1248,N_1201);
nor U1319 (N_1319,N_1211,N_1244);
or U1320 (N_1320,N_1267,N_1263);
and U1321 (N_1321,N_1309,N_1292);
and U1322 (N_1322,N_1316,N_1279);
nor U1323 (N_1323,N_1284,N_1307);
nand U1324 (N_1324,N_1269,N_1278);
or U1325 (N_1325,N_1282,N_1264);
or U1326 (N_1326,N_1297,N_1312);
nand U1327 (N_1327,N_1305,N_1262);
nand U1328 (N_1328,N_1289,N_1287);
xnor U1329 (N_1329,N_1294,N_1265);
xor U1330 (N_1330,N_1293,N_1301);
nand U1331 (N_1331,N_1261,N_1296);
nor U1332 (N_1332,N_1286,N_1304);
and U1333 (N_1333,N_1319,N_1277);
or U1334 (N_1334,N_1313,N_1276);
and U1335 (N_1335,N_1299,N_1308);
or U1336 (N_1336,N_1280,N_1314);
or U1337 (N_1337,N_1273,N_1306);
and U1338 (N_1338,N_1271,N_1311);
nor U1339 (N_1339,N_1281,N_1290);
and U1340 (N_1340,N_1300,N_1274);
nor U1341 (N_1341,N_1288,N_1268);
and U1342 (N_1342,N_1298,N_1317);
nor U1343 (N_1343,N_1285,N_1315);
nor U1344 (N_1344,N_1318,N_1283);
or U1345 (N_1345,N_1272,N_1295);
or U1346 (N_1346,N_1302,N_1310);
nand U1347 (N_1347,N_1266,N_1270);
and U1348 (N_1348,N_1260,N_1303);
or U1349 (N_1349,N_1291,N_1275);
nand U1350 (N_1350,N_1262,N_1267);
or U1351 (N_1351,N_1307,N_1264);
or U1352 (N_1352,N_1314,N_1300);
xor U1353 (N_1353,N_1294,N_1312);
nor U1354 (N_1354,N_1263,N_1318);
or U1355 (N_1355,N_1274,N_1291);
and U1356 (N_1356,N_1275,N_1316);
or U1357 (N_1357,N_1293,N_1289);
nor U1358 (N_1358,N_1318,N_1269);
or U1359 (N_1359,N_1285,N_1264);
nor U1360 (N_1360,N_1309,N_1269);
or U1361 (N_1361,N_1282,N_1300);
xnor U1362 (N_1362,N_1279,N_1265);
nand U1363 (N_1363,N_1271,N_1316);
and U1364 (N_1364,N_1280,N_1274);
or U1365 (N_1365,N_1295,N_1300);
nand U1366 (N_1366,N_1305,N_1299);
nand U1367 (N_1367,N_1279,N_1275);
xnor U1368 (N_1368,N_1296,N_1289);
or U1369 (N_1369,N_1280,N_1303);
or U1370 (N_1370,N_1283,N_1314);
or U1371 (N_1371,N_1290,N_1289);
nor U1372 (N_1372,N_1318,N_1284);
nand U1373 (N_1373,N_1277,N_1303);
and U1374 (N_1374,N_1279,N_1293);
and U1375 (N_1375,N_1277,N_1315);
or U1376 (N_1376,N_1311,N_1318);
nor U1377 (N_1377,N_1293,N_1310);
or U1378 (N_1378,N_1286,N_1314);
nor U1379 (N_1379,N_1265,N_1304);
or U1380 (N_1380,N_1335,N_1349);
and U1381 (N_1381,N_1359,N_1322);
nand U1382 (N_1382,N_1365,N_1375);
nor U1383 (N_1383,N_1351,N_1323);
and U1384 (N_1384,N_1347,N_1356);
or U1385 (N_1385,N_1350,N_1379);
or U1386 (N_1386,N_1334,N_1370);
nand U1387 (N_1387,N_1348,N_1374);
nand U1388 (N_1388,N_1326,N_1361);
and U1389 (N_1389,N_1353,N_1357);
nand U1390 (N_1390,N_1364,N_1345);
nand U1391 (N_1391,N_1362,N_1342);
and U1392 (N_1392,N_1331,N_1329);
or U1393 (N_1393,N_1378,N_1354);
or U1394 (N_1394,N_1340,N_1366);
and U1395 (N_1395,N_1355,N_1360);
nor U1396 (N_1396,N_1320,N_1352);
and U1397 (N_1397,N_1377,N_1327);
nand U1398 (N_1398,N_1338,N_1339);
nor U1399 (N_1399,N_1372,N_1332);
nand U1400 (N_1400,N_1368,N_1324);
nor U1401 (N_1401,N_1328,N_1367);
and U1402 (N_1402,N_1369,N_1376);
nor U1403 (N_1403,N_1337,N_1343);
or U1404 (N_1404,N_1325,N_1363);
nor U1405 (N_1405,N_1333,N_1336);
or U1406 (N_1406,N_1371,N_1330);
or U1407 (N_1407,N_1358,N_1373);
or U1408 (N_1408,N_1344,N_1341);
nor U1409 (N_1409,N_1346,N_1321);
nor U1410 (N_1410,N_1336,N_1329);
xor U1411 (N_1411,N_1372,N_1358);
nand U1412 (N_1412,N_1340,N_1352);
nand U1413 (N_1413,N_1328,N_1350);
and U1414 (N_1414,N_1349,N_1324);
or U1415 (N_1415,N_1328,N_1357);
nor U1416 (N_1416,N_1373,N_1349);
nand U1417 (N_1417,N_1367,N_1339);
xnor U1418 (N_1418,N_1378,N_1379);
or U1419 (N_1419,N_1350,N_1364);
and U1420 (N_1420,N_1343,N_1360);
and U1421 (N_1421,N_1347,N_1342);
nand U1422 (N_1422,N_1350,N_1363);
and U1423 (N_1423,N_1370,N_1341);
or U1424 (N_1424,N_1326,N_1343);
and U1425 (N_1425,N_1338,N_1375);
nor U1426 (N_1426,N_1328,N_1369);
nor U1427 (N_1427,N_1356,N_1377);
and U1428 (N_1428,N_1335,N_1340);
and U1429 (N_1429,N_1324,N_1363);
nand U1430 (N_1430,N_1341,N_1347);
and U1431 (N_1431,N_1349,N_1322);
or U1432 (N_1432,N_1321,N_1348);
or U1433 (N_1433,N_1336,N_1335);
nand U1434 (N_1434,N_1359,N_1338);
nor U1435 (N_1435,N_1354,N_1324);
nor U1436 (N_1436,N_1367,N_1324);
nor U1437 (N_1437,N_1327,N_1366);
nand U1438 (N_1438,N_1356,N_1375);
nor U1439 (N_1439,N_1331,N_1338);
and U1440 (N_1440,N_1400,N_1435);
or U1441 (N_1441,N_1401,N_1389);
or U1442 (N_1442,N_1416,N_1404);
nand U1443 (N_1443,N_1427,N_1411);
or U1444 (N_1444,N_1415,N_1403);
nor U1445 (N_1445,N_1428,N_1423);
and U1446 (N_1446,N_1392,N_1429);
nor U1447 (N_1447,N_1388,N_1436);
or U1448 (N_1448,N_1408,N_1387);
and U1449 (N_1449,N_1399,N_1419);
nand U1450 (N_1450,N_1384,N_1397);
nand U1451 (N_1451,N_1418,N_1433);
and U1452 (N_1452,N_1439,N_1391);
or U1453 (N_1453,N_1432,N_1426);
or U1454 (N_1454,N_1380,N_1394);
nand U1455 (N_1455,N_1409,N_1414);
or U1456 (N_1456,N_1402,N_1420);
nor U1457 (N_1457,N_1421,N_1382);
and U1458 (N_1458,N_1412,N_1407);
and U1459 (N_1459,N_1425,N_1424);
nor U1460 (N_1460,N_1430,N_1438);
nand U1461 (N_1461,N_1390,N_1395);
nor U1462 (N_1462,N_1410,N_1393);
and U1463 (N_1463,N_1437,N_1413);
or U1464 (N_1464,N_1383,N_1434);
or U1465 (N_1465,N_1381,N_1417);
nor U1466 (N_1466,N_1398,N_1405);
or U1467 (N_1467,N_1406,N_1431);
nand U1468 (N_1468,N_1385,N_1422);
nor U1469 (N_1469,N_1386,N_1396);
or U1470 (N_1470,N_1414,N_1435);
nor U1471 (N_1471,N_1411,N_1381);
and U1472 (N_1472,N_1409,N_1400);
nand U1473 (N_1473,N_1399,N_1430);
and U1474 (N_1474,N_1422,N_1426);
and U1475 (N_1475,N_1433,N_1438);
and U1476 (N_1476,N_1418,N_1434);
nand U1477 (N_1477,N_1400,N_1419);
nor U1478 (N_1478,N_1387,N_1415);
and U1479 (N_1479,N_1390,N_1422);
or U1480 (N_1480,N_1414,N_1381);
xor U1481 (N_1481,N_1398,N_1404);
or U1482 (N_1482,N_1427,N_1398);
nand U1483 (N_1483,N_1420,N_1396);
or U1484 (N_1484,N_1434,N_1391);
nand U1485 (N_1485,N_1436,N_1396);
nand U1486 (N_1486,N_1431,N_1410);
and U1487 (N_1487,N_1401,N_1404);
nor U1488 (N_1488,N_1396,N_1385);
or U1489 (N_1489,N_1398,N_1415);
and U1490 (N_1490,N_1408,N_1406);
and U1491 (N_1491,N_1438,N_1410);
or U1492 (N_1492,N_1431,N_1416);
or U1493 (N_1493,N_1415,N_1435);
or U1494 (N_1494,N_1434,N_1414);
nand U1495 (N_1495,N_1380,N_1406);
nand U1496 (N_1496,N_1408,N_1385);
nand U1497 (N_1497,N_1388,N_1419);
or U1498 (N_1498,N_1424,N_1405);
nor U1499 (N_1499,N_1437,N_1424);
or U1500 (N_1500,N_1452,N_1446);
nand U1501 (N_1501,N_1465,N_1469);
nor U1502 (N_1502,N_1491,N_1467);
or U1503 (N_1503,N_1447,N_1463);
and U1504 (N_1504,N_1461,N_1468);
nor U1505 (N_1505,N_1479,N_1451);
and U1506 (N_1506,N_1453,N_1481);
nand U1507 (N_1507,N_1485,N_1466);
and U1508 (N_1508,N_1462,N_1449);
and U1509 (N_1509,N_1477,N_1478);
nand U1510 (N_1510,N_1476,N_1494);
nor U1511 (N_1511,N_1440,N_1450);
nand U1512 (N_1512,N_1499,N_1460);
or U1513 (N_1513,N_1484,N_1483);
and U1514 (N_1514,N_1475,N_1444);
and U1515 (N_1515,N_1445,N_1480);
or U1516 (N_1516,N_1457,N_1470);
nor U1517 (N_1517,N_1486,N_1488);
and U1518 (N_1518,N_1496,N_1489);
nand U1519 (N_1519,N_1464,N_1474);
and U1520 (N_1520,N_1472,N_1441);
or U1521 (N_1521,N_1443,N_1459);
and U1522 (N_1522,N_1487,N_1471);
nand U1523 (N_1523,N_1498,N_1493);
and U1524 (N_1524,N_1442,N_1497);
and U1525 (N_1525,N_1495,N_1482);
or U1526 (N_1526,N_1448,N_1456);
and U1527 (N_1527,N_1454,N_1458);
nand U1528 (N_1528,N_1455,N_1490);
nor U1529 (N_1529,N_1473,N_1492);
or U1530 (N_1530,N_1446,N_1448);
nand U1531 (N_1531,N_1444,N_1442);
nand U1532 (N_1532,N_1466,N_1447);
nand U1533 (N_1533,N_1488,N_1443);
or U1534 (N_1534,N_1479,N_1445);
nand U1535 (N_1535,N_1460,N_1491);
or U1536 (N_1536,N_1471,N_1488);
nor U1537 (N_1537,N_1492,N_1450);
or U1538 (N_1538,N_1466,N_1443);
nor U1539 (N_1539,N_1480,N_1447);
and U1540 (N_1540,N_1469,N_1462);
nand U1541 (N_1541,N_1466,N_1445);
nand U1542 (N_1542,N_1494,N_1466);
nor U1543 (N_1543,N_1484,N_1457);
and U1544 (N_1544,N_1497,N_1456);
and U1545 (N_1545,N_1455,N_1472);
nand U1546 (N_1546,N_1493,N_1468);
and U1547 (N_1547,N_1479,N_1477);
nor U1548 (N_1548,N_1444,N_1489);
nor U1549 (N_1549,N_1492,N_1498);
nand U1550 (N_1550,N_1456,N_1470);
and U1551 (N_1551,N_1454,N_1459);
or U1552 (N_1552,N_1490,N_1474);
nor U1553 (N_1553,N_1475,N_1446);
nand U1554 (N_1554,N_1462,N_1479);
and U1555 (N_1555,N_1483,N_1496);
or U1556 (N_1556,N_1495,N_1499);
nor U1557 (N_1557,N_1450,N_1469);
nor U1558 (N_1558,N_1443,N_1474);
nand U1559 (N_1559,N_1480,N_1452);
nand U1560 (N_1560,N_1521,N_1501);
nor U1561 (N_1561,N_1528,N_1508);
nor U1562 (N_1562,N_1506,N_1524);
nor U1563 (N_1563,N_1523,N_1527);
nor U1564 (N_1564,N_1518,N_1537);
nand U1565 (N_1565,N_1500,N_1522);
nor U1566 (N_1566,N_1555,N_1543);
or U1567 (N_1567,N_1542,N_1530);
and U1568 (N_1568,N_1517,N_1549);
and U1569 (N_1569,N_1502,N_1512);
or U1570 (N_1570,N_1554,N_1547);
nor U1571 (N_1571,N_1539,N_1513);
nor U1572 (N_1572,N_1511,N_1541);
and U1573 (N_1573,N_1552,N_1558);
nand U1574 (N_1574,N_1519,N_1533);
nand U1575 (N_1575,N_1525,N_1557);
or U1576 (N_1576,N_1534,N_1514);
or U1577 (N_1577,N_1538,N_1520);
nor U1578 (N_1578,N_1544,N_1526);
or U1579 (N_1579,N_1536,N_1532);
nand U1580 (N_1580,N_1551,N_1516);
nand U1581 (N_1581,N_1553,N_1529);
nor U1582 (N_1582,N_1556,N_1515);
or U1583 (N_1583,N_1545,N_1535);
and U1584 (N_1584,N_1505,N_1531);
and U1585 (N_1585,N_1550,N_1548);
nor U1586 (N_1586,N_1507,N_1540);
and U1587 (N_1587,N_1510,N_1503);
or U1588 (N_1588,N_1509,N_1559);
nor U1589 (N_1589,N_1546,N_1504);
nor U1590 (N_1590,N_1531,N_1555);
nand U1591 (N_1591,N_1525,N_1528);
nand U1592 (N_1592,N_1510,N_1527);
or U1593 (N_1593,N_1509,N_1523);
nand U1594 (N_1594,N_1545,N_1553);
and U1595 (N_1595,N_1541,N_1553);
nand U1596 (N_1596,N_1555,N_1530);
nor U1597 (N_1597,N_1549,N_1541);
nor U1598 (N_1598,N_1514,N_1532);
or U1599 (N_1599,N_1533,N_1523);
and U1600 (N_1600,N_1527,N_1530);
nand U1601 (N_1601,N_1526,N_1550);
and U1602 (N_1602,N_1548,N_1507);
nand U1603 (N_1603,N_1502,N_1557);
nand U1604 (N_1604,N_1522,N_1548);
and U1605 (N_1605,N_1527,N_1500);
nand U1606 (N_1606,N_1514,N_1559);
and U1607 (N_1607,N_1512,N_1510);
or U1608 (N_1608,N_1514,N_1540);
nand U1609 (N_1609,N_1536,N_1537);
or U1610 (N_1610,N_1551,N_1558);
nor U1611 (N_1611,N_1510,N_1543);
or U1612 (N_1612,N_1522,N_1528);
nor U1613 (N_1613,N_1516,N_1554);
nor U1614 (N_1614,N_1544,N_1549);
nor U1615 (N_1615,N_1527,N_1519);
and U1616 (N_1616,N_1518,N_1520);
nand U1617 (N_1617,N_1501,N_1508);
and U1618 (N_1618,N_1512,N_1511);
nand U1619 (N_1619,N_1501,N_1558);
nor U1620 (N_1620,N_1609,N_1582);
nor U1621 (N_1621,N_1617,N_1611);
nor U1622 (N_1622,N_1594,N_1565);
or U1623 (N_1623,N_1568,N_1560);
and U1624 (N_1624,N_1618,N_1581);
nand U1625 (N_1625,N_1576,N_1596);
nand U1626 (N_1626,N_1602,N_1599);
nand U1627 (N_1627,N_1613,N_1606);
nand U1628 (N_1628,N_1575,N_1561);
or U1629 (N_1629,N_1590,N_1566);
nand U1630 (N_1630,N_1574,N_1588);
nor U1631 (N_1631,N_1580,N_1603);
nand U1632 (N_1632,N_1612,N_1615);
and U1633 (N_1633,N_1572,N_1579);
and U1634 (N_1634,N_1604,N_1600);
nand U1635 (N_1635,N_1605,N_1584);
nand U1636 (N_1636,N_1610,N_1564);
nand U1637 (N_1637,N_1591,N_1601);
and U1638 (N_1638,N_1567,N_1577);
nand U1639 (N_1639,N_1583,N_1597);
and U1640 (N_1640,N_1562,N_1586);
nand U1641 (N_1641,N_1563,N_1593);
nand U1642 (N_1642,N_1587,N_1619);
nand U1643 (N_1643,N_1571,N_1598);
nor U1644 (N_1644,N_1589,N_1616);
nand U1645 (N_1645,N_1614,N_1573);
or U1646 (N_1646,N_1592,N_1585);
nand U1647 (N_1647,N_1607,N_1578);
nor U1648 (N_1648,N_1569,N_1570);
nor U1649 (N_1649,N_1608,N_1595);
and U1650 (N_1650,N_1575,N_1572);
and U1651 (N_1651,N_1569,N_1584);
nand U1652 (N_1652,N_1615,N_1561);
nor U1653 (N_1653,N_1572,N_1587);
or U1654 (N_1654,N_1566,N_1613);
and U1655 (N_1655,N_1570,N_1590);
and U1656 (N_1656,N_1593,N_1609);
and U1657 (N_1657,N_1572,N_1591);
or U1658 (N_1658,N_1611,N_1574);
and U1659 (N_1659,N_1565,N_1618);
or U1660 (N_1660,N_1561,N_1583);
nand U1661 (N_1661,N_1593,N_1610);
and U1662 (N_1662,N_1565,N_1564);
nor U1663 (N_1663,N_1561,N_1577);
nand U1664 (N_1664,N_1608,N_1617);
or U1665 (N_1665,N_1610,N_1605);
and U1666 (N_1666,N_1560,N_1597);
and U1667 (N_1667,N_1601,N_1586);
and U1668 (N_1668,N_1609,N_1591);
or U1669 (N_1669,N_1576,N_1597);
or U1670 (N_1670,N_1562,N_1571);
nand U1671 (N_1671,N_1581,N_1611);
nor U1672 (N_1672,N_1581,N_1563);
and U1673 (N_1673,N_1568,N_1614);
nand U1674 (N_1674,N_1571,N_1591);
and U1675 (N_1675,N_1619,N_1596);
or U1676 (N_1676,N_1587,N_1600);
nor U1677 (N_1677,N_1600,N_1581);
nand U1678 (N_1678,N_1609,N_1610);
or U1679 (N_1679,N_1612,N_1606);
nand U1680 (N_1680,N_1621,N_1630);
or U1681 (N_1681,N_1638,N_1648);
nand U1682 (N_1682,N_1626,N_1623);
nor U1683 (N_1683,N_1667,N_1637);
or U1684 (N_1684,N_1661,N_1674);
nand U1685 (N_1685,N_1622,N_1647);
or U1686 (N_1686,N_1655,N_1669);
nand U1687 (N_1687,N_1662,N_1675);
and U1688 (N_1688,N_1665,N_1634);
and U1689 (N_1689,N_1666,N_1677);
nand U1690 (N_1690,N_1643,N_1658);
and U1691 (N_1691,N_1644,N_1660);
or U1692 (N_1692,N_1646,N_1679);
and U1693 (N_1693,N_1631,N_1672);
nand U1694 (N_1694,N_1624,N_1668);
or U1695 (N_1695,N_1663,N_1639);
and U1696 (N_1696,N_1652,N_1653);
or U1697 (N_1697,N_1651,N_1642);
nand U1698 (N_1698,N_1645,N_1627);
nand U1699 (N_1699,N_1636,N_1676);
and U1700 (N_1700,N_1620,N_1633);
nand U1701 (N_1701,N_1640,N_1670);
or U1702 (N_1702,N_1678,N_1664);
or U1703 (N_1703,N_1649,N_1650);
nor U1704 (N_1704,N_1657,N_1654);
nor U1705 (N_1705,N_1659,N_1635);
and U1706 (N_1706,N_1673,N_1632);
or U1707 (N_1707,N_1656,N_1671);
or U1708 (N_1708,N_1628,N_1641);
or U1709 (N_1709,N_1629,N_1625);
and U1710 (N_1710,N_1670,N_1638);
nor U1711 (N_1711,N_1626,N_1670);
nand U1712 (N_1712,N_1627,N_1632);
nand U1713 (N_1713,N_1674,N_1666);
nor U1714 (N_1714,N_1658,N_1635);
nor U1715 (N_1715,N_1679,N_1629);
and U1716 (N_1716,N_1633,N_1654);
nand U1717 (N_1717,N_1644,N_1667);
or U1718 (N_1718,N_1661,N_1655);
nand U1719 (N_1719,N_1665,N_1625);
or U1720 (N_1720,N_1642,N_1645);
nor U1721 (N_1721,N_1653,N_1658);
nand U1722 (N_1722,N_1669,N_1653);
and U1723 (N_1723,N_1645,N_1653);
nand U1724 (N_1724,N_1653,N_1662);
xor U1725 (N_1725,N_1653,N_1648);
and U1726 (N_1726,N_1657,N_1635);
nand U1727 (N_1727,N_1647,N_1649);
or U1728 (N_1728,N_1629,N_1637);
nor U1729 (N_1729,N_1631,N_1673);
nand U1730 (N_1730,N_1657,N_1672);
nor U1731 (N_1731,N_1633,N_1650);
nand U1732 (N_1732,N_1639,N_1634);
or U1733 (N_1733,N_1659,N_1670);
and U1734 (N_1734,N_1620,N_1675);
and U1735 (N_1735,N_1639,N_1622);
nand U1736 (N_1736,N_1634,N_1675);
nand U1737 (N_1737,N_1670,N_1678);
or U1738 (N_1738,N_1620,N_1642);
and U1739 (N_1739,N_1657,N_1662);
and U1740 (N_1740,N_1710,N_1735);
nor U1741 (N_1741,N_1717,N_1705);
or U1742 (N_1742,N_1692,N_1713);
nor U1743 (N_1743,N_1694,N_1691);
nand U1744 (N_1744,N_1681,N_1724);
nand U1745 (N_1745,N_1737,N_1708);
and U1746 (N_1746,N_1693,N_1729);
and U1747 (N_1747,N_1711,N_1726);
and U1748 (N_1748,N_1727,N_1704);
nand U1749 (N_1749,N_1697,N_1703);
nor U1750 (N_1750,N_1706,N_1687);
nand U1751 (N_1751,N_1701,N_1686);
nor U1752 (N_1752,N_1689,N_1712);
nor U1753 (N_1753,N_1736,N_1682);
and U1754 (N_1754,N_1698,N_1739);
nor U1755 (N_1755,N_1733,N_1690);
and U1756 (N_1756,N_1684,N_1732);
or U1757 (N_1757,N_1716,N_1685);
or U1758 (N_1758,N_1695,N_1699);
or U1759 (N_1759,N_1720,N_1734);
nor U1760 (N_1760,N_1728,N_1702);
nand U1761 (N_1761,N_1700,N_1709);
nor U1762 (N_1762,N_1715,N_1714);
nand U1763 (N_1763,N_1680,N_1688);
nand U1764 (N_1764,N_1730,N_1696);
and U1765 (N_1765,N_1718,N_1707);
and U1766 (N_1766,N_1719,N_1723);
nor U1767 (N_1767,N_1738,N_1722);
and U1768 (N_1768,N_1721,N_1725);
nor U1769 (N_1769,N_1731,N_1683);
xnor U1770 (N_1770,N_1731,N_1697);
nor U1771 (N_1771,N_1699,N_1717);
and U1772 (N_1772,N_1733,N_1738);
nand U1773 (N_1773,N_1691,N_1732);
and U1774 (N_1774,N_1707,N_1687);
nor U1775 (N_1775,N_1737,N_1714);
nor U1776 (N_1776,N_1715,N_1701);
and U1777 (N_1777,N_1710,N_1720);
nor U1778 (N_1778,N_1693,N_1727);
nor U1779 (N_1779,N_1728,N_1683);
and U1780 (N_1780,N_1735,N_1733);
and U1781 (N_1781,N_1703,N_1712);
nand U1782 (N_1782,N_1720,N_1728);
and U1783 (N_1783,N_1689,N_1729);
nor U1784 (N_1784,N_1689,N_1728);
or U1785 (N_1785,N_1721,N_1707);
nor U1786 (N_1786,N_1727,N_1703);
nor U1787 (N_1787,N_1691,N_1727);
or U1788 (N_1788,N_1682,N_1721);
xnor U1789 (N_1789,N_1696,N_1736);
or U1790 (N_1790,N_1718,N_1695);
nor U1791 (N_1791,N_1683,N_1680);
nand U1792 (N_1792,N_1691,N_1725);
nor U1793 (N_1793,N_1737,N_1705);
nand U1794 (N_1794,N_1695,N_1711);
nor U1795 (N_1795,N_1723,N_1682);
nand U1796 (N_1796,N_1682,N_1708);
and U1797 (N_1797,N_1701,N_1726);
or U1798 (N_1798,N_1682,N_1687);
and U1799 (N_1799,N_1695,N_1730);
nand U1800 (N_1800,N_1767,N_1760);
and U1801 (N_1801,N_1772,N_1784);
nor U1802 (N_1802,N_1783,N_1774);
nor U1803 (N_1803,N_1757,N_1749);
and U1804 (N_1804,N_1777,N_1762);
or U1805 (N_1805,N_1799,N_1752);
and U1806 (N_1806,N_1761,N_1759);
and U1807 (N_1807,N_1758,N_1765);
nor U1808 (N_1808,N_1764,N_1756);
or U1809 (N_1809,N_1743,N_1755);
nand U1810 (N_1810,N_1747,N_1795);
or U1811 (N_1811,N_1753,N_1779);
nand U1812 (N_1812,N_1776,N_1798);
or U1813 (N_1813,N_1740,N_1768);
or U1814 (N_1814,N_1778,N_1770);
and U1815 (N_1815,N_1793,N_1788);
nor U1816 (N_1816,N_1763,N_1771);
or U1817 (N_1817,N_1746,N_1750);
and U1818 (N_1818,N_1782,N_1791);
and U1819 (N_1819,N_1775,N_1773);
and U1820 (N_1820,N_1744,N_1745);
nor U1821 (N_1821,N_1796,N_1785);
and U1822 (N_1822,N_1751,N_1789);
nand U1823 (N_1823,N_1792,N_1742);
nand U1824 (N_1824,N_1741,N_1754);
nand U1825 (N_1825,N_1794,N_1766);
nand U1826 (N_1826,N_1787,N_1790);
nor U1827 (N_1827,N_1797,N_1748);
and U1828 (N_1828,N_1786,N_1780);
or U1829 (N_1829,N_1769,N_1781);
and U1830 (N_1830,N_1781,N_1794);
nor U1831 (N_1831,N_1781,N_1784);
nand U1832 (N_1832,N_1798,N_1758);
nand U1833 (N_1833,N_1798,N_1790);
or U1834 (N_1834,N_1795,N_1781);
nand U1835 (N_1835,N_1789,N_1793);
and U1836 (N_1836,N_1789,N_1795);
nor U1837 (N_1837,N_1787,N_1754);
nor U1838 (N_1838,N_1786,N_1772);
nand U1839 (N_1839,N_1783,N_1744);
nor U1840 (N_1840,N_1775,N_1777);
or U1841 (N_1841,N_1774,N_1798);
nand U1842 (N_1842,N_1771,N_1744);
and U1843 (N_1843,N_1748,N_1786);
nor U1844 (N_1844,N_1758,N_1781);
nor U1845 (N_1845,N_1778,N_1754);
nand U1846 (N_1846,N_1790,N_1767);
or U1847 (N_1847,N_1740,N_1743);
and U1848 (N_1848,N_1782,N_1754);
or U1849 (N_1849,N_1741,N_1769);
and U1850 (N_1850,N_1799,N_1778);
and U1851 (N_1851,N_1799,N_1784);
nor U1852 (N_1852,N_1779,N_1749);
nand U1853 (N_1853,N_1775,N_1778);
or U1854 (N_1854,N_1752,N_1775);
nor U1855 (N_1855,N_1794,N_1767);
and U1856 (N_1856,N_1746,N_1761);
or U1857 (N_1857,N_1796,N_1748);
nand U1858 (N_1858,N_1756,N_1775);
nand U1859 (N_1859,N_1776,N_1791);
nand U1860 (N_1860,N_1848,N_1831);
or U1861 (N_1861,N_1832,N_1836);
or U1862 (N_1862,N_1822,N_1807);
or U1863 (N_1863,N_1844,N_1814);
and U1864 (N_1864,N_1827,N_1833);
nand U1865 (N_1865,N_1828,N_1838);
and U1866 (N_1866,N_1845,N_1808);
nand U1867 (N_1867,N_1834,N_1805);
nor U1868 (N_1868,N_1847,N_1850);
and U1869 (N_1869,N_1843,N_1859);
and U1870 (N_1870,N_1830,N_1804);
and U1871 (N_1871,N_1841,N_1820);
nor U1872 (N_1872,N_1802,N_1849);
nor U1873 (N_1873,N_1812,N_1810);
nor U1874 (N_1874,N_1803,N_1800);
or U1875 (N_1875,N_1837,N_1809);
nand U1876 (N_1876,N_1819,N_1806);
and U1877 (N_1877,N_1826,N_1856);
nand U1878 (N_1878,N_1854,N_1823);
and U1879 (N_1879,N_1852,N_1817);
nand U1880 (N_1880,N_1825,N_1801);
nor U1881 (N_1881,N_1855,N_1842);
nor U1882 (N_1882,N_1853,N_1818);
nor U1883 (N_1883,N_1840,N_1813);
xor U1884 (N_1884,N_1811,N_1816);
or U1885 (N_1885,N_1824,N_1839);
or U1886 (N_1886,N_1821,N_1815);
or U1887 (N_1887,N_1829,N_1846);
or U1888 (N_1888,N_1851,N_1858);
and U1889 (N_1889,N_1857,N_1835);
and U1890 (N_1890,N_1829,N_1816);
and U1891 (N_1891,N_1814,N_1838);
or U1892 (N_1892,N_1822,N_1834);
xnor U1893 (N_1893,N_1858,N_1801);
nor U1894 (N_1894,N_1851,N_1854);
nor U1895 (N_1895,N_1811,N_1821);
or U1896 (N_1896,N_1852,N_1826);
or U1897 (N_1897,N_1835,N_1844);
or U1898 (N_1898,N_1842,N_1804);
nor U1899 (N_1899,N_1807,N_1811);
nand U1900 (N_1900,N_1831,N_1832);
or U1901 (N_1901,N_1825,N_1847);
and U1902 (N_1902,N_1804,N_1803);
or U1903 (N_1903,N_1843,N_1851);
or U1904 (N_1904,N_1840,N_1830);
nand U1905 (N_1905,N_1805,N_1855);
nor U1906 (N_1906,N_1801,N_1809);
nor U1907 (N_1907,N_1829,N_1822);
or U1908 (N_1908,N_1809,N_1854);
nor U1909 (N_1909,N_1816,N_1832);
and U1910 (N_1910,N_1813,N_1824);
or U1911 (N_1911,N_1858,N_1820);
nor U1912 (N_1912,N_1857,N_1855);
nor U1913 (N_1913,N_1841,N_1807);
nor U1914 (N_1914,N_1834,N_1852);
nor U1915 (N_1915,N_1820,N_1855);
nor U1916 (N_1916,N_1814,N_1851);
and U1917 (N_1917,N_1819,N_1803);
or U1918 (N_1918,N_1849,N_1854);
or U1919 (N_1919,N_1827,N_1828);
and U1920 (N_1920,N_1867,N_1862);
or U1921 (N_1921,N_1902,N_1919);
nor U1922 (N_1922,N_1910,N_1881);
and U1923 (N_1923,N_1875,N_1873);
nand U1924 (N_1924,N_1888,N_1864);
nand U1925 (N_1925,N_1871,N_1870);
nand U1926 (N_1926,N_1877,N_1897);
or U1927 (N_1927,N_1916,N_1904);
or U1928 (N_1928,N_1893,N_1900);
or U1929 (N_1929,N_1907,N_1917);
and U1930 (N_1930,N_1913,N_1898);
and U1931 (N_1931,N_1861,N_1887);
nand U1932 (N_1932,N_1878,N_1892);
nand U1933 (N_1933,N_1874,N_1880);
or U1934 (N_1934,N_1879,N_1918);
nand U1935 (N_1935,N_1912,N_1885);
and U1936 (N_1936,N_1905,N_1899);
xnor U1937 (N_1937,N_1896,N_1860);
nor U1938 (N_1938,N_1911,N_1914);
nand U1939 (N_1939,N_1866,N_1865);
nor U1940 (N_1940,N_1915,N_1863);
nor U1941 (N_1941,N_1889,N_1876);
nand U1942 (N_1942,N_1886,N_1908);
and U1943 (N_1943,N_1872,N_1890);
nand U1944 (N_1944,N_1884,N_1906);
nand U1945 (N_1945,N_1909,N_1882);
and U1946 (N_1946,N_1895,N_1894);
and U1947 (N_1947,N_1903,N_1883);
and U1948 (N_1948,N_1869,N_1868);
nor U1949 (N_1949,N_1901,N_1891);
and U1950 (N_1950,N_1890,N_1882);
nand U1951 (N_1951,N_1892,N_1874);
or U1952 (N_1952,N_1896,N_1871);
nor U1953 (N_1953,N_1897,N_1888);
and U1954 (N_1954,N_1893,N_1915);
nand U1955 (N_1955,N_1890,N_1900);
and U1956 (N_1956,N_1899,N_1908);
nor U1957 (N_1957,N_1909,N_1912);
or U1958 (N_1958,N_1900,N_1897);
and U1959 (N_1959,N_1899,N_1882);
or U1960 (N_1960,N_1878,N_1890);
and U1961 (N_1961,N_1864,N_1882);
or U1962 (N_1962,N_1905,N_1904);
nor U1963 (N_1963,N_1869,N_1901);
nand U1964 (N_1964,N_1917,N_1884);
nor U1965 (N_1965,N_1875,N_1897);
or U1966 (N_1966,N_1881,N_1882);
or U1967 (N_1967,N_1873,N_1904);
or U1968 (N_1968,N_1866,N_1907);
nand U1969 (N_1969,N_1885,N_1903);
nor U1970 (N_1970,N_1914,N_1861);
nand U1971 (N_1971,N_1875,N_1872);
and U1972 (N_1972,N_1915,N_1881);
or U1973 (N_1973,N_1869,N_1899);
nor U1974 (N_1974,N_1908,N_1883);
or U1975 (N_1975,N_1864,N_1860);
or U1976 (N_1976,N_1864,N_1915);
or U1977 (N_1977,N_1916,N_1872);
or U1978 (N_1978,N_1870,N_1915);
or U1979 (N_1979,N_1917,N_1897);
or U1980 (N_1980,N_1966,N_1945);
and U1981 (N_1981,N_1921,N_1934);
and U1982 (N_1982,N_1956,N_1938);
nor U1983 (N_1983,N_1940,N_1979);
nor U1984 (N_1984,N_1931,N_1930);
and U1985 (N_1985,N_1943,N_1961);
and U1986 (N_1986,N_1974,N_1926);
and U1987 (N_1987,N_1969,N_1960);
nor U1988 (N_1988,N_1967,N_1946);
nor U1989 (N_1989,N_1975,N_1948);
and U1990 (N_1990,N_1949,N_1954);
nor U1991 (N_1991,N_1959,N_1957);
and U1992 (N_1992,N_1935,N_1950);
and U1993 (N_1993,N_1972,N_1955);
nor U1994 (N_1994,N_1944,N_1965);
and U1995 (N_1995,N_1927,N_1977);
and U1996 (N_1996,N_1936,N_1925);
nor U1997 (N_1997,N_1932,N_1937);
or U1998 (N_1998,N_1922,N_1962);
nand U1999 (N_1999,N_1942,N_1928);
and U2000 (N_2000,N_1952,N_1941);
or U2001 (N_2001,N_1953,N_1923);
and U2002 (N_2002,N_1947,N_1951);
nand U2003 (N_2003,N_1968,N_1920);
xnor U2004 (N_2004,N_1978,N_1929);
and U2005 (N_2005,N_1973,N_1933);
nand U2006 (N_2006,N_1958,N_1976);
and U2007 (N_2007,N_1939,N_1964);
or U2008 (N_2008,N_1971,N_1970);
and U2009 (N_2009,N_1924,N_1963);
nor U2010 (N_2010,N_1944,N_1960);
and U2011 (N_2011,N_1922,N_1933);
nand U2012 (N_2012,N_1935,N_1931);
nand U2013 (N_2013,N_1955,N_1969);
nand U2014 (N_2014,N_1942,N_1957);
nand U2015 (N_2015,N_1924,N_1971);
or U2016 (N_2016,N_1928,N_1953);
and U2017 (N_2017,N_1950,N_1922);
or U2018 (N_2018,N_1969,N_1977);
nand U2019 (N_2019,N_1962,N_1932);
or U2020 (N_2020,N_1936,N_1922);
and U2021 (N_2021,N_1967,N_1952);
nand U2022 (N_2022,N_1932,N_1927);
and U2023 (N_2023,N_1970,N_1958);
or U2024 (N_2024,N_1928,N_1962);
and U2025 (N_2025,N_1951,N_1979);
nor U2026 (N_2026,N_1952,N_1956);
or U2027 (N_2027,N_1949,N_1926);
or U2028 (N_2028,N_1959,N_1937);
and U2029 (N_2029,N_1955,N_1926);
or U2030 (N_2030,N_1932,N_1925);
nor U2031 (N_2031,N_1954,N_1942);
nor U2032 (N_2032,N_1929,N_1941);
and U2033 (N_2033,N_1956,N_1976);
and U2034 (N_2034,N_1920,N_1928);
nor U2035 (N_2035,N_1961,N_1931);
or U2036 (N_2036,N_1975,N_1965);
or U2037 (N_2037,N_1931,N_1940);
and U2038 (N_2038,N_1928,N_1968);
nor U2039 (N_2039,N_1959,N_1955);
nor U2040 (N_2040,N_2015,N_2003);
and U2041 (N_2041,N_2022,N_2034);
nor U2042 (N_2042,N_1985,N_1982);
or U2043 (N_2043,N_1991,N_2038);
or U2044 (N_2044,N_1999,N_2006);
or U2045 (N_2045,N_2033,N_2018);
and U2046 (N_2046,N_1987,N_2024);
nand U2047 (N_2047,N_2017,N_2028);
nor U2048 (N_2048,N_1997,N_2029);
nor U2049 (N_2049,N_2014,N_2027);
and U2050 (N_2050,N_1984,N_2037);
or U2051 (N_2051,N_2013,N_2001);
and U2052 (N_2052,N_2009,N_2019);
and U2053 (N_2053,N_2012,N_2007);
xor U2054 (N_2054,N_2031,N_2004);
nand U2055 (N_2055,N_2039,N_2008);
xnor U2056 (N_2056,N_1994,N_2032);
and U2057 (N_2057,N_1990,N_2002);
nand U2058 (N_2058,N_1993,N_2030);
nand U2059 (N_2059,N_1986,N_2016);
nor U2060 (N_2060,N_1992,N_1983);
nor U2061 (N_2061,N_1981,N_2036);
nand U2062 (N_2062,N_2035,N_2021);
and U2063 (N_2063,N_2025,N_2000);
and U2064 (N_2064,N_1980,N_2020);
nor U2065 (N_2065,N_2011,N_2023);
or U2066 (N_2066,N_2010,N_2005);
nor U2067 (N_2067,N_2026,N_1998);
nor U2068 (N_2068,N_1989,N_1996);
nand U2069 (N_2069,N_1988,N_1995);
nor U2070 (N_2070,N_1987,N_2029);
nand U2071 (N_2071,N_1996,N_2003);
nand U2072 (N_2072,N_2033,N_1980);
xnor U2073 (N_2073,N_2022,N_2023);
nor U2074 (N_2074,N_2016,N_1998);
nand U2075 (N_2075,N_2023,N_2016);
nand U2076 (N_2076,N_1993,N_2011);
xor U2077 (N_2077,N_2014,N_2010);
and U2078 (N_2078,N_2001,N_2028);
and U2079 (N_2079,N_1984,N_2020);
nor U2080 (N_2080,N_2012,N_2014);
nand U2081 (N_2081,N_2027,N_2000);
nor U2082 (N_2082,N_2038,N_2018);
nor U2083 (N_2083,N_2001,N_2022);
nor U2084 (N_2084,N_1988,N_2037);
or U2085 (N_2085,N_2017,N_2037);
nor U2086 (N_2086,N_2039,N_1982);
nor U2087 (N_2087,N_1990,N_2037);
xor U2088 (N_2088,N_2002,N_2025);
or U2089 (N_2089,N_2011,N_2036);
or U2090 (N_2090,N_2034,N_2023);
and U2091 (N_2091,N_2016,N_1980);
or U2092 (N_2092,N_1981,N_2012);
nor U2093 (N_2093,N_1990,N_1984);
nor U2094 (N_2094,N_1991,N_2023);
nor U2095 (N_2095,N_2016,N_2039);
nand U2096 (N_2096,N_2035,N_2038);
nand U2097 (N_2097,N_2003,N_1994);
nor U2098 (N_2098,N_2016,N_2018);
or U2099 (N_2099,N_2028,N_2018);
nor U2100 (N_2100,N_2089,N_2058);
nand U2101 (N_2101,N_2042,N_2079);
nand U2102 (N_2102,N_2068,N_2044);
nand U2103 (N_2103,N_2056,N_2086);
nor U2104 (N_2104,N_2057,N_2049);
nand U2105 (N_2105,N_2099,N_2072);
or U2106 (N_2106,N_2055,N_2092);
nand U2107 (N_2107,N_2048,N_2053);
and U2108 (N_2108,N_2067,N_2062);
or U2109 (N_2109,N_2075,N_2045);
nand U2110 (N_2110,N_2076,N_2041);
or U2111 (N_2111,N_2081,N_2083);
nand U2112 (N_2112,N_2064,N_2043);
or U2113 (N_2113,N_2059,N_2047);
and U2114 (N_2114,N_2065,N_2080);
or U2115 (N_2115,N_2069,N_2054);
nor U2116 (N_2116,N_2098,N_2050);
nand U2117 (N_2117,N_2097,N_2061);
nor U2118 (N_2118,N_2094,N_2085);
nor U2119 (N_2119,N_2077,N_2040);
or U2120 (N_2120,N_2073,N_2087);
and U2121 (N_2121,N_2096,N_2091);
and U2122 (N_2122,N_2066,N_2082);
nor U2123 (N_2123,N_2070,N_2052);
or U2124 (N_2124,N_2071,N_2046);
nor U2125 (N_2125,N_2060,N_2074);
nand U2126 (N_2126,N_2090,N_2063);
or U2127 (N_2127,N_2095,N_2093);
nand U2128 (N_2128,N_2051,N_2088);
and U2129 (N_2129,N_2084,N_2078);
nor U2130 (N_2130,N_2076,N_2050);
nor U2131 (N_2131,N_2083,N_2041);
nor U2132 (N_2132,N_2077,N_2097);
or U2133 (N_2133,N_2084,N_2041);
nand U2134 (N_2134,N_2081,N_2085);
nor U2135 (N_2135,N_2073,N_2053);
nor U2136 (N_2136,N_2048,N_2041);
nand U2137 (N_2137,N_2092,N_2065);
nand U2138 (N_2138,N_2047,N_2099);
nand U2139 (N_2139,N_2094,N_2099);
nor U2140 (N_2140,N_2076,N_2096);
and U2141 (N_2141,N_2092,N_2089);
nand U2142 (N_2142,N_2058,N_2045);
and U2143 (N_2143,N_2061,N_2085);
and U2144 (N_2144,N_2044,N_2072);
or U2145 (N_2145,N_2053,N_2043);
and U2146 (N_2146,N_2076,N_2048);
or U2147 (N_2147,N_2051,N_2082);
or U2148 (N_2148,N_2099,N_2073);
nor U2149 (N_2149,N_2047,N_2085);
or U2150 (N_2150,N_2074,N_2087);
nand U2151 (N_2151,N_2071,N_2097);
or U2152 (N_2152,N_2080,N_2044);
and U2153 (N_2153,N_2071,N_2093);
or U2154 (N_2154,N_2049,N_2093);
or U2155 (N_2155,N_2041,N_2063);
and U2156 (N_2156,N_2056,N_2092);
and U2157 (N_2157,N_2074,N_2049);
nor U2158 (N_2158,N_2045,N_2091);
and U2159 (N_2159,N_2041,N_2040);
nor U2160 (N_2160,N_2113,N_2146);
nand U2161 (N_2161,N_2104,N_2156);
and U2162 (N_2162,N_2155,N_2153);
or U2163 (N_2163,N_2107,N_2128);
or U2164 (N_2164,N_2120,N_2114);
nor U2165 (N_2165,N_2135,N_2105);
nand U2166 (N_2166,N_2149,N_2116);
nand U2167 (N_2167,N_2102,N_2115);
and U2168 (N_2168,N_2139,N_2143);
nand U2169 (N_2169,N_2159,N_2137);
or U2170 (N_2170,N_2141,N_2132);
nand U2171 (N_2171,N_2133,N_2123);
nand U2172 (N_2172,N_2157,N_2130);
or U2173 (N_2173,N_2131,N_2122);
and U2174 (N_2174,N_2126,N_2121);
nand U2175 (N_2175,N_2150,N_2151);
nor U2176 (N_2176,N_2119,N_2127);
nor U2177 (N_2177,N_2124,N_2103);
and U2178 (N_2178,N_2110,N_2118);
nor U2179 (N_2179,N_2109,N_2138);
or U2180 (N_2180,N_2101,N_2108);
or U2181 (N_2181,N_2117,N_2140);
or U2182 (N_2182,N_2142,N_2106);
nand U2183 (N_2183,N_2145,N_2152);
nor U2184 (N_2184,N_2129,N_2134);
nor U2185 (N_2185,N_2136,N_2144);
nand U2186 (N_2186,N_2148,N_2100);
nand U2187 (N_2187,N_2125,N_2154);
or U2188 (N_2188,N_2147,N_2111);
nand U2189 (N_2189,N_2158,N_2112);
nor U2190 (N_2190,N_2114,N_2148);
and U2191 (N_2191,N_2129,N_2115);
or U2192 (N_2192,N_2119,N_2141);
nand U2193 (N_2193,N_2146,N_2119);
nand U2194 (N_2194,N_2126,N_2103);
and U2195 (N_2195,N_2156,N_2132);
nand U2196 (N_2196,N_2153,N_2122);
and U2197 (N_2197,N_2142,N_2158);
nand U2198 (N_2198,N_2144,N_2109);
or U2199 (N_2199,N_2122,N_2148);
or U2200 (N_2200,N_2126,N_2134);
and U2201 (N_2201,N_2121,N_2149);
and U2202 (N_2202,N_2136,N_2112);
or U2203 (N_2203,N_2145,N_2100);
nor U2204 (N_2204,N_2121,N_2136);
or U2205 (N_2205,N_2134,N_2147);
or U2206 (N_2206,N_2144,N_2104);
xor U2207 (N_2207,N_2152,N_2138);
nor U2208 (N_2208,N_2144,N_2159);
or U2209 (N_2209,N_2152,N_2153);
nand U2210 (N_2210,N_2124,N_2134);
or U2211 (N_2211,N_2106,N_2140);
and U2212 (N_2212,N_2100,N_2116);
or U2213 (N_2213,N_2120,N_2148);
nand U2214 (N_2214,N_2157,N_2104);
and U2215 (N_2215,N_2158,N_2151);
nor U2216 (N_2216,N_2122,N_2107);
nand U2217 (N_2217,N_2126,N_2112);
nor U2218 (N_2218,N_2122,N_2144);
nand U2219 (N_2219,N_2158,N_2136);
or U2220 (N_2220,N_2176,N_2208);
or U2221 (N_2221,N_2196,N_2199);
and U2222 (N_2222,N_2183,N_2162);
nand U2223 (N_2223,N_2170,N_2172);
or U2224 (N_2224,N_2191,N_2218);
nand U2225 (N_2225,N_2190,N_2169);
nand U2226 (N_2226,N_2205,N_2210);
nor U2227 (N_2227,N_2192,N_2175);
nand U2228 (N_2228,N_2164,N_2201);
and U2229 (N_2229,N_2194,N_2215);
and U2230 (N_2230,N_2219,N_2182);
nand U2231 (N_2231,N_2209,N_2198);
and U2232 (N_2232,N_2206,N_2163);
and U2233 (N_2233,N_2161,N_2203);
and U2234 (N_2234,N_2197,N_2160);
or U2235 (N_2235,N_2207,N_2187);
nor U2236 (N_2236,N_2213,N_2168);
nor U2237 (N_2237,N_2184,N_2202);
or U2238 (N_2238,N_2193,N_2180);
nor U2239 (N_2239,N_2174,N_2188);
nand U2240 (N_2240,N_2177,N_2217);
and U2241 (N_2241,N_2200,N_2181);
or U2242 (N_2242,N_2165,N_2214);
nand U2243 (N_2243,N_2216,N_2178);
or U2244 (N_2244,N_2166,N_2185);
and U2245 (N_2245,N_2195,N_2173);
and U2246 (N_2246,N_2186,N_2171);
nor U2247 (N_2247,N_2211,N_2189);
and U2248 (N_2248,N_2167,N_2179);
and U2249 (N_2249,N_2212,N_2204);
nand U2250 (N_2250,N_2171,N_2166);
or U2251 (N_2251,N_2193,N_2218);
or U2252 (N_2252,N_2199,N_2183);
and U2253 (N_2253,N_2180,N_2217);
and U2254 (N_2254,N_2199,N_2219);
and U2255 (N_2255,N_2177,N_2190);
or U2256 (N_2256,N_2161,N_2214);
or U2257 (N_2257,N_2218,N_2174);
and U2258 (N_2258,N_2165,N_2185);
nand U2259 (N_2259,N_2210,N_2165);
nand U2260 (N_2260,N_2177,N_2162);
xnor U2261 (N_2261,N_2178,N_2215);
nor U2262 (N_2262,N_2175,N_2217);
and U2263 (N_2263,N_2194,N_2191);
and U2264 (N_2264,N_2186,N_2205);
and U2265 (N_2265,N_2160,N_2161);
or U2266 (N_2266,N_2195,N_2160);
nand U2267 (N_2267,N_2216,N_2194);
or U2268 (N_2268,N_2183,N_2174);
nand U2269 (N_2269,N_2173,N_2217);
or U2270 (N_2270,N_2184,N_2172);
and U2271 (N_2271,N_2184,N_2213);
nor U2272 (N_2272,N_2180,N_2176);
nand U2273 (N_2273,N_2177,N_2198);
nand U2274 (N_2274,N_2201,N_2204);
and U2275 (N_2275,N_2179,N_2188);
nor U2276 (N_2276,N_2213,N_2192);
nor U2277 (N_2277,N_2219,N_2173);
or U2278 (N_2278,N_2183,N_2209);
or U2279 (N_2279,N_2191,N_2204);
or U2280 (N_2280,N_2273,N_2235);
or U2281 (N_2281,N_2249,N_2279);
and U2282 (N_2282,N_2246,N_2268);
and U2283 (N_2283,N_2259,N_2258);
or U2284 (N_2284,N_2223,N_2221);
nand U2285 (N_2285,N_2269,N_2264);
nor U2286 (N_2286,N_2265,N_2270);
nor U2287 (N_2287,N_2227,N_2247);
or U2288 (N_2288,N_2243,N_2224);
or U2289 (N_2289,N_2263,N_2239);
nand U2290 (N_2290,N_2262,N_2238);
and U2291 (N_2291,N_2255,N_2253);
and U2292 (N_2292,N_2231,N_2241);
or U2293 (N_2293,N_2242,N_2275);
or U2294 (N_2294,N_2278,N_2245);
and U2295 (N_2295,N_2254,N_2267);
or U2296 (N_2296,N_2251,N_2228);
nand U2297 (N_2297,N_2232,N_2244);
or U2298 (N_2298,N_2272,N_2248);
nor U2299 (N_2299,N_2250,N_2256);
and U2300 (N_2300,N_2222,N_2261);
and U2301 (N_2301,N_2230,N_2237);
and U2302 (N_2302,N_2220,N_2260);
nand U2303 (N_2303,N_2226,N_2229);
nand U2304 (N_2304,N_2233,N_2277);
nand U2305 (N_2305,N_2225,N_2274);
xor U2306 (N_2306,N_2271,N_2240);
nand U2307 (N_2307,N_2257,N_2234);
nor U2308 (N_2308,N_2266,N_2252);
nand U2309 (N_2309,N_2236,N_2276);
or U2310 (N_2310,N_2270,N_2239);
or U2311 (N_2311,N_2248,N_2253);
and U2312 (N_2312,N_2255,N_2227);
and U2313 (N_2313,N_2228,N_2268);
and U2314 (N_2314,N_2264,N_2254);
nor U2315 (N_2315,N_2259,N_2227);
nor U2316 (N_2316,N_2252,N_2263);
and U2317 (N_2317,N_2235,N_2261);
or U2318 (N_2318,N_2250,N_2264);
or U2319 (N_2319,N_2272,N_2231);
and U2320 (N_2320,N_2243,N_2239);
nand U2321 (N_2321,N_2261,N_2273);
nand U2322 (N_2322,N_2268,N_2248);
nor U2323 (N_2323,N_2222,N_2226);
or U2324 (N_2324,N_2232,N_2275);
or U2325 (N_2325,N_2263,N_2227);
or U2326 (N_2326,N_2254,N_2240);
and U2327 (N_2327,N_2268,N_2279);
nand U2328 (N_2328,N_2265,N_2269);
or U2329 (N_2329,N_2228,N_2260);
nor U2330 (N_2330,N_2262,N_2259);
nand U2331 (N_2331,N_2221,N_2253);
nor U2332 (N_2332,N_2229,N_2264);
or U2333 (N_2333,N_2242,N_2264);
nand U2334 (N_2334,N_2246,N_2261);
and U2335 (N_2335,N_2223,N_2257);
and U2336 (N_2336,N_2226,N_2230);
nand U2337 (N_2337,N_2240,N_2279);
or U2338 (N_2338,N_2269,N_2257);
or U2339 (N_2339,N_2260,N_2265);
or U2340 (N_2340,N_2284,N_2283);
nor U2341 (N_2341,N_2291,N_2312);
and U2342 (N_2342,N_2306,N_2317);
nand U2343 (N_2343,N_2339,N_2319);
or U2344 (N_2344,N_2316,N_2287);
and U2345 (N_2345,N_2322,N_2337);
and U2346 (N_2346,N_2320,N_2314);
and U2347 (N_2347,N_2336,N_2293);
nor U2348 (N_2348,N_2308,N_2289);
or U2349 (N_2349,N_2331,N_2338);
nor U2350 (N_2350,N_2315,N_2295);
nand U2351 (N_2351,N_2288,N_2285);
and U2352 (N_2352,N_2326,N_2334);
and U2353 (N_2353,N_2311,N_2333);
or U2354 (N_2354,N_2281,N_2325);
and U2355 (N_2355,N_2294,N_2332);
nand U2356 (N_2356,N_2321,N_2313);
nor U2357 (N_2357,N_2298,N_2310);
or U2358 (N_2358,N_2309,N_2304);
nand U2359 (N_2359,N_2286,N_2301);
nor U2360 (N_2360,N_2297,N_2307);
nor U2361 (N_2361,N_2323,N_2282);
nand U2362 (N_2362,N_2305,N_2299);
nor U2363 (N_2363,N_2303,N_2300);
and U2364 (N_2364,N_2328,N_2324);
nand U2365 (N_2365,N_2329,N_2292);
nand U2366 (N_2366,N_2327,N_2302);
nand U2367 (N_2367,N_2330,N_2290);
nor U2368 (N_2368,N_2318,N_2335);
nor U2369 (N_2369,N_2296,N_2280);
nand U2370 (N_2370,N_2300,N_2311);
or U2371 (N_2371,N_2325,N_2329);
nand U2372 (N_2372,N_2326,N_2336);
and U2373 (N_2373,N_2329,N_2337);
nand U2374 (N_2374,N_2297,N_2280);
or U2375 (N_2375,N_2291,N_2337);
or U2376 (N_2376,N_2331,N_2310);
or U2377 (N_2377,N_2307,N_2285);
or U2378 (N_2378,N_2290,N_2294);
or U2379 (N_2379,N_2293,N_2326);
or U2380 (N_2380,N_2308,N_2314);
or U2381 (N_2381,N_2286,N_2336);
and U2382 (N_2382,N_2314,N_2280);
and U2383 (N_2383,N_2319,N_2302);
or U2384 (N_2384,N_2293,N_2306);
and U2385 (N_2385,N_2332,N_2290);
nor U2386 (N_2386,N_2330,N_2308);
xor U2387 (N_2387,N_2295,N_2314);
or U2388 (N_2388,N_2323,N_2318);
and U2389 (N_2389,N_2310,N_2335);
nand U2390 (N_2390,N_2316,N_2338);
nor U2391 (N_2391,N_2295,N_2292);
or U2392 (N_2392,N_2311,N_2327);
nor U2393 (N_2393,N_2322,N_2316);
or U2394 (N_2394,N_2283,N_2307);
nor U2395 (N_2395,N_2333,N_2280);
nor U2396 (N_2396,N_2305,N_2284);
nor U2397 (N_2397,N_2329,N_2317);
nand U2398 (N_2398,N_2294,N_2283);
or U2399 (N_2399,N_2334,N_2304);
and U2400 (N_2400,N_2362,N_2370);
and U2401 (N_2401,N_2389,N_2394);
or U2402 (N_2402,N_2374,N_2384);
nor U2403 (N_2403,N_2364,N_2345);
and U2404 (N_2404,N_2381,N_2353);
and U2405 (N_2405,N_2359,N_2388);
or U2406 (N_2406,N_2399,N_2352);
nand U2407 (N_2407,N_2358,N_2350);
or U2408 (N_2408,N_2390,N_2349);
and U2409 (N_2409,N_2397,N_2377);
nand U2410 (N_2410,N_2396,N_2393);
and U2411 (N_2411,N_2355,N_2356);
and U2412 (N_2412,N_2398,N_2347);
and U2413 (N_2413,N_2342,N_2378);
nor U2414 (N_2414,N_2368,N_2382);
nand U2415 (N_2415,N_2340,N_2375);
nand U2416 (N_2416,N_2391,N_2361);
nand U2417 (N_2417,N_2371,N_2376);
xor U2418 (N_2418,N_2372,N_2341);
nand U2419 (N_2419,N_2357,N_2343);
nor U2420 (N_2420,N_2386,N_2383);
or U2421 (N_2421,N_2369,N_2373);
nor U2422 (N_2422,N_2367,N_2346);
or U2423 (N_2423,N_2354,N_2351);
nor U2424 (N_2424,N_2380,N_2348);
or U2425 (N_2425,N_2360,N_2365);
xnor U2426 (N_2426,N_2392,N_2385);
nand U2427 (N_2427,N_2344,N_2366);
or U2428 (N_2428,N_2387,N_2363);
nor U2429 (N_2429,N_2395,N_2379);
and U2430 (N_2430,N_2396,N_2394);
nor U2431 (N_2431,N_2394,N_2387);
nor U2432 (N_2432,N_2356,N_2379);
and U2433 (N_2433,N_2396,N_2363);
and U2434 (N_2434,N_2368,N_2359);
nand U2435 (N_2435,N_2397,N_2388);
and U2436 (N_2436,N_2379,N_2349);
or U2437 (N_2437,N_2360,N_2385);
or U2438 (N_2438,N_2351,N_2385);
nand U2439 (N_2439,N_2397,N_2346);
nand U2440 (N_2440,N_2399,N_2379);
nand U2441 (N_2441,N_2365,N_2353);
and U2442 (N_2442,N_2391,N_2348);
and U2443 (N_2443,N_2377,N_2356);
and U2444 (N_2444,N_2342,N_2371);
xnor U2445 (N_2445,N_2387,N_2395);
nor U2446 (N_2446,N_2375,N_2351);
nand U2447 (N_2447,N_2364,N_2353);
nand U2448 (N_2448,N_2356,N_2388);
nand U2449 (N_2449,N_2340,N_2389);
or U2450 (N_2450,N_2347,N_2394);
and U2451 (N_2451,N_2381,N_2388);
nand U2452 (N_2452,N_2388,N_2390);
and U2453 (N_2453,N_2364,N_2362);
and U2454 (N_2454,N_2383,N_2387);
and U2455 (N_2455,N_2364,N_2372);
nand U2456 (N_2456,N_2359,N_2398);
or U2457 (N_2457,N_2385,N_2383);
and U2458 (N_2458,N_2346,N_2352);
or U2459 (N_2459,N_2387,N_2399);
or U2460 (N_2460,N_2406,N_2454);
nand U2461 (N_2461,N_2427,N_2423);
or U2462 (N_2462,N_2441,N_2413);
nand U2463 (N_2463,N_2448,N_2402);
or U2464 (N_2464,N_2434,N_2449);
nand U2465 (N_2465,N_2405,N_2401);
and U2466 (N_2466,N_2424,N_2430);
and U2467 (N_2467,N_2419,N_2439);
nor U2468 (N_2468,N_2444,N_2407);
nor U2469 (N_2469,N_2410,N_2436);
or U2470 (N_2470,N_2440,N_2403);
or U2471 (N_2471,N_2435,N_2411);
and U2472 (N_2472,N_2426,N_2409);
nor U2473 (N_2473,N_2442,N_2443);
and U2474 (N_2474,N_2455,N_2428);
or U2475 (N_2475,N_2432,N_2451);
nand U2476 (N_2476,N_2447,N_2415);
or U2477 (N_2477,N_2446,N_2404);
nor U2478 (N_2478,N_2416,N_2458);
nand U2479 (N_2479,N_2438,N_2421);
nor U2480 (N_2480,N_2456,N_2400);
nor U2481 (N_2481,N_2412,N_2452);
nor U2482 (N_2482,N_2450,N_2431);
nand U2483 (N_2483,N_2422,N_2425);
nor U2484 (N_2484,N_2437,N_2414);
and U2485 (N_2485,N_2418,N_2445);
and U2486 (N_2486,N_2429,N_2417);
nand U2487 (N_2487,N_2457,N_2408);
nor U2488 (N_2488,N_2433,N_2459);
nand U2489 (N_2489,N_2420,N_2453);
nor U2490 (N_2490,N_2448,N_2454);
and U2491 (N_2491,N_2443,N_2404);
nand U2492 (N_2492,N_2427,N_2421);
and U2493 (N_2493,N_2413,N_2405);
and U2494 (N_2494,N_2408,N_2413);
xor U2495 (N_2495,N_2440,N_2401);
nor U2496 (N_2496,N_2450,N_2444);
and U2497 (N_2497,N_2417,N_2434);
nand U2498 (N_2498,N_2451,N_2459);
or U2499 (N_2499,N_2432,N_2459);
and U2500 (N_2500,N_2442,N_2422);
nand U2501 (N_2501,N_2410,N_2433);
or U2502 (N_2502,N_2444,N_2418);
or U2503 (N_2503,N_2401,N_2458);
nand U2504 (N_2504,N_2412,N_2436);
or U2505 (N_2505,N_2448,N_2432);
and U2506 (N_2506,N_2459,N_2405);
nand U2507 (N_2507,N_2420,N_2407);
and U2508 (N_2508,N_2442,N_2401);
nand U2509 (N_2509,N_2409,N_2434);
and U2510 (N_2510,N_2401,N_2402);
nand U2511 (N_2511,N_2422,N_2429);
and U2512 (N_2512,N_2405,N_2435);
or U2513 (N_2513,N_2422,N_2428);
nor U2514 (N_2514,N_2402,N_2408);
and U2515 (N_2515,N_2426,N_2415);
nor U2516 (N_2516,N_2434,N_2443);
or U2517 (N_2517,N_2424,N_2443);
and U2518 (N_2518,N_2445,N_2441);
and U2519 (N_2519,N_2407,N_2450);
nor U2520 (N_2520,N_2517,N_2465);
nand U2521 (N_2521,N_2500,N_2466);
or U2522 (N_2522,N_2469,N_2511);
nand U2523 (N_2523,N_2488,N_2468);
nor U2524 (N_2524,N_2464,N_2504);
nor U2525 (N_2525,N_2514,N_2487);
nor U2526 (N_2526,N_2478,N_2502);
or U2527 (N_2527,N_2475,N_2507);
nor U2528 (N_2528,N_2484,N_2519);
and U2529 (N_2529,N_2479,N_2508);
nand U2530 (N_2530,N_2476,N_2472);
and U2531 (N_2531,N_2512,N_2462);
and U2532 (N_2532,N_2461,N_2505);
nor U2533 (N_2533,N_2482,N_2510);
or U2534 (N_2534,N_2483,N_2460);
nand U2535 (N_2535,N_2515,N_2489);
nor U2536 (N_2536,N_2509,N_2496);
and U2537 (N_2537,N_2471,N_2481);
and U2538 (N_2538,N_2498,N_2486);
nor U2539 (N_2539,N_2499,N_2506);
nand U2540 (N_2540,N_2491,N_2516);
or U2541 (N_2541,N_2480,N_2473);
nor U2542 (N_2542,N_2493,N_2485);
nand U2543 (N_2543,N_2518,N_2470);
nand U2544 (N_2544,N_2495,N_2503);
and U2545 (N_2545,N_2494,N_2463);
and U2546 (N_2546,N_2477,N_2492);
nor U2547 (N_2547,N_2501,N_2474);
or U2548 (N_2548,N_2490,N_2497);
nand U2549 (N_2549,N_2513,N_2467);
nor U2550 (N_2550,N_2486,N_2512);
nor U2551 (N_2551,N_2471,N_2496);
nand U2552 (N_2552,N_2499,N_2473);
nor U2553 (N_2553,N_2489,N_2502);
nand U2554 (N_2554,N_2512,N_2493);
and U2555 (N_2555,N_2480,N_2496);
or U2556 (N_2556,N_2496,N_2507);
nor U2557 (N_2557,N_2475,N_2495);
nand U2558 (N_2558,N_2495,N_2504);
and U2559 (N_2559,N_2470,N_2483);
nand U2560 (N_2560,N_2516,N_2517);
nor U2561 (N_2561,N_2472,N_2503);
nand U2562 (N_2562,N_2471,N_2501);
or U2563 (N_2563,N_2507,N_2514);
nand U2564 (N_2564,N_2468,N_2476);
nor U2565 (N_2565,N_2506,N_2488);
nor U2566 (N_2566,N_2506,N_2495);
nor U2567 (N_2567,N_2481,N_2498);
nor U2568 (N_2568,N_2461,N_2466);
and U2569 (N_2569,N_2515,N_2471);
nor U2570 (N_2570,N_2474,N_2512);
or U2571 (N_2571,N_2501,N_2472);
and U2572 (N_2572,N_2488,N_2480);
or U2573 (N_2573,N_2473,N_2479);
nor U2574 (N_2574,N_2476,N_2504);
nand U2575 (N_2575,N_2511,N_2475);
or U2576 (N_2576,N_2472,N_2497);
nor U2577 (N_2577,N_2489,N_2512);
nand U2578 (N_2578,N_2465,N_2496);
nand U2579 (N_2579,N_2486,N_2515);
nand U2580 (N_2580,N_2568,N_2536);
nor U2581 (N_2581,N_2579,N_2538);
or U2582 (N_2582,N_2540,N_2542);
or U2583 (N_2583,N_2541,N_2575);
or U2584 (N_2584,N_2535,N_2537);
or U2585 (N_2585,N_2561,N_2556);
and U2586 (N_2586,N_2576,N_2523);
nor U2587 (N_2587,N_2562,N_2552);
or U2588 (N_2588,N_2543,N_2578);
or U2589 (N_2589,N_2566,N_2573);
nand U2590 (N_2590,N_2534,N_2549);
nand U2591 (N_2591,N_2555,N_2574);
or U2592 (N_2592,N_2524,N_2539);
nand U2593 (N_2593,N_2569,N_2554);
nor U2594 (N_2594,N_2529,N_2553);
or U2595 (N_2595,N_2567,N_2558);
nand U2596 (N_2596,N_2546,N_2545);
nand U2597 (N_2597,N_2533,N_2526);
and U2598 (N_2598,N_2551,N_2559);
nor U2599 (N_2599,N_2547,N_2532);
nor U2600 (N_2600,N_2525,N_2521);
or U2601 (N_2601,N_2530,N_2564);
nor U2602 (N_2602,N_2544,N_2548);
and U2603 (N_2603,N_2577,N_2528);
or U2604 (N_2604,N_2563,N_2560);
nor U2605 (N_2605,N_2522,N_2571);
and U2606 (N_2606,N_2527,N_2570);
nand U2607 (N_2607,N_2520,N_2557);
xnor U2608 (N_2608,N_2565,N_2531);
and U2609 (N_2609,N_2550,N_2572);
and U2610 (N_2610,N_2537,N_2534);
and U2611 (N_2611,N_2537,N_2533);
nand U2612 (N_2612,N_2541,N_2538);
or U2613 (N_2613,N_2551,N_2578);
and U2614 (N_2614,N_2565,N_2551);
or U2615 (N_2615,N_2539,N_2567);
nand U2616 (N_2616,N_2522,N_2539);
and U2617 (N_2617,N_2568,N_2538);
or U2618 (N_2618,N_2532,N_2564);
nand U2619 (N_2619,N_2535,N_2571);
or U2620 (N_2620,N_2577,N_2555);
nor U2621 (N_2621,N_2539,N_2564);
or U2622 (N_2622,N_2531,N_2520);
nand U2623 (N_2623,N_2549,N_2551);
or U2624 (N_2624,N_2542,N_2579);
or U2625 (N_2625,N_2520,N_2522);
xor U2626 (N_2626,N_2538,N_2544);
and U2627 (N_2627,N_2523,N_2537);
nand U2628 (N_2628,N_2577,N_2574);
and U2629 (N_2629,N_2545,N_2533);
nand U2630 (N_2630,N_2538,N_2549);
and U2631 (N_2631,N_2530,N_2523);
nand U2632 (N_2632,N_2560,N_2571);
or U2633 (N_2633,N_2569,N_2563);
and U2634 (N_2634,N_2536,N_2549);
or U2635 (N_2635,N_2548,N_2541);
nand U2636 (N_2636,N_2546,N_2541);
nor U2637 (N_2637,N_2522,N_2528);
or U2638 (N_2638,N_2560,N_2541);
nor U2639 (N_2639,N_2573,N_2559);
or U2640 (N_2640,N_2614,N_2582);
and U2641 (N_2641,N_2620,N_2587);
or U2642 (N_2642,N_2595,N_2622);
and U2643 (N_2643,N_2583,N_2591);
and U2644 (N_2644,N_2608,N_2633);
nand U2645 (N_2645,N_2600,N_2586);
or U2646 (N_2646,N_2590,N_2598);
and U2647 (N_2647,N_2631,N_2592);
or U2648 (N_2648,N_2637,N_2638);
or U2649 (N_2649,N_2635,N_2636);
or U2650 (N_2650,N_2619,N_2606);
nor U2651 (N_2651,N_2597,N_2639);
nand U2652 (N_2652,N_2613,N_2585);
nand U2653 (N_2653,N_2621,N_2623);
nand U2654 (N_2654,N_2609,N_2610);
nor U2655 (N_2655,N_2581,N_2612);
nor U2656 (N_2656,N_2627,N_2615);
nor U2657 (N_2657,N_2628,N_2632);
nor U2658 (N_2658,N_2634,N_2601);
nand U2659 (N_2659,N_2604,N_2630);
nand U2660 (N_2660,N_2580,N_2607);
nand U2661 (N_2661,N_2624,N_2596);
and U2662 (N_2662,N_2611,N_2626);
and U2663 (N_2663,N_2588,N_2616);
nor U2664 (N_2664,N_2584,N_2625);
or U2665 (N_2665,N_2599,N_2594);
or U2666 (N_2666,N_2593,N_2618);
or U2667 (N_2667,N_2629,N_2617);
nand U2668 (N_2668,N_2605,N_2602);
and U2669 (N_2669,N_2589,N_2603);
nand U2670 (N_2670,N_2608,N_2622);
or U2671 (N_2671,N_2585,N_2638);
or U2672 (N_2672,N_2595,N_2621);
nand U2673 (N_2673,N_2610,N_2584);
nand U2674 (N_2674,N_2630,N_2624);
nand U2675 (N_2675,N_2588,N_2590);
nand U2676 (N_2676,N_2613,N_2638);
nor U2677 (N_2677,N_2602,N_2599);
and U2678 (N_2678,N_2589,N_2615);
or U2679 (N_2679,N_2615,N_2637);
and U2680 (N_2680,N_2639,N_2605);
and U2681 (N_2681,N_2604,N_2612);
or U2682 (N_2682,N_2623,N_2619);
and U2683 (N_2683,N_2595,N_2626);
or U2684 (N_2684,N_2593,N_2619);
nand U2685 (N_2685,N_2616,N_2590);
nand U2686 (N_2686,N_2630,N_2600);
or U2687 (N_2687,N_2612,N_2618);
nor U2688 (N_2688,N_2635,N_2628);
nor U2689 (N_2689,N_2633,N_2620);
nand U2690 (N_2690,N_2616,N_2626);
or U2691 (N_2691,N_2601,N_2593);
nand U2692 (N_2692,N_2634,N_2614);
or U2693 (N_2693,N_2612,N_2630);
nor U2694 (N_2694,N_2582,N_2635);
and U2695 (N_2695,N_2625,N_2627);
nor U2696 (N_2696,N_2586,N_2620);
nor U2697 (N_2697,N_2625,N_2620);
nor U2698 (N_2698,N_2625,N_2619);
or U2699 (N_2699,N_2608,N_2605);
nand U2700 (N_2700,N_2659,N_2680);
nor U2701 (N_2701,N_2673,N_2686);
nand U2702 (N_2702,N_2660,N_2689);
or U2703 (N_2703,N_2646,N_2641);
nor U2704 (N_2704,N_2674,N_2640);
or U2705 (N_2705,N_2649,N_2669);
nand U2706 (N_2706,N_2672,N_2655);
or U2707 (N_2707,N_2682,N_2687);
and U2708 (N_2708,N_2652,N_2657);
or U2709 (N_2709,N_2698,N_2685);
nand U2710 (N_2710,N_2661,N_2642);
nor U2711 (N_2711,N_2694,N_2654);
and U2712 (N_2712,N_2650,N_2692);
nor U2713 (N_2713,N_2677,N_2697);
or U2714 (N_2714,N_2651,N_2671);
and U2715 (N_2715,N_2678,N_2648);
and U2716 (N_2716,N_2667,N_2647);
nand U2717 (N_2717,N_2644,N_2681);
nor U2718 (N_2718,N_2658,N_2664);
nor U2719 (N_2719,N_2670,N_2663);
xor U2720 (N_2720,N_2643,N_2695);
or U2721 (N_2721,N_2693,N_2696);
or U2722 (N_2722,N_2662,N_2665);
and U2723 (N_2723,N_2653,N_2666);
nor U2724 (N_2724,N_2688,N_2668);
or U2725 (N_2725,N_2656,N_2679);
nor U2726 (N_2726,N_2676,N_2675);
or U2727 (N_2727,N_2699,N_2645);
nor U2728 (N_2728,N_2690,N_2684);
nand U2729 (N_2729,N_2683,N_2691);
or U2730 (N_2730,N_2691,N_2674);
or U2731 (N_2731,N_2694,N_2662);
and U2732 (N_2732,N_2649,N_2650);
and U2733 (N_2733,N_2665,N_2681);
nor U2734 (N_2734,N_2692,N_2671);
or U2735 (N_2735,N_2677,N_2689);
nor U2736 (N_2736,N_2693,N_2690);
or U2737 (N_2737,N_2671,N_2654);
nand U2738 (N_2738,N_2682,N_2667);
nor U2739 (N_2739,N_2668,N_2641);
nor U2740 (N_2740,N_2679,N_2689);
nor U2741 (N_2741,N_2668,N_2693);
nor U2742 (N_2742,N_2695,N_2659);
nand U2743 (N_2743,N_2646,N_2691);
nand U2744 (N_2744,N_2650,N_2642);
and U2745 (N_2745,N_2680,N_2646);
or U2746 (N_2746,N_2675,N_2646);
nand U2747 (N_2747,N_2664,N_2665);
nand U2748 (N_2748,N_2658,N_2644);
or U2749 (N_2749,N_2649,N_2684);
nand U2750 (N_2750,N_2663,N_2666);
xor U2751 (N_2751,N_2673,N_2641);
and U2752 (N_2752,N_2684,N_2640);
nand U2753 (N_2753,N_2653,N_2660);
nand U2754 (N_2754,N_2697,N_2682);
xnor U2755 (N_2755,N_2654,N_2642);
nand U2756 (N_2756,N_2685,N_2647);
and U2757 (N_2757,N_2661,N_2646);
nand U2758 (N_2758,N_2674,N_2642);
or U2759 (N_2759,N_2656,N_2650);
and U2760 (N_2760,N_2722,N_2701);
nor U2761 (N_2761,N_2725,N_2740);
or U2762 (N_2762,N_2750,N_2723);
nor U2763 (N_2763,N_2729,N_2720);
and U2764 (N_2764,N_2742,N_2724);
or U2765 (N_2765,N_2708,N_2709);
and U2766 (N_2766,N_2739,N_2721);
or U2767 (N_2767,N_2759,N_2706);
nor U2768 (N_2768,N_2751,N_2733);
or U2769 (N_2769,N_2703,N_2714);
nand U2770 (N_2770,N_2713,N_2758);
nand U2771 (N_2771,N_2704,N_2746);
nor U2772 (N_2772,N_2741,N_2726);
nand U2773 (N_2773,N_2702,N_2748);
nand U2774 (N_2774,N_2744,N_2752);
nand U2775 (N_2775,N_2754,N_2738);
nor U2776 (N_2776,N_2727,N_2700);
nor U2777 (N_2777,N_2707,N_2728);
and U2778 (N_2778,N_2756,N_2743);
or U2779 (N_2779,N_2717,N_2749);
or U2780 (N_2780,N_2716,N_2712);
nor U2781 (N_2781,N_2719,N_2747);
nand U2782 (N_2782,N_2734,N_2718);
or U2783 (N_2783,N_2735,N_2755);
nand U2784 (N_2784,N_2705,N_2731);
nand U2785 (N_2785,N_2715,N_2736);
nand U2786 (N_2786,N_2757,N_2753);
nor U2787 (N_2787,N_2732,N_2745);
nor U2788 (N_2788,N_2711,N_2710);
and U2789 (N_2789,N_2737,N_2730);
nor U2790 (N_2790,N_2744,N_2757);
and U2791 (N_2791,N_2741,N_2704);
and U2792 (N_2792,N_2712,N_2714);
nand U2793 (N_2793,N_2739,N_2710);
and U2794 (N_2794,N_2743,N_2702);
or U2795 (N_2795,N_2726,N_2743);
nor U2796 (N_2796,N_2734,N_2713);
nor U2797 (N_2797,N_2746,N_2718);
or U2798 (N_2798,N_2726,N_2747);
and U2799 (N_2799,N_2754,N_2719);
and U2800 (N_2800,N_2759,N_2711);
and U2801 (N_2801,N_2746,N_2709);
nor U2802 (N_2802,N_2702,N_2750);
and U2803 (N_2803,N_2727,N_2713);
or U2804 (N_2804,N_2746,N_2752);
and U2805 (N_2805,N_2753,N_2706);
or U2806 (N_2806,N_2754,N_2744);
or U2807 (N_2807,N_2743,N_2720);
and U2808 (N_2808,N_2733,N_2721);
and U2809 (N_2809,N_2707,N_2742);
and U2810 (N_2810,N_2743,N_2752);
nand U2811 (N_2811,N_2715,N_2707);
or U2812 (N_2812,N_2718,N_2757);
or U2813 (N_2813,N_2732,N_2710);
nand U2814 (N_2814,N_2703,N_2737);
nand U2815 (N_2815,N_2721,N_2754);
nor U2816 (N_2816,N_2731,N_2752);
or U2817 (N_2817,N_2744,N_2742);
and U2818 (N_2818,N_2720,N_2741);
or U2819 (N_2819,N_2753,N_2728);
or U2820 (N_2820,N_2774,N_2817);
or U2821 (N_2821,N_2784,N_2786);
and U2822 (N_2822,N_2787,N_2810);
nand U2823 (N_2823,N_2760,N_2788);
nor U2824 (N_2824,N_2778,N_2780);
nor U2825 (N_2825,N_2804,N_2792);
or U2826 (N_2826,N_2776,N_2806);
or U2827 (N_2827,N_2799,N_2763);
or U2828 (N_2828,N_2771,N_2807);
and U2829 (N_2829,N_2764,N_2793);
or U2830 (N_2830,N_2781,N_2785);
nor U2831 (N_2831,N_2800,N_2766);
or U2832 (N_2832,N_2791,N_2815);
and U2833 (N_2833,N_2775,N_2762);
nor U2834 (N_2834,N_2801,N_2818);
and U2835 (N_2835,N_2809,N_2802);
nand U2836 (N_2836,N_2814,N_2768);
nand U2837 (N_2837,N_2794,N_2819);
nor U2838 (N_2838,N_2773,N_2797);
nand U2839 (N_2839,N_2765,N_2795);
nor U2840 (N_2840,N_2798,N_2770);
nand U2841 (N_2841,N_2767,N_2789);
and U2842 (N_2842,N_2790,N_2808);
nor U2843 (N_2843,N_2796,N_2811);
or U2844 (N_2844,N_2782,N_2777);
xnor U2845 (N_2845,N_2783,N_2813);
nand U2846 (N_2846,N_2812,N_2805);
nor U2847 (N_2847,N_2761,N_2803);
nor U2848 (N_2848,N_2772,N_2769);
and U2849 (N_2849,N_2779,N_2816);
nand U2850 (N_2850,N_2788,N_2782);
and U2851 (N_2851,N_2811,N_2780);
nor U2852 (N_2852,N_2818,N_2797);
nor U2853 (N_2853,N_2802,N_2819);
and U2854 (N_2854,N_2777,N_2783);
nand U2855 (N_2855,N_2769,N_2761);
or U2856 (N_2856,N_2815,N_2776);
or U2857 (N_2857,N_2793,N_2785);
and U2858 (N_2858,N_2783,N_2792);
nand U2859 (N_2859,N_2766,N_2811);
or U2860 (N_2860,N_2797,N_2768);
nor U2861 (N_2861,N_2772,N_2767);
or U2862 (N_2862,N_2815,N_2789);
nand U2863 (N_2863,N_2791,N_2808);
xor U2864 (N_2864,N_2795,N_2790);
nand U2865 (N_2865,N_2787,N_2814);
and U2866 (N_2866,N_2786,N_2801);
nand U2867 (N_2867,N_2801,N_2810);
nor U2868 (N_2868,N_2785,N_2769);
and U2869 (N_2869,N_2783,N_2815);
or U2870 (N_2870,N_2768,N_2818);
nand U2871 (N_2871,N_2766,N_2801);
and U2872 (N_2872,N_2807,N_2761);
nor U2873 (N_2873,N_2805,N_2787);
or U2874 (N_2874,N_2816,N_2772);
nand U2875 (N_2875,N_2768,N_2799);
or U2876 (N_2876,N_2819,N_2811);
or U2877 (N_2877,N_2779,N_2785);
nand U2878 (N_2878,N_2772,N_2779);
nor U2879 (N_2879,N_2764,N_2770);
nand U2880 (N_2880,N_2840,N_2855);
nor U2881 (N_2881,N_2874,N_2838);
nor U2882 (N_2882,N_2847,N_2863);
and U2883 (N_2883,N_2821,N_2824);
nand U2884 (N_2884,N_2825,N_2841);
and U2885 (N_2885,N_2850,N_2846);
nor U2886 (N_2886,N_2849,N_2869);
nor U2887 (N_2887,N_2853,N_2833);
nor U2888 (N_2888,N_2860,N_2848);
nor U2889 (N_2889,N_2870,N_2864);
nor U2890 (N_2890,N_2872,N_2822);
or U2891 (N_2891,N_2827,N_2879);
nand U2892 (N_2892,N_2830,N_2877);
nor U2893 (N_2893,N_2826,N_2823);
and U2894 (N_2894,N_2828,N_2842);
nand U2895 (N_2895,N_2829,N_2854);
nor U2896 (N_2896,N_2875,N_2873);
nand U2897 (N_2897,N_2834,N_2837);
nand U2898 (N_2898,N_2858,N_2862);
or U2899 (N_2899,N_2867,N_2876);
and U2900 (N_2900,N_2871,N_2843);
and U2901 (N_2901,N_2859,N_2868);
nor U2902 (N_2902,N_2851,N_2839);
or U2903 (N_2903,N_2832,N_2831);
and U2904 (N_2904,N_2865,N_2820);
nand U2905 (N_2905,N_2836,N_2866);
nand U2906 (N_2906,N_2861,N_2845);
nand U2907 (N_2907,N_2852,N_2857);
nor U2908 (N_2908,N_2856,N_2835);
nor U2909 (N_2909,N_2844,N_2878);
or U2910 (N_2910,N_2842,N_2878);
nor U2911 (N_2911,N_2828,N_2825);
or U2912 (N_2912,N_2879,N_2836);
nand U2913 (N_2913,N_2820,N_2850);
and U2914 (N_2914,N_2874,N_2835);
nor U2915 (N_2915,N_2869,N_2848);
nand U2916 (N_2916,N_2837,N_2860);
and U2917 (N_2917,N_2836,N_2857);
nand U2918 (N_2918,N_2833,N_2829);
and U2919 (N_2919,N_2870,N_2848);
and U2920 (N_2920,N_2852,N_2874);
nand U2921 (N_2921,N_2821,N_2852);
and U2922 (N_2922,N_2867,N_2851);
and U2923 (N_2923,N_2866,N_2872);
nand U2924 (N_2924,N_2863,N_2848);
nor U2925 (N_2925,N_2860,N_2859);
nand U2926 (N_2926,N_2833,N_2828);
nand U2927 (N_2927,N_2866,N_2861);
nand U2928 (N_2928,N_2875,N_2871);
nor U2929 (N_2929,N_2841,N_2853);
nor U2930 (N_2930,N_2842,N_2829);
nor U2931 (N_2931,N_2839,N_2868);
nand U2932 (N_2932,N_2832,N_2862);
and U2933 (N_2933,N_2850,N_2829);
nand U2934 (N_2934,N_2827,N_2820);
xnor U2935 (N_2935,N_2844,N_2857);
and U2936 (N_2936,N_2854,N_2878);
and U2937 (N_2937,N_2875,N_2861);
or U2938 (N_2938,N_2863,N_2827);
nor U2939 (N_2939,N_2821,N_2865);
nor U2940 (N_2940,N_2911,N_2930);
nor U2941 (N_2941,N_2884,N_2913);
nor U2942 (N_2942,N_2918,N_2882);
or U2943 (N_2943,N_2880,N_2914);
or U2944 (N_2944,N_2910,N_2932);
or U2945 (N_2945,N_2921,N_2939);
nor U2946 (N_2946,N_2909,N_2905);
and U2947 (N_2947,N_2888,N_2934);
nand U2948 (N_2948,N_2896,N_2916);
and U2949 (N_2949,N_2925,N_2899);
nor U2950 (N_2950,N_2912,N_2904);
and U2951 (N_2951,N_2903,N_2908);
and U2952 (N_2952,N_2886,N_2890);
or U2953 (N_2953,N_2900,N_2897);
and U2954 (N_2954,N_2928,N_2931);
nor U2955 (N_2955,N_2920,N_2933);
or U2956 (N_2956,N_2893,N_2902);
and U2957 (N_2957,N_2889,N_2926);
or U2958 (N_2958,N_2887,N_2901);
and U2959 (N_2959,N_2894,N_2938);
nand U2960 (N_2960,N_2898,N_2929);
or U2961 (N_2961,N_2923,N_2907);
nor U2962 (N_2962,N_2906,N_2881);
and U2963 (N_2963,N_2917,N_2937);
nand U2964 (N_2964,N_2885,N_2895);
nor U2965 (N_2965,N_2883,N_2922);
and U2966 (N_2966,N_2919,N_2936);
nor U2967 (N_2967,N_2892,N_2927);
or U2968 (N_2968,N_2924,N_2935);
nand U2969 (N_2969,N_2915,N_2891);
nand U2970 (N_2970,N_2926,N_2905);
or U2971 (N_2971,N_2908,N_2937);
nor U2972 (N_2972,N_2924,N_2910);
and U2973 (N_2973,N_2911,N_2898);
nand U2974 (N_2974,N_2881,N_2912);
and U2975 (N_2975,N_2917,N_2926);
nor U2976 (N_2976,N_2924,N_2934);
nand U2977 (N_2977,N_2889,N_2907);
nand U2978 (N_2978,N_2895,N_2921);
or U2979 (N_2979,N_2885,N_2924);
or U2980 (N_2980,N_2907,N_2933);
or U2981 (N_2981,N_2902,N_2935);
or U2982 (N_2982,N_2897,N_2903);
nor U2983 (N_2983,N_2939,N_2915);
nor U2984 (N_2984,N_2900,N_2920);
and U2985 (N_2985,N_2937,N_2935);
nor U2986 (N_2986,N_2907,N_2912);
and U2987 (N_2987,N_2882,N_2936);
and U2988 (N_2988,N_2927,N_2926);
nand U2989 (N_2989,N_2903,N_2929);
or U2990 (N_2990,N_2895,N_2934);
xor U2991 (N_2991,N_2887,N_2927);
nand U2992 (N_2992,N_2906,N_2933);
or U2993 (N_2993,N_2925,N_2897);
nand U2994 (N_2994,N_2937,N_2904);
nor U2995 (N_2995,N_2880,N_2915);
or U2996 (N_2996,N_2896,N_2897);
nand U2997 (N_2997,N_2935,N_2909);
nand U2998 (N_2998,N_2886,N_2908);
or U2999 (N_2999,N_2895,N_2881);
and UO_0 (O_0,N_2991,N_2969);
nor UO_1 (O_1,N_2997,N_2987);
and UO_2 (O_2,N_2965,N_2951);
nor UO_3 (O_3,N_2971,N_2977);
nor UO_4 (O_4,N_2981,N_2988);
nor UO_5 (O_5,N_2957,N_2975);
or UO_6 (O_6,N_2947,N_2954);
nand UO_7 (O_7,N_2983,N_2944);
or UO_8 (O_8,N_2945,N_2984);
nor UO_9 (O_9,N_2982,N_2990);
or UO_10 (O_10,N_2942,N_2953);
nor UO_11 (O_11,N_2979,N_2996);
nand UO_12 (O_12,N_2964,N_2995);
nand UO_13 (O_13,N_2943,N_2972);
nor UO_14 (O_14,N_2999,N_2986);
and UO_15 (O_15,N_2976,N_2959);
nand UO_16 (O_16,N_2998,N_2941);
nand UO_17 (O_17,N_2952,N_2989);
or UO_18 (O_18,N_2955,N_2940);
nand UO_19 (O_19,N_2960,N_2946);
and UO_20 (O_20,N_2980,N_2966);
xnor UO_21 (O_21,N_2994,N_2956);
and UO_22 (O_22,N_2949,N_2967);
or UO_23 (O_23,N_2993,N_2970);
and UO_24 (O_24,N_2962,N_2963);
or UO_25 (O_25,N_2961,N_2985);
or UO_26 (O_26,N_2948,N_2973);
nand UO_27 (O_27,N_2950,N_2968);
xnor UO_28 (O_28,N_2958,N_2974);
and UO_29 (O_29,N_2978,N_2992);
nor UO_30 (O_30,N_2968,N_2947);
nor UO_31 (O_31,N_2997,N_2946);
and UO_32 (O_32,N_2966,N_2969);
nand UO_33 (O_33,N_2980,N_2988);
or UO_34 (O_34,N_2977,N_2965);
and UO_35 (O_35,N_2984,N_2958);
or UO_36 (O_36,N_2970,N_2953);
nor UO_37 (O_37,N_2973,N_2975);
and UO_38 (O_38,N_2969,N_2959);
or UO_39 (O_39,N_2941,N_2978);
or UO_40 (O_40,N_2980,N_2998);
nor UO_41 (O_41,N_2946,N_2967);
or UO_42 (O_42,N_2980,N_2954);
nand UO_43 (O_43,N_2964,N_2958);
nor UO_44 (O_44,N_2972,N_2982);
nor UO_45 (O_45,N_2952,N_2988);
nor UO_46 (O_46,N_2970,N_2979);
and UO_47 (O_47,N_2974,N_2961);
nand UO_48 (O_48,N_2960,N_2984);
or UO_49 (O_49,N_2982,N_2995);
or UO_50 (O_50,N_2976,N_2974);
nand UO_51 (O_51,N_2961,N_2976);
nor UO_52 (O_52,N_2952,N_2972);
nand UO_53 (O_53,N_2969,N_2963);
nand UO_54 (O_54,N_2996,N_2975);
or UO_55 (O_55,N_2963,N_2951);
or UO_56 (O_56,N_2998,N_2948);
or UO_57 (O_57,N_2946,N_2965);
nand UO_58 (O_58,N_2958,N_2963);
nand UO_59 (O_59,N_2971,N_2944);
or UO_60 (O_60,N_2958,N_2997);
or UO_61 (O_61,N_2946,N_2986);
and UO_62 (O_62,N_2979,N_2977);
nand UO_63 (O_63,N_2957,N_2980);
nand UO_64 (O_64,N_2992,N_2968);
nor UO_65 (O_65,N_2996,N_2968);
nor UO_66 (O_66,N_2955,N_2998);
and UO_67 (O_67,N_2988,N_2998);
nand UO_68 (O_68,N_2955,N_2993);
nor UO_69 (O_69,N_2941,N_2954);
nor UO_70 (O_70,N_2950,N_2983);
nand UO_71 (O_71,N_2988,N_2957);
nand UO_72 (O_72,N_2992,N_2972);
or UO_73 (O_73,N_2964,N_2962);
or UO_74 (O_74,N_2949,N_2953);
or UO_75 (O_75,N_2953,N_2972);
nand UO_76 (O_76,N_2950,N_2972);
nor UO_77 (O_77,N_2975,N_2943);
nor UO_78 (O_78,N_2994,N_2973);
nor UO_79 (O_79,N_2943,N_2986);
and UO_80 (O_80,N_2978,N_2959);
nor UO_81 (O_81,N_2952,N_2987);
nor UO_82 (O_82,N_2982,N_2967);
or UO_83 (O_83,N_2952,N_2985);
or UO_84 (O_84,N_2982,N_2962);
nor UO_85 (O_85,N_2957,N_2999);
and UO_86 (O_86,N_2967,N_2940);
nand UO_87 (O_87,N_2990,N_2960);
or UO_88 (O_88,N_2991,N_2959);
and UO_89 (O_89,N_2983,N_2998);
or UO_90 (O_90,N_2963,N_2976);
nor UO_91 (O_91,N_2942,N_2956);
and UO_92 (O_92,N_2941,N_2959);
nand UO_93 (O_93,N_2975,N_2966);
nand UO_94 (O_94,N_2961,N_2989);
or UO_95 (O_95,N_2958,N_2975);
nor UO_96 (O_96,N_2942,N_2973);
and UO_97 (O_97,N_2994,N_2950);
or UO_98 (O_98,N_2991,N_2940);
or UO_99 (O_99,N_2960,N_2977);
nand UO_100 (O_100,N_2990,N_2948);
nand UO_101 (O_101,N_2981,N_2978);
nor UO_102 (O_102,N_2971,N_2958);
and UO_103 (O_103,N_2977,N_2975);
nand UO_104 (O_104,N_2967,N_2989);
or UO_105 (O_105,N_2947,N_2949);
or UO_106 (O_106,N_2990,N_2983);
nor UO_107 (O_107,N_2954,N_2946);
and UO_108 (O_108,N_2980,N_2994);
or UO_109 (O_109,N_2962,N_2996);
or UO_110 (O_110,N_2962,N_2945);
nand UO_111 (O_111,N_2958,N_2969);
and UO_112 (O_112,N_2979,N_2968);
or UO_113 (O_113,N_2977,N_2978);
and UO_114 (O_114,N_2982,N_2981);
nor UO_115 (O_115,N_2991,N_2996);
or UO_116 (O_116,N_2950,N_2952);
and UO_117 (O_117,N_2968,N_2944);
nand UO_118 (O_118,N_2979,N_2975);
xnor UO_119 (O_119,N_2986,N_2940);
or UO_120 (O_120,N_2971,N_2970);
nand UO_121 (O_121,N_2942,N_2961);
nand UO_122 (O_122,N_2981,N_2967);
nor UO_123 (O_123,N_2975,N_2947);
nand UO_124 (O_124,N_2944,N_2966);
nor UO_125 (O_125,N_2985,N_2994);
nand UO_126 (O_126,N_2975,N_2948);
and UO_127 (O_127,N_2941,N_2951);
or UO_128 (O_128,N_2943,N_2947);
or UO_129 (O_129,N_2972,N_2949);
or UO_130 (O_130,N_2990,N_2944);
and UO_131 (O_131,N_2966,N_2965);
and UO_132 (O_132,N_2967,N_2993);
or UO_133 (O_133,N_2954,N_2943);
nand UO_134 (O_134,N_2966,N_2993);
nand UO_135 (O_135,N_2979,N_2959);
nand UO_136 (O_136,N_2994,N_2990);
or UO_137 (O_137,N_2968,N_2985);
or UO_138 (O_138,N_2977,N_2974);
or UO_139 (O_139,N_2959,N_2963);
nand UO_140 (O_140,N_2961,N_2995);
nor UO_141 (O_141,N_2958,N_2945);
or UO_142 (O_142,N_2946,N_2971);
and UO_143 (O_143,N_2981,N_2973);
and UO_144 (O_144,N_2979,N_2966);
and UO_145 (O_145,N_2954,N_2992);
nand UO_146 (O_146,N_2969,N_2952);
and UO_147 (O_147,N_2994,N_2995);
nor UO_148 (O_148,N_2999,N_2972);
xor UO_149 (O_149,N_2956,N_2961);
or UO_150 (O_150,N_2947,N_2989);
and UO_151 (O_151,N_2946,N_2979);
nand UO_152 (O_152,N_2954,N_2955);
and UO_153 (O_153,N_2974,N_2980);
nand UO_154 (O_154,N_2988,N_2979);
and UO_155 (O_155,N_2976,N_2970);
or UO_156 (O_156,N_2979,N_2948);
nor UO_157 (O_157,N_2973,N_2983);
nand UO_158 (O_158,N_2955,N_2952);
and UO_159 (O_159,N_2965,N_2953);
nor UO_160 (O_160,N_2984,N_2975);
nand UO_161 (O_161,N_2956,N_2967);
and UO_162 (O_162,N_2970,N_2975);
nor UO_163 (O_163,N_2962,N_2955);
nand UO_164 (O_164,N_2990,N_2954);
or UO_165 (O_165,N_2979,N_2958);
nand UO_166 (O_166,N_2997,N_2994);
nor UO_167 (O_167,N_2959,N_2975);
nor UO_168 (O_168,N_2955,N_2981);
or UO_169 (O_169,N_2943,N_2945);
or UO_170 (O_170,N_2958,N_2940);
or UO_171 (O_171,N_2960,N_2943);
nand UO_172 (O_172,N_2992,N_2955);
nor UO_173 (O_173,N_2954,N_2949);
and UO_174 (O_174,N_2983,N_2994);
nor UO_175 (O_175,N_2952,N_2994);
nand UO_176 (O_176,N_2980,N_2992);
nor UO_177 (O_177,N_2963,N_2949);
and UO_178 (O_178,N_2977,N_2959);
nand UO_179 (O_179,N_2960,N_2968);
or UO_180 (O_180,N_2955,N_2999);
nor UO_181 (O_181,N_2975,N_2999);
and UO_182 (O_182,N_2983,N_2957);
and UO_183 (O_183,N_2985,N_2986);
nor UO_184 (O_184,N_2987,N_2963);
and UO_185 (O_185,N_2972,N_2951);
nand UO_186 (O_186,N_2946,N_2998);
nand UO_187 (O_187,N_2950,N_2992);
and UO_188 (O_188,N_2970,N_2957);
and UO_189 (O_189,N_2949,N_2979);
or UO_190 (O_190,N_2949,N_2985);
or UO_191 (O_191,N_2941,N_2999);
nor UO_192 (O_192,N_2979,N_2974);
or UO_193 (O_193,N_2990,N_2993);
nor UO_194 (O_194,N_2957,N_2968);
or UO_195 (O_195,N_2962,N_2965);
nor UO_196 (O_196,N_2973,N_2993);
and UO_197 (O_197,N_2955,N_2982);
nor UO_198 (O_198,N_2943,N_2998);
and UO_199 (O_199,N_2995,N_2966);
nor UO_200 (O_200,N_2984,N_2969);
or UO_201 (O_201,N_2969,N_2962);
nor UO_202 (O_202,N_2989,N_2975);
nor UO_203 (O_203,N_2993,N_2978);
and UO_204 (O_204,N_2967,N_2941);
nor UO_205 (O_205,N_2997,N_2989);
nor UO_206 (O_206,N_2958,N_2977);
or UO_207 (O_207,N_2953,N_2982);
nor UO_208 (O_208,N_2953,N_2955);
and UO_209 (O_209,N_2948,N_2967);
nand UO_210 (O_210,N_2946,N_2956);
and UO_211 (O_211,N_2954,N_2999);
nor UO_212 (O_212,N_2958,N_2995);
nand UO_213 (O_213,N_2953,N_2997);
or UO_214 (O_214,N_2957,N_2985);
nor UO_215 (O_215,N_2993,N_2950);
nor UO_216 (O_216,N_2942,N_2997);
xor UO_217 (O_217,N_2975,N_2942);
nor UO_218 (O_218,N_2947,N_2977);
nand UO_219 (O_219,N_2973,N_2989);
and UO_220 (O_220,N_2983,N_2979);
nand UO_221 (O_221,N_2992,N_2995);
or UO_222 (O_222,N_2980,N_2977);
nor UO_223 (O_223,N_2944,N_2984);
nor UO_224 (O_224,N_2999,N_2949);
xor UO_225 (O_225,N_2990,N_2976);
nor UO_226 (O_226,N_2943,N_2959);
nand UO_227 (O_227,N_2981,N_2979);
nor UO_228 (O_228,N_2952,N_2962);
nor UO_229 (O_229,N_2983,N_2960);
nand UO_230 (O_230,N_2997,N_2940);
nand UO_231 (O_231,N_2959,N_2953);
and UO_232 (O_232,N_2980,N_2940);
or UO_233 (O_233,N_2953,N_2977);
or UO_234 (O_234,N_2943,N_2984);
and UO_235 (O_235,N_2967,N_2951);
nor UO_236 (O_236,N_2954,N_2970);
nand UO_237 (O_237,N_2977,N_2967);
nand UO_238 (O_238,N_2951,N_2998);
and UO_239 (O_239,N_2969,N_2968);
or UO_240 (O_240,N_2992,N_2958);
nor UO_241 (O_241,N_2976,N_2958);
nand UO_242 (O_242,N_2985,N_2976);
or UO_243 (O_243,N_2987,N_2979);
nand UO_244 (O_244,N_2970,N_2987);
or UO_245 (O_245,N_2946,N_2962);
nand UO_246 (O_246,N_2983,N_2982);
nor UO_247 (O_247,N_2970,N_2948);
nand UO_248 (O_248,N_2979,N_2965);
nand UO_249 (O_249,N_2987,N_2980);
nand UO_250 (O_250,N_2955,N_2941);
nand UO_251 (O_251,N_2961,N_2952);
nor UO_252 (O_252,N_2997,N_2981);
and UO_253 (O_253,N_2960,N_2981);
or UO_254 (O_254,N_2984,N_2992);
and UO_255 (O_255,N_2960,N_2964);
or UO_256 (O_256,N_2959,N_2971);
nand UO_257 (O_257,N_2950,N_2988);
nand UO_258 (O_258,N_2982,N_2989);
nor UO_259 (O_259,N_2991,N_2978);
or UO_260 (O_260,N_2988,N_2956);
nor UO_261 (O_261,N_2982,N_2958);
and UO_262 (O_262,N_2966,N_2970);
nor UO_263 (O_263,N_2967,N_2944);
nor UO_264 (O_264,N_2994,N_2941);
and UO_265 (O_265,N_2961,N_2957);
nor UO_266 (O_266,N_2969,N_2988);
or UO_267 (O_267,N_2962,N_2970);
nor UO_268 (O_268,N_2993,N_2975);
nand UO_269 (O_269,N_2978,N_2951);
or UO_270 (O_270,N_2981,N_2987);
nand UO_271 (O_271,N_2954,N_2965);
or UO_272 (O_272,N_2968,N_2967);
nor UO_273 (O_273,N_2985,N_2979);
nand UO_274 (O_274,N_2972,N_2993);
and UO_275 (O_275,N_2947,N_2944);
and UO_276 (O_276,N_2969,N_2957);
and UO_277 (O_277,N_2960,N_2993);
and UO_278 (O_278,N_2988,N_2948);
nor UO_279 (O_279,N_2959,N_2996);
and UO_280 (O_280,N_2987,N_2991);
nand UO_281 (O_281,N_2981,N_2944);
nor UO_282 (O_282,N_2995,N_2940);
nand UO_283 (O_283,N_2993,N_2968);
nor UO_284 (O_284,N_2950,N_2995);
or UO_285 (O_285,N_2977,N_2988);
nor UO_286 (O_286,N_2985,N_2962);
and UO_287 (O_287,N_2969,N_2951);
or UO_288 (O_288,N_2940,N_2964);
or UO_289 (O_289,N_2965,N_2992);
or UO_290 (O_290,N_2960,N_2948);
and UO_291 (O_291,N_2970,N_2986);
and UO_292 (O_292,N_2972,N_2985);
or UO_293 (O_293,N_2985,N_2951);
nor UO_294 (O_294,N_2981,N_2964);
nand UO_295 (O_295,N_2954,N_2956);
and UO_296 (O_296,N_2954,N_2964);
and UO_297 (O_297,N_2941,N_2997);
nand UO_298 (O_298,N_2962,N_2983);
nand UO_299 (O_299,N_2963,N_2950);
nor UO_300 (O_300,N_2964,N_2941);
and UO_301 (O_301,N_2988,N_2949);
nand UO_302 (O_302,N_2967,N_2971);
nand UO_303 (O_303,N_2950,N_2974);
or UO_304 (O_304,N_2982,N_2980);
nand UO_305 (O_305,N_2999,N_2983);
and UO_306 (O_306,N_2952,N_2997);
or UO_307 (O_307,N_2964,N_2990);
and UO_308 (O_308,N_2955,N_2963);
nand UO_309 (O_309,N_2940,N_2984);
nor UO_310 (O_310,N_2984,N_2994);
or UO_311 (O_311,N_2968,N_2961);
nand UO_312 (O_312,N_2945,N_2951);
nor UO_313 (O_313,N_2983,N_2947);
nor UO_314 (O_314,N_2997,N_2970);
nor UO_315 (O_315,N_2981,N_2961);
nand UO_316 (O_316,N_2961,N_2987);
and UO_317 (O_317,N_2990,N_2949);
or UO_318 (O_318,N_2947,N_2956);
nand UO_319 (O_319,N_2940,N_2950);
or UO_320 (O_320,N_2962,N_2953);
or UO_321 (O_321,N_2951,N_2973);
or UO_322 (O_322,N_2946,N_2945);
nor UO_323 (O_323,N_2950,N_2981);
or UO_324 (O_324,N_2976,N_2943);
nor UO_325 (O_325,N_2971,N_2988);
nor UO_326 (O_326,N_2957,N_2955);
nand UO_327 (O_327,N_2959,N_2964);
nand UO_328 (O_328,N_2979,N_2956);
and UO_329 (O_329,N_2998,N_2971);
nor UO_330 (O_330,N_2949,N_2982);
nor UO_331 (O_331,N_2961,N_2940);
and UO_332 (O_332,N_2953,N_2968);
nand UO_333 (O_333,N_2982,N_2984);
or UO_334 (O_334,N_2986,N_2987);
and UO_335 (O_335,N_2958,N_2973);
nand UO_336 (O_336,N_2979,N_2995);
nand UO_337 (O_337,N_2987,N_2948);
or UO_338 (O_338,N_2982,N_2994);
or UO_339 (O_339,N_2946,N_2976);
or UO_340 (O_340,N_2962,N_2960);
nand UO_341 (O_341,N_2997,N_2944);
and UO_342 (O_342,N_2978,N_2965);
nand UO_343 (O_343,N_2993,N_2992);
nor UO_344 (O_344,N_2983,N_2980);
nor UO_345 (O_345,N_2970,N_2955);
nand UO_346 (O_346,N_2945,N_2979);
nor UO_347 (O_347,N_2982,N_2950);
nand UO_348 (O_348,N_2974,N_2946);
or UO_349 (O_349,N_2984,N_2947);
and UO_350 (O_350,N_2971,N_2985);
and UO_351 (O_351,N_2991,N_2952);
nor UO_352 (O_352,N_2953,N_2958);
and UO_353 (O_353,N_2996,N_2956);
and UO_354 (O_354,N_2981,N_2984);
or UO_355 (O_355,N_2967,N_2992);
or UO_356 (O_356,N_2966,N_2991);
or UO_357 (O_357,N_2960,N_2959);
and UO_358 (O_358,N_2957,N_2940);
nor UO_359 (O_359,N_2966,N_2940);
and UO_360 (O_360,N_2977,N_2968);
or UO_361 (O_361,N_2978,N_2989);
nor UO_362 (O_362,N_2964,N_2950);
or UO_363 (O_363,N_2976,N_2977);
nand UO_364 (O_364,N_2989,N_2960);
and UO_365 (O_365,N_2949,N_2962);
nand UO_366 (O_366,N_2984,N_2959);
and UO_367 (O_367,N_2950,N_2943);
or UO_368 (O_368,N_2953,N_2990);
nor UO_369 (O_369,N_2940,N_2971);
and UO_370 (O_370,N_2964,N_2979);
nand UO_371 (O_371,N_2998,N_2944);
nand UO_372 (O_372,N_2991,N_2963);
or UO_373 (O_373,N_2961,N_2997);
and UO_374 (O_374,N_2980,N_2967);
or UO_375 (O_375,N_2979,N_2952);
and UO_376 (O_376,N_2966,N_2971);
or UO_377 (O_377,N_2945,N_2968);
and UO_378 (O_378,N_2942,N_2992);
and UO_379 (O_379,N_2976,N_2972);
or UO_380 (O_380,N_2989,N_2996);
nor UO_381 (O_381,N_2955,N_2976);
nor UO_382 (O_382,N_2942,N_2998);
or UO_383 (O_383,N_2968,N_2994);
nand UO_384 (O_384,N_2963,N_2993);
nor UO_385 (O_385,N_2978,N_2949);
and UO_386 (O_386,N_2941,N_2943);
nor UO_387 (O_387,N_2983,N_2965);
or UO_388 (O_388,N_2977,N_2991);
nor UO_389 (O_389,N_2986,N_2994);
nand UO_390 (O_390,N_2976,N_2948);
nor UO_391 (O_391,N_2942,N_2990);
nor UO_392 (O_392,N_2960,N_2957);
or UO_393 (O_393,N_2985,N_2982);
and UO_394 (O_394,N_2980,N_2943);
and UO_395 (O_395,N_2953,N_2946);
nand UO_396 (O_396,N_2942,N_2995);
nand UO_397 (O_397,N_2997,N_2945);
and UO_398 (O_398,N_2972,N_2989);
nor UO_399 (O_399,N_2947,N_2957);
or UO_400 (O_400,N_2982,N_2976);
nand UO_401 (O_401,N_2942,N_2972);
nor UO_402 (O_402,N_2989,N_2991);
and UO_403 (O_403,N_2954,N_2971);
or UO_404 (O_404,N_2955,N_2959);
and UO_405 (O_405,N_2976,N_2996);
nor UO_406 (O_406,N_2948,N_2959);
and UO_407 (O_407,N_2942,N_2960);
and UO_408 (O_408,N_2944,N_2987);
nand UO_409 (O_409,N_2955,N_2989);
or UO_410 (O_410,N_2964,N_2944);
and UO_411 (O_411,N_2976,N_2965);
and UO_412 (O_412,N_2957,N_2951);
nand UO_413 (O_413,N_2953,N_2991);
and UO_414 (O_414,N_2953,N_2995);
or UO_415 (O_415,N_2948,N_2956);
and UO_416 (O_416,N_2996,N_2980);
and UO_417 (O_417,N_2982,N_2940);
and UO_418 (O_418,N_2979,N_2973);
or UO_419 (O_419,N_2978,N_2964);
nor UO_420 (O_420,N_2971,N_2981);
nor UO_421 (O_421,N_2945,N_2980);
nand UO_422 (O_422,N_2992,N_2985);
or UO_423 (O_423,N_2946,N_2996);
or UO_424 (O_424,N_2967,N_2999);
and UO_425 (O_425,N_2973,N_2980);
nor UO_426 (O_426,N_2948,N_2972);
nand UO_427 (O_427,N_2950,N_2985);
and UO_428 (O_428,N_2962,N_2978);
or UO_429 (O_429,N_2958,N_2948);
or UO_430 (O_430,N_2951,N_2944);
nor UO_431 (O_431,N_2953,N_2980);
and UO_432 (O_432,N_2940,N_2944);
or UO_433 (O_433,N_2998,N_2968);
nand UO_434 (O_434,N_2992,N_2940);
and UO_435 (O_435,N_2954,N_2952);
and UO_436 (O_436,N_2997,N_2968);
nor UO_437 (O_437,N_2947,N_2963);
nor UO_438 (O_438,N_2982,N_2973);
and UO_439 (O_439,N_2957,N_2978);
nand UO_440 (O_440,N_2976,N_2952);
nand UO_441 (O_441,N_2942,N_2951);
nand UO_442 (O_442,N_2989,N_2946);
and UO_443 (O_443,N_2995,N_2984);
nor UO_444 (O_444,N_2998,N_2986);
nor UO_445 (O_445,N_2948,N_2946);
nand UO_446 (O_446,N_2952,N_2993);
nor UO_447 (O_447,N_2956,N_2973);
and UO_448 (O_448,N_2964,N_2969);
or UO_449 (O_449,N_2944,N_2974);
or UO_450 (O_450,N_2983,N_2940);
and UO_451 (O_451,N_2981,N_2983);
nor UO_452 (O_452,N_2961,N_2990);
nor UO_453 (O_453,N_2968,N_2956);
and UO_454 (O_454,N_2992,N_2982);
or UO_455 (O_455,N_2951,N_2977);
nand UO_456 (O_456,N_2981,N_2970);
nand UO_457 (O_457,N_2995,N_2947);
nand UO_458 (O_458,N_2953,N_2969);
nand UO_459 (O_459,N_2989,N_2979);
or UO_460 (O_460,N_2943,N_2964);
and UO_461 (O_461,N_2999,N_2987);
or UO_462 (O_462,N_2998,N_2999);
and UO_463 (O_463,N_2947,N_2998);
and UO_464 (O_464,N_2948,N_2983);
xor UO_465 (O_465,N_2963,N_2973);
nor UO_466 (O_466,N_2972,N_2977);
and UO_467 (O_467,N_2979,N_2992);
and UO_468 (O_468,N_2949,N_2960);
nand UO_469 (O_469,N_2941,N_2982);
nor UO_470 (O_470,N_2942,N_2974);
nor UO_471 (O_471,N_2968,N_2999);
or UO_472 (O_472,N_2958,N_2941);
or UO_473 (O_473,N_2951,N_2984);
or UO_474 (O_474,N_2976,N_2980);
or UO_475 (O_475,N_2966,N_2977);
and UO_476 (O_476,N_2941,N_2973);
nand UO_477 (O_477,N_2993,N_2961);
nand UO_478 (O_478,N_2989,N_2969);
nor UO_479 (O_479,N_2974,N_2988);
and UO_480 (O_480,N_2956,N_2941);
or UO_481 (O_481,N_2972,N_2981);
or UO_482 (O_482,N_2971,N_2963);
nor UO_483 (O_483,N_2942,N_2991);
nor UO_484 (O_484,N_2944,N_2980);
or UO_485 (O_485,N_2947,N_2952);
or UO_486 (O_486,N_2974,N_2997);
nor UO_487 (O_487,N_2971,N_2961);
nand UO_488 (O_488,N_2966,N_2956);
and UO_489 (O_489,N_2970,N_2958);
nor UO_490 (O_490,N_2952,N_2996);
nor UO_491 (O_491,N_2974,N_2971);
nand UO_492 (O_492,N_2991,N_2974);
and UO_493 (O_493,N_2961,N_2960);
and UO_494 (O_494,N_2944,N_2963);
and UO_495 (O_495,N_2975,N_2967);
nand UO_496 (O_496,N_2945,N_2994);
and UO_497 (O_497,N_2985,N_2980);
or UO_498 (O_498,N_2989,N_2974);
and UO_499 (O_499,N_2972,N_2945);
endmodule