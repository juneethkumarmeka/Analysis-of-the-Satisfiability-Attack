module basic_1000_10000_1500_2_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5001,N_5002,N_5003,N_5004,N_5007,N_5008,N_5010,N_5012,N_5014,N_5015,N_5016,N_5017,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5029,N_5030,N_5031,N_5033,N_5034,N_5035,N_5036,N_5038,N_5041,N_5043,N_5044,N_5045,N_5047,N_5048,N_5050,N_5052,N_5053,N_5054,N_5055,N_5058,N_5059,N_5062,N_5063,N_5064,N_5067,N_5069,N_5070,N_5072,N_5075,N_5078,N_5079,N_5080,N_5081,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5091,N_5092,N_5093,N_5094,N_5095,N_5097,N_5099,N_5100,N_5101,N_5104,N_5105,N_5106,N_5107,N_5108,N_5111,N_5112,N_5113,N_5114,N_5115,N_5117,N_5118,N_5119,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5133,N_5137,N_5138,N_5139,N_5140,N_5143,N_5144,N_5145,N_5146,N_5149,N_5150,N_5151,N_5153,N_5154,N_5155,N_5157,N_5158,N_5159,N_5160,N_5162,N_5163,N_5164,N_5165,N_5168,N_5171,N_5173,N_5174,N_5175,N_5176,N_5177,N_5179,N_5180,N_5181,N_5182,N_5184,N_5186,N_5187,N_5191,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5202,N_5203,N_5204,N_5206,N_5207,N_5209,N_5210,N_5211,N_5212,N_5214,N_5217,N_5219,N_5220,N_5221,N_5222,N_5225,N_5226,N_5227,N_5229,N_5231,N_5232,N_5233,N_5237,N_5239,N_5240,N_5244,N_5247,N_5248,N_5250,N_5251,N_5257,N_5258,N_5261,N_5263,N_5265,N_5269,N_5273,N_5274,N_5275,N_5276,N_5279,N_5282,N_5284,N_5285,N_5288,N_5289,N_5291,N_5295,N_5296,N_5298,N_5299,N_5300,N_5301,N_5303,N_5304,N_5305,N_5306,N_5309,N_5310,N_5312,N_5314,N_5315,N_5317,N_5322,N_5324,N_5325,N_5328,N_5329,N_5331,N_5332,N_5334,N_5335,N_5336,N_5337,N_5338,N_5340,N_5343,N_5344,N_5347,N_5348,N_5349,N_5350,N_5352,N_5353,N_5354,N_5356,N_5357,N_5359,N_5361,N_5363,N_5364,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5373,N_5374,N_5377,N_5381,N_5382,N_5384,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5395,N_5398,N_5400,N_5401,N_5403,N_5404,N_5405,N_5406,N_5408,N_5410,N_5412,N_5414,N_5415,N_5417,N_5418,N_5419,N_5420,N_5422,N_5423,N_5425,N_5426,N_5427,N_5429,N_5430,N_5431,N_5432,N_5433,N_5439,N_5441,N_5443,N_5444,N_5446,N_5448,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5457,N_5458,N_5459,N_5460,N_5464,N_5465,N_5469,N_5470,N_5471,N_5472,N_5473,N_5476,N_5477,N_5480,N_5483,N_5485,N_5486,N_5492,N_5494,N_5495,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5508,N_5510,N_5511,N_5514,N_5518,N_5520,N_5522,N_5524,N_5525,N_5526,N_5527,N_5529,N_5531,N_5533,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5546,N_5548,N_5549,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5564,N_5565,N_5566,N_5567,N_5568,N_5570,N_5571,N_5573,N_5574,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5587,N_5589,N_5594,N_5595,N_5597,N_5599,N_5603,N_5604,N_5606,N_5608,N_5609,N_5612,N_5615,N_5616,N_5617,N_5623,N_5626,N_5629,N_5631,N_5632,N_5633,N_5634,N_5636,N_5638,N_5639,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5650,N_5651,N_5652,N_5654,N_5657,N_5659,N_5660,N_5662,N_5663,N_5664,N_5665,N_5666,N_5668,N_5669,N_5673,N_5674,N_5675,N_5677,N_5678,N_5679,N_5681,N_5682,N_5683,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5698,N_5700,N_5703,N_5705,N_5707,N_5710,N_5711,N_5713,N_5715,N_5716,N_5719,N_5720,N_5724,N_5725,N_5726,N_5727,N_5729,N_5730,N_5731,N_5732,N_5734,N_5736,N_5739,N_5741,N_5742,N_5743,N_5745,N_5746,N_5747,N_5750,N_5752,N_5753,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5768,N_5769,N_5771,N_5776,N_5778,N_5779,N_5785,N_5786,N_5787,N_5788,N_5789,N_5792,N_5794,N_5798,N_5799,N_5801,N_5803,N_5805,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5819,N_5821,N_5822,N_5823,N_5827,N_5829,N_5830,N_5832,N_5834,N_5835,N_5837,N_5838,N_5839,N_5840,N_5842,N_5843,N_5847,N_5849,N_5851,N_5853,N_5854,N_5857,N_5858,N_5859,N_5862,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5882,N_5883,N_5884,N_5885,N_5889,N_5890,N_5891,N_5894,N_5898,N_5899,N_5905,N_5906,N_5907,N_5910,N_5912,N_5914,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5926,N_5927,N_5928,N_5929,N_5931,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5940,N_5942,N_5943,N_5946,N_5947,N_5948,N_5952,N_5954,N_5957,N_5958,N_5959,N_5960,N_5962,N_5963,N_5964,N_5965,N_5971,N_5974,N_5975,N_5976,N_5977,N_5979,N_5981,N_5982,N_5988,N_5990,N_5993,N_5994,N_5997,N_5999,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6012,N_6013,N_6015,N_6016,N_6018,N_6021,N_6023,N_6024,N_6025,N_6027,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6040,N_6041,N_6044,N_6045,N_6046,N_6047,N_6050,N_6052,N_6054,N_6058,N_6059,N_6063,N_6065,N_6066,N_6068,N_6071,N_6072,N_6074,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6092,N_6093,N_6094,N_6097,N_6098,N_6099,N_6100,N_6101,N_6103,N_6109,N_6110,N_6111,N_6114,N_6115,N_6116,N_6119,N_6121,N_6123,N_6127,N_6128,N_6131,N_6132,N_6135,N_6136,N_6138,N_6139,N_6140,N_6142,N_6143,N_6148,N_6150,N_6154,N_6156,N_6158,N_6160,N_6161,N_6163,N_6166,N_6167,N_6169,N_6170,N_6173,N_6174,N_6175,N_6176,N_6179,N_6182,N_6185,N_6188,N_6192,N_6193,N_6195,N_6198,N_6202,N_6203,N_6204,N_6205,N_6208,N_6209,N_6211,N_6212,N_6214,N_6216,N_6217,N_6219,N_6221,N_6222,N_6224,N_6225,N_6226,N_6230,N_6232,N_6233,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6243,N_6244,N_6247,N_6248,N_6249,N_6251,N_6252,N_6254,N_6255,N_6256,N_6258,N_6259,N_6260,N_6262,N_6263,N_6266,N_6267,N_6268,N_6271,N_6273,N_6274,N_6276,N_6277,N_6279,N_6281,N_6282,N_6283,N_6287,N_6288,N_6289,N_6295,N_6296,N_6297,N_6298,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6309,N_6310,N_6312,N_6313,N_6314,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6326,N_6327,N_6328,N_6332,N_6335,N_6336,N_6338,N_6339,N_6340,N_6342,N_6346,N_6347,N_6349,N_6352,N_6354,N_6355,N_6363,N_6365,N_6366,N_6367,N_6371,N_6374,N_6375,N_6376,N_6377,N_6378,N_6381,N_6384,N_6386,N_6387,N_6389,N_6390,N_6391,N_6393,N_6395,N_6397,N_6398,N_6399,N_6402,N_6403,N_6404,N_6408,N_6409,N_6410,N_6412,N_6413,N_6414,N_6415,N_6416,N_6419,N_6422,N_6424,N_6430,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6440,N_6441,N_6442,N_6443,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6458,N_6459,N_6460,N_6462,N_6464,N_6465,N_6466,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6477,N_6479,N_6480,N_6482,N_6483,N_6485,N_6486,N_6487,N_6488,N_6491,N_6493,N_6494,N_6496,N_6498,N_6499,N_6500,N_6502,N_6504,N_6505,N_6508,N_6509,N_6511,N_6512,N_6514,N_6515,N_6516,N_6519,N_6520,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6534,N_6537,N_6538,N_6539,N_6540,N_6541,N_6543,N_6545,N_6546,N_6547,N_6549,N_6551,N_6553,N_6554,N_6555,N_6556,N_6557,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6568,N_6571,N_6574,N_6576,N_6577,N_6578,N_6581,N_6583,N_6584,N_6586,N_6587,N_6588,N_6589,N_6590,N_6594,N_6595,N_6596,N_6598,N_6601,N_6602,N_6604,N_6605,N_6606,N_6610,N_6611,N_6612,N_6614,N_6616,N_6617,N_6618,N_6619,N_6620,N_6628,N_6631,N_6634,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6643,N_6644,N_6645,N_6646,N_6647,N_6649,N_6651,N_6652,N_6653,N_6654,N_6656,N_6657,N_6658,N_6661,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6672,N_6673,N_6674,N_6676,N_6678,N_6679,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6689,N_6691,N_6694,N_6695,N_6698,N_6699,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6710,N_6711,N_6714,N_6717,N_6719,N_6724,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6735,N_6737,N_6738,N_6739,N_6740,N_6742,N_6743,N_6744,N_6745,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6757,N_6759,N_6761,N_6763,N_6765,N_6767,N_6770,N_6772,N_6774,N_6776,N_6777,N_6778,N_6780,N_6782,N_6783,N_6785,N_6788,N_6789,N_6790,N_6791,N_6794,N_6796,N_6798,N_6802,N_6803,N_6806,N_6807,N_6809,N_6813,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6824,N_6829,N_6830,N_6831,N_6832,N_6833,N_6835,N_6836,N_6837,N_6838,N_6840,N_6844,N_6845,N_6846,N_6850,N_6851,N_6852,N_6853,N_6855,N_6856,N_6858,N_6859,N_6862,N_6864,N_6865,N_6866,N_6868,N_6871,N_6872,N_6873,N_6874,N_6876,N_6877,N_6879,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6896,N_6897,N_6898,N_6900,N_6901,N_6902,N_6904,N_6905,N_6906,N_6910,N_6912,N_6916,N_6918,N_6920,N_6923,N_6928,N_6929,N_6930,N_6931,N_6932,N_6939,N_6940,N_6941,N_6942,N_6945,N_6948,N_6949,N_6950,N_6951,N_6959,N_6960,N_6962,N_6965,N_6967,N_6968,N_6969,N_6971,N_6973,N_6976,N_6977,N_6978,N_6979,N_6980,N_6983,N_6986,N_6987,N_6989,N_6990,N_6992,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7005,N_7006,N_7007,N_7011,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7024,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7033,N_7034,N_7037,N_7039,N_7040,N_7046,N_7047,N_7048,N_7051,N_7052,N_7053,N_7054,N_7056,N_7057,N_7058,N_7059,N_7060,N_7064,N_7066,N_7068,N_7071,N_7072,N_7077,N_7078,N_7080,N_7081,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7092,N_7093,N_7094,N_7095,N_7097,N_7098,N_7103,N_7106,N_7107,N_7109,N_7111,N_7112,N_7113,N_7114,N_7116,N_7121,N_7122,N_7123,N_7124,N_7126,N_7128,N_7129,N_7130,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7139,N_7145,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7161,N_7162,N_7165,N_7166,N_7169,N_7170,N_7172,N_7173,N_7175,N_7178,N_7182,N_7183,N_7184,N_7185,N_7186,N_7189,N_7190,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7200,N_7202,N_7207,N_7208,N_7210,N_7211,N_7213,N_7214,N_7215,N_7216,N_7217,N_7220,N_7221,N_7222,N_7223,N_7225,N_7226,N_7227,N_7228,N_7229,N_7231,N_7232,N_7233,N_7239,N_7240,N_7242,N_7244,N_7245,N_7246,N_7247,N_7248,N_7252,N_7253,N_7254,N_7257,N_7258,N_7259,N_7260,N_7263,N_7264,N_7266,N_7267,N_7269,N_7273,N_7276,N_7278,N_7280,N_7281,N_7282,N_7285,N_7286,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7299,N_7301,N_7302,N_7304,N_7305,N_7306,N_7307,N_7309,N_7310,N_7311,N_7312,N_7313,N_7315,N_7316,N_7317,N_7321,N_7322,N_7324,N_7325,N_7326,N_7329,N_7335,N_7340,N_7341,N_7342,N_7344,N_7347,N_7348,N_7349,N_7350,N_7352,N_7353,N_7356,N_7358,N_7362,N_7368,N_7370,N_7375,N_7376,N_7377,N_7378,N_7379,N_7382,N_7385,N_7386,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7398,N_7399,N_7400,N_7401,N_7402,N_7405,N_7409,N_7410,N_7411,N_7412,N_7413,N_7415,N_7416,N_7417,N_7420,N_7422,N_7423,N_7430,N_7431,N_7432,N_7433,N_7436,N_7437,N_7438,N_7439,N_7443,N_7444,N_7445,N_7448,N_7454,N_7455,N_7457,N_7458,N_7459,N_7461,N_7463,N_7467,N_7469,N_7471,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7486,N_7487,N_7488,N_7490,N_7492,N_7493,N_7495,N_7496,N_7497,N_7498,N_7499,N_7501,N_7502,N_7503,N_7505,N_7508,N_7510,N_7512,N_7513,N_7514,N_7515,N_7517,N_7519,N_7521,N_7522,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7533,N_7534,N_7537,N_7539,N_7540,N_7541,N_7543,N_7544,N_7548,N_7549,N_7550,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7560,N_7561,N_7562,N_7563,N_7564,N_7566,N_7569,N_7570,N_7572,N_7573,N_7574,N_7576,N_7578,N_7580,N_7581,N_7582,N_7583,N_7586,N_7588,N_7591,N_7592,N_7593,N_7594,N_7596,N_7598,N_7599,N_7600,N_7602,N_7604,N_7605,N_7608,N_7610,N_7614,N_7615,N_7616,N_7617,N_7618,N_7623,N_7626,N_7630,N_7636,N_7637,N_7638,N_7639,N_7641,N_7643,N_7645,N_7646,N_7648,N_7650,N_7651,N_7654,N_7655,N_7656,N_7658,N_7659,N_7660,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7669,N_7670,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7684,N_7685,N_7687,N_7688,N_7689,N_7694,N_7695,N_7696,N_7697,N_7699,N_7701,N_7702,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7715,N_7716,N_7717,N_7718,N_7721,N_7723,N_7724,N_7725,N_7726,N_7728,N_7729,N_7731,N_7732,N_7733,N_7734,N_7736,N_7738,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7749,N_7750,N_7753,N_7754,N_7756,N_7759,N_7760,N_7764,N_7766,N_7767,N_7771,N_7772,N_7773,N_7776,N_7777,N_7778,N_7780,N_7781,N_7782,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7793,N_7794,N_7796,N_7797,N_7798,N_7799,N_7803,N_7804,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7817,N_7819,N_7820,N_7821,N_7822,N_7823,N_7826,N_7828,N_7829,N_7830,N_7831,N_7832,N_7834,N_7835,N_7837,N_7838,N_7839,N_7840,N_7843,N_7844,N_7845,N_7846,N_7848,N_7849,N_7852,N_7853,N_7854,N_7855,N_7856,N_7859,N_7860,N_7866,N_7868,N_7869,N_7873,N_7874,N_7875,N_7877,N_7878,N_7879,N_7880,N_7882,N_7885,N_7886,N_7887,N_7889,N_7890,N_7891,N_7893,N_7894,N_7895,N_7896,N_7899,N_7902,N_7905,N_7906,N_7908,N_7911,N_7913,N_7914,N_7915,N_7919,N_7920,N_7921,N_7922,N_7924,N_7927,N_7928,N_7929,N_7930,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7939,N_7940,N_7941,N_7942,N_7943,N_7946,N_7948,N_7950,N_7952,N_7953,N_7954,N_7955,N_7956,N_7958,N_7960,N_7963,N_7965,N_7966,N_7970,N_7971,N_7975,N_7976,N_7977,N_7979,N_7981,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7992,N_7993,N_7995,N_7996,N_7998,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8011,N_8012,N_8017,N_8018,N_8019,N_8020,N_8022,N_8025,N_8026,N_8028,N_8030,N_8032,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8044,N_8046,N_8047,N_8049,N_8052,N_8053,N_8055,N_8056,N_8057,N_8059,N_8060,N_8061,N_8062,N_8063,N_8065,N_8067,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8088,N_8089,N_8093,N_8094,N_8095,N_8099,N_8100,N_8106,N_8107,N_8108,N_8110,N_8112,N_8114,N_8115,N_8117,N_8118,N_8119,N_8122,N_8123,N_8124,N_8126,N_8127,N_8129,N_8132,N_8134,N_8135,N_8141,N_8143,N_8147,N_8148,N_8149,N_8151,N_8152,N_8153,N_8155,N_8156,N_8158,N_8159,N_8161,N_8162,N_8164,N_8167,N_8169,N_8175,N_8177,N_8178,N_8179,N_8183,N_8184,N_8185,N_8187,N_8189,N_8190,N_8192,N_8193,N_8194,N_8195,N_8196,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8207,N_8208,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8219,N_8220,N_8222,N_8223,N_8224,N_8226,N_8227,N_8228,N_8232,N_8233,N_8234,N_8236,N_8237,N_8238,N_8241,N_8243,N_8245,N_8246,N_8247,N_8249,N_8250,N_8252,N_8254,N_8257,N_8258,N_8261,N_8262,N_8263,N_8264,N_8266,N_8268,N_8270,N_8272,N_8273,N_8276,N_8279,N_8282,N_8283,N_8284,N_8286,N_8287,N_8288,N_8289,N_8292,N_8294,N_8295,N_8296,N_8297,N_8298,N_8300,N_8302,N_8309,N_8310,N_8311,N_8312,N_8315,N_8316,N_8317,N_8321,N_8322,N_8325,N_8326,N_8329,N_8334,N_8335,N_8336,N_8337,N_8338,N_8340,N_8341,N_8342,N_8345,N_8346,N_8348,N_8351,N_8353,N_8357,N_8358,N_8361,N_8362,N_8363,N_8364,N_8366,N_8370,N_8371,N_8372,N_8374,N_8375,N_8376,N_8377,N_8379,N_8380,N_8381,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8394,N_8396,N_8397,N_8401,N_8404,N_8406,N_8407,N_8408,N_8410,N_8411,N_8412,N_8413,N_8415,N_8416,N_8417,N_8419,N_8420,N_8421,N_8423,N_8425,N_8427,N_8428,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8438,N_8441,N_8443,N_8444,N_8445,N_8448,N_8449,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8463,N_8464,N_8465,N_8466,N_8467,N_8469,N_8470,N_8473,N_8476,N_8478,N_8481,N_8482,N_8484,N_8487,N_8488,N_8489,N_8491,N_8492,N_8493,N_8495,N_8496,N_8497,N_8501,N_8502,N_8503,N_8504,N_8505,N_8508,N_8511,N_8512,N_8513,N_8514,N_8516,N_8517,N_8519,N_8520,N_8521,N_8522,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8535,N_8536,N_8539,N_8540,N_8541,N_8546,N_8547,N_8548,N_8549,N_8550,N_8553,N_8554,N_8557,N_8559,N_8560,N_8562,N_8564,N_8567,N_8568,N_8569,N_8570,N_8573,N_8574,N_8576,N_8577,N_8580,N_8584,N_8585,N_8588,N_8589,N_8590,N_8592,N_8595,N_8596,N_8597,N_8598,N_8600,N_8601,N_8603,N_8604,N_8606,N_8607,N_8608,N_8610,N_8613,N_8614,N_8616,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8627,N_8628,N_8629,N_8630,N_8635,N_8636,N_8637,N_8638,N_8639,N_8641,N_8642,N_8643,N_8645,N_8647,N_8648,N_8651,N_8652,N_8653,N_8654,N_8656,N_8657,N_8660,N_8663,N_8664,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8682,N_8683,N_8685,N_8686,N_8687,N_8690,N_8691,N_8694,N_8695,N_8696,N_8697,N_8701,N_8702,N_8703,N_8707,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8719,N_8720,N_8721,N_8724,N_8725,N_8726,N_8727,N_8728,N_8730,N_8732,N_8733,N_8737,N_8741,N_8743,N_8744,N_8745,N_8746,N_8747,N_8749,N_8753,N_8755,N_8756,N_8757,N_8758,N_8760,N_8763,N_8764,N_8765,N_8768,N_8769,N_8770,N_8772,N_8774,N_8776,N_8777,N_8778,N_8780,N_8781,N_8783,N_8784,N_8788,N_8789,N_8791,N_8795,N_8797,N_8800,N_8801,N_8802,N_8806,N_8807,N_8808,N_8810,N_8813,N_8814,N_8815,N_8817,N_8820,N_8821,N_8822,N_8823,N_8826,N_8827,N_8828,N_8829,N_8830,N_8832,N_8835,N_8837,N_8839,N_8841,N_8842,N_8844,N_8845,N_8846,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8858,N_8859,N_8860,N_8862,N_8863,N_8864,N_8865,N_8866,N_8869,N_8870,N_8871,N_8874,N_8875,N_8880,N_8881,N_8882,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8892,N_8893,N_8896,N_8897,N_8898,N_8901,N_8903,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8915,N_8917,N_8919,N_8921,N_8922,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8933,N_8934,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8949,N_8952,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8964,N_8965,N_8969,N_8970,N_8971,N_8972,N_8973,N_8975,N_8976,N_8977,N_8978,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8989,N_8990,N_8991,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_9000,N_9001,N_9002,N_9003,N_9006,N_9008,N_9009,N_9011,N_9013,N_9014,N_9015,N_9017,N_9019,N_9022,N_9023,N_9024,N_9027,N_9028,N_9029,N_9031,N_9033,N_9035,N_9036,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9046,N_9048,N_9049,N_9050,N_9053,N_9057,N_9060,N_9061,N_9062,N_9063,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9073,N_9074,N_9076,N_9078,N_9079,N_9080,N_9081,N_9083,N_9084,N_9086,N_9088,N_9089,N_9091,N_9092,N_9093,N_9095,N_9096,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9106,N_9110,N_9112,N_9114,N_9115,N_9116,N_9121,N_9125,N_9126,N_9127,N_9128,N_9131,N_9132,N_9133,N_9136,N_9138,N_9142,N_9146,N_9147,N_9148,N_9150,N_9153,N_9156,N_9158,N_9159,N_9161,N_9162,N_9164,N_9165,N_9167,N_9168,N_9169,N_9170,N_9171,N_9175,N_9176,N_9178,N_9179,N_9182,N_9183,N_9185,N_9186,N_9188,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9197,N_9199,N_9201,N_9202,N_9203,N_9204,N_9205,N_9207,N_9208,N_9210,N_9211,N_9212,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9222,N_9224,N_9226,N_9227,N_9229,N_9230,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9245,N_9247,N_9248,N_9250,N_9251,N_9253,N_9258,N_9260,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9279,N_9280,N_9281,N_9284,N_9285,N_9287,N_9289,N_9291,N_9293,N_9294,N_9295,N_9296,N_9297,N_9300,N_9302,N_9304,N_9306,N_9307,N_9309,N_9311,N_9313,N_9315,N_9318,N_9319,N_9320,N_9321,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9336,N_9337,N_9338,N_9340,N_9341,N_9342,N_9343,N_9353,N_9354,N_9357,N_9358,N_9360,N_9361,N_9363,N_9365,N_9366,N_9367,N_9372,N_9373,N_9374,N_9376,N_9377,N_9378,N_9380,N_9381,N_9382,N_9383,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9398,N_9399,N_9400,N_9403,N_9404,N_9406,N_9407,N_9410,N_9411,N_9414,N_9416,N_9417,N_9418,N_9419,N_9420,N_9424,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9437,N_9439,N_9440,N_9441,N_9442,N_9443,N_9445,N_9447,N_9450,N_9452,N_9453,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9466,N_9467,N_9469,N_9472,N_9473,N_9474,N_9475,N_9476,N_9478,N_9483,N_9485,N_9488,N_9491,N_9493,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9503,N_9504,N_9505,N_9506,N_9507,N_9510,N_9511,N_9512,N_9514,N_9515,N_9518,N_9519,N_9520,N_9522,N_9523,N_9525,N_9526,N_9527,N_9529,N_9531,N_9532,N_9533,N_9537,N_9539,N_9540,N_9542,N_9543,N_9545,N_9550,N_9553,N_9555,N_9556,N_9559,N_9561,N_9564,N_9565,N_9566,N_9568,N_9570,N_9571,N_9574,N_9578,N_9579,N_9580,N_9585,N_9586,N_9587,N_9588,N_9590,N_9593,N_9594,N_9596,N_9597,N_9599,N_9600,N_9603,N_9604,N_9605,N_9606,N_9608,N_9609,N_9610,N_9612,N_9614,N_9615,N_9617,N_9619,N_9621,N_9623,N_9627,N_9628,N_9629,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9639,N_9640,N_9641,N_9644,N_9647,N_9648,N_9650,N_9651,N_9652,N_9655,N_9656,N_9658,N_9660,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9672,N_9673,N_9674,N_9676,N_9677,N_9679,N_9682,N_9683,N_9684,N_9685,N_9687,N_9688,N_9689,N_9691,N_9692,N_9696,N_9697,N_9698,N_9700,N_9702,N_9703,N_9707,N_9709,N_9710,N_9713,N_9715,N_9716,N_9717,N_9719,N_9720,N_9722,N_9724,N_9725,N_9726,N_9727,N_9728,N_9731,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9742,N_9744,N_9745,N_9746,N_9748,N_9750,N_9751,N_9754,N_9756,N_9757,N_9761,N_9762,N_9763,N_9764,N_9766,N_9768,N_9769,N_9770,N_9773,N_9774,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9786,N_9790,N_9791,N_9794,N_9795,N_9796,N_9797,N_9799,N_9800,N_9801,N_9803,N_9805,N_9806,N_9808,N_9809,N_9810,N_9812,N_9813,N_9815,N_9817,N_9818,N_9819,N_9821,N_9822,N_9825,N_9826,N_9829,N_9830,N_9831,N_9832,N_9834,N_9836,N_9839,N_9840,N_9841,N_9842,N_9845,N_9846,N_9849,N_9852,N_9853,N_9854,N_9855,N_9858,N_9859,N_9862,N_9864,N_9865,N_9866,N_9868,N_9869,N_9871,N_9874,N_9877,N_9878,N_9879,N_9881,N_9883,N_9884,N_9888,N_9890,N_9892,N_9893,N_9894,N_9897,N_9901,N_9903,N_9904,N_9905,N_9907,N_9909,N_9910,N_9913,N_9915,N_9918,N_9921,N_9922,N_9923,N_9924,N_9925,N_9929,N_9930,N_9931,N_9932,N_9934,N_9936,N_9937,N_9938,N_9940,N_9942,N_9943,N_9947,N_9948,N_9949,N_9950,N_9952,N_9953,N_9954,N_9961,N_9964,N_9966,N_9969,N_9970,N_9971,N_9973,N_9975,N_9977,N_9979,N_9981,N_9982,N_9989,N_9992,N_9993,N_9995,N_9996,N_9997,N_9998;
or U0 (N_0,In_205,In_840);
xor U1 (N_1,In_367,In_528);
and U2 (N_2,In_799,In_723);
nand U3 (N_3,In_58,In_123);
nand U4 (N_4,In_970,In_547);
nand U5 (N_5,In_623,In_833);
xor U6 (N_6,In_867,In_654);
xnor U7 (N_7,In_685,In_604);
nor U8 (N_8,In_628,In_568);
and U9 (N_9,In_744,In_972);
or U10 (N_10,In_503,In_304);
nor U11 (N_11,In_688,In_736);
or U12 (N_12,In_35,In_324);
nor U13 (N_13,In_681,In_124);
and U14 (N_14,In_191,In_784);
or U15 (N_15,In_395,In_931);
or U16 (N_16,In_668,In_666);
and U17 (N_17,In_873,In_237);
nand U18 (N_18,In_834,In_612);
nor U19 (N_19,In_185,In_366);
or U20 (N_20,In_635,In_794);
or U21 (N_21,In_277,In_512);
xor U22 (N_22,In_886,In_861);
nor U23 (N_23,In_116,In_7);
nor U24 (N_24,In_117,In_542);
nand U25 (N_25,In_5,In_266);
nor U26 (N_26,In_167,In_54);
or U27 (N_27,In_426,In_935);
nor U28 (N_28,In_819,In_754);
or U29 (N_29,In_800,In_373);
nand U30 (N_30,In_53,In_435);
nand U31 (N_31,In_313,In_944);
or U32 (N_32,In_851,In_497);
nand U33 (N_33,In_118,In_221);
and U34 (N_34,In_998,In_383);
or U35 (N_35,In_730,In_283);
and U36 (N_36,In_918,In_753);
nor U37 (N_37,In_164,In_527);
nand U38 (N_38,In_691,In_619);
nand U39 (N_39,In_255,In_739);
or U40 (N_40,In_876,In_737);
and U41 (N_41,In_368,In_826);
nand U42 (N_42,In_274,In_8);
nor U43 (N_43,In_626,In_109);
and U44 (N_44,In_550,In_244);
xor U45 (N_45,In_504,In_564);
or U46 (N_46,In_629,In_22);
nand U47 (N_47,In_245,In_903);
xnor U48 (N_48,In_803,In_962);
and U49 (N_49,In_827,In_682);
and U50 (N_50,In_110,In_402);
or U51 (N_51,In_791,In_917);
xor U52 (N_52,In_536,In_76);
nor U53 (N_53,In_250,In_709);
nor U54 (N_54,In_427,In_584);
or U55 (N_55,In_694,In_756);
nand U56 (N_56,In_476,In_68);
nor U57 (N_57,In_136,In_956);
nand U58 (N_58,In_581,In_806);
or U59 (N_59,In_982,In_887);
and U60 (N_60,In_845,In_261);
xnor U61 (N_61,In_122,In_706);
nand U62 (N_62,In_717,In_423);
or U63 (N_63,In_922,In_3);
and U64 (N_64,In_575,In_501);
and U65 (N_65,In_872,In_543);
xnor U66 (N_66,In_186,In_967);
nor U67 (N_67,In_259,In_639);
or U68 (N_68,In_462,In_355);
xnor U69 (N_69,In_748,In_203);
or U70 (N_70,In_820,In_842);
or U71 (N_71,In_673,In_262);
nand U72 (N_72,In_987,In_847);
or U73 (N_73,In_190,In_286);
nor U74 (N_74,In_957,In_240);
xnor U75 (N_75,In_725,In_848);
nand U76 (N_76,In_986,In_620);
and U77 (N_77,In_144,In_65);
and U78 (N_78,In_537,In_170);
or U79 (N_79,In_563,In_151);
nor U80 (N_80,In_0,In_818);
xnor U81 (N_81,In_700,In_749);
and U82 (N_82,In_514,In_458);
nand U83 (N_83,In_621,In_273);
or U84 (N_84,In_624,In_541);
nor U85 (N_85,In_438,In_522);
nand U86 (N_86,In_448,In_659);
or U87 (N_87,In_38,In_822);
nor U88 (N_88,In_985,In_115);
or U89 (N_89,In_388,In_645);
xor U90 (N_90,In_429,In_150);
and U91 (N_91,In_807,In_863);
and U92 (N_92,In_415,In_450);
or U93 (N_93,In_582,In_643);
and U94 (N_94,In_686,In_390);
nand U95 (N_95,In_696,In_750);
xor U96 (N_96,In_955,In_483);
xor U97 (N_97,In_363,In_484);
nor U98 (N_98,In_31,In_162);
nand U99 (N_99,In_455,In_412);
and U100 (N_100,In_763,In_359);
and U101 (N_101,In_21,In_320);
and U102 (N_102,In_132,In_920);
or U103 (N_103,In_385,In_340);
nor U104 (N_104,In_11,In_413);
nor U105 (N_105,In_712,In_797);
or U106 (N_106,In_916,In_767);
xnor U107 (N_107,In_552,In_404);
and U108 (N_108,In_724,In_193);
nor U109 (N_109,In_958,In_731);
xor U110 (N_110,In_601,In_43);
nor U111 (N_111,In_263,In_318);
xnor U112 (N_112,In_896,In_408);
xnor U113 (N_113,In_921,In_94);
nand U114 (N_114,In_988,In_409);
nor U115 (N_115,In_276,In_439);
nand U116 (N_116,In_699,In_650);
and U117 (N_117,In_771,In_769);
xnor U118 (N_118,In_398,In_362);
and U119 (N_119,In_579,In_715);
nor U120 (N_120,In_460,In_303);
nor U121 (N_121,In_768,In_997);
nor U122 (N_122,In_816,In_344);
nor U123 (N_123,In_678,In_182);
nand U124 (N_124,In_502,In_393);
nand U125 (N_125,In_335,In_345);
xnor U126 (N_126,In_561,In_55);
and U127 (N_127,In_538,In_488);
and U128 (N_128,In_9,In_420);
nor U129 (N_129,In_328,In_209);
nor U130 (N_130,In_843,In_592);
nor U131 (N_131,In_672,In_984);
nand U132 (N_132,In_831,In_759);
or U133 (N_133,In_60,In_948);
or U134 (N_134,In_578,In_173);
xnor U135 (N_135,In_46,In_112);
nor U136 (N_136,In_285,In_312);
or U137 (N_137,In_101,In_422);
nor U138 (N_138,In_513,In_292);
or U139 (N_139,In_271,In_153);
nor U140 (N_140,In_583,In_95);
or U141 (N_141,In_296,In_437);
and U142 (N_142,In_70,In_837);
nor U143 (N_143,In_410,In_529);
nand U144 (N_144,In_128,In_86);
or U145 (N_145,In_134,In_350);
nor U146 (N_146,In_352,In_823);
or U147 (N_147,In_381,In_257);
nor U148 (N_148,In_157,In_26);
and U149 (N_149,In_801,In_486);
and U150 (N_150,In_49,In_877);
or U151 (N_151,In_18,In_379);
nor U152 (N_152,In_23,In_178);
nor U153 (N_153,In_498,In_399);
nor U154 (N_154,In_103,In_28);
and U155 (N_155,In_882,In_158);
xor U156 (N_156,In_589,In_338);
nand U157 (N_157,In_457,In_311);
and U158 (N_158,In_2,In_991);
xnor U159 (N_159,In_667,In_557);
xnor U160 (N_160,In_857,In_942);
or U161 (N_161,In_634,In_287);
or U162 (N_162,In_859,In_565);
or U163 (N_163,In_808,In_227);
nand U164 (N_164,In_39,In_156);
nand U165 (N_165,In_549,In_1);
and U166 (N_166,In_113,In_17);
nand U167 (N_167,In_378,In_539);
or U168 (N_168,In_135,In_371);
nor U169 (N_169,In_330,In_243);
nor U170 (N_170,In_632,In_297);
and U171 (N_171,In_33,In_661);
or U172 (N_172,In_792,In_323);
and U173 (N_173,In_855,In_108);
and U174 (N_174,In_499,In_199);
or U175 (N_175,In_228,In_992);
nand U176 (N_176,In_463,In_456);
or U177 (N_177,In_80,In_651);
and U178 (N_178,In_597,In_607);
and U179 (N_179,In_310,In_319);
nor U180 (N_180,In_71,In_941);
and U181 (N_181,In_198,In_434);
nor U182 (N_182,In_217,In_387);
nor U183 (N_183,In_111,In_946);
nor U184 (N_184,In_804,In_192);
nand U185 (N_185,In_82,In_279);
nand U186 (N_186,In_945,In_862);
nand U187 (N_187,In_571,In_770);
nand U188 (N_188,In_301,In_674);
or U189 (N_189,In_810,In_570);
nand U190 (N_190,In_252,In_614);
or U191 (N_191,In_331,In_937);
or U192 (N_192,In_644,In_779);
xnor U193 (N_193,In_953,In_690);
nor U194 (N_194,In_743,In_594);
xnor U195 (N_195,In_927,In_93);
nand U196 (N_196,In_468,In_722);
and U197 (N_197,In_732,In_159);
and U198 (N_198,In_919,In_411);
and U199 (N_199,In_47,In_817);
xnor U200 (N_200,In_852,In_990);
and U201 (N_201,In_346,In_99);
xnor U202 (N_202,In_971,In_692);
xnor U203 (N_203,In_459,In_610);
and U204 (N_204,In_289,In_830);
nor U205 (N_205,In_545,In_174);
xnor U206 (N_206,In_683,In_631);
nand U207 (N_207,In_41,In_881);
xor U208 (N_208,In_711,In_264);
nand U209 (N_209,In_532,In_442);
nand U210 (N_210,In_306,In_965);
xor U211 (N_211,In_361,In_906);
nor U212 (N_212,In_234,In_374);
nand U213 (N_213,In_235,In_689);
and U214 (N_214,In_671,In_451);
nand U215 (N_215,In_684,In_447);
and U216 (N_216,In_471,In_663);
or U217 (N_217,In_977,In_850);
nand U218 (N_218,In_282,In_148);
or U219 (N_219,In_787,In_485);
and U220 (N_220,In_161,In_87);
and U221 (N_221,In_389,In_670);
xnor U222 (N_222,In_32,In_983);
or U223 (N_223,In_464,In_652);
nor U224 (N_224,In_495,In_146);
nand U225 (N_225,In_546,In_102);
nand U226 (N_226,In_675,In_846);
or U227 (N_227,In_75,In_856);
or U228 (N_228,In_835,In_492);
and U229 (N_229,In_885,In_294);
and U230 (N_230,In_633,In_288);
nand U231 (N_231,In_30,In_951);
nand U232 (N_232,In_258,In_764);
nor U233 (N_233,In_795,In_695);
xor U234 (N_234,In_392,In_637);
or U235 (N_235,In_697,In_207);
nand U236 (N_236,In_284,In_74);
and U237 (N_237,In_106,In_314);
and U238 (N_238,In_45,In_300);
and U239 (N_239,In_641,In_275);
or U240 (N_240,In_326,In_490);
and U241 (N_241,In_56,In_473);
and U242 (N_242,In_354,In_229);
and U243 (N_243,In_175,In_556);
xnor U244 (N_244,In_577,In_915);
and U245 (N_245,In_781,In_572);
nand U246 (N_246,In_278,In_206);
nor U247 (N_247,In_200,In_883);
nand U248 (N_248,In_544,In_838);
or U249 (N_249,In_445,In_421);
and U250 (N_250,In_396,In_573);
nand U251 (N_251,In_44,In_272);
nand U252 (N_252,In_531,In_220);
nand U253 (N_253,In_940,In_926);
and U254 (N_254,In_871,In_923);
xor U255 (N_255,In_976,In_69);
nand U256 (N_256,In_865,In_231);
and U257 (N_257,In_836,In_713);
nand U258 (N_258,In_617,In_305);
or U259 (N_259,In_758,In_560);
and U260 (N_260,In_980,In_138);
or U261 (N_261,In_131,In_364);
nor U262 (N_262,In_210,In_401);
nand U263 (N_263,In_85,In_786);
and U264 (N_264,In_177,In_928);
nor U265 (N_265,In_961,In_405);
or U266 (N_266,In_593,In_290);
nand U267 (N_267,In_308,In_160);
and U268 (N_268,In_246,In_27);
nor U269 (N_269,In_126,In_899);
or U270 (N_270,In_265,In_356);
nand U271 (N_271,In_718,In_932);
nor U272 (N_272,In_357,In_765);
or U273 (N_273,In_397,In_999);
nand U274 (N_274,In_40,In_790);
nand U275 (N_275,In_981,In_521);
xnor U276 (N_276,In_630,In_660);
or U277 (N_277,In_814,In_701);
nand U278 (N_278,In_576,In_444);
nor U279 (N_279,In_107,In_774);
nor U280 (N_280,In_558,In_853);
nand U281 (N_281,In_15,In_907);
or U282 (N_282,In_34,In_798);
nor U283 (N_283,In_6,In_933);
or U284 (N_284,In_888,In_567);
or U285 (N_285,In_169,In_909);
or U286 (N_286,In_716,In_525);
nand U287 (N_287,In_912,In_595);
and U288 (N_288,In_152,In_317);
or U289 (N_289,In_902,In_254);
nand U290 (N_290,In_78,In_901);
and U291 (N_291,In_465,In_219);
or U292 (N_292,In_608,In_428);
nor U293 (N_293,In_163,In_821);
or U294 (N_294,In_327,In_226);
nand U295 (N_295,In_625,In_517);
or U296 (N_296,In_555,In_469);
nor U297 (N_297,In_50,In_394);
and U298 (N_298,In_761,In_247);
xnor U299 (N_299,In_904,In_348);
and U300 (N_300,In_936,In_119);
nor U301 (N_301,In_467,In_796);
xor U302 (N_302,In_406,In_432);
nor U303 (N_303,In_510,In_656);
or U304 (N_304,In_183,In_762);
nor U305 (N_305,In_950,In_609);
and U306 (N_306,In_494,In_802);
nor U307 (N_307,In_780,In_924);
nand U308 (N_308,In_52,In_477);
and U309 (N_309,In_214,In_238);
nand U310 (N_310,In_454,In_574);
nand U311 (N_311,In_616,In_470);
xor U312 (N_312,In_993,In_196);
nor U313 (N_313,In_51,In_964);
and U314 (N_314,In_302,In_280);
nand U315 (N_315,In_251,In_664);
and U316 (N_316,In_889,In_954);
nand U317 (N_317,In_506,In_523);
or U318 (N_318,In_714,In_230);
or U319 (N_319,In_232,In_104);
nand U320 (N_320,In_98,In_487);
nor U321 (N_321,In_548,In_647);
or U322 (N_322,In_562,In_336);
nand U323 (N_323,In_751,In_704);
nand U324 (N_324,In_59,In_375);
nand U325 (N_325,In_653,In_168);
and U326 (N_326,In_24,In_519);
nand U327 (N_327,In_599,In_526);
nand U328 (N_328,In_534,In_693);
xnor U329 (N_329,In_424,In_813);
nand U330 (N_330,In_588,In_281);
or U331 (N_331,In_365,In_551);
or U332 (N_332,In_728,In_611);
nor U333 (N_333,In_491,In_97);
nand U334 (N_334,In_868,In_211);
and U335 (N_335,In_515,In_676);
nand U336 (N_336,In_782,In_745);
and U337 (N_337,In_416,In_789);
xor U338 (N_338,In_256,In_307);
nor U339 (N_339,In_493,In_914);
nor U340 (N_340,In_309,In_213);
and U341 (N_341,In_603,In_172);
and U342 (N_342,In_880,In_755);
nor U343 (N_343,In_655,In_825);
nand U344 (N_344,In_978,In_166);
and U345 (N_345,In_79,In_740);
or U346 (N_346,In_443,In_376);
nor U347 (N_347,In_248,In_478);
nand U348 (N_348,In_475,In_241);
nor U349 (N_349,In_949,In_649);
and U350 (N_350,In_341,In_194);
nor U351 (N_351,In_249,In_403);
nor U352 (N_352,In_61,In_669);
nand U353 (N_353,In_839,In_216);
nand U354 (N_354,In_295,In_64);
nor U355 (N_355,In_329,In_893);
nor U356 (N_356,In_929,In_184);
nor U357 (N_357,In_648,In_299);
nor U358 (N_358,In_453,In_530);
and U359 (N_359,In_4,In_343);
and U360 (N_360,In_947,In_569);
or U361 (N_361,In_524,In_141);
nor U362 (N_362,In_83,In_605);
nor U363 (N_363,In_14,In_721);
xnor U364 (N_364,In_640,In_37);
nor U365 (N_365,In_702,In_316);
and U366 (N_366,In_815,In_342);
or U367 (N_367,In_377,In_298);
nor U368 (N_368,In_590,In_812);
nand U369 (N_369,In_360,In_890);
or U370 (N_370,In_900,In_96);
nor U371 (N_371,In_91,In_849);
nor U372 (N_372,In_746,In_142);
xor U373 (N_373,In_875,In_864);
nand U374 (N_374,In_975,In_996);
or U375 (N_375,In_710,In_322);
and U376 (N_376,In_508,In_878);
nand U377 (N_377,In_773,In_520);
and U378 (N_378,In_910,In_995);
or U379 (N_379,In_580,In_268);
or U380 (N_380,In_165,In_12);
and U381 (N_381,In_480,In_963);
nor U382 (N_382,In_269,In_566);
nor U383 (N_383,In_425,In_67);
nand U384 (N_384,In_130,In_188);
xnor U385 (N_385,In_325,In_29);
or U386 (N_386,In_596,In_908);
or U387 (N_387,In_707,In_658);
nand U388 (N_388,In_783,In_772);
xor U389 (N_389,In_66,In_925);
or U390 (N_390,In_766,In_858);
nand U391 (N_391,In_129,In_90);
or U392 (N_392,In_73,In_417);
nor U393 (N_393,In_989,In_418);
or U394 (N_394,In_474,In_441);
nor U395 (N_395,In_727,In_979);
nor U396 (N_396,In_741,In_496);
or U397 (N_397,In_436,In_291);
xnor U398 (N_398,In_433,In_382);
xnor U399 (N_399,In_391,In_894);
and U400 (N_400,In_636,In_77);
nand U401 (N_401,In_559,In_414);
and U402 (N_402,In_260,In_380);
nor U403 (N_403,In_913,In_334);
and U404 (N_404,In_19,In_602);
and U405 (N_405,In_233,In_48);
and U406 (N_406,In_703,In_466);
nor U407 (N_407,In_63,In_898);
nor U408 (N_408,In_100,In_642);
nand U409 (N_409,In_829,In_760);
and U410 (N_410,In_89,In_705);
or U411 (N_411,In_777,In_879);
nor U412 (N_412,In_854,In_215);
nand U413 (N_413,In_500,In_752);
or U414 (N_414,In_337,In_481);
nand U415 (N_415,In_585,In_747);
or U416 (N_416,In_472,In_20);
nor U417 (N_417,In_785,In_507);
nand U418 (N_418,In_966,In_533);
or U419 (N_419,In_137,In_25);
or U420 (N_420,In_828,In_333);
nand U421 (N_421,In_618,In_905);
and U422 (N_422,In_866,In_88);
or U423 (N_423,In_776,In_180);
nor U424 (N_424,In_969,In_844);
xnor U425 (N_425,In_242,In_934);
nor U426 (N_426,In_400,In_349);
and U427 (N_427,In_236,In_824);
nand U428 (N_428,In_930,In_84);
and U429 (N_429,In_189,In_92);
and U430 (N_430,In_622,In_778);
nand U431 (N_431,In_870,In_884);
nand U432 (N_432,In_860,In_125);
nor U433 (N_433,In_218,In_479);
xor U434 (N_434,In_253,In_729);
nor U435 (N_435,In_10,In_208);
xor U436 (N_436,In_733,In_482);
nor U437 (N_437,In_638,In_179);
nand U438 (N_438,In_145,In_793);
xnor U439 (N_439,In_738,In_339);
xor U440 (N_440,In_805,In_419);
and U441 (N_441,In_742,In_891);
and U442 (N_442,In_960,In_139);
or U443 (N_443,In_293,In_133);
or U444 (N_444,In_347,In_665);
and U445 (N_445,In_449,In_351);
xor U446 (N_446,In_315,In_720);
or U447 (N_447,In_114,In_698);
nand U448 (N_448,In_187,In_222);
nor U449 (N_449,In_897,In_452);
xnor U450 (N_450,In_646,In_509);
nor U451 (N_451,In_613,In_598);
nor U452 (N_452,In_171,In_270);
or U453 (N_453,In_757,In_994);
nor U454 (N_454,In_540,In_147);
and U455 (N_455,In_657,In_708);
or U456 (N_456,In_775,In_212);
nand U457 (N_457,In_176,In_121);
nand U458 (N_458,In_952,In_505);
nand U459 (N_459,In_81,In_939);
nor U460 (N_460,In_687,In_224);
nand U461 (N_461,In_587,In_869);
and U462 (N_462,In_407,In_726);
and U463 (N_463,In_911,In_36);
or U464 (N_464,In_841,In_679);
nor U465 (N_465,In_72,In_811);
nor U466 (N_466,In_384,In_959);
or U467 (N_467,In_446,In_195);
nor U468 (N_468,In_680,In_143);
nand U469 (N_469,In_120,In_615);
or U470 (N_470,In_627,In_719);
and U471 (N_471,In_202,In_105);
nor U472 (N_472,In_430,In_461);
or U473 (N_473,In_181,In_895);
and U474 (N_474,In_968,In_223);
nand U475 (N_475,In_239,In_606);
nor U476 (N_476,In_358,In_13);
or U477 (N_477,In_267,In_511);
or U478 (N_478,In_553,In_516);
and U479 (N_479,In_440,In_372);
xor U480 (N_480,In_535,In_734);
nor U481 (N_481,In_369,In_735);
nand U482 (N_482,In_353,In_62);
nand U483 (N_483,In_974,In_518);
and U484 (N_484,In_370,In_154);
xnor U485 (N_485,In_16,In_140);
nand U486 (N_486,In_973,In_201);
or U487 (N_487,In_943,In_832);
and U488 (N_488,In_155,In_677);
or U489 (N_489,In_489,In_600);
and U490 (N_490,In_809,In_197);
and U491 (N_491,In_127,In_149);
and U492 (N_492,In_386,In_57);
nor U493 (N_493,In_321,In_662);
or U494 (N_494,In_586,In_591);
xor U495 (N_495,In_874,In_554);
or U496 (N_496,In_225,In_938);
and U497 (N_497,In_332,In_204);
xor U498 (N_498,In_892,In_788);
and U499 (N_499,In_42,In_431);
nor U500 (N_500,In_663,In_10);
or U501 (N_501,In_557,In_260);
nor U502 (N_502,In_625,In_372);
nand U503 (N_503,In_45,In_30);
and U504 (N_504,In_3,In_316);
nor U505 (N_505,In_939,In_428);
nor U506 (N_506,In_273,In_63);
nor U507 (N_507,In_751,In_411);
nand U508 (N_508,In_124,In_112);
nand U509 (N_509,In_61,In_291);
and U510 (N_510,In_282,In_831);
or U511 (N_511,In_579,In_73);
nor U512 (N_512,In_178,In_465);
or U513 (N_513,In_178,In_824);
nor U514 (N_514,In_980,In_359);
nor U515 (N_515,In_60,In_215);
nor U516 (N_516,In_437,In_863);
or U517 (N_517,In_100,In_72);
nand U518 (N_518,In_903,In_27);
and U519 (N_519,In_492,In_10);
nand U520 (N_520,In_122,In_858);
nor U521 (N_521,In_441,In_3);
and U522 (N_522,In_643,In_43);
xnor U523 (N_523,In_642,In_256);
nor U524 (N_524,In_723,In_144);
nor U525 (N_525,In_568,In_343);
nand U526 (N_526,In_122,In_183);
nor U527 (N_527,In_487,In_886);
nand U528 (N_528,In_864,In_373);
and U529 (N_529,In_775,In_337);
nand U530 (N_530,In_532,In_13);
nor U531 (N_531,In_103,In_449);
nand U532 (N_532,In_493,In_939);
nand U533 (N_533,In_512,In_970);
and U534 (N_534,In_444,In_723);
nor U535 (N_535,In_693,In_859);
xor U536 (N_536,In_296,In_38);
nor U537 (N_537,In_261,In_244);
or U538 (N_538,In_888,In_198);
and U539 (N_539,In_854,In_71);
nand U540 (N_540,In_741,In_957);
and U541 (N_541,In_288,In_514);
nor U542 (N_542,In_461,In_909);
nand U543 (N_543,In_84,In_309);
xnor U544 (N_544,In_834,In_245);
xnor U545 (N_545,In_542,In_208);
nor U546 (N_546,In_623,In_0);
and U547 (N_547,In_702,In_567);
and U548 (N_548,In_438,In_950);
nor U549 (N_549,In_53,In_850);
xor U550 (N_550,In_262,In_577);
or U551 (N_551,In_746,In_421);
nand U552 (N_552,In_466,In_465);
or U553 (N_553,In_323,In_301);
or U554 (N_554,In_673,In_206);
and U555 (N_555,In_555,In_786);
nor U556 (N_556,In_743,In_182);
and U557 (N_557,In_703,In_471);
nand U558 (N_558,In_133,In_753);
and U559 (N_559,In_902,In_492);
xor U560 (N_560,In_628,In_631);
and U561 (N_561,In_321,In_979);
and U562 (N_562,In_761,In_395);
nand U563 (N_563,In_63,In_321);
nor U564 (N_564,In_669,In_653);
nand U565 (N_565,In_102,In_184);
xor U566 (N_566,In_908,In_835);
and U567 (N_567,In_225,In_139);
nand U568 (N_568,In_714,In_447);
or U569 (N_569,In_613,In_706);
nand U570 (N_570,In_408,In_629);
nand U571 (N_571,In_209,In_446);
or U572 (N_572,In_513,In_560);
nand U573 (N_573,In_673,In_62);
nand U574 (N_574,In_942,In_624);
nor U575 (N_575,In_930,In_87);
and U576 (N_576,In_628,In_622);
nor U577 (N_577,In_959,In_130);
nor U578 (N_578,In_978,In_889);
nand U579 (N_579,In_651,In_280);
xnor U580 (N_580,In_493,In_917);
nor U581 (N_581,In_151,In_772);
or U582 (N_582,In_194,In_415);
or U583 (N_583,In_638,In_367);
or U584 (N_584,In_628,In_946);
and U585 (N_585,In_272,In_142);
and U586 (N_586,In_175,In_620);
and U587 (N_587,In_37,In_508);
nand U588 (N_588,In_173,In_228);
nand U589 (N_589,In_658,In_634);
nor U590 (N_590,In_139,In_159);
and U591 (N_591,In_117,In_22);
or U592 (N_592,In_307,In_974);
or U593 (N_593,In_996,In_492);
and U594 (N_594,In_589,In_926);
nor U595 (N_595,In_173,In_163);
and U596 (N_596,In_712,In_29);
nand U597 (N_597,In_591,In_604);
and U598 (N_598,In_784,In_247);
or U599 (N_599,In_805,In_366);
nand U600 (N_600,In_46,In_309);
nor U601 (N_601,In_836,In_32);
and U602 (N_602,In_852,In_857);
nand U603 (N_603,In_329,In_811);
nand U604 (N_604,In_889,In_490);
and U605 (N_605,In_371,In_498);
or U606 (N_606,In_232,In_361);
nand U607 (N_607,In_439,In_834);
or U608 (N_608,In_321,In_840);
nand U609 (N_609,In_245,In_361);
nand U610 (N_610,In_980,In_531);
or U611 (N_611,In_563,In_810);
nor U612 (N_612,In_27,In_293);
nand U613 (N_613,In_656,In_943);
or U614 (N_614,In_61,In_412);
or U615 (N_615,In_704,In_98);
xor U616 (N_616,In_586,In_102);
nor U617 (N_617,In_66,In_607);
and U618 (N_618,In_897,In_152);
nand U619 (N_619,In_737,In_967);
nor U620 (N_620,In_952,In_479);
or U621 (N_621,In_0,In_38);
and U622 (N_622,In_25,In_444);
nor U623 (N_623,In_689,In_926);
nand U624 (N_624,In_23,In_520);
nand U625 (N_625,In_966,In_162);
xnor U626 (N_626,In_232,In_968);
nor U627 (N_627,In_544,In_474);
nand U628 (N_628,In_930,In_567);
or U629 (N_629,In_821,In_408);
nand U630 (N_630,In_746,In_514);
or U631 (N_631,In_331,In_740);
nand U632 (N_632,In_37,In_628);
nor U633 (N_633,In_852,In_867);
nand U634 (N_634,In_883,In_900);
nand U635 (N_635,In_41,In_236);
and U636 (N_636,In_170,In_794);
nor U637 (N_637,In_650,In_595);
nand U638 (N_638,In_215,In_744);
nor U639 (N_639,In_777,In_782);
or U640 (N_640,In_652,In_88);
xor U641 (N_641,In_157,In_875);
nand U642 (N_642,In_9,In_807);
nor U643 (N_643,In_56,In_488);
or U644 (N_644,In_487,In_735);
nor U645 (N_645,In_208,In_82);
or U646 (N_646,In_529,In_54);
nand U647 (N_647,In_530,In_914);
nand U648 (N_648,In_22,In_172);
nand U649 (N_649,In_818,In_467);
nand U650 (N_650,In_858,In_37);
nor U651 (N_651,In_519,In_509);
or U652 (N_652,In_537,In_807);
nor U653 (N_653,In_359,In_387);
and U654 (N_654,In_419,In_847);
and U655 (N_655,In_981,In_226);
nand U656 (N_656,In_590,In_687);
nor U657 (N_657,In_168,In_359);
or U658 (N_658,In_636,In_658);
or U659 (N_659,In_763,In_73);
or U660 (N_660,In_940,In_905);
nor U661 (N_661,In_655,In_96);
nand U662 (N_662,In_867,In_704);
nand U663 (N_663,In_121,In_381);
nand U664 (N_664,In_963,In_694);
and U665 (N_665,In_407,In_64);
xnor U666 (N_666,In_958,In_203);
and U667 (N_667,In_492,In_106);
nor U668 (N_668,In_722,In_69);
nand U669 (N_669,In_577,In_819);
or U670 (N_670,In_150,In_968);
and U671 (N_671,In_98,In_492);
nor U672 (N_672,In_191,In_919);
or U673 (N_673,In_374,In_155);
nor U674 (N_674,In_374,In_238);
nor U675 (N_675,In_574,In_994);
or U676 (N_676,In_222,In_869);
xnor U677 (N_677,In_541,In_448);
nor U678 (N_678,In_702,In_75);
nand U679 (N_679,In_647,In_344);
and U680 (N_680,In_508,In_934);
and U681 (N_681,In_687,In_749);
or U682 (N_682,In_814,In_773);
nand U683 (N_683,In_537,In_695);
nor U684 (N_684,In_88,In_396);
nor U685 (N_685,In_170,In_621);
nand U686 (N_686,In_402,In_903);
nor U687 (N_687,In_977,In_181);
nand U688 (N_688,In_293,In_805);
or U689 (N_689,In_69,In_724);
and U690 (N_690,In_36,In_871);
xnor U691 (N_691,In_454,In_384);
nand U692 (N_692,In_617,In_202);
or U693 (N_693,In_336,In_826);
or U694 (N_694,In_482,In_381);
nor U695 (N_695,In_514,In_888);
nor U696 (N_696,In_98,In_403);
and U697 (N_697,In_859,In_40);
nand U698 (N_698,In_249,In_550);
nor U699 (N_699,In_898,In_428);
nor U700 (N_700,In_833,In_686);
and U701 (N_701,In_39,In_311);
or U702 (N_702,In_424,In_780);
and U703 (N_703,In_237,In_150);
xnor U704 (N_704,In_176,In_75);
and U705 (N_705,In_412,In_538);
nor U706 (N_706,In_270,In_110);
nand U707 (N_707,In_647,In_460);
and U708 (N_708,In_425,In_607);
nor U709 (N_709,In_93,In_257);
nor U710 (N_710,In_557,In_698);
nor U711 (N_711,In_721,In_34);
nand U712 (N_712,In_659,In_146);
nor U713 (N_713,In_961,In_515);
nor U714 (N_714,In_463,In_782);
nand U715 (N_715,In_174,In_707);
nand U716 (N_716,In_793,In_222);
nor U717 (N_717,In_529,In_872);
nor U718 (N_718,In_631,In_922);
nor U719 (N_719,In_855,In_436);
xor U720 (N_720,In_210,In_714);
and U721 (N_721,In_652,In_450);
or U722 (N_722,In_784,In_331);
nor U723 (N_723,In_450,In_731);
and U724 (N_724,In_151,In_633);
and U725 (N_725,In_507,In_566);
and U726 (N_726,In_550,In_818);
xor U727 (N_727,In_47,In_152);
nor U728 (N_728,In_596,In_780);
nand U729 (N_729,In_309,In_809);
and U730 (N_730,In_129,In_480);
or U731 (N_731,In_442,In_52);
nand U732 (N_732,In_316,In_732);
nand U733 (N_733,In_317,In_340);
nor U734 (N_734,In_926,In_410);
nor U735 (N_735,In_682,In_896);
or U736 (N_736,In_96,In_730);
or U737 (N_737,In_142,In_351);
nand U738 (N_738,In_44,In_98);
nand U739 (N_739,In_970,In_812);
and U740 (N_740,In_153,In_350);
nor U741 (N_741,In_242,In_434);
nor U742 (N_742,In_605,In_664);
or U743 (N_743,In_522,In_147);
or U744 (N_744,In_249,In_905);
or U745 (N_745,In_319,In_813);
or U746 (N_746,In_475,In_13);
xnor U747 (N_747,In_869,In_296);
or U748 (N_748,In_936,In_564);
nor U749 (N_749,In_244,In_450);
nand U750 (N_750,In_554,In_443);
nand U751 (N_751,In_278,In_875);
and U752 (N_752,In_594,In_35);
nor U753 (N_753,In_414,In_170);
nand U754 (N_754,In_292,In_377);
nand U755 (N_755,In_689,In_344);
xnor U756 (N_756,In_166,In_644);
or U757 (N_757,In_933,In_642);
nor U758 (N_758,In_494,In_217);
nor U759 (N_759,In_934,In_735);
xnor U760 (N_760,In_431,In_911);
nor U761 (N_761,In_408,In_815);
xor U762 (N_762,In_383,In_846);
nor U763 (N_763,In_785,In_612);
and U764 (N_764,In_419,In_134);
xor U765 (N_765,In_663,In_236);
or U766 (N_766,In_222,In_837);
xnor U767 (N_767,In_435,In_819);
and U768 (N_768,In_380,In_229);
and U769 (N_769,In_301,In_358);
and U770 (N_770,In_451,In_295);
or U771 (N_771,In_221,In_457);
nor U772 (N_772,In_408,In_214);
or U773 (N_773,In_519,In_612);
xor U774 (N_774,In_302,In_699);
or U775 (N_775,In_374,In_547);
xor U776 (N_776,In_710,In_966);
nor U777 (N_777,In_794,In_94);
and U778 (N_778,In_606,In_456);
or U779 (N_779,In_540,In_515);
nand U780 (N_780,In_993,In_777);
nand U781 (N_781,In_894,In_903);
and U782 (N_782,In_619,In_40);
nor U783 (N_783,In_34,In_592);
nor U784 (N_784,In_569,In_993);
or U785 (N_785,In_139,In_62);
or U786 (N_786,In_701,In_492);
nand U787 (N_787,In_799,In_396);
or U788 (N_788,In_612,In_410);
xnor U789 (N_789,In_450,In_537);
or U790 (N_790,In_253,In_195);
and U791 (N_791,In_520,In_512);
and U792 (N_792,In_102,In_218);
xor U793 (N_793,In_614,In_220);
nor U794 (N_794,In_639,In_785);
nand U795 (N_795,In_875,In_600);
nand U796 (N_796,In_900,In_606);
nor U797 (N_797,In_498,In_162);
or U798 (N_798,In_910,In_597);
nand U799 (N_799,In_625,In_971);
xor U800 (N_800,In_785,In_695);
nand U801 (N_801,In_331,In_264);
nor U802 (N_802,In_432,In_601);
or U803 (N_803,In_690,In_224);
nand U804 (N_804,In_765,In_564);
or U805 (N_805,In_942,In_864);
nor U806 (N_806,In_341,In_263);
nand U807 (N_807,In_428,In_472);
nor U808 (N_808,In_332,In_689);
nor U809 (N_809,In_501,In_489);
and U810 (N_810,In_408,In_98);
nor U811 (N_811,In_344,In_88);
and U812 (N_812,In_242,In_451);
xor U813 (N_813,In_403,In_687);
xor U814 (N_814,In_946,In_299);
nor U815 (N_815,In_339,In_699);
or U816 (N_816,In_579,In_968);
or U817 (N_817,In_731,In_840);
or U818 (N_818,In_782,In_886);
nand U819 (N_819,In_965,In_452);
nand U820 (N_820,In_774,In_907);
or U821 (N_821,In_572,In_356);
and U822 (N_822,In_940,In_770);
nor U823 (N_823,In_979,In_135);
and U824 (N_824,In_96,In_432);
and U825 (N_825,In_995,In_237);
nand U826 (N_826,In_223,In_577);
nor U827 (N_827,In_844,In_414);
or U828 (N_828,In_943,In_659);
xor U829 (N_829,In_269,In_500);
nand U830 (N_830,In_896,In_228);
or U831 (N_831,In_831,In_217);
and U832 (N_832,In_605,In_133);
nand U833 (N_833,In_919,In_719);
or U834 (N_834,In_577,In_831);
xnor U835 (N_835,In_603,In_222);
nand U836 (N_836,In_0,In_538);
or U837 (N_837,In_995,In_580);
nand U838 (N_838,In_17,In_536);
nand U839 (N_839,In_636,In_629);
and U840 (N_840,In_467,In_214);
nand U841 (N_841,In_898,In_53);
nor U842 (N_842,In_449,In_479);
xnor U843 (N_843,In_50,In_695);
and U844 (N_844,In_836,In_762);
or U845 (N_845,In_902,In_689);
and U846 (N_846,In_508,In_797);
nor U847 (N_847,In_871,In_248);
or U848 (N_848,In_477,In_297);
or U849 (N_849,In_688,In_410);
and U850 (N_850,In_177,In_649);
or U851 (N_851,In_56,In_976);
nand U852 (N_852,In_115,In_469);
nand U853 (N_853,In_740,In_908);
nand U854 (N_854,In_3,In_748);
xor U855 (N_855,In_71,In_123);
nor U856 (N_856,In_373,In_165);
and U857 (N_857,In_706,In_859);
and U858 (N_858,In_775,In_535);
nand U859 (N_859,In_369,In_269);
or U860 (N_860,In_290,In_542);
and U861 (N_861,In_814,In_460);
or U862 (N_862,In_565,In_918);
or U863 (N_863,In_381,In_422);
nand U864 (N_864,In_388,In_496);
and U865 (N_865,In_868,In_14);
and U866 (N_866,In_426,In_53);
xor U867 (N_867,In_554,In_123);
nand U868 (N_868,In_745,In_981);
and U869 (N_869,In_91,In_596);
nand U870 (N_870,In_39,In_324);
nor U871 (N_871,In_152,In_7);
xnor U872 (N_872,In_712,In_264);
nor U873 (N_873,In_1,In_554);
xor U874 (N_874,In_6,In_941);
nor U875 (N_875,In_152,In_657);
or U876 (N_876,In_865,In_705);
nor U877 (N_877,In_958,In_763);
nor U878 (N_878,In_237,In_226);
nand U879 (N_879,In_538,In_274);
nand U880 (N_880,In_824,In_746);
nor U881 (N_881,In_798,In_300);
nor U882 (N_882,In_462,In_711);
nand U883 (N_883,In_606,In_942);
or U884 (N_884,In_912,In_500);
nand U885 (N_885,In_427,In_79);
nand U886 (N_886,In_896,In_571);
nand U887 (N_887,In_100,In_29);
nor U888 (N_888,In_615,In_42);
nor U889 (N_889,In_773,In_456);
nand U890 (N_890,In_571,In_579);
and U891 (N_891,In_40,In_633);
nor U892 (N_892,In_938,In_739);
xnor U893 (N_893,In_834,In_384);
nand U894 (N_894,In_77,In_242);
or U895 (N_895,In_93,In_869);
nor U896 (N_896,In_60,In_478);
or U897 (N_897,In_154,In_994);
or U898 (N_898,In_82,In_548);
nand U899 (N_899,In_747,In_324);
and U900 (N_900,In_280,In_512);
and U901 (N_901,In_721,In_664);
nand U902 (N_902,In_118,In_610);
nor U903 (N_903,In_39,In_424);
nand U904 (N_904,In_337,In_916);
or U905 (N_905,In_455,In_55);
nor U906 (N_906,In_486,In_794);
nor U907 (N_907,In_396,In_331);
or U908 (N_908,In_425,In_945);
xnor U909 (N_909,In_623,In_951);
xor U910 (N_910,In_392,In_597);
and U911 (N_911,In_764,In_72);
nand U912 (N_912,In_458,In_946);
or U913 (N_913,In_308,In_558);
nor U914 (N_914,In_869,In_457);
nand U915 (N_915,In_689,In_470);
xor U916 (N_916,In_597,In_18);
or U917 (N_917,In_775,In_619);
or U918 (N_918,In_359,In_918);
and U919 (N_919,In_178,In_820);
nor U920 (N_920,In_154,In_611);
and U921 (N_921,In_100,In_53);
and U922 (N_922,In_458,In_47);
nand U923 (N_923,In_76,In_206);
nor U924 (N_924,In_259,In_859);
nor U925 (N_925,In_785,In_433);
xor U926 (N_926,In_121,In_464);
and U927 (N_927,In_377,In_706);
and U928 (N_928,In_167,In_200);
xor U929 (N_929,In_179,In_417);
xor U930 (N_930,In_800,In_549);
nand U931 (N_931,In_203,In_846);
nor U932 (N_932,In_249,In_8);
and U933 (N_933,In_786,In_133);
nand U934 (N_934,In_817,In_216);
nand U935 (N_935,In_406,In_967);
nand U936 (N_936,In_922,In_177);
or U937 (N_937,In_597,In_523);
and U938 (N_938,In_624,In_935);
or U939 (N_939,In_760,In_977);
and U940 (N_940,In_976,In_315);
nor U941 (N_941,In_643,In_521);
nor U942 (N_942,In_905,In_366);
or U943 (N_943,In_404,In_695);
and U944 (N_944,In_208,In_854);
or U945 (N_945,In_562,In_933);
and U946 (N_946,In_614,In_900);
nand U947 (N_947,In_254,In_419);
xnor U948 (N_948,In_449,In_330);
nand U949 (N_949,In_250,In_726);
nor U950 (N_950,In_15,In_407);
nand U951 (N_951,In_273,In_960);
nor U952 (N_952,In_701,In_746);
xnor U953 (N_953,In_359,In_329);
nor U954 (N_954,In_538,In_233);
nand U955 (N_955,In_966,In_984);
nor U956 (N_956,In_821,In_528);
or U957 (N_957,In_473,In_616);
nand U958 (N_958,In_548,In_549);
or U959 (N_959,In_379,In_873);
nor U960 (N_960,In_529,In_49);
nor U961 (N_961,In_438,In_235);
and U962 (N_962,In_749,In_43);
nand U963 (N_963,In_699,In_952);
xnor U964 (N_964,In_211,In_252);
or U965 (N_965,In_299,In_858);
nor U966 (N_966,In_410,In_479);
or U967 (N_967,In_22,In_781);
nor U968 (N_968,In_749,In_248);
nor U969 (N_969,In_982,In_876);
nor U970 (N_970,In_932,In_384);
and U971 (N_971,In_456,In_699);
and U972 (N_972,In_760,In_622);
nand U973 (N_973,In_341,In_315);
and U974 (N_974,In_667,In_158);
nand U975 (N_975,In_871,In_586);
and U976 (N_976,In_957,In_355);
xnor U977 (N_977,In_826,In_340);
nand U978 (N_978,In_693,In_658);
nor U979 (N_979,In_666,In_864);
nand U980 (N_980,In_887,In_117);
nand U981 (N_981,In_949,In_903);
nand U982 (N_982,In_357,In_469);
nand U983 (N_983,In_419,In_659);
or U984 (N_984,In_231,In_610);
or U985 (N_985,In_443,In_861);
nand U986 (N_986,In_416,In_444);
xor U987 (N_987,In_204,In_379);
or U988 (N_988,In_748,In_986);
or U989 (N_989,In_733,In_970);
and U990 (N_990,In_463,In_605);
nand U991 (N_991,In_821,In_475);
nand U992 (N_992,In_165,In_433);
nand U993 (N_993,In_461,In_333);
nand U994 (N_994,In_141,In_587);
nand U995 (N_995,In_670,In_513);
nand U996 (N_996,In_75,In_309);
nor U997 (N_997,In_879,In_230);
nor U998 (N_998,In_969,In_320);
nor U999 (N_999,In_869,In_562);
or U1000 (N_1000,In_984,In_304);
and U1001 (N_1001,In_548,In_423);
or U1002 (N_1002,In_454,In_633);
and U1003 (N_1003,In_71,In_34);
and U1004 (N_1004,In_28,In_706);
nand U1005 (N_1005,In_482,In_556);
nor U1006 (N_1006,In_853,In_420);
xor U1007 (N_1007,In_552,In_513);
nor U1008 (N_1008,In_670,In_599);
nand U1009 (N_1009,In_667,In_899);
xnor U1010 (N_1010,In_624,In_128);
or U1011 (N_1011,In_672,In_311);
nor U1012 (N_1012,In_119,In_471);
nand U1013 (N_1013,In_104,In_447);
or U1014 (N_1014,In_413,In_407);
or U1015 (N_1015,In_880,In_483);
and U1016 (N_1016,In_136,In_932);
nand U1017 (N_1017,In_586,In_234);
nand U1018 (N_1018,In_328,In_666);
xnor U1019 (N_1019,In_745,In_359);
or U1020 (N_1020,In_89,In_187);
and U1021 (N_1021,In_933,In_370);
nor U1022 (N_1022,In_658,In_452);
nand U1023 (N_1023,In_851,In_202);
and U1024 (N_1024,In_596,In_386);
and U1025 (N_1025,In_258,In_203);
nor U1026 (N_1026,In_907,In_524);
or U1027 (N_1027,In_156,In_173);
and U1028 (N_1028,In_733,In_920);
or U1029 (N_1029,In_378,In_26);
or U1030 (N_1030,In_920,In_855);
or U1031 (N_1031,In_271,In_719);
xnor U1032 (N_1032,In_327,In_153);
nand U1033 (N_1033,In_138,In_777);
xor U1034 (N_1034,In_895,In_98);
nand U1035 (N_1035,In_530,In_587);
and U1036 (N_1036,In_982,In_381);
nor U1037 (N_1037,In_163,In_996);
or U1038 (N_1038,In_962,In_607);
or U1039 (N_1039,In_263,In_236);
and U1040 (N_1040,In_302,In_202);
xor U1041 (N_1041,In_30,In_129);
nor U1042 (N_1042,In_312,In_947);
and U1043 (N_1043,In_69,In_355);
and U1044 (N_1044,In_805,In_325);
or U1045 (N_1045,In_173,In_393);
nor U1046 (N_1046,In_229,In_618);
and U1047 (N_1047,In_15,In_367);
nand U1048 (N_1048,In_455,In_495);
nor U1049 (N_1049,In_951,In_478);
nor U1050 (N_1050,In_41,In_501);
or U1051 (N_1051,In_902,In_296);
and U1052 (N_1052,In_860,In_762);
nor U1053 (N_1053,In_142,In_664);
nor U1054 (N_1054,In_400,In_175);
or U1055 (N_1055,In_672,In_691);
nor U1056 (N_1056,In_158,In_942);
nand U1057 (N_1057,In_684,In_666);
nand U1058 (N_1058,In_617,In_736);
xnor U1059 (N_1059,In_638,In_389);
nand U1060 (N_1060,In_396,In_915);
nand U1061 (N_1061,In_320,In_471);
or U1062 (N_1062,In_611,In_352);
or U1063 (N_1063,In_861,In_547);
nor U1064 (N_1064,In_499,In_47);
xnor U1065 (N_1065,In_925,In_900);
and U1066 (N_1066,In_515,In_496);
or U1067 (N_1067,In_675,In_352);
nand U1068 (N_1068,In_510,In_983);
nand U1069 (N_1069,In_872,In_424);
and U1070 (N_1070,In_855,In_774);
xnor U1071 (N_1071,In_619,In_614);
and U1072 (N_1072,In_521,In_879);
or U1073 (N_1073,In_646,In_294);
and U1074 (N_1074,In_562,In_431);
nor U1075 (N_1075,In_731,In_878);
xnor U1076 (N_1076,In_177,In_455);
or U1077 (N_1077,In_761,In_40);
or U1078 (N_1078,In_993,In_469);
or U1079 (N_1079,In_146,In_507);
or U1080 (N_1080,In_644,In_268);
and U1081 (N_1081,In_359,In_78);
or U1082 (N_1082,In_634,In_242);
and U1083 (N_1083,In_832,In_547);
nor U1084 (N_1084,In_877,In_703);
and U1085 (N_1085,In_646,In_910);
nand U1086 (N_1086,In_194,In_206);
xnor U1087 (N_1087,In_421,In_651);
nand U1088 (N_1088,In_862,In_137);
and U1089 (N_1089,In_146,In_311);
nor U1090 (N_1090,In_195,In_307);
and U1091 (N_1091,In_126,In_922);
or U1092 (N_1092,In_606,In_698);
and U1093 (N_1093,In_45,In_242);
and U1094 (N_1094,In_399,In_712);
nor U1095 (N_1095,In_122,In_218);
nand U1096 (N_1096,In_344,In_727);
and U1097 (N_1097,In_676,In_571);
nand U1098 (N_1098,In_835,In_639);
xor U1099 (N_1099,In_35,In_485);
or U1100 (N_1100,In_343,In_506);
and U1101 (N_1101,In_102,In_8);
or U1102 (N_1102,In_511,In_286);
or U1103 (N_1103,In_826,In_490);
nand U1104 (N_1104,In_399,In_914);
or U1105 (N_1105,In_272,In_984);
and U1106 (N_1106,In_248,In_748);
nor U1107 (N_1107,In_887,In_90);
nor U1108 (N_1108,In_438,In_229);
or U1109 (N_1109,In_182,In_449);
or U1110 (N_1110,In_963,In_166);
nand U1111 (N_1111,In_9,In_809);
or U1112 (N_1112,In_730,In_475);
nor U1113 (N_1113,In_775,In_173);
or U1114 (N_1114,In_802,In_32);
nand U1115 (N_1115,In_252,In_937);
or U1116 (N_1116,In_206,In_250);
xnor U1117 (N_1117,In_874,In_79);
or U1118 (N_1118,In_970,In_319);
and U1119 (N_1119,In_644,In_940);
nor U1120 (N_1120,In_112,In_147);
and U1121 (N_1121,In_992,In_308);
and U1122 (N_1122,In_75,In_131);
and U1123 (N_1123,In_431,In_464);
and U1124 (N_1124,In_370,In_39);
nand U1125 (N_1125,In_102,In_110);
nand U1126 (N_1126,In_548,In_710);
nor U1127 (N_1127,In_605,In_756);
nand U1128 (N_1128,In_944,In_366);
nand U1129 (N_1129,In_726,In_795);
or U1130 (N_1130,In_512,In_618);
nor U1131 (N_1131,In_563,In_390);
nor U1132 (N_1132,In_998,In_619);
nand U1133 (N_1133,In_241,In_766);
and U1134 (N_1134,In_118,In_649);
nor U1135 (N_1135,In_704,In_519);
nor U1136 (N_1136,In_952,In_924);
nand U1137 (N_1137,In_24,In_497);
nand U1138 (N_1138,In_616,In_304);
nand U1139 (N_1139,In_271,In_613);
nor U1140 (N_1140,In_635,In_383);
and U1141 (N_1141,In_808,In_794);
and U1142 (N_1142,In_886,In_100);
nor U1143 (N_1143,In_41,In_868);
and U1144 (N_1144,In_682,In_554);
nand U1145 (N_1145,In_454,In_935);
nand U1146 (N_1146,In_631,In_152);
or U1147 (N_1147,In_347,In_771);
nor U1148 (N_1148,In_296,In_191);
nand U1149 (N_1149,In_115,In_34);
or U1150 (N_1150,In_288,In_808);
and U1151 (N_1151,In_474,In_303);
or U1152 (N_1152,In_594,In_512);
xnor U1153 (N_1153,In_33,In_857);
nor U1154 (N_1154,In_323,In_698);
nand U1155 (N_1155,In_94,In_335);
and U1156 (N_1156,In_825,In_513);
xnor U1157 (N_1157,In_634,In_30);
or U1158 (N_1158,In_730,In_450);
nor U1159 (N_1159,In_195,In_969);
xnor U1160 (N_1160,In_252,In_556);
and U1161 (N_1161,In_193,In_650);
xor U1162 (N_1162,In_95,In_912);
xnor U1163 (N_1163,In_975,In_805);
nand U1164 (N_1164,In_554,In_395);
nand U1165 (N_1165,In_341,In_410);
nand U1166 (N_1166,In_610,In_852);
or U1167 (N_1167,In_84,In_130);
or U1168 (N_1168,In_113,In_405);
xnor U1169 (N_1169,In_697,In_340);
and U1170 (N_1170,In_73,In_285);
xor U1171 (N_1171,In_254,In_241);
and U1172 (N_1172,In_570,In_724);
nor U1173 (N_1173,In_990,In_20);
or U1174 (N_1174,In_681,In_762);
nand U1175 (N_1175,In_967,In_676);
or U1176 (N_1176,In_682,In_326);
or U1177 (N_1177,In_318,In_235);
nand U1178 (N_1178,In_768,In_309);
or U1179 (N_1179,In_36,In_467);
and U1180 (N_1180,In_832,In_262);
nor U1181 (N_1181,In_181,In_669);
nand U1182 (N_1182,In_398,In_576);
or U1183 (N_1183,In_93,In_648);
nor U1184 (N_1184,In_34,In_862);
nand U1185 (N_1185,In_494,In_771);
and U1186 (N_1186,In_55,In_948);
and U1187 (N_1187,In_363,In_938);
xor U1188 (N_1188,In_300,In_596);
and U1189 (N_1189,In_110,In_647);
nor U1190 (N_1190,In_139,In_547);
nor U1191 (N_1191,In_830,In_469);
or U1192 (N_1192,In_560,In_842);
nand U1193 (N_1193,In_962,In_346);
nor U1194 (N_1194,In_543,In_659);
nand U1195 (N_1195,In_156,In_265);
nand U1196 (N_1196,In_610,In_582);
nor U1197 (N_1197,In_640,In_536);
or U1198 (N_1198,In_343,In_906);
and U1199 (N_1199,In_185,In_883);
and U1200 (N_1200,In_749,In_815);
nor U1201 (N_1201,In_985,In_204);
nand U1202 (N_1202,In_848,In_118);
nor U1203 (N_1203,In_403,In_753);
nand U1204 (N_1204,In_771,In_317);
or U1205 (N_1205,In_789,In_850);
nor U1206 (N_1206,In_435,In_642);
nand U1207 (N_1207,In_115,In_96);
xnor U1208 (N_1208,In_596,In_841);
nor U1209 (N_1209,In_251,In_563);
xor U1210 (N_1210,In_369,In_886);
nor U1211 (N_1211,In_326,In_262);
nor U1212 (N_1212,In_340,In_488);
and U1213 (N_1213,In_415,In_220);
nand U1214 (N_1214,In_483,In_411);
xor U1215 (N_1215,In_798,In_279);
nor U1216 (N_1216,In_210,In_480);
or U1217 (N_1217,In_941,In_236);
or U1218 (N_1218,In_888,In_624);
nor U1219 (N_1219,In_806,In_785);
or U1220 (N_1220,In_930,In_44);
xor U1221 (N_1221,In_639,In_590);
nand U1222 (N_1222,In_769,In_371);
nand U1223 (N_1223,In_231,In_715);
or U1224 (N_1224,In_301,In_714);
or U1225 (N_1225,In_231,In_107);
nand U1226 (N_1226,In_487,In_410);
nand U1227 (N_1227,In_337,In_912);
or U1228 (N_1228,In_46,In_709);
or U1229 (N_1229,In_650,In_903);
nor U1230 (N_1230,In_234,In_656);
xnor U1231 (N_1231,In_638,In_448);
and U1232 (N_1232,In_86,In_263);
or U1233 (N_1233,In_496,In_646);
xor U1234 (N_1234,In_426,In_472);
and U1235 (N_1235,In_261,In_155);
xor U1236 (N_1236,In_158,In_554);
nor U1237 (N_1237,In_17,In_504);
nand U1238 (N_1238,In_252,In_694);
and U1239 (N_1239,In_504,In_612);
nor U1240 (N_1240,In_114,In_403);
xnor U1241 (N_1241,In_300,In_911);
and U1242 (N_1242,In_453,In_354);
or U1243 (N_1243,In_829,In_45);
nand U1244 (N_1244,In_860,In_754);
nor U1245 (N_1245,In_839,In_783);
and U1246 (N_1246,In_22,In_101);
and U1247 (N_1247,In_995,In_914);
or U1248 (N_1248,In_414,In_834);
nand U1249 (N_1249,In_656,In_339);
or U1250 (N_1250,In_430,In_940);
and U1251 (N_1251,In_608,In_145);
nor U1252 (N_1252,In_885,In_663);
and U1253 (N_1253,In_731,In_162);
or U1254 (N_1254,In_303,In_978);
and U1255 (N_1255,In_394,In_788);
or U1256 (N_1256,In_942,In_810);
and U1257 (N_1257,In_82,In_882);
nand U1258 (N_1258,In_455,In_486);
nand U1259 (N_1259,In_482,In_342);
and U1260 (N_1260,In_57,In_194);
nand U1261 (N_1261,In_11,In_515);
xnor U1262 (N_1262,In_242,In_746);
nor U1263 (N_1263,In_83,In_4);
nand U1264 (N_1264,In_691,In_329);
nor U1265 (N_1265,In_667,In_226);
and U1266 (N_1266,In_945,In_949);
or U1267 (N_1267,In_200,In_187);
nand U1268 (N_1268,In_794,In_948);
nor U1269 (N_1269,In_495,In_876);
or U1270 (N_1270,In_89,In_659);
or U1271 (N_1271,In_911,In_684);
nor U1272 (N_1272,In_633,In_414);
nand U1273 (N_1273,In_141,In_152);
or U1274 (N_1274,In_169,In_740);
and U1275 (N_1275,In_152,In_240);
nor U1276 (N_1276,In_22,In_812);
or U1277 (N_1277,In_686,In_164);
nor U1278 (N_1278,In_531,In_825);
and U1279 (N_1279,In_827,In_608);
and U1280 (N_1280,In_697,In_25);
nor U1281 (N_1281,In_512,In_301);
or U1282 (N_1282,In_946,In_722);
nand U1283 (N_1283,In_623,In_11);
nor U1284 (N_1284,In_114,In_517);
nor U1285 (N_1285,In_264,In_632);
and U1286 (N_1286,In_504,In_523);
and U1287 (N_1287,In_693,In_458);
nand U1288 (N_1288,In_96,In_146);
or U1289 (N_1289,In_434,In_704);
or U1290 (N_1290,In_680,In_891);
nor U1291 (N_1291,In_411,In_40);
or U1292 (N_1292,In_557,In_753);
nand U1293 (N_1293,In_411,In_19);
xnor U1294 (N_1294,In_303,In_842);
nor U1295 (N_1295,In_822,In_809);
and U1296 (N_1296,In_933,In_870);
nand U1297 (N_1297,In_414,In_229);
xor U1298 (N_1298,In_119,In_875);
nor U1299 (N_1299,In_321,In_6);
nand U1300 (N_1300,In_397,In_351);
xnor U1301 (N_1301,In_304,In_524);
or U1302 (N_1302,In_86,In_185);
and U1303 (N_1303,In_383,In_706);
and U1304 (N_1304,In_304,In_626);
nand U1305 (N_1305,In_92,In_672);
or U1306 (N_1306,In_852,In_326);
or U1307 (N_1307,In_71,In_728);
or U1308 (N_1308,In_456,In_927);
xor U1309 (N_1309,In_908,In_326);
xnor U1310 (N_1310,In_483,In_871);
nand U1311 (N_1311,In_367,In_109);
and U1312 (N_1312,In_720,In_479);
or U1313 (N_1313,In_36,In_426);
xor U1314 (N_1314,In_153,In_668);
or U1315 (N_1315,In_749,In_427);
nor U1316 (N_1316,In_494,In_410);
and U1317 (N_1317,In_950,In_106);
or U1318 (N_1318,In_604,In_985);
or U1319 (N_1319,In_819,In_329);
nor U1320 (N_1320,In_784,In_577);
xor U1321 (N_1321,In_118,In_93);
nor U1322 (N_1322,In_621,In_631);
or U1323 (N_1323,In_526,In_172);
and U1324 (N_1324,In_143,In_737);
and U1325 (N_1325,In_945,In_992);
and U1326 (N_1326,In_707,In_330);
nor U1327 (N_1327,In_65,In_745);
nand U1328 (N_1328,In_385,In_687);
or U1329 (N_1329,In_112,In_136);
or U1330 (N_1330,In_263,In_171);
nand U1331 (N_1331,In_462,In_212);
and U1332 (N_1332,In_575,In_613);
nand U1333 (N_1333,In_380,In_356);
nor U1334 (N_1334,In_107,In_559);
xnor U1335 (N_1335,In_299,In_104);
or U1336 (N_1336,In_787,In_686);
nand U1337 (N_1337,In_514,In_524);
nand U1338 (N_1338,In_819,In_807);
or U1339 (N_1339,In_80,In_838);
nand U1340 (N_1340,In_870,In_59);
nand U1341 (N_1341,In_710,In_562);
nand U1342 (N_1342,In_651,In_686);
nand U1343 (N_1343,In_708,In_240);
nand U1344 (N_1344,In_999,In_953);
xor U1345 (N_1345,In_841,In_507);
or U1346 (N_1346,In_72,In_425);
nand U1347 (N_1347,In_995,In_152);
and U1348 (N_1348,In_443,In_25);
nand U1349 (N_1349,In_102,In_228);
and U1350 (N_1350,In_724,In_738);
nor U1351 (N_1351,In_107,In_745);
nand U1352 (N_1352,In_33,In_240);
or U1353 (N_1353,In_806,In_119);
or U1354 (N_1354,In_367,In_682);
xnor U1355 (N_1355,In_3,In_935);
nand U1356 (N_1356,In_874,In_53);
and U1357 (N_1357,In_322,In_768);
and U1358 (N_1358,In_680,In_506);
nor U1359 (N_1359,In_929,In_41);
nand U1360 (N_1360,In_101,In_542);
and U1361 (N_1361,In_157,In_77);
nor U1362 (N_1362,In_488,In_267);
nand U1363 (N_1363,In_259,In_67);
and U1364 (N_1364,In_257,In_757);
or U1365 (N_1365,In_273,In_78);
or U1366 (N_1366,In_642,In_218);
nand U1367 (N_1367,In_643,In_814);
or U1368 (N_1368,In_666,In_318);
nor U1369 (N_1369,In_6,In_585);
nor U1370 (N_1370,In_243,In_710);
nor U1371 (N_1371,In_274,In_902);
nand U1372 (N_1372,In_492,In_350);
or U1373 (N_1373,In_779,In_880);
nor U1374 (N_1374,In_661,In_584);
nor U1375 (N_1375,In_867,In_137);
and U1376 (N_1376,In_126,In_391);
or U1377 (N_1377,In_725,In_483);
or U1378 (N_1378,In_788,In_865);
and U1379 (N_1379,In_132,In_99);
and U1380 (N_1380,In_308,In_134);
or U1381 (N_1381,In_837,In_956);
and U1382 (N_1382,In_403,In_678);
or U1383 (N_1383,In_882,In_443);
or U1384 (N_1384,In_195,In_380);
xor U1385 (N_1385,In_115,In_395);
and U1386 (N_1386,In_769,In_612);
xnor U1387 (N_1387,In_770,In_562);
and U1388 (N_1388,In_694,In_354);
xor U1389 (N_1389,In_750,In_178);
nor U1390 (N_1390,In_320,In_551);
nor U1391 (N_1391,In_603,In_348);
or U1392 (N_1392,In_209,In_250);
nand U1393 (N_1393,In_44,In_591);
or U1394 (N_1394,In_104,In_147);
nor U1395 (N_1395,In_182,In_390);
or U1396 (N_1396,In_670,In_856);
xnor U1397 (N_1397,In_207,In_110);
nor U1398 (N_1398,In_524,In_956);
nand U1399 (N_1399,In_365,In_293);
nand U1400 (N_1400,In_454,In_77);
nand U1401 (N_1401,In_206,In_168);
nor U1402 (N_1402,In_409,In_867);
nand U1403 (N_1403,In_865,In_332);
nor U1404 (N_1404,In_872,In_53);
and U1405 (N_1405,In_816,In_205);
or U1406 (N_1406,In_728,In_347);
nand U1407 (N_1407,In_615,In_737);
or U1408 (N_1408,In_823,In_838);
and U1409 (N_1409,In_40,In_941);
or U1410 (N_1410,In_388,In_57);
and U1411 (N_1411,In_304,In_424);
nand U1412 (N_1412,In_277,In_183);
nor U1413 (N_1413,In_910,In_237);
or U1414 (N_1414,In_59,In_300);
or U1415 (N_1415,In_841,In_19);
nor U1416 (N_1416,In_289,In_190);
nor U1417 (N_1417,In_842,In_235);
nand U1418 (N_1418,In_357,In_901);
nor U1419 (N_1419,In_957,In_274);
nand U1420 (N_1420,In_160,In_22);
nor U1421 (N_1421,In_480,In_298);
nand U1422 (N_1422,In_287,In_547);
and U1423 (N_1423,In_923,In_61);
and U1424 (N_1424,In_213,In_407);
or U1425 (N_1425,In_276,In_640);
nand U1426 (N_1426,In_271,In_786);
or U1427 (N_1427,In_641,In_148);
and U1428 (N_1428,In_107,In_928);
nor U1429 (N_1429,In_49,In_519);
nand U1430 (N_1430,In_881,In_480);
nand U1431 (N_1431,In_909,In_851);
xnor U1432 (N_1432,In_779,In_45);
and U1433 (N_1433,In_968,In_562);
nor U1434 (N_1434,In_770,In_231);
nor U1435 (N_1435,In_416,In_999);
or U1436 (N_1436,In_790,In_446);
xnor U1437 (N_1437,In_920,In_25);
or U1438 (N_1438,In_559,In_319);
or U1439 (N_1439,In_489,In_684);
and U1440 (N_1440,In_856,In_287);
and U1441 (N_1441,In_799,In_649);
or U1442 (N_1442,In_495,In_156);
or U1443 (N_1443,In_602,In_25);
xor U1444 (N_1444,In_552,In_13);
xnor U1445 (N_1445,In_341,In_488);
nor U1446 (N_1446,In_220,In_739);
nand U1447 (N_1447,In_836,In_247);
and U1448 (N_1448,In_173,In_667);
nor U1449 (N_1449,In_808,In_714);
xnor U1450 (N_1450,In_498,In_200);
nor U1451 (N_1451,In_421,In_325);
or U1452 (N_1452,In_910,In_269);
nor U1453 (N_1453,In_671,In_447);
or U1454 (N_1454,In_402,In_584);
and U1455 (N_1455,In_328,In_815);
nand U1456 (N_1456,In_404,In_79);
nor U1457 (N_1457,In_63,In_138);
nor U1458 (N_1458,In_383,In_136);
or U1459 (N_1459,In_76,In_256);
nor U1460 (N_1460,In_982,In_699);
or U1461 (N_1461,In_104,In_943);
nand U1462 (N_1462,In_199,In_480);
nor U1463 (N_1463,In_904,In_415);
nand U1464 (N_1464,In_34,In_313);
nor U1465 (N_1465,In_571,In_888);
and U1466 (N_1466,In_31,In_122);
or U1467 (N_1467,In_733,In_885);
nand U1468 (N_1468,In_533,In_420);
and U1469 (N_1469,In_363,In_830);
or U1470 (N_1470,In_102,In_617);
and U1471 (N_1471,In_596,In_448);
and U1472 (N_1472,In_507,In_550);
or U1473 (N_1473,In_478,In_656);
xor U1474 (N_1474,In_525,In_616);
and U1475 (N_1475,In_230,In_792);
and U1476 (N_1476,In_624,In_416);
nor U1477 (N_1477,In_806,In_20);
nor U1478 (N_1478,In_871,In_235);
xor U1479 (N_1479,In_493,In_927);
and U1480 (N_1480,In_750,In_245);
and U1481 (N_1481,In_538,In_216);
and U1482 (N_1482,In_509,In_689);
xnor U1483 (N_1483,In_692,In_258);
xnor U1484 (N_1484,In_763,In_4);
and U1485 (N_1485,In_522,In_189);
or U1486 (N_1486,In_98,In_904);
and U1487 (N_1487,In_389,In_247);
nor U1488 (N_1488,In_952,In_776);
nand U1489 (N_1489,In_866,In_207);
or U1490 (N_1490,In_377,In_456);
and U1491 (N_1491,In_299,In_666);
or U1492 (N_1492,In_915,In_807);
nor U1493 (N_1493,In_993,In_781);
and U1494 (N_1494,In_761,In_912);
xor U1495 (N_1495,In_91,In_231);
and U1496 (N_1496,In_582,In_478);
nor U1497 (N_1497,In_473,In_994);
and U1498 (N_1498,In_360,In_705);
nor U1499 (N_1499,In_14,In_759);
or U1500 (N_1500,In_70,In_419);
and U1501 (N_1501,In_508,In_157);
nand U1502 (N_1502,In_605,In_641);
xnor U1503 (N_1503,In_670,In_475);
xor U1504 (N_1504,In_366,In_392);
nand U1505 (N_1505,In_199,In_264);
nand U1506 (N_1506,In_931,In_483);
nor U1507 (N_1507,In_845,In_428);
and U1508 (N_1508,In_749,In_348);
nand U1509 (N_1509,In_772,In_694);
and U1510 (N_1510,In_575,In_824);
or U1511 (N_1511,In_417,In_263);
or U1512 (N_1512,In_223,In_626);
xnor U1513 (N_1513,In_936,In_738);
nand U1514 (N_1514,In_182,In_737);
or U1515 (N_1515,In_847,In_916);
nor U1516 (N_1516,In_20,In_520);
and U1517 (N_1517,In_224,In_908);
nand U1518 (N_1518,In_307,In_116);
and U1519 (N_1519,In_991,In_503);
or U1520 (N_1520,In_602,In_992);
nor U1521 (N_1521,In_313,In_868);
nand U1522 (N_1522,In_286,In_868);
nand U1523 (N_1523,In_401,In_507);
nand U1524 (N_1524,In_475,In_71);
nor U1525 (N_1525,In_219,In_704);
nor U1526 (N_1526,In_804,In_489);
and U1527 (N_1527,In_889,In_285);
nand U1528 (N_1528,In_284,In_166);
or U1529 (N_1529,In_81,In_44);
and U1530 (N_1530,In_745,In_764);
xnor U1531 (N_1531,In_967,In_389);
or U1532 (N_1532,In_862,In_121);
nor U1533 (N_1533,In_968,In_859);
nor U1534 (N_1534,In_823,In_739);
and U1535 (N_1535,In_177,In_263);
or U1536 (N_1536,In_332,In_920);
nand U1537 (N_1537,In_890,In_184);
nor U1538 (N_1538,In_960,In_835);
or U1539 (N_1539,In_867,In_905);
nand U1540 (N_1540,In_392,In_864);
nand U1541 (N_1541,In_450,In_137);
and U1542 (N_1542,In_275,In_16);
nor U1543 (N_1543,In_947,In_938);
or U1544 (N_1544,In_733,In_770);
nor U1545 (N_1545,In_816,In_242);
xor U1546 (N_1546,In_7,In_143);
nand U1547 (N_1547,In_953,In_30);
and U1548 (N_1548,In_188,In_929);
and U1549 (N_1549,In_620,In_256);
or U1550 (N_1550,In_470,In_346);
xor U1551 (N_1551,In_627,In_912);
nor U1552 (N_1552,In_419,In_424);
nor U1553 (N_1553,In_735,In_472);
or U1554 (N_1554,In_542,In_847);
or U1555 (N_1555,In_644,In_376);
xor U1556 (N_1556,In_605,In_177);
xor U1557 (N_1557,In_837,In_228);
xnor U1558 (N_1558,In_600,In_765);
or U1559 (N_1559,In_821,In_749);
or U1560 (N_1560,In_524,In_824);
nand U1561 (N_1561,In_496,In_456);
and U1562 (N_1562,In_987,In_501);
nand U1563 (N_1563,In_302,In_624);
nand U1564 (N_1564,In_928,In_447);
and U1565 (N_1565,In_731,In_211);
nor U1566 (N_1566,In_985,In_507);
or U1567 (N_1567,In_59,In_966);
nand U1568 (N_1568,In_296,In_805);
and U1569 (N_1569,In_322,In_357);
or U1570 (N_1570,In_712,In_404);
or U1571 (N_1571,In_350,In_205);
and U1572 (N_1572,In_2,In_785);
and U1573 (N_1573,In_660,In_281);
nand U1574 (N_1574,In_702,In_182);
or U1575 (N_1575,In_315,In_32);
xor U1576 (N_1576,In_521,In_855);
nand U1577 (N_1577,In_313,In_751);
xor U1578 (N_1578,In_467,In_587);
and U1579 (N_1579,In_887,In_84);
nor U1580 (N_1580,In_677,In_506);
nand U1581 (N_1581,In_200,In_684);
nor U1582 (N_1582,In_262,In_30);
or U1583 (N_1583,In_123,In_542);
or U1584 (N_1584,In_830,In_987);
or U1585 (N_1585,In_627,In_741);
or U1586 (N_1586,In_557,In_510);
nand U1587 (N_1587,In_246,In_555);
xnor U1588 (N_1588,In_615,In_708);
nand U1589 (N_1589,In_721,In_651);
nor U1590 (N_1590,In_396,In_572);
and U1591 (N_1591,In_0,In_921);
nor U1592 (N_1592,In_993,In_596);
and U1593 (N_1593,In_737,In_636);
nor U1594 (N_1594,In_397,In_969);
nand U1595 (N_1595,In_576,In_910);
xnor U1596 (N_1596,In_364,In_913);
or U1597 (N_1597,In_393,In_516);
or U1598 (N_1598,In_592,In_706);
and U1599 (N_1599,In_90,In_920);
and U1600 (N_1600,In_40,In_248);
and U1601 (N_1601,In_965,In_774);
or U1602 (N_1602,In_386,In_114);
or U1603 (N_1603,In_916,In_380);
nand U1604 (N_1604,In_715,In_501);
and U1605 (N_1605,In_354,In_561);
and U1606 (N_1606,In_191,In_9);
or U1607 (N_1607,In_25,In_67);
nand U1608 (N_1608,In_923,In_697);
nand U1609 (N_1609,In_262,In_860);
nand U1610 (N_1610,In_445,In_342);
nand U1611 (N_1611,In_158,In_3);
and U1612 (N_1612,In_36,In_846);
and U1613 (N_1613,In_553,In_93);
and U1614 (N_1614,In_37,In_540);
nor U1615 (N_1615,In_731,In_351);
nand U1616 (N_1616,In_310,In_888);
nor U1617 (N_1617,In_24,In_111);
or U1618 (N_1618,In_497,In_178);
and U1619 (N_1619,In_260,In_115);
and U1620 (N_1620,In_772,In_833);
and U1621 (N_1621,In_349,In_608);
nor U1622 (N_1622,In_94,In_191);
nand U1623 (N_1623,In_966,In_714);
xnor U1624 (N_1624,In_879,In_943);
nand U1625 (N_1625,In_79,In_118);
nor U1626 (N_1626,In_360,In_312);
nor U1627 (N_1627,In_564,In_847);
xor U1628 (N_1628,In_795,In_13);
xnor U1629 (N_1629,In_224,In_858);
nand U1630 (N_1630,In_626,In_755);
nand U1631 (N_1631,In_356,In_223);
and U1632 (N_1632,In_516,In_90);
or U1633 (N_1633,In_36,In_352);
nand U1634 (N_1634,In_875,In_297);
nand U1635 (N_1635,In_851,In_579);
or U1636 (N_1636,In_747,In_750);
nor U1637 (N_1637,In_735,In_32);
or U1638 (N_1638,In_287,In_266);
nor U1639 (N_1639,In_859,In_269);
or U1640 (N_1640,In_709,In_850);
nand U1641 (N_1641,In_225,In_622);
or U1642 (N_1642,In_781,In_778);
nor U1643 (N_1643,In_232,In_722);
or U1644 (N_1644,In_432,In_342);
nor U1645 (N_1645,In_75,In_823);
nand U1646 (N_1646,In_335,In_707);
nand U1647 (N_1647,In_435,In_151);
and U1648 (N_1648,In_691,In_538);
or U1649 (N_1649,In_956,In_354);
and U1650 (N_1650,In_237,In_31);
or U1651 (N_1651,In_931,In_720);
and U1652 (N_1652,In_947,In_143);
and U1653 (N_1653,In_946,In_226);
nor U1654 (N_1654,In_716,In_740);
xnor U1655 (N_1655,In_893,In_739);
nor U1656 (N_1656,In_0,In_825);
or U1657 (N_1657,In_781,In_594);
and U1658 (N_1658,In_365,In_985);
or U1659 (N_1659,In_52,In_587);
nand U1660 (N_1660,In_63,In_329);
nand U1661 (N_1661,In_555,In_207);
or U1662 (N_1662,In_362,In_304);
xor U1663 (N_1663,In_495,In_466);
xnor U1664 (N_1664,In_726,In_639);
or U1665 (N_1665,In_571,In_820);
and U1666 (N_1666,In_185,In_7);
or U1667 (N_1667,In_289,In_813);
nor U1668 (N_1668,In_931,In_201);
and U1669 (N_1669,In_60,In_532);
nand U1670 (N_1670,In_602,In_935);
nand U1671 (N_1671,In_276,In_678);
or U1672 (N_1672,In_475,In_336);
nand U1673 (N_1673,In_479,In_122);
nor U1674 (N_1674,In_108,In_921);
nand U1675 (N_1675,In_458,In_922);
or U1676 (N_1676,In_611,In_722);
or U1677 (N_1677,In_841,In_962);
nand U1678 (N_1678,In_315,In_60);
or U1679 (N_1679,In_120,In_470);
xor U1680 (N_1680,In_420,In_656);
and U1681 (N_1681,In_697,In_561);
or U1682 (N_1682,In_561,In_99);
and U1683 (N_1683,In_45,In_613);
nor U1684 (N_1684,In_960,In_157);
nand U1685 (N_1685,In_569,In_117);
nor U1686 (N_1686,In_198,In_936);
and U1687 (N_1687,In_52,In_922);
nand U1688 (N_1688,In_671,In_556);
xnor U1689 (N_1689,In_959,In_104);
nand U1690 (N_1690,In_125,In_784);
or U1691 (N_1691,In_359,In_495);
nor U1692 (N_1692,In_887,In_750);
or U1693 (N_1693,In_561,In_823);
nand U1694 (N_1694,In_953,In_704);
nor U1695 (N_1695,In_101,In_433);
or U1696 (N_1696,In_891,In_997);
nand U1697 (N_1697,In_342,In_822);
xnor U1698 (N_1698,In_826,In_670);
or U1699 (N_1699,In_479,In_940);
nand U1700 (N_1700,In_22,In_456);
and U1701 (N_1701,In_458,In_544);
or U1702 (N_1702,In_263,In_924);
nand U1703 (N_1703,In_607,In_84);
or U1704 (N_1704,In_594,In_349);
nand U1705 (N_1705,In_779,In_745);
nor U1706 (N_1706,In_429,In_760);
xnor U1707 (N_1707,In_419,In_198);
nand U1708 (N_1708,In_937,In_767);
or U1709 (N_1709,In_565,In_444);
and U1710 (N_1710,In_14,In_683);
xnor U1711 (N_1711,In_620,In_124);
nor U1712 (N_1712,In_232,In_680);
nand U1713 (N_1713,In_986,In_459);
or U1714 (N_1714,In_25,In_303);
nor U1715 (N_1715,In_361,In_511);
and U1716 (N_1716,In_34,In_2);
nand U1717 (N_1717,In_650,In_349);
xnor U1718 (N_1718,In_188,In_606);
nand U1719 (N_1719,In_345,In_242);
nor U1720 (N_1720,In_652,In_839);
xor U1721 (N_1721,In_729,In_429);
or U1722 (N_1722,In_463,In_562);
and U1723 (N_1723,In_179,In_19);
and U1724 (N_1724,In_598,In_832);
nor U1725 (N_1725,In_3,In_451);
or U1726 (N_1726,In_512,In_146);
nor U1727 (N_1727,In_20,In_540);
nand U1728 (N_1728,In_940,In_560);
or U1729 (N_1729,In_232,In_424);
xor U1730 (N_1730,In_790,In_922);
and U1731 (N_1731,In_559,In_818);
nand U1732 (N_1732,In_999,In_903);
or U1733 (N_1733,In_571,In_487);
nand U1734 (N_1734,In_35,In_860);
or U1735 (N_1735,In_644,In_944);
and U1736 (N_1736,In_450,In_229);
xor U1737 (N_1737,In_779,In_446);
nand U1738 (N_1738,In_918,In_80);
or U1739 (N_1739,In_282,In_242);
or U1740 (N_1740,In_106,In_744);
and U1741 (N_1741,In_750,In_803);
and U1742 (N_1742,In_664,In_647);
xor U1743 (N_1743,In_529,In_115);
or U1744 (N_1744,In_173,In_271);
and U1745 (N_1745,In_956,In_348);
and U1746 (N_1746,In_993,In_994);
nand U1747 (N_1747,In_837,In_935);
nand U1748 (N_1748,In_396,In_426);
or U1749 (N_1749,In_760,In_159);
or U1750 (N_1750,In_164,In_660);
nand U1751 (N_1751,In_184,In_495);
or U1752 (N_1752,In_65,In_247);
nand U1753 (N_1753,In_991,In_990);
nand U1754 (N_1754,In_34,In_535);
nand U1755 (N_1755,In_248,In_645);
nor U1756 (N_1756,In_473,In_52);
and U1757 (N_1757,In_818,In_262);
or U1758 (N_1758,In_247,In_252);
nor U1759 (N_1759,In_152,In_355);
nor U1760 (N_1760,In_563,In_525);
or U1761 (N_1761,In_237,In_435);
or U1762 (N_1762,In_545,In_831);
and U1763 (N_1763,In_658,In_364);
nand U1764 (N_1764,In_829,In_378);
nand U1765 (N_1765,In_909,In_338);
nor U1766 (N_1766,In_301,In_354);
and U1767 (N_1767,In_287,In_917);
nor U1768 (N_1768,In_792,In_387);
nand U1769 (N_1769,In_786,In_201);
or U1770 (N_1770,In_92,In_455);
nand U1771 (N_1771,In_685,In_729);
nor U1772 (N_1772,In_94,In_800);
nor U1773 (N_1773,In_70,In_601);
nand U1774 (N_1774,In_989,In_226);
and U1775 (N_1775,In_27,In_521);
or U1776 (N_1776,In_283,In_280);
or U1777 (N_1777,In_618,In_217);
xor U1778 (N_1778,In_801,In_82);
and U1779 (N_1779,In_859,In_829);
and U1780 (N_1780,In_160,In_717);
and U1781 (N_1781,In_331,In_670);
and U1782 (N_1782,In_333,In_487);
nor U1783 (N_1783,In_387,In_899);
and U1784 (N_1784,In_504,In_901);
nor U1785 (N_1785,In_697,In_688);
nand U1786 (N_1786,In_584,In_840);
or U1787 (N_1787,In_466,In_274);
nor U1788 (N_1788,In_273,In_319);
or U1789 (N_1789,In_85,In_642);
and U1790 (N_1790,In_7,In_932);
or U1791 (N_1791,In_551,In_197);
or U1792 (N_1792,In_739,In_127);
nor U1793 (N_1793,In_461,In_596);
or U1794 (N_1794,In_775,In_521);
nand U1795 (N_1795,In_521,In_654);
or U1796 (N_1796,In_892,In_808);
and U1797 (N_1797,In_814,In_962);
or U1798 (N_1798,In_722,In_529);
and U1799 (N_1799,In_780,In_13);
nand U1800 (N_1800,In_726,In_961);
nand U1801 (N_1801,In_894,In_214);
nand U1802 (N_1802,In_553,In_584);
nor U1803 (N_1803,In_315,In_517);
nand U1804 (N_1804,In_779,In_614);
nand U1805 (N_1805,In_18,In_203);
nor U1806 (N_1806,In_127,In_932);
and U1807 (N_1807,In_322,In_93);
or U1808 (N_1808,In_172,In_21);
or U1809 (N_1809,In_867,In_595);
nand U1810 (N_1810,In_498,In_600);
nor U1811 (N_1811,In_400,In_325);
nor U1812 (N_1812,In_419,In_802);
xor U1813 (N_1813,In_154,In_643);
and U1814 (N_1814,In_200,In_178);
xor U1815 (N_1815,In_109,In_800);
nand U1816 (N_1816,In_387,In_757);
or U1817 (N_1817,In_958,In_22);
or U1818 (N_1818,In_780,In_232);
and U1819 (N_1819,In_765,In_145);
and U1820 (N_1820,In_970,In_471);
and U1821 (N_1821,In_386,In_518);
nand U1822 (N_1822,In_300,In_831);
and U1823 (N_1823,In_739,In_636);
nand U1824 (N_1824,In_551,In_36);
and U1825 (N_1825,In_856,In_0);
nor U1826 (N_1826,In_23,In_355);
xor U1827 (N_1827,In_992,In_728);
and U1828 (N_1828,In_401,In_154);
and U1829 (N_1829,In_267,In_70);
xnor U1830 (N_1830,In_262,In_529);
and U1831 (N_1831,In_80,In_261);
nor U1832 (N_1832,In_127,In_38);
xnor U1833 (N_1833,In_671,In_925);
xnor U1834 (N_1834,In_339,In_462);
or U1835 (N_1835,In_254,In_336);
or U1836 (N_1836,In_207,In_549);
and U1837 (N_1837,In_340,In_437);
nor U1838 (N_1838,In_675,In_911);
xor U1839 (N_1839,In_324,In_902);
nor U1840 (N_1840,In_116,In_29);
or U1841 (N_1841,In_43,In_144);
nand U1842 (N_1842,In_714,In_862);
nand U1843 (N_1843,In_313,In_822);
nor U1844 (N_1844,In_922,In_850);
nand U1845 (N_1845,In_247,In_380);
and U1846 (N_1846,In_285,In_168);
and U1847 (N_1847,In_227,In_903);
nor U1848 (N_1848,In_934,In_388);
nand U1849 (N_1849,In_868,In_812);
nand U1850 (N_1850,In_854,In_622);
nor U1851 (N_1851,In_591,In_17);
nand U1852 (N_1852,In_781,In_219);
nand U1853 (N_1853,In_707,In_492);
and U1854 (N_1854,In_398,In_875);
or U1855 (N_1855,In_906,In_432);
nor U1856 (N_1856,In_105,In_173);
and U1857 (N_1857,In_158,In_71);
and U1858 (N_1858,In_823,In_0);
nand U1859 (N_1859,In_515,In_109);
or U1860 (N_1860,In_844,In_268);
nor U1861 (N_1861,In_969,In_77);
and U1862 (N_1862,In_471,In_595);
and U1863 (N_1863,In_352,In_757);
nor U1864 (N_1864,In_553,In_720);
nor U1865 (N_1865,In_825,In_675);
or U1866 (N_1866,In_585,In_309);
and U1867 (N_1867,In_608,In_716);
and U1868 (N_1868,In_581,In_436);
and U1869 (N_1869,In_858,In_301);
xnor U1870 (N_1870,In_622,In_418);
xor U1871 (N_1871,In_650,In_682);
xnor U1872 (N_1872,In_474,In_795);
and U1873 (N_1873,In_468,In_186);
or U1874 (N_1874,In_934,In_199);
and U1875 (N_1875,In_347,In_345);
or U1876 (N_1876,In_566,In_570);
and U1877 (N_1877,In_484,In_470);
and U1878 (N_1878,In_364,In_547);
and U1879 (N_1879,In_346,In_778);
or U1880 (N_1880,In_754,In_386);
nand U1881 (N_1881,In_55,In_640);
nor U1882 (N_1882,In_123,In_814);
xnor U1883 (N_1883,In_763,In_528);
or U1884 (N_1884,In_705,In_525);
and U1885 (N_1885,In_54,In_170);
nor U1886 (N_1886,In_828,In_811);
xor U1887 (N_1887,In_691,In_684);
nand U1888 (N_1888,In_391,In_646);
and U1889 (N_1889,In_2,In_490);
nor U1890 (N_1890,In_387,In_120);
and U1891 (N_1891,In_413,In_854);
nor U1892 (N_1892,In_331,In_393);
or U1893 (N_1893,In_700,In_154);
xnor U1894 (N_1894,In_229,In_684);
xor U1895 (N_1895,In_181,In_774);
and U1896 (N_1896,In_919,In_483);
nand U1897 (N_1897,In_655,In_736);
xnor U1898 (N_1898,In_685,In_930);
and U1899 (N_1899,In_186,In_976);
or U1900 (N_1900,In_759,In_985);
nand U1901 (N_1901,In_606,In_346);
or U1902 (N_1902,In_750,In_964);
and U1903 (N_1903,In_869,In_732);
and U1904 (N_1904,In_653,In_354);
nor U1905 (N_1905,In_35,In_610);
or U1906 (N_1906,In_935,In_478);
nor U1907 (N_1907,In_555,In_729);
and U1908 (N_1908,In_494,In_346);
nand U1909 (N_1909,In_47,In_601);
or U1910 (N_1910,In_961,In_862);
xnor U1911 (N_1911,In_796,In_514);
and U1912 (N_1912,In_799,In_374);
nor U1913 (N_1913,In_526,In_927);
and U1914 (N_1914,In_543,In_874);
and U1915 (N_1915,In_721,In_748);
and U1916 (N_1916,In_948,In_329);
nand U1917 (N_1917,In_37,In_559);
and U1918 (N_1918,In_821,In_690);
and U1919 (N_1919,In_420,In_503);
nand U1920 (N_1920,In_110,In_176);
and U1921 (N_1921,In_396,In_198);
xor U1922 (N_1922,In_811,In_294);
and U1923 (N_1923,In_279,In_612);
xor U1924 (N_1924,In_434,In_593);
nor U1925 (N_1925,In_120,In_334);
nor U1926 (N_1926,In_314,In_204);
or U1927 (N_1927,In_30,In_927);
or U1928 (N_1928,In_592,In_102);
nand U1929 (N_1929,In_703,In_649);
or U1930 (N_1930,In_949,In_139);
and U1931 (N_1931,In_547,In_447);
or U1932 (N_1932,In_788,In_421);
and U1933 (N_1933,In_440,In_958);
nor U1934 (N_1934,In_898,In_498);
or U1935 (N_1935,In_419,In_962);
nor U1936 (N_1936,In_484,In_161);
nand U1937 (N_1937,In_772,In_485);
nor U1938 (N_1938,In_794,In_206);
and U1939 (N_1939,In_29,In_520);
nor U1940 (N_1940,In_634,In_124);
nand U1941 (N_1941,In_269,In_357);
nor U1942 (N_1942,In_485,In_62);
or U1943 (N_1943,In_328,In_121);
nor U1944 (N_1944,In_85,In_764);
and U1945 (N_1945,In_643,In_472);
or U1946 (N_1946,In_410,In_35);
nor U1947 (N_1947,In_471,In_205);
or U1948 (N_1948,In_579,In_174);
or U1949 (N_1949,In_83,In_634);
xor U1950 (N_1950,In_904,In_251);
or U1951 (N_1951,In_141,In_133);
or U1952 (N_1952,In_647,In_25);
or U1953 (N_1953,In_846,In_646);
and U1954 (N_1954,In_34,In_337);
nor U1955 (N_1955,In_63,In_457);
nor U1956 (N_1956,In_30,In_325);
and U1957 (N_1957,In_574,In_46);
nor U1958 (N_1958,In_9,In_115);
nand U1959 (N_1959,In_939,In_73);
xnor U1960 (N_1960,In_563,In_531);
or U1961 (N_1961,In_586,In_99);
or U1962 (N_1962,In_650,In_7);
nor U1963 (N_1963,In_7,In_189);
nor U1964 (N_1964,In_20,In_328);
nand U1965 (N_1965,In_304,In_749);
or U1966 (N_1966,In_716,In_767);
and U1967 (N_1967,In_269,In_797);
and U1968 (N_1968,In_601,In_722);
and U1969 (N_1969,In_854,In_471);
nand U1970 (N_1970,In_126,In_937);
nor U1971 (N_1971,In_21,In_875);
nand U1972 (N_1972,In_217,In_130);
nand U1973 (N_1973,In_107,In_300);
or U1974 (N_1974,In_253,In_23);
and U1975 (N_1975,In_390,In_865);
nand U1976 (N_1976,In_551,In_171);
or U1977 (N_1977,In_817,In_802);
or U1978 (N_1978,In_806,In_172);
xnor U1979 (N_1979,In_932,In_851);
nor U1980 (N_1980,In_201,In_708);
or U1981 (N_1981,In_306,In_774);
xor U1982 (N_1982,In_993,In_838);
and U1983 (N_1983,In_37,In_476);
or U1984 (N_1984,In_938,In_257);
nand U1985 (N_1985,In_438,In_109);
nand U1986 (N_1986,In_429,In_646);
nor U1987 (N_1987,In_729,In_960);
nand U1988 (N_1988,In_769,In_733);
nand U1989 (N_1989,In_209,In_713);
nand U1990 (N_1990,In_443,In_929);
nand U1991 (N_1991,In_86,In_27);
or U1992 (N_1992,In_848,In_325);
nand U1993 (N_1993,In_527,In_269);
nor U1994 (N_1994,In_840,In_438);
nor U1995 (N_1995,In_87,In_610);
or U1996 (N_1996,In_147,In_944);
and U1997 (N_1997,In_230,In_708);
and U1998 (N_1998,In_706,In_564);
nand U1999 (N_1999,In_270,In_956);
and U2000 (N_2000,In_520,In_140);
nor U2001 (N_2001,In_716,In_589);
and U2002 (N_2002,In_257,In_350);
and U2003 (N_2003,In_305,In_578);
xnor U2004 (N_2004,In_543,In_274);
nor U2005 (N_2005,In_883,In_352);
and U2006 (N_2006,In_545,In_208);
nor U2007 (N_2007,In_221,In_511);
nand U2008 (N_2008,In_20,In_721);
nor U2009 (N_2009,In_618,In_881);
nand U2010 (N_2010,In_748,In_243);
and U2011 (N_2011,In_661,In_117);
or U2012 (N_2012,In_855,In_709);
nor U2013 (N_2013,In_786,In_794);
nor U2014 (N_2014,In_655,In_222);
nor U2015 (N_2015,In_527,In_919);
nor U2016 (N_2016,In_636,In_944);
nor U2017 (N_2017,In_62,In_804);
or U2018 (N_2018,In_203,In_290);
nand U2019 (N_2019,In_23,In_543);
nand U2020 (N_2020,In_240,In_520);
nor U2021 (N_2021,In_743,In_825);
nor U2022 (N_2022,In_774,In_162);
and U2023 (N_2023,In_567,In_76);
nor U2024 (N_2024,In_426,In_47);
and U2025 (N_2025,In_230,In_960);
xnor U2026 (N_2026,In_85,In_731);
and U2027 (N_2027,In_31,In_738);
nand U2028 (N_2028,In_197,In_680);
nand U2029 (N_2029,In_336,In_964);
nand U2030 (N_2030,In_462,In_873);
and U2031 (N_2031,In_360,In_212);
and U2032 (N_2032,In_887,In_752);
and U2033 (N_2033,In_651,In_673);
or U2034 (N_2034,In_196,In_971);
nand U2035 (N_2035,In_566,In_806);
or U2036 (N_2036,In_899,In_4);
nand U2037 (N_2037,In_273,In_364);
xor U2038 (N_2038,In_667,In_660);
or U2039 (N_2039,In_68,In_435);
nand U2040 (N_2040,In_233,In_379);
and U2041 (N_2041,In_962,In_244);
nor U2042 (N_2042,In_90,In_422);
nand U2043 (N_2043,In_80,In_865);
nand U2044 (N_2044,In_949,In_450);
and U2045 (N_2045,In_235,In_203);
or U2046 (N_2046,In_901,In_273);
nand U2047 (N_2047,In_7,In_695);
xor U2048 (N_2048,In_973,In_740);
nand U2049 (N_2049,In_110,In_362);
and U2050 (N_2050,In_183,In_299);
or U2051 (N_2051,In_946,In_482);
xor U2052 (N_2052,In_250,In_71);
and U2053 (N_2053,In_309,In_262);
and U2054 (N_2054,In_240,In_449);
nor U2055 (N_2055,In_211,In_566);
nor U2056 (N_2056,In_97,In_408);
nand U2057 (N_2057,In_264,In_958);
xor U2058 (N_2058,In_475,In_822);
or U2059 (N_2059,In_335,In_825);
and U2060 (N_2060,In_69,In_503);
nor U2061 (N_2061,In_517,In_572);
and U2062 (N_2062,In_347,In_823);
xnor U2063 (N_2063,In_172,In_529);
nand U2064 (N_2064,In_95,In_473);
or U2065 (N_2065,In_394,In_176);
nor U2066 (N_2066,In_994,In_664);
xnor U2067 (N_2067,In_215,In_307);
nor U2068 (N_2068,In_583,In_515);
nor U2069 (N_2069,In_455,In_265);
nor U2070 (N_2070,In_875,In_417);
nor U2071 (N_2071,In_36,In_497);
and U2072 (N_2072,In_667,In_736);
or U2073 (N_2073,In_389,In_609);
or U2074 (N_2074,In_609,In_767);
or U2075 (N_2075,In_187,In_900);
nor U2076 (N_2076,In_451,In_682);
nand U2077 (N_2077,In_35,In_127);
or U2078 (N_2078,In_700,In_612);
and U2079 (N_2079,In_986,In_385);
or U2080 (N_2080,In_181,In_4);
and U2081 (N_2081,In_230,In_335);
nand U2082 (N_2082,In_832,In_243);
and U2083 (N_2083,In_543,In_251);
nand U2084 (N_2084,In_116,In_922);
and U2085 (N_2085,In_944,In_691);
and U2086 (N_2086,In_69,In_136);
nor U2087 (N_2087,In_628,In_362);
and U2088 (N_2088,In_269,In_667);
nor U2089 (N_2089,In_270,In_117);
nor U2090 (N_2090,In_729,In_958);
xnor U2091 (N_2091,In_165,In_95);
or U2092 (N_2092,In_605,In_508);
and U2093 (N_2093,In_160,In_422);
and U2094 (N_2094,In_151,In_748);
nor U2095 (N_2095,In_973,In_125);
or U2096 (N_2096,In_891,In_158);
or U2097 (N_2097,In_416,In_971);
or U2098 (N_2098,In_430,In_979);
nor U2099 (N_2099,In_86,In_531);
or U2100 (N_2100,In_163,In_332);
nand U2101 (N_2101,In_631,In_53);
or U2102 (N_2102,In_106,In_885);
nor U2103 (N_2103,In_628,In_752);
nor U2104 (N_2104,In_127,In_779);
nand U2105 (N_2105,In_957,In_881);
and U2106 (N_2106,In_621,In_346);
xnor U2107 (N_2107,In_871,In_986);
xor U2108 (N_2108,In_6,In_334);
and U2109 (N_2109,In_433,In_895);
or U2110 (N_2110,In_300,In_876);
or U2111 (N_2111,In_242,In_207);
nor U2112 (N_2112,In_698,In_131);
nand U2113 (N_2113,In_975,In_125);
or U2114 (N_2114,In_737,In_321);
nand U2115 (N_2115,In_905,In_642);
and U2116 (N_2116,In_930,In_338);
and U2117 (N_2117,In_902,In_404);
nand U2118 (N_2118,In_290,In_852);
or U2119 (N_2119,In_294,In_773);
or U2120 (N_2120,In_951,In_601);
xnor U2121 (N_2121,In_155,In_539);
nand U2122 (N_2122,In_104,In_99);
and U2123 (N_2123,In_147,In_404);
nand U2124 (N_2124,In_550,In_440);
or U2125 (N_2125,In_798,In_49);
nand U2126 (N_2126,In_618,In_297);
nand U2127 (N_2127,In_935,In_313);
and U2128 (N_2128,In_276,In_475);
xnor U2129 (N_2129,In_554,In_629);
or U2130 (N_2130,In_827,In_851);
nor U2131 (N_2131,In_402,In_807);
nor U2132 (N_2132,In_379,In_568);
nor U2133 (N_2133,In_318,In_918);
nand U2134 (N_2134,In_825,In_648);
and U2135 (N_2135,In_99,In_293);
or U2136 (N_2136,In_451,In_585);
or U2137 (N_2137,In_441,In_975);
nand U2138 (N_2138,In_188,In_832);
and U2139 (N_2139,In_764,In_238);
or U2140 (N_2140,In_367,In_614);
and U2141 (N_2141,In_274,In_231);
or U2142 (N_2142,In_476,In_281);
or U2143 (N_2143,In_386,In_515);
or U2144 (N_2144,In_151,In_892);
and U2145 (N_2145,In_699,In_870);
nor U2146 (N_2146,In_399,In_402);
and U2147 (N_2147,In_659,In_828);
nor U2148 (N_2148,In_925,In_553);
and U2149 (N_2149,In_58,In_852);
xnor U2150 (N_2150,In_596,In_439);
and U2151 (N_2151,In_982,In_255);
or U2152 (N_2152,In_14,In_617);
and U2153 (N_2153,In_349,In_514);
and U2154 (N_2154,In_958,In_372);
nand U2155 (N_2155,In_861,In_121);
or U2156 (N_2156,In_740,In_346);
nand U2157 (N_2157,In_820,In_95);
or U2158 (N_2158,In_963,In_742);
or U2159 (N_2159,In_882,In_670);
nand U2160 (N_2160,In_644,In_896);
and U2161 (N_2161,In_741,In_820);
and U2162 (N_2162,In_199,In_455);
and U2163 (N_2163,In_117,In_689);
and U2164 (N_2164,In_272,In_319);
nor U2165 (N_2165,In_735,In_427);
nor U2166 (N_2166,In_419,In_649);
and U2167 (N_2167,In_337,In_153);
or U2168 (N_2168,In_133,In_763);
nand U2169 (N_2169,In_457,In_778);
nor U2170 (N_2170,In_781,In_309);
nand U2171 (N_2171,In_450,In_373);
nand U2172 (N_2172,In_610,In_737);
nor U2173 (N_2173,In_213,In_488);
nand U2174 (N_2174,In_621,In_483);
and U2175 (N_2175,In_545,In_565);
nand U2176 (N_2176,In_164,In_222);
nand U2177 (N_2177,In_60,In_106);
nand U2178 (N_2178,In_303,In_820);
nand U2179 (N_2179,In_244,In_272);
nand U2180 (N_2180,In_784,In_520);
nor U2181 (N_2181,In_658,In_121);
nor U2182 (N_2182,In_505,In_799);
nand U2183 (N_2183,In_945,In_549);
and U2184 (N_2184,In_563,In_739);
or U2185 (N_2185,In_533,In_45);
nor U2186 (N_2186,In_194,In_648);
and U2187 (N_2187,In_749,In_742);
or U2188 (N_2188,In_232,In_99);
nand U2189 (N_2189,In_151,In_978);
xor U2190 (N_2190,In_593,In_777);
nor U2191 (N_2191,In_348,In_437);
nor U2192 (N_2192,In_633,In_463);
or U2193 (N_2193,In_628,In_0);
or U2194 (N_2194,In_383,In_926);
nor U2195 (N_2195,In_320,In_569);
nor U2196 (N_2196,In_173,In_825);
or U2197 (N_2197,In_511,In_672);
and U2198 (N_2198,In_755,In_784);
nand U2199 (N_2199,In_549,In_912);
nand U2200 (N_2200,In_635,In_282);
or U2201 (N_2201,In_735,In_832);
nor U2202 (N_2202,In_318,In_228);
and U2203 (N_2203,In_414,In_74);
xnor U2204 (N_2204,In_123,In_880);
and U2205 (N_2205,In_991,In_143);
or U2206 (N_2206,In_514,In_890);
nor U2207 (N_2207,In_94,In_240);
nand U2208 (N_2208,In_795,In_162);
or U2209 (N_2209,In_612,In_667);
or U2210 (N_2210,In_780,In_389);
or U2211 (N_2211,In_467,In_300);
nor U2212 (N_2212,In_217,In_577);
and U2213 (N_2213,In_884,In_412);
nor U2214 (N_2214,In_394,In_236);
or U2215 (N_2215,In_816,In_411);
nand U2216 (N_2216,In_534,In_200);
or U2217 (N_2217,In_258,In_676);
and U2218 (N_2218,In_285,In_997);
nor U2219 (N_2219,In_387,In_772);
and U2220 (N_2220,In_900,In_733);
nor U2221 (N_2221,In_607,In_166);
nor U2222 (N_2222,In_747,In_682);
nand U2223 (N_2223,In_824,In_728);
or U2224 (N_2224,In_744,In_178);
nor U2225 (N_2225,In_138,In_733);
and U2226 (N_2226,In_139,In_97);
and U2227 (N_2227,In_18,In_221);
or U2228 (N_2228,In_233,In_699);
nand U2229 (N_2229,In_308,In_987);
and U2230 (N_2230,In_622,In_635);
nor U2231 (N_2231,In_33,In_482);
and U2232 (N_2232,In_263,In_227);
or U2233 (N_2233,In_775,In_649);
xor U2234 (N_2234,In_354,In_24);
nor U2235 (N_2235,In_331,In_771);
and U2236 (N_2236,In_285,In_855);
or U2237 (N_2237,In_786,In_355);
nand U2238 (N_2238,In_528,In_0);
nand U2239 (N_2239,In_621,In_157);
or U2240 (N_2240,In_74,In_516);
nand U2241 (N_2241,In_938,In_879);
nor U2242 (N_2242,In_698,In_388);
or U2243 (N_2243,In_322,In_522);
nor U2244 (N_2244,In_907,In_349);
nand U2245 (N_2245,In_378,In_618);
or U2246 (N_2246,In_877,In_42);
and U2247 (N_2247,In_767,In_27);
or U2248 (N_2248,In_473,In_5);
or U2249 (N_2249,In_227,In_244);
nand U2250 (N_2250,In_276,In_13);
or U2251 (N_2251,In_900,In_607);
nor U2252 (N_2252,In_242,In_260);
and U2253 (N_2253,In_105,In_745);
or U2254 (N_2254,In_583,In_83);
xor U2255 (N_2255,In_957,In_414);
nor U2256 (N_2256,In_264,In_535);
nor U2257 (N_2257,In_79,In_439);
or U2258 (N_2258,In_548,In_385);
nand U2259 (N_2259,In_237,In_152);
or U2260 (N_2260,In_65,In_414);
nor U2261 (N_2261,In_320,In_361);
or U2262 (N_2262,In_418,In_899);
and U2263 (N_2263,In_813,In_22);
nand U2264 (N_2264,In_722,In_914);
nand U2265 (N_2265,In_477,In_690);
and U2266 (N_2266,In_283,In_823);
or U2267 (N_2267,In_613,In_25);
and U2268 (N_2268,In_959,In_584);
or U2269 (N_2269,In_984,In_812);
nor U2270 (N_2270,In_581,In_567);
or U2271 (N_2271,In_541,In_31);
nand U2272 (N_2272,In_16,In_299);
or U2273 (N_2273,In_256,In_35);
nand U2274 (N_2274,In_754,In_648);
and U2275 (N_2275,In_431,In_268);
nor U2276 (N_2276,In_657,In_935);
or U2277 (N_2277,In_954,In_423);
and U2278 (N_2278,In_136,In_605);
and U2279 (N_2279,In_198,In_209);
and U2280 (N_2280,In_262,In_84);
nor U2281 (N_2281,In_164,In_439);
nand U2282 (N_2282,In_139,In_72);
nand U2283 (N_2283,In_206,In_687);
nand U2284 (N_2284,In_210,In_361);
and U2285 (N_2285,In_628,In_240);
nand U2286 (N_2286,In_738,In_208);
xor U2287 (N_2287,In_753,In_543);
or U2288 (N_2288,In_703,In_307);
nand U2289 (N_2289,In_211,In_835);
nand U2290 (N_2290,In_913,In_866);
or U2291 (N_2291,In_124,In_846);
or U2292 (N_2292,In_897,In_886);
and U2293 (N_2293,In_407,In_177);
xor U2294 (N_2294,In_933,In_809);
xnor U2295 (N_2295,In_598,In_738);
nor U2296 (N_2296,In_368,In_832);
and U2297 (N_2297,In_519,In_212);
nand U2298 (N_2298,In_382,In_403);
or U2299 (N_2299,In_260,In_343);
nand U2300 (N_2300,In_652,In_283);
nand U2301 (N_2301,In_613,In_460);
nand U2302 (N_2302,In_852,In_679);
and U2303 (N_2303,In_168,In_623);
nand U2304 (N_2304,In_393,In_170);
nand U2305 (N_2305,In_363,In_980);
nor U2306 (N_2306,In_737,In_27);
or U2307 (N_2307,In_786,In_350);
nor U2308 (N_2308,In_17,In_662);
and U2309 (N_2309,In_744,In_247);
nor U2310 (N_2310,In_968,In_254);
xnor U2311 (N_2311,In_999,In_325);
nand U2312 (N_2312,In_870,In_109);
nand U2313 (N_2313,In_848,In_929);
xnor U2314 (N_2314,In_714,In_602);
xor U2315 (N_2315,In_649,In_599);
nor U2316 (N_2316,In_104,In_968);
nor U2317 (N_2317,In_506,In_926);
or U2318 (N_2318,In_451,In_732);
xnor U2319 (N_2319,In_847,In_156);
and U2320 (N_2320,In_80,In_970);
or U2321 (N_2321,In_462,In_8);
or U2322 (N_2322,In_929,In_793);
nand U2323 (N_2323,In_695,In_728);
and U2324 (N_2324,In_856,In_10);
nand U2325 (N_2325,In_456,In_916);
and U2326 (N_2326,In_739,In_47);
and U2327 (N_2327,In_582,In_177);
or U2328 (N_2328,In_380,In_423);
nand U2329 (N_2329,In_386,In_364);
xor U2330 (N_2330,In_97,In_949);
or U2331 (N_2331,In_97,In_291);
and U2332 (N_2332,In_727,In_903);
nor U2333 (N_2333,In_837,In_989);
and U2334 (N_2334,In_187,In_168);
nand U2335 (N_2335,In_328,In_941);
nand U2336 (N_2336,In_754,In_563);
xnor U2337 (N_2337,In_639,In_70);
or U2338 (N_2338,In_24,In_841);
nand U2339 (N_2339,In_969,In_873);
or U2340 (N_2340,In_305,In_827);
nand U2341 (N_2341,In_894,In_212);
and U2342 (N_2342,In_144,In_23);
nand U2343 (N_2343,In_862,In_363);
nor U2344 (N_2344,In_14,In_153);
and U2345 (N_2345,In_528,In_625);
nor U2346 (N_2346,In_0,In_277);
or U2347 (N_2347,In_325,In_953);
nor U2348 (N_2348,In_33,In_326);
or U2349 (N_2349,In_632,In_75);
and U2350 (N_2350,In_607,In_799);
or U2351 (N_2351,In_540,In_904);
or U2352 (N_2352,In_363,In_668);
nor U2353 (N_2353,In_406,In_782);
nand U2354 (N_2354,In_93,In_57);
or U2355 (N_2355,In_372,In_432);
and U2356 (N_2356,In_972,In_127);
nand U2357 (N_2357,In_29,In_297);
or U2358 (N_2358,In_521,In_571);
or U2359 (N_2359,In_201,In_401);
nor U2360 (N_2360,In_633,In_491);
nand U2361 (N_2361,In_720,In_761);
or U2362 (N_2362,In_737,In_187);
or U2363 (N_2363,In_620,In_26);
and U2364 (N_2364,In_24,In_367);
nand U2365 (N_2365,In_408,In_854);
nor U2366 (N_2366,In_402,In_966);
and U2367 (N_2367,In_327,In_569);
or U2368 (N_2368,In_485,In_550);
xor U2369 (N_2369,In_185,In_511);
nand U2370 (N_2370,In_959,In_164);
nor U2371 (N_2371,In_770,In_534);
and U2372 (N_2372,In_710,In_806);
or U2373 (N_2373,In_588,In_598);
and U2374 (N_2374,In_854,In_844);
nand U2375 (N_2375,In_991,In_668);
or U2376 (N_2376,In_407,In_28);
and U2377 (N_2377,In_51,In_298);
nor U2378 (N_2378,In_282,In_875);
nor U2379 (N_2379,In_723,In_335);
xor U2380 (N_2380,In_740,In_758);
nand U2381 (N_2381,In_118,In_688);
or U2382 (N_2382,In_348,In_215);
and U2383 (N_2383,In_694,In_29);
nor U2384 (N_2384,In_75,In_148);
nand U2385 (N_2385,In_958,In_818);
nor U2386 (N_2386,In_407,In_424);
and U2387 (N_2387,In_999,In_438);
and U2388 (N_2388,In_913,In_249);
nand U2389 (N_2389,In_481,In_550);
nand U2390 (N_2390,In_657,In_972);
nor U2391 (N_2391,In_256,In_438);
and U2392 (N_2392,In_127,In_159);
and U2393 (N_2393,In_41,In_278);
nor U2394 (N_2394,In_203,In_721);
or U2395 (N_2395,In_911,In_25);
nor U2396 (N_2396,In_452,In_430);
or U2397 (N_2397,In_900,In_884);
or U2398 (N_2398,In_78,In_574);
or U2399 (N_2399,In_688,In_348);
nor U2400 (N_2400,In_925,In_979);
or U2401 (N_2401,In_584,In_104);
nand U2402 (N_2402,In_706,In_624);
nand U2403 (N_2403,In_997,In_244);
nor U2404 (N_2404,In_81,In_976);
nor U2405 (N_2405,In_798,In_302);
xnor U2406 (N_2406,In_624,In_778);
xnor U2407 (N_2407,In_462,In_988);
nor U2408 (N_2408,In_233,In_352);
nand U2409 (N_2409,In_521,In_231);
nor U2410 (N_2410,In_668,In_867);
nand U2411 (N_2411,In_317,In_338);
and U2412 (N_2412,In_970,In_224);
or U2413 (N_2413,In_730,In_281);
and U2414 (N_2414,In_619,In_504);
xor U2415 (N_2415,In_919,In_297);
nor U2416 (N_2416,In_610,In_990);
and U2417 (N_2417,In_410,In_417);
or U2418 (N_2418,In_167,In_236);
and U2419 (N_2419,In_254,In_969);
nand U2420 (N_2420,In_908,In_946);
or U2421 (N_2421,In_789,In_547);
nand U2422 (N_2422,In_482,In_258);
xnor U2423 (N_2423,In_301,In_292);
or U2424 (N_2424,In_268,In_995);
nand U2425 (N_2425,In_457,In_66);
and U2426 (N_2426,In_365,In_562);
or U2427 (N_2427,In_238,In_647);
nor U2428 (N_2428,In_235,In_564);
nor U2429 (N_2429,In_534,In_504);
nand U2430 (N_2430,In_479,In_455);
nor U2431 (N_2431,In_991,In_485);
or U2432 (N_2432,In_641,In_457);
and U2433 (N_2433,In_440,In_419);
nand U2434 (N_2434,In_199,In_669);
or U2435 (N_2435,In_245,In_844);
nand U2436 (N_2436,In_215,In_613);
and U2437 (N_2437,In_839,In_471);
nand U2438 (N_2438,In_36,In_303);
or U2439 (N_2439,In_535,In_305);
or U2440 (N_2440,In_256,In_340);
or U2441 (N_2441,In_595,In_53);
or U2442 (N_2442,In_693,In_193);
and U2443 (N_2443,In_308,In_294);
and U2444 (N_2444,In_153,In_662);
or U2445 (N_2445,In_860,In_777);
and U2446 (N_2446,In_543,In_738);
nand U2447 (N_2447,In_871,In_55);
or U2448 (N_2448,In_244,In_248);
and U2449 (N_2449,In_387,In_381);
nand U2450 (N_2450,In_945,In_931);
or U2451 (N_2451,In_935,In_354);
or U2452 (N_2452,In_225,In_459);
and U2453 (N_2453,In_362,In_440);
or U2454 (N_2454,In_522,In_819);
and U2455 (N_2455,In_557,In_263);
nor U2456 (N_2456,In_833,In_816);
nor U2457 (N_2457,In_255,In_851);
nor U2458 (N_2458,In_594,In_289);
xor U2459 (N_2459,In_914,In_804);
nand U2460 (N_2460,In_560,In_105);
and U2461 (N_2461,In_973,In_769);
and U2462 (N_2462,In_392,In_772);
or U2463 (N_2463,In_749,In_715);
nand U2464 (N_2464,In_971,In_249);
nor U2465 (N_2465,In_162,In_424);
xor U2466 (N_2466,In_645,In_485);
or U2467 (N_2467,In_158,In_611);
or U2468 (N_2468,In_554,In_653);
nor U2469 (N_2469,In_751,In_258);
and U2470 (N_2470,In_753,In_613);
and U2471 (N_2471,In_202,In_472);
nor U2472 (N_2472,In_387,In_988);
nand U2473 (N_2473,In_308,In_408);
or U2474 (N_2474,In_866,In_710);
nand U2475 (N_2475,In_265,In_967);
nand U2476 (N_2476,In_39,In_437);
xor U2477 (N_2477,In_629,In_478);
nand U2478 (N_2478,In_710,In_570);
nor U2479 (N_2479,In_276,In_788);
or U2480 (N_2480,In_343,In_361);
or U2481 (N_2481,In_490,In_760);
or U2482 (N_2482,In_22,In_515);
and U2483 (N_2483,In_1,In_231);
or U2484 (N_2484,In_942,In_532);
and U2485 (N_2485,In_876,In_345);
nand U2486 (N_2486,In_581,In_633);
nand U2487 (N_2487,In_300,In_874);
and U2488 (N_2488,In_242,In_867);
or U2489 (N_2489,In_935,In_979);
nand U2490 (N_2490,In_199,In_907);
and U2491 (N_2491,In_32,In_63);
or U2492 (N_2492,In_66,In_39);
nor U2493 (N_2493,In_784,In_394);
nor U2494 (N_2494,In_777,In_47);
and U2495 (N_2495,In_41,In_311);
or U2496 (N_2496,In_258,In_440);
and U2497 (N_2497,In_279,In_57);
nand U2498 (N_2498,In_439,In_494);
or U2499 (N_2499,In_263,In_603);
and U2500 (N_2500,In_803,In_335);
or U2501 (N_2501,In_937,In_327);
and U2502 (N_2502,In_457,In_64);
or U2503 (N_2503,In_570,In_777);
or U2504 (N_2504,In_463,In_204);
nand U2505 (N_2505,In_148,In_509);
xnor U2506 (N_2506,In_482,In_931);
nor U2507 (N_2507,In_629,In_727);
xor U2508 (N_2508,In_222,In_555);
and U2509 (N_2509,In_313,In_214);
or U2510 (N_2510,In_815,In_161);
and U2511 (N_2511,In_430,In_988);
nand U2512 (N_2512,In_314,In_922);
and U2513 (N_2513,In_148,In_816);
nor U2514 (N_2514,In_695,In_932);
nand U2515 (N_2515,In_998,In_734);
or U2516 (N_2516,In_628,In_490);
nand U2517 (N_2517,In_640,In_503);
xnor U2518 (N_2518,In_532,In_543);
xnor U2519 (N_2519,In_295,In_126);
nand U2520 (N_2520,In_568,In_292);
nor U2521 (N_2521,In_158,In_576);
nand U2522 (N_2522,In_484,In_115);
and U2523 (N_2523,In_292,In_832);
nor U2524 (N_2524,In_282,In_225);
and U2525 (N_2525,In_410,In_366);
nor U2526 (N_2526,In_171,In_478);
xnor U2527 (N_2527,In_693,In_780);
or U2528 (N_2528,In_473,In_435);
and U2529 (N_2529,In_436,In_924);
or U2530 (N_2530,In_581,In_382);
nand U2531 (N_2531,In_170,In_292);
and U2532 (N_2532,In_44,In_497);
and U2533 (N_2533,In_966,In_848);
or U2534 (N_2534,In_243,In_388);
nand U2535 (N_2535,In_318,In_887);
xor U2536 (N_2536,In_558,In_425);
nand U2537 (N_2537,In_707,In_10);
nand U2538 (N_2538,In_812,In_790);
nor U2539 (N_2539,In_873,In_311);
xor U2540 (N_2540,In_226,In_406);
and U2541 (N_2541,In_759,In_919);
nor U2542 (N_2542,In_480,In_862);
nand U2543 (N_2543,In_454,In_579);
nor U2544 (N_2544,In_275,In_611);
and U2545 (N_2545,In_826,In_178);
nor U2546 (N_2546,In_424,In_770);
nor U2547 (N_2547,In_757,In_101);
nand U2548 (N_2548,In_173,In_542);
or U2549 (N_2549,In_812,In_432);
nor U2550 (N_2550,In_608,In_191);
nor U2551 (N_2551,In_212,In_367);
nand U2552 (N_2552,In_842,In_934);
or U2553 (N_2553,In_174,In_312);
and U2554 (N_2554,In_694,In_955);
or U2555 (N_2555,In_768,In_299);
or U2556 (N_2556,In_460,In_866);
nand U2557 (N_2557,In_355,In_272);
nor U2558 (N_2558,In_101,In_87);
or U2559 (N_2559,In_776,In_378);
xnor U2560 (N_2560,In_149,In_952);
nand U2561 (N_2561,In_168,In_420);
and U2562 (N_2562,In_344,In_760);
nor U2563 (N_2563,In_169,In_372);
and U2564 (N_2564,In_643,In_789);
or U2565 (N_2565,In_715,In_393);
nor U2566 (N_2566,In_477,In_230);
nand U2567 (N_2567,In_48,In_890);
or U2568 (N_2568,In_759,In_468);
nand U2569 (N_2569,In_93,In_552);
or U2570 (N_2570,In_931,In_135);
nor U2571 (N_2571,In_774,In_485);
and U2572 (N_2572,In_412,In_457);
and U2573 (N_2573,In_674,In_985);
and U2574 (N_2574,In_819,In_423);
xor U2575 (N_2575,In_69,In_158);
nor U2576 (N_2576,In_128,In_825);
nor U2577 (N_2577,In_858,In_121);
and U2578 (N_2578,In_527,In_20);
and U2579 (N_2579,In_226,In_761);
or U2580 (N_2580,In_136,In_494);
xnor U2581 (N_2581,In_186,In_371);
or U2582 (N_2582,In_777,In_984);
nand U2583 (N_2583,In_749,In_853);
nand U2584 (N_2584,In_2,In_724);
and U2585 (N_2585,In_666,In_759);
nor U2586 (N_2586,In_175,In_705);
or U2587 (N_2587,In_524,In_199);
and U2588 (N_2588,In_673,In_740);
nor U2589 (N_2589,In_24,In_660);
nand U2590 (N_2590,In_699,In_842);
xor U2591 (N_2591,In_132,In_179);
nand U2592 (N_2592,In_401,In_237);
nand U2593 (N_2593,In_156,In_984);
or U2594 (N_2594,In_677,In_788);
nand U2595 (N_2595,In_387,In_29);
nor U2596 (N_2596,In_739,In_361);
xor U2597 (N_2597,In_882,In_913);
or U2598 (N_2598,In_51,In_464);
or U2599 (N_2599,In_610,In_518);
or U2600 (N_2600,In_621,In_563);
or U2601 (N_2601,In_535,In_115);
or U2602 (N_2602,In_416,In_589);
and U2603 (N_2603,In_551,In_377);
or U2604 (N_2604,In_453,In_355);
nand U2605 (N_2605,In_807,In_40);
nor U2606 (N_2606,In_965,In_564);
nor U2607 (N_2607,In_930,In_462);
and U2608 (N_2608,In_6,In_902);
nor U2609 (N_2609,In_731,In_433);
xnor U2610 (N_2610,In_522,In_118);
or U2611 (N_2611,In_371,In_408);
nand U2612 (N_2612,In_695,In_463);
and U2613 (N_2613,In_777,In_9);
nor U2614 (N_2614,In_875,In_477);
or U2615 (N_2615,In_455,In_861);
nor U2616 (N_2616,In_96,In_330);
nor U2617 (N_2617,In_945,In_647);
xor U2618 (N_2618,In_172,In_737);
nand U2619 (N_2619,In_348,In_717);
and U2620 (N_2620,In_581,In_985);
nand U2621 (N_2621,In_809,In_280);
nand U2622 (N_2622,In_833,In_614);
or U2623 (N_2623,In_640,In_616);
or U2624 (N_2624,In_181,In_483);
or U2625 (N_2625,In_584,In_710);
or U2626 (N_2626,In_92,In_554);
nand U2627 (N_2627,In_259,In_253);
or U2628 (N_2628,In_562,In_966);
nor U2629 (N_2629,In_636,In_893);
and U2630 (N_2630,In_882,In_604);
and U2631 (N_2631,In_321,In_658);
xnor U2632 (N_2632,In_370,In_761);
xor U2633 (N_2633,In_191,In_332);
xnor U2634 (N_2634,In_173,In_270);
xnor U2635 (N_2635,In_510,In_770);
or U2636 (N_2636,In_197,In_467);
and U2637 (N_2637,In_192,In_863);
and U2638 (N_2638,In_331,In_203);
or U2639 (N_2639,In_212,In_517);
nand U2640 (N_2640,In_774,In_19);
nand U2641 (N_2641,In_709,In_54);
or U2642 (N_2642,In_541,In_268);
xnor U2643 (N_2643,In_981,In_439);
xor U2644 (N_2644,In_723,In_495);
and U2645 (N_2645,In_336,In_658);
xor U2646 (N_2646,In_856,In_152);
and U2647 (N_2647,In_316,In_82);
and U2648 (N_2648,In_676,In_45);
nor U2649 (N_2649,In_197,In_150);
and U2650 (N_2650,In_561,In_549);
or U2651 (N_2651,In_665,In_62);
and U2652 (N_2652,In_579,In_272);
xor U2653 (N_2653,In_479,In_747);
nor U2654 (N_2654,In_21,In_88);
nand U2655 (N_2655,In_622,In_300);
or U2656 (N_2656,In_696,In_261);
nand U2657 (N_2657,In_82,In_928);
xnor U2658 (N_2658,In_806,In_549);
or U2659 (N_2659,In_534,In_380);
nor U2660 (N_2660,In_275,In_601);
xor U2661 (N_2661,In_169,In_856);
nor U2662 (N_2662,In_601,In_428);
or U2663 (N_2663,In_999,In_197);
and U2664 (N_2664,In_333,In_425);
or U2665 (N_2665,In_646,In_399);
and U2666 (N_2666,In_248,In_613);
xnor U2667 (N_2667,In_166,In_498);
or U2668 (N_2668,In_570,In_804);
nor U2669 (N_2669,In_807,In_194);
and U2670 (N_2670,In_392,In_239);
or U2671 (N_2671,In_246,In_852);
or U2672 (N_2672,In_350,In_33);
and U2673 (N_2673,In_836,In_236);
nand U2674 (N_2674,In_911,In_589);
nor U2675 (N_2675,In_378,In_549);
or U2676 (N_2676,In_175,In_440);
xor U2677 (N_2677,In_989,In_434);
and U2678 (N_2678,In_649,In_406);
nor U2679 (N_2679,In_988,In_278);
nand U2680 (N_2680,In_452,In_487);
and U2681 (N_2681,In_984,In_429);
nand U2682 (N_2682,In_285,In_72);
or U2683 (N_2683,In_225,In_415);
and U2684 (N_2684,In_894,In_119);
or U2685 (N_2685,In_348,In_685);
nor U2686 (N_2686,In_969,In_184);
nand U2687 (N_2687,In_455,In_380);
nand U2688 (N_2688,In_584,In_168);
or U2689 (N_2689,In_959,In_685);
or U2690 (N_2690,In_357,In_840);
nor U2691 (N_2691,In_71,In_148);
nor U2692 (N_2692,In_271,In_281);
or U2693 (N_2693,In_388,In_418);
nor U2694 (N_2694,In_212,In_285);
xnor U2695 (N_2695,In_582,In_137);
nand U2696 (N_2696,In_687,In_173);
nand U2697 (N_2697,In_180,In_463);
and U2698 (N_2698,In_270,In_848);
or U2699 (N_2699,In_457,In_363);
xor U2700 (N_2700,In_354,In_381);
xnor U2701 (N_2701,In_7,In_716);
or U2702 (N_2702,In_319,In_194);
and U2703 (N_2703,In_304,In_650);
nand U2704 (N_2704,In_74,In_333);
or U2705 (N_2705,In_579,In_255);
nand U2706 (N_2706,In_729,In_716);
nor U2707 (N_2707,In_384,In_502);
and U2708 (N_2708,In_410,In_731);
xor U2709 (N_2709,In_63,In_464);
or U2710 (N_2710,In_514,In_206);
nor U2711 (N_2711,In_63,In_260);
nand U2712 (N_2712,In_387,In_759);
or U2713 (N_2713,In_431,In_535);
nand U2714 (N_2714,In_751,In_834);
nor U2715 (N_2715,In_862,In_302);
or U2716 (N_2716,In_441,In_56);
and U2717 (N_2717,In_102,In_196);
nor U2718 (N_2718,In_335,In_95);
nor U2719 (N_2719,In_427,In_859);
nand U2720 (N_2720,In_3,In_534);
or U2721 (N_2721,In_743,In_712);
and U2722 (N_2722,In_328,In_827);
nor U2723 (N_2723,In_820,In_335);
nor U2724 (N_2724,In_601,In_205);
nor U2725 (N_2725,In_268,In_449);
nand U2726 (N_2726,In_77,In_752);
xnor U2727 (N_2727,In_513,In_803);
xor U2728 (N_2728,In_892,In_191);
xnor U2729 (N_2729,In_729,In_785);
xnor U2730 (N_2730,In_700,In_742);
xnor U2731 (N_2731,In_609,In_333);
and U2732 (N_2732,In_469,In_353);
or U2733 (N_2733,In_746,In_723);
and U2734 (N_2734,In_223,In_440);
nand U2735 (N_2735,In_33,In_589);
xnor U2736 (N_2736,In_151,In_903);
nand U2737 (N_2737,In_622,In_176);
nand U2738 (N_2738,In_201,In_220);
and U2739 (N_2739,In_678,In_551);
or U2740 (N_2740,In_147,In_103);
xor U2741 (N_2741,In_730,In_855);
xor U2742 (N_2742,In_141,In_432);
xor U2743 (N_2743,In_611,In_455);
and U2744 (N_2744,In_993,In_140);
nand U2745 (N_2745,In_52,In_787);
and U2746 (N_2746,In_79,In_785);
nor U2747 (N_2747,In_859,In_879);
nor U2748 (N_2748,In_864,In_777);
nand U2749 (N_2749,In_862,In_828);
or U2750 (N_2750,In_797,In_624);
and U2751 (N_2751,In_832,In_791);
nand U2752 (N_2752,In_832,In_568);
nor U2753 (N_2753,In_8,In_829);
nor U2754 (N_2754,In_497,In_873);
and U2755 (N_2755,In_467,In_737);
and U2756 (N_2756,In_584,In_594);
nor U2757 (N_2757,In_991,In_683);
or U2758 (N_2758,In_977,In_782);
and U2759 (N_2759,In_792,In_603);
nor U2760 (N_2760,In_414,In_82);
nor U2761 (N_2761,In_71,In_533);
nand U2762 (N_2762,In_94,In_173);
nor U2763 (N_2763,In_861,In_842);
nand U2764 (N_2764,In_679,In_115);
or U2765 (N_2765,In_785,In_290);
nand U2766 (N_2766,In_689,In_883);
or U2767 (N_2767,In_535,In_37);
nand U2768 (N_2768,In_870,In_346);
and U2769 (N_2769,In_307,In_326);
and U2770 (N_2770,In_86,In_328);
or U2771 (N_2771,In_799,In_685);
nand U2772 (N_2772,In_459,In_158);
xnor U2773 (N_2773,In_374,In_70);
nand U2774 (N_2774,In_226,In_986);
nand U2775 (N_2775,In_636,In_504);
nand U2776 (N_2776,In_190,In_66);
and U2777 (N_2777,In_825,In_106);
nand U2778 (N_2778,In_140,In_531);
xnor U2779 (N_2779,In_593,In_941);
or U2780 (N_2780,In_832,In_565);
and U2781 (N_2781,In_359,In_770);
and U2782 (N_2782,In_177,In_226);
and U2783 (N_2783,In_743,In_464);
nor U2784 (N_2784,In_942,In_865);
nand U2785 (N_2785,In_616,In_315);
nand U2786 (N_2786,In_894,In_686);
xor U2787 (N_2787,In_956,In_203);
and U2788 (N_2788,In_639,In_555);
or U2789 (N_2789,In_295,In_556);
or U2790 (N_2790,In_870,In_936);
or U2791 (N_2791,In_529,In_913);
and U2792 (N_2792,In_660,In_430);
nor U2793 (N_2793,In_141,In_640);
nor U2794 (N_2794,In_926,In_662);
or U2795 (N_2795,In_400,In_911);
xor U2796 (N_2796,In_573,In_931);
or U2797 (N_2797,In_454,In_819);
or U2798 (N_2798,In_479,In_631);
and U2799 (N_2799,In_584,In_817);
or U2800 (N_2800,In_107,In_959);
xnor U2801 (N_2801,In_380,In_15);
nand U2802 (N_2802,In_440,In_511);
nor U2803 (N_2803,In_659,In_719);
nor U2804 (N_2804,In_611,In_281);
or U2805 (N_2805,In_402,In_800);
xnor U2806 (N_2806,In_278,In_543);
nand U2807 (N_2807,In_767,In_486);
or U2808 (N_2808,In_245,In_432);
or U2809 (N_2809,In_4,In_112);
or U2810 (N_2810,In_225,In_276);
nand U2811 (N_2811,In_102,In_97);
xnor U2812 (N_2812,In_259,In_943);
and U2813 (N_2813,In_875,In_323);
or U2814 (N_2814,In_641,In_291);
nor U2815 (N_2815,In_536,In_102);
or U2816 (N_2816,In_184,In_557);
xnor U2817 (N_2817,In_128,In_437);
nor U2818 (N_2818,In_646,In_500);
or U2819 (N_2819,In_292,In_651);
nor U2820 (N_2820,In_134,In_436);
and U2821 (N_2821,In_911,In_642);
nor U2822 (N_2822,In_530,In_579);
nor U2823 (N_2823,In_910,In_992);
nand U2824 (N_2824,In_402,In_354);
nand U2825 (N_2825,In_999,In_772);
nor U2826 (N_2826,In_309,In_216);
nand U2827 (N_2827,In_296,In_992);
and U2828 (N_2828,In_943,In_815);
nor U2829 (N_2829,In_932,In_558);
and U2830 (N_2830,In_872,In_953);
and U2831 (N_2831,In_939,In_382);
or U2832 (N_2832,In_784,In_322);
or U2833 (N_2833,In_335,In_770);
xnor U2834 (N_2834,In_385,In_93);
xor U2835 (N_2835,In_289,In_776);
nand U2836 (N_2836,In_429,In_731);
or U2837 (N_2837,In_93,In_241);
nand U2838 (N_2838,In_203,In_586);
or U2839 (N_2839,In_26,In_771);
nor U2840 (N_2840,In_848,In_733);
xnor U2841 (N_2841,In_371,In_298);
or U2842 (N_2842,In_860,In_543);
or U2843 (N_2843,In_212,In_171);
or U2844 (N_2844,In_755,In_381);
or U2845 (N_2845,In_724,In_438);
or U2846 (N_2846,In_685,In_403);
nand U2847 (N_2847,In_356,In_995);
nand U2848 (N_2848,In_828,In_302);
nor U2849 (N_2849,In_872,In_442);
nor U2850 (N_2850,In_238,In_588);
and U2851 (N_2851,In_695,In_466);
and U2852 (N_2852,In_155,In_820);
nand U2853 (N_2853,In_464,In_760);
and U2854 (N_2854,In_379,In_200);
nand U2855 (N_2855,In_705,In_845);
nor U2856 (N_2856,In_789,In_7);
or U2857 (N_2857,In_978,In_844);
nand U2858 (N_2858,In_594,In_998);
nand U2859 (N_2859,In_668,In_674);
nand U2860 (N_2860,In_159,In_641);
nand U2861 (N_2861,In_257,In_19);
nand U2862 (N_2862,In_228,In_714);
nor U2863 (N_2863,In_610,In_1);
nor U2864 (N_2864,In_261,In_563);
nand U2865 (N_2865,In_281,In_446);
nand U2866 (N_2866,In_356,In_899);
or U2867 (N_2867,In_558,In_98);
xnor U2868 (N_2868,In_447,In_732);
nor U2869 (N_2869,In_673,In_822);
or U2870 (N_2870,In_424,In_303);
nor U2871 (N_2871,In_965,In_17);
and U2872 (N_2872,In_707,In_31);
or U2873 (N_2873,In_365,In_902);
nor U2874 (N_2874,In_276,In_140);
and U2875 (N_2875,In_395,In_310);
nand U2876 (N_2876,In_546,In_657);
xor U2877 (N_2877,In_933,In_221);
nand U2878 (N_2878,In_587,In_623);
or U2879 (N_2879,In_62,In_399);
nand U2880 (N_2880,In_583,In_902);
or U2881 (N_2881,In_421,In_931);
nand U2882 (N_2882,In_87,In_899);
nor U2883 (N_2883,In_672,In_322);
nand U2884 (N_2884,In_257,In_27);
nand U2885 (N_2885,In_202,In_848);
nor U2886 (N_2886,In_426,In_892);
and U2887 (N_2887,In_109,In_388);
nor U2888 (N_2888,In_227,In_757);
nor U2889 (N_2889,In_73,In_685);
and U2890 (N_2890,In_562,In_613);
xor U2891 (N_2891,In_230,In_784);
nand U2892 (N_2892,In_950,In_818);
nor U2893 (N_2893,In_411,In_50);
nand U2894 (N_2894,In_25,In_963);
nand U2895 (N_2895,In_834,In_629);
xnor U2896 (N_2896,In_845,In_322);
or U2897 (N_2897,In_682,In_324);
and U2898 (N_2898,In_268,In_469);
or U2899 (N_2899,In_694,In_245);
nor U2900 (N_2900,In_121,In_144);
and U2901 (N_2901,In_285,In_545);
nor U2902 (N_2902,In_298,In_651);
or U2903 (N_2903,In_991,In_395);
nor U2904 (N_2904,In_528,In_425);
xor U2905 (N_2905,In_369,In_88);
nor U2906 (N_2906,In_347,In_540);
or U2907 (N_2907,In_395,In_117);
nor U2908 (N_2908,In_909,In_433);
nor U2909 (N_2909,In_849,In_360);
or U2910 (N_2910,In_908,In_238);
nor U2911 (N_2911,In_376,In_380);
or U2912 (N_2912,In_148,In_198);
nand U2913 (N_2913,In_642,In_584);
and U2914 (N_2914,In_866,In_632);
nor U2915 (N_2915,In_924,In_307);
nand U2916 (N_2916,In_853,In_201);
and U2917 (N_2917,In_173,In_867);
or U2918 (N_2918,In_306,In_474);
nor U2919 (N_2919,In_704,In_615);
and U2920 (N_2920,In_22,In_761);
and U2921 (N_2921,In_14,In_588);
or U2922 (N_2922,In_992,In_787);
and U2923 (N_2923,In_836,In_435);
and U2924 (N_2924,In_19,In_701);
and U2925 (N_2925,In_999,In_81);
and U2926 (N_2926,In_388,In_283);
nand U2927 (N_2927,In_141,In_352);
or U2928 (N_2928,In_252,In_613);
or U2929 (N_2929,In_38,In_98);
nor U2930 (N_2930,In_625,In_144);
xor U2931 (N_2931,In_795,In_329);
and U2932 (N_2932,In_244,In_785);
nor U2933 (N_2933,In_740,In_161);
and U2934 (N_2934,In_335,In_416);
or U2935 (N_2935,In_599,In_703);
nor U2936 (N_2936,In_833,In_857);
nand U2937 (N_2937,In_471,In_102);
nand U2938 (N_2938,In_761,In_865);
and U2939 (N_2939,In_526,In_323);
or U2940 (N_2940,In_983,In_624);
and U2941 (N_2941,In_721,In_297);
nand U2942 (N_2942,In_838,In_934);
xnor U2943 (N_2943,In_80,In_268);
and U2944 (N_2944,In_373,In_312);
or U2945 (N_2945,In_366,In_868);
xor U2946 (N_2946,In_165,In_948);
nand U2947 (N_2947,In_456,In_432);
and U2948 (N_2948,In_204,In_466);
nand U2949 (N_2949,In_479,In_637);
nand U2950 (N_2950,In_991,In_843);
or U2951 (N_2951,In_806,In_115);
nand U2952 (N_2952,In_676,In_131);
or U2953 (N_2953,In_528,In_994);
xnor U2954 (N_2954,In_951,In_865);
nor U2955 (N_2955,In_924,In_81);
nand U2956 (N_2956,In_609,In_149);
and U2957 (N_2957,In_687,In_192);
nor U2958 (N_2958,In_362,In_168);
nand U2959 (N_2959,In_873,In_888);
nand U2960 (N_2960,In_502,In_877);
nand U2961 (N_2961,In_466,In_133);
xnor U2962 (N_2962,In_906,In_593);
nor U2963 (N_2963,In_685,In_400);
nand U2964 (N_2964,In_70,In_604);
or U2965 (N_2965,In_119,In_678);
nor U2966 (N_2966,In_301,In_250);
nor U2967 (N_2967,In_716,In_451);
nand U2968 (N_2968,In_655,In_74);
and U2969 (N_2969,In_335,In_231);
nand U2970 (N_2970,In_969,In_688);
or U2971 (N_2971,In_157,In_405);
or U2972 (N_2972,In_259,In_370);
xor U2973 (N_2973,In_6,In_996);
nand U2974 (N_2974,In_352,In_473);
or U2975 (N_2975,In_322,In_795);
nand U2976 (N_2976,In_652,In_336);
and U2977 (N_2977,In_194,In_245);
nand U2978 (N_2978,In_768,In_420);
nand U2979 (N_2979,In_730,In_537);
xnor U2980 (N_2980,In_885,In_613);
nand U2981 (N_2981,In_238,In_606);
and U2982 (N_2982,In_586,In_357);
and U2983 (N_2983,In_606,In_399);
xnor U2984 (N_2984,In_36,In_318);
nor U2985 (N_2985,In_335,In_366);
or U2986 (N_2986,In_299,In_99);
nor U2987 (N_2987,In_749,In_93);
and U2988 (N_2988,In_423,In_654);
or U2989 (N_2989,In_2,In_330);
or U2990 (N_2990,In_851,In_64);
and U2991 (N_2991,In_219,In_997);
or U2992 (N_2992,In_532,In_552);
nor U2993 (N_2993,In_369,In_914);
and U2994 (N_2994,In_308,In_740);
nand U2995 (N_2995,In_48,In_617);
xor U2996 (N_2996,In_358,In_489);
xor U2997 (N_2997,In_440,In_140);
and U2998 (N_2998,In_678,In_756);
nand U2999 (N_2999,In_520,In_720);
nor U3000 (N_3000,In_942,In_479);
and U3001 (N_3001,In_519,In_998);
nand U3002 (N_3002,In_193,In_507);
or U3003 (N_3003,In_311,In_751);
or U3004 (N_3004,In_995,In_355);
or U3005 (N_3005,In_294,In_944);
or U3006 (N_3006,In_277,In_491);
nor U3007 (N_3007,In_913,In_928);
or U3008 (N_3008,In_829,In_599);
nand U3009 (N_3009,In_512,In_843);
xor U3010 (N_3010,In_832,In_405);
nor U3011 (N_3011,In_126,In_728);
nand U3012 (N_3012,In_176,In_425);
or U3013 (N_3013,In_183,In_301);
and U3014 (N_3014,In_508,In_518);
nor U3015 (N_3015,In_840,In_208);
nand U3016 (N_3016,In_379,In_971);
or U3017 (N_3017,In_117,In_791);
or U3018 (N_3018,In_908,In_821);
nor U3019 (N_3019,In_631,In_965);
and U3020 (N_3020,In_740,In_418);
and U3021 (N_3021,In_940,In_221);
nand U3022 (N_3022,In_730,In_947);
nor U3023 (N_3023,In_776,In_411);
or U3024 (N_3024,In_952,In_420);
or U3025 (N_3025,In_188,In_718);
nand U3026 (N_3026,In_439,In_159);
and U3027 (N_3027,In_389,In_146);
or U3028 (N_3028,In_466,In_251);
or U3029 (N_3029,In_285,In_316);
xor U3030 (N_3030,In_81,In_180);
nor U3031 (N_3031,In_420,In_95);
or U3032 (N_3032,In_753,In_717);
and U3033 (N_3033,In_607,In_737);
or U3034 (N_3034,In_781,In_117);
or U3035 (N_3035,In_203,In_978);
or U3036 (N_3036,In_408,In_326);
nand U3037 (N_3037,In_76,In_55);
nand U3038 (N_3038,In_398,In_669);
nand U3039 (N_3039,In_647,In_581);
and U3040 (N_3040,In_992,In_218);
nor U3041 (N_3041,In_300,In_412);
nor U3042 (N_3042,In_935,In_235);
or U3043 (N_3043,In_382,In_933);
nor U3044 (N_3044,In_322,In_892);
and U3045 (N_3045,In_688,In_163);
and U3046 (N_3046,In_88,In_79);
nor U3047 (N_3047,In_103,In_567);
nand U3048 (N_3048,In_209,In_715);
nor U3049 (N_3049,In_663,In_481);
nand U3050 (N_3050,In_8,In_576);
and U3051 (N_3051,In_191,In_952);
and U3052 (N_3052,In_742,In_71);
xnor U3053 (N_3053,In_448,In_280);
xor U3054 (N_3054,In_610,In_148);
or U3055 (N_3055,In_420,In_879);
nor U3056 (N_3056,In_256,In_507);
or U3057 (N_3057,In_770,In_337);
nand U3058 (N_3058,In_914,In_733);
nand U3059 (N_3059,In_83,In_770);
or U3060 (N_3060,In_876,In_215);
xor U3061 (N_3061,In_900,In_653);
or U3062 (N_3062,In_698,In_649);
nor U3063 (N_3063,In_27,In_731);
or U3064 (N_3064,In_589,In_56);
nor U3065 (N_3065,In_913,In_920);
and U3066 (N_3066,In_337,In_636);
and U3067 (N_3067,In_95,In_891);
and U3068 (N_3068,In_171,In_91);
nor U3069 (N_3069,In_121,In_774);
xor U3070 (N_3070,In_636,In_485);
nand U3071 (N_3071,In_454,In_462);
nand U3072 (N_3072,In_893,In_103);
or U3073 (N_3073,In_565,In_795);
and U3074 (N_3074,In_428,In_146);
and U3075 (N_3075,In_342,In_963);
and U3076 (N_3076,In_908,In_60);
nand U3077 (N_3077,In_638,In_166);
nor U3078 (N_3078,In_696,In_812);
or U3079 (N_3079,In_97,In_305);
and U3080 (N_3080,In_576,In_161);
and U3081 (N_3081,In_101,In_517);
and U3082 (N_3082,In_766,In_770);
nand U3083 (N_3083,In_865,In_19);
xnor U3084 (N_3084,In_979,In_454);
and U3085 (N_3085,In_288,In_932);
nand U3086 (N_3086,In_650,In_985);
nor U3087 (N_3087,In_530,In_138);
or U3088 (N_3088,In_194,In_478);
nor U3089 (N_3089,In_164,In_578);
or U3090 (N_3090,In_181,In_562);
or U3091 (N_3091,In_85,In_734);
nand U3092 (N_3092,In_96,In_166);
nand U3093 (N_3093,In_579,In_469);
xnor U3094 (N_3094,In_182,In_328);
and U3095 (N_3095,In_705,In_409);
nand U3096 (N_3096,In_518,In_700);
xor U3097 (N_3097,In_533,In_42);
nor U3098 (N_3098,In_819,In_596);
and U3099 (N_3099,In_487,In_239);
nor U3100 (N_3100,In_293,In_508);
or U3101 (N_3101,In_99,In_914);
nand U3102 (N_3102,In_532,In_362);
and U3103 (N_3103,In_879,In_276);
nor U3104 (N_3104,In_267,In_101);
nor U3105 (N_3105,In_575,In_691);
nand U3106 (N_3106,In_474,In_764);
nand U3107 (N_3107,In_47,In_169);
nor U3108 (N_3108,In_16,In_533);
or U3109 (N_3109,In_946,In_780);
nand U3110 (N_3110,In_651,In_314);
nand U3111 (N_3111,In_890,In_94);
nand U3112 (N_3112,In_767,In_772);
or U3113 (N_3113,In_24,In_213);
nand U3114 (N_3114,In_594,In_0);
xnor U3115 (N_3115,In_490,In_516);
and U3116 (N_3116,In_22,In_340);
nand U3117 (N_3117,In_531,In_274);
and U3118 (N_3118,In_659,In_542);
and U3119 (N_3119,In_647,In_733);
xor U3120 (N_3120,In_716,In_488);
nand U3121 (N_3121,In_792,In_811);
nor U3122 (N_3122,In_813,In_64);
nor U3123 (N_3123,In_67,In_9);
or U3124 (N_3124,In_140,In_766);
xor U3125 (N_3125,In_57,In_973);
xnor U3126 (N_3126,In_145,In_398);
nand U3127 (N_3127,In_70,In_448);
nand U3128 (N_3128,In_501,In_996);
or U3129 (N_3129,In_574,In_993);
nor U3130 (N_3130,In_494,In_845);
or U3131 (N_3131,In_195,In_774);
and U3132 (N_3132,In_646,In_747);
or U3133 (N_3133,In_694,In_500);
or U3134 (N_3134,In_588,In_723);
nand U3135 (N_3135,In_821,In_831);
nand U3136 (N_3136,In_350,In_853);
nor U3137 (N_3137,In_708,In_504);
or U3138 (N_3138,In_951,In_327);
and U3139 (N_3139,In_858,In_18);
or U3140 (N_3140,In_604,In_362);
nor U3141 (N_3141,In_768,In_396);
and U3142 (N_3142,In_720,In_980);
nor U3143 (N_3143,In_136,In_109);
nor U3144 (N_3144,In_402,In_913);
nor U3145 (N_3145,In_464,In_210);
nor U3146 (N_3146,In_219,In_424);
nand U3147 (N_3147,In_633,In_530);
or U3148 (N_3148,In_377,In_693);
nor U3149 (N_3149,In_30,In_316);
nor U3150 (N_3150,In_617,In_752);
and U3151 (N_3151,In_222,In_649);
and U3152 (N_3152,In_345,In_919);
and U3153 (N_3153,In_607,In_75);
or U3154 (N_3154,In_260,In_628);
nor U3155 (N_3155,In_199,In_311);
nand U3156 (N_3156,In_100,In_357);
and U3157 (N_3157,In_132,In_994);
nor U3158 (N_3158,In_585,In_413);
nor U3159 (N_3159,In_525,In_181);
nand U3160 (N_3160,In_786,In_967);
or U3161 (N_3161,In_762,In_91);
and U3162 (N_3162,In_376,In_456);
xnor U3163 (N_3163,In_624,In_583);
nor U3164 (N_3164,In_917,In_333);
nand U3165 (N_3165,In_995,In_429);
xor U3166 (N_3166,In_334,In_558);
nand U3167 (N_3167,In_833,In_954);
nor U3168 (N_3168,In_67,In_862);
nand U3169 (N_3169,In_293,In_882);
or U3170 (N_3170,In_82,In_865);
nand U3171 (N_3171,In_493,In_743);
or U3172 (N_3172,In_957,In_404);
nand U3173 (N_3173,In_967,In_946);
nor U3174 (N_3174,In_886,In_29);
or U3175 (N_3175,In_316,In_20);
and U3176 (N_3176,In_313,In_513);
or U3177 (N_3177,In_772,In_790);
nor U3178 (N_3178,In_44,In_389);
or U3179 (N_3179,In_235,In_632);
or U3180 (N_3180,In_892,In_487);
or U3181 (N_3181,In_310,In_619);
nand U3182 (N_3182,In_224,In_13);
nand U3183 (N_3183,In_885,In_469);
nand U3184 (N_3184,In_191,In_821);
or U3185 (N_3185,In_221,In_53);
nand U3186 (N_3186,In_573,In_523);
and U3187 (N_3187,In_795,In_911);
and U3188 (N_3188,In_1,In_747);
nand U3189 (N_3189,In_851,In_573);
nand U3190 (N_3190,In_186,In_491);
xnor U3191 (N_3191,In_915,In_953);
xnor U3192 (N_3192,In_380,In_238);
nand U3193 (N_3193,In_562,In_997);
nor U3194 (N_3194,In_83,In_986);
xor U3195 (N_3195,In_213,In_534);
or U3196 (N_3196,In_958,In_393);
and U3197 (N_3197,In_90,In_190);
or U3198 (N_3198,In_484,In_594);
or U3199 (N_3199,In_95,In_854);
or U3200 (N_3200,In_126,In_40);
nand U3201 (N_3201,In_550,In_88);
nor U3202 (N_3202,In_150,In_595);
or U3203 (N_3203,In_697,In_289);
xnor U3204 (N_3204,In_209,In_835);
xor U3205 (N_3205,In_743,In_202);
and U3206 (N_3206,In_17,In_91);
and U3207 (N_3207,In_873,In_785);
nor U3208 (N_3208,In_80,In_842);
nor U3209 (N_3209,In_427,In_21);
nor U3210 (N_3210,In_824,In_7);
nor U3211 (N_3211,In_265,In_575);
or U3212 (N_3212,In_835,In_942);
or U3213 (N_3213,In_472,In_655);
nand U3214 (N_3214,In_26,In_388);
or U3215 (N_3215,In_149,In_974);
and U3216 (N_3216,In_210,In_700);
nand U3217 (N_3217,In_537,In_505);
and U3218 (N_3218,In_155,In_439);
nand U3219 (N_3219,In_131,In_259);
and U3220 (N_3220,In_501,In_957);
nand U3221 (N_3221,In_545,In_758);
and U3222 (N_3222,In_760,In_27);
nor U3223 (N_3223,In_122,In_443);
nor U3224 (N_3224,In_616,In_112);
and U3225 (N_3225,In_863,In_218);
nand U3226 (N_3226,In_813,In_443);
and U3227 (N_3227,In_341,In_409);
xnor U3228 (N_3228,In_527,In_730);
or U3229 (N_3229,In_762,In_134);
and U3230 (N_3230,In_998,In_852);
and U3231 (N_3231,In_922,In_876);
xnor U3232 (N_3232,In_233,In_541);
and U3233 (N_3233,In_25,In_757);
and U3234 (N_3234,In_5,In_524);
nor U3235 (N_3235,In_551,In_969);
nand U3236 (N_3236,In_75,In_197);
nand U3237 (N_3237,In_614,In_226);
nand U3238 (N_3238,In_897,In_340);
and U3239 (N_3239,In_68,In_686);
xnor U3240 (N_3240,In_447,In_934);
or U3241 (N_3241,In_395,In_244);
nand U3242 (N_3242,In_274,In_605);
nand U3243 (N_3243,In_532,In_191);
nand U3244 (N_3244,In_644,In_68);
nor U3245 (N_3245,In_573,In_434);
nand U3246 (N_3246,In_339,In_725);
xor U3247 (N_3247,In_800,In_408);
nand U3248 (N_3248,In_879,In_685);
nor U3249 (N_3249,In_421,In_251);
or U3250 (N_3250,In_573,In_545);
nor U3251 (N_3251,In_873,In_89);
nor U3252 (N_3252,In_956,In_116);
nor U3253 (N_3253,In_966,In_394);
nor U3254 (N_3254,In_989,In_323);
nor U3255 (N_3255,In_455,In_829);
and U3256 (N_3256,In_792,In_979);
nand U3257 (N_3257,In_558,In_557);
or U3258 (N_3258,In_282,In_718);
nor U3259 (N_3259,In_604,In_619);
or U3260 (N_3260,In_831,In_635);
nand U3261 (N_3261,In_374,In_611);
nor U3262 (N_3262,In_366,In_869);
nand U3263 (N_3263,In_995,In_861);
or U3264 (N_3264,In_997,In_792);
nand U3265 (N_3265,In_211,In_419);
nor U3266 (N_3266,In_192,In_287);
nand U3267 (N_3267,In_153,In_752);
or U3268 (N_3268,In_925,In_705);
nor U3269 (N_3269,In_564,In_921);
and U3270 (N_3270,In_634,In_115);
nand U3271 (N_3271,In_915,In_356);
and U3272 (N_3272,In_587,In_720);
or U3273 (N_3273,In_896,In_389);
nor U3274 (N_3274,In_905,In_523);
nor U3275 (N_3275,In_763,In_885);
xor U3276 (N_3276,In_772,In_829);
nand U3277 (N_3277,In_21,In_615);
and U3278 (N_3278,In_116,In_970);
and U3279 (N_3279,In_42,In_254);
nand U3280 (N_3280,In_93,In_92);
nor U3281 (N_3281,In_319,In_231);
or U3282 (N_3282,In_569,In_513);
or U3283 (N_3283,In_113,In_299);
or U3284 (N_3284,In_16,In_714);
and U3285 (N_3285,In_650,In_33);
and U3286 (N_3286,In_348,In_678);
or U3287 (N_3287,In_970,In_756);
and U3288 (N_3288,In_548,In_139);
nor U3289 (N_3289,In_537,In_238);
nand U3290 (N_3290,In_504,In_687);
and U3291 (N_3291,In_587,In_498);
and U3292 (N_3292,In_357,In_283);
nand U3293 (N_3293,In_278,In_173);
nand U3294 (N_3294,In_658,In_233);
nand U3295 (N_3295,In_953,In_848);
xnor U3296 (N_3296,In_50,In_702);
or U3297 (N_3297,In_172,In_613);
nor U3298 (N_3298,In_699,In_917);
nor U3299 (N_3299,In_39,In_527);
or U3300 (N_3300,In_841,In_328);
xnor U3301 (N_3301,In_952,In_351);
xnor U3302 (N_3302,In_869,In_220);
and U3303 (N_3303,In_700,In_101);
or U3304 (N_3304,In_537,In_289);
or U3305 (N_3305,In_85,In_542);
nand U3306 (N_3306,In_408,In_548);
nand U3307 (N_3307,In_446,In_535);
xor U3308 (N_3308,In_691,In_805);
or U3309 (N_3309,In_499,In_901);
or U3310 (N_3310,In_101,In_328);
nor U3311 (N_3311,In_390,In_49);
or U3312 (N_3312,In_227,In_651);
nand U3313 (N_3313,In_349,In_198);
or U3314 (N_3314,In_210,In_454);
nand U3315 (N_3315,In_625,In_153);
nand U3316 (N_3316,In_253,In_640);
nand U3317 (N_3317,In_629,In_538);
nand U3318 (N_3318,In_776,In_277);
nor U3319 (N_3319,In_138,In_118);
or U3320 (N_3320,In_283,In_987);
and U3321 (N_3321,In_71,In_385);
and U3322 (N_3322,In_833,In_267);
or U3323 (N_3323,In_924,In_123);
nand U3324 (N_3324,In_979,In_834);
and U3325 (N_3325,In_553,In_27);
nand U3326 (N_3326,In_220,In_841);
nor U3327 (N_3327,In_296,In_251);
nand U3328 (N_3328,In_563,In_394);
or U3329 (N_3329,In_396,In_817);
and U3330 (N_3330,In_561,In_619);
nand U3331 (N_3331,In_942,In_25);
nand U3332 (N_3332,In_874,In_579);
nor U3333 (N_3333,In_448,In_784);
or U3334 (N_3334,In_425,In_197);
nor U3335 (N_3335,In_566,In_561);
nand U3336 (N_3336,In_429,In_436);
and U3337 (N_3337,In_952,In_586);
xor U3338 (N_3338,In_226,In_456);
and U3339 (N_3339,In_634,In_344);
and U3340 (N_3340,In_325,In_588);
nor U3341 (N_3341,In_981,In_938);
nor U3342 (N_3342,In_578,In_990);
nand U3343 (N_3343,In_90,In_761);
and U3344 (N_3344,In_267,In_260);
and U3345 (N_3345,In_554,In_229);
or U3346 (N_3346,In_917,In_85);
nor U3347 (N_3347,In_553,In_693);
or U3348 (N_3348,In_763,In_966);
nand U3349 (N_3349,In_70,In_989);
and U3350 (N_3350,In_892,In_969);
or U3351 (N_3351,In_718,In_799);
or U3352 (N_3352,In_11,In_930);
nand U3353 (N_3353,In_272,In_960);
nor U3354 (N_3354,In_931,In_498);
nand U3355 (N_3355,In_342,In_244);
xnor U3356 (N_3356,In_574,In_763);
and U3357 (N_3357,In_661,In_138);
nor U3358 (N_3358,In_206,In_995);
or U3359 (N_3359,In_77,In_285);
or U3360 (N_3360,In_592,In_116);
nor U3361 (N_3361,In_277,In_276);
xnor U3362 (N_3362,In_957,In_247);
nand U3363 (N_3363,In_585,In_545);
nand U3364 (N_3364,In_449,In_646);
nand U3365 (N_3365,In_852,In_727);
nor U3366 (N_3366,In_729,In_660);
nand U3367 (N_3367,In_478,In_136);
or U3368 (N_3368,In_545,In_182);
or U3369 (N_3369,In_591,In_53);
and U3370 (N_3370,In_313,In_102);
xnor U3371 (N_3371,In_809,In_169);
nor U3372 (N_3372,In_835,In_596);
nor U3373 (N_3373,In_125,In_681);
or U3374 (N_3374,In_552,In_598);
nor U3375 (N_3375,In_308,In_572);
and U3376 (N_3376,In_674,In_461);
and U3377 (N_3377,In_618,In_966);
xnor U3378 (N_3378,In_473,In_962);
nor U3379 (N_3379,In_646,In_853);
and U3380 (N_3380,In_807,In_303);
and U3381 (N_3381,In_873,In_876);
nor U3382 (N_3382,In_901,In_34);
xnor U3383 (N_3383,In_470,In_985);
and U3384 (N_3384,In_803,In_239);
and U3385 (N_3385,In_356,In_571);
xnor U3386 (N_3386,In_42,In_797);
nor U3387 (N_3387,In_915,In_860);
nor U3388 (N_3388,In_747,In_255);
or U3389 (N_3389,In_381,In_81);
or U3390 (N_3390,In_268,In_0);
nand U3391 (N_3391,In_252,In_662);
xnor U3392 (N_3392,In_646,In_463);
nor U3393 (N_3393,In_903,In_964);
nor U3394 (N_3394,In_160,In_21);
nor U3395 (N_3395,In_775,In_876);
and U3396 (N_3396,In_223,In_57);
nand U3397 (N_3397,In_867,In_554);
or U3398 (N_3398,In_224,In_568);
nor U3399 (N_3399,In_310,In_494);
and U3400 (N_3400,In_187,In_993);
nor U3401 (N_3401,In_894,In_646);
and U3402 (N_3402,In_130,In_341);
or U3403 (N_3403,In_471,In_165);
xor U3404 (N_3404,In_753,In_1);
or U3405 (N_3405,In_176,In_738);
nand U3406 (N_3406,In_153,In_289);
nand U3407 (N_3407,In_179,In_807);
nor U3408 (N_3408,In_525,In_655);
and U3409 (N_3409,In_821,In_890);
nor U3410 (N_3410,In_933,In_305);
xor U3411 (N_3411,In_280,In_409);
nand U3412 (N_3412,In_209,In_778);
or U3413 (N_3413,In_844,In_870);
nand U3414 (N_3414,In_805,In_125);
or U3415 (N_3415,In_778,In_914);
and U3416 (N_3416,In_273,In_173);
nor U3417 (N_3417,In_894,In_155);
xnor U3418 (N_3418,In_708,In_479);
xnor U3419 (N_3419,In_514,In_971);
and U3420 (N_3420,In_216,In_276);
nand U3421 (N_3421,In_614,In_434);
or U3422 (N_3422,In_742,In_131);
nor U3423 (N_3423,In_636,In_946);
nor U3424 (N_3424,In_747,In_807);
nand U3425 (N_3425,In_22,In_381);
nor U3426 (N_3426,In_946,In_833);
or U3427 (N_3427,In_689,In_136);
nand U3428 (N_3428,In_680,In_855);
xnor U3429 (N_3429,In_358,In_325);
and U3430 (N_3430,In_90,In_492);
nand U3431 (N_3431,In_446,In_212);
nor U3432 (N_3432,In_442,In_852);
nand U3433 (N_3433,In_796,In_436);
and U3434 (N_3434,In_260,In_8);
and U3435 (N_3435,In_824,In_510);
nor U3436 (N_3436,In_275,In_972);
nor U3437 (N_3437,In_273,In_417);
nor U3438 (N_3438,In_863,In_295);
nor U3439 (N_3439,In_965,In_856);
nor U3440 (N_3440,In_396,In_474);
or U3441 (N_3441,In_875,In_792);
or U3442 (N_3442,In_235,In_337);
and U3443 (N_3443,In_371,In_206);
or U3444 (N_3444,In_294,In_29);
nor U3445 (N_3445,In_876,In_544);
xnor U3446 (N_3446,In_857,In_323);
xnor U3447 (N_3447,In_518,In_903);
and U3448 (N_3448,In_433,In_525);
nand U3449 (N_3449,In_363,In_829);
xor U3450 (N_3450,In_499,In_324);
and U3451 (N_3451,In_696,In_406);
nor U3452 (N_3452,In_559,In_446);
or U3453 (N_3453,In_923,In_677);
nor U3454 (N_3454,In_31,In_311);
and U3455 (N_3455,In_532,In_275);
and U3456 (N_3456,In_9,In_727);
and U3457 (N_3457,In_28,In_878);
nand U3458 (N_3458,In_238,In_90);
nor U3459 (N_3459,In_840,In_423);
nand U3460 (N_3460,In_384,In_288);
nor U3461 (N_3461,In_22,In_235);
xnor U3462 (N_3462,In_904,In_335);
or U3463 (N_3463,In_896,In_226);
and U3464 (N_3464,In_814,In_402);
or U3465 (N_3465,In_906,In_475);
nor U3466 (N_3466,In_491,In_769);
or U3467 (N_3467,In_394,In_42);
or U3468 (N_3468,In_188,In_584);
nand U3469 (N_3469,In_708,In_466);
and U3470 (N_3470,In_902,In_237);
and U3471 (N_3471,In_796,In_434);
or U3472 (N_3472,In_465,In_162);
xnor U3473 (N_3473,In_134,In_258);
and U3474 (N_3474,In_400,In_280);
or U3475 (N_3475,In_494,In_26);
nor U3476 (N_3476,In_834,In_745);
nand U3477 (N_3477,In_510,In_860);
xnor U3478 (N_3478,In_143,In_310);
and U3479 (N_3479,In_212,In_229);
and U3480 (N_3480,In_95,In_708);
and U3481 (N_3481,In_599,In_688);
xor U3482 (N_3482,In_22,In_49);
nand U3483 (N_3483,In_36,In_333);
or U3484 (N_3484,In_612,In_617);
and U3485 (N_3485,In_197,In_313);
or U3486 (N_3486,In_956,In_88);
nor U3487 (N_3487,In_874,In_810);
nand U3488 (N_3488,In_891,In_877);
and U3489 (N_3489,In_327,In_343);
and U3490 (N_3490,In_319,In_735);
nand U3491 (N_3491,In_818,In_460);
nor U3492 (N_3492,In_85,In_134);
or U3493 (N_3493,In_109,In_287);
nor U3494 (N_3494,In_307,In_861);
or U3495 (N_3495,In_6,In_647);
nand U3496 (N_3496,In_858,In_870);
nand U3497 (N_3497,In_883,In_30);
nand U3498 (N_3498,In_425,In_152);
and U3499 (N_3499,In_580,In_850);
nor U3500 (N_3500,In_955,In_728);
xnor U3501 (N_3501,In_711,In_467);
nand U3502 (N_3502,In_570,In_742);
and U3503 (N_3503,In_954,In_375);
and U3504 (N_3504,In_989,In_368);
or U3505 (N_3505,In_944,In_676);
or U3506 (N_3506,In_906,In_723);
nand U3507 (N_3507,In_240,In_87);
xnor U3508 (N_3508,In_856,In_364);
and U3509 (N_3509,In_897,In_471);
and U3510 (N_3510,In_511,In_745);
nand U3511 (N_3511,In_598,In_14);
and U3512 (N_3512,In_958,In_212);
or U3513 (N_3513,In_757,In_712);
or U3514 (N_3514,In_722,In_83);
nand U3515 (N_3515,In_842,In_813);
nand U3516 (N_3516,In_604,In_487);
and U3517 (N_3517,In_957,In_650);
xor U3518 (N_3518,In_338,In_370);
xnor U3519 (N_3519,In_391,In_344);
or U3520 (N_3520,In_663,In_497);
nor U3521 (N_3521,In_28,In_50);
nand U3522 (N_3522,In_415,In_337);
and U3523 (N_3523,In_841,In_646);
and U3524 (N_3524,In_924,In_466);
or U3525 (N_3525,In_931,In_560);
nand U3526 (N_3526,In_198,In_436);
nand U3527 (N_3527,In_580,In_75);
or U3528 (N_3528,In_201,In_252);
nor U3529 (N_3529,In_912,In_137);
nand U3530 (N_3530,In_380,In_786);
and U3531 (N_3531,In_245,In_343);
nand U3532 (N_3532,In_286,In_906);
or U3533 (N_3533,In_653,In_251);
or U3534 (N_3534,In_760,In_308);
nor U3535 (N_3535,In_891,In_853);
or U3536 (N_3536,In_158,In_190);
nand U3537 (N_3537,In_354,In_899);
xnor U3538 (N_3538,In_121,In_725);
nor U3539 (N_3539,In_301,In_872);
and U3540 (N_3540,In_550,In_378);
or U3541 (N_3541,In_74,In_120);
nand U3542 (N_3542,In_41,In_761);
nor U3543 (N_3543,In_405,In_309);
and U3544 (N_3544,In_730,In_432);
nand U3545 (N_3545,In_545,In_860);
and U3546 (N_3546,In_7,In_677);
nor U3547 (N_3547,In_343,In_272);
nor U3548 (N_3548,In_501,In_266);
nand U3549 (N_3549,In_271,In_835);
and U3550 (N_3550,In_835,In_475);
and U3551 (N_3551,In_97,In_856);
xnor U3552 (N_3552,In_166,In_286);
or U3553 (N_3553,In_800,In_879);
and U3554 (N_3554,In_767,In_979);
and U3555 (N_3555,In_38,In_857);
and U3556 (N_3556,In_0,In_173);
nor U3557 (N_3557,In_714,In_830);
nor U3558 (N_3558,In_758,In_43);
nor U3559 (N_3559,In_444,In_684);
xor U3560 (N_3560,In_472,In_264);
nor U3561 (N_3561,In_657,In_79);
or U3562 (N_3562,In_272,In_719);
nand U3563 (N_3563,In_259,In_242);
or U3564 (N_3564,In_889,In_206);
nor U3565 (N_3565,In_225,In_567);
nor U3566 (N_3566,In_456,In_95);
or U3567 (N_3567,In_165,In_381);
nand U3568 (N_3568,In_858,In_368);
nor U3569 (N_3569,In_153,In_825);
or U3570 (N_3570,In_315,In_159);
nand U3571 (N_3571,In_878,In_311);
and U3572 (N_3572,In_404,In_877);
nor U3573 (N_3573,In_804,In_59);
or U3574 (N_3574,In_773,In_275);
or U3575 (N_3575,In_380,In_270);
xor U3576 (N_3576,In_720,In_354);
and U3577 (N_3577,In_299,In_350);
xor U3578 (N_3578,In_620,In_330);
nand U3579 (N_3579,In_791,In_894);
nand U3580 (N_3580,In_169,In_76);
nand U3581 (N_3581,In_136,In_231);
nand U3582 (N_3582,In_571,In_8);
and U3583 (N_3583,In_342,In_425);
or U3584 (N_3584,In_821,In_394);
xnor U3585 (N_3585,In_730,In_850);
xnor U3586 (N_3586,In_902,In_885);
and U3587 (N_3587,In_638,In_711);
nand U3588 (N_3588,In_325,In_226);
nor U3589 (N_3589,In_442,In_491);
nor U3590 (N_3590,In_223,In_50);
or U3591 (N_3591,In_798,In_213);
nand U3592 (N_3592,In_868,In_469);
and U3593 (N_3593,In_909,In_521);
nor U3594 (N_3594,In_926,In_568);
nor U3595 (N_3595,In_556,In_644);
nand U3596 (N_3596,In_495,In_802);
and U3597 (N_3597,In_233,In_748);
nand U3598 (N_3598,In_447,In_221);
and U3599 (N_3599,In_348,In_792);
or U3600 (N_3600,In_737,In_808);
or U3601 (N_3601,In_580,In_530);
nor U3602 (N_3602,In_494,In_261);
or U3603 (N_3603,In_212,In_682);
and U3604 (N_3604,In_259,In_898);
nor U3605 (N_3605,In_830,In_178);
or U3606 (N_3606,In_101,In_168);
or U3607 (N_3607,In_672,In_99);
xnor U3608 (N_3608,In_795,In_984);
and U3609 (N_3609,In_82,In_233);
nand U3610 (N_3610,In_569,In_50);
nor U3611 (N_3611,In_72,In_703);
xnor U3612 (N_3612,In_29,In_658);
or U3613 (N_3613,In_870,In_210);
nor U3614 (N_3614,In_726,In_25);
nand U3615 (N_3615,In_856,In_80);
nand U3616 (N_3616,In_369,In_95);
and U3617 (N_3617,In_304,In_43);
nand U3618 (N_3618,In_147,In_666);
or U3619 (N_3619,In_454,In_697);
nor U3620 (N_3620,In_90,In_291);
and U3621 (N_3621,In_572,In_987);
nand U3622 (N_3622,In_393,In_889);
xor U3623 (N_3623,In_936,In_835);
nor U3624 (N_3624,In_833,In_279);
nor U3625 (N_3625,In_898,In_893);
nand U3626 (N_3626,In_881,In_650);
nor U3627 (N_3627,In_92,In_552);
and U3628 (N_3628,In_109,In_570);
xor U3629 (N_3629,In_107,In_490);
or U3630 (N_3630,In_535,In_993);
nand U3631 (N_3631,In_595,In_707);
nor U3632 (N_3632,In_86,In_336);
or U3633 (N_3633,In_338,In_327);
or U3634 (N_3634,In_441,In_708);
or U3635 (N_3635,In_372,In_695);
or U3636 (N_3636,In_740,In_111);
nand U3637 (N_3637,In_792,In_190);
or U3638 (N_3638,In_669,In_552);
xnor U3639 (N_3639,In_452,In_77);
or U3640 (N_3640,In_784,In_904);
and U3641 (N_3641,In_153,In_274);
and U3642 (N_3642,In_168,In_883);
or U3643 (N_3643,In_937,In_204);
or U3644 (N_3644,In_40,In_932);
or U3645 (N_3645,In_173,In_50);
nor U3646 (N_3646,In_105,In_936);
nor U3647 (N_3647,In_483,In_607);
nor U3648 (N_3648,In_600,In_191);
or U3649 (N_3649,In_139,In_79);
or U3650 (N_3650,In_255,In_666);
nor U3651 (N_3651,In_487,In_564);
nor U3652 (N_3652,In_975,In_613);
xor U3653 (N_3653,In_984,In_784);
xnor U3654 (N_3654,In_138,In_536);
nor U3655 (N_3655,In_706,In_193);
nand U3656 (N_3656,In_128,In_601);
nor U3657 (N_3657,In_539,In_866);
or U3658 (N_3658,In_896,In_265);
nor U3659 (N_3659,In_601,In_183);
or U3660 (N_3660,In_221,In_255);
or U3661 (N_3661,In_850,In_96);
nand U3662 (N_3662,In_20,In_404);
or U3663 (N_3663,In_718,In_649);
nand U3664 (N_3664,In_304,In_55);
or U3665 (N_3665,In_892,In_796);
and U3666 (N_3666,In_220,In_12);
or U3667 (N_3667,In_822,In_232);
nor U3668 (N_3668,In_451,In_23);
and U3669 (N_3669,In_150,In_447);
nor U3670 (N_3670,In_666,In_895);
nand U3671 (N_3671,In_801,In_60);
and U3672 (N_3672,In_25,In_492);
nor U3673 (N_3673,In_149,In_735);
nand U3674 (N_3674,In_820,In_459);
or U3675 (N_3675,In_672,In_595);
nand U3676 (N_3676,In_422,In_463);
nor U3677 (N_3677,In_350,In_417);
or U3678 (N_3678,In_658,In_106);
and U3679 (N_3679,In_13,In_698);
or U3680 (N_3680,In_2,In_667);
and U3681 (N_3681,In_964,In_726);
or U3682 (N_3682,In_571,In_40);
nor U3683 (N_3683,In_258,In_161);
or U3684 (N_3684,In_48,In_113);
nand U3685 (N_3685,In_184,In_555);
or U3686 (N_3686,In_803,In_969);
or U3687 (N_3687,In_143,In_225);
and U3688 (N_3688,In_936,In_355);
or U3689 (N_3689,In_67,In_687);
nand U3690 (N_3690,In_349,In_617);
nand U3691 (N_3691,In_496,In_635);
xor U3692 (N_3692,In_604,In_637);
nor U3693 (N_3693,In_249,In_875);
or U3694 (N_3694,In_376,In_978);
nand U3695 (N_3695,In_891,In_558);
and U3696 (N_3696,In_940,In_21);
nand U3697 (N_3697,In_942,In_490);
and U3698 (N_3698,In_976,In_141);
or U3699 (N_3699,In_52,In_756);
nor U3700 (N_3700,In_230,In_487);
nand U3701 (N_3701,In_585,In_351);
nand U3702 (N_3702,In_587,In_182);
or U3703 (N_3703,In_913,In_260);
nand U3704 (N_3704,In_647,In_83);
nand U3705 (N_3705,In_700,In_588);
nor U3706 (N_3706,In_591,In_933);
or U3707 (N_3707,In_688,In_774);
nor U3708 (N_3708,In_130,In_284);
xnor U3709 (N_3709,In_383,In_413);
and U3710 (N_3710,In_675,In_158);
nor U3711 (N_3711,In_749,In_673);
nand U3712 (N_3712,In_149,In_567);
nand U3713 (N_3713,In_460,In_253);
nor U3714 (N_3714,In_721,In_130);
xor U3715 (N_3715,In_244,In_723);
nor U3716 (N_3716,In_337,In_41);
nand U3717 (N_3717,In_514,In_622);
nor U3718 (N_3718,In_875,In_607);
nor U3719 (N_3719,In_297,In_21);
xnor U3720 (N_3720,In_24,In_422);
and U3721 (N_3721,In_900,In_631);
or U3722 (N_3722,In_137,In_106);
nand U3723 (N_3723,In_153,In_902);
nor U3724 (N_3724,In_102,In_58);
and U3725 (N_3725,In_390,In_974);
xnor U3726 (N_3726,In_304,In_404);
nor U3727 (N_3727,In_563,In_158);
or U3728 (N_3728,In_141,In_713);
or U3729 (N_3729,In_809,In_646);
or U3730 (N_3730,In_884,In_339);
nand U3731 (N_3731,In_661,In_937);
nor U3732 (N_3732,In_995,In_927);
and U3733 (N_3733,In_686,In_310);
and U3734 (N_3734,In_448,In_345);
or U3735 (N_3735,In_416,In_661);
nor U3736 (N_3736,In_511,In_700);
nor U3737 (N_3737,In_59,In_77);
nor U3738 (N_3738,In_362,In_167);
nand U3739 (N_3739,In_169,In_40);
nand U3740 (N_3740,In_911,In_567);
xor U3741 (N_3741,In_114,In_438);
or U3742 (N_3742,In_157,In_836);
nor U3743 (N_3743,In_796,In_223);
nand U3744 (N_3744,In_871,In_317);
nand U3745 (N_3745,In_766,In_516);
or U3746 (N_3746,In_24,In_744);
and U3747 (N_3747,In_616,In_998);
xor U3748 (N_3748,In_891,In_700);
or U3749 (N_3749,In_208,In_187);
nand U3750 (N_3750,In_259,In_715);
nor U3751 (N_3751,In_263,In_192);
or U3752 (N_3752,In_128,In_491);
nand U3753 (N_3753,In_171,In_617);
nand U3754 (N_3754,In_450,In_543);
or U3755 (N_3755,In_532,In_984);
and U3756 (N_3756,In_62,In_37);
nor U3757 (N_3757,In_577,In_738);
nor U3758 (N_3758,In_912,In_338);
and U3759 (N_3759,In_560,In_605);
nor U3760 (N_3760,In_159,In_958);
nor U3761 (N_3761,In_612,In_3);
or U3762 (N_3762,In_889,In_99);
xnor U3763 (N_3763,In_11,In_763);
and U3764 (N_3764,In_372,In_653);
nand U3765 (N_3765,In_532,In_414);
nor U3766 (N_3766,In_919,In_229);
xnor U3767 (N_3767,In_314,In_886);
nor U3768 (N_3768,In_271,In_553);
nor U3769 (N_3769,In_599,In_418);
nor U3770 (N_3770,In_412,In_849);
xor U3771 (N_3771,In_242,In_80);
nor U3772 (N_3772,In_582,In_424);
nor U3773 (N_3773,In_30,In_753);
nand U3774 (N_3774,In_696,In_375);
and U3775 (N_3775,In_944,In_684);
or U3776 (N_3776,In_905,In_470);
and U3777 (N_3777,In_557,In_163);
nand U3778 (N_3778,In_221,In_41);
nor U3779 (N_3779,In_300,In_943);
or U3780 (N_3780,In_696,In_483);
or U3781 (N_3781,In_397,In_812);
and U3782 (N_3782,In_138,In_994);
or U3783 (N_3783,In_344,In_891);
nand U3784 (N_3784,In_274,In_391);
nand U3785 (N_3785,In_398,In_799);
xnor U3786 (N_3786,In_151,In_440);
or U3787 (N_3787,In_740,In_763);
xor U3788 (N_3788,In_986,In_413);
nand U3789 (N_3789,In_270,In_630);
or U3790 (N_3790,In_273,In_387);
nor U3791 (N_3791,In_682,In_23);
xor U3792 (N_3792,In_579,In_274);
nand U3793 (N_3793,In_26,In_956);
and U3794 (N_3794,In_710,In_577);
xor U3795 (N_3795,In_460,In_322);
or U3796 (N_3796,In_423,In_470);
or U3797 (N_3797,In_964,In_926);
nor U3798 (N_3798,In_433,In_15);
or U3799 (N_3799,In_198,In_930);
or U3800 (N_3800,In_677,In_244);
nand U3801 (N_3801,In_727,In_369);
and U3802 (N_3802,In_833,In_908);
and U3803 (N_3803,In_462,In_43);
or U3804 (N_3804,In_659,In_569);
nor U3805 (N_3805,In_613,In_715);
xor U3806 (N_3806,In_21,In_889);
xor U3807 (N_3807,In_911,In_323);
or U3808 (N_3808,In_294,In_321);
xnor U3809 (N_3809,In_531,In_374);
nor U3810 (N_3810,In_104,In_8);
and U3811 (N_3811,In_171,In_996);
and U3812 (N_3812,In_476,In_497);
or U3813 (N_3813,In_708,In_491);
nor U3814 (N_3814,In_493,In_343);
and U3815 (N_3815,In_118,In_735);
or U3816 (N_3816,In_269,In_91);
nand U3817 (N_3817,In_699,In_418);
and U3818 (N_3818,In_869,In_511);
nand U3819 (N_3819,In_145,In_788);
nand U3820 (N_3820,In_855,In_222);
xnor U3821 (N_3821,In_467,In_438);
xor U3822 (N_3822,In_70,In_615);
and U3823 (N_3823,In_666,In_186);
nor U3824 (N_3824,In_730,In_559);
nor U3825 (N_3825,In_903,In_785);
xnor U3826 (N_3826,In_588,In_862);
or U3827 (N_3827,In_510,In_26);
nand U3828 (N_3828,In_869,In_851);
or U3829 (N_3829,In_439,In_810);
and U3830 (N_3830,In_599,In_881);
and U3831 (N_3831,In_288,In_404);
and U3832 (N_3832,In_268,In_850);
nand U3833 (N_3833,In_784,In_494);
nand U3834 (N_3834,In_390,In_852);
nand U3835 (N_3835,In_218,In_229);
nor U3836 (N_3836,In_693,In_23);
and U3837 (N_3837,In_635,In_538);
nand U3838 (N_3838,In_383,In_608);
and U3839 (N_3839,In_644,In_947);
or U3840 (N_3840,In_968,In_953);
nor U3841 (N_3841,In_925,In_460);
nand U3842 (N_3842,In_699,In_374);
and U3843 (N_3843,In_259,In_678);
nor U3844 (N_3844,In_353,In_29);
and U3845 (N_3845,In_765,In_871);
nor U3846 (N_3846,In_562,In_93);
and U3847 (N_3847,In_960,In_891);
and U3848 (N_3848,In_138,In_677);
nor U3849 (N_3849,In_836,In_126);
nand U3850 (N_3850,In_815,In_145);
or U3851 (N_3851,In_641,In_871);
xor U3852 (N_3852,In_604,In_898);
nor U3853 (N_3853,In_322,In_831);
or U3854 (N_3854,In_622,In_961);
nand U3855 (N_3855,In_466,In_244);
nor U3856 (N_3856,In_853,In_526);
or U3857 (N_3857,In_465,In_449);
nand U3858 (N_3858,In_423,In_494);
xor U3859 (N_3859,In_36,In_107);
nor U3860 (N_3860,In_709,In_666);
nor U3861 (N_3861,In_655,In_996);
and U3862 (N_3862,In_406,In_865);
nand U3863 (N_3863,In_993,In_933);
nor U3864 (N_3864,In_252,In_863);
or U3865 (N_3865,In_424,In_549);
and U3866 (N_3866,In_971,In_649);
and U3867 (N_3867,In_372,In_2);
xor U3868 (N_3868,In_165,In_814);
nor U3869 (N_3869,In_369,In_57);
and U3870 (N_3870,In_983,In_500);
nor U3871 (N_3871,In_184,In_906);
and U3872 (N_3872,In_78,In_586);
xnor U3873 (N_3873,In_137,In_647);
xor U3874 (N_3874,In_830,In_59);
or U3875 (N_3875,In_948,In_482);
and U3876 (N_3876,In_548,In_680);
nor U3877 (N_3877,In_223,In_658);
or U3878 (N_3878,In_6,In_769);
and U3879 (N_3879,In_376,In_930);
nand U3880 (N_3880,In_411,In_882);
nand U3881 (N_3881,In_612,In_507);
nor U3882 (N_3882,In_232,In_919);
and U3883 (N_3883,In_674,In_557);
and U3884 (N_3884,In_680,In_10);
nand U3885 (N_3885,In_812,In_141);
nor U3886 (N_3886,In_399,In_966);
or U3887 (N_3887,In_208,In_493);
and U3888 (N_3888,In_609,In_529);
nand U3889 (N_3889,In_507,In_275);
nor U3890 (N_3890,In_606,In_183);
nor U3891 (N_3891,In_993,In_511);
and U3892 (N_3892,In_830,In_322);
nand U3893 (N_3893,In_522,In_92);
and U3894 (N_3894,In_494,In_215);
or U3895 (N_3895,In_957,In_977);
nor U3896 (N_3896,In_560,In_713);
or U3897 (N_3897,In_58,In_908);
nor U3898 (N_3898,In_357,In_225);
nand U3899 (N_3899,In_684,In_457);
xor U3900 (N_3900,In_605,In_662);
nor U3901 (N_3901,In_62,In_470);
xnor U3902 (N_3902,In_699,In_608);
nand U3903 (N_3903,In_665,In_476);
or U3904 (N_3904,In_833,In_308);
or U3905 (N_3905,In_284,In_446);
xnor U3906 (N_3906,In_156,In_716);
and U3907 (N_3907,In_601,In_218);
and U3908 (N_3908,In_91,In_625);
nand U3909 (N_3909,In_121,In_822);
nand U3910 (N_3910,In_303,In_694);
nand U3911 (N_3911,In_777,In_526);
or U3912 (N_3912,In_223,In_661);
nor U3913 (N_3913,In_353,In_256);
or U3914 (N_3914,In_792,In_892);
nand U3915 (N_3915,In_154,In_505);
and U3916 (N_3916,In_267,In_760);
nand U3917 (N_3917,In_11,In_391);
or U3918 (N_3918,In_515,In_970);
or U3919 (N_3919,In_943,In_144);
nor U3920 (N_3920,In_219,In_468);
and U3921 (N_3921,In_125,In_249);
nand U3922 (N_3922,In_798,In_750);
or U3923 (N_3923,In_196,In_73);
nor U3924 (N_3924,In_505,In_662);
nor U3925 (N_3925,In_52,In_518);
and U3926 (N_3926,In_204,In_990);
and U3927 (N_3927,In_734,In_201);
or U3928 (N_3928,In_517,In_163);
nor U3929 (N_3929,In_855,In_882);
nor U3930 (N_3930,In_30,In_949);
or U3931 (N_3931,In_455,In_851);
and U3932 (N_3932,In_145,In_346);
nand U3933 (N_3933,In_442,In_798);
nand U3934 (N_3934,In_143,In_926);
and U3935 (N_3935,In_902,In_37);
nand U3936 (N_3936,In_940,In_897);
or U3937 (N_3937,In_587,In_788);
nor U3938 (N_3938,In_67,In_141);
nand U3939 (N_3939,In_812,In_831);
nor U3940 (N_3940,In_22,In_839);
xor U3941 (N_3941,In_38,In_55);
and U3942 (N_3942,In_485,In_629);
nand U3943 (N_3943,In_264,In_89);
or U3944 (N_3944,In_822,In_907);
or U3945 (N_3945,In_922,In_302);
xor U3946 (N_3946,In_98,In_532);
or U3947 (N_3947,In_330,In_708);
and U3948 (N_3948,In_368,In_81);
xnor U3949 (N_3949,In_539,In_971);
nor U3950 (N_3950,In_26,In_68);
and U3951 (N_3951,In_402,In_517);
or U3952 (N_3952,In_146,In_881);
or U3953 (N_3953,In_706,In_178);
nand U3954 (N_3954,In_844,In_584);
or U3955 (N_3955,In_855,In_553);
and U3956 (N_3956,In_666,In_94);
nor U3957 (N_3957,In_611,In_845);
xor U3958 (N_3958,In_748,In_936);
or U3959 (N_3959,In_542,In_378);
nor U3960 (N_3960,In_226,In_132);
or U3961 (N_3961,In_565,In_690);
nand U3962 (N_3962,In_913,In_1);
or U3963 (N_3963,In_838,In_944);
xnor U3964 (N_3964,In_81,In_845);
nand U3965 (N_3965,In_608,In_429);
nand U3966 (N_3966,In_922,In_42);
nor U3967 (N_3967,In_104,In_116);
nand U3968 (N_3968,In_386,In_276);
nand U3969 (N_3969,In_474,In_266);
xor U3970 (N_3970,In_773,In_21);
and U3971 (N_3971,In_103,In_173);
or U3972 (N_3972,In_781,In_620);
and U3973 (N_3973,In_205,In_730);
and U3974 (N_3974,In_181,In_384);
nand U3975 (N_3975,In_167,In_330);
nand U3976 (N_3976,In_470,In_147);
nand U3977 (N_3977,In_816,In_741);
or U3978 (N_3978,In_265,In_672);
nor U3979 (N_3979,In_724,In_874);
and U3980 (N_3980,In_92,In_322);
or U3981 (N_3981,In_945,In_142);
or U3982 (N_3982,In_953,In_655);
or U3983 (N_3983,In_615,In_365);
xnor U3984 (N_3984,In_744,In_742);
xnor U3985 (N_3985,In_352,In_821);
nor U3986 (N_3986,In_514,In_142);
and U3987 (N_3987,In_447,In_438);
or U3988 (N_3988,In_516,In_48);
nor U3989 (N_3989,In_685,In_388);
nand U3990 (N_3990,In_326,In_253);
nand U3991 (N_3991,In_61,In_911);
or U3992 (N_3992,In_329,In_404);
nor U3993 (N_3993,In_35,In_253);
or U3994 (N_3994,In_474,In_622);
nor U3995 (N_3995,In_607,In_330);
and U3996 (N_3996,In_487,In_869);
nor U3997 (N_3997,In_8,In_437);
or U3998 (N_3998,In_936,In_769);
nand U3999 (N_3999,In_866,In_976);
or U4000 (N_4000,In_722,In_975);
xnor U4001 (N_4001,In_505,In_50);
or U4002 (N_4002,In_181,In_955);
and U4003 (N_4003,In_189,In_645);
and U4004 (N_4004,In_7,In_649);
and U4005 (N_4005,In_155,In_915);
nor U4006 (N_4006,In_188,In_273);
xor U4007 (N_4007,In_946,In_718);
nand U4008 (N_4008,In_915,In_127);
and U4009 (N_4009,In_476,In_442);
xnor U4010 (N_4010,In_548,In_411);
nor U4011 (N_4011,In_90,In_145);
and U4012 (N_4012,In_756,In_881);
nor U4013 (N_4013,In_843,In_82);
nor U4014 (N_4014,In_701,In_433);
nor U4015 (N_4015,In_549,In_433);
nor U4016 (N_4016,In_952,In_725);
nor U4017 (N_4017,In_397,In_700);
nand U4018 (N_4018,In_465,In_549);
nor U4019 (N_4019,In_738,In_906);
nand U4020 (N_4020,In_771,In_268);
and U4021 (N_4021,In_694,In_332);
nor U4022 (N_4022,In_752,In_86);
nor U4023 (N_4023,In_54,In_552);
or U4024 (N_4024,In_525,In_447);
nand U4025 (N_4025,In_895,In_55);
nand U4026 (N_4026,In_640,In_633);
xor U4027 (N_4027,In_92,In_753);
or U4028 (N_4028,In_367,In_772);
xnor U4029 (N_4029,In_51,In_814);
nand U4030 (N_4030,In_269,In_762);
nor U4031 (N_4031,In_762,In_100);
and U4032 (N_4032,In_942,In_570);
nand U4033 (N_4033,In_694,In_563);
and U4034 (N_4034,In_730,In_258);
and U4035 (N_4035,In_452,In_332);
nand U4036 (N_4036,In_180,In_679);
or U4037 (N_4037,In_636,In_648);
nand U4038 (N_4038,In_848,In_882);
nand U4039 (N_4039,In_188,In_80);
or U4040 (N_4040,In_947,In_728);
nand U4041 (N_4041,In_824,In_579);
nor U4042 (N_4042,In_173,In_359);
nand U4043 (N_4043,In_500,In_170);
nand U4044 (N_4044,In_855,In_207);
or U4045 (N_4045,In_493,In_576);
and U4046 (N_4046,In_608,In_635);
nand U4047 (N_4047,In_268,In_311);
nor U4048 (N_4048,In_542,In_402);
or U4049 (N_4049,In_167,In_497);
and U4050 (N_4050,In_48,In_574);
or U4051 (N_4051,In_208,In_788);
nor U4052 (N_4052,In_109,In_424);
and U4053 (N_4053,In_523,In_884);
nor U4054 (N_4054,In_116,In_644);
or U4055 (N_4055,In_3,In_926);
or U4056 (N_4056,In_227,In_215);
nor U4057 (N_4057,In_237,In_117);
nand U4058 (N_4058,In_968,In_39);
and U4059 (N_4059,In_619,In_827);
and U4060 (N_4060,In_198,In_384);
or U4061 (N_4061,In_261,In_330);
nor U4062 (N_4062,In_326,In_804);
xnor U4063 (N_4063,In_291,In_46);
or U4064 (N_4064,In_752,In_612);
nand U4065 (N_4065,In_617,In_38);
nor U4066 (N_4066,In_595,In_985);
nand U4067 (N_4067,In_425,In_992);
xnor U4068 (N_4068,In_479,In_147);
and U4069 (N_4069,In_253,In_188);
or U4070 (N_4070,In_888,In_692);
or U4071 (N_4071,In_223,In_337);
or U4072 (N_4072,In_753,In_978);
nor U4073 (N_4073,In_398,In_832);
nor U4074 (N_4074,In_692,In_501);
xor U4075 (N_4075,In_557,In_216);
and U4076 (N_4076,In_345,In_862);
or U4077 (N_4077,In_134,In_497);
nand U4078 (N_4078,In_638,In_836);
nand U4079 (N_4079,In_430,In_841);
and U4080 (N_4080,In_392,In_342);
nor U4081 (N_4081,In_610,In_604);
or U4082 (N_4082,In_972,In_927);
or U4083 (N_4083,In_622,In_230);
and U4084 (N_4084,In_328,In_598);
nor U4085 (N_4085,In_694,In_981);
nand U4086 (N_4086,In_207,In_60);
and U4087 (N_4087,In_199,In_35);
nand U4088 (N_4088,In_378,In_662);
or U4089 (N_4089,In_322,In_367);
xor U4090 (N_4090,In_367,In_793);
or U4091 (N_4091,In_881,In_484);
nand U4092 (N_4092,In_230,In_255);
nand U4093 (N_4093,In_314,In_731);
nand U4094 (N_4094,In_478,In_95);
nor U4095 (N_4095,In_759,In_977);
or U4096 (N_4096,In_586,In_892);
and U4097 (N_4097,In_472,In_550);
nand U4098 (N_4098,In_338,In_109);
or U4099 (N_4099,In_834,In_964);
nand U4100 (N_4100,In_932,In_827);
xor U4101 (N_4101,In_222,In_593);
xor U4102 (N_4102,In_535,In_407);
nor U4103 (N_4103,In_156,In_981);
or U4104 (N_4104,In_546,In_74);
and U4105 (N_4105,In_89,In_904);
or U4106 (N_4106,In_411,In_860);
nor U4107 (N_4107,In_337,In_848);
or U4108 (N_4108,In_443,In_991);
xnor U4109 (N_4109,In_133,In_231);
nand U4110 (N_4110,In_973,In_377);
and U4111 (N_4111,In_326,In_333);
nand U4112 (N_4112,In_750,In_663);
and U4113 (N_4113,In_74,In_291);
nor U4114 (N_4114,In_512,In_439);
nand U4115 (N_4115,In_14,In_943);
and U4116 (N_4116,In_79,In_503);
nor U4117 (N_4117,In_158,In_119);
nor U4118 (N_4118,In_939,In_684);
or U4119 (N_4119,In_535,In_440);
or U4120 (N_4120,In_840,In_861);
or U4121 (N_4121,In_374,In_847);
nand U4122 (N_4122,In_924,In_8);
nand U4123 (N_4123,In_750,In_813);
and U4124 (N_4124,In_468,In_990);
nand U4125 (N_4125,In_707,In_229);
xor U4126 (N_4126,In_453,In_636);
and U4127 (N_4127,In_475,In_977);
and U4128 (N_4128,In_12,In_658);
nor U4129 (N_4129,In_790,In_338);
or U4130 (N_4130,In_175,In_519);
or U4131 (N_4131,In_91,In_63);
nand U4132 (N_4132,In_97,In_339);
nand U4133 (N_4133,In_993,In_308);
or U4134 (N_4134,In_350,In_20);
nor U4135 (N_4135,In_204,In_382);
nand U4136 (N_4136,In_897,In_327);
nor U4137 (N_4137,In_139,In_698);
nor U4138 (N_4138,In_937,In_394);
or U4139 (N_4139,In_585,In_274);
or U4140 (N_4140,In_311,In_426);
nand U4141 (N_4141,In_78,In_251);
and U4142 (N_4142,In_458,In_627);
or U4143 (N_4143,In_521,In_548);
nor U4144 (N_4144,In_809,In_69);
and U4145 (N_4145,In_117,In_54);
or U4146 (N_4146,In_500,In_657);
or U4147 (N_4147,In_234,In_418);
and U4148 (N_4148,In_393,In_450);
nor U4149 (N_4149,In_629,In_586);
nor U4150 (N_4150,In_600,In_940);
nand U4151 (N_4151,In_959,In_539);
nor U4152 (N_4152,In_466,In_815);
or U4153 (N_4153,In_143,In_715);
or U4154 (N_4154,In_93,In_203);
nand U4155 (N_4155,In_822,In_444);
xor U4156 (N_4156,In_916,In_910);
nor U4157 (N_4157,In_960,In_193);
xnor U4158 (N_4158,In_241,In_151);
or U4159 (N_4159,In_707,In_638);
nand U4160 (N_4160,In_733,In_147);
nand U4161 (N_4161,In_772,In_126);
or U4162 (N_4162,In_167,In_822);
nor U4163 (N_4163,In_570,In_319);
or U4164 (N_4164,In_469,In_641);
xnor U4165 (N_4165,In_49,In_96);
and U4166 (N_4166,In_615,In_958);
nor U4167 (N_4167,In_76,In_802);
and U4168 (N_4168,In_876,In_375);
nand U4169 (N_4169,In_929,In_472);
or U4170 (N_4170,In_326,In_730);
xor U4171 (N_4171,In_422,In_525);
and U4172 (N_4172,In_300,In_658);
or U4173 (N_4173,In_120,In_96);
or U4174 (N_4174,In_586,In_232);
nand U4175 (N_4175,In_609,In_39);
nand U4176 (N_4176,In_730,In_905);
nor U4177 (N_4177,In_897,In_760);
or U4178 (N_4178,In_238,In_365);
nor U4179 (N_4179,In_734,In_577);
nand U4180 (N_4180,In_356,In_958);
xnor U4181 (N_4181,In_327,In_87);
nand U4182 (N_4182,In_636,In_28);
nor U4183 (N_4183,In_784,In_937);
or U4184 (N_4184,In_522,In_354);
nor U4185 (N_4185,In_306,In_573);
nor U4186 (N_4186,In_552,In_350);
xnor U4187 (N_4187,In_25,In_58);
or U4188 (N_4188,In_627,In_230);
nand U4189 (N_4189,In_18,In_155);
xor U4190 (N_4190,In_627,In_892);
nand U4191 (N_4191,In_381,In_329);
nor U4192 (N_4192,In_575,In_484);
nor U4193 (N_4193,In_855,In_237);
nor U4194 (N_4194,In_943,In_363);
nor U4195 (N_4195,In_541,In_320);
xnor U4196 (N_4196,In_805,In_102);
or U4197 (N_4197,In_483,In_913);
xnor U4198 (N_4198,In_570,In_873);
or U4199 (N_4199,In_866,In_503);
nand U4200 (N_4200,In_711,In_561);
xnor U4201 (N_4201,In_524,In_604);
and U4202 (N_4202,In_96,In_217);
nand U4203 (N_4203,In_578,In_572);
nor U4204 (N_4204,In_28,In_683);
nor U4205 (N_4205,In_162,In_658);
xnor U4206 (N_4206,In_497,In_435);
nor U4207 (N_4207,In_889,In_405);
or U4208 (N_4208,In_14,In_599);
xor U4209 (N_4209,In_398,In_682);
or U4210 (N_4210,In_947,In_693);
nand U4211 (N_4211,In_493,In_957);
nor U4212 (N_4212,In_208,In_784);
nand U4213 (N_4213,In_118,In_656);
nor U4214 (N_4214,In_837,In_580);
nor U4215 (N_4215,In_219,In_33);
nand U4216 (N_4216,In_731,In_927);
and U4217 (N_4217,In_154,In_269);
xnor U4218 (N_4218,In_772,In_193);
xnor U4219 (N_4219,In_475,In_198);
xor U4220 (N_4220,In_720,In_991);
nor U4221 (N_4221,In_596,In_953);
xor U4222 (N_4222,In_888,In_810);
or U4223 (N_4223,In_27,In_153);
and U4224 (N_4224,In_456,In_30);
nor U4225 (N_4225,In_492,In_6);
nand U4226 (N_4226,In_869,In_275);
and U4227 (N_4227,In_337,In_185);
nand U4228 (N_4228,In_4,In_993);
nand U4229 (N_4229,In_778,In_662);
nand U4230 (N_4230,In_805,In_232);
or U4231 (N_4231,In_700,In_716);
or U4232 (N_4232,In_320,In_452);
nor U4233 (N_4233,In_524,In_172);
and U4234 (N_4234,In_516,In_600);
nor U4235 (N_4235,In_902,In_767);
and U4236 (N_4236,In_569,In_361);
nor U4237 (N_4237,In_519,In_336);
or U4238 (N_4238,In_540,In_873);
or U4239 (N_4239,In_584,In_266);
or U4240 (N_4240,In_770,In_956);
or U4241 (N_4241,In_939,In_918);
or U4242 (N_4242,In_532,In_239);
nor U4243 (N_4243,In_600,In_738);
nand U4244 (N_4244,In_178,In_442);
nand U4245 (N_4245,In_643,In_833);
nand U4246 (N_4246,In_242,In_838);
nand U4247 (N_4247,In_765,In_739);
nand U4248 (N_4248,In_410,In_989);
or U4249 (N_4249,In_365,In_7);
xor U4250 (N_4250,In_215,In_72);
nor U4251 (N_4251,In_418,In_475);
nand U4252 (N_4252,In_198,In_147);
or U4253 (N_4253,In_726,In_565);
or U4254 (N_4254,In_864,In_217);
or U4255 (N_4255,In_979,In_233);
nor U4256 (N_4256,In_10,In_26);
xor U4257 (N_4257,In_745,In_59);
and U4258 (N_4258,In_567,In_294);
or U4259 (N_4259,In_122,In_669);
or U4260 (N_4260,In_452,In_877);
nand U4261 (N_4261,In_655,In_467);
nor U4262 (N_4262,In_950,In_956);
nand U4263 (N_4263,In_782,In_400);
nor U4264 (N_4264,In_231,In_733);
and U4265 (N_4265,In_392,In_924);
and U4266 (N_4266,In_717,In_733);
nor U4267 (N_4267,In_407,In_504);
nand U4268 (N_4268,In_388,In_637);
nand U4269 (N_4269,In_715,In_117);
or U4270 (N_4270,In_131,In_576);
or U4271 (N_4271,In_2,In_210);
nor U4272 (N_4272,In_112,In_122);
xnor U4273 (N_4273,In_778,In_413);
nor U4274 (N_4274,In_583,In_730);
or U4275 (N_4275,In_836,In_336);
and U4276 (N_4276,In_488,In_844);
nand U4277 (N_4277,In_822,In_626);
nand U4278 (N_4278,In_284,In_740);
nand U4279 (N_4279,In_170,In_703);
nor U4280 (N_4280,In_699,In_937);
nor U4281 (N_4281,In_873,In_227);
and U4282 (N_4282,In_726,In_245);
nor U4283 (N_4283,In_111,In_376);
or U4284 (N_4284,In_52,In_381);
nor U4285 (N_4285,In_416,In_916);
nand U4286 (N_4286,In_621,In_676);
nand U4287 (N_4287,In_660,In_799);
or U4288 (N_4288,In_849,In_167);
nand U4289 (N_4289,In_133,In_434);
xor U4290 (N_4290,In_493,In_19);
and U4291 (N_4291,In_133,In_504);
and U4292 (N_4292,In_144,In_950);
nand U4293 (N_4293,In_198,In_681);
or U4294 (N_4294,In_386,In_792);
nor U4295 (N_4295,In_440,In_377);
nor U4296 (N_4296,In_294,In_589);
nor U4297 (N_4297,In_345,In_497);
nand U4298 (N_4298,In_501,In_235);
xor U4299 (N_4299,In_664,In_940);
and U4300 (N_4300,In_829,In_78);
and U4301 (N_4301,In_423,In_737);
nor U4302 (N_4302,In_285,In_89);
nor U4303 (N_4303,In_88,In_250);
or U4304 (N_4304,In_145,In_594);
or U4305 (N_4305,In_308,In_928);
nand U4306 (N_4306,In_248,In_431);
nand U4307 (N_4307,In_555,In_621);
nor U4308 (N_4308,In_872,In_131);
nor U4309 (N_4309,In_657,In_990);
xor U4310 (N_4310,In_987,In_571);
nand U4311 (N_4311,In_346,In_384);
and U4312 (N_4312,In_169,In_188);
or U4313 (N_4313,In_492,In_405);
and U4314 (N_4314,In_906,In_904);
nand U4315 (N_4315,In_955,In_133);
nand U4316 (N_4316,In_269,In_732);
nand U4317 (N_4317,In_497,In_188);
nor U4318 (N_4318,In_502,In_672);
or U4319 (N_4319,In_187,In_198);
nand U4320 (N_4320,In_134,In_322);
or U4321 (N_4321,In_189,In_86);
and U4322 (N_4322,In_547,In_958);
nand U4323 (N_4323,In_48,In_584);
nand U4324 (N_4324,In_862,In_366);
nand U4325 (N_4325,In_471,In_928);
or U4326 (N_4326,In_643,In_946);
or U4327 (N_4327,In_466,In_498);
and U4328 (N_4328,In_147,In_454);
nor U4329 (N_4329,In_212,In_532);
or U4330 (N_4330,In_723,In_663);
nor U4331 (N_4331,In_176,In_848);
or U4332 (N_4332,In_180,In_496);
nand U4333 (N_4333,In_275,In_901);
or U4334 (N_4334,In_277,In_916);
or U4335 (N_4335,In_202,In_648);
xnor U4336 (N_4336,In_379,In_30);
nor U4337 (N_4337,In_153,In_924);
and U4338 (N_4338,In_761,In_185);
nand U4339 (N_4339,In_633,In_39);
and U4340 (N_4340,In_530,In_503);
xnor U4341 (N_4341,In_95,In_595);
or U4342 (N_4342,In_659,In_6);
and U4343 (N_4343,In_191,In_204);
or U4344 (N_4344,In_668,In_693);
nor U4345 (N_4345,In_77,In_681);
and U4346 (N_4346,In_151,In_236);
xor U4347 (N_4347,In_341,In_920);
nand U4348 (N_4348,In_445,In_530);
nor U4349 (N_4349,In_344,In_620);
and U4350 (N_4350,In_796,In_559);
or U4351 (N_4351,In_911,In_89);
or U4352 (N_4352,In_723,In_750);
and U4353 (N_4353,In_971,In_465);
xor U4354 (N_4354,In_540,In_575);
or U4355 (N_4355,In_7,In_691);
nand U4356 (N_4356,In_948,In_524);
and U4357 (N_4357,In_400,In_790);
and U4358 (N_4358,In_23,In_20);
or U4359 (N_4359,In_699,In_763);
and U4360 (N_4360,In_547,In_620);
or U4361 (N_4361,In_995,In_586);
xnor U4362 (N_4362,In_443,In_667);
or U4363 (N_4363,In_846,In_426);
or U4364 (N_4364,In_153,In_728);
and U4365 (N_4365,In_194,In_885);
or U4366 (N_4366,In_465,In_374);
nand U4367 (N_4367,In_41,In_107);
xnor U4368 (N_4368,In_803,In_410);
nand U4369 (N_4369,In_97,In_723);
or U4370 (N_4370,In_820,In_713);
nor U4371 (N_4371,In_154,In_740);
or U4372 (N_4372,In_352,In_368);
or U4373 (N_4373,In_205,In_225);
or U4374 (N_4374,In_129,In_930);
or U4375 (N_4375,In_374,In_554);
nor U4376 (N_4376,In_111,In_523);
or U4377 (N_4377,In_158,In_797);
or U4378 (N_4378,In_298,In_180);
and U4379 (N_4379,In_879,In_951);
nor U4380 (N_4380,In_900,In_777);
nand U4381 (N_4381,In_113,In_195);
or U4382 (N_4382,In_162,In_220);
or U4383 (N_4383,In_469,In_986);
nand U4384 (N_4384,In_445,In_24);
or U4385 (N_4385,In_584,In_862);
nor U4386 (N_4386,In_410,In_374);
and U4387 (N_4387,In_984,In_679);
nand U4388 (N_4388,In_148,In_505);
or U4389 (N_4389,In_211,In_711);
and U4390 (N_4390,In_360,In_845);
or U4391 (N_4391,In_547,In_331);
nor U4392 (N_4392,In_233,In_141);
nand U4393 (N_4393,In_80,In_601);
nand U4394 (N_4394,In_297,In_119);
and U4395 (N_4395,In_641,In_840);
nor U4396 (N_4396,In_937,In_660);
or U4397 (N_4397,In_442,In_777);
and U4398 (N_4398,In_315,In_758);
nand U4399 (N_4399,In_519,In_890);
xnor U4400 (N_4400,In_283,In_243);
or U4401 (N_4401,In_439,In_832);
or U4402 (N_4402,In_235,In_213);
nor U4403 (N_4403,In_117,In_735);
xor U4404 (N_4404,In_730,In_374);
or U4405 (N_4405,In_727,In_813);
nor U4406 (N_4406,In_932,In_940);
and U4407 (N_4407,In_355,In_0);
and U4408 (N_4408,In_403,In_177);
or U4409 (N_4409,In_485,In_347);
or U4410 (N_4410,In_872,In_788);
nor U4411 (N_4411,In_17,In_371);
nand U4412 (N_4412,In_73,In_350);
or U4413 (N_4413,In_860,In_521);
nand U4414 (N_4414,In_890,In_393);
nor U4415 (N_4415,In_439,In_989);
nand U4416 (N_4416,In_176,In_27);
and U4417 (N_4417,In_704,In_623);
nor U4418 (N_4418,In_105,In_407);
and U4419 (N_4419,In_138,In_830);
nor U4420 (N_4420,In_486,In_493);
and U4421 (N_4421,In_777,In_18);
nand U4422 (N_4422,In_842,In_549);
xnor U4423 (N_4423,In_943,In_769);
and U4424 (N_4424,In_75,In_786);
nand U4425 (N_4425,In_665,In_921);
and U4426 (N_4426,In_623,In_193);
and U4427 (N_4427,In_339,In_370);
nand U4428 (N_4428,In_770,In_448);
xor U4429 (N_4429,In_707,In_517);
nor U4430 (N_4430,In_213,In_948);
or U4431 (N_4431,In_128,In_908);
nand U4432 (N_4432,In_138,In_34);
and U4433 (N_4433,In_775,In_352);
nand U4434 (N_4434,In_48,In_6);
or U4435 (N_4435,In_851,In_113);
nand U4436 (N_4436,In_951,In_449);
or U4437 (N_4437,In_844,In_926);
nor U4438 (N_4438,In_911,In_225);
or U4439 (N_4439,In_131,In_541);
nor U4440 (N_4440,In_793,In_35);
nand U4441 (N_4441,In_470,In_127);
nand U4442 (N_4442,In_669,In_408);
nand U4443 (N_4443,In_46,In_592);
nand U4444 (N_4444,In_524,In_970);
nand U4445 (N_4445,In_321,In_244);
nor U4446 (N_4446,In_221,In_706);
nor U4447 (N_4447,In_917,In_95);
or U4448 (N_4448,In_365,In_283);
nor U4449 (N_4449,In_679,In_788);
and U4450 (N_4450,In_127,In_37);
nand U4451 (N_4451,In_141,In_667);
nand U4452 (N_4452,In_854,In_238);
nand U4453 (N_4453,In_547,In_121);
or U4454 (N_4454,In_109,In_77);
or U4455 (N_4455,In_548,In_90);
nor U4456 (N_4456,In_381,In_206);
and U4457 (N_4457,In_827,In_468);
xor U4458 (N_4458,In_397,In_66);
nand U4459 (N_4459,In_515,In_194);
and U4460 (N_4460,In_137,In_391);
nor U4461 (N_4461,In_825,In_244);
or U4462 (N_4462,In_55,In_617);
nor U4463 (N_4463,In_908,In_56);
nor U4464 (N_4464,In_94,In_26);
nand U4465 (N_4465,In_172,In_816);
nor U4466 (N_4466,In_292,In_277);
nor U4467 (N_4467,In_868,In_63);
or U4468 (N_4468,In_278,In_933);
and U4469 (N_4469,In_733,In_678);
nand U4470 (N_4470,In_863,In_30);
and U4471 (N_4471,In_297,In_404);
or U4472 (N_4472,In_338,In_32);
or U4473 (N_4473,In_299,In_999);
and U4474 (N_4474,In_468,In_563);
xor U4475 (N_4475,In_42,In_99);
nor U4476 (N_4476,In_464,In_896);
and U4477 (N_4477,In_305,In_511);
xnor U4478 (N_4478,In_778,In_85);
and U4479 (N_4479,In_866,In_354);
xor U4480 (N_4480,In_758,In_281);
nor U4481 (N_4481,In_400,In_541);
nor U4482 (N_4482,In_996,In_480);
nand U4483 (N_4483,In_192,In_842);
and U4484 (N_4484,In_200,In_119);
xnor U4485 (N_4485,In_537,In_866);
and U4486 (N_4486,In_53,In_291);
nand U4487 (N_4487,In_254,In_85);
or U4488 (N_4488,In_751,In_216);
nand U4489 (N_4489,In_341,In_811);
nand U4490 (N_4490,In_119,In_95);
xor U4491 (N_4491,In_125,In_870);
or U4492 (N_4492,In_93,In_861);
nor U4493 (N_4493,In_29,In_306);
or U4494 (N_4494,In_256,In_191);
nor U4495 (N_4495,In_965,In_237);
and U4496 (N_4496,In_834,In_147);
or U4497 (N_4497,In_414,In_998);
nand U4498 (N_4498,In_649,In_846);
or U4499 (N_4499,In_238,In_408);
xor U4500 (N_4500,In_692,In_67);
or U4501 (N_4501,In_494,In_613);
nand U4502 (N_4502,In_644,In_238);
and U4503 (N_4503,In_525,In_491);
and U4504 (N_4504,In_972,In_603);
or U4505 (N_4505,In_658,In_936);
xnor U4506 (N_4506,In_813,In_884);
nor U4507 (N_4507,In_710,In_384);
nand U4508 (N_4508,In_595,In_25);
nor U4509 (N_4509,In_698,In_747);
nor U4510 (N_4510,In_519,In_235);
or U4511 (N_4511,In_900,In_25);
or U4512 (N_4512,In_469,In_320);
nor U4513 (N_4513,In_833,In_658);
nor U4514 (N_4514,In_502,In_430);
and U4515 (N_4515,In_24,In_350);
xor U4516 (N_4516,In_867,In_420);
and U4517 (N_4517,In_104,In_481);
nor U4518 (N_4518,In_966,In_702);
nor U4519 (N_4519,In_215,In_462);
nor U4520 (N_4520,In_891,In_189);
or U4521 (N_4521,In_848,In_5);
or U4522 (N_4522,In_149,In_115);
and U4523 (N_4523,In_279,In_116);
and U4524 (N_4524,In_604,In_111);
xor U4525 (N_4525,In_954,In_977);
and U4526 (N_4526,In_353,In_548);
xnor U4527 (N_4527,In_347,In_214);
or U4528 (N_4528,In_727,In_256);
nor U4529 (N_4529,In_862,In_888);
nand U4530 (N_4530,In_486,In_633);
nor U4531 (N_4531,In_901,In_876);
nand U4532 (N_4532,In_110,In_811);
or U4533 (N_4533,In_494,In_953);
nor U4534 (N_4534,In_869,In_839);
nor U4535 (N_4535,In_737,In_783);
or U4536 (N_4536,In_542,In_846);
nor U4537 (N_4537,In_221,In_713);
nand U4538 (N_4538,In_279,In_922);
or U4539 (N_4539,In_558,In_598);
xnor U4540 (N_4540,In_636,In_345);
nand U4541 (N_4541,In_930,In_746);
and U4542 (N_4542,In_638,In_441);
nor U4543 (N_4543,In_918,In_608);
or U4544 (N_4544,In_409,In_0);
nand U4545 (N_4545,In_436,In_701);
or U4546 (N_4546,In_472,In_18);
and U4547 (N_4547,In_954,In_334);
nor U4548 (N_4548,In_196,In_43);
or U4549 (N_4549,In_432,In_65);
and U4550 (N_4550,In_808,In_581);
xor U4551 (N_4551,In_998,In_177);
or U4552 (N_4552,In_827,In_454);
and U4553 (N_4553,In_556,In_976);
and U4554 (N_4554,In_702,In_682);
nor U4555 (N_4555,In_390,In_291);
nand U4556 (N_4556,In_695,In_364);
and U4557 (N_4557,In_790,In_585);
and U4558 (N_4558,In_304,In_375);
nand U4559 (N_4559,In_70,In_497);
nand U4560 (N_4560,In_568,In_532);
or U4561 (N_4561,In_652,In_932);
nor U4562 (N_4562,In_370,In_633);
nor U4563 (N_4563,In_765,In_371);
nand U4564 (N_4564,In_612,In_965);
nor U4565 (N_4565,In_807,In_68);
and U4566 (N_4566,In_579,In_848);
and U4567 (N_4567,In_608,In_215);
nand U4568 (N_4568,In_293,In_54);
or U4569 (N_4569,In_102,In_511);
and U4570 (N_4570,In_149,In_649);
nand U4571 (N_4571,In_151,In_208);
or U4572 (N_4572,In_225,In_64);
xor U4573 (N_4573,In_657,In_537);
nand U4574 (N_4574,In_435,In_532);
nand U4575 (N_4575,In_445,In_772);
nor U4576 (N_4576,In_777,In_778);
and U4577 (N_4577,In_891,In_204);
nor U4578 (N_4578,In_236,In_346);
nor U4579 (N_4579,In_797,In_529);
or U4580 (N_4580,In_232,In_341);
and U4581 (N_4581,In_384,In_641);
nand U4582 (N_4582,In_159,In_742);
nand U4583 (N_4583,In_480,In_826);
and U4584 (N_4584,In_297,In_676);
or U4585 (N_4585,In_489,In_820);
nor U4586 (N_4586,In_492,In_760);
nor U4587 (N_4587,In_82,In_727);
and U4588 (N_4588,In_457,In_12);
and U4589 (N_4589,In_744,In_655);
or U4590 (N_4590,In_313,In_111);
nand U4591 (N_4591,In_520,In_881);
nand U4592 (N_4592,In_769,In_520);
or U4593 (N_4593,In_681,In_996);
or U4594 (N_4594,In_717,In_852);
and U4595 (N_4595,In_185,In_221);
or U4596 (N_4596,In_119,In_504);
and U4597 (N_4597,In_132,In_726);
nand U4598 (N_4598,In_984,In_868);
and U4599 (N_4599,In_669,In_582);
nand U4600 (N_4600,In_676,In_249);
nand U4601 (N_4601,In_501,In_668);
nor U4602 (N_4602,In_675,In_597);
or U4603 (N_4603,In_308,In_127);
xor U4604 (N_4604,In_456,In_264);
nor U4605 (N_4605,In_883,In_54);
or U4606 (N_4606,In_310,In_35);
nor U4607 (N_4607,In_110,In_946);
or U4608 (N_4608,In_343,In_390);
or U4609 (N_4609,In_139,In_590);
nor U4610 (N_4610,In_16,In_563);
nand U4611 (N_4611,In_554,In_457);
nor U4612 (N_4612,In_387,In_163);
and U4613 (N_4613,In_261,In_854);
or U4614 (N_4614,In_656,In_78);
and U4615 (N_4615,In_415,In_587);
xor U4616 (N_4616,In_610,In_809);
xor U4617 (N_4617,In_157,In_467);
or U4618 (N_4618,In_580,In_723);
nor U4619 (N_4619,In_699,In_170);
or U4620 (N_4620,In_442,In_160);
xor U4621 (N_4621,In_289,In_56);
nand U4622 (N_4622,In_997,In_563);
nand U4623 (N_4623,In_124,In_821);
nor U4624 (N_4624,In_361,In_250);
nor U4625 (N_4625,In_780,In_182);
nor U4626 (N_4626,In_409,In_767);
nor U4627 (N_4627,In_703,In_543);
nor U4628 (N_4628,In_490,In_194);
or U4629 (N_4629,In_408,In_907);
and U4630 (N_4630,In_108,In_84);
or U4631 (N_4631,In_914,In_928);
or U4632 (N_4632,In_541,In_971);
and U4633 (N_4633,In_493,In_566);
or U4634 (N_4634,In_250,In_464);
and U4635 (N_4635,In_769,In_242);
nor U4636 (N_4636,In_194,In_357);
or U4637 (N_4637,In_772,In_700);
and U4638 (N_4638,In_319,In_181);
and U4639 (N_4639,In_632,In_537);
or U4640 (N_4640,In_860,In_136);
or U4641 (N_4641,In_640,In_31);
nand U4642 (N_4642,In_838,In_409);
nor U4643 (N_4643,In_86,In_587);
or U4644 (N_4644,In_451,In_388);
nor U4645 (N_4645,In_980,In_881);
and U4646 (N_4646,In_499,In_572);
xnor U4647 (N_4647,In_711,In_188);
nand U4648 (N_4648,In_454,In_589);
or U4649 (N_4649,In_833,In_238);
and U4650 (N_4650,In_395,In_232);
nor U4651 (N_4651,In_364,In_71);
nand U4652 (N_4652,In_915,In_725);
or U4653 (N_4653,In_810,In_30);
and U4654 (N_4654,In_524,In_781);
xor U4655 (N_4655,In_659,In_833);
and U4656 (N_4656,In_607,In_334);
nor U4657 (N_4657,In_467,In_24);
nand U4658 (N_4658,In_742,In_428);
or U4659 (N_4659,In_810,In_234);
and U4660 (N_4660,In_646,In_957);
nor U4661 (N_4661,In_769,In_895);
or U4662 (N_4662,In_761,In_78);
nor U4663 (N_4663,In_517,In_880);
nand U4664 (N_4664,In_953,In_479);
or U4665 (N_4665,In_847,In_181);
nor U4666 (N_4666,In_215,In_968);
nor U4667 (N_4667,In_332,In_55);
xnor U4668 (N_4668,In_484,In_874);
or U4669 (N_4669,In_919,In_332);
or U4670 (N_4670,In_503,In_46);
nor U4671 (N_4671,In_985,In_31);
nand U4672 (N_4672,In_183,In_669);
or U4673 (N_4673,In_606,In_723);
nor U4674 (N_4674,In_168,In_535);
nor U4675 (N_4675,In_676,In_235);
and U4676 (N_4676,In_954,In_103);
or U4677 (N_4677,In_895,In_879);
nor U4678 (N_4678,In_470,In_598);
nand U4679 (N_4679,In_681,In_472);
nand U4680 (N_4680,In_868,In_2);
xor U4681 (N_4681,In_372,In_489);
nor U4682 (N_4682,In_358,In_459);
and U4683 (N_4683,In_28,In_679);
nand U4684 (N_4684,In_763,In_525);
and U4685 (N_4685,In_438,In_915);
and U4686 (N_4686,In_297,In_755);
nand U4687 (N_4687,In_892,In_490);
nand U4688 (N_4688,In_488,In_406);
nor U4689 (N_4689,In_611,In_882);
or U4690 (N_4690,In_237,In_221);
nand U4691 (N_4691,In_872,In_950);
xor U4692 (N_4692,In_685,In_422);
xor U4693 (N_4693,In_428,In_692);
or U4694 (N_4694,In_344,In_317);
nor U4695 (N_4695,In_677,In_811);
nor U4696 (N_4696,In_618,In_852);
or U4697 (N_4697,In_753,In_943);
and U4698 (N_4698,In_282,In_937);
or U4699 (N_4699,In_579,In_958);
or U4700 (N_4700,In_843,In_386);
nand U4701 (N_4701,In_127,In_630);
xnor U4702 (N_4702,In_936,In_541);
nor U4703 (N_4703,In_387,In_465);
and U4704 (N_4704,In_652,In_319);
and U4705 (N_4705,In_89,In_547);
nand U4706 (N_4706,In_780,In_848);
nor U4707 (N_4707,In_603,In_478);
xnor U4708 (N_4708,In_200,In_384);
and U4709 (N_4709,In_447,In_627);
nand U4710 (N_4710,In_185,In_431);
nand U4711 (N_4711,In_253,In_70);
nor U4712 (N_4712,In_208,In_700);
and U4713 (N_4713,In_968,In_250);
and U4714 (N_4714,In_943,In_513);
or U4715 (N_4715,In_441,In_473);
or U4716 (N_4716,In_317,In_721);
or U4717 (N_4717,In_336,In_825);
nand U4718 (N_4718,In_310,In_159);
nor U4719 (N_4719,In_984,In_779);
and U4720 (N_4720,In_430,In_56);
nand U4721 (N_4721,In_924,In_502);
or U4722 (N_4722,In_24,In_979);
nor U4723 (N_4723,In_327,In_984);
nand U4724 (N_4724,In_581,In_408);
or U4725 (N_4725,In_393,In_116);
nor U4726 (N_4726,In_831,In_612);
nand U4727 (N_4727,In_663,In_681);
or U4728 (N_4728,In_152,In_174);
nor U4729 (N_4729,In_320,In_326);
nor U4730 (N_4730,In_887,In_262);
nor U4731 (N_4731,In_348,In_589);
xor U4732 (N_4732,In_621,In_467);
nand U4733 (N_4733,In_963,In_476);
nand U4734 (N_4734,In_715,In_435);
and U4735 (N_4735,In_874,In_726);
nor U4736 (N_4736,In_972,In_14);
nand U4737 (N_4737,In_645,In_193);
nand U4738 (N_4738,In_634,In_766);
and U4739 (N_4739,In_594,In_462);
or U4740 (N_4740,In_663,In_956);
or U4741 (N_4741,In_761,In_232);
and U4742 (N_4742,In_312,In_906);
and U4743 (N_4743,In_822,In_414);
nor U4744 (N_4744,In_80,In_765);
nor U4745 (N_4745,In_185,In_908);
and U4746 (N_4746,In_69,In_668);
and U4747 (N_4747,In_575,In_21);
xor U4748 (N_4748,In_93,In_662);
or U4749 (N_4749,In_68,In_454);
or U4750 (N_4750,In_746,In_387);
nand U4751 (N_4751,In_351,In_458);
nor U4752 (N_4752,In_151,In_964);
nand U4753 (N_4753,In_122,In_67);
nor U4754 (N_4754,In_893,In_939);
nand U4755 (N_4755,In_557,In_205);
nand U4756 (N_4756,In_673,In_574);
xor U4757 (N_4757,In_450,In_847);
or U4758 (N_4758,In_930,In_295);
nor U4759 (N_4759,In_21,In_904);
xor U4760 (N_4760,In_644,In_94);
xnor U4761 (N_4761,In_687,In_96);
nand U4762 (N_4762,In_587,In_939);
nor U4763 (N_4763,In_249,In_648);
nor U4764 (N_4764,In_942,In_266);
or U4765 (N_4765,In_186,In_446);
nor U4766 (N_4766,In_545,In_646);
nor U4767 (N_4767,In_346,In_1);
and U4768 (N_4768,In_786,In_708);
or U4769 (N_4769,In_810,In_375);
nor U4770 (N_4770,In_628,In_118);
or U4771 (N_4771,In_179,In_919);
nand U4772 (N_4772,In_705,In_416);
and U4773 (N_4773,In_489,In_9);
or U4774 (N_4774,In_987,In_165);
or U4775 (N_4775,In_516,In_802);
xor U4776 (N_4776,In_308,In_784);
or U4777 (N_4777,In_140,In_937);
nand U4778 (N_4778,In_857,In_740);
nand U4779 (N_4779,In_358,In_514);
and U4780 (N_4780,In_259,In_403);
nand U4781 (N_4781,In_634,In_574);
xor U4782 (N_4782,In_91,In_917);
nand U4783 (N_4783,In_587,In_930);
nand U4784 (N_4784,In_998,In_8);
xor U4785 (N_4785,In_948,In_638);
nor U4786 (N_4786,In_604,In_333);
nand U4787 (N_4787,In_239,In_963);
or U4788 (N_4788,In_539,In_814);
xor U4789 (N_4789,In_744,In_229);
and U4790 (N_4790,In_203,In_112);
or U4791 (N_4791,In_556,In_495);
nor U4792 (N_4792,In_499,In_544);
nor U4793 (N_4793,In_356,In_526);
xnor U4794 (N_4794,In_418,In_99);
nand U4795 (N_4795,In_434,In_93);
xor U4796 (N_4796,In_740,In_391);
nor U4797 (N_4797,In_296,In_426);
and U4798 (N_4798,In_25,In_125);
nor U4799 (N_4799,In_106,In_927);
nand U4800 (N_4800,In_226,In_555);
or U4801 (N_4801,In_375,In_546);
nand U4802 (N_4802,In_779,In_656);
nor U4803 (N_4803,In_967,In_114);
and U4804 (N_4804,In_918,In_157);
nand U4805 (N_4805,In_616,In_498);
nand U4806 (N_4806,In_384,In_14);
nand U4807 (N_4807,In_278,In_647);
or U4808 (N_4808,In_147,In_725);
nand U4809 (N_4809,In_862,In_601);
xnor U4810 (N_4810,In_937,In_634);
and U4811 (N_4811,In_953,In_365);
and U4812 (N_4812,In_449,In_442);
or U4813 (N_4813,In_79,In_75);
nor U4814 (N_4814,In_807,In_958);
nand U4815 (N_4815,In_651,In_982);
nand U4816 (N_4816,In_583,In_279);
nand U4817 (N_4817,In_75,In_849);
nand U4818 (N_4818,In_819,In_670);
nand U4819 (N_4819,In_326,In_6);
or U4820 (N_4820,In_67,In_612);
and U4821 (N_4821,In_330,In_605);
and U4822 (N_4822,In_494,In_822);
nor U4823 (N_4823,In_43,In_357);
nor U4824 (N_4824,In_201,In_129);
and U4825 (N_4825,In_823,In_400);
and U4826 (N_4826,In_328,In_725);
nor U4827 (N_4827,In_851,In_177);
and U4828 (N_4828,In_208,In_578);
nor U4829 (N_4829,In_386,In_94);
and U4830 (N_4830,In_200,In_56);
nor U4831 (N_4831,In_439,In_441);
and U4832 (N_4832,In_415,In_250);
and U4833 (N_4833,In_238,In_400);
or U4834 (N_4834,In_204,In_35);
and U4835 (N_4835,In_26,In_531);
or U4836 (N_4836,In_671,In_492);
or U4837 (N_4837,In_502,In_821);
or U4838 (N_4838,In_741,In_486);
and U4839 (N_4839,In_432,In_143);
nand U4840 (N_4840,In_365,In_539);
and U4841 (N_4841,In_28,In_690);
xor U4842 (N_4842,In_95,In_132);
or U4843 (N_4843,In_949,In_138);
xor U4844 (N_4844,In_637,In_421);
and U4845 (N_4845,In_925,In_907);
xor U4846 (N_4846,In_351,In_875);
nand U4847 (N_4847,In_274,In_733);
nor U4848 (N_4848,In_254,In_555);
or U4849 (N_4849,In_461,In_634);
or U4850 (N_4850,In_384,In_357);
nand U4851 (N_4851,In_205,In_851);
or U4852 (N_4852,In_329,In_382);
and U4853 (N_4853,In_60,In_97);
nand U4854 (N_4854,In_199,In_357);
nand U4855 (N_4855,In_5,In_236);
nor U4856 (N_4856,In_603,In_487);
or U4857 (N_4857,In_367,In_774);
nor U4858 (N_4858,In_359,In_491);
or U4859 (N_4859,In_310,In_259);
nand U4860 (N_4860,In_993,In_206);
or U4861 (N_4861,In_381,In_866);
xor U4862 (N_4862,In_141,In_857);
xnor U4863 (N_4863,In_878,In_366);
nand U4864 (N_4864,In_632,In_893);
nor U4865 (N_4865,In_692,In_193);
and U4866 (N_4866,In_40,In_697);
and U4867 (N_4867,In_134,In_472);
or U4868 (N_4868,In_645,In_580);
and U4869 (N_4869,In_181,In_776);
and U4870 (N_4870,In_62,In_570);
nand U4871 (N_4871,In_245,In_625);
and U4872 (N_4872,In_754,In_129);
nor U4873 (N_4873,In_40,In_401);
and U4874 (N_4874,In_369,In_973);
and U4875 (N_4875,In_476,In_942);
nand U4876 (N_4876,In_589,In_501);
and U4877 (N_4877,In_0,In_900);
xnor U4878 (N_4878,In_755,In_867);
nand U4879 (N_4879,In_888,In_464);
and U4880 (N_4880,In_922,In_453);
or U4881 (N_4881,In_783,In_212);
nor U4882 (N_4882,In_267,In_3);
nor U4883 (N_4883,In_934,In_558);
nor U4884 (N_4884,In_552,In_35);
or U4885 (N_4885,In_367,In_192);
nor U4886 (N_4886,In_279,In_861);
and U4887 (N_4887,In_992,In_924);
and U4888 (N_4888,In_104,In_759);
nor U4889 (N_4889,In_903,In_141);
and U4890 (N_4890,In_568,In_861);
nor U4891 (N_4891,In_646,In_420);
nand U4892 (N_4892,In_239,In_470);
nor U4893 (N_4893,In_683,In_557);
xnor U4894 (N_4894,In_659,In_940);
nor U4895 (N_4895,In_574,In_736);
and U4896 (N_4896,In_409,In_10);
and U4897 (N_4897,In_656,In_652);
or U4898 (N_4898,In_570,In_423);
or U4899 (N_4899,In_324,In_399);
or U4900 (N_4900,In_913,In_636);
or U4901 (N_4901,In_650,In_919);
nand U4902 (N_4902,In_218,In_623);
or U4903 (N_4903,In_90,In_700);
nor U4904 (N_4904,In_675,In_366);
nand U4905 (N_4905,In_367,In_36);
xor U4906 (N_4906,In_828,In_65);
nor U4907 (N_4907,In_260,In_336);
nand U4908 (N_4908,In_771,In_694);
nor U4909 (N_4909,In_315,In_146);
and U4910 (N_4910,In_23,In_563);
nand U4911 (N_4911,In_762,In_583);
nand U4912 (N_4912,In_977,In_702);
nand U4913 (N_4913,In_101,In_527);
xor U4914 (N_4914,In_132,In_484);
nor U4915 (N_4915,In_481,In_797);
and U4916 (N_4916,In_606,In_811);
or U4917 (N_4917,In_812,In_876);
and U4918 (N_4918,In_584,In_706);
nor U4919 (N_4919,In_592,In_719);
nor U4920 (N_4920,In_931,In_973);
and U4921 (N_4921,In_130,In_237);
nor U4922 (N_4922,In_874,In_858);
nor U4923 (N_4923,In_229,In_861);
nand U4924 (N_4924,In_780,In_459);
or U4925 (N_4925,In_7,In_837);
and U4926 (N_4926,In_69,In_727);
and U4927 (N_4927,In_987,In_161);
nor U4928 (N_4928,In_166,In_410);
nor U4929 (N_4929,In_471,In_223);
nand U4930 (N_4930,In_707,In_635);
nor U4931 (N_4931,In_247,In_638);
xnor U4932 (N_4932,In_782,In_543);
nand U4933 (N_4933,In_218,In_830);
nand U4934 (N_4934,In_181,In_637);
and U4935 (N_4935,In_378,In_945);
nor U4936 (N_4936,In_188,In_620);
nand U4937 (N_4937,In_931,In_991);
nand U4938 (N_4938,In_578,In_807);
nand U4939 (N_4939,In_539,In_927);
and U4940 (N_4940,In_9,In_260);
nand U4941 (N_4941,In_493,In_654);
nand U4942 (N_4942,In_491,In_333);
or U4943 (N_4943,In_473,In_350);
or U4944 (N_4944,In_322,In_370);
or U4945 (N_4945,In_689,In_472);
nor U4946 (N_4946,In_770,In_708);
and U4947 (N_4947,In_351,In_626);
and U4948 (N_4948,In_302,In_18);
or U4949 (N_4949,In_988,In_441);
nand U4950 (N_4950,In_938,In_58);
nand U4951 (N_4951,In_157,In_761);
nand U4952 (N_4952,In_185,In_1);
and U4953 (N_4953,In_357,In_658);
nand U4954 (N_4954,In_501,In_554);
and U4955 (N_4955,In_240,In_109);
nand U4956 (N_4956,In_398,In_418);
nor U4957 (N_4957,In_259,In_499);
nand U4958 (N_4958,In_419,In_861);
and U4959 (N_4959,In_311,In_163);
and U4960 (N_4960,In_684,In_239);
nor U4961 (N_4961,In_313,In_699);
xnor U4962 (N_4962,In_703,In_830);
nand U4963 (N_4963,In_680,In_469);
nor U4964 (N_4964,In_378,In_274);
nor U4965 (N_4965,In_237,In_193);
nand U4966 (N_4966,In_669,In_303);
nand U4967 (N_4967,In_683,In_398);
or U4968 (N_4968,In_10,In_725);
or U4969 (N_4969,In_764,In_679);
nor U4970 (N_4970,In_918,In_892);
and U4971 (N_4971,In_591,In_412);
nand U4972 (N_4972,In_981,In_535);
xnor U4973 (N_4973,In_727,In_441);
nand U4974 (N_4974,In_723,In_179);
nor U4975 (N_4975,In_976,In_268);
and U4976 (N_4976,In_85,In_391);
nand U4977 (N_4977,In_508,In_404);
and U4978 (N_4978,In_138,In_467);
nor U4979 (N_4979,In_797,In_532);
or U4980 (N_4980,In_588,In_234);
xnor U4981 (N_4981,In_300,In_58);
nor U4982 (N_4982,In_693,In_436);
and U4983 (N_4983,In_158,In_313);
or U4984 (N_4984,In_225,In_0);
and U4985 (N_4985,In_640,In_648);
nor U4986 (N_4986,In_742,In_626);
xnor U4987 (N_4987,In_411,In_968);
nand U4988 (N_4988,In_516,In_395);
or U4989 (N_4989,In_843,In_318);
nand U4990 (N_4990,In_654,In_848);
nand U4991 (N_4991,In_86,In_11);
nand U4992 (N_4992,In_568,In_770);
nor U4993 (N_4993,In_826,In_454);
nor U4994 (N_4994,In_380,In_196);
or U4995 (N_4995,In_509,In_541);
nand U4996 (N_4996,In_678,In_899);
or U4997 (N_4997,In_443,In_572);
or U4998 (N_4998,In_625,In_412);
nor U4999 (N_4999,In_833,In_195);
xnor U5000 (N_5000,N_4141,N_4790);
or U5001 (N_5001,N_1643,N_1290);
or U5002 (N_5002,N_2694,N_3601);
or U5003 (N_5003,N_227,N_4789);
nor U5004 (N_5004,N_1983,N_2673);
or U5005 (N_5005,N_1667,N_3783);
or U5006 (N_5006,N_1442,N_1517);
nor U5007 (N_5007,N_51,N_914);
nand U5008 (N_5008,N_967,N_702);
nand U5009 (N_5009,N_1619,N_4546);
or U5010 (N_5010,N_4022,N_1977);
or U5011 (N_5011,N_4753,N_1483);
and U5012 (N_5012,N_4286,N_735);
nor U5013 (N_5013,N_2716,N_167);
nor U5014 (N_5014,N_4669,N_1536);
nand U5015 (N_5015,N_624,N_2642);
xor U5016 (N_5016,N_3703,N_4820);
nand U5017 (N_5017,N_3850,N_3643);
and U5018 (N_5018,N_4493,N_4545);
and U5019 (N_5019,N_4154,N_1408);
and U5020 (N_5020,N_4876,N_2895);
and U5021 (N_5021,N_378,N_2789);
nor U5022 (N_5022,N_2674,N_2986);
or U5023 (N_5023,N_3003,N_4948);
nand U5024 (N_5024,N_1644,N_3539);
xnor U5025 (N_5025,N_2560,N_1836);
xor U5026 (N_5026,N_1126,N_779);
nand U5027 (N_5027,N_1671,N_4391);
nand U5028 (N_5028,N_2045,N_682);
and U5029 (N_5029,N_262,N_3002);
and U5030 (N_5030,N_1469,N_949);
and U5031 (N_5031,N_2484,N_3927);
nor U5032 (N_5032,N_1832,N_41);
and U5033 (N_5033,N_4702,N_2593);
or U5034 (N_5034,N_2918,N_1268);
nor U5035 (N_5035,N_3588,N_3335);
nor U5036 (N_5036,N_486,N_115);
nand U5037 (N_5037,N_132,N_2960);
xor U5038 (N_5038,N_2909,N_2878);
and U5039 (N_5039,N_672,N_2393);
nand U5040 (N_5040,N_3397,N_4288);
or U5041 (N_5041,N_739,N_4840);
nand U5042 (N_5042,N_286,N_3647);
nand U5043 (N_5043,N_4394,N_1681);
nor U5044 (N_5044,N_1169,N_3175);
or U5045 (N_5045,N_222,N_4745);
nand U5046 (N_5046,N_1295,N_2815);
or U5047 (N_5047,N_4728,N_279);
nor U5048 (N_5048,N_57,N_4479);
nor U5049 (N_5049,N_1645,N_148);
xor U5050 (N_5050,N_1436,N_2804);
nand U5051 (N_5051,N_3879,N_398);
and U5052 (N_5052,N_368,N_1621);
or U5053 (N_5053,N_442,N_4256);
nor U5054 (N_5054,N_4945,N_4017);
and U5055 (N_5055,N_542,N_1624);
or U5056 (N_5056,N_601,N_135);
nor U5057 (N_5057,N_2559,N_1500);
and U5058 (N_5058,N_2355,N_1754);
nand U5059 (N_5059,N_3457,N_891);
or U5060 (N_5060,N_3293,N_3901);
or U5061 (N_5061,N_1273,N_1193);
nand U5062 (N_5062,N_2055,N_3764);
and U5063 (N_5063,N_2582,N_900);
xor U5064 (N_5064,N_2380,N_817);
nor U5065 (N_5065,N_3646,N_1715);
and U5066 (N_5066,N_2797,N_3091);
xnor U5067 (N_5067,N_736,N_4796);
nand U5068 (N_5068,N_3395,N_4240);
or U5069 (N_5069,N_3778,N_1808);
and U5070 (N_5070,N_2759,N_4261);
nand U5071 (N_5071,N_3219,N_2284);
nor U5072 (N_5072,N_2607,N_1630);
and U5073 (N_5073,N_4102,N_4881);
nor U5074 (N_5074,N_800,N_2390);
or U5075 (N_5075,N_3722,N_884);
or U5076 (N_5076,N_1368,N_1209);
nand U5077 (N_5077,N_1385,N_4140);
or U5078 (N_5078,N_358,N_1838);
or U5079 (N_5079,N_694,N_1943);
nor U5080 (N_5080,N_4594,N_4826);
nor U5081 (N_5081,N_3208,N_4041);
xor U5082 (N_5082,N_1378,N_4424);
and U5083 (N_5083,N_1131,N_4720);
nand U5084 (N_5084,N_677,N_1192);
and U5085 (N_5085,N_2760,N_4848);
nand U5086 (N_5086,N_1197,N_1758);
xnor U5087 (N_5087,N_1661,N_1902);
or U5088 (N_5088,N_487,N_1918);
nand U5089 (N_5089,N_1297,N_3960);
or U5090 (N_5090,N_1354,N_2128);
and U5091 (N_5091,N_4201,N_3987);
nand U5092 (N_5092,N_669,N_313);
xnor U5093 (N_5093,N_341,N_3076);
nand U5094 (N_5094,N_3887,N_3513);
xnor U5095 (N_5095,N_942,N_3865);
nor U5096 (N_5096,N_4588,N_2719);
and U5097 (N_5097,N_4356,N_4606);
nor U5098 (N_5098,N_307,N_2268);
nand U5099 (N_5099,N_3873,N_2339);
nand U5100 (N_5100,N_372,N_2098);
and U5101 (N_5101,N_1413,N_1646);
nand U5102 (N_5102,N_4412,N_1694);
or U5103 (N_5103,N_3109,N_49);
or U5104 (N_5104,N_1708,N_4455);
nand U5105 (N_5105,N_1878,N_2327);
xnor U5106 (N_5106,N_1560,N_646);
or U5107 (N_5107,N_929,N_1084);
or U5108 (N_5108,N_314,N_4747);
or U5109 (N_5109,N_274,N_3518);
and U5110 (N_5110,N_4451,N_3436);
xor U5111 (N_5111,N_3452,N_4647);
nor U5112 (N_5112,N_2876,N_4111);
or U5113 (N_5113,N_614,N_4856);
nor U5114 (N_5114,N_724,N_1805);
nand U5115 (N_5115,N_2467,N_4862);
xnor U5116 (N_5116,N_1405,N_4711);
nor U5117 (N_5117,N_1157,N_3123);
nor U5118 (N_5118,N_4357,N_4683);
and U5119 (N_5119,N_4536,N_2584);
xor U5120 (N_5120,N_3692,N_4408);
nand U5121 (N_5121,N_3027,N_4020);
and U5122 (N_5122,N_4272,N_3822);
and U5123 (N_5123,N_3507,N_1831);
nand U5124 (N_5124,N_937,N_2325);
nor U5125 (N_5125,N_1230,N_3196);
and U5126 (N_5126,N_4957,N_3502);
nand U5127 (N_5127,N_880,N_3306);
nand U5128 (N_5128,N_3762,N_3939);
xor U5129 (N_5129,N_2225,N_4136);
nand U5130 (N_5130,N_3500,N_3311);
nand U5131 (N_5131,N_367,N_2419);
or U5132 (N_5132,N_1728,N_3754);
or U5133 (N_5133,N_2509,N_3991);
nand U5134 (N_5134,N_4284,N_3970);
nand U5135 (N_5135,N_4153,N_1925);
and U5136 (N_5136,N_342,N_3357);
and U5137 (N_5137,N_4215,N_4322);
and U5138 (N_5138,N_2323,N_2476);
nor U5139 (N_5139,N_3984,N_2839);
nor U5140 (N_5140,N_2254,N_4997);
nand U5141 (N_5141,N_2543,N_2326);
and U5142 (N_5142,N_3679,N_3508);
and U5143 (N_5143,N_23,N_4822);
nand U5144 (N_5144,N_1716,N_2309);
nor U5145 (N_5145,N_1050,N_2657);
and U5146 (N_5146,N_64,N_3134);
and U5147 (N_5147,N_553,N_1799);
nand U5148 (N_5148,N_3283,N_360);
nand U5149 (N_5149,N_3654,N_2258);
nor U5150 (N_5150,N_4057,N_3444);
or U5151 (N_5151,N_1244,N_4797);
nor U5152 (N_5152,N_3857,N_4828);
nor U5153 (N_5153,N_3846,N_1916);
xor U5154 (N_5154,N_4315,N_1402);
nand U5155 (N_5155,N_1870,N_2205);
nor U5156 (N_5156,N_4704,N_4506);
nand U5157 (N_5157,N_232,N_861);
or U5158 (N_5158,N_3463,N_1818);
and U5159 (N_5159,N_3586,N_4331);
and U5160 (N_5160,N_4898,N_3828);
or U5161 (N_5161,N_4459,N_275);
nor U5162 (N_5162,N_837,N_1574);
nand U5163 (N_5163,N_4958,N_2247);
and U5164 (N_5164,N_3303,N_43);
nand U5165 (N_5165,N_44,N_3845);
nand U5166 (N_5166,N_1163,N_3354);
and U5167 (N_5167,N_4395,N_1038);
or U5168 (N_5168,N_1830,N_4043);
or U5169 (N_5169,N_4398,N_4842);
nor U5170 (N_5170,N_4879,N_3182);
nand U5171 (N_5171,N_3920,N_1276);
nand U5172 (N_5172,N_48,N_2293);
or U5173 (N_5173,N_2793,N_1480);
or U5174 (N_5174,N_2084,N_2880);
and U5175 (N_5175,N_261,N_4837);
nand U5176 (N_5176,N_2670,N_670);
and U5177 (N_5177,N_4120,N_3267);
nand U5178 (N_5178,N_2852,N_3936);
nor U5179 (N_5179,N_490,N_2538);
nor U5180 (N_5180,N_3995,N_1837);
nor U5181 (N_5181,N_4283,N_2263);
or U5182 (N_5182,N_4280,N_4819);
and U5183 (N_5183,N_2978,N_2398);
xnor U5184 (N_5184,N_3546,N_3766);
or U5185 (N_5185,N_2611,N_2154);
and U5186 (N_5186,N_4426,N_632);
nor U5187 (N_5187,N_3514,N_3565);
nand U5188 (N_5188,N_2495,N_3593);
nand U5189 (N_5189,N_4882,N_1284);
nand U5190 (N_5190,N_532,N_1550);
nand U5191 (N_5191,N_4291,N_747);
nand U5192 (N_5192,N_1872,N_2099);
and U5193 (N_5193,N_2302,N_893);
and U5194 (N_5194,N_4860,N_3009);
nand U5195 (N_5195,N_4608,N_1191);
nor U5196 (N_5196,N_1583,N_306);
and U5197 (N_5197,N_3810,N_3046);
and U5198 (N_5198,N_3435,N_328);
and U5199 (N_5199,N_3363,N_2540);
xnor U5200 (N_5200,N_4325,N_462);
nand U5201 (N_5201,N_4192,N_500);
nor U5202 (N_5202,N_2157,N_4962);
nor U5203 (N_5203,N_242,N_2028);
and U5204 (N_5204,N_4213,N_2342);
nor U5205 (N_5205,N_3569,N_895);
and U5206 (N_5206,N_1357,N_2596);
nor U5207 (N_5207,N_1121,N_3524);
nor U5208 (N_5208,N_4501,N_4562);
nand U5209 (N_5209,N_1729,N_475);
xnor U5210 (N_5210,N_1589,N_16);
nand U5211 (N_5211,N_2452,N_2022);
and U5212 (N_5212,N_1320,N_2563);
nor U5213 (N_5213,N_1425,N_656);
and U5214 (N_5214,N_1102,N_1665);
and U5215 (N_5215,N_1961,N_457);
xor U5216 (N_5216,N_158,N_928);
or U5217 (N_5217,N_1374,N_3305);
nand U5218 (N_5218,N_4760,N_3634);
and U5219 (N_5219,N_325,N_740);
xnor U5220 (N_5220,N_449,N_3202);
and U5221 (N_5221,N_2070,N_1675);
or U5222 (N_5222,N_224,N_2828);
or U5223 (N_5223,N_2234,N_3759);
nand U5224 (N_5224,N_2021,N_3146);
nand U5225 (N_5225,N_17,N_2542);
and U5226 (N_5226,N_3087,N_2358);
and U5227 (N_5227,N_4666,N_4089);
nand U5228 (N_5228,N_1924,N_2048);
nand U5229 (N_5229,N_4973,N_4337);
or U5230 (N_5230,N_2615,N_750);
nor U5231 (N_5231,N_2438,N_1492);
nand U5232 (N_5232,N_2377,N_4684);
and U5233 (N_5233,N_3730,N_828);
nand U5234 (N_5234,N_506,N_3256);
nand U5235 (N_5235,N_3536,N_1825);
xnor U5236 (N_5236,N_145,N_4260);
or U5237 (N_5237,N_3095,N_906);
nand U5238 (N_5238,N_4134,N_1979);
nand U5239 (N_5239,N_2466,N_4067);
nor U5240 (N_5240,N_1265,N_2241);
nor U5241 (N_5241,N_4338,N_4174);
nor U5242 (N_5242,N_3434,N_4276);
nor U5243 (N_5243,N_3125,N_533);
nand U5244 (N_5244,N_2117,N_3322);
and U5245 (N_5245,N_221,N_1605);
and U5246 (N_5246,N_1108,N_1835);
or U5247 (N_5247,N_2279,N_1228);
or U5248 (N_5248,N_4094,N_1850);
nor U5249 (N_5249,N_4904,N_968);
and U5250 (N_5250,N_3605,N_2822);
xor U5251 (N_5251,N_2250,N_4891);
and U5252 (N_5252,N_776,N_2262);
and U5253 (N_5253,N_4661,N_4919);
or U5254 (N_5254,N_4777,N_4155);
nand U5255 (N_5255,N_4574,N_777);
nand U5256 (N_5256,N_4734,N_3408);
nor U5257 (N_5257,N_4540,N_2100);
xor U5258 (N_5258,N_3742,N_822);
xnor U5259 (N_5259,N_3054,N_4042);
nor U5260 (N_5260,N_3410,N_4183);
nor U5261 (N_5261,N_821,N_304);
nor U5262 (N_5262,N_4964,N_4034);
nor U5263 (N_5263,N_876,N_1557);
and U5264 (N_5264,N_2330,N_4393);
nand U5265 (N_5265,N_155,N_3271);
nand U5266 (N_5266,N_4248,N_4610);
nand U5267 (N_5267,N_416,N_2827);
nand U5268 (N_5268,N_4477,N_3542);
xor U5269 (N_5269,N_1148,N_3616);
xor U5270 (N_5270,N_3460,N_3250);
nand U5271 (N_5271,N_3420,N_4653);
nand U5272 (N_5272,N_4524,N_4385);
nor U5273 (N_5273,N_1967,N_1321);
and U5274 (N_5274,N_4366,N_2388);
or U5275 (N_5275,N_1648,N_1606);
nand U5276 (N_5276,N_3118,N_4432);
nand U5277 (N_5277,N_948,N_1972);
and U5278 (N_5278,N_4643,N_4214);
nand U5279 (N_5279,N_3983,N_1366);
and U5280 (N_5280,N_1988,N_4895);
and U5281 (N_5281,N_4399,N_4145);
nor U5282 (N_5282,N_3906,N_2744);
nand U5283 (N_5283,N_3346,N_1781);
nand U5284 (N_5284,N_3674,N_2905);
nand U5285 (N_5285,N_3607,N_288);
and U5286 (N_5286,N_105,N_1501);
nor U5287 (N_5287,N_2619,N_2078);
nand U5288 (N_5288,N_3060,N_1474);
or U5289 (N_5289,N_4347,N_4763);
nand U5290 (N_5290,N_1670,N_1677);
nand U5291 (N_5291,N_3682,N_4770);
nand U5292 (N_5292,N_3882,N_433);
and U5293 (N_5293,N_947,N_3177);
and U5294 (N_5294,N_992,N_1003);
nor U5295 (N_5295,N_1072,N_4090);
and U5296 (N_5296,N_4285,N_4795);
or U5297 (N_5297,N_4269,N_760);
nand U5298 (N_5298,N_1515,N_2979);
and U5299 (N_5299,N_4780,N_2981);
nor U5300 (N_5300,N_4488,N_2965);
or U5301 (N_5301,N_2465,N_390);
and U5302 (N_5302,N_2057,N_756);
nand U5303 (N_5303,N_4405,N_2901);
and U5304 (N_5304,N_2230,N_50);
nor U5305 (N_5305,N_63,N_933);
or U5306 (N_5306,N_2949,N_3467);
nand U5307 (N_5307,N_188,N_3688);
nand U5308 (N_5308,N_4060,N_4026);
nor U5309 (N_5309,N_1327,N_3591);
or U5310 (N_5310,N_1945,N_576);
and U5311 (N_5311,N_3409,N_4100);
and U5312 (N_5312,N_160,N_4474);
nand U5313 (N_5313,N_2816,N_365);
and U5314 (N_5314,N_4465,N_2726);
nor U5315 (N_5315,N_4314,N_4362);
or U5316 (N_5316,N_4457,N_4645);
nor U5317 (N_5317,N_1778,N_1032);
nor U5318 (N_5318,N_4952,N_4577);
and U5319 (N_5319,N_1100,N_1154);
nand U5320 (N_5320,N_4438,N_3347);
xnor U5321 (N_5321,N_3568,N_2591);
nor U5322 (N_5322,N_2303,N_2718);
nor U5323 (N_5323,N_1426,N_3505);
nand U5324 (N_5324,N_2900,N_3401);
and U5325 (N_5325,N_2491,N_693);
xnor U5326 (N_5326,N_3008,N_2191);
or U5327 (N_5327,N_1172,N_1793);
and U5328 (N_5328,N_1308,N_137);
or U5329 (N_5329,N_1625,N_2005);
nor U5330 (N_5330,N_1748,N_2654);
nand U5331 (N_5331,N_1067,N_419);
nor U5332 (N_5332,N_4230,N_1203);
nor U5333 (N_5333,N_4496,N_4107);
or U5334 (N_5334,N_1790,N_3615);
and U5335 (N_5335,N_3221,N_3900);
and U5336 (N_5336,N_2834,N_996);
nor U5337 (N_5337,N_4494,N_271);
or U5338 (N_5338,N_4482,N_1543);
nor U5339 (N_5339,N_4625,N_1356);
nand U5340 (N_5340,N_4264,N_4278);
or U5341 (N_5341,N_2031,N_872);
nor U5342 (N_5342,N_572,N_2842);
or U5343 (N_5343,N_4939,N_259);
or U5344 (N_5344,N_428,N_2568);
or U5345 (N_5345,N_345,N_4676);
and U5346 (N_5346,N_978,N_1942);
and U5347 (N_5347,N_3344,N_4656);
nor U5348 (N_5348,N_4859,N_2516);
or U5349 (N_5349,N_2308,N_2885);
nand U5350 (N_5350,N_1887,N_97);
nor U5351 (N_5351,N_2032,N_1948);
xor U5352 (N_5352,N_201,N_1208);
nand U5353 (N_5353,N_4658,N_2938);
nand U5354 (N_5354,N_1238,N_1957);
and U5355 (N_5355,N_4596,N_19);
nand U5356 (N_5356,N_2104,N_1705);
xnor U5357 (N_5357,N_1745,N_1651);
nand U5358 (N_5358,N_482,N_4148);
nand U5359 (N_5359,N_1390,N_1787);
and U5360 (N_5360,N_3932,N_1343);
or U5361 (N_5361,N_3486,N_1188);
or U5362 (N_5362,N_2518,N_4023);
and U5363 (N_5363,N_4146,N_1083);
nand U5364 (N_5364,N_432,N_3331);
xnor U5365 (N_5365,N_3661,N_241);
nor U5366 (N_5366,N_1264,N_1987);
or U5367 (N_5367,N_1636,N_1164);
or U5368 (N_5368,N_91,N_1615);
and U5369 (N_5369,N_2210,N_293);
nor U5370 (N_5370,N_612,N_2149);
and U5371 (N_5371,N_517,N_1575);
and U5372 (N_5372,N_1212,N_1305);
or U5373 (N_5373,N_391,N_2713);
or U5374 (N_5374,N_4374,N_1666);
and U5375 (N_5375,N_3971,N_855);
nand U5376 (N_5376,N_4088,N_4887);
or U5377 (N_5377,N_2894,N_3242);
nand U5378 (N_5378,N_3416,N_2734);
nor U5379 (N_5379,N_2026,N_379);
or U5380 (N_5380,N_4342,N_4270);
xor U5381 (N_5381,N_3281,N_889);
nor U5382 (N_5382,N_4360,N_754);
or U5383 (N_5383,N_722,N_3245);
nor U5384 (N_5384,N_2482,N_4951);
nand U5385 (N_5385,N_2232,N_3114);
nor U5386 (N_5386,N_4363,N_4406);
nand U5387 (N_5387,N_1056,N_1658);
and U5388 (N_5388,N_3547,N_1029);
nor U5389 (N_5389,N_2817,N_3890);
or U5390 (N_5390,N_1272,N_194);
xnor U5391 (N_5391,N_3482,N_4470);
nand U5392 (N_5392,N_4975,N_396);
nand U5393 (N_5393,N_4581,N_3288);
nand U5394 (N_5394,N_1250,N_2093);
and U5395 (N_5395,N_42,N_885);
nor U5396 (N_5396,N_4924,N_2521);
and U5397 (N_5397,N_705,N_2075);
or U5398 (N_5398,N_3360,N_2397);
nor U5399 (N_5399,N_732,N_4323);
or U5400 (N_5400,N_3774,N_4985);
nand U5401 (N_5401,N_2984,N_123);
nand U5402 (N_5402,N_1246,N_3537);
and U5403 (N_5403,N_3138,N_1037);
and U5404 (N_5404,N_3868,N_2110);
or U5405 (N_5405,N_1770,N_2081);
nor U5406 (N_5406,N_1706,N_618);
or U5407 (N_5407,N_2790,N_4007);
and U5408 (N_5408,N_4851,N_3907);
nor U5409 (N_5409,N_3299,N_1472);
nand U5410 (N_5410,N_4452,N_1296);
nor U5411 (N_5411,N_2599,N_3617);
or U5412 (N_5412,N_3244,N_954);
nand U5413 (N_5413,N_406,N_2228);
or U5414 (N_5414,N_698,N_2993);
xnor U5415 (N_5415,N_3328,N_676);
xnor U5416 (N_5416,N_2146,N_2411);
or U5417 (N_5417,N_2576,N_4724);
nor U5418 (N_5418,N_4708,N_3213);
and U5419 (N_5419,N_3998,N_3628);
nor U5420 (N_5420,N_4103,N_4693);
nand U5421 (N_5421,N_1608,N_2427);
nor U5422 (N_5422,N_1846,N_1464);
xor U5423 (N_5423,N_710,N_3205);
and U5424 (N_5424,N_3701,N_2025);
nor U5425 (N_5425,N_300,N_901);
nor U5426 (N_5426,N_3665,N_2150);
nand U5427 (N_5427,N_661,N_2689);
nor U5428 (N_5428,N_1933,N_1444);
and U5429 (N_5429,N_1855,N_3950);
nand U5430 (N_5430,N_1668,N_4810);
nand U5431 (N_5431,N_4492,N_3997);
nand U5432 (N_5432,N_1047,N_1481);
nor U5433 (N_5433,N_2211,N_4304);
or U5434 (N_5434,N_4204,N_1155);
and U5435 (N_5435,N_1069,N_2366);
or U5436 (N_5436,N_603,N_4361);
and U5437 (N_5437,N_4871,N_1427);
or U5438 (N_5438,N_1819,N_4462);
nand U5439 (N_5439,N_2964,N_3375);
nor U5440 (N_5440,N_1281,N_3919);
and U5441 (N_5441,N_1095,N_4458);
xor U5442 (N_5442,N_3384,N_413);
and U5443 (N_5443,N_470,N_3449);
nand U5444 (N_5444,N_4222,N_2068);
and U5445 (N_5445,N_1842,N_712);
nor U5446 (N_5446,N_899,N_4650);
or U5447 (N_5447,N_3585,N_2983);
or U5448 (N_5448,N_294,N_263);
or U5449 (N_5449,N_2620,N_4127);
nor U5450 (N_5450,N_1704,N_4138);
nand U5451 (N_5451,N_82,N_3749);
and U5452 (N_5452,N_4101,N_3272);
nand U5453 (N_5453,N_3642,N_443);
or U5454 (N_5454,N_2526,N_205);
nand U5455 (N_5455,N_4239,N_420);
and U5456 (N_5456,N_1487,N_1210);
or U5457 (N_5457,N_4755,N_3222);
xor U5458 (N_5458,N_1657,N_574);
xnor U5459 (N_5459,N_1586,N_3402);
nand U5460 (N_5460,N_169,N_4227);
nor U5461 (N_5461,N_2317,N_2001);
xor U5462 (N_5462,N_2209,N_2875);
nor U5463 (N_5463,N_960,N_3657);
nor U5464 (N_5464,N_2687,N_1847);
nand U5465 (N_5465,N_3162,N_1314);
nand U5466 (N_5466,N_1007,N_3956);
nand U5467 (N_5467,N_886,N_374);
or U5468 (N_5468,N_4265,N_3558);
nand U5469 (N_5469,N_2945,N_1400);
nor U5470 (N_5470,N_2387,N_3494);
nor U5471 (N_5471,N_1404,N_4626);
nand U5472 (N_5472,N_383,N_18);
and U5473 (N_5473,N_630,N_2396);
nand U5474 (N_5474,N_3317,N_2982);
xor U5475 (N_5475,N_25,N_4460);
nand U5476 (N_5476,N_680,N_1291);
nor U5477 (N_5477,N_2315,N_1269);
and U5478 (N_5478,N_3512,N_478);
or U5479 (N_5479,N_1386,N_2162);
xnor U5480 (N_5480,N_4427,N_361);
and U5481 (N_5481,N_61,N_2089);
and U5482 (N_5482,N_1361,N_2679);
nand U5483 (N_5483,N_3072,N_3116);
nor U5484 (N_5484,N_3613,N_2490);
and U5485 (N_5485,N_1399,N_439);
or U5486 (N_5486,N_708,N_2548);
and U5487 (N_5487,N_1490,N_2635);
and U5488 (N_5488,N_679,N_4803);
or U5489 (N_5489,N_589,N_2818);
or U5490 (N_5490,N_2376,N_2043);
xor U5491 (N_5491,N_2450,N_1616);
or U5492 (N_5492,N_969,N_3127);
nand U5493 (N_5493,N_1289,N_793);
nor U5494 (N_5494,N_931,N_4933);
nand U5495 (N_5495,N_4420,N_4909);
nor U5496 (N_5496,N_3724,N_1422);
nor U5497 (N_5497,N_647,N_3578);
xnor U5498 (N_5498,N_4422,N_2101);
nand U5499 (N_5499,N_3117,N_788);
or U5500 (N_5500,N_2318,N_2989);
nor U5501 (N_5501,N_2115,N_3740);
and U5502 (N_5502,N_184,N_1590);
nand U5503 (N_5503,N_4317,N_4124);
and U5504 (N_5504,N_4838,N_1617);
and U5505 (N_5505,N_1075,N_1762);
and U5506 (N_5506,N_1759,N_1952);
and U5507 (N_5507,N_3230,N_4805);
nand U5508 (N_5508,N_2264,N_2547);
nand U5509 (N_5509,N_29,N_1719);
nand U5510 (N_5510,N_4994,N_4274);
or U5511 (N_5511,N_761,N_231);
and U5512 (N_5512,N_2752,N_849);
nor U5513 (N_5513,N_2190,N_493);
xor U5514 (N_5514,N_4984,N_1053);
and U5515 (N_5515,N_2737,N_4311);
or U5516 (N_5516,N_1479,N_2893);
and U5517 (N_5517,N_1329,N_4055);
or U5518 (N_5518,N_2200,N_3902);
nor U5519 (N_5519,N_4671,N_1485);
and U5520 (N_5520,N_1982,N_2215);
or U5521 (N_5521,N_1755,N_2931);
nand U5522 (N_5522,N_4530,N_4431);
or U5523 (N_5523,N_187,N_2610);
and U5524 (N_5524,N_2248,N_3496);
xnor U5525 (N_5525,N_4814,N_3019);
nand U5526 (N_5526,N_1410,N_2567);
nor U5527 (N_5527,N_1457,N_3240);
or U5528 (N_5528,N_4762,N_2928);
or U5529 (N_5529,N_1546,N_4350);
nand U5530 (N_5530,N_448,N_3619);
nor U5531 (N_5531,N_3816,N_2275);
or U5532 (N_5532,N_3470,N_1798);
nand U5533 (N_5533,N_4371,N_270);
xor U5534 (N_5534,N_308,N_4097);
nor U5535 (N_5535,N_1824,N_4677);
nor U5536 (N_5536,N_317,N_4813);
nand U5537 (N_5537,N_4231,N_4950);
xnor U5538 (N_5538,N_13,N_3993);
nand U5539 (N_5539,N_3308,N_3430);
nor U5540 (N_5540,N_1683,N_3455);
or U5541 (N_5541,N_3789,N_4093);
nor U5542 (N_5542,N_1727,N_3479);
or U5543 (N_5543,N_2823,N_3119);
nand U5544 (N_5544,N_3122,N_3057);
or U5545 (N_5545,N_1350,N_198);
and U5546 (N_5546,N_2972,N_4247);
nand U5547 (N_5547,N_4687,N_2936);
and U5548 (N_5548,N_2090,N_1672);
or U5549 (N_5549,N_1304,N_2870);
and U5550 (N_5550,N_4212,N_58);
nor U5551 (N_5551,N_3655,N_4742);
or U5552 (N_5552,N_4792,N_728);
or U5553 (N_5553,N_650,N_2196);
or U5554 (N_5554,N_798,N_797);
xor U5555 (N_5555,N_1865,N_2629);
or U5556 (N_5556,N_4232,N_806);
or U5557 (N_5557,N_1332,N_3492);
and U5558 (N_5558,N_27,N_2757);
or U5559 (N_5559,N_741,N_719);
nor U5560 (N_5560,N_4965,N_1226);
and U5561 (N_5561,N_1372,N_1937);
or U5562 (N_5562,N_30,N_2939);
nor U5563 (N_5563,N_1449,N_1080);
or U5564 (N_5564,N_1691,N_3911);
nand U5565 (N_5565,N_2036,N_2356);
nand U5566 (N_5566,N_4392,N_329);
or U5567 (N_5567,N_1851,N_1507);
and U5568 (N_5568,N_3753,N_749);
and U5569 (N_5569,N_1496,N_823);
xnor U5570 (N_5570,N_3946,N_2785);
nor U5571 (N_5571,N_3632,N_1534);
nand U5572 (N_5572,N_2430,N_1774);
or U5573 (N_5573,N_878,N_3115);
xnor U5574 (N_5574,N_512,N_2217);
nor U5575 (N_5575,N_762,N_3398);
or U5576 (N_5576,N_236,N_3336);
and U5577 (N_5577,N_2172,N_1392);
and U5578 (N_5578,N_3179,N_4870);
nand U5579 (N_5579,N_2261,N_2227);
and U5580 (N_5580,N_3968,N_3501);
nor U5581 (N_5581,N_562,N_423);
nand U5582 (N_5582,N_303,N_4833);
nand U5583 (N_5583,N_790,N_2189);
and U5584 (N_5584,N_375,N_2016);
and U5585 (N_5585,N_2848,N_530);
nand U5586 (N_5586,N_2201,N_2522);
and U5587 (N_5587,N_4396,N_2130);
and U5588 (N_5588,N_1712,N_592);
or U5589 (N_5589,N_2754,N_4365);
nor U5590 (N_5590,N_1877,N_1883);
nand U5591 (N_5591,N_3650,N_4397);
or U5592 (N_5592,N_2410,N_1690);
or U5593 (N_5593,N_4599,N_4794);
nor U5594 (N_5594,N_3071,N_1741);
nor U5595 (N_5595,N_3814,N_608);
xor U5596 (N_5596,N_441,N_2766);
nand U5597 (N_5597,N_2237,N_2923);
nor U5598 (N_5598,N_2158,N_2708);
nand U5599 (N_5599,N_3007,N_3652);
xnor U5600 (N_5600,N_4852,N_3768);
and U5601 (N_5601,N_3349,N_3247);
and U5602 (N_5602,N_3419,N_84);
nor U5603 (N_5603,N_2056,N_2202);
nand U5604 (N_5604,N_1214,N_4998);
or U5605 (N_5605,N_1247,N_1581);
and U5606 (N_5606,N_3270,N_3421);
nor U5607 (N_5607,N_3041,N_2866);
nand U5608 (N_5608,N_1213,N_3790);
nand U5609 (N_5609,N_875,N_3566);
nand U5610 (N_5610,N_3135,N_3698);
nand U5611 (N_5611,N_794,N_2943);
nand U5612 (N_5612,N_3387,N_600);
nor U5613 (N_5613,N_1827,N_1090);
and U5614 (N_5614,N_1511,N_874);
nor U5615 (N_5615,N_4597,N_1739);
xnor U5616 (N_5616,N_780,N_2144);
and U5617 (N_5617,N_3251,N_28);
xor U5618 (N_5618,N_2681,N_3760);
and U5619 (N_5619,N_2120,N_848);
and U5620 (N_5620,N_191,N_3105);
nor U5621 (N_5621,N_3437,N_1724);
nor U5622 (N_5622,N_4639,N_3464);
nand U5623 (N_5623,N_4611,N_472);
nor U5624 (N_5624,N_3191,N_1696);
nor U5625 (N_5625,N_3068,N_1985);
nor U5626 (N_5626,N_4176,N_255);
or U5627 (N_5627,N_56,N_4378);
and U5628 (N_5628,N_3713,N_284);
and U5629 (N_5629,N_322,N_2824);
or U5630 (N_5630,N_4341,N_2932);
nand U5631 (N_5631,N_2532,N_464);
or U5632 (N_5632,N_3049,N_2922);
nor U5633 (N_5633,N_2626,N_4857);
or U5634 (N_5634,N_2770,N_4386);
and U5635 (N_5635,N_3083,N_2456);
or U5636 (N_5636,N_2494,N_2997);
nor U5637 (N_5637,N_3090,N_723);
or U5638 (N_5638,N_1020,N_3029);
and U5639 (N_5639,N_4733,N_1005);
xnor U5640 (N_5640,N_3450,N_104);
xor U5641 (N_5641,N_153,N_1176);
and U5642 (N_5642,N_4052,N_311);
and U5643 (N_5643,N_2697,N_3793);
nand U5644 (N_5644,N_3274,N_4955);
or U5645 (N_5645,N_2855,N_3173);
xnor U5646 (N_5646,N_966,N_1954);
nand U5647 (N_5647,N_3711,N_2821);
nor U5648 (N_5648,N_1565,N_197);
or U5649 (N_5649,N_2577,N_22);
xnor U5650 (N_5650,N_718,N_1242);
xnor U5651 (N_5651,N_2954,N_4632);
and U5652 (N_5652,N_4818,N_3280);
xor U5653 (N_5653,N_2590,N_258);
nor U5654 (N_5654,N_4657,N_62);
or U5655 (N_5655,N_3567,N_4085);
and U5656 (N_5656,N_4539,N_4886);
and U5657 (N_5657,N_1377,N_3301);
and U5658 (N_5658,N_0,N_2585);
nand U5659 (N_5659,N_1124,N_4947);
and U5660 (N_5660,N_3459,N_4915);
nor U5661 (N_5661,N_497,N_295);
xor U5662 (N_5662,N_611,N_3192);
xor U5663 (N_5663,N_2840,N_1941);
nand U5664 (N_5664,N_1577,N_4642);
nand U5665 (N_5665,N_4938,N_3772);
nand U5666 (N_5666,N_219,N_2595);
nand U5667 (N_5667,N_2544,N_4220);
nand U5668 (N_5668,N_3266,N_2240);
nor U5669 (N_5669,N_2700,N_585);
nand U5670 (N_5670,N_3587,N_4104);
and U5671 (N_5671,N_4246,N_4108);
nand U5672 (N_5672,N_3326,N_1077);
or U5673 (N_5673,N_516,N_369);
and U5674 (N_5674,N_1876,N_2507);
nor U5675 (N_5675,N_2420,N_3268);
and U5676 (N_5676,N_1736,N_769);
nor U5677 (N_5677,N_3697,N_4487);
nand U5678 (N_5678,N_3757,N_1919);
or U5679 (N_5679,N_3595,N_4224);
nand U5680 (N_5680,N_3214,N_1432);
nor U5681 (N_5681,N_3294,N_4646);
and U5682 (N_5682,N_2433,N_440);
and U5683 (N_5683,N_4772,N_1735);
and U5684 (N_5684,N_3581,N_4765);
xor U5685 (N_5685,N_364,N_2589);
nor U5686 (N_5686,N_1593,N_2648);
or U5687 (N_5687,N_2738,N_1391);
nand U5688 (N_5688,N_3394,N_3499);
and U5689 (N_5689,N_1528,N_3338);
or U5690 (N_5690,N_883,N_1415);
and U5691 (N_5691,N_4132,N_4567);
nand U5692 (N_5692,N_3745,N_4709);
and U5693 (N_5693,N_2957,N_3709);
and U5694 (N_5694,N_4816,N_214);
nor U5695 (N_5695,N_3443,N_4066);
nor U5696 (N_5696,N_3487,N_1347);
nor U5697 (N_5697,N_1733,N_956);
xor U5698 (N_5698,N_2235,N_4197);
nor U5699 (N_5699,N_3073,N_1508);
nor U5700 (N_5700,N_1471,N_1917);
nor U5701 (N_5701,N_4015,N_3238);
nor U5702 (N_5702,N_3325,N_1530);
or U5703 (N_5703,N_2238,N_932);
and U5704 (N_5704,N_1506,N_557);
xor U5705 (N_5705,N_925,N_249);
and U5706 (N_5706,N_2271,N_3819);
or U5707 (N_5707,N_2063,N_3184);
nand U5708 (N_5708,N_3836,N_4699);
nor U5709 (N_5709,N_3893,N_72);
nor U5710 (N_5710,N_2702,N_130);
nor U5711 (N_5711,N_2354,N_3880);
nor U5712 (N_5712,N_4723,N_3037);
nand U5713 (N_5713,N_3018,N_4379);
and U5714 (N_5714,N_2699,N_2486);
and U5715 (N_5715,N_1167,N_4968);
nand U5716 (N_5716,N_504,N_1939);
xor U5717 (N_5717,N_629,N_3241);
nor U5718 (N_5718,N_2343,N_540);
xnor U5719 (N_5719,N_2600,N_3702);
xor U5720 (N_5720,N_2664,N_4651);
xor U5721 (N_5721,N_2801,N_1359);
nand U5722 (N_5722,N_2669,N_4786);
xnor U5723 (N_5723,N_4453,N_3781);
nand U5724 (N_5724,N_210,N_4375);
or U5725 (N_5725,N_812,N_3916);
nand U5726 (N_5726,N_1239,N_3400);
or U5727 (N_5727,N_1312,N_2155);
or U5728 (N_5728,N_2083,N_639);
and U5729 (N_5729,N_386,N_2638);
or U5730 (N_5730,N_1240,N_3686);
nor U5731 (N_5731,N_2017,N_4351);
nor U5732 (N_5732,N_4116,N_791);
nand U5733 (N_5733,N_1303,N_1910);
and U5734 (N_5734,N_213,N_165);
nor U5735 (N_5735,N_4177,N_4552);
and U5736 (N_5736,N_3198,N_2087);
nand U5737 (N_5737,N_1599,N_112);
nand U5738 (N_5738,N_1260,N_1815);
nand U5739 (N_5739,N_1211,N_3432);
and U5740 (N_5740,N_1267,N_626);
nor U5741 (N_5741,N_1430,N_2352);
or U5742 (N_5742,N_3744,N_1027);
or U5743 (N_5743,N_1603,N_4980);
and U5744 (N_5744,N_1369,N_2274);
or U5745 (N_5745,N_3942,N_1074);
nand U5746 (N_5746,N_1179,N_4358);
nor U5747 (N_5747,N_2616,N_2985);
nand U5748 (N_5748,N_2399,N_3653);
or U5749 (N_5749,N_1375,N_3896);
nor U5750 (N_5750,N_1009,N_2423);
or U5751 (N_5751,N_816,N_1771);
or U5752 (N_5752,N_2136,N_1253);
nand U5753 (N_5753,N_2429,N_1491);
or U5754 (N_5754,N_554,N_352);
or U5755 (N_5755,N_3621,N_309);
and U5756 (N_5756,N_3447,N_79);
and U5757 (N_5757,N_2289,N_3779);
nor U5758 (N_5758,N_3441,N_845);
or U5759 (N_5759,N_4614,N_3478);
nor U5760 (N_5760,N_1725,N_3314);
or U5761 (N_5761,N_1088,N_910);
or U5762 (N_5762,N_1236,N_1904);
or U5763 (N_5763,N_2168,N_2375);
nor U5764 (N_5764,N_4205,N_4039);
nor U5765 (N_5765,N_1417,N_1828);
and U5766 (N_5766,N_4696,N_437);
and U5767 (N_5767,N_1039,N_958);
nor U5768 (N_5768,N_2027,N_4196);
and U5769 (N_5769,N_2292,N_4198);
nor U5770 (N_5770,N_2000,N_1489);
nand U5771 (N_5771,N_2572,N_335);
nor U5772 (N_5772,N_2963,N_4618);
or U5773 (N_5773,N_4931,N_1597);
or U5774 (N_5774,N_4144,N_287);
nor U5775 (N_5775,N_3120,N_2550);
or U5776 (N_5776,N_1138,N_4376);
nor U5777 (N_5777,N_896,N_2373);
nor U5778 (N_5778,N_4769,N_3031);
and U5779 (N_5779,N_3818,N_1235);
nand U5780 (N_5780,N_438,N_2379);
nor U5781 (N_5781,N_59,N_2469);
and U5782 (N_5782,N_569,N_1523);
or U5783 (N_5783,N_1044,N_999);
nand U5784 (N_5784,N_4099,N_1010);
and U5785 (N_5785,N_3925,N_3366);
nor U5786 (N_5786,N_1149,N_2704);
nand U5787 (N_5787,N_2774,N_4849);
nand U5788 (N_5788,N_4268,N_3433);
and U5789 (N_5789,N_302,N_4981);
nor U5790 (N_5790,N_4517,N_974);
and U5791 (N_5791,N_1255,N_597);
or U5792 (N_5792,N_3260,N_4555);
nor U5793 (N_5793,N_39,N_4251);
or U5794 (N_5794,N_2039,N_3871);
and U5795 (N_5795,N_2701,N_887);
nor U5796 (N_5796,N_4324,N_582);
nand U5797 (N_5797,N_4685,N_1016);
xnor U5798 (N_5798,N_3318,N_3549);
and U5799 (N_5799,N_2703,N_4827);
nor U5800 (N_5800,N_2627,N_2883);
or U5801 (N_5801,N_1997,N_2749);
or U5802 (N_5802,N_3065,N_3491);
or U5803 (N_5803,N_2511,N_4434);
or U5804 (N_5804,N_4532,N_578);
xor U5805 (N_5805,N_3705,N_4208);
nor U5806 (N_5806,N_2363,N_80);
xor U5807 (N_5807,N_4463,N_3693);
and U5808 (N_5808,N_836,N_4173);
xnor U5809 (N_5809,N_3963,N_4564);
nor U5810 (N_5810,N_4025,N_4091);
or U5811 (N_5811,N_2384,N_2449);
nand U5812 (N_5812,N_21,N_427);
and U5813 (N_5813,N_489,N_4682);
or U5814 (N_5814,N_518,N_211);
nand U5815 (N_5815,N_2019,N_3284);
or U5816 (N_5816,N_2361,N_1600);
and U5817 (N_5817,N_1618,N_2462);
and U5818 (N_5818,N_4035,N_1763);
nand U5819 (N_5819,N_4754,N_1222);
and U5820 (N_5820,N_2468,N_4718);
and U5821 (N_5821,N_3488,N_4255);
nand U5822 (N_5822,N_2510,N_260);
or U5823 (N_5823,N_3673,N_3209);
nor U5824 (N_5824,N_4834,N_455);
nor U5825 (N_5825,N_4743,N_1894);
and U5826 (N_5826,N_3275,N_4051);
and U5827 (N_5827,N_913,N_727);
or U5828 (N_5828,N_959,N_2134);
and U5829 (N_5829,N_3377,N_4259);
nand U5830 (N_5830,N_1453,N_4572);
and U5831 (N_5831,N_1928,N_3648);
and U5832 (N_5832,N_3700,N_1306);
and U5833 (N_5833,N_4498,N_498);
nor U5834 (N_5834,N_2097,N_1156);
nand U5835 (N_5835,N_1757,N_3570);
or U5836 (N_5836,N_2333,N_2811);
or U5837 (N_5837,N_3747,N_2249);
nor U5838 (N_5838,N_2077,N_4221);
and U5839 (N_5839,N_805,N_881);
xor U5840 (N_5840,N_1578,N_445);
nor U5841 (N_5841,N_4313,N_140);
xor U5842 (N_5842,N_1946,N_4774);
nor U5843 (N_5843,N_3645,N_1207);
nand U5844 (N_5844,N_3515,N_3922);
and U5845 (N_5845,N_1526,N_2473);
or U5846 (N_5846,N_4996,N_1363);
nor U5847 (N_5847,N_2447,N_621);
nor U5848 (N_5848,N_2446,N_3912);
xor U5849 (N_5849,N_1697,N_4686);
or U5850 (N_5850,N_4150,N_1166);
nand U5851 (N_5851,N_1460,N_4732);
nand U5852 (N_5852,N_565,N_1726);
nor U5853 (N_5853,N_1656,N_220);
nor U5854 (N_5854,N_4731,N_4171);
nand U5855 (N_5855,N_2748,N_3368);
or U5856 (N_5856,N_2601,N_256);
or U5857 (N_5857,N_936,N_1834);
and U5858 (N_5858,N_6,N_4817);
or U5859 (N_5859,N_3941,N_99);
and U5860 (N_5860,N_1620,N_3867);
xnor U5861 (N_5861,N_994,N_1150);
and U5862 (N_5862,N_2745,N_3848);
nor U5863 (N_5863,N_1510,N_3898);
nor U5864 (N_5864,N_2437,N_2505);
or U5865 (N_5865,N_32,N_832);
nor U5866 (N_5866,N_3255,N_3881);
xnor U5867 (N_5867,N_2329,N_2846);
nor U5868 (N_5868,N_1545,N_2860);
or U5869 (N_5869,N_508,N_691);
nor U5870 (N_5870,N_2877,N_2843);
and U5871 (N_5871,N_1897,N_894);
and U5872 (N_5872,N_4429,N_4308);
or U5873 (N_5873,N_4497,N_2386);
or U5874 (N_5874,N_1768,N_2403);
nand U5875 (N_5875,N_2138,N_535);
xor U5876 (N_5876,N_2605,N_2395);
or U5877 (N_5877,N_1494,N_2529);
and U5878 (N_5878,N_3715,N_3315);
and U5879 (N_5879,N_2054,N_4179);
nor U5880 (N_5880,N_759,N_3429);
or U5881 (N_5881,N_4435,N_3390);
nand U5882 (N_5882,N_1202,N_768);
nand U5883 (N_5883,N_2685,N_1001);
and U5884 (N_5884,N_460,N_152);
nor U5885 (N_5885,N_654,N_2050);
nand U5886 (N_5886,N_2058,N_3089);
and U5887 (N_5887,N_2948,N_726);
nand U5888 (N_5888,N_1714,N_1927);
xnor U5889 (N_5889,N_3298,N_3752);
xor U5890 (N_5890,N_4844,N_2961);
xor U5891 (N_5891,N_1279,N_1613);
nor U5892 (N_5892,N_1968,N_4649);
nor U5893 (N_5893,N_3951,N_3626);
or U5894 (N_5894,N_3142,N_3872);
and U5895 (N_5895,N_3714,N_552);
or U5896 (N_5896,N_436,N_4419);
nand U5897 (N_5897,N_2735,N_207);
or U5898 (N_5898,N_684,N_3580);
or U5899 (N_5899,N_3637,N_3098);
xnor U5900 (N_5900,N_2892,N_1596);
nor U5901 (N_5901,N_382,N_2621);
nor U5902 (N_5902,N_984,N_4812);
nor U5903 (N_5903,N_4162,N_505);
xor U5904 (N_5904,N_1,N_2222);
nor U5905 (N_5905,N_2992,N_4903);
nand U5906 (N_5906,N_3796,N_3933);
or U5907 (N_5907,N_869,N_4267);
nand U5908 (N_5908,N_4409,N_688);
nor U5909 (N_5909,N_3782,N_1564);
or U5910 (N_5910,N_4929,N_3100);
nand U5911 (N_5911,N_4890,N_2773);
nand U5912 (N_5912,N_2623,N_660);
or U5913 (N_5913,N_3074,N_2562);
nor U5914 (N_5914,N_2257,N_2187);
nand U5915 (N_5915,N_2176,N_1106);
or U5916 (N_5916,N_835,N_208);
or U5917 (N_5917,N_1806,N_4634);
nand U5918 (N_5918,N_4992,N_1401);
nor U5919 (N_5919,N_4400,N_4130);
nor U5920 (N_5920,N_4535,N_980);
or U5921 (N_5921,N_1637,N_2108);
nand U5922 (N_5922,N_841,N_551);
nor U5923 (N_5923,N_3220,N_3506);
nor U5924 (N_5924,N_2369,N_1521);
and U5925 (N_5925,N_2071,N_4575);
xnor U5926 (N_5926,N_4510,N_4953);
nand U5927 (N_5927,N_3839,N_3340);
nand U5928 (N_5928,N_3124,N_3548);
nor U5929 (N_5929,N_1127,N_3350);
and U5930 (N_5930,N_4219,N_3086);
and U5931 (N_5931,N_149,N_4125);
or U5932 (N_5932,N_2304,N_3930);
and U5933 (N_5933,N_1689,N_1161);
nand U5934 (N_5934,N_4003,N_453);
nand U5935 (N_5935,N_2780,N_2709);
and U5936 (N_5936,N_3949,N_3174);
nand U5937 (N_5937,N_3393,N_1205);
nand U5938 (N_5938,N_3597,N_1522);
or U5939 (N_5939,N_575,N_4172);
nand U5940 (N_5940,N_3448,N_1720);
or U5941 (N_5941,N_2066,N_1731);
or U5942 (N_5942,N_1186,N_1257);
nor U5943 (N_5943,N_1004,N_2051);
xor U5944 (N_5944,N_3150,N_4062);
nand U5945 (N_5945,N_521,N_640);
xor U5946 (N_5946,N_1502,N_538);
and U5947 (N_5947,N_3042,N_2470);
and U5948 (N_5948,N_4585,N_3269);
nand U5949 (N_5949,N_2808,N_1693);
and U5950 (N_5950,N_842,N_1760);
nand U5951 (N_5951,N_1567,N_395);
or U5952 (N_5952,N_2109,N_1403);
nor U5953 (N_5953,N_2166,N_1991);
and U5954 (N_5954,N_272,N_4863);
nand U5955 (N_5955,N_4692,N_3461);
nand U5956 (N_5956,N_1896,N_253);
and U5957 (N_5957,N_2836,N_73);
nor U5958 (N_5958,N_3555,N_2006);
nor U5959 (N_5959,N_4044,N_3594);
and U5960 (N_5960,N_4005,N_4697);
nor U5961 (N_5961,N_3719,N_3957);
and U5962 (N_5962,N_1540,N_1109);
nand U5963 (N_5963,N_4716,N_2581);
or U5964 (N_5964,N_4925,N_468);
nand U5965 (N_5965,N_4105,N_3382);
nand U5966 (N_5966,N_3641,N_4628);
and U5967 (N_5967,N_1558,N_2564);
and U5968 (N_5968,N_985,N_4430);
nor U5969 (N_5969,N_3102,N_2503);
and U5970 (N_5970,N_594,N_4670);
xor U5971 (N_5971,N_831,N_2644);
nor U5972 (N_5972,N_3035,N_2862);
or U5973 (N_5973,N_1816,N_3466);
nand U5974 (N_5974,N_3870,N_3801);
or U5975 (N_5975,N_4128,N_617);
nand U5976 (N_5976,N_3696,N_3823);
xor U5977 (N_5977,N_4615,N_2416);
and U5978 (N_5978,N_742,N_4740);
nor U5979 (N_5979,N_4877,N_1178);
nand U5980 (N_5980,N_4715,N_4075);
nand U5981 (N_5981,N_3608,N_2229);
nor U5982 (N_5982,N_174,N_2740);
nor U5983 (N_5983,N_3550,N_1655);
xnor U5984 (N_5984,N_463,N_1062);
or U5985 (N_5985,N_2717,N_1965);
nand U5986 (N_5986,N_3216,N_2994);
nor U5987 (N_5987,N_643,N_4509);
nor U5988 (N_5988,N_771,N_4714);
nor U5989 (N_5989,N_2871,N_1468);
nand U5990 (N_5990,N_4525,N_3319);
and U5991 (N_5991,N_2183,N_1049);
nor U5992 (N_5992,N_4040,N_133);
nor U5993 (N_5993,N_4353,N_3367);
and U5994 (N_5994,N_3660,N_2182);
nor U5995 (N_5995,N_1886,N_3780);
or U5996 (N_5996,N_3663,N_2273);
xnor U5997 (N_5997,N_2265,N_4071);
xor U5998 (N_5998,N_3052,N_2859);
or U5999 (N_5999,N_3994,N_2312);
or U6000 (N_6000,N_3915,N_171);
nand U6001 (N_6001,N_4087,N_930);
nor U6002 (N_6002,N_709,N_2667);
or U6003 (N_6003,N_2266,N_3807);
nand U6004 (N_6004,N_1822,N_3835);
xnor U6005 (N_6005,N_473,N_4045);
or U6006 (N_6006,N_3940,N_4336);
or U6007 (N_6007,N_3928,N_4748);
nand U6008 (N_6008,N_1455,N_494);
nand U6009 (N_6009,N_2171,N_2825);
or U6010 (N_6010,N_1962,N_4793);
xnor U6011 (N_6011,N_2786,N_2504);
or U6012 (N_6012,N_78,N_4110);
and U6013 (N_6013,N_903,N_550);
nand U6014 (N_6014,N_584,N_349);
nor U6015 (N_6015,N_3168,N_3576);
or U6016 (N_6016,N_4046,N_2408);
nor U6017 (N_6017,N_4223,N_1091);
and U6018 (N_6018,N_4281,N_69);
nand U6019 (N_6019,N_4292,N_2612);
nor U6020 (N_6020,N_4515,N_4783);
or U6021 (N_6021,N_4617,N_3620);
nor U6022 (N_6022,N_501,N_1182);
xnor U6023 (N_6023,N_2530,N_3088);
and U6024 (N_6024,N_1014,N_3736);
nand U6025 (N_6025,N_246,N_37);
nand U6026 (N_6026,N_2173,N_298);
nor U6027 (N_6027,N_2925,N_2671);
or U6028 (N_6028,N_452,N_919);
or U6029 (N_6029,N_1076,N_4756);
and U6030 (N_6030,N_1352,N_4855);
nand U6031 (N_6031,N_4158,N_2742);
nand U6032 (N_6032,N_3304,N_1862);
nand U6033 (N_6033,N_47,N_3342);
nand U6034 (N_6034,N_2125,N_2847);
and U6035 (N_6035,N_3909,N_2884);
nand U6036 (N_6036,N_3428,N_4526);
nor U6037 (N_6037,N_1256,N_2208);
or U6038 (N_6038,N_3140,N_2003);
and U6039 (N_6039,N_106,N_2908);
and U6040 (N_6040,N_666,N_3838);
or U6041 (N_6041,N_1811,N_3170);
nor U6042 (N_6042,N_799,N_2747);
xor U6043 (N_6043,N_2461,N_3510);
nand U6044 (N_6044,N_4293,N_4168);
or U6045 (N_6045,N_509,N_3529);
xnor U6046 (N_6046,N_3462,N_1418);
or U6047 (N_6047,N_3078,N_2142);
and U6048 (N_6048,N_344,N_4305);
nand U6049 (N_6049,N_1863,N_4316);
or U6050 (N_6050,N_2813,N_1145);
and U6051 (N_6051,N_1899,N_2203);
nor U6052 (N_6052,N_1198,N_4563);
and U6053 (N_6053,N_2281,N_4142);
or U6054 (N_6054,N_312,N_4678);
and U6055 (N_6055,N_858,N_963);
and U6056 (N_6056,N_267,N_1434);
nor U6057 (N_6057,N_534,N_4959);
or U6058 (N_6058,N_176,N_1542);
or U6059 (N_6059,N_765,N_854);
xnor U6060 (N_6060,N_1199,N_3039);
nand U6061 (N_6061,N_4832,N_3161);
nor U6062 (N_6062,N_1662,N_2221);
nand U6063 (N_6063,N_3473,N_918);
or U6064 (N_6064,N_1995,N_3264);
nor U6065 (N_6065,N_4262,N_4674);
and U6066 (N_6066,N_1848,N_1101);
nor U6067 (N_6067,N_2069,N_159);
and U6068 (N_6068,N_658,N_2357);
and U6069 (N_6069,N_200,N_752);
or U6070 (N_6070,N_4547,N_3431);
nor U6071 (N_6071,N_4694,N_3225);
nand U6072 (N_6072,N_488,N_3842);
nand U6073 (N_6073,N_252,N_3381);
nand U6074 (N_6074,N_804,N_2278);
or U6075 (N_6075,N_2291,N_3493);
and U6076 (N_6076,N_4949,N_590);
and U6077 (N_6077,N_3561,N_4629);
or U6078 (N_6078,N_1459,N_634);
nand U6079 (N_6079,N_3636,N_1387);
and U6080 (N_6080,N_1627,N_356);
nor U6081 (N_6081,N_1165,N_4149);
or U6082 (N_6082,N_3690,N_3372);
nor U6083 (N_6083,N_4751,N_690);
nand U6084 (N_6084,N_90,N_1786);
and U6085 (N_6085,N_2729,N_2316);
or U6086 (N_6086,N_3577,N_2286);
or U6087 (N_6087,N_330,N_3273);
nand U6088 (N_6088,N_3337,N_4914);
nand U6089 (N_6089,N_2692,N_3147);
xor U6090 (N_6090,N_758,N_2038);
or U6091 (N_6091,N_1913,N_721);
nor U6092 (N_6092,N_3531,N_1817);
nand U6093 (N_6093,N_1424,N_96);
and U6094 (N_6094,N_3021,N_492);
xor U6095 (N_6095,N_897,N_922);
nand U6096 (N_6096,N_3938,N_1998);
and U6097 (N_6097,N_3889,N_87);
or U6098 (N_6098,N_770,N_1700);
nor U6099 (N_6099,N_4413,N_1984);
nand U6100 (N_6100,N_1042,N_1602);
nand U6101 (N_6101,N_1275,N_4982);
nand U6102 (N_6102,N_1398,N_2792);
nor U6103 (N_6103,N_4352,N_2322);
or U6104 (N_6104,N_952,N_4554);
and U6105 (N_6105,N_2820,N_2609);
xnor U6106 (N_6106,N_1341,N_1298);
nor U6107 (N_6107,N_182,N_338);
nor U6108 (N_6108,N_531,N_3407);
and U6109 (N_6109,N_83,N_2661);
xor U6110 (N_6110,N_435,N_204);
or U6111 (N_6111,N_2370,N_4328);
nand U6112 (N_6112,N_2064,N_3053);
nor U6113 (N_6113,N_4354,N_2444);
nand U6114 (N_6114,N_662,N_1857);
nor U6115 (N_6115,N_628,N_3803);
or U6116 (N_6116,N_4086,N_987);
nand U6117 (N_6117,N_2457,N_399);
xor U6118 (N_6118,N_4038,N_904);
and U6119 (N_6119,N_1331,N_2244);
xor U6120 (N_6120,N_1120,N_89);
or U6121 (N_6121,N_3329,N_2112);
or U6122 (N_6122,N_2480,N_507);
nor U6123 (N_6123,N_3787,N_2508);
or U6124 (N_6124,N_1119,N_3856);
nor U6125 (N_6125,N_292,N_3080);
nand U6126 (N_6126,N_2181,N_2499);
xnor U6127 (N_6127,N_1092,N_1019);
or U6128 (N_6128,N_4764,N_2574);
and U6129 (N_6129,N_715,N_4956);
nand U6130 (N_6130,N_2874,N_1068);
nand U6131 (N_6131,N_107,N_3633);
and U6132 (N_6132,N_3257,N_4976);
and U6133 (N_6133,N_2336,N_2310);
or U6134 (N_6134,N_1730,N_1930);
nor U6135 (N_6135,N_2314,N_2514);
or U6136 (N_6136,N_3980,N_4511);
and U6137 (N_6137,N_2536,N_3291);
nor U6138 (N_6138,N_1905,N_1990);
xor U6139 (N_6139,N_515,N_917);
nor U6140 (N_6140,N_4387,N_3332);
or U6141 (N_6141,N_451,N_3897);
nand U6142 (N_6142,N_4989,N_2835);
nand U6143 (N_6143,N_1259,N_1607);
and U6144 (N_6144,N_2245,N_4960);
and U6145 (N_6145,N_3237,N_2052);
and U6146 (N_6146,N_1497,N_4364);
nor U6147 (N_6147,N_3101,N_2633);
nand U6148 (N_6148,N_3604,N_3552);
nand U6149 (N_6149,N_2371,N_2914);
xor U6150 (N_6150,N_4845,N_2971);
and U6151 (N_6151,N_4339,N_3563);
nor U6152 (N_6152,N_2448,N_1792);
xor U6153 (N_6153,N_701,N_3624);
or U6154 (N_6154,N_3718,N_4236);
nor U6155 (N_6155,N_2065,N_3476);
nor U6156 (N_6156,N_2904,N_1419);
and U6157 (N_6157,N_4636,N_350);
and U6158 (N_6158,N_3355,N_502);
and U6159 (N_6159,N_3,N_2400);
nand U6160 (N_6160,N_2223,N_3223);
nand U6161 (N_6161,N_2338,N_1215);
nor U6162 (N_6162,N_2285,N_2658);
nor U6163 (N_6163,N_2085,N_2389);
and U6164 (N_6164,N_4414,N_2553);
xor U6165 (N_6165,N_407,N_2520);
or U6166 (N_6166,N_1159,N_2781);
nor U6167 (N_6167,N_3199,N_782);
or U6168 (N_6168,N_3425,N_3468);
or U6169 (N_6169,N_111,N_1566);
or U6170 (N_6170,N_683,N_4073);
or U6171 (N_6171,N_873,N_3422);
nand U6172 (N_6172,N_4712,N_3726);
and U6173 (N_6173,N_190,N_3575);
nor U6174 (N_6174,N_3152,N_1438);
or U6175 (N_6175,N_3954,N_566);
nand U6176 (N_6176,N_3154,N_2641);
nand U6177 (N_6177,N_3943,N_3126);
nand U6178 (N_6178,N_3976,N_795);
or U6179 (N_6179,N_4846,N_737);
xnor U6180 (N_6180,N_4402,N_4115);
nor U6181 (N_6181,N_4746,N_4730);
nor U6182 (N_6182,N_233,N_1307);
and U6183 (N_6183,N_3725,N_1873);
nor U6184 (N_6184,N_644,N_1318);
nand U6185 (N_6185,N_4184,N_555);
or U6186 (N_6186,N_1996,N_2712);
nor U6187 (N_6187,N_1135,N_3706);
and U6188 (N_6188,N_2121,N_3944);
nand U6189 (N_6189,N_4443,N_402);
nand U6190 (N_6190,N_2167,N_774);
nand U6191 (N_6191,N_1923,N_1310);
nand U6192 (N_6192,N_4767,N_2741);
and U6193 (N_6193,N_3584,N_2);
or U6194 (N_6194,N_1110,N_3364);
and U6195 (N_6195,N_4578,N_2103);
and U6196 (N_6196,N_4403,N_2831);
nor U6197 (N_6197,N_4448,N_1475);
nor U6198 (N_6198,N_4273,N_3526);
or U6199 (N_6199,N_4013,N_496);
and U6200 (N_6200,N_4668,N_3413);
nor U6201 (N_6201,N_2018,N_4444);
and U6202 (N_6202,N_4894,N_3376);
or U6203 (N_6203,N_2647,N_591);
nand U6204 (N_6204,N_3024,N_1845);
nand U6205 (N_6205,N_4139,N_2652);
and U6206 (N_6206,N_4469,N_753);
nor U6207 (N_6207,N_2650,N_4126);
and U6208 (N_6208,N_1065,N_3612);
nor U6209 (N_6209,N_2133,N_142);
nor U6210 (N_6210,N_4622,N_388);
nand U6211 (N_6211,N_2756,N_3130);
nand U6212 (N_6212,N_2873,N_1698);
nor U6213 (N_6213,N_3036,N_3990);
or U6214 (N_6214,N_1262,N_571);
and U6215 (N_6215,N_2034,N_3439);
or U6216 (N_6216,N_944,N_4612);
nor U6217 (N_6217,N_2498,N_3201);
or U6218 (N_6218,N_2412,N_4445);
nor U6219 (N_6219,N_3862,N_3136);
nand U6220 (N_6220,N_4872,N_2854);
and U6221 (N_6221,N_1537,N_1325);
nor U6222 (N_6222,N_495,N_2193);
and U6223 (N_6223,N_610,N_4602);
and U6224 (N_6224,N_1875,N_4489);
nor U6225 (N_6225,N_4587,N_2515);
nand U6226 (N_6226,N_3635,N_1940);
and U6227 (N_6227,N_2119,N_907);
or U6228 (N_6228,N_2096,N_4112);
nand U6229 (N_6229,N_1330,N_127);
and U6230 (N_6230,N_4464,N_3735);
xor U6231 (N_6231,N_2506,N_3704);
nor U6232 (N_6232,N_4592,N_74);
or U6233 (N_6233,N_4436,N_291);
nor U6234 (N_6234,N_154,N_2464);
or U6235 (N_6235,N_3092,N_4638);
and U6236 (N_6236,N_2500,N_4190);
and U6237 (N_6237,N_3186,N_2812);
xor U6238 (N_6238,N_278,N_1949);
nor U6239 (N_6239,N_920,N_2999);
nor U6240 (N_6240,N_4566,N_1133);
or U6241 (N_6241,N_4163,N_2406);
nor U6242 (N_6242,N_3844,N_2739);
and U6243 (N_6243,N_4735,N_3472);
nor U6244 (N_6244,N_1448,N_3369);
and U6245 (N_6245,N_4186,N_4908);
nor U6246 (N_6246,N_738,N_3171);
and U6247 (N_6247,N_2207,N_3535);
and U6248 (N_6248,N_4570,N_2276);
nor U6249 (N_6249,N_2344,N_139);
nor U6250 (N_6250,N_481,N_4521);
nor U6251 (N_6251,N_2040,N_477);
and U6252 (N_6252,N_4513,N_1659);
or U6253 (N_6253,N_2256,N_4064);
nand U6254 (N_6254,N_2483,N_4332);
nor U6255 (N_6255,N_3831,N_696);
and U6256 (N_6256,N_1175,N_4560);
and U6257 (N_6257,N_2942,N_4084);
xor U6258 (N_6258,N_3817,N_2631);
nor U6259 (N_6259,N_40,N_979);
and U6260 (N_6260,N_2865,N_131);
nor U6261 (N_6261,N_2184,N_4081);
and U6262 (N_6262,N_3006,N_2147);
nand U6263 (N_6263,N_3287,N_357);
nor U6264 (N_6264,N_281,N_4326);
or U6265 (N_6265,N_2242,N_1750);
or U6266 (N_6266,N_4290,N_915);
nor U6267 (N_6267,N_1647,N_4969);
xnor U6268 (N_6268,N_1324,N_784);
nand U6269 (N_6269,N_3187,N_1971);
nor U6270 (N_6270,N_265,N_2118);
nand U6271 (N_6271,N_1346,N_4503);
and U6272 (N_6272,N_484,N_2662);
and U6273 (N_6273,N_1096,N_1926);
and U6274 (N_6274,N_3876,N_4033);
and U6275 (N_6275,N_637,N_2042);
nor U6276 (N_6276,N_3689,N_36);
xnor U6277 (N_6277,N_4002,N_1338);
or U6278 (N_6278,N_1895,N_2721);
or U6279 (N_6279,N_2958,N_3471);
nand U6280 (N_6280,N_2137,N_2837);
or U6281 (N_6281,N_1554,N_2123);
nor U6282 (N_6282,N_1761,N_975);
nor U6283 (N_6283,N_3670,N_957);
and U6284 (N_6284,N_3252,N_4627);
nand U6285 (N_6285,N_4505,N_1033);
or U6286 (N_6286,N_196,N_4902);
nor U6287 (N_6287,N_3877,N_4934);
and U6288 (N_6288,N_1901,N_720);
and U6289 (N_6289,N_2080,N_3979);
nand U6290 (N_6290,N_3458,N_3668);
xor U6291 (N_6291,N_3320,N_45);
xor U6292 (N_6292,N_3855,N_953);
and U6293 (N_6293,N_526,N_882);
and U6294 (N_6294,N_1465,N_3684);
and U6295 (N_6295,N_422,N_4410);
and U6296 (N_6296,N_4815,N_4922);
nand U6297 (N_6297,N_4800,N_1947);
nand U6298 (N_6298,N_305,N_4118);
nand U6299 (N_6299,N_4229,N_3618);
nor U6300 (N_6300,N_2975,N_1414);
and U6301 (N_6301,N_3767,N_3574);
nand U6302 (N_6302,N_4519,N_1880);
or U6303 (N_6303,N_636,N_333);
nor U6304 (N_6304,N_3721,N_2067);
nor U6305 (N_6305,N_1254,N_1775);
nand U6306 (N_6306,N_2951,N_1283);
nor U6307 (N_6307,N_354,N_3541);
or U6308 (N_6308,N_1553,N_92);
nor U6309 (N_6309,N_4495,N_4468);
nand U6310 (N_6310,N_3278,N_1225);
nor U6311 (N_6311,N_2698,N_409);
or U6312 (N_6312,N_3069,N_3785);
or U6313 (N_6313,N_814,N_2152);
or U6314 (N_6314,N_2680,N_1796);
or U6315 (N_6315,N_4181,N_1852);
nand U6316 (N_6316,N_909,N_622);
or U6317 (N_6317,N_2653,N_4446);
nand U6318 (N_6318,N_4415,N_3233);
or U6319 (N_6319,N_2970,N_1123);
or U6320 (N_6320,N_2451,N_1000);
nor U6321 (N_6321,N_1421,N_767);
and U6322 (N_6322,N_392,N_3859);
or U6323 (N_6323,N_748,N_659);
or U6324 (N_6324,N_4202,N_1116);
nor U6325 (N_6325,N_85,N_178);
nor U6326 (N_6326,N_3955,N_3834);
nand U6327 (N_6327,N_1300,N_2851);
and U6328 (N_6328,N_2571,N_3727);
nor U6329 (N_6329,N_3014,N_1974);
nand U6330 (N_6330,N_2707,N_3851);
and U6331 (N_6331,N_1234,N_4476);
nor U6332 (N_6332,N_3583,N_1173);
nand U6333 (N_6333,N_4241,N_1311);
nor U6334 (N_6334,N_3276,N_1934);
nand U6335 (N_6335,N_3111,N_4589);
xnor U6336 (N_6336,N_1456,N_2910);
nor U6337 (N_6337,N_548,N_102);
nand U6338 (N_6338,N_1516,N_3824);
nor U6339 (N_6339,N_1584,N_3799);
nor U6340 (N_6340,N_1467,N_3379);
or U6341 (N_6341,N_2485,N_4277);
xor U6342 (N_6342,N_1285,N_1376);
or U6343 (N_6343,N_3921,N_625);
nor U6344 (N_6344,N_4030,N_4048);
nand U6345 (N_6345,N_4889,N_257);
nor U6346 (N_6346,N_847,N_3026);
and U6347 (N_6347,N_1932,N_1034);
and U6348 (N_6348,N_2382,N_1160);
or U6349 (N_6349,N_3353,N_729);
and U6350 (N_6350,N_1052,N_1556);
nand U6351 (N_6351,N_2777,N_2492);
xnor U6352 (N_6352,N_1721,N_180);
nand U6353 (N_6353,N_2331,N_2243);
nand U6354 (N_6354,N_3456,N_161);
and U6355 (N_6355,N_3863,N_675);
nand U6356 (N_6356,N_1858,N_1488);
or U6357 (N_6357,N_704,N_1051);
or U6358 (N_6358,N_2321,N_1966);
nand U6359 (N_6359,N_2177,N_1660);
or U6360 (N_6360,N_4550,N_4533);
or U6361 (N_6361,N_4355,N_510);
nand U6362 (N_6362,N_86,N_4544);
nor U6363 (N_6363,N_3025,N_4920);
and U6364 (N_6364,N_4912,N_2906);
xnor U6365 (N_6365,N_2710,N_351);
nor U6366 (N_6366,N_404,N_4785);
nand U6367 (N_6367,N_635,N_250);
nand U6368 (N_6368,N_2459,N_1185);
nand U6369 (N_6369,N_3423,N_1684);
nand U6370 (N_6370,N_2049,N_4979);
nor U6371 (N_6371,N_733,N_4717);
xor U6372 (N_6372,N_1609,N_2614);
nand U6373 (N_6373,N_4843,N_3699);
nor U6374 (N_6374,N_2417,N_417);
nand U6375 (N_6375,N_3720,N_2758);
or U6376 (N_6376,N_4738,N_3180);
xor U6377 (N_6377,N_3649,N_935);
or U6378 (N_6378,N_1993,N_3048);
nand U6379 (N_6379,N_4801,N_921);
xnor U6380 (N_6380,N_997,N_1429);
or U6381 (N_6381,N_1478,N_4472);
or U6382 (N_6382,N_2502,N_2630);
or U6383 (N_6383,N_3226,N_3631);
xnor U6384 (N_6384,N_2795,N_3528);
nand U6385 (N_6385,N_3427,N_581);
nand U6386 (N_6386,N_394,N_2161);
nor U6387 (N_6387,N_2102,N_558);
or U6388 (N_6388,N_4508,N_3734);
and U6389 (N_6389,N_1107,N_4050);
nor U6390 (N_6390,N_3522,N_2912);
nor U6391 (N_6391,N_1388,N_3112);
nand U6392 (N_6392,N_3981,N_3892);
and U6393 (N_6393,N_2415,N_4916);
and U6394 (N_6394,N_3370,N_2887);
or U6395 (N_6395,N_3756,N_2132);
and U6396 (N_6396,N_3013,N_3348);
nor U6397 (N_6397,N_1958,N_1216);
or U6398 (N_6398,N_1921,N_1008);
and U6399 (N_6399,N_397,N_4079);
and U6400 (N_6400,N_4211,N_3926);
nor U6401 (N_6401,N_3878,N_239);
or U6402 (N_6402,N_3923,N_3066);
xor U6403 (N_6403,N_4831,N_499);
nor U6404 (N_6404,N_4404,N_1395);
nor U6405 (N_6405,N_1856,N_2720);
and U6406 (N_6406,N_2106,N_2409);
or U6407 (N_6407,N_4407,N_2513);
or U6408 (N_6408,N_4302,N_3864);
xnor U6409 (N_6409,N_2849,N_2407);
and U6410 (N_6410,N_2082,N_3207);
nand U6411 (N_6411,N_3986,N_2280);
nor U6412 (N_6412,N_4151,N_4621);
nor U6413 (N_6413,N_4779,N_4787);
and U6414 (N_6414,N_1898,N_2236);
or U6415 (N_6415,N_4679,N_4250);
xnor U6416 (N_6416,N_1409,N_4913);
xor U6417 (N_6417,N_3858,N_3743);
nor U6418 (N_6418,N_3935,N_1649);
or U6419 (N_6419,N_587,N_2830);
or U6420 (N_6420,N_1703,N_166);
nand U6421 (N_6421,N_1476,N_567);
nand U6422 (N_6422,N_469,N_1869);
nor U6423 (N_6423,N_381,N_1679);
nor U6424 (N_6424,N_1174,N_2645);
nand U6425 (N_6425,N_3530,N_4775);
and U6426 (N_6426,N_1673,N_3490);
and U6427 (N_6427,N_4143,N_4899);
or U6428 (N_6428,N_615,N_1512);
xnor U6429 (N_6429,N_101,N_1821);
and U6430 (N_6430,N_2477,N_4388);
nor U6431 (N_6431,N_124,N_347);
xor U6432 (N_6432,N_3312,N_3253);
or U6433 (N_6433,N_1277,N_4335);
and U6434 (N_6434,N_1060,N_2967);
or U6435 (N_6435,N_3239,N_3775);
nand U6436 (N_6436,N_3469,N_1539);
and U6437 (N_6437,N_3543,N_4254);
and U6438 (N_6438,N_3343,N_2933);
nand U6439 (N_6439,N_4971,N_1524);
and U6440 (N_6440,N_3755,N_1843);
and U6441 (N_6441,N_3978,N_1292);
nor U6442 (N_6442,N_1580,N_3962);
nor U6443 (N_6443,N_4773,N_2665);
or U6444 (N_6444,N_1964,N_3952);
nor U6445 (N_6445,N_3292,N_857);
nand U6446 (N_6446,N_1734,N_1527);
or U6447 (N_6447,N_1309,N_772);
nor U6448 (N_6448,N_2129,N_1685);
nor U6449 (N_6449,N_3874,N_4320);
nor U6450 (N_6450,N_524,N_2214);
and U6451 (N_6451,N_1335,N_940);
and U6452 (N_6452,N_3323,N_1231);
nand U6453 (N_6453,N_4076,N_1389);
nor U6454 (N_6454,N_3309,N_4811);
or U6455 (N_6455,N_4652,N_3412);
and U6456 (N_6456,N_2192,N_4927);
nand U6457 (N_6457,N_192,N_4907);
or U6458 (N_6458,N_1301,N_403);
nor U6459 (N_6459,N_2362,N_2974);
nor U6460 (N_6460,N_183,N_1015);
or U6461 (N_6461,N_3204,N_2185);
and U6462 (N_6462,N_998,N_5);
and U6463 (N_6463,N_2140,N_1622);
xnor U6464 (N_6464,N_2455,N_4527);
or U6465 (N_6465,N_665,N_2139);
and U6466 (N_6466,N_678,N_206);
and U6467 (N_6467,N_3728,N_3121);
or U6468 (N_6468,N_348,N_1093);
nor U6469 (N_6469,N_1911,N_4607);
nand U6470 (N_6470,N_1953,N_4203);
or U6471 (N_6471,N_3804,N_2294);
and U6472 (N_6472,N_3016,N_332);
or U6473 (N_6473,N_2007,N_4681);
xnor U6474 (N_6474,N_1013,N_2583);
nand U6475 (N_6475,N_801,N_2639);
xor U6476 (N_6476,N_1769,N_570);
or U6477 (N_6477,N_3133,N_177);
nor U6478 (N_6478,N_3334,N_4741);
and U6479 (N_6479,N_1807,N_3279);
and U6480 (N_6480,N_1840,N_2527);
or U6481 (N_6481,N_189,N_2844);
and U6482 (N_6482,N_1345,N_1804);
and U6483 (N_6483,N_3143,N_2383);
nand U6484 (N_6484,N_1407,N_520);
xnor U6485 (N_6485,N_1323,N_3167);
or U6486 (N_6486,N_938,N_1674);
nand U6487 (N_6487,N_3671,N_3045);
nor U6488 (N_6488,N_2198,N_1626);
or U6489 (N_6489,N_826,N_927);
and U6490 (N_6490,N_3989,N_4823);
nor U6491 (N_6491,N_7,N_2135);
nor U6492 (N_6492,N_4641,N_1340);
or U6493 (N_6493,N_4601,N_4940);
nor U6494 (N_6494,N_4421,N_4576);
nand U6495 (N_6495,N_1454,N_4425);
and U6496 (N_6496,N_865,N_3218);
or U6497 (N_6497,N_2428,N_3235);
nor U6498 (N_6498,N_385,N_2479);
xnor U6499 (N_6499,N_1099,N_4416);
nand U6500 (N_6500,N_4189,N_934);
nand U6501 (N_6501,N_1336,N_1737);
and U6502 (N_6502,N_4873,N_3999);
nor U6503 (N_6503,N_456,N_1058);
and U6504 (N_6504,N_1859,N_4159);
xor U6505 (N_6505,N_4456,N_2711);
nor U6506 (N_6506,N_2272,N_3023);
nor U6507 (N_6507,N_1866,N_4768);
xnor U6508 (N_6508,N_1420,N_426);
nand U6509 (N_6509,N_2695,N_989);
nand U6510 (N_6510,N_4478,N_3883);
xnor U6511 (N_6511,N_3051,N_4867);
nor U6512 (N_6512,N_652,N_4541);
and U6513 (N_6513,N_4070,N_4106);
and U6514 (N_6514,N_4635,N_430);
xor U6515 (N_6515,N_3380,N_4037);
nor U6516 (N_6516,N_877,N_4377);
xnor U6517 (N_6517,N_2035,N_4188);
nand U6518 (N_6518,N_450,N_3481);
and U6519 (N_6519,N_3075,N_2332);
nor U6520 (N_6520,N_645,N_3033);
nor U6521 (N_6521,N_2231,N_2004);
nor U6522 (N_6522,N_4225,N_1975);
and U6523 (N_6523,N_234,N_4129);
nand U6524 (N_6524,N_2517,N_4884);
and U6525 (N_6525,N_977,N_1315);
nand U6526 (N_6526,N_380,N_1533);
and U6527 (N_6527,N_26,N_4340);
nand U6528 (N_6528,N_2608,N_479);
or U6529 (N_6529,N_4194,N_4600);
or U6530 (N_6530,N_1710,N_4707);
or U6531 (N_6531,N_4175,N_853);
or U6532 (N_6532,N_981,N_3059);
nor U6533 (N_6533,N_852,N_4516);
and U6534 (N_6534,N_1903,N_474);
or U6535 (N_6535,N_1196,N_898);
xnor U6536 (N_6536,N_2029,N_1079);
nand U6537 (N_6537,N_2460,N_2803);
or U6538 (N_6538,N_1252,N_2806);
and U6539 (N_6539,N_3302,N_1742);
nor U6540 (N_6540,N_2935,N_3603);
nor U6541 (N_6541,N_2145,N_254);
nand U6542 (N_6542,N_1462,N_3820);
and U6543 (N_6543,N_3424,N_905);
and U6544 (N_6544,N_65,N_3680);
or U6545 (N_6545,N_4941,N_3908);
nor U6546 (N_6546,N_3139,N_3333);
nand U6547 (N_6547,N_4514,N_4122);
nor U6548 (N_6548,N_4910,N_1779);
or U6549 (N_6549,N_2351,N_1073);
or U6550 (N_6550,N_119,N_862);
nand U6551 (N_6551,N_2328,N_4109);
or U6552 (N_6552,N_1355,N_4054);
and U6553 (N_6553,N_1125,N_3788);
or U6554 (N_6554,N_3234,N_3389);
or U6555 (N_6555,N_4932,N_3517);
and U6556 (N_6556,N_851,N_2968);
xor U6557 (N_6557,N_775,N_4032);
nand U6558 (N_6558,N_446,N_4561);
or U6559 (N_6559,N_2845,N_2659);
or U6560 (N_6560,N_2324,N_3383);
or U6561 (N_6561,N_3610,N_2287);
and U6562 (N_6562,N_1187,N_3644);
nor U6563 (N_6563,N_2558,N_4294);
nand U6564 (N_6564,N_1652,N_3206);
and U6565 (N_6565,N_2349,N_560);
and U6566 (N_6566,N_1950,N_2037);
or U6567 (N_6567,N_3451,N_318);
nand U6568 (N_6568,N_46,N_3295);
xor U6569 (N_6569,N_4593,N_4296);
nor U6570 (N_6570,N_2690,N_117);
nor U6571 (N_6571,N_1765,N_4069);
nand U6572 (N_6572,N_681,N_4688);
or U6573 (N_6573,N_1406,N_2374);
and U6574 (N_6574,N_1529,N_150);
or U6575 (N_6575,N_2122,N_3067);
nor U6576 (N_6576,N_138,N_3832);
nand U6577 (N_6577,N_3843,N_1365);
nor U6578 (N_6578,N_3249,N_577);
nor U6579 (N_6579,N_563,N_1002);
or U6580 (N_6580,N_144,N_3417);
or U6581 (N_6581,N_2872,N_129);
and U6582 (N_6582,N_519,N_3043);
and U6583 (N_6583,N_2092,N_3200);
nand U6584 (N_6584,N_3061,N_4401);
nand U6585 (N_6585,N_3144,N_4147);
nand U6586 (N_6586,N_2545,N_4868);
nor U6587 (N_6587,N_1428,N_3729);
or U6588 (N_6588,N_34,N_1431);
nor U6589 (N_6589,N_2864,N_2917);
nand U6590 (N_6590,N_8,N_2911);
nand U6591 (N_6591,N_674,N_971);
xnor U6592 (N_6592,N_1833,N_3532);
xor U6593 (N_6593,N_1411,N_245);
or U6594 (N_6594,N_1592,N_700);
and U6595 (N_6595,N_1773,N_866);
xnor U6596 (N_6596,N_2832,N_4664);
nand U6597 (N_6597,N_4161,N_2546);
nor U6598 (N_6598,N_3776,N_4518);
xnor U6599 (N_6599,N_12,N_2772);
nor U6600 (N_6600,N_3445,N_4896);
nand U6601 (N_6601,N_2478,N_55);
nand U6602 (N_6602,N_3662,N_1484);
nor U6603 (N_6603,N_588,N_1118);
or U6604 (N_6604,N_1063,N_1782);
nor U6605 (N_6605,N_3261,N_3454);
nor U6606 (N_6606,N_4559,N_1702);
or U6607 (N_6607,N_2151,N_2637);
or U6608 (N_6608,N_4974,N_336);
nor U6609 (N_6609,N_3286,N_2771);
and U6610 (N_6610,N_976,N_2833);
nand U6611 (N_6611,N_14,N_1766);
nand U6612 (N_6612,N_20,N_4334);
or U6613 (N_6613,N_3625,N_4700);
or U6614 (N_6614,N_945,N_3732);
and U6615 (N_6615,N_833,N_4993);
and U6616 (N_6616,N_3131,N_4466);
and U6617 (N_6617,N_1604,N_4228);
and U6618 (N_6618,N_2141,N_3913);
or U6619 (N_6619,N_1707,N_151);
and U6620 (N_6620,N_1089,N_3108);
nand U6621 (N_6621,N_412,N_10);
or U6622 (N_6622,N_1881,N_4440);
or U6623 (N_6623,N_2753,N_2443);
nor U6624 (N_6624,N_1669,N_1168);
xnor U6625 (N_6625,N_4942,N_3160);
or U6626 (N_6626,N_264,N_3571);
nand U6627 (N_6627,N_2613,N_4058);
nor U6628 (N_6628,N_3910,N_1054);
or U6629 (N_6629,N_2725,N_4368);
and U6630 (N_6630,N_716,N_4878);
or U6631 (N_6631,N_1360,N_1709);
nand U6632 (N_6632,N_2886,N_3521);
and U6633 (N_6633,N_2311,N_3321);
or U6634 (N_6634,N_1141,N_950);
and U6635 (N_6635,N_3047,N_3485);
nand U6636 (N_6636,N_4906,N_2091);
nand U6637 (N_6637,N_970,N_134);
nand U6638 (N_6638,N_1143,N_607);
nand U6639 (N_6639,N_3560,N_1028);
nor U6640 (N_6640,N_2643,N_3683);
nand U6641 (N_6641,N_604,N_2731);
nor U6642 (N_6642,N_2853,N_2441);
and U6643 (N_6643,N_673,N_3676);
nand U6644 (N_6644,N_4135,N_1470);
or U6645 (N_6645,N_4943,N_1914);
nor U6646 (N_6646,N_2794,N_3811);
nor U6647 (N_6647,N_3861,N_2898);
or U6648 (N_6648,N_4031,N_2784);
nor U6649 (N_6649,N_1103,N_243);
nor U6650 (N_6650,N_4330,N_1224);
nand U6651 (N_6651,N_4303,N_2472);
or U6652 (N_6652,N_671,N_3359);
nor U6653 (N_6653,N_2297,N_2769);
or U6654 (N_6654,N_3784,N_2990);
and U6655 (N_6655,N_3777,N_4729);
nand U6656 (N_6656,N_1504,N_2947);
nor U6657 (N_6657,N_2751,N_2030);
and U6658 (N_6658,N_1229,N_3151);
nor U6659 (N_6659,N_2002,N_2131);
or U6660 (N_6660,N_3217,N_1906);
xnor U6661 (N_6661,N_4381,N_4018);
or U6662 (N_6662,N_1111,N_1217);
nand U6663 (N_6663,N_38,N_4345);
nand U6664 (N_6664,N_2188,N_225);
or U6665 (N_6665,N_2946,N_2454);
and U6666 (N_6666,N_2907,N_2810);
or U6667 (N_6667,N_24,N_4766);
nor U6668 (N_6668,N_1132,N_3903);
or U6669 (N_6669,N_3669,N_181);
or U6670 (N_6670,N_327,N_4182);
and U6671 (N_6671,N_4152,N_4928);
nor U6672 (N_6672,N_3277,N_2364);
nand U6673 (N_6673,N_2861,N_3362);
or U6674 (N_6674,N_4719,N_1353);
or U6675 (N_6675,N_2660,N_3623);
nand U6676 (N_6676,N_4660,N_1435);
xor U6677 (N_6677,N_649,N_631);
nand U6678 (N_6678,N_3263,N_3096);
or U6679 (N_6679,N_983,N_3596);
or U6680 (N_6680,N_4926,N_1844);
xnor U6681 (N_6681,N_4117,N_1680);
xnor U6682 (N_6682,N_3614,N_1867);
and U6683 (N_6683,N_703,N_4776);
nor U6684 (N_6684,N_122,N_3093);
nor U6685 (N_6685,N_2497,N_943);
nor U6686 (N_6686,N_1358,N_2306);
xor U6687 (N_6687,N_1788,N_2475);
xor U6688 (N_6688,N_4987,N_1153);
nand U6689 (N_6689,N_4437,N_4866);
or U6690 (N_6690,N_1158,N_4701);
nand U6691 (N_6691,N_3852,N_4157);
xnor U6692 (N_6692,N_1535,N_3918);
nor U6693 (N_6693,N_955,N_1261);
and U6694 (N_6694,N_3629,N_2764);
or U6695 (N_6695,N_834,N_3169);
xnor U6696 (N_6696,N_4486,N_1041);
or U6697 (N_6697,N_1632,N_4131);
and U6698 (N_6698,N_2684,N_128);
xnor U6699 (N_6699,N_2672,N_3572);
and U6700 (N_6700,N_4226,N_4967);
nor U6701 (N_6701,N_3934,N_2175);
and U6702 (N_6702,N_1861,N_3640);
xnor U6703 (N_6703,N_1891,N_1251);
nand U6704 (N_6704,N_4137,N_2869);
or U6705 (N_6705,N_2124,N_2204);
and U6706 (N_6706,N_1664,N_1752);
and U6707 (N_6707,N_277,N_2392);
nand U6708 (N_6708,N_2775,N_892);
nor U6709 (N_6709,N_3638,N_3770);
nor U6710 (N_6710,N_172,N_2587);
or U6711 (N_6711,N_2348,N_2728);
and U6712 (N_6712,N_467,N_4306);
nor U6713 (N_6713,N_1944,N_3516);
or U6714 (N_6714,N_2788,N_4888);
and U6715 (N_6715,N_4538,N_1814);
and U6716 (N_6716,N_4558,N_4944);
and U6717 (N_6717,N_3573,N_2952);
xnor U6718 (N_6718,N_4892,N_863);
or U6719 (N_6719,N_1722,N_4199);
nand U6720 (N_6720,N_2290,N_528);
nor U6721 (N_6721,N_596,N_1319);
or U6722 (N_6722,N_844,N_1519);
nor U6723 (N_6723,N_459,N_3678);
nor U6724 (N_6724,N_4252,N_4549);
and U6725 (N_6725,N_421,N_2212);
or U6726 (N_6726,N_2733,N_1756);
and U6727 (N_6727,N_4383,N_573);
nand U6728 (N_6728,N_1641,N_2226);
or U6729 (N_6729,N_1440,N_3953);
and U6730 (N_6730,N_1931,N_1433);
nand U6731 (N_6731,N_3914,N_1999);
and U6732 (N_6732,N_641,N_3386);
or U6733 (N_6733,N_4242,N_3544);
or U6734 (N_6734,N_3011,N_2675);
and U6735 (N_6735,N_2915,N_1333);
or U6736 (N_6736,N_4631,N_4935);
and U6737 (N_6737,N_4243,N_3996);
nand U6738 (N_6738,N_4167,N_3924);
nor U6739 (N_6739,N_1302,N_2424);
and U6740 (N_6740,N_3695,N_4966);
or U6741 (N_6741,N_3677,N_2159);
nor U6742 (N_6742,N_110,N_1482);
and U6743 (N_6743,N_2360,N_734);
nor U6744 (N_6744,N_3438,N_3082);
nand U6745 (N_6745,N_995,N_3190);
xor U6746 (N_6746,N_120,N_4901);
and U6747 (N_6747,N_1571,N_4782);
and U6748 (N_6748,N_580,N_1849);
nor U6749 (N_6749,N_890,N_3254);
and U6750 (N_6750,N_3391,N_2622);
and U6751 (N_6751,N_4584,N_3854);
or U6752 (N_6752,N_4605,N_4282);
and U6753 (N_6753,N_1908,N_511);
and U6754 (N_6754,N_3948,N_3966);
nor U6755 (N_6755,N_3005,N_434);
or U6756 (N_6756,N_4725,N_3070);
nand U6757 (N_6757,N_4972,N_860);
xnor U6758 (N_6758,N_3480,N_2761);
nand U6759 (N_6759,N_3030,N_1040);
or U6760 (N_6760,N_1639,N_2440);
or U6761 (N_6761,N_4418,N_3538);
and U6762 (N_6762,N_2239,N_2528);
nor U6763 (N_6763,N_1784,N_2732);
or U6764 (N_6764,N_3352,N_1509);
or U6765 (N_6765,N_2763,N_789);
nand U6766 (N_6766,N_3533,N_2882);
and U6767 (N_6767,N_1992,N_2857);
and U6768 (N_6768,N_1441,N_2575);
xor U6769 (N_6769,N_4372,N_121);
nand U6770 (N_6770,N_3094,N_4078);
or U6771 (N_6771,N_3884,N_2778);
nand U6772 (N_6772,N_1879,N_4850);
and U6773 (N_6773,N_3786,N_355);
or U6774 (N_6774,N_4307,N_53);
and U6775 (N_6775,N_1113,N_1140);
or U6776 (N_6776,N_1551,N_1829);
or U6777 (N_6777,N_986,N_4579);
or U6778 (N_6778,N_1628,N_4077);
and U6779 (N_6779,N_3992,N_4689);
nand U6780 (N_6780,N_175,N_3378);
or U6781 (N_6781,N_4921,N_3582);
nor U6782 (N_6782,N_4082,N_4911);
or U6783 (N_6783,N_3128,N_4191);
nand U6784 (N_6784,N_2651,N_1785);
nor U6785 (N_6785,N_3232,N_1764);
nand U6786 (N_6786,N_1115,N_4507);
or U6787 (N_6787,N_2573,N_807);
nand U6788 (N_6788,N_4349,N_1147);
nor U6789 (N_6789,N_393,N_1791);
and U6790 (N_6790,N_993,N_408);
nand U6791 (N_6791,N_2588,N_1337);
or U6792 (N_6792,N_3590,N_4869);
xor U6793 (N_6793,N_1130,N_4727);
or U6794 (N_6794,N_4502,N_3974);
nor U6795 (N_6795,N_3675,N_2381);
xnor U6796 (N_6796,N_2079,N_4237);
nor U6797 (N_6797,N_2169,N_1772);
and U6798 (N_6798,N_366,N_3155);
or U6799 (N_6799,N_972,N_1678);
and U6800 (N_6800,N_1367,N_4946);
nand U6801 (N_6801,N_2481,N_217);
nor U6802 (N_6802,N_2955,N_4011);
and U6803 (N_6803,N_2625,N_4008);
nor U6804 (N_6804,N_3285,N_619);
and U6805 (N_6805,N_141,N_1278);
or U6806 (N_6806,N_125,N_4586);
nand U6807 (N_6807,N_546,N_4001);
nor U6808 (N_6808,N_2246,N_1841);
nand U6809 (N_6809,N_3969,N_4802);
and U6810 (N_6810,N_2706,N_209);
and U6811 (N_6811,N_763,N_2296);
and U6812 (N_6812,N_3183,N_605);
or U6813 (N_6813,N_529,N_3498);
and U6814 (N_6814,N_2251,N_2569);
xnor U6815 (N_6815,N_68,N_4565);
or U6816 (N_6816,N_547,N_4083);
nor U6817 (N_6817,N_4373,N_2153);
nor U6818 (N_6818,N_1094,N_757);
and U6819 (N_6819,N_4447,N_2059);
and U6820 (N_6820,N_4004,N_4648);
or U6821 (N_6821,N_3611,N_1629);
nand U6822 (N_6822,N_939,N_4061);
and U6823 (N_6823,N_94,N_2787);
nor U6824 (N_6824,N_4333,N_3079);
or U6825 (N_6825,N_4238,N_3860);
and U6826 (N_6826,N_3917,N_1495);
and U6827 (N_6827,N_1653,N_4543);
nor U6828 (N_6828,N_1206,N_4824);
or U6829 (N_6829,N_633,N_4279);
and U6830 (N_6830,N_1043,N_2941);
nor U6831 (N_6831,N_2926,N_54);
and U6832 (N_6832,N_651,N_2487);
nor U6833 (N_6833,N_1614,N_4295);
xnor U6834 (N_6834,N_2020,N_3345);
and U6835 (N_6835,N_4263,N_802);
or U6836 (N_6836,N_1864,N_4442);
xnor U6837 (N_6837,N_3658,N_3651);
nand U6838 (N_6838,N_2164,N_743);
nand U6839 (N_6839,N_751,N_586);
or U6840 (N_6840,N_2604,N_2730);
nand U6841 (N_6841,N_248,N_4900);
nor U6842 (N_6842,N_4865,N_1888);
nand U6843 (N_6843,N_3188,N_3826);
nor U6844 (N_6844,N_1458,N_4359);
nor U6845 (N_6845,N_3982,N_3189);
xor U6846 (N_6846,N_1920,N_4327);
or U6847 (N_6847,N_2445,N_2160);
nand U6848 (N_6848,N_843,N_1853);
nand U6849 (N_6849,N_3763,N_4164);
nand U6850 (N_6850,N_1576,N_2723);
xnor U6851 (N_6851,N_2073,N_3153);
or U6852 (N_6852,N_1266,N_2867);
or U6853 (N_6853,N_4123,N_1642);
nor U6854 (N_6854,N_1287,N_1348);
nand U6855 (N_6855,N_146,N_297);
and U6856 (N_6856,N_2597,N_2163);
or U6857 (N_6857,N_2524,N_2439);
and U6858 (N_6858,N_4454,N_4113);
xnor U6859 (N_6859,N_4875,N_2298);
or U6860 (N_6860,N_1048,N_4195);
and U6861 (N_6861,N_3483,N_4737);
and U6862 (N_6862,N_2334,N_4160);
xor U6863 (N_6863,N_1087,N_923);
nand U6864 (N_6864,N_2060,N_3426);
or U6865 (N_6865,N_988,N_3741);
and U6866 (N_6866,N_1549,N_1183);
xor U6867 (N_6867,N_1699,N_247);
nor U6868 (N_6868,N_359,N_3414);
and U6869 (N_6869,N_4839,N_4551);
or U6870 (N_6870,N_4672,N_4473);
nand U6871 (N_6871,N_4244,N_4835);
nand U6872 (N_6872,N_3001,N_1711);
nand U6873 (N_6873,N_3330,N_2677);
or U6874 (N_6874,N_4178,N_4758);
or U6875 (N_6875,N_447,N_4016);
and U6876 (N_6876,N_4603,N_1097);
and U6877 (N_6877,N_4289,N_2525);
nor U6878 (N_6878,N_3058,N_2554);
nor U6879 (N_6879,N_4,N_4791);
nand U6880 (N_6880,N_290,N_3809);
nor U6881 (N_6881,N_717,N_4207);
or U6882 (N_6882,N_4528,N_2715);
nor U6883 (N_6883,N_3894,N_3110);
nand U6884 (N_6884,N_1280,N_4348);
xnor U6885 (N_6885,N_536,N_2618);
nand U6886 (N_6886,N_3771,N_1885);
nand U6887 (N_6887,N_902,N_1744);
or U6888 (N_6888,N_3056,N_2033);
nand U6889 (N_6889,N_4312,N_2186);
and U6890 (N_6890,N_2765,N_3717);
nor U6891 (N_6891,N_2682,N_3606);
nand U6892 (N_6892,N_1612,N_3511);
nand U6893 (N_6893,N_2959,N_4977);
nor U6894 (N_6894,N_1370,N_1826);
and U6895 (N_6895,N_362,N_3710);
or U6896 (N_6896,N_4675,N_1447);
nor U6897 (N_6897,N_3519,N_991);
nor U6898 (N_6898,N_2998,N_2678);
xor U6899 (N_6899,N_2197,N_4995);
xor U6900 (N_6900,N_3967,N_3837);
or U6901 (N_6901,N_598,N_4778);
nand U6902 (N_6902,N_4710,N_4534);
nor U6903 (N_6903,N_1463,N_4739);
and U6904 (N_6904,N_2696,N_4218);
nand U6905 (N_6905,N_2534,N_2252);
or U6906 (N_6906,N_4637,N_228);
or U6907 (N_6907,N_2976,N_1220);
or U6908 (N_6908,N_4344,N_1045);
nor U6909 (N_6909,N_820,N_425);
nand U6910 (N_6910,N_2586,N_411);
or U6911 (N_6911,N_3044,N_4963);
nand U6912 (N_6912,N_2549,N_3875);
nand U6913 (N_6913,N_1200,N_113);
and U6914 (N_6914,N_4056,N_2496);
xnor U6915 (N_6915,N_4423,N_2156);
or U6916 (N_6916,N_3977,N_911);
or U6917 (N_6917,N_3540,N_1219);
and U6918 (N_6918,N_523,N_808);
or U6919 (N_6919,N_4258,N_2746);
and U6920 (N_6920,N_4788,N_965);
and U6921 (N_6921,N_2656,N_3985);
xor U6922 (N_6922,N_2023,N_4761);
nor U6923 (N_6923,N_3600,N_2277);
or U6924 (N_6924,N_4923,N_321);
nor U6925 (N_6925,N_4858,N_3296);
nor U6926 (N_6926,N_3687,N_4591);
nor U6927 (N_6927,N_4781,N_706);
xor U6928 (N_6928,N_1122,N_871);
nor U6929 (N_6929,N_195,N_1956);
nand U6930 (N_6930,N_3739,N_1610);
and U6931 (N_6931,N_4571,N_838);
or U6932 (N_6932,N_3310,N_2819);
or U6933 (N_6933,N_2074,N_1874);
nand U6934 (N_6934,N_803,N_4504);
nor U6935 (N_6935,N_3813,N_1381);
xnor U6936 (N_6936,N_3149,N_4483);
and U6937 (N_6937,N_216,N_1573);
nand U6938 (N_6938,N_3885,N_4499);
nor U6939 (N_6939,N_3972,N_787);
nor U6940 (N_6940,N_4449,N_3829);
nor U6941 (N_6941,N_4680,N_3895);
and U6942 (N_6942,N_2555,N_70);
nand U6943 (N_6943,N_1594,N_3195);
nand U6944 (N_6944,N_237,N_3891);
nor U6945 (N_6945,N_792,N_2891);
or U6946 (N_6946,N_3509,N_1112);
or U6947 (N_6947,N_1969,N_2404);
xnor U6948 (N_6948,N_2233,N_840);
or U6949 (N_6949,N_431,N_1889);
xnor U6950 (N_6950,N_2944,N_2953);
and U6951 (N_6951,N_4522,N_1373);
and U6952 (N_6952,N_2194,N_1362);
nor U6953 (N_6953,N_1802,N_1732);
or U6954 (N_6954,N_1012,N_88);
nand U6955 (N_6955,N_2782,N_4759);
nor U6956 (N_6956,N_2809,N_3503);
or U6957 (N_6957,N_3194,N_3403);
xnor U6958 (N_6958,N_4417,N_642);
nand U6959 (N_6959,N_4806,N_4990);
nor U6960 (N_6960,N_4705,N_3795);
and U6961 (N_6961,N_109,N_471);
xor U6962 (N_6962,N_3231,N_1349);
nand U6963 (N_6963,N_114,N_2934);
or U6964 (N_6964,N_2305,N_4166);
and U6965 (N_6965,N_9,N_2402);
nand U6966 (N_6966,N_4609,N_1623);
nand U6967 (N_6967,N_1025,N_1687);
xor U6968 (N_6968,N_4604,N_218);
and U6969 (N_6969,N_3731,N_2180);
nand U6970 (N_6970,N_2570,N_4121);
and U6971 (N_6971,N_2008,N_4854);
nor U6972 (N_6972,N_2628,N_1151);
xor U6973 (N_6973,N_4620,N_514);
nand U6974 (N_6974,N_773,N_2365);
and U6975 (N_6975,N_1503,N_1221);
nand U6976 (N_6976,N_3385,N_1650);
or U6977 (N_6977,N_2165,N_2566);
nand U6978 (N_6978,N_3341,N_1525);
or U6979 (N_6979,N_3224,N_1451);
or U6980 (N_6980,N_4441,N_3589);
nand U6981 (N_6981,N_1854,N_389);
or U6982 (N_6982,N_1860,N_1258);
and U6983 (N_6983,N_4024,N_3020);
and U6984 (N_6984,N_3805,N_202);
nor U6985 (N_6985,N_1380,N_3691);
and U6986 (N_6986,N_1316,N_4119);
or U6987 (N_6987,N_3737,N_1777);
and U6988 (N_6988,N_3557,N_4978);
or U6989 (N_6989,N_1871,N_2453);
nor U6990 (N_6990,N_98,N_4012);
nand U6991 (N_6991,N_2346,N_2047);
xor U6992 (N_6992,N_2624,N_1587);
and U6993 (N_6993,N_337,N_1342);
nand U6994 (N_6994,N_3886,N_4467);
and U6995 (N_6995,N_2649,N_4553);
or U6996 (N_6996,N_1572,N_3484);
xnor U6997 (N_6997,N_2693,N_2580);
nor U6998 (N_6998,N_1326,N_2216);
or U6999 (N_6999,N_3551,N_522);
nor U7000 (N_7000,N_1562,N_3246);
or U7001 (N_7001,N_108,N_4654);
and U7002 (N_7002,N_2858,N_2755);
nor U7003 (N_7003,N_2646,N_2044);
nand U7004 (N_7004,N_384,N_81);
and U7005 (N_7005,N_1317,N_2950);
nand U7006 (N_7006,N_3630,N_3520);
and U7007 (N_7007,N_2474,N_3609);
and U7008 (N_7008,N_4662,N_324);
nand U7009 (N_7009,N_3525,N_870);
or U7010 (N_7010,N_4266,N_2259);
nor U7011 (N_7011,N_3107,N_4829);
xor U7012 (N_7012,N_4623,N_525);
nand U7013 (N_7013,N_2889,N_315);
nand U7014 (N_7014,N_3773,N_4523);
nor U7015 (N_7015,N_4798,N_3000);
and U7016 (N_7016,N_667,N_3808);
xor U7017 (N_7017,N_3371,N_1994);
xnor U7018 (N_7018,N_4809,N_2434);
and U7019 (N_7019,N_1241,N_4703);
nand U7020 (N_7020,N_1393,N_2602);
xor U7021 (N_7021,N_1532,N_1893);
nand U7022 (N_7022,N_3418,N_2736);
or U7023 (N_7023,N_2899,N_2578);
and U7024 (N_7024,N_343,N_1951);
xnor U7025 (N_7025,N_4000,N_2353);
nor U7026 (N_7026,N_3077,N_173);
nand U7027 (N_7027,N_52,N_2683);
and U7028 (N_7028,N_226,N_1177);
xor U7029 (N_7029,N_583,N_2688);
or U7030 (N_7030,N_4180,N_4590);
or U7031 (N_7031,N_1129,N_3553);
nor U7032 (N_7032,N_3961,N_4485);
nor U7033 (N_7033,N_549,N_458);
nand U7034 (N_7034,N_4991,N_4021);
or U7035 (N_7035,N_3685,N_1249);
nor U7036 (N_7036,N_3840,N_3442);
or U7037 (N_7037,N_1136,N_2414);
nor U7038 (N_7038,N_2937,N_2686);
or U7039 (N_7039,N_2372,N_4883);
nand U7040 (N_7040,N_1981,N_2401);
nand U7041 (N_7041,N_346,N_376);
nand U7042 (N_7042,N_2902,N_2531);
and U7043 (N_7043,N_3748,N_946);
or U7044 (N_7044,N_3905,N_2267);
nand U7045 (N_7045,N_3815,N_1450);
nand U7046 (N_7046,N_2762,N_4029);
nor U7047 (N_7047,N_2727,N_3806);
nor U7048 (N_7048,N_340,N_4640);
nor U7049 (N_7049,N_1986,N_4200);
nor U7050 (N_7050,N_1640,N_1713);
or U7051 (N_7051,N_405,N_1839);
or U7052 (N_7052,N_3163,N_4389);
and U7053 (N_7053,N_4185,N_3399);
and U7054 (N_7054,N_2269,N_3022);
nor U7055 (N_7055,N_1548,N_2319);
xor U7056 (N_7056,N_4569,N_4065);
and U7057 (N_7057,N_1144,N_377);
or U7058 (N_7058,N_1579,N_825);
nand U7059 (N_7059,N_4624,N_1086);
nor U7060 (N_7060,N_2805,N_3639);
and U7061 (N_7061,N_1717,N_1723);
or U7062 (N_7062,N_3141,N_387);
or U7063 (N_7063,N_1559,N_323);
xor U7064 (N_7064,N_2255,N_3064);
xor U7065 (N_7065,N_1486,N_3830);
or U7066 (N_7066,N_1114,N_2061);
and U7067 (N_7067,N_1227,N_1935);
nand U7068 (N_7068,N_1397,N_3849);
nand U7069 (N_7069,N_1800,N_951);
or U7070 (N_7070,N_3798,N_1288);
nor U7071 (N_7071,N_235,N_1989);
nor U7072 (N_7072,N_2458,N_2920);
nand U7073 (N_7073,N_3062,N_3228);
or U7074 (N_7074,N_2378,N_2053);
nor U7075 (N_7075,N_2841,N_2940);
xnor U7076 (N_7076,N_3945,N_363);
nand U7077 (N_7077,N_2561,N_3929);
nor U7078 (N_7078,N_164,N_4752);
xor U7079 (N_7079,N_2488,N_461);
nand U7080 (N_7080,N_1591,N_289);
nand U7081 (N_7081,N_1098,N_4014);
nor U7082 (N_7082,N_4234,N_962);
nor U7083 (N_7083,N_4665,N_3038);
nand U7084 (N_7084,N_699,N_990);
nand U7085 (N_7085,N_1812,N_4206);
nor U7086 (N_7086,N_1180,N_2768);
and U7087 (N_7087,N_2013,N_1085);
or U7088 (N_7088,N_3106,N_3869);
and U7089 (N_7089,N_3666,N_1531);
and U7090 (N_7090,N_4049,N_1882);
nor U7091 (N_7091,N_3290,N_2391);
or U7092 (N_7092,N_695,N_1006);
and U7093 (N_7093,N_1237,N_4329);
nor U7094 (N_7094,N_3800,N_1547);
or U7095 (N_7095,N_2385,N_3159);
and U7096 (N_7096,N_168,N_2691);
and U7097 (N_7097,N_3404,N_1190);
nand U7098 (N_7098,N_1017,N_2340);
nand U7099 (N_7099,N_1520,N_1493);
or U7100 (N_7100,N_2107,N_786);
nand U7101 (N_7101,N_4382,N_1344);
xor U7102 (N_7102,N_4529,N_2807);
nand U7103 (N_7103,N_414,N_1963);
and U7104 (N_7104,N_1585,N_2888);
nand U7105 (N_7105,N_4450,N_1595);
and U7106 (N_7106,N_2552,N_4053);
nand U7107 (N_7107,N_4961,N_118);
nor U7108 (N_7108,N_4068,N_1938);
and U7109 (N_7109,N_4807,N_1189);
and U7110 (N_7110,N_339,N_1638);
nand U7111 (N_7111,N_3599,N_4897);
nand U7112 (N_7112,N_537,N_476);
nand U7113 (N_7113,N_3388,N_1538);
xor U7114 (N_7114,N_418,N_3050);
and U7115 (N_7115,N_2127,N_4744);
nand U7116 (N_7116,N_664,N_3193);
or U7117 (N_7117,N_1071,N_4853);
or U7118 (N_7118,N_170,N_244);
and U7119 (N_7119,N_4114,N_266);
or U7120 (N_7120,N_2838,N_1955);
nand U7121 (N_7121,N_4613,N_212);
nor U7122 (N_7122,N_4690,N_4930);
xnor U7123 (N_7123,N_1907,N_1676);
or U7124 (N_7124,N_503,N_1915);
and U7125 (N_7125,N_35,N_1201);
nand U7126 (N_7126,N_1021,N_595);
or U7127 (N_7127,N_4036,N_2010);
nor U7128 (N_7128,N_2493,N_2512);
or U7129 (N_7129,N_3017,N_2556);
nand U7130 (N_7130,N_4369,N_31);
xor U7131 (N_7131,N_2088,N_2283);
nand U7132 (N_7132,N_2405,N_3672);
nor U7133 (N_7133,N_2663,N_1635);
and U7134 (N_7134,N_818,N_867);
nand U7135 (N_7135,N_2598,N_2094);
or U7136 (N_7136,N_711,N_1601);
nand U7137 (N_7137,N_3504,N_964);
nor U7138 (N_7138,N_1171,N_1789);
xnor U7139 (N_7139,N_2313,N_1018);
nor U7140 (N_7140,N_229,N_2105);
nand U7141 (N_7141,N_3579,N_755);
nor U7142 (N_7142,N_2431,N_1569);
xor U7143 (N_7143,N_1243,N_1466);
or U7144 (N_7144,N_4667,N_2802);
and U7145 (N_7145,N_2987,N_4918);
and U7146 (N_7146,N_2148,N_1382);
nand U7147 (N_7147,N_2041,N_781);
xor U7148 (N_7148,N_725,N_2114);
nor U7149 (N_7149,N_4847,N_539);
nor U7150 (N_7150,N_370,N_3339);
or U7151 (N_7151,N_1797,N_692);
nor U7152 (N_7152,N_4633,N_4804);
nor U7153 (N_7153,N_301,N_1024);
nand U7154 (N_7154,N_4905,N_3324);
and U7155 (N_7155,N_4092,N_3973);
nor U7156 (N_7156,N_4936,N_1282);
nand U7157 (N_7157,N_4080,N_75);
nor U7158 (N_7158,N_1383,N_3289);
and U7159 (N_7159,N_67,N_4297);
nor U7160 (N_7160,N_2991,N_3523);
nand U7161 (N_7161,N_3229,N_4028);
nand U7162 (N_7162,N_4287,N_564);
and U7163 (N_7163,N_3406,N_60);
nor U7164 (N_7164,N_76,N_1795);
nand U7165 (N_7165,N_3028,N_4556);
nand U7166 (N_7166,N_783,N_1117);
nor U7167 (N_7167,N_1064,N_4983);
nor U7168 (N_7168,N_3262,N_3440);
nor U7169 (N_7169,N_2632,N_429);
xor U7170 (N_7170,N_707,N_2295);
and U7171 (N_7171,N_593,N_2916);
nor U7172 (N_7172,N_764,N_4663);
nor U7173 (N_7173,N_1978,N_4655);
nor U7174 (N_7174,N_731,N_1443);
nand U7175 (N_7175,N_4706,N_2015);
and U7176 (N_7176,N_1980,N_2413);
nor U7177 (N_7177,N_2705,N_2435);
nor U7178 (N_7178,N_2174,N_785);
nor U7179 (N_7179,N_609,N_2523);
nor U7180 (N_7180,N_1611,N_3708);
or U7181 (N_7181,N_4210,N_809);
nand U7182 (N_7182,N_2422,N_4390);
and U7183 (N_7183,N_3792,N_1313);
xor U7184 (N_7184,N_2260,N_4861);
nor U7185 (N_7185,N_1104,N_1416);
nor U7186 (N_7186,N_2881,N_4999);
or U7187 (N_7187,N_2966,N_1505);
nor U7188 (N_7188,N_4343,N_1514);
or U7189 (N_7189,N_269,N_71);
nand U7190 (N_7190,N_1082,N_4072);
and U7191 (N_7191,N_819,N_4808);
and U7192 (N_7192,N_4300,N_2829);
nand U7193 (N_7193,N_2345,N_3694);
nand U7194 (N_7194,N_2724,N_627);
nor U7195 (N_7195,N_4799,N_3351);
nor U7196 (N_7196,N_1695,N_2776);
and U7197 (N_7197,N_1170,N_4491);
or U7198 (N_7198,N_941,N_4298);
nor U7199 (N_7199,N_3602,N_982);
and U7200 (N_7200,N_296,N_1751);
nand U7201 (N_7201,N_4582,N_2541);
or U7202 (N_7202,N_2367,N_2539);
nand U7203 (N_7203,N_3716,N_276);
nand U7204 (N_7204,N_559,N_2800);
or U7205 (N_7205,N_3148,N_1328);
and U7206 (N_7206,N_1134,N_1513);
and U7207 (N_7207,N_3081,N_2418);
nand U7208 (N_7208,N_2076,N_2634);
nor U7209 (N_7209,N_116,N_2195);
nand U7210 (N_7210,N_1245,N_3750);
nor U7211 (N_7211,N_3712,N_3282);
or U7212 (N_7212,N_2535,N_1078);
nor U7213 (N_7213,N_3158,N_3988);
nand U7214 (N_7214,N_3738,N_273);
xnor U7215 (N_7215,N_4841,N_1162);
and U7216 (N_7216,N_3012,N_4380);
and U7217 (N_7217,N_606,N_1059);
and U7218 (N_7218,N_3534,N_3769);
and U7219 (N_7219,N_2421,N_2113);
nand U7220 (N_7220,N_3899,N_3733);
nor U7221 (N_7221,N_3103,N_2432);
or U7222 (N_7222,N_2919,N_839);
nor U7223 (N_7223,N_2519,N_1929);
xnor U7224 (N_7224,N_1813,N_4165);
and U7225 (N_7225,N_3185,N_623);
nand U7226 (N_7226,N_4821,N_744);
nor U7227 (N_7227,N_280,N_2347);
or U7228 (N_7228,N_3564,N_1767);
and U7229 (N_7229,N_827,N_4698);
nand U7230 (N_7230,N_4095,N_686);
xnor U7231 (N_7231,N_480,N_2337);
nor U7232 (N_7232,N_3853,N_373);
nand U7233 (N_7233,N_310,N_4006);
xor U7234 (N_7234,N_4257,N_491);
nand U7235 (N_7235,N_2170,N_1322);
nor U7236 (N_7236,N_2307,N_400);
or U7237 (N_7237,N_4471,N_730);
or U7238 (N_7238,N_2927,N_1682);
nor U7239 (N_7239,N_4583,N_713);
and U7240 (N_7240,N_850,N_1139);
nor U7241 (N_7241,N_4235,N_1663);
nor U7242 (N_7242,N_2850,N_4249);
and U7243 (N_7243,N_2980,N_4096);
xor U7244 (N_7244,N_2116,N_1184);
xor U7245 (N_7245,N_3562,N_126);
or U7246 (N_7246,N_162,N_3055);
nand U7247 (N_7247,N_3084,N_2750);
nor U7248 (N_7248,N_912,N_3527);
nand U7249 (N_7249,N_4318,N_4187);
nor U7250 (N_7250,N_973,N_1031);
nand U7251 (N_7251,N_2359,N_2533);
nand U7252 (N_7252,N_4480,N_3178);
and U7253 (N_7253,N_1890,N_3761);
nand U7254 (N_7254,N_1137,N_193);
or U7255 (N_7255,N_2668,N_745);
or U7256 (N_7256,N_2896,N_100);
nand U7257 (N_7257,N_1634,N_3667);
or U7258 (N_7258,N_2111,N_616);
or U7259 (N_7259,N_2014,N_4749);
nand U7260 (N_7260,N_4428,N_2126);
nor U7261 (N_7261,N_3258,N_811);
or U7262 (N_7262,N_1274,N_4520);
nand U7263 (N_7263,N_4573,N_3211);
nor U7264 (N_7264,N_3937,N_3243);
nand U7265 (N_7265,N_2863,N_1446);
or U7266 (N_7266,N_4954,N_268);
and U7267 (N_7267,N_830,N_1552);
and U7268 (N_7268,N_2814,N_3248);
nand U7269 (N_7269,N_4490,N_2913);
nor U7270 (N_7270,N_3300,N_1922);
and U7271 (N_7271,N_3365,N_1498);
and U7272 (N_7272,N_2463,N_2929);
or U7273 (N_7273,N_3888,N_3165);
and U7274 (N_7274,N_2012,N_1293);
nand U7275 (N_7275,N_4830,N_1286);
and U7276 (N_7276,N_103,N_3015);
or U7277 (N_7277,N_2335,N_657);
or U7278 (N_7278,N_203,N_1900);
nand U7279 (N_7279,N_2977,N_4253);
and U7280 (N_7280,N_3411,N_485);
and U7281 (N_7281,N_3559,N_3032);
and U7282 (N_7282,N_3097,N_3556);
or U7283 (N_7283,N_1026,N_1371);
nor U7284 (N_7284,N_3866,N_3132);
or U7285 (N_7285,N_3453,N_334);
and U7286 (N_7286,N_3137,N_4059);
nand U7287 (N_7287,N_1263,N_4836);
or U7288 (N_7288,N_3313,N_1688);
and U7289 (N_7289,N_3197,N_4009);
or U7290 (N_7290,N_283,N_4193);
and U7291 (N_7291,N_926,N_746);
nand U7292 (N_7292,N_199,N_1582);
nand U7293 (N_7293,N_2655,N_714);
and U7294 (N_7294,N_4461,N_3099);
or U7295 (N_7295,N_655,N_4616);
or U7296 (N_7296,N_4695,N_320);
xor U7297 (N_7297,N_1046,N_3113);
xnor U7298 (N_7298,N_2826,N_3975);
nand U7299 (N_7299,N_868,N_1142);
nor U7300 (N_7300,N_11,N_66);
xnor U7301 (N_7301,N_1633,N_3812);
nor U7302 (N_7302,N_3361,N_1976);
or U7303 (N_7303,N_3622,N_613);
nand U7304 (N_7304,N_157,N_685);
and U7305 (N_7305,N_2962,N_1718);
or U7306 (N_7306,N_147,N_3034);
or U7307 (N_7307,N_1204,N_544);
nor U7308 (N_7308,N_4500,N_4384);
or U7309 (N_7309,N_3156,N_3758);
and U7310 (N_7310,N_856,N_3004);
or U7311 (N_7311,N_879,N_3707);
xor U7312 (N_7312,N_4771,N_136);
and U7313 (N_7313,N_916,N_908);
and U7314 (N_7314,N_2988,N_3358);
or U7315 (N_7315,N_251,N_3821);
nand U7316 (N_7316,N_2606,N_3307);
or U7317 (N_7317,N_2956,N_2062);
and U7318 (N_7318,N_1692,N_3181);
xnor U7319 (N_7319,N_4986,N_2537);
nand U7320 (N_7320,N_1747,N_1248);
and U7321 (N_7321,N_3212,N_3373);
nand U7322 (N_7322,N_2072,N_3010);
nand U7323 (N_7323,N_223,N_2218);
or U7324 (N_7324,N_1746,N_1563);
xnor U7325 (N_7325,N_2095,N_353);
and U7326 (N_7326,N_4970,N_4367);
or U7327 (N_7327,N_2779,N_2924);
or U7328 (N_7328,N_240,N_4542);
nor U7329 (N_7329,N_2009,N_3297);
nor U7330 (N_7330,N_3446,N_1011);
nand U7331 (N_7331,N_2179,N_2594);
or U7332 (N_7332,N_2969,N_2995);
nor U7333 (N_7333,N_1749,N_215);
and U7334 (N_7334,N_4169,N_1588);
and U7335 (N_7335,N_864,N_2489);
nand U7336 (N_7336,N_1066,N_3166);
and U7337 (N_7337,N_4568,N_3791);
and U7338 (N_7338,N_1218,N_3958);
and U7339 (N_7339,N_2442,N_4047);
nor U7340 (N_7340,N_3847,N_3392);
nor U7341 (N_7341,N_2557,N_620);
or U7342 (N_7342,N_846,N_2282);
and U7343 (N_7343,N_185,N_3681);
or U7344 (N_7344,N_4864,N_1061);
nor U7345 (N_7345,N_1561,N_3227);
nand U7346 (N_7346,N_401,N_1912);
and U7347 (N_7347,N_1544,N_4757);
and U7348 (N_7348,N_2767,N_2799);
nand U7349 (N_7349,N_1499,N_2636);
and U7350 (N_7350,N_2714,N_93);
or U7351 (N_7351,N_1823,N_1452);
xnor U7352 (N_7352,N_4475,N_466);
nor U7353 (N_7353,N_4275,N_1233);
nand U7354 (N_7354,N_4673,N_4481);
nor U7355 (N_7355,N_282,N_3794);
or U7356 (N_7356,N_2046,N_568);
nor U7357 (N_7357,N_961,N_2011);
and U7358 (N_7358,N_3259,N_2206);
nand U7359 (N_7359,N_2301,N_3489);
xor U7360 (N_7360,N_2425,N_2666);
nor U7361 (N_7361,N_230,N_3825);
nor U7362 (N_7362,N_4209,N_3415);
and U7363 (N_7363,N_1181,N_1461);
nor U7364 (N_7364,N_2603,N_2024);
and U7365 (N_7365,N_1070,N_3236);
or U7366 (N_7366,N_4557,N_3176);
nor U7367 (N_7367,N_2220,N_3931);
or U7368 (N_7368,N_668,N_2617);
or U7369 (N_7369,N_4010,N_1541);
xnor U7370 (N_7370,N_1743,N_4722);
xnor U7371 (N_7371,N_3627,N_3659);
nand U7372 (N_7372,N_2676,N_4537);
nand U7373 (N_7373,N_4874,N_2178);
and U7374 (N_7374,N_3465,N_3356);
nand U7375 (N_7375,N_4531,N_527);
or U7376 (N_7376,N_1820,N_829);
nor U7377 (N_7377,N_331,N_1810);
or U7378 (N_7378,N_1686,N_4644);
nand U7379 (N_7379,N_2879,N_541);
or U7380 (N_7380,N_3396,N_2213);
xnor U7381 (N_7381,N_4580,N_1412);
or U7382 (N_7382,N_810,N_4310);
xor U7383 (N_7383,N_77,N_3765);
or U7384 (N_7384,N_1396,N_1794);
or U7385 (N_7385,N_2394,N_1146);
nand U7386 (N_7386,N_4512,N_4893);
or U7387 (N_7387,N_3797,N_371);
and U7388 (N_7388,N_2791,N_4170);
nand U7389 (N_7389,N_4937,N_1598);
and U7390 (N_7390,N_1568,N_4411);
nor U7391 (N_7391,N_653,N_1081);
and U7392 (N_7392,N_1477,N_1753);
nand U7393 (N_7393,N_1654,N_3841);
nor U7394 (N_7394,N_2973,N_1518);
nor U7395 (N_7395,N_2300,N_815);
xor U7396 (N_7396,N_3145,N_1740);
nand U7397 (N_7397,N_3802,N_143);
or U7398 (N_7398,N_1036,N_3664);
nand U7399 (N_7399,N_179,N_3172);
xor U7400 (N_7400,N_1030,N_3965);
or U7401 (N_7401,N_543,N_4271);
and U7402 (N_7402,N_2592,N_1351);
or U7403 (N_7403,N_2341,N_3497);
and U7404 (N_7404,N_3656,N_3085);
and U7405 (N_7405,N_3327,N_4825);
nand U7406 (N_7406,N_4301,N_648);
nor U7407 (N_7407,N_697,N_2288);
and U7408 (N_7408,N_1128,N_4027);
xnor U7409 (N_7409,N_602,N_1022);
nor U7410 (N_7410,N_1339,N_2996);
xor U7411 (N_7411,N_859,N_1299);
and U7412 (N_7412,N_1023,N_1936);
and U7413 (N_7413,N_454,N_1055);
and U7414 (N_7414,N_561,N_1035);
nand U7415 (N_7415,N_2743,N_1909);
and U7416 (N_7416,N_3947,N_1960);
and U7417 (N_7417,N_3964,N_1631);
or U7418 (N_7418,N_2299,N_4133);
nor U7419 (N_7419,N_4917,N_444);
nor U7420 (N_7420,N_3040,N_3203);
and U7421 (N_7421,N_4156,N_4885);
and U7422 (N_7422,N_1195,N_4630);
nor U7423 (N_7423,N_579,N_1270);
nor U7424 (N_7424,N_3904,N_163);
xor U7425 (N_7425,N_2890,N_3598);
or U7426 (N_7426,N_3265,N_2086);
nand U7427 (N_7427,N_2903,N_3474);
nor U7428 (N_7428,N_156,N_813);
nor U7429 (N_7429,N_1959,N_285);
nand U7430 (N_7430,N_2219,N_4484);
xnor U7431 (N_7431,N_2722,N_3374);
nand U7432 (N_7432,N_1555,N_1423);
or U7433 (N_7433,N_1776,N_4299);
nand U7434 (N_7434,N_4691,N_3063);
or U7435 (N_7435,N_4321,N_545);
nand U7436 (N_7436,N_3405,N_687);
nor U7437 (N_7437,N_3495,N_1473);
nor U7438 (N_7438,N_1152,N_1973);
nor U7439 (N_7439,N_4063,N_1780);
nor U7440 (N_7440,N_663,N_3164);
and U7441 (N_7441,N_2921,N_4074);
and U7442 (N_7442,N_3129,N_1294);
and U7443 (N_7443,N_3959,N_2320);
and U7444 (N_7444,N_2579,N_778);
or U7445 (N_7445,N_2868,N_4721);
nand U7446 (N_7446,N_1364,N_2501);
and U7447 (N_7447,N_513,N_556);
nor U7448 (N_7448,N_4370,N_689);
nor U7449 (N_7449,N_1570,N_2253);
nand U7450 (N_7450,N_4619,N_2551);
and U7451 (N_7451,N_1232,N_2796);
or U7452 (N_7452,N_1194,N_4548);
nand U7453 (N_7453,N_2270,N_15);
and U7454 (N_7454,N_4439,N_2897);
nor U7455 (N_7455,N_4433,N_316);
and U7456 (N_7456,N_1884,N_1970);
nand U7457 (N_7457,N_4784,N_3316);
nor U7458 (N_7458,N_3554,N_2350);
nand U7459 (N_7459,N_4245,N_824);
or U7460 (N_7460,N_1783,N_1334);
nor U7461 (N_7461,N_3746,N_4750);
nor U7462 (N_7462,N_3723,N_1057);
nand U7463 (N_7463,N_2426,N_4595);
nand U7464 (N_7464,N_1868,N_465);
nor U7465 (N_7465,N_238,N_415);
nor U7466 (N_7466,N_3104,N_1701);
and U7467 (N_7467,N_2224,N_2471);
and U7468 (N_7468,N_4216,N_1105);
or U7469 (N_7469,N_4880,N_3157);
nor U7470 (N_7470,N_2143,N_1271);
xor U7471 (N_7471,N_3592,N_924);
xor U7472 (N_7472,N_410,N_4019);
nor U7473 (N_7473,N_2640,N_2368);
nor U7474 (N_7474,N_3215,N_1437);
xnor U7475 (N_7475,N_3827,N_2930);
and U7476 (N_7476,N_1439,N_4233);
nor U7477 (N_7477,N_483,N_888);
xnor U7478 (N_7478,N_3545,N_3477);
or U7479 (N_7479,N_4988,N_2199);
or U7480 (N_7480,N_1223,N_4346);
nor U7481 (N_7481,N_1379,N_3475);
nor U7482 (N_7482,N_4598,N_186);
xnor U7483 (N_7483,N_4217,N_638);
or U7484 (N_7484,N_2783,N_1394);
or U7485 (N_7485,N_766,N_4736);
or U7486 (N_7486,N_1384,N_1892);
xor U7487 (N_7487,N_33,N_796);
nor U7488 (N_7488,N_319,N_4713);
and U7489 (N_7489,N_326,N_599);
and U7490 (N_7490,N_1445,N_1738);
or U7491 (N_7491,N_4659,N_1803);
or U7492 (N_7492,N_4098,N_4319);
or U7493 (N_7493,N_3833,N_1809);
or U7494 (N_7494,N_95,N_2798);
nor U7495 (N_7495,N_3210,N_299);
nor U7496 (N_7496,N_4726,N_4309);
and U7497 (N_7497,N_1801,N_424);
nand U7498 (N_7498,N_2565,N_2856);
or U7499 (N_7499,N_3751,N_2436);
nor U7500 (N_7500,N_1815,N_2516);
or U7501 (N_7501,N_4897,N_4380);
or U7502 (N_7502,N_2773,N_4539);
and U7503 (N_7503,N_1152,N_2223);
nand U7504 (N_7504,N_3277,N_4841);
xnor U7505 (N_7505,N_2805,N_2680);
and U7506 (N_7506,N_2691,N_1619);
xnor U7507 (N_7507,N_28,N_2159);
xor U7508 (N_7508,N_2789,N_1812);
and U7509 (N_7509,N_3787,N_3629);
and U7510 (N_7510,N_2332,N_297);
nor U7511 (N_7511,N_2252,N_1542);
nor U7512 (N_7512,N_4384,N_2785);
or U7513 (N_7513,N_2183,N_3956);
or U7514 (N_7514,N_265,N_4141);
xor U7515 (N_7515,N_3391,N_1507);
nand U7516 (N_7516,N_2895,N_2492);
xor U7517 (N_7517,N_2364,N_874);
or U7518 (N_7518,N_4953,N_2727);
xor U7519 (N_7519,N_130,N_2608);
nand U7520 (N_7520,N_3178,N_1321);
and U7521 (N_7521,N_2158,N_1014);
nand U7522 (N_7522,N_3100,N_3879);
nand U7523 (N_7523,N_4587,N_4143);
nand U7524 (N_7524,N_238,N_3891);
and U7525 (N_7525,N_1784,N_4479);
xnor U7526 (N_7526,N_181,N_2360);
or U7527 (N_7527,N_2687,N_50);
nand U7528 (N_7528,N_1586,N_4958);
nor U7529 (N_7529,N_4005,N_3226);
nand U7530 (N_7530,N_4516,N_4871);
nand U7531 (N_7531,N_423,N_1067);
and U7532 (N_7532,N_335,N_486);
and U7533 (N_7533,N_1673,N_2250);
nand U7534 (N_7534,N_1452,N_2166);
or U7535 (N_7535,N_4218,N_4619);
nand U7536 (N_7536,N_4071,N_4803);
nor U7537 (N_7537,N_4851,N_1725);
and U7538 (N_7538,N_30,N_1251);
nor U7539 (N_7539,N_1270,N_1055);
nand U7540 (N_7540,N_2038,N_4541);
nor U7541 (N_7541,N_3550,N_3451);
or U7542 (N_7542,N_2086,N_4617);
and U7543 (N_7543,N_2548,N_1231);
or U7544 (N_7544,N_1863,N_3927);
nand U7545 (N_7545,N_2596,N_4266);
nor U7546 (N_7546,N_1666,N_1960);
or U7547 (N_7547,N_456,N_3587);
or U7548 (N_7548,N_349,N_4885);
nand U7549 (N_7549,N_3124,N_670);
nor U7550 (N_7550,N_2981,N_1416);
or U7551 (N_7551,N_3678,N_4977);
nand U7552 (N_7552,N_3583,N_3120);
nand U7553 (N_7553,N_3753,N_550);
nor U7554 (N_7554,N_2141,N_3419);
nand U7555 (N_7555,N_3019,N_3324);
nor U7556 (N_7556,N_1414,N_3111);
nor U7557 (N_7557,N_2944,N_604);
nand U7558 (N_7558,N_1366,N_2788);
or U7559 (N_7559,N_991,N_4090);
nor U7560 (N_7560,N_1179,N_1122);
or U7561 (N_7561,N_1675,N_3934);
xor U7562 (N_7562,N_1469,N_676);
nor U7563 (N_7563,N_4041,N_3487);
or U7564 (N_7564,N_509,N_4276);
or U7565 (N_7565,N_674,N_2466);
nand U7566 (N_7566,N_3251,N_4390);
xor U7567 (N_7567,N_769,N_3948);
or U7568 (N_7568,N_1857,N_4885);
or U7569 (N_7569,N_2643,N_4595);
nand U7570 (N_7570,N_721,N_3483);
nand U7571 (N_7571,N_1847,N_2801);
nor U7572 (N_7572,N_1203,N_3108);
or U7573 (N_7573,N_3168,N_341);
nand U7574 (N_7574,N_3553,N_1833);
or U7575 (N_7575,N_2829,N_4956);
xor U7576 (N_7576,N_3786,N_1818);
and U7577 (N_7577,N_1519,N_1482);
nand U7578 (N_7578,N_1099,N_2502);
nand U7579 (N_7579,N_3997,N_532);
nor U7580 (N_7580,N_2179,N_906);
and U7581 (N_7581,N_1884,N_2445);
or U7582 (N_7582,N_4208,N_4850);
or U7583 (N_7583,N_1518,N_1224);
nand U7584 (N_7584,N_2779,N_3665);
and U7585 (N_7585,N_3814,N_4824);
or U7586 (N_7586,N_3569,N_1815);
or U7587 (N_7587,N_910,N_1533);
or U7588 (N_7588,N_2766,N_91);
or U7589 (N_7589,N_1713,N_2915);
nand U7590 (N_7590,N_1809,N_151);
nor U7591 (N_7591,N_4158,N_1387);
xor U7592 (N_7592,N_371,N_4024);
or U7593 (N_7593,N_3617,N_159);
nor U7594 (N_7594,N_2009,N_3202);
nor U7595 (N_7595,N_2669,N_1728);
or U7596 (N_7596,N_2130,N_885);
and U7597 (N_7597,N_2005,N_2437);
nor U7598 (N_7598,N_3630,N_2186);
xor U7599 (N_7599,N_71,N_1241);
xor U7600 (N_7600,N_3600,N_2904);
and U7601 (N_7601,N_1412,N_2733);
nand U7602 (N_7602,N_2022,N_2532);
or U7603 (N_7603,N_3550,N_25);
or U7604 (N_7604,N_2962,N_1703);
nand U7605 (N_7605,N_362,N_1185);
or U7606 (N_7606,N_482,N_803);
nor U7607 (N_7607,N_4334,N_1830);
and U7608 (N_7608,N_3802,N_4503);
nand U7609 (N_7609,N_4203,N_3808);
nand U7610 (N_7610,N_2179,N_736);
xor U7611 (N_7611,N_613,N_1647);
xor U7612 (N_7612,N_1281,N_2331);
nor U7613 (N_7613,N_1596,N_105);
nand U7614 (N_7614,N_2789,N_4273);
or U7615 (N_7615,N_4333,N_747);
and U7616 (N_7616,N_4283,N_1790);
nand U7617 (N_7617,N_4241,N_2890);
and U7618 (N_7618,N_1766,N_2424);
and U7619 (N_7619,N_305,N_942);
or U7620 (N_7620,N_3712,N_2018);
nand U7621 (N_7621,N_533,N_3235);
and U7622 (N_7622,N_4863,N_4795);
nor U7623 (N_7623,N_2987,N_1892);
and U7624 (N_7624,N_1056,N_3386);
or U7625 (N_7625,N_1784,N_4108);
or U7626 (N_7626,N_4177,N_4836);
and U7627 (N_7627,N_840,N_2474);
and U7628 (N_7628,N_2988,N_494);
nor U7629 (N_7629,N_728,N_2901);
nor U7630 (N_7630,N_1777,N_1783);
and U7631 (N_7631,N_2346,N_718);
and U7632 (N_7632,N_4686,N_519);
or U7633 (N_7633,N_248,N_3387);
nand U7634 (N_7634,N_1397,N_4429);
nor U7635 (N_7635,N_3924,N_3991);
and U7636 (N_7636,N_382,N_1303);
nand U7637 (N_7637,N_4344,N_2287);
xnor U7638 (N_7638,N_3539,N_4690);
and U7639 (N_7639,N_3130,N_4272);
or U7640 (N_7640,N_4815,N_1488);
or U7641 (N_7641,N_705,N_2586);
or U7642 (N_7642,N_1190,N_2276);
or U7643 (N_7643,N_4517,N_753);
nand U7644 (N_7644,N_569,N_2541);
nor U7645 (N_7645,N_3736,N_2499);
or U7646 (N_7646,N_2466,N_4325);
xnor U7647 (N_7647,N_4057,N_743);
and U7648 (N_7648,N_1493,N_1912);
nor U7649 (N_7649,N_4113,N_1519);
and U7650 (N_7650,N_1214,N_1882);
or U7651 (N_7651,N_896,N_795);
or U7652 (N_7652,N_4031,N_2949);
and U7653 (N_7653,N_4559,N_1716);
nor U7654 (N_7654,N_2203,N_3163);
and U7655 (N_7655,N_3163,N_4647);
and U7656 (N_7656,N_3348,N_66);
nor U7657 (N_7657,N_1763,N_4964);
nor U7658 (N_7658,N_4945,N_110);
nand U7659 (N_7659,N_3976,N_4277);
or U7660 (N_7660,N_2726,N_3330);
nor U7661 (N_7661,N_2564,N_1157);
and U7662 (N_7662,N_4890,N_1200);
nor U7663 (N_7663,N_4953,N_2255);
nand U7664 (N_7664,N_1880,N_1703);
nor U7665 (N_7665,N_3592,N_1656);
and U7666 (N_7666,N_1570,N_4991);
and U7667 (N_7667,N_4095,N_2523);
xnor U7668 (N_7668,N_1823,N_351);
and U7669 (N_7669,N_3132,N_864);
or U7670 (N_7670,N_412,N_4147);
or U7671 (N_7671,N_172,N_1453);
nor U7672 (N_7672,N_3857,N_2239);
nand U7673 (N_7673,N_4573,N_4882);
nand U7674 (N_7674,N_167,N_4171);
xnor U7675 (N_7675,N_2225,N_3680);
or U7676 (N_7676,N_3358,N_4526);
and U7677 (N_7677,N_3353,N_1468);
and U7678 (N_7678,N_1027,N_449);
nand U7679 (N_7679,N_4910,N_4992);
nor U7680 (N_7680,N_2769,N_2886);
nor U7681 (N_7681,N_608,N_1157);
or U7682 (N_7682,N_2714,N_173);
or U7683 (N_7683,N_2606,N_4739);
and U7684 (N_7684,N_78,N_712);
nand U7685 (N_7685,N_2653,N_1826);
or U7686 (N_7686,N_849,N_3197);
and U7687 (N_7687,N_2345,N_1129);
nor U7688 (N_7688,N_3102,N_4728);
and U7689 (N_7689,N_1725,N_1513);
nand U7690 (N_7690,N_2534,N_85);
nor U7691 (N_7691,N_4608,N_2023);
nand U7692 (N_7692,N_4707,N_269);
xnor U7693 (N_7693,N_2731,N_3861);
nor U7694 (N_7694,N_2388,N_3902);
nor U7695 (N_7695,N_4929,N_2850);
or U7696 (N_7696,N_3187,N_3609);
and U7697 (N_7697,N_4688,N_4701);
and U7698 (N_7698,N_2325,N_1781);
nor U7699 (N_7699,N_4345,N_3304);
nor U7700 (N_7700,N_104,N_2721);
and U7701 (N_7701,N_1956,N_3323);
nand U7702 (N_7702,N_3460,N_1220);
and U7703 (N_7703,N_1797,N_4257);
xnor U7704 (N_7704,N_3544,N_2698);
nand U7705 (N_7705,N_3077,N_3584);
or U7706 (N_7706,N_3150,N_4863);
nand U7707 (N_7707,N_498,N_3641);
nand U7708 (N_7708,N_2744,N_3467);
and U7709 (N_7709,N_708,N_382);
nand U7710 (N_7710,N_2451,N_1379);
nor U7711 (N_7711,N_4161,N_1609);
nand U7712 (N_7712,N_1515,N_3879);
nor U7713 (N_7713,N_468,N_270);
and U7714 (N_7714,N_495,N_4319);
nor U7715 (N_7715,N_2472,N_2348);
nor U7716 (N_7716,N_619,N_4503);
or U7717 (N_7717,N_1725,N_3848);
and U7718 (N_7718,N_4056,N_3392);
nor U7719 (N_7719,N_3552,N_2249);
and U7720 (N_7720,N_2650,N_1053);
xnor U7721 (N_7721,N_1427,N_155);
nand U7722 (N_7722,N_2019,N_558);
nand U7723 (N_7723,N_4582,N_202);
or U7724 (N_7724,N_2645,N_2331);
nand U7725 (N_7725,N_3793,N_3174);
nand U7726 (N_7726,N_1577,N_4855);
and U7727 (N_7727,N_194,N_1474);
xor U7728 (N_7728,N_1587,N_2906);
nand U7729 (N_7729,N_1343,N_2160);
nand U7730 (N_7730,N_755,N_2041);
nand U7731 (N_7731,N_2458,N_4357);
nor U7732 (N_7732,N_527,N_899);
and U7733 (N_7733,N_3781,N_622);
nand U7734 (N_7734,N_1819,N_4786);
nand U7735 (N_7735,N_4887,N_3665);
xor U7736 (N_7736,N_4588,N_2867);
and U7737 (N_7737,N_1920,N_2252);
nand U7738 (N_7738,N_3226,N_3680);
or U7739 (N_7739,N_3600,N_2481);
or U7740 (N_7740,N_1403,N_1284);
and U7741 (N_7741,N_16,N_2980);
or U7742 (N_7742,N_3409,N_4294);
or U7743 (N_7743,N_1442,N_4291);
nor U7744 (N_7744,N_3008,N_4085);
nor U7745 (N_7745,N_4039,N_4165);
or U7746 (N_7746,N_2457,N_1562);
and U7747 (N_7747,N_2657,N_3364);
xor U7748 (N_7748,N_620,N_1031);
and U7749 (N_7749,N_4018,N_2835);
and U7750 (N_7750,N_378,N_302);
or U7751 (N_7751,N_2560,N_1683);
nor U7752 (N_7752,N_3932,N_3148);
or U7753 (N_7753,N_2654,N_4382);
nand U7754 (N_7754,N_3491,N_1340);
or U7755 (N_7755,N_573,N_3437);
or U7756 (N_7756,N_306,N_3153);
nand U7757 (N_7757,N_2395,N_918);
or U7758 (N_7758,N_1320,N_4150);
or U7759 (N_7759,N_2396,N_2854);
or U7760 (N_7760,N_2622,N_3981);
xor U7761 (N_7761,N_3825,N_27);
xor U7762 (N_7762,N_3860,N_49);
or U7763 (N_7763,N_2945,N_632);
nor U7764 (N_7764,N_181,N_710);
or U7765 (N_7765,N_1606,N_3130);
or U7766 (N_7766,N_1678,N_3886);
nand U7767 (N_7767,N_4733,N_3239);
xnor U7768 (N_7768,N_2536,N_2184);
nand U7769 (N_7769,N_3488,N_4769);
nand U7770 (N_7770,N_1785,N_4343);
nand U7771 (N_7771,N_1753,N_1945);
and U7772 (N_7772,N_82,N_4681);
and U7773 (N_7773,N_3025,N_2471);
nor U7774 (N_7774,N_1768,N_1870);
and U7775 (N_7775,N_1210,N_721);
nor U7776 (N_7776,N_3144,N_338);
nand U7777 (N_7777,N_3211,N_333);
nand U7778 (N_7778,N_4537,N_2563);
and U7779 (N_7779,N_4039,N_675);
or U7780 (N_7780,N_4312,N_42);
or U7781 (N_7781,N_3280,N_388);
nor U7782 (N_7782,N_4238,N_4956);
or U7783 (N_7783,N_4961,N_3609);
nor U7784 (N_7784,N_1501,N_3003);
and U7785 (N_7785,N_2245,N_2497);
and U7786 (N_7786,N_4209,N_3358);
and U7787 (N_7787,N_4531,N_943);
or U7788 (N_7788,N_961,N_1597);
or U7789 (N_7789,N_2561,N_862);
nand U7790 (N_7790,N_3727,N_772);
or U7791 (N_7791,N_4442,N_4163);
nor U7792 (N_7792,N_2517,N_2395);
or U7793 (N_7793,N_489,N_298);
xor U7794 (N_7794,N_1980,N_3863);
nand U7795 (N_7795,N_3163,N_3621);
or U7796 (N_7796,N_658,N_2665);
and U7797 (N_7797,N_2186,N_3729);
or U7798 (N_7798,N_4234,N_4822);
nor U7799 (N_7799,N_4942,N_3837);
nand U7800 (N_7800,N_3015,N_4519);
xnor U7801 (N_7801,N_4999,N_1088);
nand U7802 (N_7802,N_3183,N_2503);
or U7803 (N_7803,N_2041,N_2099);
nor U7804 (N_7804,N_2989,N_85);
xor U7805 (N_7805,N_4412,N_1297);
nor U7806 (N_7806,N_2231,N_704);
or U7807 (N_7807,N_3044,N_3421);
nand U7808 (N_7808,N_644,N_3434);
nand U7809 (N_7809,N_2043,N_2811);
nand U7810 (N_7810,N_4692,N_2107);
or U7811 (N_7811,N_1777,N_1734);
xnor U7812 (N_7812,N_2123,N_2873);
or U7813 (N_7813,N_2553,N_2294);
or U7814 (N_7814,N_4959,N_3761);
nor U7815 (N_7815,N_1752,N_1610);
or U7816 (N_7816,N_3969,N_3992);
nor U7817 (N_7817,N_2287,N_1199);
and U7818 (N_7818,N_4268,N_4344);
nand U7819 (N_7819,N_3616,N_3990);
or U7820 (N_7820,N_2634,N_2974);
nand U7821 (N_7821,N_1686,N_3629);
and U7822 (N_7822,N_909,N_3154);
xor U7823 (N_7823,N_3864,N_765);
xnor U7824 (N_7824,N_577,N_960);
nand U7825 (N_7825,N_614,N_2881);
or U7826 (N_7826,N_3351,N_2083);
or U7827 (N_7827,N_2047,N_2509);
nand U7828 (N_7828,N_934,N_560);
and U7829 (N_7829,N_2788,N_4101);
xor U7830 (N_7830,N_1830,N_3407);
or U7831 (N_7831,N_2685,N_2511);
nor U7832 (N_7832,N_4922,N_3674);
xor U7833 (N_7833,N_4849,N_680);
and U7834 (N_7834,N_4797,N_2093);
nand U7835 (N_7835,N_2922,N_3429);
and U7836 (N_7836,N_3255,N_358);
nand U7837 (N_7837,N_2143,N_4781);
or U7838 (N_7838,N_2115,N_4384);
nand U7839 (N_7839,N_4077,N_4531);
nor U7840 (N_7840,N_2011,N_612);
or U7841 (N_7841,N_1550,N_3698);
nand U7842 (N_7842,N_1061,N_497);
xnor U7843 (N_7843,N_3427,N_4355);
xor U7844 (N_7844,N_2631,N_2220);
nor U7845 (N_7845,N_348,N_4728);
nand U7846 (N_7846,N_4944,N_4871);
nor U7847 (N_7847,N_370,N_1844);
nand U7848 (N_7848,N_228,N_4622);
and U7849 (N_7849,N_229,N_3108);
nor U7850 (N_7850,N_2065,N_1748);
nor U7851 (N_7851,N_2179,N_3958);
nor U7852 (N_7852,N_3275,N_33);
xnor U7853 (N_7853,N_4971,N_2985);
or U7854 (N_7854,N_1779,N_2412);
nand U7855 (N_7855,N_2814,N_2455);
nor U7856 (N_7856,N_1495,N_4549);
nand U7857 (N_7857,N_4533,N_3718);
nor U7858 (N_7858,N_3820,N_4192);
nand U7859 (N_7859,N_4659,N_2252);
or U7860 (N_7860,N_1654,N_1483);
and U7861 (N_7861,N_2234,N_1387);
and U7862 (N_7862,N_2494,N_668);
nor U7863 (N_7863,N_882,N_4388);
and U7864 (N_7864,N_2235,N_434);
or U7865 (N_7865,N_3926,N_2459);
nand U7866 (N_7866,N_2684,N_2460);
nor U7867 (N_7867,N_2083,N_1445);
nand U7868 (N_7868,N_1484,N_3563);
nand U7869 (N_7869,N_411,N_405);
nand U7870 (N_7870,N_114,N_2881);
xnor U7871 (N_7871,N_4040,N_2247);
nand U7872 (N_7872,N_4952,N_2559);
and U7873 (N_7873,N_4771,N_86);
nor U7874 (N_7874,N_882,N_3933);
nand U7875 (N_7875,N_2941,N_4264);
nor U7876 (N_7876,N_4325,N_2392);
and U7877 (N_7877,N_670,N_2702);
or U7878 (N_7878,N_2288,N_43);
nand U7879 (N_7879,N_4473,N_2128);
xnor U7880 (N_7880,N_1054,N_1844);
nor U7881 (N_7881,N_4574,N_1987);
nand U7882 (N_7882,N_3659,N_2587);
xor U7883 (N_7883,N_304,N_3937);
nand U7884 (N_7884,N_4120,N_3944);
or U7885 (N_7885,N_4509,N_2644);
xnor U7886 (N_7886,N_1797,N_4009);
or U7887 (N_7887,N_637,N_1243);
nand U7888 (N_7888,N_1223,N_3692);
and U7889 (N_7889,N_2272,N_1587);
nand U7890 (N_7890,N_2224,N_3094);
and U7891 (N_7891,N_627,N_3477);
xor U7892 (N_7892,N_20,N_4944);
nor U7893 (N_7893,N_3872,N_3672);
or U7894 (N_7894,N_151,N_4666);
or U7895 (N_7895,N_1903,N_4163);
and U7896 (N_7896,N_4438,N_3425);
or U7897 (N_7897,N_2091,N_2079);
nand U7898 (N_7898,N_1344,N_3582);
nand U7899 (N_7899,N_3441,N_1823);
nand U7900 (N_7900,N_4320,N_4023);
and U7901 (N_7901,N_979,N_673);
xor U7902 (N_7902,N_248,N_2455);
and U7903 (N_7903,N_859,N_715);
nor U7904 (N_7904,N_1855,N_449);
or U7905 (N_7905,N_1472,N_784);
or U7906 (N_7906,N_2443,N_2751);
and U7907 (N_7907,N_4048,N_4896);
or U7908 (N_7908,N_3270,N_4560);
nand U7909 (N_7909,N_3993,N_4616);
and U7910 (N_7910,N_4742,N_1209);
nand U7911 (N_7911,N_2321,N_1152);
or U7912 (N_7912,N_2229,N_4724);
xnor U7913 (N_7913,N_934,N_3191);
and U7914 (N_7914,N_4281,N_1627);
or U7915 (N_7915,N_2793,N_3792);
or U7916 (N_7916,N_2723,N_3086);
and U7917 (N_7917,N_2658,N_4867);
xor U7918 (N_7918,N_900,N_4109);
and U7919 (N_7919,N_2556,N_1120);
or U7920 (N_7920,N_1354,N_778);
nor U7921 (N_7921,N_2989,N_2637);
and U7922 (N_7922,N_1960,N_2889);
nand U7923 (N_7923,N_897,N_725);
and U7924 (N_7924,N_1501,N_1703);
and U7925 (N_7925,N_3726,N_3007);
nor U7926 (N_7926,N_1911,N_1490);
nand U7927 (N_7927,N_144,N_2230);
and U7928 (N_7928,N_1213,N_3147);
nand U7929 (N_7929,N_2093,N_869);
and U7930 (N_7930,N_3211,N_3613);
nor U7931 (N_7931,N_545,N_1205);
nor U7932 (N_7932,N_4661,N_1455);
or U7933 (N_7933,N_1181,N_3277);
and U7934 (N_7934,N_2386,N_4799);
and U7935 (N_7935,N_2589,N_3482);
nor U7936 (N_7936,N_1665,N_111);
nor U7937 (N_7937,N_1969,N_900);
nand U7938 (N_7938,N_820,N_1971);
or U7939 (N_7939,N_1308,N_3391);
and U7940 (N_7940,N_1500,N_4930);
nor U7941 (N_7941,N_1932,N_4669);
nor U7942 (N_7942,N_2470,N_3901);
and U7943 (N_7943,N_4210,N_3381);
nand U7944 (N_7944,N_4375,N_3748);
and U7945 (N_7945,N_1936,N_4319);
xnor U7946 (N_7946,N_3986,N_3982);
and U7947 (N_7947,N_3883,N_2570);
xor U7948 (N_7948,N_3436,N_598);
nor U7949 (N_7949,N_1392,N_2381);
nand U7950 (N_7950,N_3045,N_421);
nor U7951 (N_7951,N_2862,N_2180);
nand U7952 (N_7952,N_283,N_721);
and U7953 (N_7953,N_3367,N_4327);
nor U7954 (N_7954,N_3370,N_4630);
or U7955 (N_7955,N_541,N_2325);
nand U7956 (N_7956,N_3639,N_811);
nand U7957 (N_7957,N_423,N_1554);
nand U7958 (N_7958,N_2940,N_85);
nor U7959 (N_7959,N_3802,N_3771);
and U7960 (N_7960,N_460,N_2018);
nor U7961 (N_7961,N_3362,N_307);
and U7962 (N_7962,N_386,N_1950);
nor U7963 (N_7963,N_3598,N_2078);
nand U7964 (N_7964,N_3812,N_4334);
nor U7965 (N_7965,N_4,N_4761);
nor U7966 (N_7966,N_2879,N_602);
or U7967 (N_7967,N_1696,N_2332);
nand U7968 (N_7968,N_131,N_4058);
and U7969 (N_7969,N_3706,N_2620);
nand U7970 (N_7970,N_1767,N_3546);
nand U7971 (N_7971,N_4076,N_2946);
nand U7972 (N_7972,N_178,N_3183);
nand U7973 (N_7973,N_3078,N_439);
nor U7974 (N_7974,N_1723,N_789);
and U7975 (N_7975,N_4616,N_267);
or U7976 (N_7976,N_2855,N_2013);
nand U7977 (N_7977,N_9,N_234);
nand U7978 (N_7978,N_2106,N_629);
nand U7979 (N_7979,N_1749,N_3402);
nor U7980 (N_7980,N_3232,N_2526);
xor U7981 (N_7981,N_54,N_3582);
or U7982 (N_7982,N_1784,N_1995);
and U7983 (N_7983,N_4622,N_771);
and U7984 (N_7984,N_3052,N_4889);
or U7985 (N_7985,N_838,N_2389);
xnor U7986 (N_7986,N_306,N_4060);
nand U7987 (N_7987,N_1703,N_3173);
or U7988 (N_7988,N_4067,N_4891);
nor U7989 (N_7989,N_1166,N_2643);
and U7990 (N_7990,N_3349,N_2317);
nand U7991 (N_7991,N_1073,N_2985);
xnor U7992 (N_7992,N_419,N_1102);
nor U7993 (N_7993,N_3412,N_2371);
nand U7994 (N_7994,N_768,N_1215);
and U7995 (N_7995,N_2420,N_2969);
nand U7996 (N_7996,N_623,N_3195);
and U7997 (N_7997,N_711,N_907);
or U7998 (N_7998,N_4602,N_3539);
or U7999 (N_7999,N_448,N_4285);
nand U8000 (N_8000,N_3307,N_4587);
and U8001 (N_8001,N_203,N_2008);
xnor U8002 (N_8002,N_3462,N_386);
nor U8003 (N_8003,N_4793,N_4624);
nand U8004 (N_8004,N_1200,N_1838);
nand U8005 (N_8005,N_545,N_4471);
nor U8006 (N_8006,N_1137,N_1468);
nand U8007 (N_8007,N_2473,N_3438);
and U8008 (N_8008,N_908,N_842);
and U8009 (N_8009,N_3215,N_3025);
xnor U8010 (N_8010,N_2904,N_4214);
nand U8011 (N_8011,N_2021,N_3463);
nand U8012 (N_8012,N_2540,N_4067);
and U8013 (N_8013,N_745,N_2260);
and U8014 (N_8014,N_4325,N_1060);
xnor U8015 (N_8015,N_623,N_3388);
nor U8016 (N_8016,N_3440,N_3885);
nor U8017 (N_8017,N_3067,N_1749);
or U8018 (N_8018,N_714,N_4402);
nand U8019 (N_8019,N_4495,N_943);
or U8020 (N_8020,N_3243,N_1412);
nor U8021 (N_8021,N_343,N_3571);
nor U8022 (N_8022,N_2140,N_4321);
xnor U8023 (N_8023,N_4138,N_2921);
nor U8024 (N_8024,N_1046,N_4539);
and U8025 (N_8025,N_4650,N_2429);
or U8026 (N_8026,N_1808,N_2039);
or U8027 (N_8027,N_2769,N_1871);
nand U8028 (N_8028,N_4459,N_1160);
or U8029 (N_8029,N_1030,N_4395);
nand U8030 (N_8030,N_272,N_4661);
nand U8031 (N_8031,N_4240,N_3826);
nand U8032 (N_8032,N_2412,N_3878);
nor U8033 (N_8033,N_4717,N_3983);
xnor U8034 (N_8034,N_473,N_2333);
nand U8035 (N_8035,N_1662,N_2956);
and U8036 (N_8036,N_3167,N_1835);
nand U8037 (N_8037,N_3251,N_1800);
xnor U8038 (N_8038,N_909,N_2313);
or U8039 (N_8039,N_3110,N_849);
nor U8040 (N_8040,N_2819,N_2074);
and U8041 (N_8041,N_2065,N_776);
xor U8042 (N_8042,N_4259,N_1854);
and U8043 (N_8043,N_3808,N_2055);
and U8044 (N_8044,N_538,N_1374);
and U8045 (N_8045,N_529,N_911);
nand U8046 (N_8046,N_601,N_941);
nor U8047 (N_8047,N_4251,N_3845);
nor U8048 (N_8048,N_2392,N_3986);
and U8049 (N_8049,N_3890,N_2011);
nand U8050 (N_8050,N_2565,N_2343);
nand U8051 (N_8051,N_1279,N_3531);
or U8052 (N_8052,N_4042,N_1285);
or U8053 (N_8053,N_2511,N_4988);
nor U8054 (N_8054,N_4062,N_2884);
nor U8055 (N_8055,N_4371,N_429);
nor U8056 (N_8056,N_2906,N_1942);
nand U8057 (N_8057,N_3786,N_3135);
or U8058 (N_8058,N_81,N_4392);
nand U8059 (N_8059,N_3496,N_518);
and U8060 (N_8060,N_1567,N_4708);
and U8061 (N_8061,N_4903,N_3798);
nor U8062 (N_8062,N_4372,N_2786);
nor U8063 (N_8063,N_4187,N_2087);
nor U8064 (N_8064,N_1948,N_3115);
or U8065 (N_8065,N_2523,N_1694);
nand U8066 (N_8066,N_3483,N_1770);
or U8067 (N_8067,N_4322,N_4152);
nand U8068 (N_8068,N_2419,N_883);
xnor U8069 (N_8069,N_2890,N_2259);
or U8070 (N_8070,N_2210,N_4775);
or U8071 (N_8071,N_4816,N_4793);
nor U8072 (N_8072,N_2776,N_4974);
or U8073 (N_8073,N_347,N_1401);
nand U8074 (N_8074,N_3668,N_2270);
or U8075 (N_8075,N_958,N_3409);
xor U8076 (N_8076,N_3727,N_4036);
nor U8077 (N_8077,N_2519,N_430);
xor U8078 (N_8078,N_4368,N_4029);
and U8079 (N_8079,N_707,N_2977);
and U8080 (N_8080,N_3258,N_3438);
and U8081 (N_8081,N_947,N_1019);
and U8082 (N_8082,N_135,N_2389);
nor U8083 (N_8083,N_1317,N_782);
and U8084 (N_8084,N_3812,N_1659);
nor U8085 (N_8085,N_2921,N_647);
nor U8086 (N_8086,N_181,N_2934);
nor U8087 (N_8087,N_3780,N_1374);
nor U8088 (N_8088,N_4184,N_1829);
nand U8089 (N_8089,N_2288,N_2814);
and U8090 (N_8090,N_1334,N_445);
and U8091 (N_8091,N_1945,N_3455);
and U8092 (N_8092,N_4187,N_3913);
nand U8093 (N_8093,N_174,N_4055);
and U8094 (N_8094,N_4813,N_3757);
and U8095 (N_8095,N_91,N_2578);
nor U8096 (N_8096,N_3624,N_2756);
nor U8097 (N_8097,N_3664,N_3705);
nand U8098 (N_8098,N_2786,N_2028);
xnor U8099 (N_8099,N_1206,N_1942);
nor U8100 (N_8100,N_2070,N_1222);
nand U8101 (N_8101,N_4349,N_4696);
nand U8102 (N_8102,N_2993,N_3036);
nand U8103 (N_8103,N_4842,N_4152);
nand U8104 (N_8104,N_4711,N_4524);
or U8105 (N_8105,N_3644,N_121);
and U8106 (N_8106,N_3067,N_2605);
xnor U8107 (N_8107,N_3967,N_4560);
nor U8108 (N_8108,N_3696,N_292);
and U8109 (N_8109,N_3185,N_2737);
or U8110 (N_8110,N_4165,N_4930);
nand U8111 (N_8111,N_1700,N_4155);
xnor U8112 (N_8112,N_1798,N_314);
nor U8113 (N_8113,N_3193,N_2556);
and U8114 (N_8114,N_3814,N_2099);
or U8115 (N_8115,N_2050,N_2525);
nor U8116 (N_8116,N_4797,N_2700);
and U8117 (N_8117,N_2689,N_3024);
nor U8118 (N_8118,N_4758,N_2369);
xnor U8119 (N_8119,N_3054,N_2455);
nand U8120 (N_8120,N_1471,N_1361);
nor U8121 (N_8121,N_424,N_2407);
xor U8122 (N_8122,N_1915,N_3082);
and U8123 (N_8123,N_4397,N_845);
or U8124 (N_8124,N_2174,N_405);
or U8125 (N_8125,N_2631,N_784);
or U8126 (N_8126,N_4680,N_2898);
nand U8127 (N_8127,N_900,N_844);
xor U8128 (N_8128,N_206,N_1315);
nor U8129 (N_8129,N_171,N_1830);
nor U8130 (N_8130,N_93,N_2648);
and U8131 (N_8131,N_1535,N_3916);
nand U8132 (N_8132,N_3367,N_2463);
nand U8133 (N_8133,N_4177,N_823);
or U8134 (N_8134,N_3952,N_3688);
or U8135 (N_8135,N_976,N_3914);
and U8136 (N_8136,N_3358,N_2236);
or U8137 (N_8137,N_2598,N_1819);
nand U8138 (N_8138,N_2770,N_3194);
nand U8139 (N_8139,N_4316,N_1837);
nand U8140 (N_8140,N_3390,N_4768);
or U8141 (N_8141,N_4165,N_4596);
nand U8142 (N_8142,N_2032,N_1036);
nor U8143 (N_8143,N_4468,N_4812);
xnor U8144 (N_8144,N_4063,N_2657);
nand U8145 (N_8145,N_4049,N_1384);
nand U8146 (N_8146,N_4238,N_848);
or U8147 (N_8147,N_1240,N_4518);
nand U8148 (N_8148,N_2186,N_4598);
nor U8149 (N_8149,N_2791,N_4341);
nand U8150 (N_8150,N_1841,N_2998);
or U8151 (N_8151,N_2563,N_2408);
and U8152 (N_8152,N_4331,N_2757);
and U8153 (N_8153,N_1491,N_1596);
nor U8154 (N_8154,N_3189,N_1805);
or U8155 (N_8155,N_2299,N_4634);
and U8156 (N_8156,N_4742,N_3582);
nand U8157 (N_8157,N_2803,N_565);
or U8158 (N_8158,N_3522,N_4584);
or U8159 (N_8159,N_4573,N_3076);
or U8160 (N_8160,N_1211,N_3963);
and U8161 (N_8161,N_2270,N_4518);
nor U8162 (N_8162,N_4185,N_2354);
nand U8163 (N_8163,N_3181,N_3443);
or U8164 (N_8164,N_1826,N_4745);
and U8165 (N_8165,N_3371,N_444);
nor U8166 (N_8166,N_4268,N_3551);
or U8167 (N_8167,N_3693,N_3756);
or U8168 (N_8168,N_4001,N_3904);
or U8169 (N_8169,N_4946,N_4284);
and U8170 (N_8170,N_4431,N_113);
and U8171 (N_8171,N_4424,N_3522);
nor U8172 (N_8172,N_2121,N_4533);
nand U8173 (N_8173,N_22,N_2404);
and U8174 (N_8174,N_51,N_4375);
and U8175 (N_8175,N_1300,N_3401);
and U8176 (N_8176,N_693,N_2877);
and U8177 (N_8177,N_1831,N_970);
nand U8178 (N_8178,N_1790,N_1541);
xor U8179 (N_8179,N_4615,N_3677);
or U8180 (N_8180,N_4787,N_1639);
nor U8181 (N_8181,N_4794,N_4704);
nor U8182 (N_8182,N_3780,N_4659);
nor U8183 (N_8183,N_1744,N_4871);
and U8184 (N_8184,N_695,N_1749);
nor U8185 (N_8185,N_4369,N_3818);
and U8186 (N_8186,N_3713,N_1206);
and U8187 (N_8187,N_462,N_3232);
nand U8188 (N_8188,N_4310,N_3946);
and U8189 (N_8189,N_4882,N_3845);
and U8190 (N_8190,N_521,N_568);
or U8191 (N_8191,N_3725,N_3225);
nand U8192 (N_8192,N_714,N_3555);
xnor U8193 (N_8193,N_4731,N_4377);
or U8194 (N_8194,N_1967,N_3495);
nor U8195 (N_8195,N_3724,N_1343);
nor U8196 (N_8196,N_2254,N_4782);
nand U8197 (N_8197,N_2653,N_3559);
or U8198 (N_8198,N_4274,N_1830);
and U8199 (N_8199,N_4820,N_3191);
and U8200 (N_8200,N_2541,N_2157);
nor U8201 (N_8201,N_618,N_4972);
or U8202 (N_8202,N_3923,N_1472);
nor U8203 (N_8203,N_4821,N_2736);
nor U8204 (N_8204,N_4023,N_1723);
nand U8205 (N_8205,N_2989,N_328);
and U8206 (N_8206,N_3830,N_4198);
nand U8207 (N_8207,N_3464,N_2004);
or U8208 (N_8208,N_4728,N_1777);
nand U8209 (N_8209,N_2211,N_3246);
and U8210 (N_8210,N_2248,N_2681);
xor U8211 (N_8211,N_2244,N_1847);
or U8212 (N_8212,N_4399,N_928);
and U8213 (N_8213,N_1488,N_4161);
or U8214 (N_8214,N_1337,N_1916);
nor U8215 (N_8215,N_2999,N_276);
or U8216 (N_8216,N_2112,N_2330);
xor U8217 (N_8217,N_2794,N_1597);
or U8218 (N_8218,N_1346,N_4154);
nor U8219 (N_8219,N_2797,N_4761);
nor U8220 (N_8220,N_38,N_4425);
nand U8221 (N_8221,N_4147,N_1743);
nor U8222 (N_8222,N_2120,N_252);
nor U8223 (N_8223,N_61,N_3158);
and U8224 (N_8224,N_3009,N_1807);
or U8225 (N_8225,N_1025,N_1380);
or U8226 (N_8226,N_468,N_4106);
xnor U8227 (N_8227,N_1214,N_3366);
or U8228 (N_8228,N_2294,N_80);
or U8229 (N_8229,N_3262,N_2013);
nor U8230 (N_8230,N_1080,N_3152);
or U8231 (N_8231,N_4720,N_2351);
or U8232 (N_8232,N_871,N_3621);
nor U8233 (N_8233,N_2898,N_581);
and U8234 (N_8234,N_241,N_629);
xor U8235 (N_8235,N_2971,N_1628);
and U8236 (N_8236,N_2684,N_3086);
nand U8237 (N_8237,N_1632,N_769);
nand U8238 (N_8238,N_2672,N_4667);
or U8239 (N_8239,N_1178,N_3683);
nor U8240 (N_8240,N_336,N_3379);
nand U8241 (N_8241,N_2611,N_2724);
nand U8242 (N_8242,N_3406,N_1015);
nand U8243 (N_8243,N_1961,N_1733);
and U8244 (N_8244,N_4172,N_291);
nand U8245 (N_8245,N_606,N_198);
nor U8246 (N_8246,N_2883,N_4043);
and U8247 (N_8247,N_3919,N_3262);
nor U8248 (N_8248,N_1446,N_3405);
xnor U8249 (N_8249,N_806,N_518);
xor U8250 (N_8250,N_2371,N_3630);
and U8251 (N_8251,N_3702,N_743);
nand U8252 (N_8252,N_577,N_4182);
or U8253 (N_8253,N_4198,N_3186);
nor U8254 (N_8254,N_2031,N_4226);
or U8255 (N_8255,N_298,N_1412);
nand U8256 (N_8256,N_2811,N_2096);
and U8257 (N_8257,N_733,N_3940);
or U8258 (N_8258,N_740,N_3973);
nor U8259 (N_8259,N_4437,N_1652);
or U8260 (N_8260,N_4796,N_4469);
or U8261 (N_8261,N_4846,N_4674);
or U8262 (N_8262,N_2263,N_4348);
xor U8263 (N_8263,N_794,N_541);
nand U8264 (N_8264,N_1974,N_572);
and U8265 (N_8265,N_4696,N_2658);
nand U8266 (N_8266,N_3890,N_1317);
and U8267 (N_8267,N_2891,N_2288);
and U8268 (N_8268,N_1683,N_3182);
or U8269 (N_8269,N_4248,N_3423);
nor U8270 (N_8270,N_4923,N_593);
nand U8271 (N_8271,N_1772,N_782);
and U8272 (N_8272,N_2040,N_1290);
nor U8273 (N_8273,N_2811,N_4321);
nor U8274 (N_8274,N_1492,N_3240);
nor U8275 (N_8275,N_2143,N_2983);
xnor U8276 (N_8276,N_3826,N_4263);
or U8277 (N_8277,N_3789,N_3582);
and U8278 (N_8278,N_2158,N_1423);
nand U8279 (N_8279,N_2377,N_2648);
nand U8280 (N_8280,N_1165,N_735);
nor U8281 (N_8281,N_4074,N_2420);
nand U8282 (N_8282,N_4237,N_1082);
and U8283 (N_8283,N_4140,N_1473);
xor U8284 (N_8284,N_4823,N_2518);
or U8285 (N_8285,N_4325,N_4715);
and U8286 (N_8286,N_4561,N_2033);
or U8287 (N_8287,N_525,N_3840);
nand U8288 (N_8288,N_1849,N_1527);
nand U8289 (N_8289,N_2243,N_4972);
or U8290 (N_8290,N_4336,N_4899);
nand U8291 (N_8291,N_4538,N_3234);
nor U8292 (N_8292,N_4277,N_664);
and U8293 (N_8293,N_4249,N_1756);
and U8294 (N_8294,N_2389,N_500);
or U8295 (N_8295,N_278,N_3236);
or U8296 (N_8296,N_1433,N_3487);
nand U8297 (N_8297,N_1650,N_3420);
and U8298 (N_8298,N_552,N_185);
nand U8299 (N_8299,N_4707,N_123);
and U8300 (N_8300,N_4801,N_4365);
and U8301 (N_8301,N_924,N_4844);
or U8302 (N_8302,N_4871,N_4433);
nor U8303 (N_8303,N_185,N_3890);
or U8304 (N_8304,N_1940,N_935);
or U8305 (N_8305,N_2018,N_3385);
and U8306 (N_8306,N_4872,N_1702);
and U8307 (N_8307,N_352,N_1053);
or U8308 (N_8308,N_1032,N_4094);
or U8309 (N_8309,N_4297,N_175);
nand U8310 (N_8310,N_1971,N_3632);
nand U8311 (N_8311,N_321,N_3794);
and U8312 (N_8312,N_899,N_755);
and U8313 (N_8313,N_4640,N_670);
and U8314 (N_8314,N_3633,N_1513);
and U8315 (N_8315,N_2137,N_271);
nand U8316 (N_8316,N_3848,N_2968);
and U8317 (N_8317,N_2581,N_2137);
xnor U8318 (N_8318,N_718,N_1976);
or U8319 (N_8319,N_1980,N_2754);
and U8320 (N_8320,N_4246,N_2300);
xor U8321 (N_8321,N_4187,N_1544);
or U8322 (N_8322,N_813,N_1039);
and U8323 (N_8323,N_1558,N_0);
nor U8324 (N_8324,N_4990,N_67);
nor U8325 (N_8325,N_1424,N_2116);
or U8326 (N_8326,N_4564,N_2306);
nor U8327 (N_8327,N_3339,N_4063);
nor U8328 (N_8328,N_3596,N_2815);
or U8329 (N_8329,N_251,N_304);
and U8330 (N_8330,N_3911,N_3691);
xor U8331 (N_8331,N_2462,N_128);
nand U8332 (N_8332,N_1095,N_4085);
nand U8333 (N_8333,N_2644,N_2514);
nor U8334 (N_8334,N_2681,N_721);
or U8335 (N_8335,N_195,N_442);
or U8336 (N_8336,N_450,N_2532);
and U8337 (N_8337,N_342,N_147);
nor U8338 (N_8338,N_757,N_3893);
nand U8339 (N_8339,N_1241,N_1534);
nor U8340 (N_8340,N_4796,N_1062);
and U8341 (N_8341,N_552,N_4578);
and U8342 (N_8342,N_4241,N_59);
nor U8343 (N_8343,N_4934,N_1841);
nor U8344 (N_8344,N_4679,N_3947);
or U8345 (N_8345,N_3618,N_4889);
and U8346 (N_8346,N_3906,N_2888);
nor U8347 (N_8347,N_3905,N_3553);
xor U8348 (N_8348,N_2806,N_2866);
nor U8349 (N_8349,N_3268,N_1823);
and U8350 (N_8350,N_938,N_4051);
nand U8351 (N_8351,N_397,N_1369);
xor U8352 (N_8352,N_3731,N_4718);
nand U8353 (N_8353,N_993,N_1608);
nor U8354 (N_8354,N_1088,N_4874);
nor U8355 (N_8355,N_1058,N_284);
or U8356 (N_8356,N_146,N_2630);
nor U8357 (N_8357,N_4596,N_642);
nand U8358 (N_8358,N_1493,N_268);
nand U8359 (N_8359,N_3483,N_3413);
or U8360 (N_8360,N_2678,N_3250);
or U8361 (N_8361,N_4878,N_806);
nor U8362 (N_8362,N_1787,N_3507);
xnor U8363 (N_8363,N_3550,N_3768);
or U8364 (N_8364,N_2355,N_1321);
nor U8365 (N_8365,N_1006,N_2158);
nand U8366 (N_8366,N_2044,N_4750);
nor U8367 (N_8367,N_2384,N_4893);
and U8368 (N_8368,N_684,N_3643);
nand U8369 (N_8369,N_2489,N_3310);
nand U8370 (N_8370,N_3287,N_1261);
xor U8371 (N_8371,N_4194,N_3033);
or U8372 (N_8372,N_327,N_1305);
nor U8373 (N_8373,N_771,N_4548);
nor U8374 (N_8374,N_1755,N_3759);
nand U8375 (N_8375,N_1753,N_225);
and U8376 (N_8376,N_478,N_1914);
or U8377 (N_8377,N_4309,N_1580);
nand U8378 (N_8378,N_4393,N_1731);
or U8379 (N_8379,N_2986,N_1064);
xnor U8380 (N_8380,N_4542,N_544);
nand U8381 (N_8381,N_680,N_4163);
nand U8382 (N_8382,N_3545,N_1944);
xor U8383 (N_8383,N_1675,N_2485);
xnor U8384 (N_8384,N_4882,N_4878);
nor U8385 (N_8385,N_723,N_2456);
or U8386 (N_8386,N_832,N_1016);
nor U8387 (N_8387,N_3371,N_2026);
nand U8388 (N_8388,N_2172,N_1143);
and U8389 (N_8389,N_2495,N_1725);
nor U8390 (N_8390,N_3269,N_2420);
and U8391 (N_8391,N_559,N_4520);
and U8392 (N_8392,N_2833,N_813);
and U8393 (N_8393,N_3533,N_3244);
and U8394 (N_8394,N_4371,N_1570);
nand U8395 (N_8395,N_1574,N_4661);
xor U8396 (N_8396,N_3252,N_1699);
nand U8397 (N_8397,N_251,N_3175);
or U8398 (N_8398,N_3964,N_3940);
nand U8399 (N_8399,N_2299,N_4789);
nor U8400 (N_8400,N_3896,N_1006);
nand U8401 (N_8401,N_2324,N_934);
or U8402 (N_8402,N_4524,N_2371);
and U8403 (N_8403,N_4203,N_2555);
nand U8404 (N_8404,N_3387,N_4767);
or U8405 (N_8405,N_1407,N_2923);
nor U8406 (N_8406,N_3256,N_4655);
nand U8407 (N_8407,N_4647,N_3057);
nor U8408 (N_8408,N_4629,N_3183);
or U8409 (N_8409,N_1327,N_1302);
or U8410 (N_8410,N_261,N_1423);
or U8411 (N_8411,N_3479,N_3390);
xnor U8412 (N_8412,N_4321,N_2881);
nor U8413 (N_8413,N_3998,N_3694);
or U8414 (N_8414,N_2836,N_4610);
xor U8415 (N_8415,N_4757,N_987);
nand U8416 (N_8416,N_3812,N_951);
nor U8417 (N_8417,N_4461,N_2912);
and U8418 (N_8418,N_1608,N_692);
and U8419 (N_8419,N_390,N_3120);
xor U8420 (N_8420,N_2171,N_4323);
or U8421 (N_8421,N_1934,N_4817);
nor U8422 (N_8422,N_463,N_3606);
or U8423 (N_8423,N_1168,N_4283);
nand U8424 (N_8424,N_1532,N_3379);
or U8425 (N_8425,N_1054,N_4742);
nand U8426 (N_8426,N_1746,N_3929);
and U8427 (N_8427,N_2189,N_3056);
or U8428 (N_8428,N_1208,N_4980);
nor U8429 (N_8429,N_370,N_4321);
nand U8430 (N_8430,N_435,N_1072);
xnor U8431 (N_8431,N_272,N_3536);
nand U8432 (N_8432,N_1961,N_4737);
xnor U8433 (N_8433,N_3302,N_942);
nor U8434 (N_8434,N_4527,N_4593);
nor U8435 (N_8435,N_862,N_4584);
nand U8436 (N_8436,N_1243,N_1448);
or U8437 (N_8437,N_3968,N_1347);
nand U8438 (N_8438,N_2314,N_3400);
xnor U8439 (N_8439,N_2153,N_4129);
nand U8440 (N_8440,N_549,N_4837);
nand U8441 (N_8441,N_579,N_3287);
or U8442 (N_8442,N_248,N_3782);
nand U8443 (N_8443,N_3670,N_3039);
or U8444 (N_8444,N_3448,N_137);
xnor U8445 (N_8445,N_4290,N_2049);
nand U8446 (N_8446,N_4160,N_121);
nand U8447 (N_8447,N_1068,N_3015);
and U8448 (N_8448,N_4300,N_2007);
nor U8449 (N_8449,N_803,N_4102);
nand U8450 (N_8450,N_4287,N_950);
or U8451 (N_8451,N_1542,N_2466);
or U8452 (N_8452,N_2035,N_3931);
nand U8453 (N_8453,N_1636,N_4763);
nor U8454 (N_8454,N_2616,N_260);
and U8455 (N_8455,N_1402,N_1351);
nor U8456 (N_8456,N_4091,N_4408);
and U8457 (N_8457,N_1967,N_2239);
xnor U8458 (N_8458,N_971,N_4830);
nor U8459 (N_8459,N_2575,N_4882);
nor U8460 (N_8460,N_4123,N_2030);
or U8461 (N_8461,N_3512,N_3909);
or U8462 (N_8462,N_4163,N_1915);
nand U8463 (N_8463,N_281,N_4502);
and U8464 (N_8464,N_796,N_1337);
xor U8465 (N_8465,N_4578,N_3097);
nand U8466 (N_8466,N_1707,N_3786);
and U8467 (N_8467,N_3361,N_4015);
and U8468 (N_8468,N_1661,N_3541);
nor U8469 (N_8469,N_2747,N_4471);
nor U8470 (N_8470,N_3281,N_3466);
and U8471 (N_8471,N_4453,N_3292);
nor U8472 (N_8472,N_4755,N_4584);
nand U8473 (N_8473,N_993,N_2582);
xnor U8474 (N_8474,N_2463,N_8);
nand U8475 (N_8475,N_1653,N_4373);
or U8476 (N_8476,N_3252,N_4608);
or U8477 (N_8477,N_4927,N_1834);
or U8478 (N_8478,N_1976,N_2342);
nand U8479 (N_8479,N_4276,N_3115);
xor U8480 (N_8480,N_2680,N_2884);
and U8481 (N_8481,N_4770,N_3006);
and U8482 (N_8482,N_3844,N_2378);
or U8483 (N_8483,N_1692,N_3739);
nor U8484 (N_8484,N_2332,N_1158);
nor U8485 (N_8485,N_3748,N_2629);
or U8486 (N_8486,N_3804,N_4939);
xnor U8487 (N_8487,N_1711,N_2664);
nand U8488 (N_8488,N_4600,N_4234);
and U8489 (N_8489,N_4459,N_3466);
or U8490 (N_8490,N_849,N_2521);
or U8491 (N_8491,N_2191,N_1409);
nor U8492 (N_8492,N_702,N_3388);
xnor U8493 (N_8493,N_4289,N_971);
xor U8494 (N_8494,N_1269,N_872);
or U8495 (N_8495,N_3404,N_1383);
and U8496 (N_8496,N_2179,N_2499);
and U8497 (N_8497,N_1781,N_2817);
and U8498 (N_8498,N_642,N_931);
or U8499 (N_8499,N_1995,N_4645);
and U8500 (N_8500,N_156,N_4729);
xor U8501 (N_8501,N_3220,N_3612);
nand U8502 (N_8502,N_4157,N_1849);
nor U8503 (N_8503,N_1795,N_835);
nor U8504 (N_8504,N_3789,N_787);
xnor U8505 (N_8505,N_4535,N_4412);
nand U8506 (N_8506,N_73,N_2280);
nor U8507 (N_8507,N_2656,N_265);
or U8508 (N_8508,N_1538,N_3180);
nor U8509 (N_8509,N_877,N_3880);
nor U8510 (N_8510,N_2003,N_512);
or U8511 (N_8511,N_1122,N_3233);
or U8512 (N_8512,N_2909,N_2370);
nand U8513 (N_8513,N_3604,N_829);
nor U8514 (N_8514,N_2933,N_3471);
nand U8515 (N_8515,N_4494,N_4146);
nand U8516 (N_8516,N_729,N_1182);
nor U8517 (N_8517,N_2294,N_1895);
and U8518 (N_8518,N_244,N_3298);
nand U8519 (N_8519,N_4904,N_118);
and U8520 (N_8520,N_3979,N_1846);
nand U8521 (N_8521,N_3502,N_4303);
nor U8522 (N_8522,N_4338,N_2500);
nor U8523 (N_8523,N_2493,N_4178);
and U8524 (N_8524,N_3575,N_1867);
nand U8525 (N_8525,N_2387,N_1628);
and U8526 (N_8526,N_899,N_4288);
and U8527 (N_8527,N_794,N_690);
nor U8528 (N_8528,N_2278,N_3340);
nand U8529 (N_8529,N_1342,N_2495);
or U8530 (N_8530,N_518,N_266);
nor U8531 (N_8531,N_1307,N_1443);
or U8532 (N_8532,N_2561,N_1821);
and U8533 (N_8533,N_3699,N_3938);
and U8534 (N_8534,N_1603,N_1103);
nor U8535 (N_8535,N_4305,N_3652);
or U8536 (N_8536,N_2824,N_2744);
or U8537 (N_8537,N_763,N_497);
or U8538 (N_8538,N_784,N_4656);
nand U8539 (N_8539,N_1690,N_3000);
or U8540 (N_8540,N_2296,N_4817);
nand U8541 (N_8541,N_1625,N_2017);
or U8542 (N_8542,N_4108,N_4011);
nor U8543 (N_8543,N_957,N_4248);
nand U8544 (N_8544,N_2169,N_3771);
xnor U8545 (N_8545,N_3828,N_2925);
or U8546 (N_8546,N_3997,N_3397);
nor U8547 (N_8547,N_3809,N_3981);
nand U8548 (N_8548,N_3074,N_2963);
xor U8549 (N_8549,N_1564,N_1340);
nor U8550 (N_8550,N_3597,N_870);
and U8551 (N_8551,N_2869,N_2664);
nand U8552 (N_8552,N_390,N_401);
and U8553 (N_8553,N_1493,N_137);
or U8554 (N_8554,N_1908,N_1689);
nor U8555 (N_8555,N_2950,N_590);
nand U8556 (N_8556,N_4411,N_4034);
nand U8557 (N_8557,N_1924,N_200);
nor U8558 (N_8558,N_2812,N_4365);
nand U8559 (N_8559,N_4447,N_2484);
nor U8560 (N_8560,N_182,N_1190);
nor U8561 (N_8561,N_3661,N_1800);
or U8562 (N_8562,N_3745,N_3655);
or U8563 (N_8563,N_3173,N_2186);
nand U8564 (N_8564,N_3661,N_2477);
nand U8565 (N_8565,N_3476,N_4215);
nor U8566 (N_8566,N_2862,N_2381);
and U8567 (N_8567,N_4017,N_1146);
and U8568 (N_8568,N_2346,N_2516);
xor U8569 (N_8569,N_4750,N_969);
nand U8570 (N_8570,N_3541,N_2337);
nand U8571 (N_8571,N_1842,N_2849);
or U8572 (N_8572,N_4252,N_2738);
nor U8573 (N_8573,N_3148,N_3887);
or U8574 (N_8574,N_4718,N_1237);
and U8575 (N_8575,N_675,N_333);
nand U8576 (N_8576,N_3723,N_1117);
nand U8577 (N_8577,N_3346,N_3194);
nand U8578 (N_8578,N_1295,N_2996);
and U8579 (N_8579,N_2747,N_3057);
and U8580 (N_8580,N_3741,N_4194);
nand U8581 (N_8581,N_1868,N_2202);
or U8582 (N_8582,N_4328,N_4588);
nor U8583 (N_8583,N_2329,N_1585);
nor U8584 (N_8584,N_3566,N_165);
and U8585 (N_8585,N_1938,N_476);
nor U8586 (N_8586,N_4448,N_2929);
nand U8587 (N_8587,N_616,N_129);
nor U8588 (N_8588,N_3029,N_1700);
nor U8589 (N_8589,N_10,N_2102);
or U8590 (N_8590,N_2926,N_2552);
nand U8591 (N_8591,N_3203,N_4695);
nand U8592 (N_8592,N_3191,N_2348);
and U8593 (N_8593,N_56,N_3342);
or U8594 (N_8594,N_3230,N_2586);
and U8595 (N_8595,N_3802,N_1933);
and U8596 (N_8596,N_121,N_3642);
nand U8597 (N_8597,N_203,N_4711);
nand U8598 (N_8598,N_2423,N_1938);
or U8599 (N_8599,N_31,N_4705);
and U8600 (N_8600,N_249,N_2383);
nor U8601 (N_8601,N_2504,N_2391);
nand U8602 (N_8602,N_137,N_778);
nand U8603 (N_8603,N_4841,N_1532);
or U8604 (N_8604,N_696,N_4644);
nand U8605 (N_8605,N_3817,N_3307);
nand U8606 (N_8606,N_3595,N_2228);
xnor U8607 (N_8607,N_178,N_603);
nand U8608 (N_8608,N_214,N_2533);
nor U8609 (N_8609,N_3802,N_4596);
nand U8610 (N_8610,N_2571,N_3442);
or U8611 (N_8611,N_1757,N_2717);
xor U8612 (N_8612,N_1435,N_2124);
nor U8613 (N_8613,N_1363,N_4192);
nor U8614 (N_8614,N_2326,N_1530);
nor U8615 (N_8615,N_3087,N_2704);
or U8616 (N_8616,N_2485,N_621);
nand U8617 (N_8617,N_3107,N_4140);
nor U8618 (N_8618,N_1476,N_1370);
nor U8619 (N_8619,N_948,N_2717);
nor U8620 (N_8620,N_1470,N_2798);
nand U8621 (N_8621,N_122,N_1621);
and U8622 (N_8622,N_3412,N_751);
or U8623 (N_8623,N_3070,N_4000);
nand U8624 (N_8624,N_2789,N_3870);
or U8625 (N_8625,N_1715,N_1122);
xnor U8626 (N_8626,N_1443,N_2208);
nor U8627 (N_8627,N_549,N_98);
nand U8628 (N_8628,N_486,N_833);
and U8629 (N_8629,N_334,N_3698);
and U8630 (N_8630,N_3292,N_4742);
nor U8631 (N_8631,N_1998,N_3640);
xnor U8632 (N_8632,N_4894,N_2131);
or U8633 (N_8633,N_4314,N_409);
or U8634 (N_8634,N_2978,N_799);
nor U8635 (N_8635,N_1439,N_2586);
and U8636 (N_8636,N_4449,N_2063);
and U8637 (N_8637,N_3585,N_3947);
and U8638 (N_8638,N_1024,N_4666);
nand U8639 (N_8639,N_1263,N_2099);
xnor U8640 (N_8640,N_2108,N_1696);
and U8641 (N_8641,N_1311,N_3581);
and U8642 (N_8642,N_2544,N_1264);
or U8643 (N_8643,N_3505,N_1653);
nand U8644 (N_8644,N_3761,N_2239);
nor U8645 (N_8645,N_3635,N_4574);
or U8646 (N_8646,N_2160,N_2616);
nand U8647 (N_8647,N_2463,N_3803);
nand U8648 (N_8648,N_4805,N_4696);
or U8649 (N_8649,N_3999,N_2067);
nand U8650 (N_8650,N_2262,N_1306);
nand U8651 (N_8651,N_4046,N_626);
nor U8652 (N_8652,N_544,N_1878);
nand U8653 (N_8653,N_786,N_2790);
or U8654 (N_8654,N_4343,N_2884);
xor U8655 (N_8655,N_4496,N_189);
or U8656 (N_8656,N_3427,N_4029);
and U8657 (N_8657,N_2408,N_272);
or U8658 (N_8658,N_3568,N_1880);
nand U8659 (N_8659,N_3765,N_4803);
and U8660 (N_8660,N_3841,N_1572);
nand U8661 (N_8661,N_2619,N_103);
and U8662 (N_8662,N_2141,N_3803);
or U8663 (N_8663,N_3348,N_1574);
or U8664 (N_8664,N_2453,N_2476);
nand U8665 (N_8665,N_2418,N_1410);
xnor U8666 (N_8666,N_3537,N_847);
nor U8667 (N_8667,N_2913,N_731);
nor U8668 (N_8668,N_4126,N_1050);
and U8669 (N_8669,N_18,N_893);
nor U8670 (N_8670,N_2419,N_298);
nand U8671 (N_8671,N_3315,N_4350);
nand U8672 (N_8672,N_1296,N_3586);
and U8673 (N_8673,N_1243,N_4365);
and U8674 (N_8674,N_639,N_4439);
or U8675 (N_8675,N_1102,N_2551);
xor U8676 (N_8676,N_1696,N_3735);
nor U8677 (N_8677,N_3991,N_3507);
nand U8678 (N_8678,N_2755,N_1705);
and U8679 (N_8679,N_2376,N_2932);
nor U8680 (N_8680,N_945,N_2858);
and U8681 (N_8681,N_2022,N_2569);
or U8682 (N_8682,N_3081,N_3961);
nor U8683 (N_8683,N_4158,N_1671);
nor U8684 (N_8684,N_1235,N_3945);
xor U8685 (N_8685,N_2870,N_260);
and U8686 (N_8686,N_1174,N_603);
and U8687 (N_8687,N_732,N_3396);
nor U8688 (N_8688,N_1393,N_318);
nand U8689 (N_8689,N_426,N_1198);
and U8690 (N_8690,N_376,N_917);
or U8691 (N_8691,N_4749,N_4773);
and U8692 (N_8692,N_1673,N_4124);
or U8693 (N_8693,N_138,N_4368);
nor U8694 (N_8694,N_232,N_2931);
nand U8695 (N_8695,N_3797,N_4404);
and U8696 (N_8696,N_3114,N_2017);
nand U8697 (N_8697,N_3862,N_4887);
and U8698 (N_8698,N_3452,N_4097);
nand U8699 (N_8699,N_4463,N_4618);
nand U8700 (N_8700,N_3029,N_3432);
nor U8701 (N_8701,N_3331,N_958);
or U8702 (N_8702,N_4702,N_4291);
xnor U8703 (N_8703,N_4254,N_1405);
nand U8704 (N_8704,N_4363,N_1913);
and U8705 (N_8705,N_4435,N_3464);
and U8706 (N_8706,N_4177,N_307);
and U8707 (N_8707,N_1825,N_4854);
or U8708 (N_8708,N_2560,N_339);
nor U8709 (N_8709,N_771,N_4275);
nor U8710 (N_8710,N_1816,N_4458);
nand U8711 (N_8711,N_2825,N_3334);
xor U8712 (N_8712,N_3247,N_3883);
nand U8713 (N_8713,N_3308,N_3068);
or U8714 (N_8714,N_2402,N_3691);
nor U8715 (N_8715,N_2449,N_4388);
nor U8716 (N_8716,N_3879,N_29);
nand U8717 (N_8717,N_4808,N_3616);
nand U8718 (N_8718,N_4037,N_386);
or U8719 (N_8719,N_3835,N_4649);
nand U8720 (N_8720,N_3317,N_606);
and U8721 (N_8721,N_356,N_3587);
nor U8722 (N_8722,N_591,N_4334);
nor U8723 (N_8723,N_2548,N_550);
nand U8724 (N_8724,N_3989,N_1324);
xnor U8725 (N_8725,N_4913,N_1702);
and U8726 (N_8726,N_3484,N_3732);
xor U8727 (N_8727,N_2791,N_2715);
nand U8728 (N_8728,N_4910,N_702);
or U8729 (N_8729,N_2913,N_444);
and U8730 (N_8730,N_4117,N_4684);
or U8731 (N_8731,N_1819,N_4981);
xor U8732 (N_8732,N_1953,N_985);
or U8733 (N_8733,N_3717,N_4006);
or U8734 (N_8734,N_4008,N_3126);
nor U8735 (N_8735,N_929,N_3951);
or U8736 (N_8736,N_3600,N_1695);
or U8737 (N_8737,N_2848,N_2589);
or U8738 (N_8738,N_826,N_4400);
nand U8739 (N_8739,N_4434,N_1816);
and U8740 (N_8740,N_511,N_4803);
nand U8741 (N_8741,N_4172,N_4791);
xnor U8742 (N_8742,N_186,N_2151);
nor U8743 (N_8743,N_1533,N_2429);
nand U8744 (N_8744,N_2722,N_2383);
or U8745 (N_8745,N_4899,N_3611);
nand U8746 (N_8746,N_3187,N_878);
and U8747 (N_8747,N_1793,N_4370);
and U8748 (N_8748,N_1559,N_1604);
nor U8749 (N_8749,N_1571,N_1390);
nor U8750 (N_8750,N_1459,N_2952);
nand U8751 (N_8751,N_1745,N_1598);
nand U8752 (N_8752,N_260,N_43);
and U8753 (N_8753,N_951,N_3732);
nor U8754 (N_8754,N_4204,N_643);
nand U8755 (N_8755,N_3152,N_215);
nand U8756 (N_8756,N_2496,N_1661);
nand U8757 (N_8757,N_4416,N_988);
and U8758 (N_8758,N_2928,N_4608);
or U8759 (N_8759,N_757,N_612);
nand U8760 (N_8760,N_3422,N_2329);
xnor U8761 (N_8761,N_4534,N_1055);
xnor U8762 (N_8762,N_1687,N_2981);
nor U8763 (N_8763,N_610,N_4041);
nand U8764 (N_8764,N_2103,N_2631);
xnor U8765 (N_8765,N_4002,N_2777);
nor U8766 (N_8766,N_304,N_918);
and U8767 (N_8767,N_4813,N_3239);
nor U8768 (N_8768,N_4449,N_388);
or U8769 (N_8769,N_1829,N_2722);
nand U8770 (N_8770,N_1178,N_1057);
or U8771 (N_8771,N_2264,N_1504);
xor U8772 (N_8772,N_2149,N_765);
xnor U8773 (N_8773,N_2201,N_650);
and U8774 (N_8774,N_4126,N_3550);
and U8775 (N_8775,N_985,N_4067);
or U8776 (N_8776,N_1271,N_4072);
or U8777 (N_8777,N_1336,N_1881);
and U8778 (N_8778,N_1362,N_2354);
and U8779 (N_8779,N_3709,N_2475);
xor U8780 (N_8780,N_4318,N_158);
and U8781 (N_8781,N_4953,N_1780);
and U8782 (N_8782,N_281,N_2404);
nor U8783 (N_8783,N_4406,N_1705);
or U8784 (N_8784,N_2239,N_486);
nor U8785 (N_8785,N_3149,N_2077);
nor U8786 (N_8786,N_22,N_2653);
or U8787 (N_8787,N_902,N_2226);
or U8788 (N_8788,N_1047,N_3536);
nand U8789 (N_8789,N_4662,N_2069);
nor U8790 (N_8790,N_2190,N_630);
or U8791 (N_8791,N_1354,N_476);
or U8792 (N_8792,N_3394,N_1815);
nand U8793 (N_8793,N_4112,N_1343);
or U8794 (N_8794,N_2985,N_3419);
or U8795 (N_8795,N_542,N_3692);
nor U8796 (N_8796,N_1527,N_3861);
and U8797 (N_8797,N_4044,N_2123);
and U8798 (N_8798,N_98,N_702);
nand U8799 (N_8799,N_2067,N_2715);
or U8800 (N_8800,N_1839,N_4783);
and U8801 (N_8801,N_2547,N_3530);
nor U8802 (N_8802,N_1715,N_1115);
xor U8803 (N_8803,N_3974,N_2276);
or U8804 (N_8804,N_2636,N_347);
or U8805 (N_8805,N_4454,N_43);
and U8806 (N_8806,N_3849,N_1533);
and U8807 (N_8807,N_595,N_2573);
xor U8808 (N_8808,N_2537,N_2937);
xor U8809 (N_8809,N_1687,N_4290);
nor U8810 (N_8810,N_2079,N_3484);
or U8811 (N_8811,N_3790,N_915);
nor U8812 (N_8812,N_2548,N_2127);
or U8813 (N_8813,N_3204,N_1217);
nor U8814 (N_8814,N_1525,N_4075);
nand U8815 (N_8815,N_3856,N_1782);
nor U8816 (N_8816,N_4203,N_4280);
or U8817 (N_8817,N_4375,N_1649);
and U8818 (N_8818,N_686,N_2120);
or U8819 (N_8819,N_1515,N_3902);
or U8820 (N_8820,N_3090,N_1566);
xor U8821 (N_8821,N_3123,N_4355);
nand U8822 (N_8822,N_2916,N_236);
xor U8823 (N_8823,N_611,N_1069);
or U8824 (N_8824,N_1446,N_3773);
or U8825 (N_8825,N_690,N_2072);
nand U8826 (N_8826,N_3915,N_4446);
and U8827 (N_8827,N_411,N_2173);
or U8828 (N_8828,N_2925,N_2982);
xor U8829 (N_8829,N_446,N_3429);
and U8830 (N_8830,N_2458,N_3273);
nor U8831 (N_8831,N_1711,N_1072);
or U8832 (N_8832,N_895,N_4646);
and U8833 (N_8833,N_2650,N_3525);
or U8834 (N_8834,N_1724,N_733);
xnor U8835 (N_8835,N_3719,N_4931);
and U8836 (N_8836,N_1118,N_4864);
nand U8837 (N_8837,N_1946,N_4225);
nand U8838 (N_8838,N_4644,N_2250);
xnor U8839 (N_8839,N_229,N_111);
and U8840 (N_8840,N_2943,N_3706);
and U8841 (N_8841,N_4085,N_1794);
nor U8842 (N_8842,N_3933,N_263);
nand U8843 (N_8843,N_1524,N_4956);
nand U8844 (N_8844,N_3334,N_1842);
nand U8845 (N_8845,N_2020,N_2578);
nand U8846 (N_8846,N_2023,N_4688);
or U8847 (N_8847,N_1221,N_3276);
nor U8848 (N_8848,N_2798,N_128);
nand U8849 (N_8849,N_841,N_3054);
nand U8850 (N_8850,N_2253,N_4703);
nand U8851 (N_8851,N_3704,N_4827);
xnor U8852 (N_8852,N_869,N_3610);
and U8853 (N_8853,N_4328,N_3041);
or U8854 (N_8854,N_2348,N_2170);
nand U8855 (N_8855,N_4105,N_4621);
or U8856 (N_8856,N_4233,N_2998);
or U8857 (N_8857,N_4445,N_2439);
and U8858 (N_8858,N_1897,N_3014);
and U8859 (N_8859,N_3115,N_3415);
xnor U8860 (N_8860,N_4542,N_1389);
nor U8861 (N_8861,N_3365,N_1455);
nand U8862 (N_8862,N_414,N_3870);
nand U8863 (N_8863,N_828,N_4032);
nand U8864 (N_8864,N_3967,N_1624);
or U8865 (N_8865,N_4550,N_512);
nor U8866 (N_8866,N_1804,N_3466);
and U8867 (N_8867,N_897,N_3381);
nor U8868 (N_8868,N_1536,N_1327);
and U8869 (N_8869,N_2211,N_996);
and U8870 (N_8870,N_3967,N_1907);
nand U8871 (N_8871,N_1229,N_4989);
nor U8872 (N_8872,N_675,N_456);
nand U8873 (N_8873,N_2489,N_1841);
or U8874 (N_8874,N_4767,N_3797);
nand U8875 (N_8875,N_1031,N_2149);
or U8876 (N_8876,N_2227,N_4130);
and U8877 (N_8877,N_3319,N_1291);
nand U8878 (N_8878,N_358,N_4789);
or U8879 (N_8879,N_872,N_4968);
and U8880 (N_8880,N_2695,N_3070);
nor U8881 (N_8881,N_2356,N_2048);
and U8882 (N_8882,N_1698,N_3636);
xnor U8883 (N_8883,N_4477,N_2377);
nand U8884 (N_8884,N_1176,N_4408);
or U8885 (N_8885,N_2175,N_4977);
nor U8886 (N_8886,N_1269,N_2496);
nand U8887 (N_8887,N_2384,N_436);
or U8888 (N_8888,N_3704,N_4084);
nand U8889 (N_8889,N_591,N_1261);
xor U8890 (N_8890,N_4441,N_2540);
or U8891 (N_8891,N_2031,N_1023);
and U8892 (N_8892,N_4172,N_2569);
or U8893 (N_8893,N_707,N_4497);
and U8894 (N_8894,N_2427,N_1145);
and U8895 (N_8895,N_1407,N_1107);
or U8896 (N_8896,N_1239,N_612);
nand U8897 (N_8897,N_4314,N_2521);
and U8898 (N_8898,N_1500,N_4743);
nand U8899 (N_8899,N_3186,N_1988);
nor U8900 (N_8900,N_2623,N_4761);
and U8901 (N_8901,N_2344,N_3823);
xor U8902 (N_8902,N_436,N_2282);
or U8903 (N_8903,N_2486,N_3139);
nand U8904 (N_8904,N_510,N_4348);
or U8905 (N_8905,N_3489,N_1087);
nor U8906 (N_8906,N_3751,N_4222);
or U8907 (N_8907,N_2894,N_4759);
nor U8908 (N_8908,N_3532,N_4793);
or U8909 (N_8909,N_2788,N_1734);
or U8910 (N_8910,N_4043,N_681);
nor U8911 (N_8911,N_842,N_3864);
nand U8912 (N_8912,N_2123,N_3182);
nand U8913 (N_8913,N_2810,N_3607);
or U8914 (N_8914,N_4504,N_2665);
and U8915 (N_8915,N_230,N_1626);
nor U8916 (N_8916,N_807,N_3937);
and U8917 (N_8917,N_1201,N_3337);
and U8918 (N_8918,N_2286,N_838);
or U8919 (N_8919,N_4429,N_4703);
nand U8920 (N_8920,N_2563,N_2317);
or U8921 (N_8921,N_4777,N_4165);
nand U8922 (N_8922,N_4870,N_2649);
or U8923 (N_8923,N_928,N_4435);
xnor U8924 (N_8924,N_4028,N_273);
nand U8925 (N_8925,N_2996,N_3783);
nand U8926 (N_8926,N_7,N_3272);
and U8927 (N_8927,N_1716,N_1730);
and U8928 (N_8928,N_4767,N_3042);
and U8929 (N_8929,N_2051,N_4818);
and U8930 (N_8930,N_1708,N_2015);
nor U8931 (N_8931,N_2703,N_122);
nand U8932 (N_8932,N_2111,N_2001);
nor U8933 (N_8933,N_4054,N_2129);
nor U8934 (N_8934,N_4943,N_3374);
xor U8935 (N_8935,N_4800,N_3477);
nor U8936 (N_8936,N_4876,N_1264);
or U8937 (N_8937,N_4062,N_1815);
or U8938 (N_8938,N_1855,N_1037);
or U8939 (N_8939,N_3667,N_1953);
nor U8940 (N_8940,N_2632,N_4208);
nand U8941 (N_8941,N_1474,N_3653);
and U8942 (N_8942,N_3456,N_4284);
or U8943 (N_8943,N_2448,N_305);
nand U8944 (N_8944,N_2844,N_4269);
or U8945 (N_8945,N_3597,N_3713);
nand U8946 (N_8946,N_3735,N_3112);
and U8947 (N_8947,N_2560,N_4580);
nor U8948 (N_8948,N_1808,N_3945);
or U8949 (N_8949,N_153,N_4478);
nand U8950 (N_8950,N_416,N_3154);
or U8951 (N_8951,N_2666,N_4125);
nand U8952 (N_8952,N_4441,N_2291);
nor U8953 (N_8953,N_3273,N_1358);
or U8954 (N_8954,N_3886,N_4779);
or U8955 (N_8955,N_2087,N_2905);
nor U8956 (N_8956,N_3962,N_770);
nand U8957 (N_8957,N_3100,N_810);
and U8958 (N_8958,N_3383,N_2510);
nor U8959 (N_8959,N_4910,N_1385);
nor U8960 (N_8960,N_3503,N_3857);
xor U8961 (N_8961,N_3003,N_57);
nor U8962 (N_8962,N_4790,N_1987);
or U8963 (N_8963,N_4743,N_400);
nor U8964 (N_8964,N_871,N_574);
nor U8965 (N_8965,N_1689,N_354);
nor U8966 (N_8966,N_3154,N_702);
nand U8967 (N_8967,N_3952,N_1622);
nor U8968 (N_8968,N_275,N_4223);
nand U8969 (N_8969,N_1893,N_395);
xnor U8970 (N_8970,N_1117,N_1589);
or U8971 (N_8971,N_4532,N_68);
nor U8972 (N_8972,N_4762,N_4008);
nand U8973 (N_8973,N_1621,N_750);
nand U8974 (N_8974,N_3374,N_3806);
nor U8975 (N_8975,N_4390,N_725);
and U8976 (N_8976,N_4981,N_4909);
nand U8977 (N_8977,N_4510,N_3879);
nor U8978 (N_8978,N_359,N_4553);
nor U8979 (N_8979,N_3848,N_609);
nor U8980 (N_8980,N_3339,N_1567);
and U8981 (N_8981,N_2701,N_1561);
nor U8982 (N_8982,N_118,N_3556);
nand U8983 (N_8983,N_2201,N_3675);
or U8984 (N_8984,N_4259,N_872);
and U8985 (N_8985,N_3147,N_525);
and U8986 (N_8986,N_1685,N_2093);
nand U8987 (N_8987,N_3974,N_372);
nor U8988 (N_8988,N_1624,N_4272);
and U8989 (N_8989,N_2862,N_2368);
nor U8990 (N_8990,N_3730,N_1250);
nand U8991 (N_8991,N_921,N_2229);
nand U8992 (N_8992,N_373,N_3524);
or U8993 (N_8993,N_2927,N_879);
and U8994 (N_8994,N_4693,N_3190);
nor U8995 (N_8995,N_2826,N_2841);
and U8996 (N_8996,N_3890,N_3163);
nand U8997 (N_8997,N_1616,N_829);
and U8998 (N_8998,N_2448,N_4248);
nand U8999 (N_8999,N_4429,N_3477);
nand U9000 (N_9000,N_3431,N_1254);
xnor U9001 (N_9001,N_3394,N_2345);
and U9002 (N_9002,N_3453,N_2512);
nand U9003 (N_9003,N_780,N_2855);
or U9004 (N_9004,N_1611,N_709);
or U9005 (N_9005,N_233,N_4648);
nand U9006 (N_9006,N_620,N_302);
nor U9007 (N_9007,N_66,N_2403);
nand U9008 (N_9008,N_4854,N_1099);
or U9009 (N_9009,N_4483,N_224);
xor U9010 (N_9010,N_664,N_1165);
and U9011 (N_9011,N_4985,N_874);
nor U9012 (N_9012,N_3376,N_172);
and U9013 (N_9013,N_395,N_2744);
or U9014 (N_9014,N_984,N_465);
nand U9015 (N_9015,N_735,N_2355);
or U9016 (N_9016,N_3696,N_2242);
xor U9017 (N_9017,N_4794,N_4630);
xnor U9018 (N_9018,N_2858,N_838);
nand U9019 (N_9019,N_4998,N_2722);
and U9020 (N_9020,N_3359,N_1259);
or U9021 (N_9021,N_344,N_3974);
and U9022 (N_9022,N_3981,N_4008);
and U9023 (N_9023,N_168,N_3213);
and U9024 (N_9024,N_4724,N_143);
and U9025 (N_9025,N_4219,N_4218);
nand U9026 (N_9026,N_4947,N_2084);
nor U9027 (N_9027,N_997,N_3052);
or U9028 (N_9028,N_1972,N_206);
nor U9029 (N_9029,N_1725,N_4057);
and U9030 (N_9030,N_2139,N_505);
nand U9031 (N_9031,N_1076,N_3606);
nor U9032 (N_9032,N_934,N_3885);
or U9033 (N_9033,N_4573,N_704);
nor U9034 (N_9034,N_1212,N_3439);
nor U9035 (N_9035,N_795,N_2585);
and U9036 (N_9036,N_4240,N_4146);
and U9037 (N_9037,N_2059,N_4346);
or U9038 (N_9038,N_1856,N_754);
or U9039 (N_9039,N_1693,N_1279);
nor U9040 (N_9040,N_4760,N_2296);
nand U9041 (N_9041,N_4113,N_2439);
and U9042 (N_9042,N_253,N_3598);
xor U9043 (N_9043,N_4364,N_2605);
xnor U9044 (N_9044,N_2040,N_4696);
nand U9045 (N_9045,N_3326,N_61);
or U9046 (N_9046,N_4585,N_2663);
and U9047 (N_9047,N_1223,N_3515);
or U9048 (N_9048,N_4157,N_4578);
nand U9049 (N_9049,N_3599,N_1589);
and U9050 (N_9050,N_3585,N_2815);
nand U9051 (N_9051,N_333,N_4173);
nand U9052 (N_9052,N_4521,N_2569);
or U9053 (N_9053,N_3757,N_1956);
or U9054 (N_9054,N_618,N_2183);
and U9055 (N_9055,N_733,N_777);
nor U9056 (N_9056,N_3798,N_3938);
and U9057 (N_9057,N_4761,N_359);
nand U9058 (N_9058,N_3452,N_4616);
nor U9059 (N_9059,N_2929,N_1324);
or U9060 (N_9060,N_1677,N_328);
and U9061 (N_9061,N_95,N_4102);
and U9062 (N_9062,N_4693,N_3994);
and U9063 (N_9063,N_1691,N_3429);
nand U9064 (N_9064,N_4334,N_286);
and U9065 (N_9065,N_4347,N_2664);
or U9066 (N_9066,N_535,N_2101);
nor U9067 (N_9067,N_2669,N_4680);
nor U9068 (N_9068,N_368,N_3626);
and U9069 (N_9069,N_1504,N_2402);
xnor U9070 (N_9070,N_4336,N_3514);
nor U9071 (N_9071,N_1286,N_4983);
nand U9072 (N_9072,N_688,N_3215);
and U9073 (N_9073,N_2207,N_1560);
or U9074 (N_9074,N_1350,N_3285);
nor U9075 (N_9075,N_4029,N_2813);
and U9076 (N_9076,N_4148,N_2868);
nand U9077 (N_9077,N_2418,N_114);
nor U9078 (N_9078,N_3744,N_751);
nand U9079 (N_9079,N_102,N_1741);
and U9080 (N_9080,N_4600,N_2052);
xnor U9081 (N_9081,N_4266,N_4141);
nor U9082 (N_9082,N_959,N_1109);
and U9083 (N_9083,N_1568,N_1550);
nand U9084 (N_9084,N_4098,N_1147);
xor U9085 (N_9085,N_3193,N_4025);
xor U9086 (N_9086,N_4002,N_5);
nand U9087 (N_9087,N_3939,N_3364);
nand U9088 (N_9088,N_4570,N_3695);
and U9089 (N_9089,N_705,N_269);
and U9090 (N_9090,N_3661,N_3745);
or U9091 (N_9091,N_2892,N_2705);
or U9092 (N_9092,N_520,N_4617);
xnor U9093 (N_9093,N_1063,N_4810);
nand U9094 (N_9094,N_2763,N_4889);
and U9095 (N_9095,N_255,N_4445);
and U9096 (N_9096,N_3056,N_2247);
and U9097 (N_9097,N_3076,N_2408);
or U9098 (N_9098,N_4181,N_1458);
and U9099 (N_9099,N_3307,N_3828);
and U9100 (N_9100,N_2680,N_4335);
nor U9101 (N_9101,N_265,N_994);
and U9102 (N_9102,N_4509,N_668);
and U9103 (N_9103,N_3392,N_3295);
nand U9104 (N_9104,N_3972,N_4599);
nand U9105 (N_9105,N_680,N_1225);
nand U9106 (N_9106,N_2491,N_4237);
nand U9107 (N_9107,N_2616,N_1714);
nand U9108 (N_9108,N_4844,N_325);
nor U9109 (N_9109,N_3784,N_3409);
and U9110 (N_9110,N_4656,N_1043);
nand U9111 (N_9111,N_4735,N_1894);
or U9112 (N_9112,N_2525,N_3019);
nor U9113 (N_9113,N_1307,N_2955);
or U9114 (N_9114,N_1429,N_2001);
nand U9115 (N_9115,N_1600,N_103);
nand U9116 (N_9116,N_3729,N_1363);
or U9117 (N_9117,N_2668,N_1570);
nor U9118 (N_9118,N_4004,N_122);
and U9119 (N_9119,N_3618,N_2363);
nand U9120 (N_9120,N_2296,N_918);
or U9121 (N_9121,N_4862,N_3880);
or U9122 (N_9122,N_4160,N_2726);
nor U9123 (N_9123,N_3554,N_227);
and U9124 (N_9124,N_2242,N_2960);
nor U9125 (N_9125,N_2564,N_4398);
nand U9126 (N_9126,N_2605,N_3111);
or U9127 (N_9127,N_1918,N_1816);
or U9128 (N_9128,N_1649,N_3905);
nand U9129 (N_9129,N_2572,N_4552);
nor U9130 (N_9130,N_3810,N_2165);
or U9131 (N_9131,N_396,N_1056);
and U9132 (N_9132,N_4016,N_3608);
nand U9133 (N_9133,N_599,N_1573);
nand U9134 (N_9134,N_940,N_238);
nand U9135 (N_9135,N_3902,N_694);
and U9136 (N_9136,N_698,N_2542);
nand U9137 (N_9137,N_3222,N_1823);
nor U9138 (N_9138,N_1237,N_1130);
and U9139 (N_9139,N_2191,N_3642);
nor U9140 (N_9140,N_179,N_2839);
nor U9141 (N_9141,N_3857,N_1073);
nor U9142 (N_9142,N_655,N_1348);
or U9143 (N_9143,N_389,N_709);
nor U9144 (N_9144,N_3829,N_3483);
xor U9145 (N_9145,N_4838,N_1975);
and U9146 (N_9146,N_2274,N_4742);
nand U9147 (N_9147,N_1787,N_4737);
and U9148 (N_9148,N_3236,N_274);
nand U9149 (N_9149,N_80,N_2780);
nand U9150 (N_9150,N_1690,N_2869);
nor U9151 (N_9151,N_3162,N_2586);
or U9152 (N_9152,N_1473,N_2082);
or U9153 (N_9153,N_3165,N_1205);
or U9154 (N_9154,N_3714,N_4268);
and U9155 (N_9155,N_1650,N_4304);
nor U9156 (N_9156,N_4089,N_4961);
nor U9157 (N_9157,N_4657,N_1400);
and U9158 (N_9158,N_510,N_3017);
nor U9159 (N_9159,N_1027,N_760);
and U9160 (N_9160,N_791,N_2832);
nor U9161 (N_9161,N_4477,N_2258);
or U9162 (N_9162,N_53,N_1295);
and U9163 (N_9163,N_4510,N_3643);
xnor U9164 (N_9164,N_2742,N_2762);
or U9165 (N_9165,N_1852,N_995);
nor U9166 (N_9166,N_4868,N_3025);
or U9167 (N_9167,N_1360,N_990);
xnor U9168 (N_9168,N_1001,N_3548);
nand U9169 (N_9169,N_4092,N_2341);
and U9170 (N_9170,N_3968,N_1578);
nor U9171 (N_9171,N_2499,N_3219);
or U9172 (N_9172,N_3525,N_2511);
or U9173 (N_9173,N_3680,N_3146);
and U9174 (N_9174,N_1518,N_1558);
or U9175 (N_9175,N_180,N_4046);
and U9176 (N_9176,N_1334,N_1425);
or U9177 (N_9177,N_3850,N_1786);
and U9178 (N_9178,N_3952,N_1030);
xor U9179 (N_9179,N_1778,N_3008);
nand U9180 (N_9180,N_4056,N_594);
nor U9181 (N_9181,N_1565,N_3162);
and U9182 (N_9182,N_2415,N_4807);
and U9183 (N_9183,N_179,N_3986);
nand U9184 (N_9184,N_3418,N_541);
or U9185 (N_9185,N_2125,N_1708);
nor U9186 (N_9186,N_1770,N_2392);
xnor U9187 (N_9187,N_3181,N_1791);
and U9188 (N_9188,N_326,N_1305);
or U9189 (N_9189,N_2255,N_2129);
nor U9190 (N_9190,N_814,N_252);
or U9191 (N_9191,N_3569,N_1924);
nand U9192 (N_9192,N_4489,N_3737);
and U9193 (N_9193,N_1949,N_843);
or U9194 (N_9194,N_1631,N_2634);
nor U9195 (N_9195,N_307,N_417);
or U9196 (N_9196,N_1954,N_1473);
nor U9197 (N_9197,N_1427,N_1240);
nand U9198 (N_9198,N_1646,N_3608);
nand U9199 (N_9199,N_3853,N_159);
nor U9200 (N_9200,N_1690,N_3014);
or U9201 (N_9201,N_1607,N_3420);
and U9202 (N_9202,N_1468,N_2325);
nor U9203 (N_9203,N_1215,N_2278);
and U9204 (N_9204,N_3801,N_4119);
nand U9205 (N_9205,N_86,N_1308);
nand U9206 (N_9206,N_337,N_1047);
nor U9207 (N_9207,N_2500,N_3390);
nand U9208 (N_9208,N_2285,N_3987);
or U9209 (N_9209,N_4212,N_441);
or U9210 (N_9210,N_1368,N_1995);
and U9211 (N_9211,N_3573,N_3710);
nand U9212 (N_9212,N_3037,N_203);
and U9213 (N_9213,N_2218,N_2513);
or U9214 (N_9214,N_1517,N_1157);
and U9215 (N_9215,N_1544,N_4747);
xnor U9216 (N_9216,N_4116,N_4947);
or U9217 (N_9217,N_1456,N_861);
xnor U9218 (N_9218,N_2250,N_2338);
nand U9219 (N_9219,N_2124,N_2412);
nand U9220 (N_9220,N_1677,N_4460);
nand U9221 (N_9221,N_625,N_4447);
or U9222 (N_9222,N_2904,N_595);
or U9223 (N_9223,N_1621,N_1713);
xor U9224 (N_9224,N_4560,N_2063);
or U9225 (N_9225,N_1436,N_4430);
nand U9226 (N_9226,N_1784,N_714);
nand U9227 (N_9227,N_169,N_2159);
nor U9228 (N_9228,N_2062,N_2294);
nand U9229 (N_9229,N_4352,N_4414);
nor U9230 (N_9230,N_4532,N_3962);
nor U9231 (N_9231,N_692,N_3319);
and U9232 (N_9232,N_4656,N_4963);
and U9233 (N_9233,N_2988,N_4386);
nand U9234 (N_9234,N_3767,N_3257);
xor U9235 (N_9235,N_842,N_3636);
xor U9236 (N_9236,N_2693,N_398);
nand U9237 (N_9237,N_962,N_303);
or U9238 (N_9238,N_3873,N_1172);
nor U9239 (N_9239,N_2684,N_204);
nand U9240 (N_9240,N_3564,N_1162);
nor U9241 (N_9241,N_3218,N_3593);
xnor U9242 (N_9242,N_4390,N_2617);
and U9243 (N_9243,N_1333,N_989);
nor U9244 (N_9244,N_2024,N_4390);
nand U9245 (N_9245,N_983,N_3512);
or U9246 (N_9246,N_4045,N_4055);
or U9247 (N_9247,N_3610,N_1560);
nor U9248 (N_9248,N_2459,N_4150);
or U9249 (N_9249,N_2510,N_1088);
nand U9250 (N_9250,N_4764,N_1186);
xor U9251 (N_9251,N_4236,N_486);
and U9252 (N_9252,N_855,N_1241);
nand U9253 (N_9253,N_4398,N_3018);
nor U9254 (N_9254,N_416,N_2496);
and U9255 (N_9255,N_4531,N_1694);
nor U9256 (N_9256,N_2524,N_4736);
or U9257 (N_9257,N_1634,N_4933);
nand U9258 (N_9258,N_1580,N_4483);
nand U9259 (N_9259,N_4960,N_1745);
and U9260 (N_9260,N_1617,N_3160);
nor U9261 (N_9261,N_1183,N_631);
xor U9262 (N_9262,N_3090,N_3972);
nor U9263 (N_9263,N_2076,N_4472);
nand U9264 (N_9264,N_2295,N_4946);
and U9265 (N_9265,N_1779,N_4609);
and U9266 (N_9266,N_4433,N_2151);
nor U9267 (N_9267,N_1840,N_3858);
nand U9268 (N_9268,N_4882,N_166);
xor U9269 (N_9269,N_2550,N_4529);
and U9270 (N_9270,N_2085,N_3797);
nor U9271 (N_9271,N_3571,N_4525);
or U9272 (N_9272,N_1774,N_1916);
xor U9273 (N_9273,N_736,N_2192);
nor U9274 (N_9274,N_3664,N_116);
and U9275 (N_9275,N_4090,N_3303);
or U9276 (N_9276,N_2453,N_1659);
or U9277 (N_9277,N_1532,N_1848);
nand U9278 (N_9278,N_4339,N_2380);
nor U9279 (N_9279,N_2031,N_2817);
xnor U9280 (N_9280,N_4811,N_1472);
xnor U9281 (N_9281,N_2993,N_4322);
nor U9282 (N_9282,N_3975,N_1645);
nor U9283 (N_9283,N_2885,N_1445);
or U9284 (N_9284,N_347,N_2609);
or U9285 (N_9285,N_1608,N_4270);
nor U9286 (N_9286,N_2406,N_2487);
or U9287 (N_9287,N_2017,N_4570);
nand U9288 (N_9288,N_1586,N_1729);
nand U9289 (N_9289,N_4893,N_28);
or U9290 (N_9290,N_3455,N_2051);
nand U9291 (N_9291,N_3036,N_1400);
and U9292 (N_9292,N_642,N_3571);
xnor U9293 (N_9293,N_3437,N_3923);
or U9294 (N_9294,N_2247,N_1001);
nand U9295 (N_9295,N_1721,N_2644);
nor U9296 (N_9296,N_1720,N_4534);
and U9297 (N_9297,N_291,N_690);
or U9298 (N_9298,N_960,N_3934);
nand U9299 (N_9299,N_2577,N_1223);
or U9300 (N_9300,N_3285,N_4176);
xnor U9301 (N_9301,N_502,N_1151);
nor U9302 (N_9302,N_765,N_3544);
nor U9303 (N_9303,N_1020,N_157);
and U9304 (N_9304,N_3908,N_3992);
and U9305 (N_9305,N_3202,N_2791);
nor U9306 (N_9306,N_3602,N_1782);
or U9307 (N_9307,N_4765,N_118);
nor U9308 (N_9308,N_2502,N_4816);
or U9309 (N_9309,N_1134,N_800);
nand U9310 (N_9310,N_4038,N_1150);
and U9311 (N_9311,N_4691,N_2149);
or U9312 (N_9312,N_2746,N_729);
nand U9313 (N_9313,N_2349,N_2736);
nand U9314 (N_9314,N_3602,N_3294);
and U9315 (N_9315,N_4832,N_3143);
and U9316 (N_9316,N_4361,N_100);
xor U9317 (N_9317,N_4732,N_2047);
nand U9318 (N_9318,N_1944,N_113);
nand U9319 (N_9319,N_4590,N_3783);
and U9320 (N_9320,N_4633,N_4445);
or U9321 (N_9321,N_2346,N_4389);
and U9322 (N_9322,N_4928,N_1908);
or U9323 (N_9323,N_1802,N_4613);
and U9324 (N_9324,N_4099,N_174);
or U9325 (N_9325,N_1510,N_1752);
nor U9326 (N_9326,N_78,N_4114);
or U9327 (N_9327,N_2557,N_2998);
or U9328 (N_9328,N_1549,N_1011);
xor U9329 (N_9329,N_2540,N_4128);
xor U9330 (N_9330,N_652,N_1487);
and U9331 (N_9331,N_875,N_2029);
or U9332 (N_9332,N_1160,N_97);
nor U9333 (N_9333,N_133,N_3533);
and U9334 (N_9334,N_1680,N_2034);
and U9335 (N_9335,N_2764,N_2277);
nor U9336 (N_9336,N_3262,N_434);
and U9337 (N_9337,N_4610,N_1843);
or U9338 (N_9338,N_2817,N_4941);
and U9339 (N_9339,N_1450,N_4077);
nor U9340 (N_9340,N_2503,N_1086);
xor U9341 (N_9341,N_1987,N_2495);
and U9342 (N_9342,N_2728,N_4050);
nand U9343 (N_9343,N_2787,N_2600);
nor U9344 (N_9344,N_243,N_1865);
nand U9345 (N_9345,N_711,N_2503);
nor U9346 (N_9346,N_378,N_4789);
and U9347 (N_9347,N_1342,N_2139);
nand U9348 (N_9348,N_1415,N_915);
and U9349 (N_9349,N_1072,N_1930);
nor U9350 (N_9350,N_3269,N_4856);
nand U9351 (N_9351,N_2072,N_4277);
and U9352 (N_9352,N_3882,N_2799);
or U9353 (N_9353,N_48,N_3060);
xor U9354 (N_9354,N_2349,N_3411);
nor U9355 (N_9355,N_1222,N_1114);
or U9356 (N_9356,N_4643,N_2734);
and U9357 (N_9357,N_2241,N_1293);
or U9358 (N_9358,N_1737,N_4009);
and U9359 (N_9359,N_585,N_1477);
xor U9360 (N_9360,N_606,N_2671);
nand U9361 (N_9361,N_4,N_217);
nor U9362 (N_9362,N_2780,N_3207);
nor U9363 (N_9363,N_4369,N_2167);
nor U9364 (N_9364,N_1605,N_4801);
and U9365 (N_9365,N_4232,N_4252);
nand U9366 (N_9366,N_1186,N_2365);
or U9367 (N_9367,N_4760,N_4539);
nor U9368 (N_9368,N_4569,N_727);
nand U9369 (N_9369,N_4932,N_1055);
xor U9370 (N_9370,N_3727,N_4723);
xnor U9371 (N_9371,N_1904,N_1752);
or U9372 (N_9372,N_1504,N_4513);
and U9373 (N_9373,N_1764,N_361);
nand U9374 (N_9374,N_642,N_667);
nand U9375 (N_9375,N_2023,N_1889);
and U9376 (N_9376,N_1731,N_2580);
nor U9377 (N_9377,N_2251,N_2421);
nand U9378 (N_9378,N_3719,N_1521);
nor U9379 (N_9379,N_4092,N_2356);
and U9380 (N_9380,N_1168,N_1216);
and U9381 (N_9381,N_4627,N_4699);
nor U9382 (N_9382,N_189,N_3688);
xnor U9383 (N_9383,N_3013,N_1095);
and U9384 (N_9384,N_392,N_319);
nand U9385 (N_9385,N_3162,N_2856);
or U9386 (N_9386,N_2147,N_3175);
nand U9387 (N_9387,N_1013,N_4789);
nand U9388 (N_9388,N_1505,N_2611);
nand U9389 (N_9389,N_4089,N_2550);
or U9390 (N_9390,N_396,N_2405);
nor U9391 (N_9391,N_1193,N_103);
or U9392 (N_9392,N_621,N_1149);
and U9393 (N_9393,N_2169,N_3763);
and U9394 (N_9394,N_2943,N_3895);
and U9395 (N_9395,N_3749,N_4047);
and U9396 (N_9396,N_549,N_3865);
or U9397 (N_9397,N_4354,N_1547);
xor U9398 (N_9398,N_1840,N_2610);
and U9399 (N_9399,N_4463,N_3509);
nor U9400 (N_9400,N_4104,N_4658);
nand U9401 (N_9401,N_556,N_910);
nand U9402 (N_9402,N_4615,N_4796);
or U9403 (N_9403,N_3989,N_14);
and U9404 (N_9404,N_3671,N_3302);
nand U9405 (N_9405,N_575,N_4409);
nor U9406 (N_9406,N_1360,N_3986);
xor U9407 (N_9407,N_116,N_1544);
and U9408 (N_9408,N_1468,N_2573);
and U9409 (N_9409,N_2352,N_3583);
nand U9410 (N_9410,N_278,N_1928);
nor U9411 (N_9411,N_4568,N_3553);
or U9412 (N_9412,N_2533,N_2767);
nand U9413 (N_9413,N_1527,N_1521);
nor U9414 (N_9414,N_4473,N_2259);
or U9415 (N_9415,N_908,N_3136);
nand U9416 (N_9416,N_1169,N_3665);
nor U9417 (N_9417,N_748,N_4979);
and U9418 (N_9418,N_4003,N_3658);
nor U9419 (N_9419,N_3366,N_3162);
and U9420 (N_9420,N_3045,N_2750);
nand U9421 (N_9421,N_2274,N_2493);
or U9422 (N_9422,N_3831,N_1037);
and U9423 (N_9423,N_542,N_2139);
and U9424 (N_9424,N_1538,N_1992);
nand U9425 (N_9425,N_4429,N_4329);
nor U9426 (N_9426,N_4083,N_2910);
nor U9427 (N_9427,N_1323,N_1139);
and U9428 (N_9428,N_4433,N_2942);
nand U9429 (N_9429,N_3185,N_3389);
nand U9430 (N_9430,N_2819,N_3327);
nor U9431 (N_9431,N_326,N_63);
nand U9432 (N_9432,N_1130,N_2601);
nand U9433 (N_9433,N_3967,N_2924);
xnor U9434 (N_9434,N_1607,N_4067);
or U9435 (N_9435,N_1140,N_3765);
nand U9436 (N_9436,N_2106,N_3175);
or U9437 (N_9437,N_279,N_2080);
or U9438 (N_9438,N_464,N_1995);
nand U9439 (N_9439,N_132,N_4928);
xor U9440 (N_9440,N_4174,N_114);
or U9441 (N_9441,N_2381,N_164);
xnor U9442 (N_9442,N_2349,N_3673);
nor U9443 (N_9443,N_480,N_2144);
and U9444 (N_9444,N_465,N_3283);
nand U9445 (N_9445,N_2997,N_646);
nor U9446 (N_9446,N_459,N_2554);
xor U9447 (N_9447,N_4557,N_3630);
nand U9448 (N_9448,N_121,N_4424);
xnor U9449 (N_9449,N_3317,N_1655);
nand U9450 (N_9450,N_135,N_4344);
nor U9451 (N_9451,N_1424,N_3490);
and U9452 (N_9452,N_3505,N_4350);
and U9453 (N_9453,N_1057,N_1880);
or U9454 (N_9454,N_3430,N_1698);
xor U9455 (N_9455,N_4786,N_4338);
or U9456 (N_9456,N_362,N_3098);
or U9457 (N_9457,N_992,N_2194);
nand U9458 (N_9458,N_3694,N_1379);
nand U9459 (N_9459,N_3536,N_4720);
nor U9460 (N_9460,N_1288,N_4467);
nor U9461 (N_9461,N_3151,N_1519);
nand U9462 (N_9462,N_1420,N_3221);
nor U9463 (N_9463,N_1634,N_2224);
or U9464 (N_9464,N_3607,N_1715);
nor U9465 (N_9465,N_4687,N_2657);
and U9466 (N_9466,N_2103,N_1923);
nand U9467 (N_9467,N_3732,N_3655);
and U9468 (N_9468,N_2274,N_688);
or U9469 (N_9469,N_4534,N_3513);
xor U9470 (N_9470,N_4236,N_1889);
nor U9471 (N_9471,N_657,N_1756);
nor U9472 (N_9472,N_321,N_1601);
and U9473 (N_9473,N_1849,N_4721);
xnor U9474 (N_9474,N_63,N_4035);
nand U9475 (N_9475,N_3346,N_492);
nand U9476 (N_9476,N_3281,N_2064);
nor U9477 (N_9477,N_3617,N_4931);
nor U9478 (N_9478,N_3573,N_2174);
nor U9479 (N_9479,N_2688,N_4548);
and U9480 (N_9480,N_4868,N_1552);
and U9481 (N_9481,N_4733,N_1629);
xnor U9482 (N_9482,N_76,N_1173);
nand U9483 (N_9483,N_2863,N_2921);
nand U9484 (N_9484,N_830,N_2751);
nand U9485 (N_9485,N_1041,N_4244);
or U9486 (N_9486,N_1118,N_2232);
and U9487 (N_9487,N_2813,N_1973);
and U9488 (N_9488,N_597,N_1490);
and U9489 (N_9489,N_2399,N_1155);
nor U9490 (N_9490,N_1554,N_774);
nor U9491 (N_9491,N_1894,N_606);
nand U9492 (N_9492,N_537,N_218);
nand U9493 (N_9493,N_3956,N_2369);
nor U9494 (N_9494,N_4805,N_3631);
or U9495 (N_9495,N_4676,N_2435);
and U9496 (N_9496,N_4809,N_3666);
nand U9497 (N_9497,N_2608,N_584);
and U9498 (N_9498,N_2014,N_4798);
and U9499 (N_9499,N_3797,N_50);
and U9500 (N_9500,N_2132,N_2178);
nor U9501 (N_9501,N_4223,N_3828);
nor U9502 (N_9502,N_4442,N_2611);
nand U9503 (N_9503,N_1569,N_2428);
and U9504 (N_9504,N_1338,N_3155);
nor U9505 (N_9505,N_2215,N_1459);
and U9506 (N_9506,N_444,N_1759);
nor U9507 (N_9507,N_920,N_3998);
or U9508 (N_9508,N_3023,N_1747);
or U9509 (N_9509,N_3731,N_1848);
or U9510 (N_9510,N_1129,N_4366);
nand U9511 (N_9511,N_2987,N_1098);
nor U9512 (N_9512,N_22,N_2913);
nand U9513 (N_9513,N_2341,N_1077);
nor U9514 (N_9514,N_247,N_781);
or U9515 (N_9515,N_2519,N_850);
nor U9516 (N_9516,N_3345,N_4265);
or U9517 (N_9517,N_704,N_1815);
nand U9518 (N_9518,N_333,N_4092);
or U9519 (N_9519,N_4830,N_1325);
xor U9520 (N_9520,N_711,N_643);
nor U9521 (N_9521,N_1219,N_3875);
nor U9522 (N_9522,N_1048,N_1169);
or U9523 (N_9523,N_1198,N_1533);
and U9524 (N_9524,N_2609,N_3615);
and U9525 (N_9525,N_4870,N_4314);
and U9526 (N_9526,N_1482,N_1417);
and U9527 (N_9527,N_1902,N_3870);
nor U9528 (N_9528,N_3081,N_4173);
or U9529 (N_9529,N_3055,N_2080);
and U9530 (N_9530,N_1407,N_701);
xor U9531 (N_9531,N_1371,N_1777);
nor U9532 (N_9532,N_608,N_4687);
nor U9533 (N_9533,N_2257,N_3417);
nand U9534 (N_9534,N_4775,N_3706);
nand U9535 (N_9535,N_634,N_3225);
or U9536 (N_9536,N_217,N_195);
nand U9537 (N_9537,N_4502,N_4849);
and U9538 (N_9538,N_3336,N_2670);
xnor U9539 (N_9539,N_3042,N_1033);
nand U9540 (N_9540,N_4617,N_2167);
and U9541 (N_9541,N_4919,N_1478);
nand U9542 (N_9542,N_943,N_238);
and U9543 (N_9543,N_4254,N_1685);
or U9544 (N_9544,N_1447,N_4942);
and U9545 (N_9545,N_4940,N_2305);
nand U9546 (N_9546,N_4411,N_1557);
or U9547 (N_9547,N_4350,N_3881);
and U9548 (N_9548,N_1554,N_2420);
and U9549 (N_9549,N_1634,N_3705);
nor U9550 (N_9550,N_1401,N_4411);
nor U9551 (N_9551,N_2758,N_3628);
nand U9552 (N_9552,N_1022,N_3987);
nand U9553 (N_9553,N_4838,N_4139);
and U9554 (N_9554,N_1489,N_2922);
xor U9555 (N_9555,N_651,N_4804);
nand U9556 (N_9556,N_978,N_2967);
nand U9557 (N_9557,N_2587,N_1422);
xor U9558 (N_9558,N_1130,N_4400);
and U9559 (N_9559,N_1821,N_3500);
nand U9560 (N_9560,N_3460,N_2236);
nor U9561 (N_9561,N_2010,N_4891);
and U9562 (N_9562,N_1083,N_4334);
nand U9563 (N_9563,N_4885,N_1379);
xor U9564 (N_9564,N_3175,N_4020);
nor U9565 (N_9565,N_4503,N_2835);
and U9566 (N_9566,N_1718,N_4752);
or U9567 (N_9567,N_4209,N_1088);
or U9568 (N_9568,N_2873,N_2465);
and U9569 (N_9569,N_1114,N_66);
or U9570 (N_9570,N_2692,N_499);
and U9571 (N_9571,N_1909,N_2216);
nor U9572 (N_9572,N_3796,N_488);
nor U9573 (N_9573,N_4294,N_1027);
or U9574 (N_9574,N_1451,N_161);
or U9575 (N_9575,N_2633,N_2250);
nand U9576 (N_9576,N_4660,N_2146);
or U9577 (N_9577,N_343,N_2986);
nor U9578 (N_9578,N_4411,N_4873);
nor U9579 (N_9579,N_2548,N_4253);
nand U9580 (N_9580,N_2695,N_3914);
nand U9581 (N_9581,N_4385,N_4310);
nand U9582 (N_9582,N_1019,N_480);
xnor U9583 (N_9583,N_3291,N_2231);
or U9584 (N_9584,N_607,N_3578);
nand U9585 (N_9585,N_556,N_224);
nand U9586 (N_9586,N_4317,N_4135);
or U9587 (N_9587,N_3353,N_4054);
or U9588 (N_9588,N_4604,N_35);
xor U9589 (N_9589,N_182,N_896);
nand U9590 (N_9590,N_3160,N_510);
or U9591 (N_9591,N_3852,N_1735);
and U9592 (N_9592,N_869,N_4755);
xnor U9593 (N_9593,N_269,N_510);
or U9594 (N_9594,N_4162,N_3800);
and U9595 (N_9595,N_4180,N_511);
nor U9596 (N_9596,N_4286,N_284);
and U9597 (N_9597,N_2071,N_4080);
nor U9598 (N_9598,N_4748,N_938);
nand U9599 (N_9599,N_2464,N_2894);
nor U9600 (N_9600,N_2344,N_508);
nor U9601 (N_9601,N_189,N_2685);
nand U9602 (N_9602,N_2610,N_4848);
nor U9603 (N_9603,N_314,N_4588);
nor U9604 (N_9604,N_527,N_3895);
nor U9605 (N_9605,N_3206,N_691);
nand U9606 (N_9606,N_1088,N_4991);
xor U9607 (N_9607,N_4164,N_4371);
and U9608 (N_9608,N_3786,N_4645);
nand U9609 (N_9609,N_4702,N_1976);
or U9610 (N_9610,N_1429,N_311);
nand U9611 (N_9611,N_3558,N_1403);
and U9612 (N_9612,N_1381,N_4591);
nand U9613 (N_9613,N_3083,N_1476);
and U9614 (N_9614,N_2832,N_1662);
and U9615 (N_9615,N_3390,N_4995);
or U9616 (N_9616,N_1613,N_683);
nand U9617 (N_9617,N_717,N_52);
and U9618 (N_9618,N_1187,N_4828);
nor U9619 (N_9619,N_2802,N_395);
nor U9620 (N_9620,N_143,N_4057);
and U9621 (N_9621,N_4055,N_1959);
or U9622 (N_9622,N_4113,N_1301);
or U9623 (N_9623,N_1941,N_3586);
xor U9624 (N_9624,N_3059,N_3561);
nor U9625 (N_9625,N_630,N_4895);
or U9626 (N_9626,N_1107,N_4730);
and U9627 (N_9627,N_3195,N_2154);
or U9628 (N_9628,N_2848,N_1026);
nand U9629 (N_9629,N_4719,N_4980);
or U9630 (N_9630,N_3176,N_1786);
nor U9631 (N_9631,N_1748,N_2549);
nor U9632 (N_9632,N_2816,N_2911);
nor U9633 (N_9633,N_1784,N_1620);
nor U9634 (N_9634,N_96,N_3505);
xor U9635 (N_9635,N_1990,N_2568);
nor U9636 (N_9636,N_2073,N_265);
nor U9637 (N_9637,N_1123,N_2018);
nand U9638 (N_9638,N_1752,N_3642);
or U9639 (N_9639,N_469,N_1477);
nand U9640 (N_9640,N_385,N_2472);
xor U9641 (N_9641,N_36,N_3558);
or U9642 (N_9642,N_1679,N_2356);
nand U9643 (N_9643,N_3329,N_2635);
nand U9644 (N_9644,N_4441,N_4634);
or U9645 (N_9645,N_4830,N_3342);
and U9646 (N_9646,N_1133,N_926);
or U9647 (N_9647,N_1293,N_2385);
nor U9648 (N_9648,N_360,N_833);
and U9649 (N_9649,N_1996,N_838);
nand U9650 (N_9650,N_4724,N_2494);
xnor U9651 (N_9651,N_3372,N_2789);
or U9652 (N_9652,N_2912,N_4020);
nor U9653 (N_9653,N_4966,N_3674);
nor U9654 (N_9654,N_1402,N_983);
and U9655 (N_9655,N_2566,N_740);
nand U9656 (N_9656,N_2751,N_3918);
xor U9657 (N_9657,N_4192,N_2200);
nor U9658 (N_9658,N_2219,N_3142);
nor U9659 (N_9659,N_2558,N_1893);
nand U9660 (N_9660,N_2033,N_2653);
nand U9661 (N_9661,N_3262,N_4498);
and U9662 (N_9662,N_449,N_1794);
nor U9663 (N_9663,N_4354,N_3434);
xor U9664 (N_9664,N_3486,N_4372);
nand U9665 (N_9665,N_1093,N_4300);
xnor U9666 (N_9666,N_3972,N_4570);
nand U9667 (N_9667,N_3144,N_4754);
and U9668 (N_9668,N_3927,N_2029);
nor U9669 (N_9669,N_160,N_1376);
xnor U9670 (N_9670,N_370,N_2567);
or U9671 (N_9671,N_690,N_1295);
and U9672 (N_9672,N_3163,N_2133);
and U9673 (N_9673,N_3025,N_1038);
nand U9674 (N_9674,N_3106,N_1790);
xnor U9675 (N_9675,N_775,N_3343);
nor U9676 (N_9676,N_572,N_1393);
xor U9677 (N_9677,N_3258,N_3154);
and U9678 (N_9678,N_1676,N_1589);
and U9679 (N_9679,N_4713,N_3829);
and U9680 (N_9680,N_4397,N_4615);
nand U9681 (N_9681,N_957,N_933);
and U9682 (N_9682,N_426,N_4894);
and U9683 (N_9683,N_2772,N_322);
or U9684 (N_9684,N_4068,N_1910);
nand U9685 (N_9685,N_3263,N_3502);
or U9686 (N_9686,N_1870,N_2629);
and U9687 (N_9687,N_583,N_2496);
and U9688 (N_9688,N_1474,N_659);
or U9689 (N_9689,N_4635,N_3451);
or U9690 (N_9690,N_4753,N_3635);
nor U9691 (N_9691,N_3949,N_4510);
nand U9692 (N_9692,N_254,N_3555);
xor U9693 (N_9693,N_3112,N_1088);
nor U9694 (N_9694,N_296,N_4751);
nand U9695 (N_9695,N_1907,N_3200);
nor U9696 (N_9696,N_4177,N_1665);
nor U9697 (N_9697,N_1654,N_4275);
or U9698 (N_9698,N_1187,N_1651);
nand U9699 (N_9699,N_4156,N_3923);
and U9700 (N_9700,N_3293,N_1602);
nor U9701 (N_9701,N_4540,N_4611);
nand U9702 (N_9702,N_656,N_1962);
nor U9703 (N_9703,N_2335,N_1231);
nand U9704 (N_9704,N_4367,N_3885);
xnor U9705 (N_9705,N_1227,N_4601);
and U9706 (N_9706,N_4944,N_2866);
nand U9707 (N_9707,N_2298,N_4035);
nand U9708 (N_9708,N_1795,N_209);
nor U9709 (N_9709,N_4958,N_4647);
nor U9710 (N_9710,N_4471,N_2937);
or U9711 (N_9711,N_28,N_1417);
or U9712 (N_9712,N_1800,N_4791);
xnor U9713 (N_9713,N_2169,N_3716);
and U9714 (N_9714,N_1338,N_4574);
or U9715 (N_9715,N_3793,N_3881);
nand U9716 (N_9716,N_1043,N_37);
and U9717 (N_9717,N_4567,N_295);
and U9718 (N_9718,N_3955,N_1940);
or U9719 (N_9719,N_1590,N_3108);
xnor U9720 (N_9720,N_3535,N_1983);
and U9721 (N_9721,N_879,N_1586);
nand U9722 (N_9722,N_2933,N_4755);
nand U9723 (N_9723,N_538,N_987);
and U9724 (N_9724,N_1616,N_1491);
xnor U9725 (N_9725,N_4236,N_1163);
nand U9726 (N_9726,N_3425,N_3342);
or U9727 (N_9727,N_848,N_1662);
or U9728 (N_9728,N_231,N_4454);
and U9729 (N_9729,N_3720,N_608);
nor U9730 (N_9730,N_4052,N_4846);
or U9731 (N_9731,N_3506,N_1583);
or U9732 (N_9732,N_3878,N_1078);
and U9733 (N_9733,N_3401,N_240);
and U9734 (N_9734,N_2580,N_3862);
xnor U9735 (N_9735,N_4940,N_3166);
and U9736 (N_9736,N_1424,N_949);
or U9737 (N_9737,N_814,N_1189);
and U9738 (N_9738,N_4069,N_3012);
or U9739 (N_9739,N_2198,N_4377);
or U9740 (N_9740,N_2676,N_4207);
and U9741 (N_9741,N_516,N_1373);
or U9742 (N_9742,N_936,N_1830);
and U9743 (N_9743,N_4463,N_1094);
nor U9744 (N_9744,N_1854,N_1028);
and U9745 (N_9745,N_4797,N_2073);
nand U9746 (N_9746,N_3381,N_72);
nand U9747 (N_9747,N_2126,N_4213);
nand U9748 (N_9748,N_534,N_4046);
and U9749 (N_9749,N_1827,N_2466);
nor U9750 (N_9750,N_284,N_4216);
nor U9751 (N_9751,N_206,N_20);
or U9752 (N_9752,N_3112,N_4315);
xnor U9753 (N_9753,N_2798,N_2445);
nand U9754 (N_9754,N_3766,N_881);
nor U9755 (N_9755,N_4033,N_1979);
nor U9756 (N_9756,N_785,N_2593);
nand U9757 (N_9757,N_245,N_987);
nor U9758 (N_9758,N_2314,N_781);
and U9759 (N_9759,N_4485,N_2026);
nand U9760 (N_9760,N_2217,N_3111);
nor U9761 (N_9761,N_534,N_1254);
or U9762 (N_9762,N_2886,N_3861);
or U9763 (N_9763,N_1234,N_3967);
nor U9764 (N_9764,N_1442,N_3978);
or U9765 (N_9765,N_2495,N_3727);
and U9766 (N_9766,N_4228,N_1590);
or U9767 (N_9767,N_4029,N_3240);
nor U9768 (N_9768,N_884,N_1106);
xnor U9769 (N_9769,N_4814,N_4789);
nor U9770 (N_9770,N_2410,N_4103);
nor U9771 (N_9771,N_1998,N_1665);
and U9772 (N_9772,N_608,N_3846);
nor U9773 (N_9773,N_2717,N_4843);
and U9774 (N_9774,N_2906,N_3896);
nand U9775 (N_9775,N_258,N_3140);
and U9776 (N_9776,N_1938,N_3551);
and U9777 (N_9777,N_1043,N_2471);
nor U9778 (N_9778,N_604,N_551);
or U9779 (N_9779,N_4,N_3265);
xnor U9780 (N_9780,N_803,N_1786);
or U9781 (N_9781,N_3580,N_2612);
and U9782 (N_9782,N_3970,N_2245);
nand U9783 (N_9783,N_2892,N_326);
nor U9784 (N_9784,N_2826,N_4310);
and U9785 (N_9785,N_4127,N_663);
or U9786 (N_9786,N_1690,N_315);
nand U9787 (N_9787,N_1397,N_544);
xnor U9788 (N_9788,N_1649,N_875);
nor U9789 (N_9789,N_3159,N_4145);
and U9790 (N_9790,N_4792,N_2530);
nand U9791 (N_9791,N_1521,N_2342);
and U9792 (N_9792,N_2394,N_692);
or U9793 (N_9793,N_642,N_4296);
nor U9794 (N_9794,N_3927,N_648);
nor U9795 (N_9795,N_2285,N_3774);
nor U9796 (N_9796,N_243,N_3728);
and U9797 (N_9797,N_2467,N_4991);
or U9798 (N_9798,N_969,N_3723);
and U9799 (N_9799,N_3715,N_4494);
nor U9800 (N_9800,N_3436,N_1428);
nor U9801 (N_9801,N_2431,N_856);
and U9802 (N_9802,N_446,N_2737);
nand U9803 (N_9803,N_2333,N_1010);
or U9804 (N_9804,N_1967,N_3543);
or U9805 (N_9805,N_2265,N_1874);
nand U9806 (N_9806,N_1703,N_3924);
or U9807 (N_9807,N_473,N_1208);
and U9808 (N_9808,N_2325,N_4897);
nor U9809 (N_9809,N_2289,N_1630);
or U9810 (N_9810,N_3928,N_1591);
nor U9811 (N_9811,N_3271,N_3399);
nand U9812 (N_9812,N_3175,N_3918);
and U9813 (N_9813,N_3957,N_2564);
nor U9814 (N_9814,N_3001,N_2772);
xor U9815 (N_9815,N_322,N_3079);
nand U9816 (N_9816,N_2701,N_3174);
xor U9817 (N_9817,N_3136,N_3564);
and U9818 (N_9818,N_1240,N_4041);
or U9819 (N_9819,N_260,N_2196);
nor U9820 (N_9820,N_4543,N_4468);
and U9821 (N_9821,N_3957,N_612);
and U9822 (N_9822,N_2750,N_134);
nor U9823 (N_9823,N_4159,N_3859);
xnor U9824 (N_9824,N_849,N_1994);
or U9825 (N_9825,N_1405,N_319);
and U9826 (N_9826,N_2358,N_3257);
and U9827 (N_9827,N_69,N_810);
or U9828 (N_9828,N_952,N_3712);
and U9829 (N_9829,N_3655,N_1695);
and U9830 (N_9830,N_4292,N_2664);
nor U9831 (N_9831,N_1632,N_4640);
or U9832 (N_9832,N_1469,N_3655);
and U9833 (N_9833,N_2262,N_1198);
nand U9834 (N_9834,N_845,N_4908);
nor U9835 (N_9835,N_346,N_3878);
nand U9836 (N_9836,N_1573,N_2280);
and U9837 (N_9837,N_1798,N_4146);
or U9838 (N_9838,N_3498,N_2423);
or U9839 (N_9839,N_3121,N_4666);
nor U9840 (N_9840,N_4308,N_2221);
nor U9841 (N_9841,N_1827,N_2426);
or U9842 (N_9842,N_1875,N_943);
and U9843 (N_9843,N_4624,N_3375);
nor U9844 (N_9844,N_3892,N_4);
and U9845 (N_9845,N_534,N_2765);
nand U9846 (N_9846,N_3236,N_2369);
nor U9847 (N_9847,N_1627,N_1566);
nand U9848 (N_9848,N_1411,N_4186);
and U9849 (N_9849,N_4228,N_1337);
xnor U9850 (N_9850,N_28,N_3112);
nor U9851 (N_9851,N_3409,N_4929);
or U9852 (N_9852,N_3903,N_949);
and U9853 (N_9853,N_1334,N_3501);
nand U9854 (N_9854,N_218,N_3416);
xnor U9855 (N_9855,N_1915,N_4780);
nand U9856 (N_9856,N_377,N_3556);
or U9857 (N_9857,N_1455,N_4551);
nand U9858 (N_9858,N_2912,N_1534);
or U9859 (N_9859,N_4804,N_4463);
or U9860 (N_9860,N_3111,N_4816);
nand U9861 (N_9861,N_4383,N_3721);
nor U9862 (N_9862,N_1008,N_744);
or U9863 (N_9863,N_1791,N_2435);
and U9864 (N_9864,N_1668,N_4171);
or U9865 (N_9865,N_2157,N_1270);
and U9866 (N_9866,N_4620,N_3085);
xnor U9867 (N_9867,N_4639,N_2609);
nor U9868 (N_9868,N_3791,N_1164);
or U9869 (N_9869,N_1889,N_1671);
or U9870 (N_9870,N_2865,N_398);
nor U9871 (N_9871,N_2982,N_3124);
nor U9872 (N_9872,N_302,N_2912);
and U9873 (N_9873,N_4877,N_2173);
nand U9874 (N_9874,N_2251,N_4999);
xnor U9875 (N_9875,N_1780,N_3759);
or U9876 (N_9876,N_2629,N_2134);
xor U9877 (N_9877,N_3394,N_4781);
or U9878 (N_9878,N_164,N_3241);
nand U9879 (N_9879,N_331,N_2994);
or U9880 (N_9880,N_4011,N_1348);
and U9881 (N_9881,N_936,N_1649);
nor U9882 (N_9882,N_1344,N_1917);
nand U9883 (N_9883,N_2644,N_557);
nor U9884 (N_9884,N_2529,N_4750);
nor U9885 (N_9885,N_2590,N_4880);
or U9886 (N_9886,N_2975,N_1415);
or U9887 (N_9887,N_3283,N_4912);
xor U9888 (N_9888,N_2488,N_2571);
or U9889 (N_9889,N_792,N_274);
xor U9890 (N_9890,N_490,N_4882);
xor U9891 (N_9891,N_2464,N_4577);
and U9892 (N_9892,N_1872,N_4485);
nand U9893 (N_9893,N_4066,N_1246);
or U9894 (N_9894,N_4199,N_3102);
nand U9895 (N_9895,N_3823,N_4000);
nor U9896 (N_9896,N_2564,N_4840);
and U9897 (N_9897,N_2855,N_4927);
nand U9898 (N_9898,N_2771,N_995);
nor U9899 (N_9899,N_2395,N_2600);
or U9900 (N_9900,N_2852,N_567);
and U9901 (N_9901,N_1605,N_900);
nand U9902 (N_9902,N_376,N_1852);
nor U9903 (N_9903,N_3971,N_2478);
nand U9904 (N_9904,N_2094,N_1733);
nand U9905 (N_9905,N_1730,N_443);
nor U9906 (N_9906,N_3304,N_4467);
and U9907 (N_9907,N_91,N_1545);
nand U9908 (N_9908,N_2535,N_1872);
nand U9909 (N_9909,N_4281,N_4);
or U9910 (N_9910,N_1728,N_4984);
or U9911 (N_9911,N_1402,N_1733);
nor U9912 (N_9912,N_1022,N_940);
nor U9913 (N_9913,N_2928,N_2144);
xnor U9914 (N_9914,N_2061,N_86);
and U9915 (N_9915,N_1246,N_4661);
nor U9916 (N_9916,N_4890,N_1924);
nand U9917 (N_9917,N_4487,N_4613);
nor U9918 (N_9918,N_1286,N_3048);
nor U9919 (N_9919,N_4333,N_4755);
nand U9920 (N_9920,N_3983,N_1952);
and U9921 (N_9921,N_1620,N_897);
and U9922 (N_9922,N_4482,N_4088);
and U9923 (N_9923,N_4162,N_2444);
nand U9924 (N_9924,N_1473,N_4661);
xor U9925 (N_9925,N_3037,N_2779);
nor U9926 (N_9926,N_4113,N_4338);
nand U9927 (N_9927,N_2245,N_4821);
nand U9928 (N_9928,N_3891,N_2480);
nand U9929 (N_9929,N_4978,N_2282);
nand U9930 (N_9930,N_4515,N_1133);
nand U9931 (N_9931,N_2755,N_2850);
and U9932 (N_9932,N_1995,N_3780);
and U9933 (N_9933,N_4417,N_895);
nand U9934 (N_9934,N_2954,N_1067);
nand U9935 (N_9935,N_424,N_2864);
and U9936 (N_9936,N_978,N_4693);
nor U9937 (N_9937,N_243,N_516);
and U9938 (N_9938,N_1032,N_2088);
nand U9939 (N_9939,N_829,N_119);
or U9940 (N_9940,N_1933,N_4403);
nor U9941 (N_9941,N_4128,N_3345);
nor U9942 (N_9942,N_1602,N_2385);
or U9943 (N_9943,N_3339,N_229);
nand U9944 (N_9944,N_4546,N_3846);
nand U9945 (N_9945,N_3320,N_2220);
and U9946 (N_9946,N_1628,N_327);
or U9947 (N_9947,N_2361,N_3753);
xnor U9948 (N_9948,N_3732,N_1149);
xor U9949 (N_9949,N_2376,N_1297);
xnor U9950 (N_9950,N_2110,N_771);
xor U9951 (N_9951,N_1062,N_3765);
or U9952 (N_9952,N_4299,N_3027);
nor U9953 (N_9953,N_2809,N_3777);
nor U9954 (N_9954,N_3962,N_4998);
nand U9955 (N_9955,N_4982,N_271);
nand U9956 (N_9956,N_4774,N_4335);
or U9957 (N_9957,N_4323,N_3840);
nor U9958 (N_9958,N_8,N_2026);
nand U9959 (N_9959,N_2156,N_3901);
nand U9960 (N_9960,N_3895,N_2528);
and U9961 (N_9961,N_1855,N_4582);
nor U9962 (N_9962,N_4686,N_2121);
nand U9963 (N_9963,N_2515,N_2216);
xnor U9964 (N_9964,N_4209,N_4094);
nand U9965 (N_9965,N_870,N_3371);
or U9966 (N_9966,N_4899,N_2215);
and U9967 (N_9967,N_813,N_2265);
xor U9968 (N_9968,N_4670,N_2127);
nor U9969 (N_9969,N_3221,N_3604);
nand U9970 (N_9970,N_1110,N_4798);
nor U9971 (N_9971,N_2785,N_4435);
xor U9972 (N_9972,N_1117,N_4291);
or U9973 (N_9973,N_1175,N_3412);
or U9974 (N_9974,N_731,N_291);
nor U9975 (N_9975,N_4202,N_2663);
or U9976 (N_9976,N_3485,N_4161);
xnor U9977 (N_9977,N_3999,N_1650);
nand U9978 (N_9978,N_846,N_2645);
and U9979 (N_9979,N_4130,N_2935);
xnor U9980 (N_9980,N_3387,N_3103);
nor U9981 (N_9981,N_1481,N_1280);
nand U9982 (N_9982,N_4866,N_4063);
nor U9983 (N_9983,N_4194,N_4923);
nand U9984 (N_9984,N_542,N_926);
nor U9985 (N_9985,N_3621,N_686);
or U9986 (N_9986,N_1923,N_471);
or U9987 (N_9987,N_1340,N_1512);
or U9988 (N_9988,N_3144,N_1900);
nor U9989 (N_9989,N_4312,N_3972);
or U9990 (N_9990,N_1810,N_947);
nor U9991 (N_9991,N_3161,N_677);
xor U9992 (N_9992,N_4480,N_1970);
and U9993 (N_9993,N_1064,N_4011);
or U9994 (N_9994,N_4125,N_1552);
nor U9995 (N_9995,N_1957,N_4358);
nor U9996 (N_9996,N_2006,N_1494);
xnor U9997 (N_9997,N_4461,N_1998);
nor U9998 (N_9998,N_2531,N_2946);
or U9999 (N_9999,N_1280,N_118);
or UO_0 (O_0,N_7986,N_6305);
and UO_1 (O_1,N_9365,N_5937);
and UO_2 (O_2,N_9996,N_7646);
xnor UO_3 (O_3,N_9403,N_5165);
nand UO_4 (O_4,N_8936,N_7155);
and UO_5 (O_5,N_5432,N_8783);
nor UO_6 (O_6,N_6433,N_8730);
or UO_7 (O_7,N_5314,N_9304);
or UO_8 (O_8,N_8025,N_5045);
and UO_9 (O_9,N_6044,N_5544);
xor UO_10 (O_10,N_9378,N_8404);
or UO_11 (O_11,N_6866,N_8100);
nand UO_12 (O_12,N_6244,N_5187);
nor UO_13 (O_13,N_5125,N_7915);
nand UO_14 (O_14,N_7477,N_5679);
nand UO_15 (O_15,N_8830,N_6040);
or UO_16 (O_16,N_7310,N_5050);
and UO_17 (O_17,N_6386,N_7689);
and UO_18 (O_18,N_8427,N_9381);
and UO_19 (O_19,N_8727,N_9442);
and UO_20 (O_20,N_9083,N_6637);
nor UO_21 (O_21,N_8715,N_6589);
nor UO_22 (O_22,N_5483,N_9071);
or UO_23 (O_23,N_8801,N_5920);
nor UO_24 (O_24,N_5979,N_9404);
xor UO_25 (O_25,N_5473,N_7885);
or UO_26 (O_26,N_8135,N_7097);
and UO_27 (O_27,N_6994,N_6742);
nand UO_28 (O_28,N_8854,N_6666);
or UO_29 (O_29,N_7391,N_6004);
nand UO_30 (O_30,N_9266,N_7588);
nand UO_31 (O_31,N_9073,N_8264);
xor UO_32 (O_32,N_5459,N_9253);
nor UO_33 (O_33,N_6932,N_7392);
nor UO_34 (O_34,N_5016,N_9048);
or UO_35 (O_35,N_9641,N_9542);
nand UO_36 (O_36,N_6240,N_8067);
and UO_37 (O_37,N_8263,N_9337);
or UO_38 (O_38,N_7458,N_8348);
and UO_39 (O_39,N_8608,N_7878);
nand UO_40 (O_40,N_8588,N_5002);
or UO_41 (O_41,N_5650,N_7846);
nand UO_42 (O_42,N_5768,N_8669);
and UO_43 (O_43,N_6032,N_7060);
xnor UO_44 (O_44,N_7868,N_6169);
or UO_45 (O_45,N_6989,N_8329);
nor UO_46 (O_46,N_7172,N_9636);
and UO_47 (O_47,N_7183,N_6233);
nand UO_48 (O_48,N_7195,N_7002);
nor UO_49 (O_49,N_8636,N_9499);
or UO_50 (O_50,N_6339,N_9098);
xor UO_51 (O_51,N_8618,N_5211);
nor UO_52 (O_52,N_8514,N_8421);
and UO_53 (O_53,N_5085,N_7051);
or UO_54 (O_54,N_9296,N_8554);
and UO_55 (O_55,N_6996,N_9050);
or UO_56 (O_56,N_8297,N_5651);
and UO_57 (O_57,N_8026,N_6813);
nand UO_58 (O_58,N_9383,N_8892);
nand UO_59 (O_59,N_5500,N_6460);
or UO_60 (O_60,N_6404,N_9410);
and UO_61 (O_61,N_7541,N_7189);
xnor UO_62 (O_62,N_5763,N_6740);
or UO_63 (O_63,N_7231,N_7190);
nand UO_64 (O_64,N_8580,N_6997);
nor UO_65 (O_65,N_6374,N_8822);
nor UO_66 (O_66,N_6066,N_9801);
or UO_67 (O_67,N_7960,N_7680);
or UO_68 (O_68,N_8697,N_7018);
and UO_69 (O_69,N_7431,N_6471);
nor UO_70 (O_70,N_8908,N_8887);
nor UO_71 (O_71,N_7781,N_6319);
or UO_72 (O_72,N_6346,N_6415);
nand UO_73 (O_73,N_9836,N_5606);
or UO_74 (O_74,N_5388,N_5964);
and UO_75 (O_75,N_6204,N_5633);
and UO_76 (O_76,N_7252,N_6185);
nand UO_77 (O_77,N_8826,N_9165);
xnor UO_78 (O_78,N_9190,N_5647);
and UO_79 (O_79,N_7197,N_8397);
nor UO_80 (O_80,N_7522,N_6601);
nor UO_81 (O_81,N_5117,N_6219);
and UO_82 (O_82,N_5454,N_8034);
nand UO_83 (O_83,N_7809,N_7749);
and UO_84 (O_84,N_8315,N_6886);
or UO_85 (O_85,N_7660,N_5526);
and UO_86 (O_86,N_8598,N_9605);
and UO_87 (O_87,N_6906,N_5069);
or UO_88 (O_88,N_7016,N_9762);
nand UO_89 (O_89,N_8012,N_7077);
and UO_90 (O_90,N_6789,N_5822);
nor UO_91 (O_91,N_9407,N_9336);
or UO_92 (O_92,N_9901,N_7293);
xor UO_93 (O_93,N_6384,N_6035);
nand UO_94 (O_94,N_5401,N_5693);
nor UO_95 (O_95,N_7121,N_9565);
or UO_96 (O_96,N_8585,N_9388);
or UO_97 (O_97,N_5206,N_8484);
nor UO_98 (O_98,N_6889,N_7799);
or UO_99 (O_99,N_8316,N_5209);
nor UO_100 (O_100,N_9002,N_8412);
nand UO_101 (O_101,N_8453,N_5222);
nand UO_102 (O_102,N_5752,N_7151);
nor UO_103 (O_103,N_8152,N_5872);
nand UO_104 (O_104,N_8725,N_7210);
nand UO_105 (O_105,N_7906,N_8317);
or UO_106 (O_106,N_8396,N_5531);
and UO_107 (O_107,N_5374,N_7728);
xor UO_108 (O_108,N_5097,N_7313);
nand UO_109 (O_109,N_7670,N_5952);
nand UO_110 (O_110,N_5639,N_8774);
or UO_111 (O_111,N_5244,N_5151);
and UO_112 (O_112,N_8246,N_7178);
nor UO_113 (O_113,N_5636,N_6992);
nand UO_114 (O_114,N_5710,N_6036);
or UO_115 (O_115,N_8247,N_8270);
or UO_116 (O_116,N_5021,N_6598);
nor UO_117 (O_117,N_7020,N_6486);
nor UO_118 (O_118,N_6730,N_7732);
nand UO_119 (O_119,N_7665,N_9062);
nor UO_120 (O_120,N_5834,N_9069);
or UO_121 (O_121,N_9529,N_7596);
and UO_122 (O_122,N_5999,N_6777);
nor UO_123 (O_123,N_9342,N_5279);
nor UO_124 (O_124,N_8455,N_8546);
nor UO_125 (O_125,N_8757,N_7985);
or UO_126 (O_126,N_9966,N_6818);
and UO_127 (O_127,N_9248,N_6496);
nand UO_128 (O_128,N_6321,N_5458);
nor UO_129 (O_129,N_8158,N_5741);
and UO_130 (O_130,N_8547,N_7860);
xor UO_131 (O_131,N_8930,N_6549);
or UO_132 (O_132,N_8712,N_7390);
and UO_133 (O_133,N_5832,N_7717);
and UO_134 (O_134,N_6135,N_9586);
xor UO_135 (O_135,N_5162,N_9869);
nand UO_136 (O_136,N_8889,N_6313);
or UO_137 (O_137,N_9979,N_5047);
and UO_138 (O_138,N_8651,N_9101);
xor UO_139 (O_139,N_9640,N_6493);
or UO_140 (O_140,N_7794,N_7113);
or UO_141 (O_141,N_7352,N_5734);
xor UO_142 (O_142,N_7281,N_9281);
nor UO_143 (O_143,N_8119,N_6689);
nor UO_144 (O_144,N_6951,N_6188);
nand UO_145 (O_145,N_8298,N_5419);
and UO_146 (O_146,N_6656,N_8419);
and UO_147 (O_147,N_9761,N_6525);
or UO_148 (O_148,N_8732,N_9091);
nand UO_149 (O_149,N_8311,N_9340);
nor UO_150 (O_150,N_6638,N_7479);
xor UO_151 (O_151,N_9862,N_6034);
nor UO_152 (O_152,N_7412,N_8952);
nor UO_153 (O_153,N_8880,N_8234);
nor UO_154 (O_154,N_5386,N_8261);
and UO_155 (O_155,N_8232,N_8074);
nor UO_156 (O_156,N_9507,N_6796);
nor UO_157 (O_157,N_9416,N_5276);
xor UO_158 (O_158,N_9938,N_5564);
nor UO_159 (O_159,N_8466,N_9881);
nor UO_160 (O_160,N_5384,N_5858);
and UO_161 (O_161,N_8147,N_7659);
nor UO_162 (O_162,N_6076,N_6322);
and UO_163 (O_163,N_9376,N_6002);
or UO_164 (O_164,N_9627,N_8858);
nor UO_165 (O_165,N_6892,N_5332);
or UO_166 (O_166,N_7220,N_6574);
nor UO_167 (O_167,N_5750,N_8888);
nor UO_168 (O_168,N_9210,N_8020);
nand UO_169 (O_169,N_5929,N_9319);
and UO_170 (O_170,N_8549,N_7305);
nor UO_171 (O_171,N_9164,N_6332);
nor UO_172 (O_172,N_5168,N_6086);
xor UO_173 (O_173,N_9750,N_7090);
or UO_174 (O_174,N_7086,N_6077);
nor UO_175 (O_175,N_9488,N_8379);
or UO_176 (O_176,N_5193,N_8513);
nor UO_177 (O_177,N_8813,N_8036);
and UO_178 (O_178,N_8028,N_6868);
nand UO_179 (O_179,N_7615,N_6464);
nor UO_180 (O_180,N_8800,N_7202);
or UO_181 (O_181,N_8022,N_8371);
nor UO_182 (O_182,N_5787,N_8390);
or UO_183 (O_183,N_7297,N_7987);
and UO_184 (O_184,N_5030,N_8569);
or UO_185 (O_185,N_9568,N_7285);
nor UO_186 (O_186,N_7716,N_5014);
or UO_187 (O_187,N_7843,N_8215);
and UO_188 (O_188,N_8082,N_5119);
nor UO_189 (O_189,N_6912,N_9398);
nand UO_190 (O_190,N_6023,N_6883);
xor UO_191 (O_191,N_6990,N_9053);
nand UO_192 (O_192,N_5199,N_9543);
xor UO_193 (O_193,N_8201,N_6973);
or UO_194 (O_194,N_5003,N_7028);
and UO_195 (O_195,N_7707,N_8155);
nand UO_196 (O_196,N_6820,N_6256);
or UO_197 (O_197,N_5502,N_7094);
xnor UO_198 (O_198,N_8079,N_9918);
and UO_199 (O_199,N_5041,N_8179);
nor UO_200 (O_200,N_6393,N_6545);
nor UO_201 (O_201,N_8570,N_8874);
and UO_202 (O_202,N_8997,N_9854);
or UO_203 (O_203,N_5177,N_9931);
or UO_204 (O_204,N_5334,N_9267);
or UO_205 (O_205,N_8407,N_9865);
nor UO_206 (O_206,N_5038,N_9070);
nor UO_207 (O_207,N_7582,N_5448);
or UO_208 (O_208,N_7444,N_7655);
nor UO_209 (O_209,N_5356,N_9800);
xor UO_210 (O_210,N_5729,N_8057);
and UO_211 (O_211,N_7388,N_5004);
nor UO_212 (O_212,N_5113,N_7849);
xnor UO_213 (O_213,N_8502,N_7695);
nor UO_214 (O_214,N_8907,N_7875);
and UO_215 (O_215,N_8184,N_8252);
or UO_216 (O_216,N_9832,N_9922);
nor UO_217 (O_217,N_5203,N_7696);
xor UO_218 (O_218,N_5815,N_6170);
and UO_219 (O_219,N_8567,N_7153);
nand UO_220 (O_220,N_6413,N_8749);
nand UO_221 (O_221,N_7578,N_9623);
nand UO_222 (O_222,N_8664,N_8214);
nor UO_223 (O_223,N_5155,N_6306);
nand UO_224 (O_224,N_9937,N_9430);
and UO_225 (O_225,N_6378,N_7750);
nor UO_226 (O_226,N_6297,N_8449);
xnor UO_227 (O_227,N_5928,N_8832);
nor UO_228 (O_228,N_8070,N_7529);
and UO_229 (O_229,N_8678,N_8702);
nand UO_230 (O_230,N_5511,N_5265);
or UO_231 (O_231,N_8497,N_7258);
nor UO_232 (O_232,N_9424,N_6084);
nand UO_233 (O_233,N_5492,N_7658);
and UO_234 (O_234,N_8743,N_5471);
or UO_235 (O_235,N_9178,N_5347);
and UO_236 (O_236,N_9495,N_8210);
nor UO_237 (O_237,N_6565,N_9331);
and UO_238 (O_238,N_5583,N_9930);
xor UO_239 (O_239,N_5798,N_9024);
nand UO_240 (O_240,N_9450,N_9453);
nor UO_241 (O_241,N_9326,N_6283);
nor UO_242 (O_242,N_9116,N_5799);
xnor UO_243 (O_243,N_5404,N_6962);
and UO_244 (O_244,N_8521,N_7493);
and UO_245 (O_245,N_5731,N_5441);
and UO_246 (O_246,N_7834,N_6163);
or UO_247 (O_247,N_6555,N_8380);
nor UO_248 (O_248,N_9890,N_9545);
or UO_249 (O_249,N_8465,N_6375);
or UO_250 (O_250,N_9081,N_5727);
nand UO_251 (O_251,N_8719,N_6705);
nor UO_252 (O_252,N_9555,N_5785);
or UO_253 (O_253,N_7650,N_6161);
nor UO_254 (O_254,N_5446,N_5540);
and UO_255 (O_255,N_5931,N_5890);
nor UO_256 (O_256,N_8094,N_7015);
nor UO_257 (O_257,N_9230,N_7786);
nand UO_258 (O_258,N_7602,N_6538);
or UO_259 (O_259,N_9969,N_5274);
nor UO_260 (O_260,N_9561,N_5644);
or UO_261 (O_261,N_8487,N_9910);
or UO_262 (O_262,N_7771,N_7159);
or UO_263 (O_263,N_9115,N_9504);
or UO_264 (O_264,N_6902,N_8562);
nor UO_265 (O_265,N_5617,N_6618);
and UO_266 (O_266,N_5558,N_6098);
xor UO_267 (O_267,N_7026,N_5289);
nand UO_268 (O_268,N_8668,N_7349);
nor UO_269 (O_269,N_7919,N_8835);
nand UO_270 (O_270,N_6327,N_6682);
and UO_271 (O_271,N_8577,N_9447);
nor UO_272 (O_272,N_5367,N_5150);
nand UO_273 (O_273,N_5873,N_7278);
or UO_274 (O_274,N_6695,N_9272);
and UO_275 (O_275,N_5747,N_6765);
xor UO_276 (O_276,N_6114,N_6647);
nand UO_277 (O_277,N_7734,N_5144);
or UO_278 (O_278,N_6142,N_8040);
xor UO_279 (O_279,N_7382,N_6046);
and UO_280 (O_280,N_5417,N_9089);
nor UO_281 (O_281,N_8980,N_7515);
and UO_282 (O_282,N_9205,N_9698);
nor UO_283 (O_283,N_5059,N_5934);
nor UO_284 (O_284,N_5760,N_8342);
or UO_285 (O_285,N_7299,N_9859);
and UO_286 (O_286,N_8222,N_9736);
nor UO_287 (O_287,N_5058,N_9485);
nand UO_288 (O_288,N_9126,N_9658);
or UO_289 (O_289,N_6759,N_5582);
and UO_290 (O_290,N_7499,N_7263);
nor UO_291 (O_291,N_5912,N_6512);
and UO_292 (O_292,N_8820,N_6232);
or UO_293 (O_293,N_8017,N_9515);
nor UO_294 (O_294,N_5008,N_9574);
or UO_295 (O_295,N_5083,N_7400);
nand UO_296 (O_296,N_7242,N_9770);
nand UO_297 (O_297,N_7992,N_9707);
nand UO_298 (O_298,N_6749,N_8123);
or UO_299 (O_299,N_5810,N_8806);
nor UO_300 (O_300,N_7721,N_8842);
nand UO_301 (O_301,N_7244,N_5295);
nor UO_302 (O_302,N_8501,N_5285);
nor UO_303 (O_303,N_9136,N_6942);
nand UO_304 (O_304,N_9571,N_5423);
nand UO_305 (O_305,N_8912,N_9973);
or UO_306 (O_306,N_9321,N_6455);
and UO_307 (O_307,N_7685,N_6873);
nor UO_308 (O_308,N_8797,N_9722);
nand UO_309 (O_309,N_9883,N_5443);
nor UO_310 (O_310,N_8282,N_9455);
and UO_311 (O_311,N_7550,N_5549);
and UO_312 (O_312,N_5195,N_5975);
or UO_313 (O_313,N_9651,N_7756);
or UO_314 (O_314,N_5043,N_5344);
nand UO_315 (O_315,N_5288,N_8682);
nand UO_316 (O_316,N_9778,N_6788);
or UO_317 (O_317,N_6885,N_7718);
or UO_318 (O_318,N_8808,N_7152);
xor UO_319 (O_319,N_9022,N_5974);
and UO_320 (O_320,N_6414,N_5072);
or UO_321 (O_321,N_6307,N_7760);
nand UO_322 (O_322,N_7674,N_5357);
nor UO_323 (O_323,N_8624,N_8524);
or UO_324 (O_324,N_7594,N_7702);
nor UO_325 (O_325,N_5322,N_7759);
or UO_326 (O_326,N_7741,N_5158);
or UO_327 (O_327,N_9462,N_9280);
nand UO_328 (O_328,N_9783,N_5425);
and UO_329 (O_329,N_6898,N_8983);
and UO_330 (O_330,N_7139,N_8452);
nor UO_331 (O_331,N_5353,N_7304);
xor UO_332 (O_332,N_5317,N_8294);
and UO_333 (O_333,N_8853,N_7389);
xnor UO_334 (O_334,N_8340,N_8929);
nor UO_335 (O_335,N_8714,N_6717);
or UO_336 (O_336,N_5198,N_7548);
nand UO_337 (O_337,N_5954,N_7478);
and UO_338 (O_338,N_5715,N_9146);
nand UO_339 (O_339,N_5089,N_7560);
nor UO_340 (O_340,N_9697,N_8869);
nor UO_341 (O_341,N_9773,N_5240);
nor UO_342 (O_342,N_6469,N_7935);
or UO_343 (O_343,N_7954,N_5694);
or UO_344 (O_344,N_9170,N_8504);
nand UO_345 (O_345,N_8072,N_6888);
and UO_346 (O_346,N_7928,N_6217);
and UO_347 (O_347,N_5498,N_8747);
nor UO_348 (O_348,N_8233,N_7296);
xnor UO_349 (O_349,N_8503,N_6477);
or UO_350 (O_350,N_7514,N_5088);
and UO_351 (O_351,N_9127,N_9289);
nor UO_352 (O_352,N_7095,N_7232);
nor UO_353 (O_353,N_8928,N_9234);
nand UO_354 (O_354,N_8753,N_9182);
nand UO_355 (O_355,N_5499,N_7953);
xor UO_356 (O_356,N_6335,N_9372);
and UO_357 (O_357,N_7469,N_8167);
nand UO_358 (O_358,N_7733,N_7071);
nand UO_359 (O_359,N_8129,N_9619);
and UO_360 (O_360,N_7017,N_5786);
or UO_361 (O_361,N_8610,N_7651);
nor UO_362 (O_362,N_9841,N_6422);
or UO_363 (O_363,N_7859,N_8467);
nor UO_364 (O_364,N_8648,N_6881);
xor UO_365 (O_365,N_6727,N_5812);
xor UO_366 (O_366,N_5933,N_8175);
or UO_367 (O_367,N_6222,N_5173);
nand UO_368 (O_368,N_9806,N_7948);
nor UO_369 (O_369,N_5464,N_5174);
and UO_370 (O_370,N_5349,N_8394);
and UO_371 (O_371,N_5067,N_6442);
nor UO_372 (O_372,N_6728,N_5576);
nand UO_373 (O_373,N_8245,N_6459);
xnor UO_374 (O_374,N_8941,N_5093);
nor UO_375 (O_375,N_6710,N_8037);
xor UO_376 (O_376,N_6277,N_8647);
nor UO_377 (O_377,N_6751,N_6879);
and UO_378 (O_378,N_6083,N_5476);
nand UO_379 (O_379,N_9104,N_6838);
and UO_380 (O_380,N_5581,N_9294);
nand UO_381 (O_381,N_6528,N_8643);
or UO_382 (O_382,N_9500,N_6167);
or UO_383 (O_383,N_5250,N_7630);
nand UO_384 (O_384,N_9834,N_6221);
nor UO_385 (O_385,N_5854,N_5159);
or UO_386 (O_386,N_6753,N_7981);
nand UO_387 (O_387,N_9068,N_8211);
nor UO_388 (O_388,N_7826,N_6571);
or UO_389 (O_389,N_8529,N_8511);
nand UO_390 (O_390,N_5126,N_8226);
nor UO_391 (O_391,N_9276,N_5666);
nand UO_392 (O_392,N_8720,N_5343);
nand UO_393 (O_393,N_5541,N_6085);
and UO_394 (O_394,N_7486,N_9514);
nor UO_395 (O_395,N_7998,N_5108);
nor UO_396 (O_396,N_9799,N_6063);
xnor UO_397 (O_397,N_9647,N_6617);
xnor UO_398 (O_398,N_9271,N_8860);
and UO_399 (O_399,N_7820,N_6918);
or UO_400 (O_400,N_7979,N_5457);
nor UO_401 (O_401,N_9815,N_7553);
and UO_402 (O_402,N_8065,N_8674);
and UO_403 (O_403,N_7368,N_5762);
or UO_404 (O_404,N_5853,N_7064);
nand UO_405 (O_405,N_7123,N_8370);
nor UO_406 (O_406,N_9360,N_7637);
and UO_407 (O_407,N_9604,N_6195);
nand UO_408 (O_408,N_6588,N_6071);
and UO_409 (O_409,N_7672,N_9419);
nor UO_410 (O_410,N_6465,N_5363);
nor UO_411 (O_411,N_8053,N_5348);
and UO_412 (O_412,N_8954,N_9496);
nand UO_413 (O_413,N_8837,N_6882);
and UO_414 (O_414,N_8185,N_7185);
and UO_415 (O_415,N_5309,N_9217);
nor UO_416 (O_416,N_8127,N_7157);
and UO_417 (O_417,N_8220,N_9874);
nand UO_418 (O_418,N_9380,N_8159);
nor UO_419 (O_419,N_7221,N_6547);
or UO_420 (O_420,N_5765,N_8003);
xnor UO_421 (O_421,N_7742,N_5609);
nor UO_422 (O_422,N_9540,N_6871);
or UO_423 (O_423,N_7745,N_9395);
nor UO_424 (O_424,N_9110,N_8124);
nand UO_425 (O_425,N_8238,N_5927);
nand UO_426 (O_426,N_6336,N_9386);
or UO_427 (O_427,N_6488,N_7324);
nor UO_428 (O_428,N_8828,N_8676);
nor UO_429 (O_429,N_5652,N_8959);
nand UO_430 (O_430,N_9858,N_7024);
or UO_431 (O_431,N_7533,N_7226);
nor UO_432 (O_432,N_8638,N_7699);
nor UO_433 (O_433,N_9904,N_6097);
nand UO_434 (O_434,N_5976,N_8196);
nor UO_435 (O_435,N_7812,N_5273);
nor UO_436 (O_436,N_7481,N_9700);
nand UO_437 (O_437,N_6479,N_5063);
and UO_438 (O_438,N_7598,N_9669);
nor UO_439 (O_439,N_7704,N_7413);
nor UO_440 (O_440,N_7092,N_5632);
nand UO_441 (O_441,N_8641,N_8321);
or UO_442 (O_442,N_8385,N_7513);
or UO_443 (O_443,N_7975,N_7498);
and UO_444 (O_444,N_9125,N_5567);
nand UO_445 (O_445,N_8976,N_5191);
nor UO_446 (O_446,N_7965,N_9580);
or UO_447 (O_447,N_8451,N_9733);
nor UO_448 (O_448,N_6109,N_5392);
nand UO_449 (O_449,N_8434,N_9274);
nand UO_450 (O_450,N_9092,N_7080);
or UO_451 (O_451,N_6419,N_5137);
nor UO_452 (O_452,N_5692,N_7467);
nor UO_453 (O_453,N_7914,N_8746);
or UO_454 (O_454,N_6977,N_8906);
nor UO_455 (O_455,N_5139,N_7193);
or UO_456 (O_456,N_7423,N_7879);
or UO_457 (O_457,N_5660,N_9458);
and UO_458 (O_458,N_9737,N_5641);
and UO_459 (O_459,N_5739,N_8219);
and UO_460 (O_460,N_8389,N_9279);
nand UO_461 (O_461,N_7564,N_7687);
and UO_462 (O_462,N_8721,N_5231);
and UO_463 (O_463,N_7977,N_5111);
xor UO_464 (O_464,N_7817,N_8982);
and UO_465 (O_465,N_5210,N_6639);
nand UO_466 (O_466,N_7302,N_7823);
and UO_467 (O_467,N_5084,N_9614);
and UO_468 (O_468,N_5300,N_5204);
nor UO_469 (O_469,N_6584,N_5114);
and UO_470 (O_470,N_5548,N_8814);
or UO_471 (O_471,N_9269,N_8769);
nor UO_472 (O_472,N_6110,N_5128);
or UO_473 (O_473,N_6683,N_6176);
or UO_474 (O_474,N_6829,N_6856);
or UO_475 (O_475,N_7136,N_8841);
and UO_476 (O_476,N_8055,N_9818);
nand UO_477 (O_477,N_9731,N_9719);
nand UO_478 (O_478,N_8574,N_8292);
or UO_479 (O_479,N_8059,N_6225);
nor UO_480 (O_480,N_8778,N_6612);
or UO_481 (O_481,N_7639,N_6424);
nor UO_482 (O_482,N_6651,N_6965);
and UO_483 (O_483,N_8780,N_9909);
nand UO_484 (O_484,N_8823,N_6983);
xor UO_485 (O_485,N_7886,N_8363);
and UO_486 (O_486,N_9777,N_6139);
nand UO_487 (O_487,N_7326,N_7107);
nand UO_488 (O_488,N_9273,N_5426);
xor UO_489 (O_489,N_7798,N_9556);
and UO_490 (O_490,N_9406,N_5537);
and UO_491 (O_491,N_8527,N_5788);
nor UO_492 (O_492,N_9879,N_8459);
and UO_493 (O_493,N_9309,N_7072);
nor UO_494 (O_494,N_7645,N_7169);
and UO_495 (O_495,N_9724,N_9796);
nand UO_496 (O_496,N_7887,N_6731);
and UO_497 (O_497,N_8326,N_5217);
and UO_498 (O_498,N_5337,N_5095);
or UO_499 (O_499,N_5081,N_5801);
nor UO_500 (O_500,N_6858,N_7029);
or UO_501 (O_501,N_8408,N_9389);
nor UO_502 (O_502,N_7254,N_5603);
and UO_503 (O_503,N_7269,N_6416);
or UO_504 (O_504,N_8286,N_7929);
nand UO_505 (O_505,N_8093,N_7891);
nand UO_506 (O_506,N_7996,N_7726);
nand UO_507 (O_507,N_9790,N_8685);
xor UO_508 (O_508,N_6338,N_7656);
nand UO_509 (O_509,N_5398,N_7785);
xor UO_510 (O_510,N_6516,N_6672);
or UO_511 (O_511,N_9672,N_8216);
nand UO_512 (O_512,N_5070,N_6485);
nand UO_513 (O_513,N_6209,N_6235);
and UO_514 (O_514,N_9211,N_5884);
nand UO_515 (O_515,N_9420,N_7484);
nor UO_516 (O_516,N_5839,N_9343);
or UO_517 (O_517,N_8493,N_8890);
and UO_518 (O_518,N_6830,N_8223);
xor UO_519 (O_519,N_7112,N_5698);
and UO_520 (O_520,N_9167,N_7943);
or UO_521 (O_521,N_7889,N_9921);
or UO_522 (O_522,N_7995,N_8273);
or UO_523 (O_523,N_6273,N_5055);
nand UO_524 (O_524,N_8162,N_7663);
or UO_525 (O_525,N_7215,N_6101);
nor UO_526 (O_526,N_9674,N_6175);
nor UO_527 (O_527,N_6391,N_8673);
nand UO_528 (O_528,N_9692,N_9297);
nand UO_529 (O_529,N_8430,N_8859);
nand UO_530 (O_530,N_6326,N_7196);
or UO_531 (O_531,N_7788,N_8606);
or UO_532 (O_532,N_7766,N_9506);
or UO_533 (O_533,N_6340,N_8004);
or UO_534 (O_534,N_5659,N_8114);
and UO_535 (O_535,N_7052,N_7554);
or UO_536 (O_536,N_6365,N_7927);
and UO_537 (O_537,N_9277,N_8844);
nor UO_538 (O_538,N_5412,N_9997);
and UO_539 (O_539,N_8441,N_6676);
or UO_540 (O_540,N_9138,N_7081);
nand UO_541 (O_541,N_9615,N_6398);
and UO_542 (O_542,N_9460,N_9925);
nor UO_543 (O_543,N_5371,N_9964);
and UO_544 (O_544,N_7040,N_7000);
nor UO_545 (O_545,N_8336,N_6668);
or UO_546 (O_546,N_9726,N_9216);
nand UO_547 (O_547,N_5538,N_7666);
or UO_548 (O_548,N_5453,N_6397);
nor UO_549 (O_549,N_9893,N_8901);
and UO_550 (O_550,N_5556,N_6747);
or UO_551 (O_551,N_9742,N_8073);
or UO_552 (O_552,N_6267,N_8663);
and UO_553 (O_553,N_9265,N_7821);
nand UO_554 (O_554,N_8335,N_5874);
or UO_555 (O_555,N_9734,N_7398);
nor UO_556 (O_556,N_7566,N_7087);
nor UO_557 (O_557,N_8897,N_8287);
and UO_558 (O_558,N_7030,N_8660);
xor UO_559 (O_559,N_9948,N_8915);
and UO_560 (O_560,N_6685,N_8203);
and UO_561 (O_561,N_8153,N_8357);
nor UO_562 (O_562,N_6470,N_5634);
or UO_563 (O_563,N_8194,N_8236);
or UO_564 (O_564,N_8548,N_6817);
and UO_565 (O_565,N_6604,N_9656);
and UO_566 (O_566,N_9474,N_7729);
and UO_567 (O_567,N_6214,N_7225);
and UO_568 (O_568,N_7311,N_7705);
nor UO_569 (O_569,N_9932,N_7161);
nand UO_570 (O_570,N_9539,N_9207);
and UO_571 (O_571,N_8884,N_8597);
nand UO_572 (O_572,N_7618,N_7409);
and UO_573 (O_573,N_5450,N_8288);
or UO_574 (O_574,N_9559,N_7329);
xor UO_575 (O_575,N_5364,N_8134);
nand UO_576 (O_576,N_7001,N_5328);
nand UO_577 (O_577,N_8448,N_6568);
or UO_578 (O_578,N_8085,N_9940);
nand UO_579 (O_579,N_7317,N_6123);
or UO_580 (O_580,N_9235,N_9000);
xor UO_581 (O_581,N_7563,N_9594);
or UO_582 (O_582,N_5732,N_6318);
xnor UO_583 (O_583,N_7677,N_9142);
nor UO_584 (O_584,N_9830,N_6752);
and UO_585 (O_585,N_9245,N_7066);
nand UO_586 (O_586,N_6905,N_9754);
nand UO_587 (O_587,N_7617,N_9781);
nand UO_588 (O_588,N_6399,N_8955);
nand UO_589 (O_589,N_7162,N_8550);
nand UO_590 (O_590,N_8788,N_7894);
nand UO_591 (O_591,N_5368,N_9315);
xor UO_592 (O_592,N_8886,N_8254);
or UO_593 (O_593,N_6853,N_5164);
xnor UO_594 (O_594,N_5451,N_9897);
and UO_595 (O_595,N_7600,N_9185);
or UO_596 (O_596,N_7093,N_6704);
nand UO_597 (O_597,N_5719,N_9426);
xnor UO_598 (O_598,N_9275,N_9720);
nand UO_599 (O_599,N_7605,N_7342);
nand UO_600 (O_600,N_7106,N_9794);
or UO_601 (O_601,N_5145,N_7130);
nand UO_602 (O_602,N_9553,N_5275);
xor UO_603 (O_603,N_9840,N_7530);
or UO_604 (O_604,N_5905,N_8433);
or UO_605 (O_605,N_9466,N_9285);
xor UO_606 (O_606,N_9435,N_5510);
xnor UO_607 (O_607,N_5186,N_7527);
nand UO_608 (O_608,N_9763,N_7773);
xnor UO_609 (O_609,N_8564,N_7006);
or UO_610 (O_610,N_9478,N_5112);
xor UO_611 (O_611,N_8387,N_8670);
nand UO_612 (O_612,N_5303,N_5921);
or UO_613 (O_613,N_7239,N_6969);
and UO_614 (O_614,N_7544,N_5100);
and UO_615 (O_615,N_8622,N_9293);
and UO_616 (O_616,N_6045,N_5689);
and UO_617 (O_617,N_8512,N_6546);
nor UO_618 (O_618,N_6116,N_7895);
xor UO_619 (O_619,N_6087,N_7170);
or UO_620 (O_620,N_7348,N_6500);
nand UO_621 (O_621,N_7743,N_8656);
nor UO_622 (O_622,N_9483,N_8081);
nor UO_623 (O_623,N_9764,N_9201);
or UO_624 (O_624,N_6509,N_9440);
and UO_625 (O_625,N_6248,N_8559);
and UO_626 (O_626,N_6583,N_7913);
xnor UO_627 (O_627,N_5078,N_9247);
nor UO_628 (O_628,N_5557,N_8089);
nand UO_629 (O_629,N_8106,N_6778);
and UO_630 (O_630,N_6006,N_6041);
or UO_631 (O_631,N_5127,N_7681);
nor UO_632 (O_632,N_7521,N_7793);
nor UO_633 (O_633,N_8169,N_6602);
and UO_634 (O_634,N_8458,N_7307);
nor UO_635 (O_635,N_7708,N_6619);
or UO_636 (O_636,N_5720,N_7455);
and UO_637 (O_637,N_7993,N_7145);
or UO_638 (O_638,N_9725,N_9510);
nand UO_639 (O_639,N_7483,N_9511);
xor UO_640 (O_640,N_8667,N_7068);
xor UO_641 (O_641,N_5118,N_9307);
or UO_642 (O_642,N_7562,N_6498);
or UO_643 (O_643,N_5599,N_5315);
nand UO_644 (O_644,N_5665,N_9808);
or UO_645 (O_645,N_6502,N_8683);
or UO_646 (O_646,N_7011,N_9467);
nor UO_647 (O_647,N_8741,N_8083);
nand UO_648 (O_648,N_9040,N_7555);
xor UO_649 (O_649,N_5623,N_5052);
nand UO_650 (O_650,N_8309,N_8084);
xor UO_651 (O_651,N_6910,N_8996);
and UO_652 (O_652,N_9970,N_6448);
nand UO_653 (O_653,N_8381,N_6212);
nand UO_654 (O_654,N_9603,N_6349);
nor UO_655 (O_655,N_7989,N_8965);
or UO_656 (O_656,N_6514,N_9078);
and UO_657 (O_657,N_9564,N_5390);
nor UO_658 (O_658,N_7593,N_6143);
or UO_659 (O_659,N_5196,N_8030);
nand UO_660 (O_660,N_6980,N_8614);
nand UO_661 (O_661,N_6136,N_8312);
or UO_662 (O_662,N_7454,N_6435);
nand UO_663 (O_663,N_5580,N_5225);
nor UO_664 (O_664,N_9952,N_9666);
nand UO_665 (O_665,N_6995,N_9065);
or UO_666 (O_666,N_9036,N_5875);
and UO_667 (O_667,N_5646,N_7233);
nor UO_668 (O_668,N_9612,N_6729);
nand UO_669 (O_669,N_6024,N_9805);
nor UO_670 (O_670,N_7688,N_7014);
or UO_671 (O_671,N_7950,N_9947);
or UO_672 (O_672,N_5184,N_6347);
and UO_673 (O_673,N_8846,N_7222);
or UO_674 (O_674,N_6074,N_8204);
nand UO_675 (O_675,N_9670,N_9644);
nand UO_676 (O_676,N_9665,N_5389);
or UO_677 (O_677,N_7921,N_5261);
nor UO_678 (O_678,N_5664,N_5962);
and UO_679 (O_679,N_6450,N_6408);
xnor UO_680 (O_680,N_6610,N_7616);
xnor UO_681 (O_681,N_5918,N_5143);
xor UO_682 (O_682,N_6998,N_9006);
or UO_683 (O_683,N_6694,N_5965);
nor UO_684 (O_684,N_8118,N_6526);
nor UO_685 (O_685,N_7266,N_5044);
and UO_686 (O_686,N_7840,N_5988);
and UO_687 (O_687,N_5331,N_5361);
nor UO_688 (O_688,N_6928,N_6249);
or UO_689 (O_689,N_8266,N_9768);
or UO_690 (O_690,N_9300,N_8733);
and UO_691 (O_691,N_7753,N_9427);
nor UO_692 (O_692,N_5761,N_5520);
or UO_693 (O_693,N_6897,N_6744);
nor UO_694 (O_694,N_9060,N_6454);
xnor UO_695 (O_695,N_9472,N_9099);
and UO_696 (O_696,N_5101,N_8491);
or UO_697 (O_697,N_8063,N_6821);
or UO_698 (O_698,N_5690,N_6037);
xor UO_699 (O_699,N_9354,N_5868);
and UO_700 (O_700,N_9810,N_8038);
or UO_701 (O_701,N_7420,N_9093);
nand UO_702 (O_702,N_8132,N_8653);
nor UO_703 (O_703,N_9652,N_7335);
nand UO_704 (O_704,N_8536,N_8909);
nand UO_705 (O_705,N_6737,N_7508);
nand UO_706 (O_706,N_6081,N_6276);
nand UO_707 (O_707,N_5263,N_7934);
or UO_708 (O_708,N_8080,N_9713);
nand UO_709 (O_709,N_9593,N_6390);
or UO_710 (O_710,N_7273,N_5202);
and UO_711 (O_711,N_8056,N_6352);
nand UO_712 (O_712,N_7056,N_6641);
or UO_713 (O_713,N_8925,N_8590);
nor UO_714 (O_714,N_6986,N_8946);
or UO_715 (O_715,N_6363,N_8463);
nor UO_716 (O_716,N_9392,N_8374);
or UO_717 (O_717,N_9738,N_5010);
xnor UO_718 (O_718,N_7260,N_9497);
or UO_719 (O_719,N_6475,N_6757);
xor UO_720 (O_720,N_9148,N_7312);
or UO_721 (O_721,N_7031,N_7524);
or UO_722 (O_722,N_5565,N_7088);
nand UO_723 (O_723,N_6999,N_7706);
xnor UO_724 (O_724,N_6193,N_6395);
nand UO_725 (O_725,N_9633,N_9744);
and UO_726 (O_726,N_6462,N_6686);
nand UO_727 (O_727,N_6891,N_7316);
nand UO_728 (O_728,N_9203,N_9191);
xor UO_729 (O_729,N_5284,N_9512);
and UO_730 (O_730,N_7976,N_6080);
nand UO_731 (O_731,N_8784,N_9147);
or UO_732 (O_732,N_5472,N_5866);
or UO_733 (O_733,N_6776,N_9934);
nor UO_734 (O_734,N_9169,N_6296);
nand UO_735 (O_735,N_7937,N_8926);
nand UO_736 (O_736,N_7264,N_6540);
or UO_737 (O_737,N_8875,N_5851);
nor UO_738 (O_738,N_6355,N_7819);
or UO_739 (O_739,N_5324,N_6628);
nand UO_740 (O_740,N_6472,N_5405);
xor UO_741 (O_741,N_7956,N_9393);
and UO_742 (O_742,N_7321,N_7135);
and UO_743 (O_743,N_7614,N_5947);
nor UO_744 (O_744,N_5631,N_9433);
and UO_745 (O_745,N_6312,N_6480);
xnor UO_746 (O_746,N_8657,N_6530);
or UO_747 (O_747,N_8049,N_6711);
nor UO_748 (O_748,N_9702,N_9913);
nor UO_749 (O_749,N_6703,N_7154);
xor UO_750 (O_750,N_9756,N_8679);
and UO_751 (O_751,N_8110,N_6150);
or UO_752 (O_752,N_5431,N_7830);
or UO_753 (O_753,N_8492,N_5176);
nor UO_754 (O_754,N_9688,N_6287);
and UO_755 (O_755,N_5305,N_6783);
and UO_756 (O_756,N_9153,N_9617);
and UO_757 (O_757,N_6466,N_5794);
nor UO_758 (O_758,N_6835,N_9817);
nand UO_759 (O_759,N_5906,N_8829);
nand UO_760 (O_760,N_8539,N_8112);
nand UO_761 (O_761,N_5140,N_5304);
and UO_762 (O_762,N_7540,N_6634);
and UO_763 (O_763,N_6968,N_8553);
and UO_764 (O_764,N_7228,N_7902);
and UO_765 (O_765,N_9498,N_5682);
or UO_766 (O_766,N_6366,N_8600);
nand UO_767 (O_767,N_9132,N_8827);
or UO_768 (O_768,N_9786,N_5977);
and UO_769 (O_769,N_7033,N_5157);
xnor UO_770 (O_770,N_5724,N_9043);
or UO_771 (O_771,N_5212,N_8972);
xor UO_772 (O_772,N_5891,N_8366);
xor UO_773 (O_773,N_8413,N_7970);
and UO_774 (O_774,N_8376,N_7643);
nor UO_775 (O_775,N_6551,N_9655);
nand UO_776 (O_776,N_5574,N_7610);
nand UO_777 (O_777,N_8770,N_5034);
xor UO_778 (O_778,N_6658,N_9599);
nor UO_779 (O_779,N_8995,N_5465);
or UO_780 (O_780,N_8690,N_7490);
xor UO_781 (O_781,N_5877,N_8002);
nand UO_782 (O_782,N_9096,N_9431);
nor UO_783 (O_783,N_5247,N_9320);
or UO_784 (O_784,N_7776,N_9079);
nor UO_785 (O_785,N_9179,N_5420);
and UO_786 (O_786,N_7347,N_5485);
or UO_787 (O_787,N_9387,N_7166);
xnor UO_788 (O_788,N_7501,N_8377);
or UO_789 (O_789,N_7531,N_6260);
nand UO_790 (O_790,N_5562,N_6674);
nand UO_791 (O_791,N_9673,N_5220);
or UO_792 (O_792,N_9982,N_8864);
nor UO_793 (O_793,N_6559,N_7838);
nand UO_794 (O_794,N_9766,N_9456);
and UO_795 (O_795,N_7182,N_6877);
nor UO_796 (O_796,N_8019,N_6819);
nor UO_797 (O_797,N_6534,N_7844);
or UO_798 (O_798,N_8469,N_7604);
xnor UO_799 (O_799,N_5758,N_9849);
and UO_800 (O_800,N_5703,N_7430);
nand UO_801 (O_801,N_8071,N_8645);
and UO_802 (O_802,N_7667,N_8528);
xor UO_803 (O_803,N_6643,N_7229);
or UO_804 (O_804,N_7257,N_5514);
nand UO_805 (O_805,N_9588,N_5430);
nand UO_806 (O_806,N_5391,N_6791);
nand UO_807 (O_807,N_5948,N_9825);
or UO_808 (O_808,N_8199,N_6491);
nor UO_809 (O_809,N_5811,N_7880);
xor UO_810 (O_810,N_5677,N_9046);
nor UO_811 (O_811,N_7245,N_8241);
nor UO_812 (O_812,N_8272,N_5865);
and UO_813 (O_813,N_7754,N_7259);
nand UO_814 (O_814,N_7583,N_5823);
and UO_815 (O_815,N_7126,N_5663);
and UO_816 (O_816,N_9520,N_9197);
xor UO_817 (O_817,N_5589,N_6979);
xnor UO_818 (O_818,N_9218,N_9570);
and UO_819 (O_819,N_6458,N_6631);
nor UO_820 (O_820,N_6605,N_8445);
xnor UO_821 (O_821,N_8117,N_8596);
nand UO_822 (O_822,N_6111,N_7623);
and UO_823 (O_823,N_7089,N_8845);
nor UO_824 (O_824,N_9532,N_7709);
nor UO_825 (O_825,N_7911,N_9791);
and UO_826 (O_826,N_7350,N_6904);
nand UO_827 (O_827,N_6453,N_6309);
xnor UO_828 (O_828,N_9067,N_5214);
nor UO_829 (O_829,N_5814,N_7134);
nor UO_830 (O_830,N_5695,N_9628);
nand UO_831 (O_831,N_6001,N_9358);
nor UO_832 (O_832,N_6896,N_6452);
nand UO_833 (O_833,N_6468,N_8044);
nor UO_834 (O_834,N_6794,N_6173);
xor UO_835 (O_835,N_9751,N_9585);
nor UO_836 (O_836,N_7291,N_6815);
xor UO_837 (O_837,N_5373,N_6376);
nand UO_838 (O_838,N_6262,N_8994);
and UO_839 (O_839,N_6761,N_5497);
nor UO_840 (O_840,N_9168,N_8005);
nor UO_841 (O_841,N_8401,N_7109);
or UO_842 (O_842,N_9106,N_5594);
nor UO_843 (O_843,N_5298,N_9035);
and UO_844 (O_844,N_8724,N_5577);
nor UO_845 (O_845,N_9329,N_5919);
nor UO_846 (O_846,N_8619,N_6901);
and UO_847 (O_847,N_7848,N_8866);
nor UO_848 (O_848,N_9667,N_5771);
nor UO_849 (O_849,N_7417,N_8361);
xor UO_850 (O_850,N_7217,N_5237);
nand UO_851 (O_851,N_9682,N_5048);
or UO_852 (O_852,N_8353,N_5239);
nand UO_853 (O_853,N_9353,N_8224);
nor UO_854 (O_854,N_6259,N_5700);
nor UO_855 (O_855,N_7608,N_7158);
or UO_856 (O_856,N_6483,N_6430);
xnor UO_857 (O_857,N_9503,N_6837);
nor UO_858 (O_858,N_8592,N_7866);
nand UO_859 (O_859,N_9629,N_8202);
or UO_860 (O_860,N_8060,N_5745);
nand UO_861 (O_861,N_9258,N_7476);
xor UO_862 (O_862,N_9905,N_8910);
nor UO_863 (O_863,N_6920,N_6328);
nand UO_864 (O_864,N_8964,N_7488);
or UO_865 (O_865,N_6303,N_6301);
and UO_866 (O_866,N_8865,N_9716);
xor UO_867 (O_867,N_7213,N_6698);
xnor UO_868 (O_868,N_5857,N_6976);
or UO_869 (O_869,N_8971,N_7626);
nand UO_870 (O_870,N_5938,N_9009);
and UO_871 (O_871,N_8969,N_6050);
or UO_872 (O_872,N_7280,N_9236);
and UO_873 (O_873,N_6706,N_6099);
nor UO_874 (O_874,N_8258,N_8616);
and UO_875 (O_875,N_7344,N_5444);
or UO_876 (O_876,N_8707,N_5778);
or UO_877 (O_877,N_9031,N_6078);
nor UO_878 (O_878,N_9212,N_5669);
or UO_879 (O_879,N_5870,N_9687);
or UO_880 (O_880,N_6743,N_8981);
nor UO_881 (O_881,N_8576,N_7697);
nor UO_882 (O_882,N_7057,N_5153);
or UO_883 (O_883,N_9748,N_7301);
xnor UO_884 (O_884,N_6930,N_5579);
or UO_885 (O_885,N_5258,N_8126);
nand UO_886 (O_886,N_8420,N_9033);
xnor UO_887 (O_887,N_9663,N_6093);
xnor UO_888 (O_888,N_9417,N_8489);
or UO_889 (O_889,N_9954,N_6931);
xor UO_890 (O_890,N_8584,N_9923);
or UO_891 (O_891,N_5946,N_5725);
or UO_892 (O_892,N_8517,N_7810);
or UO_893 (O_893,N_6121,N_5555);
nand UO_894 (O_894,N_6237,N_5764);
nor UO_895 (O_895,N_5616,N_5648);
xor UO_896 (O_896,N_7963,N_7370);
or UO_897 (O_897,N_6216,N_8675);
nor UO_898 (O_898,N_5711,N_5674);
xnor UO_899 (O_899,N_8302,N_7340);
or UO_900 (O_900,N_7411,N_9121);
nor UO_901 (O_901,N_6140,N_8522);
xor UO_902 (O_902,N_5124,N_5612);
nor UO_903 (O_903,N_9295,N_6669);
nor UO_904 (O_904,N_7253,N_8710);
or UO_905 (O_905,N_6198,N_6872);
and UO_906 (O_906,N_5296,N_9441);
nand UO_907 (O_907,N_9668,N_7552);
xnor UO_908 (O_908,N_5025,N_6192);
nand UO_909 (O_909,N_5518,N_8776);
or UO_910 (O_910,N_5849,N_5336);
nor UO_911 (O_911,N_5480,N_8195);
nor UO_912 (O_912,N_6499,N_9076);
nor UO_913 (O_913,N_6103,N_9188);
nor UO_914 (O_914,N_9311,N_8289);
or UO_915 (O_915,N_6059,N_7480);
xor UO_916 (O_916,N_6884,N_6941);
and UO_917 (O_917,N_5053,N_5023);
and UO_918 (O_918,N_9240,N_8508);
xnor UO_919 (O_919,N_5146,N_7294);
and UO_920 (O_920,N_6527,N_5813);
and UO_921 (O_921,N_8970,N_8939);
or UO_922 (O_922,N_6515,N_9219);
xor UO_923 (O_923,N_6987,N_8470);
nor UO_924 (O_924,N_9892,N_6809);
or UO_925 (O_925,N_6645,N_6665);
or UO_926 (O_926,N_6562,N_6179);
nor UO_927 (O_927,N_8560,N_6699);
and UO_928 (O_928,N_9457,N_5163);
xnor UO_929 (O_929,N_6774,N_7059);
nor UO_930 (O_930,N_8193,N_7856);
nor UO_931 (O_931,N_8985,N_6158);
or UO_932 (O_932,N_8885,N_6594);
nor UO_933 (O_933,N_7433,N_6595);
or UO_934 (O_934,N_6556,N_8635);
and UO_935 (O_935,N_5427,N_6255);
nand UO_936 (O_936,N_5382,N_9437);
and UO_937 (O_937,N_8903,N_6058);
nor UO_938 (O_938,N_7122,N_9533);
nand UO_939 (O_939,N_5418,N_7971);
nor UO_940 (O_940,N_9894,N_6929);
nand UO_941 (O_941,N_8691,N_9057);
nand UO_942 (O_942,N_9600,N_7438);
nor UO_943 (O_943,N_5883,N_9476);
or UO_944 (O_944,N_9414,N_6266);
and UO_945 (O_945,N_8141,N_7738);
or UO_946 (O_946,N_6611,N_9676);
nand UO_947 (O_947,N_6289,N_7128);
xnor UO_948 (O_948,N_9023,N_8086);
nand UO_949 (O_949,N_8410,N_5707);
nand UO_950 (O_950,N_9049,N_5923);
nand UO_951 (O_951,N_5410,N_6816);
or UO_952 (O_952,N_6094,N_6681);
nor UO_953 (O_953,N_8764,N_7576);
nor UO_954 (O_954,N_5359,N_7315);
and UO_955 (O_955,N_7505,N_7111);
nor UO_956 (O_956,N_9015,N_9445);
or UO_957 (O_957,N_9992,N_6288);
nor UO_958 (O_958,N_9648,N_8279);
nor UO_959 (O_959,N_8334,N_6054);
nor UO_960 (O_960,N_8975,N_8919);
xor UO_961 (O_961,N_5054,N_5899);
and UO_962 (O_962,N_6068,N_5370);
or UO_963 (O_963,N_5452,N_8695);
nor UO_964 (O_964,N_5180,N_6576);
xnor UO_965 (O_965,N_8345,N_6371);
nand UO_966 (O_966,N_9639,N_7586);
nor UO_967 (O_967,N_9685,N_5924);
nor UO_968 (O_968,N_8745,N_7207);
nor UO_969 (O_969,N_7216,N_5830);
or UO_970 (O_970,N_6864,N_6437);
and UO_971 (O_971,N_8604,N_9150);
xnor UO_972 (O_972,N_6590,N_9608);
nand UO_973 (O_973,N_7022,N_9238);
or UO_974 (O_974,N_7736,N_7306);
nor UO_975 (O_975,N_9845,N_6876);
and UO_976 (O_976,N_6948,N_9112);
nor UO_977 (O_977,N_6806,N_5460);
xnor UO_978 (O_978,N_6714,N_7855);
and UO_979 (O_979,N_7946,N_9400);
and UO_980 (O_980,N_6005,N_9013);
nand UO_981 (O_981,N_8444,N_5736);
nor UO_982 (O_982,N_5064,N_5662);
and UO_983 (O_983,N_9660,N_6831);
and UO_984 (O_984,N_5578,N_8183);
or UO_985 (O_985,N_9522,N_6432);
and UO_986 (O_986,N_6726,N_7214);
and UO_987 (O_987,N_5559,N_6845);
or UO_988 (O_988,N_9493,N_5817);
or UO_989 (O_989,N_7459,N_9237);
xor UO_990 (O_990,N_9527,N_5027);
and UO_991 (O_991,N_5608,N_7358);
nand UO_992 (O_992,N_9128,N_8108);
nand UO_993 (O_993,N_9977,N_9745);
xnor UO_994 (O_994,N_7715,N_9100);
nor UO_995 (O_995,N_5422,N_6367);
nand UO_996 (O_996,N_8423,N_6560);
or UO_997 (O_997,N_7116,N_8046);
nand UO_998 (O_998,N_6282,N_9439);
and UO_999 (O_999,N_7678,N_9868);
nor UO_1000 (O_1000,N_8993,N_8810);
nand UO_1001 (O_1001,N_8435,N_7648);
or UO_1002 (O_1002,N_6247,N_9715);
nor UO_1003 (O_1003,N_8464,N_8944);
nor UO_1004 (O_1004,N_5233,N_6950);
and UO_1005 (O_1005,N_9377,N_8755);
nand UO_1006 (O_1006,N_7941,N_6100);
nand UO_1007 (O_1007,N_6131,N_7787);
xnor UO_1008 (O_1008,N_8341,N_7448);
nor UO_1009 (O_1009,N_8530,N_7379);
nor UO_1010 (O_1010,N_8726,N_6504);
nor UO_1011 (O_1011,N_5007,N_6949);
and UO_1012 (O_1012,N_7526,N_6258);
and UO_1013 (O_1013,N_6088,N_5232);
and UO_1014 (O_1014,N_5091,N_8006);
or UO_1015 (O_1015,N_9936,N_6939);
nor UO_1016 (O_1016,N_9038,N_8870);
nand UO_1017 (O_1017,N_7007,N_6780);
nor UO_1018 (O_1018,N_9907,N_5194);
and UO_1019 (O_1019,N_9989,N_9193);
xnor UO_1020 (O_1020,N_5227,N_9159);
nor UO_1021 (O_1021,N_7839,N_9366);
and UO_1022 (O_1022,N_9459,N_8629);
or UO_1023 (O_1023,N_6554,N_9434);
or UO_1024 (O_1024,N_6916,N_5080);
or UO_1025 (O_1025,N_9864,N_5248);
nand UO_1026 (O_1026,N_7966,N_7537);
or UO_1027 (O_1027,N_8375,N_8417);
and UO_1028 (O_1028,N_7194,N_7804);
nor UO_1029 (O_1029,N_9949,N_8262);
or UO_1030 (O_1030,N_8933,N_7932);
and UO_1031 (O_1031,N_7247,N_8871);
and UO_1032 (O_1032,N_9443,N_5971);
or UO_1033 (O_1033,N_9709,N_7701);
xor UO_1034 (O_1034,N_7557,N_6563);
or UO_1035 (O_1035,N_7083,N_9429);
nand UO_1036 (O_1036,N_6724,N_9942);
nor UO_1037 (O_1037,N_6447,N_5543);
nor UO_1038 (O_1038,N_7325,N_7573);
nand UO_1039 (O_1039,N_5312,N_7831);
and UO_1040 (O_1040,N_9981,N_8677);
nor UO_1041 (O_1041,N_8243,N_7664);
and UO_1042 (O_1042,N_9635,N_9428);
nand UO_1043 (O_1043,N_7039,N_5958);
and UO_1044 (O_1044,N_6033,N_9374);
nor UO_1045 (O_1045,N_7027,N_6616);
nand UO_1046 (O_1046,N_5154,N_8817);
or UO_1047 (O_1047,N_6798,N_7744);
and UO_1048 (O_1048,N_6679,N_6887);
or UO_1049 (O_1049,N_7309,N_7534);
nor UO_1050 (O_1050,N_5062,N_7636);
nand UO_1051 (O_1051,N_5350,N_7574);
or UO_1052 (O_1052,N_5696,N_5403);
nor UO_1053 (O_1053,N_6279,N_9884);
xnor UO_1054 (O_1054,N_9903,N_7103);
and UO_1055 (O_1055,N_5325,N_7378);
nor UO_1056 (O_1056,N_8148,N_5079);
nand UO_1057 (O_1057,N_6646,N_8189);
or UO_1058 (O_1058,N_7673,N_8519);
xnor UO_1059 (O_1059,N_7457,N_6012);
and UO_1060 (O_1060,N_5415,N_6844);
xor UO_1061 (O_1061,N_7276,N_8099);
or UO_1062 (O_1062,N_8095,N_6443);
nor UO_1063 (O_1063,N_5433,N_6719);
nor UO_1064 (O_1064,N_7767,N_8850);
nand UO_1065 (O_1065,N_6323,N_7746);
or UO_1066 (O_1066,N_5838,N_7539);
nand UO_1067 (O_1067,N_6239,N_8526);
and UO_1068 (O_1068,N_7837,N_5486);
xor UO_1069 (O_1069,N_8061,N_8207);
nor UO_1070 (O_1070,N_5837,N_6678);
nor UO_1071 (O_1071,N_7399,N_7439);
or UO_1072 (O_1072,N_9757,N_8384);
and UO_1073 (O_1073,N_8781,N_8488);
and UO_1074 (O_1074,N_8187,N_9590);
nor UO_1075 (O_1075,N_8627,N_7808);
or UO_1076 (O_1076,N_9634,N_9871);
and UO_1077 (O_1077,N_5776,N_8496);
nand UO_1078 (O_1078,N_7723,N_6833);
nor UO_1079 (O_1079,N_7133,N_6127);
nand UO_1080 (O_1080,N_8283,N_8934);
or UO_1081 (O_1081,N_8977,N_9014);
xnor UO_1082 (O_1082,N_5769,N_5821);
nand UO_1083 (O_1083,N_8115,N_9821);
nor UO_1084 (O_1084,N_7676,N_7731);
and UO_1085 (O_1085,N_5882,N_9961);
nand UO_1086 (O_1086,N_5753,N_8852);
and UO_1087 (O_1087,N_8942,N_9327);
or UO_1088 (O_1088,N_7899,N_6802);
and UO_1089 (O_1089,N_7098,N_5138);
or UO_1090 (O_1090,N_5963,N_7561);
nor UO_1091 (O_1091,N_6940,N_6978);
and UO_1092 (O_1092,N_6733,N_9382);
and UO_1093 (O_1093,N_9171,N_5847);
nand UO_1094 (O_1094,N_5553,N_5179);
nand UO_1095 (O_1095,N_6661,N_8107);
nor UO_1096 (O_1096,N_9473,N_5942);
and UO_1097 (O_1097,N_9518,N_9710);
xor UO_1098 (O_1098,N_8338,N_6438);
or UO_1099 (O_1099,N_6564,N_7777);
nor UO_1100 (O_1100,N_5455,N_7772);
nand UO_1101 (O_1101,N_6553,N_5086);
or UO_1102 (O_1102,N_5257,N_5221);
xnor UO_1103 (O_1103,N_5094,N_8481);
nand UO_1104 (O_1104,N_6205,N_7223);
and UO_1105 (O_1105,N_6387,N_7019);
or UO_1106 (O_1106,N_9995,N_8943);
nand UO_1107 (O_1107,N_5104,N_9831);
nand UO_1108 (O_1108,N_6487,N_5092);
or UO_1109 (O_1109,N_9302,N_7813);
and UO_1110 (O_1110,N_8250,N_8018);
nand UO_1111 (O_1111,N_6015,N_6652);
or UO_1112 (O_1112,N_9367,N_5654);
and UO_1113 (O_1113,N_8744,N_5638);
or UO_1114 (O_1114,N_7512,N_6636);
xnor UO_1115 (O_1115,N_5560,N_6342);
nand UO_1116 (O_1116,N_7286,N_8208);
nand UO_1117 (O_1117,N_7495,N_9993);
nor UO_1118 (O_1118,N_7790,N_8881);
nor UO_1119 (O_1119,N_6208,N_5024);
and UO_1120 (O_1120,N_8703,N_9464);
or UO_1121 (O_1121,N_8911,N_5981);
and UO_1122 (O_1122,N_6224,N_7955);
nor UO_1123 (O_1123,N_7835,N_7497);
and UO_1124 (O_1124,N_6508,N_8438);
nand UO_1125 (O_1125,N_8391,N_8763);
nor UO_1126 (O_1126,N_7461,N_6505);
and UO_1127 (O_1127,N_5524,N_8937);
or UO_1128 (O_1128,N_6520,N_6226);
or UO_1129 (O_1129,N_9391,N_8454);
nand UO_1130 (O_1130,N_9162,N_7496);
nand UO_1131 (O_1131,N_9915,N_5889);
nor UO_1132 (O_1132,N_8296,N_7924);
nand UO_1133 (O_1133,N_8161,N_5022);
and UO_1134 (O_1134,N_8035,N_7463);
and UO_1135 (O_1135,N_7186,N_6310);
nand UO_1136 (O_1136,N_6236,N_7638);
nand UO_1137 (O_1137,N_5477,N_7599);
nor UO_1138 (O_1138,N_7797,N_8156);
and UO_1139 (O_1139,N_6402,N_8192);
or UO_1140 (O_1140,N_9011,N_7240);
or UO_1141 (O_1141,N_5400,N_8520);
xnor UO_1142 (O_1142,N_5789,N_5926);
xor UO_1143 (O_1143,N_6320,N_8346);
and UO_1144 (O_1144,N_7549,N_6959);
or UO_1145 (O_1145,N_9156,N_6025);
and UO_1146 (O_1146,N_6511,N_6673);
or UO_1147 (O_1147,N_5429,N_6654);
and UO_1148 (O_1148,N_6251,N_5864);
or UO_1149 (O_1149,N_6016,N_6667);
nor UO_1150 (O_1150,N_8637,N_7822);
nand UO_1151 (O_1151,N_8642,N_6166);
nor UO_1152 (O_1152,N_6412,N_6852);
and UO_1153 (O_1153,N_7034,N_7525);
xor UO_1154 (O_1154,N_6640,N_6664);
nor UO_1155 (O_1155,N_6065,N_5387);
or UO_1156 (O_1156,N_9325,N_5219);
xnor UO_1157 (O_1157,N_7432,N_9208);
xor UO_1158 (O_1158,N_7988,N_5566);
nand UO_1159 (O_1159,N_8694,N_8768);
nand UO_1160 (O_1160,N_9632,N_9727);
or UO_1161 (O_1161,N_6519,N_9039);
or UO_1162 (O_1162,N_5229,N_5759);
nor UO_1163 (O_1163,N_8716,N_8672);
and UO_1164 (O_1164,N_6859,N_5029);
or UO_1165 (O_1165,N_7517,N_5075);
and UO_1166 (O_1166,N_5335,N_9696);
or UO_1167 (O_1167,N_7475,N_6687);
and UO_1168 (O_1168,N_6243,N_5668);
nor UO_1169 (O_1169,N_6072,N_5015);
nand UO_1170 (O_1170,N_8457,N_7654);
and UO_1171 (O_1171,N_6862,N_9224);
nor UO_1172 (O_1172,N_9027,N_9813);
nand UO_1173 (O_1173,N_8337,N_5149);
and UO_1174 (O_1174,N_5743,N_9609);
or UO_1175 (O_1175,N_7814,N_5107);
and UO_1176 (O_1176,N_7796,N_9215);
xnor UO_1177 (O_1177,N_6770,N_9042);
xor UO_1178 (O_1178,N_6441,N_5885);
and UO_1179 (O_1179,N_7811,N_6967);
or UO_1180 (O_1180,N_6449,N_8212);
and UO_1181 (O_1181,N_8756,N_6434);
nand UO_1182 (O_1182,N_5291,N_5033);
nand UO_1183 (O_1183,N_9853,N_7132);
and UO_1184 (O_1184,N_5705,N_8143);
xor UO_1185 (O_1185,N_9779,N_8973);
and UO_1186 (O_1186,N_8795,N_5529);
and UO_1187 (O_1187,N_8525,N_8573);
nor UO_1188 (O_1188,N_8737,N_7940);
nor UO_1189 (O_1189,N_7211,N_6436);
nor UO_1190 (O_1190,N_9268,N_6295);
nor UO_1191 (O_1191,N_5835,N_6900);
nand UO_1192 (O_1192,N_6684,N_5469);
and UO_1193 (O_1193,N_9998,N_8978);
or UO_1194 (O_1194,N_5713,N_7669);
nand UO_1195 (O_1195,N_9679,N_6281);
nand UO_1196 (O_1196,N_7984,N_7854);
and UO_1197 (O_1197,N_9017,N_8077);
and UO_1198 (O_1198,N_8701,N_8495);
xnor UO_1199 (O_1199,N_9357,N_5726);
nand UO_1200 (O_1200,N_9287,N_9746);
xor UO_1201 (O_1201,N_9411,N_9803);
or UO_1202 (O_1202,N_8432,N_9610);
nor UO_1203 (O_1203,N_9452,N_9637);
and UO_1204 (O_1204,N_9597,N_7295);
nand UO_1205 (O_1205,N_7474,N_9194);
or UO_1206 (O_1206,N_7852,N_8711);
nand UO_1207 (O_1207,N_7422,N_9222);
or UO_1208 (O_1208,N_7046,N_5681);
nand UO_1209 (O_1209,N_8249,N_6865);
nand UO_1210 (O_1210,N_8957,N_8039);
nor UO_1211 (O_1211,N_8595,N_5017);
nand UO_1212 (O_1212,N_9505,N_6735);
or UO_1213 (O_1213,N_6596,N_7502);
and UO_1214 (O_1214,N_8227,N_9924);
nor UO_1215 (O_1215,N_8443,N_8789);
or UO_1216 (O_1216,N_8268,N_6182);
or UO_1217 (O_1217,N_7443,N_6298);
and UO_1218 (O_1218,N_8415,N_9809);
nand UO_1219 (O_1219,N_7874,N_9852);
nor UO_1220 (O_1220,N_5742,N_6824);
or UO_1221 (O_1221,N_6271,N_8386);
or UO_1222 (O_1222,N_8686,N_6013);
or UO_1223 (O_1223,N_5395,N_8411);
nor UO_1224 (O_1224,N_7682,N_8807);
or UO_1225 (O_1225,N_9239,N_9780);
or UO_1226 (O_1226,N_5827,N_8535);
nor UO_1227 (O_1227,N_9029,N_6785);
and UO_1228 (O_1228,N_7764,N_5001);
and UO_1229 (O_1229,N_5031,N_5994);
nand UO_1230 (O_1230,N_5546,N_6782);
or UO_1231 (O_1231,N_8372,N_8295);
or UO_1232 (O_1232,N_5105,N_8200);
nor UO_1233 (O_1233,N_7487,N_7789);
or UO_1234 (O_1234,N_7047,N_7436);
xor UO_1235 (O_1235,N_5960,N_8011);
and UO_1236 (O_1236,N_9074,N_7005);
xor UO_1237 (O_1237,N_7377,N_8406);
nor UO_1238 (O_1238,N_5087,N_6836);
nor UO_1239 (O_1239,N_9877,N_8839);
nor UO_1240 (O_1240,N_5542,N_8007);
or UO_1241 (O_1241,N_5251,N_8652);
nor UO_1242 (O_1242,N_8945,N_6850);
nand UO_1243 (O_1243,N_5035,N_5843);
nor UO_1244 (O_1244,N_8516,N_9776);
nor UO_1245 (O_1245,N_7353,N_6578);
nor UO_1246 (O_1246,N_5414,N_7592);
nand UO_1247 (O_1247,N_7580,N_7356);
nor UO_1248 (O_1248,N_7641,N_6252);
or UO_1249 (O_1249,N_7930,N_8990);
xor UO_1250 (O_1250,N_9080,N_7725);
and UO_1251 (O_1251,N_7873,N_8300);
xnor UO_1252 (O_1252,N_9088,N_5936);
or UO_1253 (O_1253,N_5508,N_7200);
and UO_1254 (O_1254,N_6874,N_9839);
or UO_1255 (O_1255,N_8228,N_7556);
nor UO_1256 (O_1256,N_5366,N_7394);
or UO_1257 (O_1257,N_7292,N_7684);
nand UO_1258 (O_1258,N_5352,N_5012);
nor UO_1259 (O_1259,N_6557,N_9819);
nand UO_1260 (O_1260,N_5746,N_9328);
and UO_1261 (O_1261,N_6079,N_9728);
nor UO_1262 (O_1262,N_5917,N_5642);
nand UO_1263 (O_1263,N_8639,N_5122);
nor UO_1264 (O_1264,N_6154,N_7694);
xnor UO_1265 (O_1265,N_5160,N_9133);
xnor UO_1266 (O_1266,N_9202,N_8625);
nor UO_1267 (O_1267,N_9606,N_6620);
nand UO_1268 (O_1268,N_7933,N_8284);
nor UO_1269 (O_1269,N_5779,N_6649);
nand UO_1270 (O_1270,N_8589,N_6772);
nand UO_1271 (O_1271,N_5175,N_5792);
or UO_1272 (O_1272,N_9250,N_7078);
or UO_1273 (O_1273,N_7173,N_6018);
nand UO_1274 (O_1274,N_7267,N_8728);
or UO_1275 (O_1275,N_5536,N_7882);
nand UO_1276 (O_1276,N_8456,N_5197);
or UO_1277 (O_1277,N_7415,N_9044);
or UO_1278 (O_1278,N_8758,N_6971);
and UO_1279 (O_1279,N_7510,N_5730);
nand UO_1280 (O_1280,N_9204,N_8557);
or UO_1281 (O_1281,N_7184,N_5959);
nand UO_1282 (O_1282,N_5643,N_8075);
nor UO_1283 (O_1283,N_8940,N_8922);
or UO_1284 (O_1284,N_6138,N_9161);
nor UO_1285 (O_1285,N_6440,N_7869);
nor UO_1286 (O_1286,N_8696,N_7492);
xnor UO_1287 (O_1287,N_9183,N_9519);
or UO_1288 (O_1288,N_5819,N_8654);
nor UO_1289 (O_1289,N_8149,N_5026);
or UO_1290 (O_1290,N_6539,N_8687);
and UO_1291 (O_1291,N_8164,N_9664);
xor UO_1292 (O_1292,N_7803,N_8772);
nand UO_1293 (O_1293,N_8921,N_8760);
or UO_1294 (O_1294,N_5533,N_7570);
xnor UO_1295 (O_1295,N_7362,N_8568);
nand UO_1296 (O_1296,N_5036,N_7227);
nand UO_1297 (O_1297,N_5503,N_9717);
nor UO_1298 (O_1298,N_6132,N_9432);
nand UO_1299 (O_1299,N_5993,N_7990);
nand UO_1300 (O_1300,N_5182,N_7471);
and UO_1301 (O_1301,N_6923,N_6606);
nand UO_1302 (O_1302,N_7890,N_9691);
nand UO_1303 (O_1303,N_6840,N_9846);
or UO_1304 (O_1304,N_8821,N_5990);
nor UO_1305 (O_1305,N_5997,N_8791);
and UO_1306 (O_1306,N_9812,N_5408);
nor UO_1307 (O_1307,N_7791,N_8851);
nor UO_1308 (O_1308,N_7405,N_8388);
xor UO_1309 (O_1309,N_7084,N_7156);
and UO_1310 (O_1310,N_7782,N_9782);
nor UO_1311 (O_1311,N_8613,N_5673);
nand UO_1312 (O_1312,N_7175,N_5306);
nor UO_1313 (O_1313,N_9950,N_5716);
xor UO_1314 (O_1314,N_8623,N_7572);
nor UO_1315 (O_1315,N_7675,N_5377);
or UO_1316 (O_1316,N_8917,N_9041);
or UO_1317 (O_1317,N_7410,N_9131);
and UO_1318 (O_1318,N_6410,N_5568);
and UO_1319 (O_1319,N_5816,N_5869);
nand UO_1320 (O_1320,N_9330,N_8276);
nor UO_1321 (O_1321,N_8893,N_9842);
nor UO_1322 (O_1322,N_5957,N_5805);
nand UO_1323 (O_1323,N_9684,N_5629);
nand UO_1324 (O_1324,N_6702,N_9826);
or UO_1325 (O_1325,N_7710,N_8991);
nand UO_1326 (O_1326,N_7828,N_8383);
nand UO_1327 (O_1327,N_9220,N_5495);
or UO_1328 (O_1328,N_6403,N_7958);
nor UO_1329 (O_1329,N_5645,N_8540);
nor UO_1330 (O_1330,N_5470,N_8358);
or UO_1331 (O_1331,N_6531,N_6732);
and UO_1332 (O_1332,N_9175,N_9784);
and UO_1333 (O_1333,N_5561,N_7114);
nand UO_1334 (O_1334,N_9214,N_8777);
or UO_1335 (O_1335,N_5299,N_5678);
nor UO_1336 (O_1336,N_8882,N_8310);
nor UO_1337 (O_1337,N_6577,N_8986);
and UO_1338 (O_1338,N_9975,N_9363);
or UO_1339 (O_1339,N_9263,N_9284);
nor UO_1340 (O_1340,N_8607,N_9086);
or UO_1341 (O_1341,N_9229,N_8237);
and UO_1342 (O_1342,N_6657,N_9929);
and UO_1343 (O_1343,N_5597,N_8621);
and UO_1344 (O_1344,N_8257,N_7385);
nand UO_1345 (O_1345,N_8989,N_6537);
xnor UO_1346 (O_1346,N_5226,N_7952);
nor UO_1347 (O_1347,N_6128,N_5859);
or UO_1348 (O_1348,N_8476,N_9855);
or UO_1349 (O_1349,N_5406,N_8213);
and UO_1350 (O_1350,N_6855,N_5840);
and UO_1351 (O_1351,N_5329,N_6803);
or UO_1352 (O_1352,N_5922,N_7248);
or UO_1353 (O_1353,N_6409,N_9596);
and UO_1354 (O_1354,N_9677,N_8362);
or UO_1355 (O_1355,N_7282,N_6586);
nand UO_1356 (O_1356,N_8938,N_7341);
nor UO_1357 (O_1357,N_9526,N_5595);
xor UO_1358 (O_1358,N_5570,N_7829);
or UO_1359 (O_1359,N_9103,N_8088);
nand UO_1360 (O_1360,N_8815,N_8998);
nand UO_1361 (O_1361,N_5940,N_9795);
nor UO_1362 (O_1362,N_5181,N_6474);
nand UO_1363 (O_1363,N_8151,N_7853);
nand UO_1364 (O_1364,N_7780,N_8364);
nor UO_1365 (O_1365,N_9291,N_5691);
and UO_1366 (O_1366,N_5115,N_8713);
nor UO_1367 (O_1367,N_5862,N_8601);
nand UO_1368 (O_1368,N_7778,N_5910);
xnor UO_1369 (O_1369,N_7053,N_6846);
nand UO_1370 (O_1370,N_7905,N_9525);
nor UO_1371 (O_1371,N_7581,N_9878);
or UO_1372 (O_1372,N_6945,N_9469);
nand UO_1373 (O_1373,N_9550,N_7037);
or UO_1374 (O_1374,N_5439,N_9971);
nand UO_1375 (O_1375,N_5914,N_9537);
nor UO_1376 (O_1376,N_6541,N_9822);
nand UO_1377 (O_1377,N_6960,N_9063);
or UO_1378 (O_1378,N_9579,N_7807);
xor UO_1379 (O_1379,N_6304,N_5539);
nand UO_1380 (O_1380,N_9418,N_9095);
nor UO_1381 (O_1381,N_9621,N_7679);
and UO_1382 (O_1382,N_6174,N_9176);
nor UO_1383 (O_1383,N_5604,N_7942);
nand UO_1384 (O_1384,N_7437,N_6653);
nor UO_1385 (O_1385,N_7192,N_8898);
and UO_1386 (O_1386,N_5829,N_8603);
and UO_1387 (O_1387,N_6274,N_8416);
nor UO_1388 (O_1388,N_7129,N_6119);
and UO_1389 (O_1389,N_7893,N_7503);
and UO_1390 (O_1390,N_8478,N_6314);
nor UO_1391 (O_1391,N_5207,N_6354);
nand UO_1392 (O_1392,N_7845,N_5876);
nand UO_1393 (O_1393,N_5907,N_5675);
nand UO_1394 (O_1394,N_7445,N_6750);
nor UO_1395 (O_1395,N_5935,N_8671);
nor UO_1396 (O_1396,N_9523,N_6230);
or UO_1397 (O_1397,N_5898,N_7569);
nand UO_1398 (O_1398,N_9226,N_6052);
nor UO_1399 (O_1399,N_5133,N_6473);
nor UO_1400 (O_1400,N_7246,N_8052);
or UO_1401 (O_1401,N_7591,N_6115);
or UO_1402 (O_1402,N_7021,N_7085);
and UO_1403 (O_1403,N_9829,N_5867);
or UO_1404 (O_1404,N_5527,N_7908);
or UO_1405 (O_1405,N_5123,N_7724);
nor UO_1406 (O_1406,N_9003,N_9186);
and UO_1407 (O_1407,N_7939,N_7386);
nand UO_1408 (O_1408,N_8896,N_5381);
and UO_1409 (O_1409,N_9475,N_6807);
nand UO_1410 (O_1410,N_8190,N_6482);
or UO_1411 (O_1411,N_9587,N_6763);
and UO_1412 (O_1412,N_5571,N_6027);
nor UO_1413 (O_1413,N_6021,N_6587);
nand UO_1414 (O_1414,N_7896,N_9866);
and UO_1415 (O_1415,N_8078,N_8177);
nor UO_1416 (O_1416,N_5809,N_7393);
nor UO_1417 (O_1417,N_5369,N_5099);
and UO_1418 (O_1418,N_6890,N_7528);
or UO_1419 (O_1419,N_9390,N_6148);
nor UO_1420 (O_1420,N_7482,N_9385);
xor UO_1421 (O_1421,N_6644,N_6739);
or UO_1422 (O_1422,N_6381,N_8122);
nand UO_1423 (O_1423,N_8178,N_6748);
and UO_1424 (O_1424,N_5269,N_8541);
and UO_1425 (O_1425,N_9650,N_9306);
xnor UO_1426 (O_1426,N_9888,N_7054);
and UO_1427 (O_1427,N_8765,N_5310);
nand UO_1428 (O_1428,N_6670,N_9341);
nand UO_1429 (O_1429,N_5803,N_9318);
or UO_1430 (O_1430,N_5626,N_5683);
nand UO_1431 (O_1431,N_8505,N_9943);
or UO_1432 (O_1432,N_6160,N_6561);
nand UO_1433 (O_1433,N_8856,N_5354);
and UO_1434 (O_1434,N_8322,N_9260);
or UO_1435 (O_1435,N_9373,N_8628);
and UO_1436 (O_1436,N_6529,N_8032);
nand UO_1437 (O_1437,N_8958,N_8482);
nand UO_1438 (O_1438,N_8862,N_5657);
and UO_1439 (O_1439,N_6790,N_5615);
xor UO_1440 (O_1440,N_6238,N_6543);
or UO_1441 (O_1441,N_9774,N_9114);
nor UO_1442 (O_1442,N_6701,N_7137);
or UO_1443 (O_1443,N_7416,N_7832);
and UO_1444 (O_1444,N_7395,N_8863);
xnor UO_1445 (O_1445,N_9953,N_6451);
nor UO_1446 (O_1446,N_7662,N_5171);
nand UO_1447 (O_1447,N_6614,N_7322);
nand UO_1448 (O_1448,N_7920,N_9735);
and UO_1449 (O_1449,N_7877,N_6047);
and UO_1450 (O_1450,N_5282,N_5943);
or UO_1451 (O_1451,N_9394,N_5894);
nand UO_1452 (O_1452,N_7048,N_8620);
or UO_1453 (O_1453,N_8351,N_7375);
nor UO_1454 (O_1454,N_5525,N_6851);
nor UO_1455 (O_1455,N_8956,N_6377);
xor UO_1456 (O_1456,N_5338,N_8325);
nand UO_1457 (O_1457,N_7922,N_9361);
and UO_1458 (O_1458,N_9338,N_9084);
nor UO_1459 (O_1459,N_6302,N_6254);
and UO_1460 (O_1460,N_8984,N_7519);
nor UO_1461 (O_1461,N_8630,N_6494);
or UO_1462 (O_1462,N_9061,N_8855);
nand UO_1463 (O_1463,N_9199,N_9461);
nor UO_1464 (O_1464,N_5573,N_7124);
nor UO_1465 (O_1465,N_6832,N_6389);
and UO_1466 (O_1466,N_9578,N_6007);
nor UO_1467 (O_1467,N_9192,N_9797);
nand UO_1468 (O_1468,N_9566,N_9158);
nor UO_1469 (O_1469,N_7376,N_5982);
nand UO_1470 (O_1470,N_7401,N_9689);
nand UO_1471 (O_1471,N_8473,N_8062);
nor UO_1472 (O_1472,N_5587,N_8428);
or UO_1473 (O_1473,N_5842,N_9066);
or UO_1474 (O_1474,N_9313,N_5340);
and UO_1475 (O_1475,N_6581,N_9769);
nor UO_1476 (O_1476,N_7936,N_6767);
or UO_1477 (O_1477,N_7208,N_6745);
and UO_1478 (O_1478,N_9264,N_7402);
nor UO_1479 (O_1479,N_9008,N_9463);
and UO_1480 (O_1480,N_8425,N_8431);
or UO_1481 (O_1481,N_9195,N_9001);
nand UO_1482 (O_1482,N_6202,N_6003);
or UO_1483 (O_1483,N_6738,N_9631);
and UO_1484 (O_1484,N_9251,N_8927);
nor UO_1485 (O_1485,N_9227,N_5494);
xnor UO_1486 (O_1486,N_9028,N_9399);
xor UO_1487 (O_1487,N_8949,N_6268);
nor UO_1488 (O_1488,N_6263,N_9683);
and UO_1489 (O_1489,N_5501,N_6156);
and UO_1490 (O_1490,N_6211,N_5106);
nand UO_1491 (O_1491,N_6092,N_5522);
or UO_1492 (O_1492,N_6203,N_7543);
nor UO_1493 (O_1493,N_5301,N_9531);
nor UO_1494 (O_1494,N_7058,N_7165);
nand UO_1495 (O_1495,N_8047,N_6691);
nand UO_1496 (O_1496,N_9102,N_8802);
or UO_1497 (O_1497,N_9019,N_9703);
nor UO_1498 (O_1498,N_7003,N_8008);
or UO_1499 (O_1499,N_9491,N_5554);
endmodule