module basic_3000_30000_3500_6_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_1439,In_1797);
nor U1 (N_1,In_1718,In_2759);
or U2 (N_2,In_2967,In_1498);
xor U3 (N_3,In_499,In_1568);
nand U4 (N_4,In_2447,In_2979);
xnor U5 (N_5,In_393,In_2550);
xor U6 (N_6,In_2687,In_454);
and U7 (N_7,In_509,In_2364);
nand U8 (N_8,In_561,In_457);
or U9 (N_9,In_2171,In_1944);
nor U10 (N_10,In_2668,In_217);
xor U11 (N_11,In_2213,In_140);
xnor U12 (N_12,In_672,In_2869);
nor U13 (N_13,In_643,In_221);
xnor U14 (N_14,In_1099,In_2441);
and U15 (N_15,In_2525,In_2038);
nor U16 (N_16,In_648,In_2341);
nand U17 (N_17,In_621,In_712);
or U18 (N_18,In_1359,In_1759);
and U19 (N_19,In_1722,In_742);
nand U20 (N_20,In_163,In_965);
xor U21 (N_21,In_622,In_735);
or U22 (N_22,In_2340,In_529);
nand U23 (N_23,In_663,In_1689);
nand U24 (N_24,In_2893,In_1122);
xnor U25 (N_25,In_629,In_2480);
or U26 (N_26,In_932,In_1915);
and U27 (N_27,In_2512,In_1199);
nor U28 (N_28,In_2702,In_2253);
and U29 (N_29,In_2453,In_1593);
nand U30 (N_30,In_530,In_2673);
nand U31 (N_31,In_189,In_1173);
nor U32 (N_32,In_1336,In_2634);
nand U33 (N_33,In_758,In_146);
or U34 (N_34,In_2238,In_1539);
nand U35 (N_35,In_689,In_1303);
xnor U36 (N_36,In_2137,In_2663);
or U37 (N_37,In_946,In_394);
nor U38 (N_38,In_2800,In_2083);
xnor U39 (N_39,In_1928,In_1633);
and U40 (N_40,In_1367,In_485);
nor U41 (N_41,In_1550,In_805);
xnor U42 (N_42,In_2763,In_2022);
nand U43 (N_43,In_653,In_1136);
xnor U44 (N_44,In_327,In_2944);
nand U45 (N_45,In_102,In_1662);
nor U46 (N_46,In_2335,In_626);
xor U47 (N_47,In_2460,In_1117);
or U48 (N_48,In_2089,In_1644);
and U49 (N_49,In_1046,In_746);
nor U50 (N_50,In_972,In_1030);
and U51 (N_51,In_1396,In_2991);
nor U52 (N_52,In_1618,In_1570);
nor U53 (N_53,In_2294,In_2913);
xor U54 (N_54,In_97,In_1461);
xnor U55 (N_55,In_1636,In_577);
or U56 (N_56,In_249,In_649);
and U57 (N_57,In_1112,In_83);
nand U58 (N_58,In_2692,In_1007);
or U59 (N_59,In_2555,In_1160);
nand U60 (N_60,In_1673,In_696);
xnor U61 (N_61,In_537,In_1666);
xor U62 (N_62,In_585,In_1577);
nand U63 (N_63,In_2515,In_107);
nand U64 (N_64,In_63,In_1992);
nand U65 (N_65,In_761,In_2570);
nor U66 (N_66,In_2844,In_1398);
or U67 (N_67,In_595,In_1419);
nor U68 (N_68,In_2006,In_2632);
or U69 (N_69,In_2675,In_2355);
and U70 (N_70,In_2354,In_1067);
and U71 (N_71,In_2464,In_2533);
xnor U72 (N_72,In_195,In_2313);
and U73 (N_73,In_1588,In_474);
nor U74 (N_74,In_2943,In_2385);
and U75 (N_75,In_2191,In_166);
xor U76 (N_76,In_329,In_1225);
xnor U77 (N_77,In_1228,In_1925);
xnor U78 (N_78,In_2193,In_1346);
or U79 (N_79,In_274,In_695);
nor U80 (N_80,In_1860,In_2620);
and U81 (N_81,In_1532,In_2109);
xnor U82 (N_82,In_1516,In_1485);
xor U83 (N_83,In_278,In_1170);
nor U84 (N_84,In_920,In_2283);
and U85 (N_85,In_747,In_2314);
nand U86 (N_86,In_243,In_1014);
and U87 (N_87,In_1563,In_541);
nand U88 (N_88,In_368,In_2851);
and U89 (N_89,In_1765,In_2579);
nor U90 (N_90,In_2788,In_460);
or U91 (N_91,In_2141,In_2931);
nand U92 (N_92,In_2823,In_2155);
xor U93 (N_93,In_2474,In_871);
and U94 (N_94,In_1247,In_1653);
or U95 (N_95,In_2771,In_2228);
xor U96 (N_96,In_2431,In_2619);
xor U97 (N_97,In_1163,In_567);
nand U98 (N_98,In_2119,In_2523);
xor U99 (N_99,In_1569,In_1056);
and U100 (N_100,In_2066,In_478);
xor U101 (N_101,In_416,In_1839);
and U102 (N_102,In_2451,In_2592);
and U103 (N_103,In_1310,In_358);
nor U104 (N_104,In_1754,In_366);
or U105 (N_105,In_2754,In_706);
and U106 (N_106,In_1592,In_950);
nand U107 (N_107,In_1863,In_253);
or U108 (N_108,In_2279,In_2093);
xor U109 (N_109,In_344,In_1276);
nor U110 (N_110,In_2998,In_2172);
and U111 (N_111,In_2027,In_1183);
nand U112 (N_112,In_2573,In_1930);
nor U113 (N_113,In_1409,In_1105);
and U114 (N_114,In_898,In_2516);
or U115 (N_115,In_2130,In_988);
nor U116 (N_116,In_936,In_1637);
nand U117 (N_117,In_1148,In_318);
nor U118 (N_118,In_2802,In_2725);
nor U119 (N_119,In_1833,In_439);
or U120 (N_120,In_1541,In_799);
or U121 (N_121,In_106,In_1251);
and U122 (N_122,In_1273,In_1741);
xor U123 (N_123,In_1190,In_808);
xor U124 (N_124,In_100,In_429);
or U125 (N_125,In_1040,In_2617);
nor U126 (N_126,In_2973,In_2747);
or U127 (N_127,In_232,In_1203);
xnor U128 (N_128,In_828,In_598);
and U129 (N_129,In_999,In_1055);
and U130 (N_130,In_1172,In_208);
nor U131 (N_131,In_612,In_1442);
or U132 (N_132,In_2816,In_2121);
xnor U133 (N_133,In_1238,In_1942);
and U134 (N_134,In_558,In_2189);
or U135 (N_135,In_875,In_2566);
xor U136 (N_136,In_66,In_152);
nor U137 (N_137,In_795,In_673);
nand U138 (N_138,In_1536,In_2491);
or U139 (N_139,In_2285,In_555);
nand U140 (N_140,In_2930,In_1265);
nor U141 (N_141,In_1631,In_2960);
and U142 (N_142,In_2380,In_1427);
nor U143 (N_143,In_1425,In_284);
xnor U144 (N_144,In_780,In_1213);
xnor U145 (N_145,In_519,In_2072);
nand U146 (N_146,In_28,In_513);
xor U147 (N_147,In_188,In_588);
and U148 (N_148,In_1590,In_1406);
or U149 (N_149,In_2704,In_667);
and U150 (N_150,In_1240,In_1282);
and U151 (N_151,In_313,In_2607);
and U152 (N_152,In_660,In_929);
nor U153 (N_153,In_296,In_526);
nand U154 (N_154,In_586,In_989);
or U155 (N_155,In_2300,In_1481);
xor U156 (N_156,In_760,In_2809);
nand U157 (N_157,In_2418,In_1413);
nor U158 (N_158,In_2030,In_1432);
xnor U159 (N_159,In_2440,In_641);
nand U160 (N_160,In_2925,In_2985);
and U161 (N_161,In_2321,In_2654);
or U162 (N_162,In_2105,In_2195);
nand U163 (N_163,In_1076,In_908);
and U164 (N_164,In_3,In_2848);
or U165 (N_165,In_1298,In_2409);
or U166 (N_166,In_443,In_1808);
and U167 (N_167,In_1855,In_2002);
or U168 (N_168,In_1377,In_82);
nand U169 (N_169,In_973,In_1189);
and U170 (N_170,In_1913,In_2400);
xor U171 (N_171,In_105,In_763);
or U172 (N_172,In_456,In_1374);
nand U173 (N_173,In_2551,In_183);
xnor U174 (N_174,In_79,In_831);
nor U175 (N_175,In_882,In_919);
nor U176 (N_176,In_2974,In_1278);
and U177 (N_177,In_2527,In_173);
or U178 (N_178,In_914,In_1756);
nor U179 (N_179,In_7,In_560);
nor U180 (N_180,In_1482,In_844);
nand U181 (N_181,In_1285,In_126);
and U182 (N_182,In_2173,In_593);
xnor U183 (N_183,In_2317,In_2686);
nand U184 (N_184,In_354,In_2589);
nand U185 (N_185,In_231,In_2237);
nand U186 (N_186,In_1943,In_353);
nand U187 (N_187,In_227,In_450);
nor U188 (N_188,In_1953,In_1380);
xor U189 (N_189,In_1916,In_2520);
nor U190 (N_190,In_2125,In_2830);
and U191 (N_191,In_1341,In_1693);
nand U192 (N_192,In_983,In_1993);
xnor U193 (N_193,In_1640,In_2707);
nor U194 (N_194,In_809,In_2582);
or U195 (N_195,In_2475,In_1312);
nand U196 (N_196,In_2631,In_1392);
xnor U197 (N_197,In_2138,In_553);
nor U198 (N_198,In_1975,In_91);
nand U199 (N_199,In_120,In_2009);
xnor U200 (N_200,In_2733,In_2234);
or U201 (N_201,In_2588,In_1522);
xor U202 (N_202,In_1039,In_178);
and U203 (N_203,In_1186,In_687);
nand U204 (N_204,In_2067,In_1558);
xnor U205 (N_205,In_2184,In_2047);
or U206 (N_206,In_2787,In_1772);
nor U207 (N_207,In_1082,In_782);
nor U208 (N_208,In_2946,In_938);
nor U209 (N_209,In_1876,In_963);
nand U210 (N_210,In_2458,In_1834);
xor U211 (N_211,In_128,In_1331);
xor U212 (N_212,In_4,In_1260);
or U213 (N_213,In_2495,In_1467);
nand U214 (N_214,In_1580,In_1033);
nor U215 (N_215,In_321,In_1776);
or U216 (N_216,In_1524,In_2194);
xnor U217 (N_217,In_2102,In_2466);
and U218 (N_218,In_86,In_741);
xor U219 (N_219,In_240,In_571);
and U220 (N_220,In_1243,In_315);
nand U221 (N_221,In_1687,In_1429);
nor U222 (N_222,In_2059,In_1668);
and U223 (N_223,In_2628,In_1921);
xnor U224 (N_224,In_2674,In_76);
or U225 (N_225,In_901,In_543);
or U226 (N_226,In_1037,In_1441);
and U227 (N_227,In_1527,In_1678);
or U228 (N_228,In_2423,In_915);
xnor U229 (N_229,In_258,In_1297);
and U230 (N_230,In_1326,In_897);
and U231 (N_231,In_469,In_1496);
xor U232 (N_232,In_1700,In_2572);
or U233 (N_233,In_2199,In_2270);
nor U234 (N_234,In_2698,In_468);
nand U235 (N_235,In_2945,In_1459);
xnor U236 (N_236,In_2357,In_1691);
nand U237 (N_237,In_2996,In_1702);
xor U238 (N_238,In_975,In_1500);
or U239 (N_239,In_2282,In_1624);
and U240 (N_240,In_2815,In_2114);
and U241 (N_241,In_866,In_1089);
nor U242 (N_242,In_566,In_2150);
nor U243 (N_243,In_2084,In_820);
nand U244 (N_244,In_1462,In_1463);
xnor U245 (N_245,In_873,In_1308);
or U246 (N_246,In_281,In_135);
nand U247 (N_247,In_878,In_1224);
nor U248 (N_248,In_359,In_2837);
or U249 (N_249,In_1403,In_62);
xnor U250 (N_250,In_2835,In_838);
and U251 (N_251,In_1683,In_88);
nand U252 (N_252,In_273,In_1692);
or U253 (N_253,In_2372,In_1023);
nor U254 (N_254,In_1074,In_930);
nand U255 (N_255,In_2874,In_1383);
or U256 (N_256,In_13,In_2583);
and U257 (N_257,In_2894,In_1779);
nand U258 (N_258,In_2404,In_969);
nor U259 (N_259,In_471,In_874);
nand U260 (N_260,In_582,In_430);
or U261 (N_261,In_190,In_2118);
or U262 (N_262,In_2750,In_1946);
nor U263 (N_263,In_2478,In_320);
xnor U264 (N_264,In_1342,In_705);
or U265 (N_265,In_2263,In_2261);
and U266 (N_266,In_1529,In_2057);
xor U267 (N_267,In_1535,In_1284);
and U268 (N_268,In_2266,In_1865);
nor U269 (N_269,In_1845,In_2405);
and U270 (N_270,In_9,In_1514);
nor U271 (N_271,In_204,In_497);
xnor U272 (N_272,In_2697,In_1017);
nor U273 (N_273,In_2088,In_1674);
nand U274 (N_274,In_2770,In_1645);
nand U275 (N_275,In_2638,In_2268);
or U276 (N_276,In_36,In_350);
nor U277 (N_277,In_1837,In_1824);
or U278 (N_278,In_1068,In_1766);
nor U279 (N_279,In_2500,In_1329);
and U280 (N_280,In_1620,In_532);
xor U281 (N_281,In_2581,In_418);
xor U282 (N_282,In_1339,In_2483);
xor U283 (N_283,In_1245,In_1307);
or U284 (N_284,In_2262,In_2965);
xnor U285 (N_285,In_2627,In_2711);
nand U286 (N_286,In_444,In_2370);
nand U287 (N_287,In_821,In_56);
xnor U288 (N_288,In_1399,In_565);
nand U289 (N_289,In_2056,In_2330);
or U290 (N_290,In_2861,In_382);
or U291 (N_291,In_2855,In_1426);
xnor U292 (N_292,In_2021,In_299);
or U293 (N_293,In_583,In_2929);
and U294 (N_294,In_2752,In_2232);
and U295 (N_295,In_2514,In_1446);
xor U296 (N_296,In_2188,In_2406);
nand U297 (N_297,In_576,In_293);
or U298 (N_298,In_786,In_853);
and U299 (N_299,In_515,In_1609);
xor U300 (N_300,In_2645,In_528);
xnor U301 (N_301,In_1574,In_12);
xor U302 (N_302,In_1156,In_2274);
xor U303 (N_303,In_2537,In_2806);
nor U304 (N_304,In_1748,In_1242);
xnor U305 (N_305,In_1275,In_1319);
xor U306 (N_306,In_951,In_592);
xnor U307 (N_307,In_1706,In_647);
nand U308 (N_308,In_1192,In_548);
or U309 (N_309,In_2124,In_710);
nor U310 (N_310,In_72,In_1422);
nor U311 (N_311,In_2329,In_522);
xnor U312 (N_312,In_2110,In_779);
and U313 (N_313,In_2653,In_804);
and U314 (N_314,In_248,In_1787);
nor U315 (N_315,In_2726,In_2046);
xnor U316 (N_316,In_1761,In_2896);
nor U317 (N_317,In_1447,In_993);
xnor U318 (N_318,In_1100,In_230);
or U319 (N_319,In_1635,In_493);
or U320 (N_320,In_1233,In_2981);
nor U321 (N_321,In_1801,In_916);
nor U322 (N_322,In_1230,In_2033);
xnor U323 (N_323,In_54,In_2966);
nor U324 (N_324,In_1982,In_1841);
or U325 (N_325,In_2769,In_2135);
xor U326 (N_326,In_2304,In_1826);
nor U327 (N_327,In_1113,In_171);
nand U328 (N_328,In_2510,In_373);
xnor U329 (N_329,In_408,In_1384);
nor U330 (N_330,In_899,In_1083);
nor U331 (N_331,In_542,In_235);
or U332 (N_332,In_856,In_399);
nor U333 (N_333,In_2459,In_1850);
and U334 (N_334,In_1875,In_1817);
xnor U335 (N_335,In_1200,In_1544);
nand U336 (N_336,In_1013,In_1395);
nand U337 (N_337,In_1231,In_255);
nor U338 (N_338,In_1026,In_2644);
nand U339 (N_339,In_2269,In_1065);
nor U340 (N_340,In_2684,In_650);
nor U341 (N_341,In_841,In_1862);
nand U342 (N_342,In_196,In_2338);
nor U343 (N_343,In_2328,In_992);
and U344 (N_344,In_2739,In_2741);
xnor U345 (N_345,In_1474,In_2486);
xor U346 (N_346,In_1153,In_2361);
nor U347 (N_347,In_214,In_2097);
nand U348 (N_348,In_2876,In_772);
xor U349 (N_349,In_2158,In_2889);
xnor U350 (N_350,In_2443,In_340);
or U351 (N_351,In_2103,In_1878);
nand U352 (N_352,In_1651,In_467);
nand U353 (N_353,In_1932,In_45);
or U354 (N_354,In_1729,In_2362);
nor U355 (N_355,In_1965,In_1445);
nor U356 (N_356,In_1132,In_1330);
xnor U357 (N_357,In_187,In_209);
xor U358 (N_358,In_2461,In_2014);
or U359 (N_359,In_1911,In_788);
xnor U360 (N_360,In_1047,In_1137);
and U361 (N_361,In_848,In_974);
or U362 (N_362,In_968,In_697);
or U363 (N_363,In_682,In_1545);
nand U364 (N_364,In_19,In_27);
and U365 (N_365,In_378,In_2153);
nand U366 (N_366,In_2374,In_2899);
or U367 (N_367,In_2,In_2319);
and U368 (N_368,In_1941,In_2111);
nand U369 (N_369,In_1891,In_2174);
xnor U370 (N_370,In_2571,In_316);
nor U371 (N_371,In_291,In_1052);
nand U372 (N_372,In_2968,In_60);
and U373 (N_373,In_2933,In_2614);
nor U374 (N_374,In_2530,In_1881);
xor U375 (N_375,In_698,In_1239);
nor U376 (N_376,In_1910,In_889);
nor U377 (N_377,In_1456,In_2558);
and U378 (N_378,In_219,In_1643);
nor U379 (N_379,In_2467,In_2856);
nand U380 (N_380,In_757,In_880);
nor U381 (N_381,In_1387,In_1733);
and U382 (N_382,In_1513,In_2753);
or U383 (N_383,In_265,In_1106);
nor U384 (N_384,In_1281,In_192);
or U385 (N_385,In_958,In_10);
and U386 (N_386,In_2498,In_421);
nor U387 (N_387,In_1300,In_2226);
xnor U388 (N_388,In_159,In_266);
nand U389 (N_389,In_417,In_2576);
and U390 (N_390,In_2358,In_2011);
or U391 (N_391,In_1742,In_169);
and U392 (N_392,In_618,In_716);
and U393 (N_393,In_1174,In_1011);
nand U394 (N_394,In_2288,In_412);
and U395 (N_395,In_1489,In_5);
nor U396 (N_396,In_2389,In_1652);
nand U397 (N_397,In_1378,In_2049);
nor U398 (N_398,In_2618,In_2951);
nand U399 (N_399,In_1010,In_1370);
nand U400 (N_400,In_818,In_1904);
or U401 (N_401,In_2356,In_2434);
nand U402 (N_402,In_2200,In_1110);
nand U403 (N_403,In_1505,In_317);
or U404 (N_404,In_386,In_372);
or U405 (N_405,In_381,In_489);
and U406 (N_406,In_367,In_2780);
xor U407 (N_407,In_1115,In_1139);
and U408 (N_408,In_1453,In_546);
nand U409 (N_409,In_686,In_16);
nor U410 (N_410,In_807,In_2688);
xnor U411 (N_411,In_55,In_700);
nor U412 (N_412,In_1149,In_2168);
nor U413 (N_413,In_851,In_2323);
nand U414 (N_414,In_2120,In_2371);
nor U415 (N_415,In_1080,In_2792);
nor U416 (N_416,In_237,In_338);
xnor U417 (N_417,In_1193,In_978);
or U418 (N_418,In_994,In_1546);
nor U419 (N_419,In_402,In_2902);
and U420 (N_420,In_1730,In_1185);
xnor U421 (N_421,In_2136,In_1);
xor U422 (N_422,In_1428,In_2594);
xor U423 (N_423,In_2610,In_314);
nor U424 (N_424,In_1716,In_2701);
nor U425 (N_425,In_1220,In_632);
nand U426 (N_426,In_1502,In_1882);
and U427 (N_427,In_1760,In_1176);
nand U428 (N_428,In_2696,In_596);
nand U429 (N_429,In_642,In_285);
and U430 (N_430,In_1709,In_199);
xor U431 (N_431,In_2148,In_148);
nor U432 (N_432,In_466,In_2834);
or U433 (N_433,In_22,In_986);
nor U434 (N_434,In_2322,In_945);
or U435 (N_435,In_572,In_2852);
nor U436 (N_436,In_1057,In_644);
nand U437 (N_437,In_2430,In_440);
nand U438 (N_438,In_2764,In_864);
nand U439 (N_439,In_43,In_1263);
or U440 (N_440,In_603,In_1101);
xor U441 (N_441,In_1092,In_1090);
nor U442 (N_442,In_110,In_2079);
and U443 (N_443,In_1968,In_1988);
nor U444 (N_444,In_2100,In_960);
and U445 (N_445,In_310,In_1901);
nand U446 (N_446,In_1671,In_2783);
or U447 (N_447,In_2801,In_1713);
nor U448 (N_448,In_2567,In_1034);
nor U449 (N_449,In_477,In_42);
nor U450 (N_450,In_677,In_1663);
xnor U451 (N_451,In_2660,In_1704);
or U452 (N_452,In_370,In_2470);
and U453 (N_453,In_1484,In_1438);
nor U454 (N_454,In_554,In_616);
or U455 (N_455,In_1191,In_1884);
and U456 (N_456,In_2363,In_691);
and U457 (N_457,In_405,In_1368);
xor U458 (N_458,In_1471,In_1218);
xor U459 (N_459,In_2235,In_2108);
nand U460 (N_460,In_1789,In_815);
nand U461 (N_461,In_2846,In_1021);
and U462 (N_462,In_1261,In_1867);
or U463 (N_463,In_2730,In_1825);
nor U464 (N_464,In_2432,In_2161);
nor U465 (N_465,In_2126,In_465);
or U466 (N_466,In_2828,In_1000);
and U467 (N_467,In_723,In_1274);
nor U468 (N_468,In_2553,In_2394);
nand U469 (N_469,In_2517,In_1045);
and U470 (N_470,In_1880,In_2518);
nand U471 (N_471,In_1216,In_1957);
and U472 (N_472,In_85,In_2252);
or U473 (N_473,In_1929,In_1361);
or U474 (N_474,In_2101,In_1466);
xnor U475 (N_475,In_2035,In_2647);
nand U476 (N_476,In_910,In_819);
or U477 (N_477,In_2069,In_2403);
and U478 (N_478,In_1736,In_2648);
or U479 (N_479,In_922,In_1177);
and U480 (N_480,In_1042,In_1894);
xnor U481 (N_481,In_2877,In_2908);
xnor U482 (N_482,In_200,In_2821);
xor U483 (N_483,In_2842,In_180);
nor U484 (N_484,In_693,In_89);
nor U485 (N_485,In_2482,In_711);
and U486 (N_486,In_638,In_1515);
nand U487 (N_487,In_1480,In_980);
or U488 (N_488,In_2492,In_2871);
and U489 (N_489,In_491,In_1695);
and U490 (N_490,In_2712,In_568);
nor U491 (N_491,In_1940,In_2600);
nand U492 (N_492,In_2909,In_486);
xor U493 (N_493,In_441,In_1254);
and U494 (N_494,In_2457,In_2920);
xor U495 (N_495,In_1168,In_2207);
nor U496 (N_496,In_481,In_2337);
xnor U497 (N_497,In_656,In_2840);
and U498 (N_498,In_2422,In_604);
xnor U499 (N_499,In_933,In_2302);
and U500 (N_500,In_2705,In_2157);
nor U501 (N_501,In_2490,In_2845);
and U502 (N_502,In_438,In_2671);
and U503 (N_503,In_1071,In_1927);
nor U504 (N_504,In_817,In_2822);
nand U505 (N_505,In_751,In_1317);
nand U506 (N_506,In_1997,In_2343);
and U507 (N_507,In_1443,In_275);
or U508 (N_508,In_2664,In_1158);
nand U509 (N_509,In_1133,In_488);
xnor U510 (N_510,In_2165,In_1495);
nor U511 (N_511,In_2078,In_2849);
xor U512 (N_512,In_2230,In_1559);
nand U513 (N_513,In_847,In_1194);
xor U514 (N_514,In_234,In_1141);
nor U515 (N_515,In_573,In_2142);
or U516 (N_516,In_2156,In_1657);
and U517 (N_517,In_2015,In_1134);
and U518 (N_518,In_722,In_2924);
nor U519 (N_519,In_2824,In_2164);
or U520 (N_520,In_215,In_830);
xnor U521 (N_521,In_2324,In_279);
xnor U522 (N_522,In_1490,In_1188);
xor U523 (N_523,In_2504,In_1737);
xnor U524 (N_524,In_2298,In_510);
nor U525 (N_525,In_521,In_401);
nor U526 (N_526,In_2182,In_610);
nand U527 (N_527,In_2106,In_617);
xor U528 (N_528,In_426,In_2229);
nor U529 (N_529,In_64,In_1126);
and U530 (N_530,In_1041,In_1152);
xnor U531 (N_531,In_1764,In_2216);
and U532 (N_532,In_2580,In_1267);
nand U533 (N_533,In_2336,In_2254);
nor U534 (N_534,In_348,In_1816);
and U535 (N_535,In_2503,In_1084);
nor U536 (N_536,In_991,In_1154);
xnor U537 (N_537,In_2352,In_2604);
nand U538 (N_538,In_692,In_1049);
nand U539 (N_539,In_2782,In_1807);
or U540 (N_540,In_1364,In_2519);
and U541 (N_541,In_2315,In_1348);
nor U542 (N_542,In_1596,In_1108);
nand U543 (N_543,In_1209,In_896);
nor U544 (N_544,In_2536,In_1397);
nand U545 (N_545,In_2393,In_2190);
and U546 (N_546,In_1743,In_1411);
nand U547 (N_547,In_1005,In_2587);
xor U548 (N_548,In_1264,In_458);
and U549 (N_549,In_2387,In_2095);
xor U550 (N_550,In_2767,In_1530);
xor U551 (N_551,In_494,In_1972);
xor U552 (N_552,In_2599,In_32);
and U553 (N_553,In_361,In_21);
nor U554 (N_554,In_400,In_1622);
nor U555 (N_555,In_211,In_1151);
or U556 (N_556,In_2679,In_2411);
or U557 (N_557,In_2133,In_1871);
and U558 (N_558,In_301,In_2825);
or U559 (N_559,In_1400,In_1433);
nand U560 (N_560,In_392,In_2887);
and U561 (N_561,In_1362,In_2112);
and U562 (N_562,In_1688,In_784);
nand U563 (N_563,In_2421,In_319);
and U564 (N_564,In_886,In_2528);
nand U565 (N_565,In_2736,In_2318);
nor U566 (N_566,In_1236,In_2773);
xor U567 (N_567,In_14,In_1950);
or U568 (N_568,In_1805,In_2728);
or U569 (N_569,In_1520,In_229);
and U570 (N_570,In_1585,In_134);
nand U571 (N_571,In_590,In_2071);
nand U572 (N_572,In_2048,In_1914);
or U573 (N_573,In_2416,In_646);
or U574 (N_574,In_551,In_2596);
or U575 (N_575,In_1939,In_1676);
nor U576 (N_576,In_2905,In_404);
nand U577 (N_577,In_225,In_1896);
nand U578 (N_578,In_924,In_112);
xnor U579 (N_579,In_2473,In_2000);
and U580 (N_580,In_563,In_155);
or U581 (N_581,In_286,In_2542);
or U582 (N_582,In_2774,In_2429);
xnor U583 (N_583,In_58,In_132);
and U584 (N_584,In_2751,In_245);
or U585 (N_585,In_1198,In_324);
nor U586 (N_586,In_942,In_2376);
xor U587 (N_587,In_1135,In_51);
xor U588 (N_588,In_1829,In_2737);
xor U589 (N_589,In_445,In_47);
and U590 (N_590,In_887,In_351);
or U591 (N_591,In_552,In_1542);
nand U592 (N_592,In_52,In_2613);
nor U593 (N_593,In_507,In_768);
and U594 (N_594,In_1523,In_2170);
or U595 (N_595,In_2936,In_2176);
nor U596 (N_596,In_1828,In_2786);
nor U597 (N_597,In_1605,In_952);
nor U598 (N_598,In_2008,In_2958);
nand U599 (N_599,In_1707,In_2297);
or U600 (N_600,In_1424,In_1451);
nand U601 (N_601,In_688,In_628);
and U602 (N_602,In_1181,In_1820);
xnor U603 (N_603,In_2428,In_161);
nor U604 (N_604,In_1338,In_2963);
and U605 (N_605,In_1821,In_1081);
xor U606 (N_606,In_41,In_1680);
xnor U607 (N_607,In_2850,In_959);
nor U608 (N_608,In_2868,In_1320);
or U609 (N_609,In_718,In_2209);
or U610 (N_610,In_1164,In_224);
and U611 (N_611,In_1210,In_1323);
xor U612 (N_612,In_2921,In_2522);
nor U613 (N_613,In_420,In_2472);
nand U614 (N_614,In_407,In_2144);
xnor U615 (N_615,In_1120,In_2999);
nand U616 (N_616,In_1698,In_1720);
nor U617 (N_617,In_1917,In_913);
nor U618 (N_618,In_455,In_852);
nor U619 (N_619,In_1431,In_1079);
nor U620 (N_620,In_2099,In_2259);
and U621 (N_621,In_1567,In_2146);
xnor U622 (N_622,In_2972,In_1318);
nor U623 (N_623,In_297,In_2183);
xnor U624 (N_624,In_432,In_1121);
and U625 (N_625,In_61,In_790);
nand U626 (N_626,In_2847,In_1985);
nor U627 (N_627,In_342,In_2452);
nand U628 (N_628,In_2192,In_2390);
and U629 (N_629,In_294,In_2020);
nand U630 (N_630,In_84,In_1464);
nand U631 (N_631,In_2107,In_1290);
nor U632 (N_632,In_2327,In_1372);
xor U633 (N_633,In_2672,In_2493);
xor U634 (N_634,In_733,In_295);
xnor U635 (N_635,In_1058,In_1479);
nand U636 (N_636,In_2681,In_18);
or U637 (N_637,In_2064,In_1404);
and U638 (N_638,In_1311,In_926);
nor U639 (N_639,In_2621,In_403);
nand U640 (N_640,In_1976,In_2938);
and U641 (N_641,In_1601,In_2063);
nand U642 (N_642,In_2666,In_2777);
nor U643 (N_643,In_1376,In_570);
xnor U644 (N_644,In_726,In_2310);
nor U645 (N_645,In_671,In_2658);
nand U646 (N_646,In_167,In_309);
nor U647 (N_647,In_1145,In_289);
and U648 (N_648,In_912,In_812);
and U649 (N_649,In_2025,In_1775);
nor U650 (N_650,In_2646,In_781);
xor U651 (N_651,In_2937,In_184);
nand U652 (N_652,In_2977,In_824);
or U653 (N_653,In_2031,In_87);
nor U654 (N_654,In_1036,In_2694);
xor U655 (N_655,In_156,In_2700);
nand U656 (N_656,In_664,In_2346);
nor U657 (N_657,In_766,In_2303);
and U658 (N_658,In_1949,In_1169);
nand U659 (N_659,In_731,In_2742);
and U660 (N_660,In_842,In_2880);
and U661 (N_661,In_1969,In_1363);
or U662 (N_662,In_2805,In_2070);
nand U663 (N_663,In_881,In_1256);
or U664 (N_664,In_2652,In_1385);
nor U665 (N_665,In_2061,In_765);
or U666 (N_666,In_2231,In_2034);
xnor U667 (N_667,In_1769,In_1119);
or U668 (N_668,In_1931,In_137);
xor U669 (N_669,In_533,In_1371);
nand U670 (N_670,In_1954,In_2575);
or U671 (N_671,In_1140,In_2167);
nor U672 (N_672,In_550,In_101);
nor U673 (N_673,In_1548,In_1142);
and U674 (N_674,In_484,In_222);
and U675 (N_675,In_1098,In_1258);
and U676 (N_676,In_802,In_2641);
nor U677 (N_677,In_435,In_1842);
nor U678 (N_678,In_1534,In_1259);
nor U679 (N_679,In_304,In_2602);
nor U680 (N_680,In_1612,In_1015);
or U681 (N_681,In_153,In_1024);
and U682 (N_682,In_1924,In_1444);
xor U683 (N_683,In_422,In_759);
nand U684 (N_684,In_298,In_1227);
xor U685 (N_685,In_1002,In_2122);
nor U686 (N_686,In_2489,In_1872);
nor U687 (N_687,In_1621,In_719);
nand U688 (N_688,In_2286,In_362);
xnor U689 (N_689,In_307,In_535);
nor U690 (N_690,In_662,In_2595);
xnor U691 (N_691,In_2399,In_1266);
nor U692 (N_692,In_2147,In_1253);
or U693 (N_693,In_1864,In_1814);
nand U694 (N_694,In_1501,In_2584);
xnor U695 (N_695,In_182,In_2560);
nand U696 (N_696,In_1767,In_774);
and U697 (N_697,In_383,In_1417);
and U698 (N_698,In_1606,In_1519);
nor U699 (N_699,In_339,In_1069);
nor U700 (N_700,In_1561,In_862);
or U701 (N_701,In_2563,In_1313);
and U702 (N_702,In_1614,In_2163);
nor U703 (N_703,In_158,In_2865);
and U704 (N_704,In_1352,In_2506);
nand U705 (N_705,In_1998,In_984);
xor U706 (N_706,In_794,In_428);
or U707 (N_707,In_2134,In_2717);
nor U708 (N_708,In_355,In_1977);
and U709 (N_709,In_2507,In_447);
and U710 (N_710,In_2791,In_1549);
nand U711 (N_711,In_2221,In_1212);
xor U712 (N_712,In_2559,In_1728);
xor U713 (N_713,In_1096,In_1719);
or U714 (N_714,In_2636,In_2028);
or U715 (N_715,In_1877,In_206);
xor U716 (N_716,In_1187,In_2236);
nand U717 (N_717,In_2804,In_1391);
and U718 (N_718,In_1771,In_720);
nand U719 (N_719,In_2026,In_431);
xnor U720 (N_720,In_1229,In_2185);
nand U721 (N_721,In_2935,In_1747);
and U722 (N_722,In_1452,In_2629);
and U723 (N_723,In_753,In_2857);
and U724 (N_724,In_1540,In_2826);
nand U725 (N_725,In_2060,In_1554);
nor U726 (N_726,In_2415,In_756);
or U727 (N_727,In_413,In_449);
xor U728 (N_728,In_1684,In_2922);
or U729 (N_729,In_332,In_2957);
nand U730 (N_730,In_2597,In_2549);
nor U731 (N_731,In_1751,In_2152);
or U732 (N_732,In_2179,In_2839);
and U733 (N_733,In_160,In_836);
or U734 (N_734,In_1050,In_1204);
nand U735 (N_735,In_2342,In_1866);
nor U736 (N_736,In_981,In_1301);
xor U737 (N_737,In_1059,In_1478);
nand U738 (N_738,In_690,In_2218);
nor U739 (N_739,In_330,In_1533);
xor U740 (N_740,In_1739,In_2345);
and U741 (N_741,In_1356,In_2331);
nand U742 (N_742,In_1470,In_1292);
nand U743 (N_743,In_2484,In_1843);
xor U744 (N_744,In_2368,In_1511);
xor U745 (N_745,In_23,In_654);
nand U746 (N_746,In_678,In_2305);
and U747 (N_747,In_1610,In_1564);
nand U748 (N_748,In_2886,In_1314);
and U749 (N_749,In_1116,In_549);
xnor U750 (N_750,In_2982,In_228);
nand U751 (N_751,In_1270,In_2569);
nor U752 (N_752,In_652,In_1232);
nor U753 (N_753,In_1727,In_424);
or U754 (N_754,In_1712,In_792);
or U755 (N_755,In_1130,In_2412);
xnor U756 (N_756,In_594,In_205);
nor U757 (N_757,In_2039,In_1966);
xnor U758 (N_758,In_2713,In_2496);
nand U759 (N_759,In_2369,In_260);
or U760 (N_760,In_271,In_2398);
and U761 (N_761,In_2265,In_2917);
nand U762 (N_762,In_2012,In_268);
nor U763 (N_763,In_498,In_1708);
and U764 (N_764,In_2598,In_1922);
nand U765 (N_765,In_303,In_452);
nor U766 (N_766,In_241,In_2662);
xnor U767 (N_767,In_1804,In_637);
and U768 (N_768,In_2204,In_2250);
and U769 (N_769,In_2578,In_2326);
nor U770 (N_770,In_668,In_2831);
nand U771 (N_771,In_2454,In_1619);
or U772 (N_772,In_410,In_2561);
xor U773 (N_773,In_349,In_1009);
nand U774 (N_774,In_1822,In_81);
nor U775 (N_775,In_1104,In_1085);
nand U776 (N_776,In_894,In_1858);
or U777 (N_777,In_1967,In_738);
xor U778 (N_778,In_2676,In_2131);
nor U779 (N_779,In_987,In_1214);
nand U780 (N_780,In_136,In_2699);
xnor U781 (N_781,In_2051,In_2984);
nand U782 (N_782,In_858,In_2351);
and U783 (N_783,In_1935,In_1437);
nand U784 (N_784,In_1937,In_2339);
nand U785 (N_785,In_149,In_2593);
and U786 (N_786,In_1799,In_1382);
and U787 (N_787,In_116,In_801);
or U788 (N_788,In_1770,In_2127);
or U789 (N_789,In_2843,In_2292);
and U790 (N_790,In_1027,In_246);
and U791 (N_791,In_1847,In_175);
nor U792 (N_792,In_1215,In_1094);
or U793 (N_793,In_904,In_2187);
xor U794 (N_794,In_2586,In_1525);
or U795 (N_795,In_174,In_50);
nand U796 (N_796,In_20,In_11);
and U797 (N_797,In_556,In_854);
or U798 (N_798,In_903,In_2058);
xor U799 (N_799,In_1632,In_1711);
nor U800 (N_800,In_1848,In_415);
xnor U801 (N_801,In_1249,In_843);
nor U802 (N_802,In_1682,In_1032);
or U803 (N_803,In_845,In_2927);
xor U804 (N_804,In_2590,In_2104);
xnor U805 (N_805,In_2827,In_1241);
xnor U806 (N_806,In_108,In_29);
nand U807 (N_807,In_2819,In_1898);
xor U808 (N_808,In_798,In_2863);
nor U809 (N_809,In_1890,In_15);
or U810 (N_810,In_138,In_1857);
or U811 (N_811,In_835,In_26);
and U812 (N_812,In_703,In_931);
nand U813 (N_813,In_1603,In_1262);
nor U814 (N_814,In_2833,In_627);
and U815 (N_815,In_2275,In_2543);
nor U816 (N_816,In_2987,In_1369);
xnor U817 (N_817,In_2867,In_966);
xnor U818 (N_818,In_2746,In_2145);
xnor U819 (N_819,In_263,In_1607);
and U820 (N_820,In_816,In_683);
or U821 (N_821,In_832,In_2724);
nor U822 (N_822,In_2154,In_1617);
nor U823 (N_823,In_2299,In_2437);
or U824 (N_824,In_2635,In_797);
xnor U825 (N_825,In_1180,In_1868);
xor U826 (N_826,In_709,In_1781);
or U827 (N_827,In_1963,In_2969);
nor U828 (N_828,In_384,In_288);
xnor U829 (N_829,In_520,In_982);
xor U830 (N_830,In_524,In_1686);
nor U831 (N_831,In_1460,In_755);
xor U832 (N_832,In_811,In_1660);
nor U833 (N_833,In_1288,In_1469);
xor U834 (N_834,In_144,In_1150);
nand U835 (N_835,In_1726,In_2284);
nor U836 (N_836,In_1960,In_2196);
xnor U837 (N_837,In_326,In_1956);
and U838 (N_838,In_2715,In_150);
nor U839 (N_839,In_1681,In_1809);
nand U840 (N_840,In_2426,In_754);
or U841 (N_841,In_517,In_2651);
and U842 (N_842,In_2637,In_462);
nor U843 (N_843,In_2219,In_1086);
nor U844 (N_844,In_2776,In_1022);
nor U845 (N_845,In_2075,In_2906);
nand U846 (N_846,In_725,In_311);
nor U847 (N_847,In_1572,In_2912);
nor U848 (N_848,In_306,In_1393);
and U849 (N_849,In_1827,In_909);
nand U850 (N_850,In_892,In_1749);
nand U851 (N_851,In_1576,In_473);
xor U852 (N_852,In_1604,In_1357);
or U853 (N_853,In_2743,In_2085);
xnor U854 (N_854,In_927,In_2273);
or U855 (N_855,In_1685,In_1195);
and U856 (N_856,In_2024,In_1611);
nand U857 (N_857,In_907,In_1492);
xnor U858 (N_858,In_1818,In_943);
nor U859 (N_859,In_1667,In_911);
nor U860 (N_860,In_1244,In_2360);
nand U861 (N_861,In_2469,In_2813);
nand U862 (N_862,In_1344,In_2878);
nor U863 (N_863,In_1768,In_2115);
or U864 (N_864,In_1745,In_944);
nor U865 (N_865,In_721,In_1740);
xnor U866 (N_866,In_1073,In_238);
or U867 (N_867,In_1366,In_203);
xor U868 (N_868,In_2577,In_2690);
nor U869 (N_869,In_749,In_2895);
xnor U870 (N_870,In_1486,In_142);
nand U871 (N_871,In_1354,In_863);
or U872 (N_872,In_822,In_639);
nand U873 (N_873,In_2923,In_623);
xnor U874 (N_874,In_732,In_803);
xor U875 (N_875,In_1746,In_2291);
xor U876 (N_876,In_940,In_773);
or U877 (N_877,In_1127,In_506);
nor U878 (N_878,In_1476,In_1724);
or U879 (N_879,In_1211,In_1517);
and U880 (N_880,In_800,In_463);
and U881 (N_881,In_272,In_2344);
and U882 (N_882,In_1715,In_2749);
nor U883 (N_883,In_1386,In_448);
nor U884 (N_884,In_345,In_2914);
xnor U885 (N_885,In_2695,In_1886);
or U886 (N_886,In_290,In_2016);
xor U887 (N_887,In_2290,In_2117);
nand U888 (N_888,In_480,In_2564);
or U889 (N_889,In_1646,In_1744);
and U890 (N_890,In_1165,In_2392);
or U891 (N_891,In_147,In_1182);
nand U892 (N_892,In_2332,In_2463);
or U893 (N_893,In_579,In_614);
nor U894 (N_894,In_244,In_1020);
and U895 (N_895,In_1454,In_2565);
or U896 (N_896,In_2540,In_343);
and U897 (N_897,In_1048,In_282);
and U898 (N_898,In_2781,In_2554);
or U899 (N_899,In_2205,In_1647);
or U900 (N_900,In_33,In_1638);
nor U901 (N_901,In_264,In_2487);
nand U902 (N_902,In_1526,In_1472);
or U903 (N_903,In_1347,In_2622);
xnor U904 (N_904,In_2383,In_2950);
nand U905 (N_905,In_657,In_2402);
and U906 (N_906,In_302,In_1016);
nor U907 (N_907,In_739,In_308);
nor U908 (N_908,In_2446,In_1892);
nand U909 (N_909,In_2320,In_1811);
xor U910 (N_910,In_1054,In_2870);
nor U911 (N_911,In_2086,In_1794);
or U912 (N_912,In_1512,In_176);
nor U913 (N_913,In_633,In_1345);
and U914 (N_914,In_2128,In_1823);
xor U915 (N_915,In_2087,In_103);
nor U916 (N_916,In_764,In_1995);
xnor U917 (N_917,In_1309,In_1343);
or U918 (N_918,In_2760,In_262);
nor U919 (N_919,In_67,In_2901);
xor U920 (N_920,In_1066,In_2436);
nand U921 (N_921,In_1035,In_2708);
nand U922 (N_922,In_928,In_655);
or U923 (N_923,In_937,In_939);
xnor U924 (N_924,In_369,In_2419);
and U925 (N_925,In_2928,In_98);
xnor U926 (N_926,In_2433,In_1412);
nand U927 (N_927,In_934,In_2612);
xor U928 (N_928,In_201,In_2820);
or U929 (N_929,In_2438,In_876);
xor U930 (N_930,In_2626,In_918);
xnor U931 (N_931,In_1785,In_728);
nand U932 (N_932,In_834,In_1118);
or U933 (N_933,In_2417,In_2890);
nor U934 (N_934,In_2211,In_357);
xnor U935 (N_935,In_2488,In_2227);
nand U936 (N_936,In_1038,In_69);
xor U937 (N_937,In_2395,In_1897);
nor U938 (N_938,In_1752,In_388);
or U939 (N_939,In_111,In_823);
xor U940 (N_940,In_813,In_1507);
or U941 (N_941,In_385,In_2448);
or U942 (N_942,In_1457,In_2693);
and U943 (N_943,In_2220,In_917);
nor U944 (N_944,In_2818,In_1302);
and U945 (N_945,In_2444,In_323);
xor U946 (N_946,In_2214,In_1029);
nor U947 (N_947,In_704,In_1670);
nor U948 (N_948,In_261,In_1962);
nor U949 (N_949,In_569,In_2241);
and U950 (N_950,In_2388,In_1293);
nand U951 (N_951,In_487,In_123);
or U952 (N_952,In_826,In_1800);
and U953 (N_953,In_2803,In_979);
nor U954 (N_954,In_961,In_377);
nor U955 (N_955,In_2062,In_2986);
nor U956 (N_956,In_998,In_396);
nor U957 (N_957,In_1091,In_2243);
xor U958 (N_958,In_867,In_1655);
nor U959 (N_959,In_1885,In_1543);
and U960 (N_960,In_1219,In_775);
nand U961 (N_961,In_789,In_1974);
xnor U962 (N_962,In_1531,In_2680);
xor U963 (N_963,In_2623,In_1978);
and U964 (N_964,In_1553,In_216);
nand U965 (N_965,In_1415,In_1271);
or U966 (N_966,In_2888,In_750);
xnor U967 (N_967,In_37,In_1201);
xor U968 (N_968,In_1324,In_1421);
and U969 (N_969,In_1315,In_2797);
or U970 (N_970,In_2005,In_1510);
or U971 (N_971,In_1582,In_1171);
xnor U972 (N_972,In_1547,In_2916);
nand U973 (N_973,In_870,In_1594);
or U974 (N_974,In_1389,In_2656);
or U975 (N_975,In_78,In_1088);
nor U976 (N_976,In_1129,In_869);
and U977 (N_977,In_1252,In_2858);
nor U978 (N_978,In_1948,In_503);
xor U979 (N_979,In_1677,In_1591);
or U980 (N_980,In_2795,In_75);
or U981 (N_981,In_1790,In_2603);
and U982 (N_982,In_2907,In_2970);
and U983 (N_983,In_2948,In_514);
nor U984 (N_984,In_2789,In_2396);
or U985 (N_985,In_2465,In_971);
nand U986 (N_986,In_2042,In_2281);
and U987 (N_987,In_2481,In_1983);
or U988 (N_988,In_674,In_328);
and U989 (N_989,In_53,In_2479);
nand U990 (N_990,In_96,In_2256);
xnor U991 (N_991,In_1961,In_2689);
xor U992 (N_992,In_2468,In_2898);
or U993 (N_993,In_1473,In_2098);
or U994 (N_994,In_2609,In_411);
xnor U995 (N_995,In_433,In_59);
nand U996 (N_996,In_1555,In_1815);
nor U997 (N_997,In_748,In_1235);
nand U998 (N_998,In_186,In_2247);
nand U999 (N_999,In_1184,In_352);
nand U1000 (N_1000,In_1327,In_1179);
xor U1001 (N_1001,In_2420,In_218);
or U1002 (N_1002,In_2260,In_2976);
nor U1003 (N_1003,In_1287,In_1861);
and U1004 (N_1004,In_2574,In_1388);
nor U1005 (N_1005,In_1044,In_713);
or U1006 (N_1006,In_1322,In_670);
nand U1007 (N_1007,In_2993,In_502);
nor U1008 (N_1008,In_1025,In_837);
nand U1009 (N_1009,In_2139,In_2375);
nor U1010 (N_1010,In_2040,In_17);
and U1011 (N_1011,In_1414,In_996);
nand U1012 (N_1012,In_46,In_2410);
nand U1013 (N_1013,In_220,In_574);
xor U1014 (N_1014,In_954,In_2081);
nor U1015 (N_1015,In_181,In_2201);
nand U1016 (N_1016,In_2731,In_1306);
xnor U1017 (N_1017,In_2552,In_2810);
or U1018 (N_1018,In_1279,In_2347);
nor U1019 (N_1019,In_2169,In_459);
nor U1020 (N_1020,In_1796,In_906);
and U1021 (N_1021,In_1613,In_1207);
nand U1022 (N_1022,In_736,In_2720);
and U1023 (N_1023,In_483,In_2900);
xor U1024 (N_1024,In_2531,In_346);
nand U1025 (N_1025,In_2556,In_547);
and U1026 (N_1026,In_2642,In_31);
xor U1027 (N_1027,In_1321,In_534);
and U1028 (N_1028,In_865,In_955);
nand U1029 (N_1029,In_223,In_2233);
xnor U1030 (N_1030,In_1900,In_1889);
xnor U1031 (N_1031,In_287,In_2624);
and U1032 (N_1032,In_1283,In_806);
and U1033 (N_1033,In_2755,In_2885);
nand U1034 (N_1034,In_2854,In_1731);
or U1035 (N_1035,In_2384,In_337);
xnor U1036 (N_1036,In_661,In_1903);
nor U1037 (N_1037,In_949,In_1938);
nor U1038 (N_1038,In_2013,In_2691);
and U1039 (N_1039,In_545,In_962);
or U1040 (N_1040,In_651,In_902);
nand U1041 (N_1041,In_2044,In_1629);
or U1042 (N_1042,In_1124,In_540);
nor U1043 (N_1043,In_1095,In_1696);
and U1044 (N_1044,In_2442,In_1763);
or U1045 (N_1045,In_145,In_2544);
and U1046 (N_1046,In_2775,In_2414);
nand U1047 (N_1047,In_2956,In_210);
xnor U1048 (N_1048,In_1497,In_38);
and U1049 (N_1049,In_162,In_1102);
xnor U1050 (N_1050,In_2217,In_109);
and U1051 (N_1051,In_1206,In_1475);
xor U1052 (N_1052,In_1167,In_2978);
and U1053 (N_1053,In_77,In_1328);
xnor U1054 (N_1054,In_2073,In_270);
nand U1055 (N_1055,In_2539,In_1373);
or U1056 (N_1056,In_2796,In_427);
nor U1057 (N_1057,In_855,In_2601);
and U1058 (N_1058,In_1075,In_1870);
nor U1059 (N_1059,In_796,In_636);
or U1060 (N_1060,In_2257,In_877);
or U1061 (N_1061,In_165,In_94);
or U1062 (N_1062,In_905,In_2740);
or U1063 (N_1063,In_2308,In_1465);
or U1064 (N_1064,In_508,In_2003);
and U1065 (N_1065,In_970,In_1286);
xor U1066 (N_1066,In_564,In_602);
nand U1067 (N_1067,In_714,In_2267);
xnor U1068 (N_1068,In_2080,In_1888);
or U1069 (N_1069,In_990,In_380);
xor U1070 (N_1070,In_2942,In_1221);
or U1071 (N_1071,In_1131,In_2639);
or U1072 (N_1072,In_631,In_1355);
and U1073 (N_1073,In_2670,In_2239);
and U1074 (N_1074,In_1883,In_170);
nor U1075 (N_1075,In_2718,In_49);
and U1076 (N_1076,In_2023,In_1793);
and U1077 (N_1077,In_1051,In_2222);
or U1078 (N_1078,In_1909,In_1205);
nand U1079 (N_1079,In_2373,In_390);
nor U1080 (N_1080,In_2019,In_2659);
and U1081 (N_1081,In_1757,In_2811);
and U1082 (N_1082,In_2949,In_2975);
nand U1083 (N_1083,In_2677,In_1595);
nor U1084 (N_1084,In_1587,In_857);
and U1085 (N_1085,In_1926,In_1291);
or U1086 (N_1086,In_1873,In_2732);
or U1087 (N_1087,In_2316,In_2961);
nor U1088 (N_1088,In_2761,In_2997);
nand U1089 (N_1089,In_776,In_2734);
and U1090 (N_1090,In_2745,In_1365);
nand U1091 (N_1091,In_1143,In_2832);
or U1092 (N_1092,In_921,In_745);
nor U1093 (N_1093,In_2683,In_1556);
xnor U1094 (N_1094,In_985,In_777);
or U1095 (N_1095,In_1669,In_707);
and U1096 (N_1096,In_2980,In_2606);
xnor U1097 (N_1097,In_2272,In_406);
or U1098 (N_1098,In_1390,In_2212);
or U1099 (N_1099,In_1060,In_624);
xnor U1100 (N_1100,In_1608,In_1335);
or U1101 (N_1101,In_1358,In_133);
nor U1102 (N_1102,In_1448,In_2181);
nor U1103 (N_1103,In_1337,In_925);
nand U1104 (N_1104,In_1869,In_2065);
or U1105 (N_1105,In_334,In_236);
nand U1106 (N_1106,In_669,In_1773);
nand U1107 (N_1107,In_2794,In_239);
or U1108 (N_1108,In_2862,In_1031);
xnor U1109 (N_1109,In_2224,In_2784);
and U1110 (N_1110,In_482,In_157);
xnor U1111 (N_1111,In_365,In_2915);
nand U1112 (N_1112,In_1879,In_1381);
or U1113 (N_1113,In_2758,In_1874);
nor U1114 (N_1114,In_770,In_2068);
or U1115 (N_1115,In_1202,In_2123);
nor U1116 (N_1116,In_376,In_1053);
nor U1117 (N_1117,In_2159,In_511);
nand U1118 (N_1118,In_2864,In_1934);
nor U1119 (N_1119,In_2729,In_1832);
or U1120 (N_1120,In_1402,In_778);
nand U1121 (N_1121,In_2667,In_2245);
nand U1122 (N_1122,In_2640,In_168);
or U1123 (N_1123,In_767,In_374);
and U1124 (N_1124,In_1951,In_2508);
nor U1125 (N_1125,In_895,In_119);
and U1126 (N_1126,In_504,In_2249);
and U1127 (N_1127,In_2175,In_997);
or U1128 (N_1128,In_2521,In_2177);
or U1129 (N_1129,In_1146,In_2223);
nand U1130 (N_1130,In_1831,In_2379);
xnor U1131 (N_1131,In_1738,In_1899);
nor U1132 (N_1132,In_527,In_1907);
xnor U1133 (N_1133,In_1701,In_587);
or U1134 (N_1134,In_893,In_2785);
or U1135 (N_1135,In_2911,In_606);
and U1136 (N_1136,In_1008,In_2882);
xnor U1137 (N_1137,In_143,In_2166);
and U1138 (N_1138,In_2709,In_2427);
nand U1139 (N_1139,In_194,In_2939);
or U1140 (N_1140,In_95,In_2904);
or U1141 (N_1141,In_2650,In_2244);
or U1142 (N_1142,In_2255,In_2716);
and U1143 (N_1143,In_872,In_2206);
and U1144 (N_1144,In_1226,In_2287);
nand U1145 (N_1145,In_1902,In_2215);
or U1146 (N_1146,In_2162,In_2509);
and U1147 (N_1147,In_676,In_333);
nand U1148 (N_1148,In_280,In_525);
nand U1149 (N_1149,In_1434,In_1615);
xnor U1150 (N_1150,In_1077,In_947);
nor U1151 (N_1151,In_1999,In_923);
xor U1152 (N_1152,In_2476,In_1455);
or U1153 (N_1153,In_1717,In_2814);
nand U1154 (N_1154,In_496,In_1628);
nand U1155 (N_1155,In_387,In_2947);
or U1156 (N_1156,In_724,In_2359);
and U1157 (N_1157,In_744,In_1360);
and U1158 (N_1158,In_1923,In_141);
or U1159 (N_1159,In_1714,In_1518);
or U1160 (N_1160,In_479,In_2004);
or U1161 (N_1161,In_1004,In_1571);
and U1162 (N_1162,In_269,In_1508);
xnor U1163 (N_1163,In_599,In_442);
xnor U1164 (N_1164,In_476,In_2010);
or U1165 (N_1165,In_2203,In_2293);
nand U1166 (N_1166,In_2892,In_1097);
nor U1167 (N_1167,In_1325,In_538);
xnor U1168 (N_1168,In_1161,In_1675);
xor U1169 (N_1169,In_769,In_1001);
and U1170 (N_1170,In_1070,In_2891);
xor U1171 (N_1171,In_2178,In_589);
xnor U1172 (N_1172,In_151,In_1538);
or U1173 (N_1173,In_363,In_1420);
or U1174 (N_1174,In_122,In_1710);
and U1175 (N_1175,In_1565,In_2585);
nand U1176 (N_1176,In_2661,In_1642);
nor U1177 (N_1177,In_375,In_1589);
xor U1178 (N_1178,In_1435,In_2407);
or U1179 (N_1179,In_2382,In_1844);
nand U1180 (N_1180,In_1316,In_1665);
nand U1181 (N_1181,In_2449,In_2198);
nor U1182 (N_1182,In_1394,In_2301);
and U1183 (N_1183,In_2538,In_785);
xnor U1184 (N_1184,In_1597,In_495);
nor U1185 (N_1185,In_1006,In_212);
and U1186 (N_1186,In_250,In_1217);
nand U1187 (N_1187,In_1735,In_2149);
nor U1188 (N_1188,In_539,In_743);
xor U1189 (N_1189,In_730,In_2995);
nor U1190 (N_1190,In_1537,In_1852);
and U1191 (N_1191,In_879,In_1859);
nand U1192 (N_1192,In_2669,In_1803);
nand U1193 (N_1193,In_198,In_2113);
or U1194 (N_1194,In_2605,In_2271);
xor U1195 (N_1195,In_341,In_659);
or U1196 (N_1196,In_1269,In_600);
xor U1197 (N_1197,In_1672,In_2955);
xor U1198 (N_1198,In_2029,In_256);
nand U1199 (N_1199,In_2765,In_2910);
or U1200 (N_1200,In_2378,In_575);
nand U1201 (N_1201,In_849,In_2366);
or U1202 (N_1202,In_1197,In_829);
nor U1203 (N_1203,In_737,In_2225);
xnor U1204 (N_1204,In_619,In_2445);
xor U1205 (N_1205,In_1918,In_25);
xor U1206 (N_1206,In_581,In_1552);
nand U1207 (N_1207,In_65,In_2045);
nor U1208 (N_1208,In_708,In_276);
nor U1209 (N_1209,In_1450,In_1333);
nand U1210 (N_1210,In_74,In_2325);
nor U1211 (N_1211,In_810,In_409);
xnor U1212 (N_1212,In_1654,In_1562);
nor U1213 (N_1213,In_2397,In_325);
and U1214 (N_1214,In_2471,In_665);
nor U1215 (N_1215,In_715,In_2524);
or U1216 (N_1216,In_2744,In_839);
xor U1217 (N_1217,In_1295,In_1690);
nand U1218 (N_1218,In_2608,In_1583);
or U1219 (N_1219,In_666,In_1246);
nand U1220 (N_1220,In_2768,In_207);
xor U1221 (N_1221,In_2934,In_118);
xnor U1222 (N_1222,In_1012,In_941);
nand U1223 (N_1223,In_257,In_557);
or U1224 (N_1224,In_2703,In_1959);
and U1225 (N_1225,In_2477,In_1980);
or U1226 (N_1226,In_1078,In_1128);
xnor U1227 (N_1227,In_562,In_1792);
xor U1228 (N_1228,In_2450,In_312);
nor U1229 (N_1229,In_1920,In_48);
nand U1230 (N_1230,In_1103,In_1854);
xor U1231 (N_1231,In_1586,In_425);
and U1232 (N_1232,In_701,In_685);
or U1233 (N_1233,In_300,In_434);
and U1234 (N_1234,In_1851,In_2532);
and U1235 (N_1235,In_2710,In_850);
and U1236 (N_1236,In_2499,In_1043);
xor U1237 (N_1237,In_99,In_2959);
or U1238 (N_1238,In_1971,In_2264);
or U1239 (N_1239,In_1819,In_1494);
xnor U1240 (N_1240,In_1723,In_559);
nand U1241 (N_1241,In_2665,In_827);
or U1242 (N_1242,In_2391,In_71);
nand U1243 (N_1243,In_2251,In_360);
or U1244 (N_1244,In_202,In_1996);
and U1245 (N_1245,In_191,In_953);
nand U1246 (N_1246,In_1304,In_2151);
and U1247 (N_1247,In_791,In_2990);
xor U1248 (N_1248,In_900,In_1623);
or U1249 (N_1249,In_1332,In_2772);
xnor U1250 (N_1250,In_1970,In_73);
nor U1251 (N_1251,In_2799,In_681);
and U1252 (N_1252,In_2853,In_2353);
or U1253 (N_1253,In_1147,In_2307);
nand U1254 (N_1254,In_2798,In_2591);
nand U1255 (N_1255,In_2334,In_1774);
xnor U1256 (N_1256,In_2727,In_2180);
or U1257 (N_1257,In_2872,In_2197);
or U1258 (N_1258,In_1649,In_2076);
and U1259 (N_1259,In_2425,In_584);
xor U1260 (N_1260,In_1234,In_2954);
xnor U1261 (N_1261,In_2836,In_490);
nor U1262 (N_1262,In_1581,In_948);
nand U1263 (N_1263,In_1755,In_861);
or U1264 (N_1264,In_2050,In_1699);
xnor U1265 (N_1265,In_2762,In_868);
or U1266 (N_1266,In_2766,In_423);
xor U1267 (N_1267,In_2037,In_1506);
nand U1268 (N_1268,In_2952,In_336);
or U1269 (N_1269,In_523,In_39);
and U1270 (N_1270,In_2649,In_2875);
xnor U1271 (N_1271,In_331,In_347);
and U1272 (N_1272,In_1107,In_115);
nor U1273 (N_1273,In_2903,In_8);
nand U1274 (N_1274,In_2807,In_883);
nand U1275 (N_1275,In_57,In_1791);
nor U1276 (N_1276,In_2278,In_127);
nor U1277 (N_1277,In_1812,In_536);
or U1278 (N_1278,In_2657,In_1721);
and U1279 (N_1279,In_1138,In_1477);
or U1280 (N_1280,In_70,In_1560);
and U1281 (N_1281,In_762,In_2041);
or U1282 (N_1282,In_2018,In_1458);
or U1283 (N_1283,In_0,In_1641);
nand U1284 (N_1284,In_1836,In_1353);
and U1285 (N_1285,In_125,In_1958);
xnor U1286 (N_1286,In_2615,In_740);
nand U1287 (N_1287,In_859,In_884);
nor U1288 (N_1288,In_2873,In_2932);
or U1289 (N_1289,In_1697,In_1616);
or U1290 (N_1290,In_2719,In_1003);
xnor U1291 (N_1291,In_2511,In_1705);
or U1292 (N_1292,In_2208,In_2548);
nand U1293 (N_1293,In_1579,In_1483);
or U1294 (N_1294,In_2377,In_634);
nand U1295 (N_1295,In_1178,In_684);
nand U1296 (N_1296,In_259,In_1991);
nand U1297 (N_1297,In_1578,In_2424);
nand U1298 (N_1298,In_620,In_2401);
or U1299 (N_1299,In_1416,In_292);
and U1300 (N_1300,In_2611,In_833);
nor U1301 (N_1301,In_2140,In_2757);
xor U1302 (N_1302,In_1893,In_335);
and U1303 (N_1303,In_2860,In_1499);
nor U1304 (N_1304,In_2557,In_1379);
nand U1305 (N_1305,In_90,In_1375);
or U1306 (N_1306,In_2534,In_1945);
or U1307 (N_1307,In_935,In_2829);
nor U1308 (N_1308,In_2616,In_2309);
nand U1309 (N_1309,In_771,In_1125);
or U1310 (N_1310,In_793,In_1289);
and U1311 (N_1311,In_1990,In_1166);
nand U1312 (N_1312,In_1340,In_2502);
xnor U1313 (N_1313,In_242,In_2547);
nor U1314 (N_1314,In_1734,In_2879);
and U1315 (N_1315,In_2036,In_121);
nor U1316 (N_1316,In_1750,In_1294);
and U1317 (N_1317,In_1028,In_658);
nand U1318 (N_1318,In_1786,In_702);
and U1319 (N_1319,In_1599,In_1196);
and U1320 (N_1320,In_601,In_2143);
nand U1321 (N_1321,In_2859,In_2296);
and U1322 (N_1322,In_2381,In_154);
and U1323 (N_1323,In_1272,In_605);
nor U1324 (N_1324,In_2408,In_1981);
and U1325 (N_1325,In_2643,In_2884);
or U1326 (N_1326,In_252,In_1895);
xor U1327 (N_1327,In_1986,In_185);
xnor U1328 (N_1328,In_1753,In_609);
xor U1329 (N_1329,In_1973,In_1795);
nor U1330 (N_1330,In_1277,In_1087);
xor U1331 (N_1331,In_699,In_1813);
xor U1332 (N_1332,In_1114,In_1758);
or U1333 (N_1333,In_492,In_436);
nor U1334 (N_1334,In_518,In_1810);
xor U1335 (N_1335,In_1853,In_2545);
nor U1336 (N_1336,In_675,In_129);
and U1337 (N_1337,In_995,In_752);
xor U1338 (N_1338,In_1908,In_254);
nand U1339 (N_1339,In_2964,In_131);
xor U1340 (N_1340,In_1661,In_717);
xnor U1341 (N_1341,In_578,In_1573);
or U1342 (N_1342,In_472,In_2289);
and U1343 (N_1343,In_2032,In_1856);
xnor U1344 (N_1344,In_1802,In_1064);
nor U1345 (N_1345,In_2280,In_1630);
nor U1346 (N_1346,In_104,In_531);
nand U1347 (N_1347,In_1063,In_130);
and U1348 (N_1348,In_1627,In_1248);
xor U1349 (N_1349,In_1111,In_607);
and U1350 (N_1350,In_597,In_2306);
or U1351 (N_1351,In_2160,In_2054);
nor U1352 (N_1352,In_1528,In_1504);
nor U1353 (N_1353,In_2082,In_1656);
or U1354 (N_1354,In_615,In_2248);
xor U1355 (N_1355,In_2685,In_611);
nand U1356 (N_1356,In_2348,In_885);
xor U1357 (N_1357,In_2240,In_2439);
nand U1358 (N_1358,In_734,In_1487);
nand U1359 (N_1359,In_2714,In_2485);
and U1360 (N_1360,In_1351,In_1694);
and U1361 (N_1361,In_680,In_44);
xnor U1362 (N_1362,In_2630,In_2919);
xnor U1363 (N_1363,In_139,In_1639);
nand U1364 (N_1364,In_117,In_2655);
or U1365 (N_1365,In_1952,In_2413);
nor U1366 (N_1366,In_1994,In_1509);
or U1367 (N_1367,In_1208,In_1835);
or U1368 (N_1368,In_1250,In_379);
nor U1369 (N_1369,In_172,In_2918);
nand U1370 (N_1370,In_251,In_976);
nor U1371 (N_1371,In_2129,In_2295);
nand U1372 (N_1372,In_2722,In_860);
and U1373 (N_1373,In_2721,In_179);
nand U1374 (N_1374,In_356,In_2678);
xor U1375 (N_1375,In_1410,In_1430);
nand U1376 (N_1376,In_1109,In_2817);
nand U1377 (N_1377,In_1919,In_1019);
xor U1378 (N_1378,In_2096,In_2090);
nor U1379 (N_1379,In_727,In_1602);
xor U1380 (N_1380,In_2526,In_679);
or U1381 (N_1381,In_1780,In_1788);
xnor U1382 (N_1382,In_1987,In_446);
and U1383 (N_1383,In_395,In_2808);
nor U1384 (N_1384,In_1849,In_1223);
xnor U1385 (N_1385,In_1846,In_1407);
xnor U1386 (N_1386,In_2116,In_1625);
or U1387 (N_1387,In_2748,In_2312);
and U1388 (N_1388,In_625,In_891);
nand U1389 (N_1389,In_30,In_93);
nand U1390 (N_1390,In_389,In_1782);
and U1391 (N_1391,In_193,In_1989);
and U1392 (N_1392,In_2494,In_2562);
and U1393 (N_1393,In_608,In_1401);
xnor U1394 (N_1394,In_2633,In_1551);
or U1395 (N_1395,In_35,In_1440);
xor U1396 (N_1396,In_957,In_2277);
nor U1397 (N_1397,In_113,In_645);
xnor U1398 (N_1398,In_501,In_1155);
nor U1399 (N_1399,In_2881,In_1305);
nor U1400 (N_1400,In_2435,In_461);
xnor U1401 (N_1401,In_197,In_1806);
and U1402 (N_1402,In_888,In_1299);
nor U1403 (N_1403,In_2349,In_233);
or U1404 (N_1404,In_640,In_437);
nor U1405 (N_1405,In_1093,In_825);
xnor U1406 (N_1406,In_1598,In_840);
or U1407 (N_1407,In_1280,In_213);
nand U1408 (N_1408,In_2202,In_2092);
nor U1409 (N_1409,In_2497,In_1840);
or U1410 (N_1410,In_787,In_516);
nor U1411 (N_1411,In_1979,In_2926);
and U1412 (N_1412,In_2838,In_267);
xor U1413 (N_1413,In_2941,In_1600);
nor U1414 (N_1414,In_1449,In_1493);
or U1415 (N_1415,In_1350,In_470);
or U1416 (N_1416,In_1784,In_1584);
xor U1417 (N_1417,In_397,In_2738);
or U1418 (N_1418,In_814,In_1162);
nand U1419 (N_1419,In_2883,In_2094);
and U1420 (N_1420,In_1018,In_1157);
or U1421 (N_1421,In_2625,In_2074);
or U1422 (N_1422,In_1648,In_2055);
nor U1423 (N_1423,In_1503,In_2333);
xor U1424 (N_1424,In_2246,In_2365);
nor U1425 (N_1425,In_1783,In_1838);
and U1426 (N_1426,In_630,In_2350);
xor U1427 (N_1427,In_1732,In_1072);
nand U1428 (N_1428,In_580,In_1575);
or U1429 (N_1429,In_635,In_967);
or U1430 (N_1430,In_694,In_1955);
or U1431 (N_1431,In_451,In_2017);
nand U1432 (N_1432,In_2052,In_2971);
and U1433 (N_1433,In_1423,In_177);
and U1434 (N_1434,In_1725,In_1255);
and U1435 (N_1435,In_2812,In_1175);
nor U1436 (N_1436,In_2541,In_2513);
xor U1437 (N_1437,In_1159,In_283);
and U1438 (N_1438,In_2866,In_2779);
nor U1439 (N_1439,In_1830,In_1468);
and U1440 (N_1440,In_2001,In_1566);
xor U1441 (N_1441,In_80,In_2505);
or U1442 (N_1442,In_2007,In_247);
or U1443 (N_1443,In_2258,In_1798);
xnor U1444 (N_1444,In_591,In_1777);
and U1445 (N_1445,In_2456,In_2989);
or U1446 (N_1446,In_2311,In_2793);
nand U1447 (N_1447,In_1144,In_226);
nor U1448 (N_1448,In_1964,In_277);
nor U1449 (N_1449,In_1062,In_1905);
and U1450 (N_1450,In_2077,In_890);
nand U1451 (N_1451,In_1912,In_2735);
xor U1452 (N_1452,In_40,In_371);
nor U1453 (N_1453,In_964,In_2186);
or U1454 (N_1454,In_977,In_1626);
nor U1455 (N_1455,In_1984,In_2242);
nand U1456 (N_1456,In_956,In_364);
xnor U1457 (N_1457,In_1650,In_2940);
or U1458 (N_1458,In_322,In_391);
nand U1459 (N_1459,In_1703,In_1521);
nor U1460 (N_1460,In_419,In_2756);
and U1461 (N_1461,In_1349,In_1296);
xor U1462 (N_1462,In_24,In_1658);
or U1463 (N_1463,In_124,In_1679);
and U1464 (N_1464,In_2992,In_500);
nand U1465 (N_1465,In_2455,In_305);
nand U1466 (N_1466,In_1557,In_2053);
or U1467 (N_1467,In_2682,In_68);
nand U1468 (N_1468,In_2043,In_2994);
xnor U1469 (N_1469,In_2276,In_1936);
or U1470 (N_1470,In_1418,In_398);
nor U1471 (N_1471,In_613,In_1334);
or U1472 (N_1472,In_2462,In_2723);
nor U1473 (N_1473,In_1257,In_512);
nor U1474 (N_1474,In_1123,In_1778);
and U1475 (N_1475,In_414,In_2988);
and U1476 (N_1476,In_846,In_2983);
and U1477 (N_1477,In_1436,In_1887);
nand U1478 (N_1478,In_1659,In_2706);
or U1479 (N_1479,In_1237,In_114);
nor U1480 (N_1480,In_2962,In_1634);
nand U1481 (N_1481,In_2367,In_2501);
or U1482 (N_1482,In_464,In_453);
or U1483 (N_1483,In_2132,In_1061);
nor U1484 (N_1484,In_505,In_1408);
xor U1485 (N_1485,In_475,In_2897);
xor U1486 (N_1486,In_6,In_2568);
nor U1487 (N_1487,In_1405,In_1933);
or U1488 (N_1488,In_1268,In_2841);
xnor U1489 (N_1489,In_2210,In_92);
or U1490 (N_1490,In_1947,In_2091);
nand U1491 (N_1491,In_1762,In_34);
xor U1492 (N_1492,In_2535,In_2386);
and U1493 (N_1493,In_1664,In_1906);
nor U1494 (N_1494,In_2546,In_1491);
xnor U1495 (N_1495,In_2790,In_1222);
nand U1496 (N_1496,In_2778,In_783);
or U1497 (N_1497,In_164,In_729);
nand U1498 (N_1498,In_2953,In_2529);
nor U1499 (N_1499,In_544,In_1488);
nor U1500 (N_1500,In_2077,In_2843);
and U1501 (N_1501,In_2062,In_1538);
xor U1502 (N_1502,In_1211,In_1745);
or U1503 (N_1503,In_1388,In_289);
nor U1504 (N_1504,In_2456,In_1609);
xnor U1505 (N_1505,In_2181,In_2863);
nand U1506 (N_1506,In_250,In_2656);
or U1507 (N_1507,In_27,In_2091);
nor U1508 (N_1508,In_1965,In_555);
nand U1509 (N_1509,In_1346,In_181);
or U1510 (N_1510,In_2336,In_2266);
nor U1511 (N_1511,In_1251,In_1813);
nand U1512 (N_1512,In_254,In_668);
or U1513 (N_1513,In_2267,In_1481);
xnor U1514 (N_1514,In_2815,In_2623);
and U1515 (N_1515,In_1790,In_1954);
nand U1516 (N_1516,In_1077,In_2619);
or U1517 (N_1517,In_2542,In_406);
xor U1518 (N_1518,In_125,In_864);
xor U1519 (N_1519,In_1490,In_1427);
nand U1520 (N_1520,In_2658,In_6);
and U1521 (N_1521,In_426,In_694);
or U1522 (N_1522,In_1913,In_1264);
nor U1523 (N_1523,In_2603,In_2291);
nand U1524 (N_1524,In_1588,In_635);
and U1525 (N_1525,In_2710,In_420);
xor U1526 (N_1526,In_2350,In_544);
and U1527 (N_1527,In_1012,In_2300);
or U1528 (N_1528,In_1752,In_656);
xor U1529 (N_1529,In_2900,In_24);
or U1530 (N_1530,In_1996,In_894);
and U1531 (N_1531,In_632,In_684);
xnor U1532 (N_1532,In_184,In_608);
or U1533 (N_1533,In_2261,In_353);
nand U1534 (N_1534,In_2917,In_2881);
nor U1535 (N_1535,In_2357,In_1478);
xnor U1536 (N_1536,In_2734,In_947);
and U1537 (N_1537,In_686,In_2996);
xor U1538 (N_1538,In_982,In_2506);
nor U1539 (N_1539,In_2320,In_1041);
nand U1540 (N_1540,In_2486,In_2626);
xor U1541 (N_1541,In_1641,In_1318);
nor U1542 (N_1542,In_1499,In_543);
nor U1543 (N_1543,In_478,In_232);
or U1544 (N_1544,In_2248,In_2725);
xor U1545 (N_1545,In_574,In_591);
or U1546 (N_1546,In_1793,In_2332);
nor U1547 (N_1547,In_1994,In_286);
or U1548 (N_1548,In_301,In_314);
xor U1549 (N_1549,In_1808,In_1000);
or U1550 (N_1550,In_689,In_2163);
nor U1551 (N_1551,In_236,In_679);
and U1552 (N_1552,In_485,In_455);
or U1553 (N_1553,In_2292,In_1990);
nor U1554 (N_1554,In_2059,In_2885);
xor U1555 (N_1555,In_1475,In_1094);
or U1556 (N_1556,In_1092,In_2385);
xnor U1557 (N_1557,In_683,In_1312);
xnor U1558 (N_1558,In_422,In_6);
xor U1559 (N_1559,In_434,In_2509);
nand U1560 (N_1560,In_1656,In_2723);
xor U1561 (N_1561,In_201,In_298);
or U1562 (N_1562,In_538,In_2069);
nand U1563 (N_1563,In_1409,In_187);
and U1564 (N_1564,In_308,In_1018);
xor U1565 (N_1565,In_31,In_1714);
nor U1566 (N_1566,In_465,In_1270);
and U1567 (N_1567,In_1996,In_604);
and U1568 (N_1568,In_643,In_1115);
xor U1569 (N_1569,In_2842,In_831);
nor U1570 (N_1570,In_30,In_2789);
xnor U1571 (N_1571,In_1961,In_2358);
xnor U1572 (N_1572,In_1202,In_509);
nand U1573 (N_1573,In_2472,In_1753);
xor U1574 (N_1574,In_1435,In_2117);
or U1575 (N_1575,In_1517,In_1215);
nand U1576 (N_1576,In_2023,In_1014);
nor U1577 (N_1577,In_1898,In_1674);
or U1578 (N_1578,In_451,In_410);
xor U1579 (N_1579,In_2579,In_1581);
or U1580 (N_1580,In_1697,In_2923);
xnor U1581 (N_1581,In_1488,In_2388);
or U1582 (N_1582,In_374,In_2562);
xnor U1583 (N_1583,In_2248,In_1237);
xor U1584 (N_1584,In_1708,In_2839);
nor U1585 (N_1585,In_1223,In_989);
and U1586 (N_1586,In_1264,In_2575);
xor U1587 (N_1587,In_732,In_386);
nor U1588 (N_1588,In_1886,In_190);
xor U1589 (N_1589,In_2810,In_929);
or U1590 (N_1590,In_2206,In_2444);
nor U1591 (N_1591,In_2413,In_1864);
nand U1592 (N_1592,In_2512,In_2151);
and U1593 (N_1593,In_374,In_158);
nand U1594 (N_1594,In_41,In_963);
xnor U1595 (N_1595,In_2718,In_1370);
or U1596 (N_1596,In_1350,In_526);
nand U1597 (N_1597,In_1538,In_2411);
nor U1598 (N_1598,In_494,In_1481);
nand U1599 (N_1599,In_1746,In_2305);
and U1600 (N_1600,In_605,In_2185);
and U1601 (N_1601,In_2960,In_197);
or U1602 (N_1602,In_2585,In_631);
nor U1603 (N_1603,In_1068,In_1667);
or U1604 (N_1604,In_294,In_1173);
or U1605 (N_1605,In_1288,In_2361);
and U1606 (N_1606,In_569,In_2970);
xor U1607 (N_1607,In_2812,In_693);
nand U1608 (N_1608,In_5,In_2812);
xnor U1609 (N_1609,In_865,In_1773);
and U1610 (N_1610,In_479,In_1231);
xor U1611 (N_1611,In_1875,In_808);
nor U1612 (N_1612,In_1959,In_59);
and U1613 (N_1613,In_1856,In_1456);
nand U1614 (N_1614,In_1252,In_1337);
nand U1615 (N_1615,In_511,In_1243);
or U1616 (N_1616,In_2761,In_1291);
and U1617 (N_1617,In_2384,In_1355);
or U1618 (N_1618,In_1901,In_1804);
nor U1619 (N_1619,In_691,In_2880);
nand U1620 (N_1620,In_366,In_480);
nand U1621 (N_1621,In_2998,In_1065);
and U1622 (N_1622,In_65,In_1083);
or U1623 (N_1623,In_388,In_1597);
and U1624 (N_1624,In_2688,In_543);
xnor U1625 (N_1625,In_1239,In_2308);
xor U1626 (N_1626,In_624,In_235);
nor U1627 (N_1627,In_1757,In_928);
or U1628 (N_1628,In_1429,In_1291);
xor U1629 (N_1629,In_494,In_352);
xnor U1630 (N_1630,In_2389,In_2805);
nor U1631 (N_1631,In_628,In_336);
nor U1632 (N_1632,In_1739,In_378);
or U1633 (N_1633,In_341,In_1855);
xnor U1634 (N_1634,In_1004,In_2139);
nand U1635 (N_1635,In_2930,In_2123);
or U1636 (N_1636,In_1163,In_481);
nand U1637 (N_1637,In_122,In_895);
or U1638 (N_1638,In_2138,In_528);
and U1639 (N_1639,In_2904,In_2983);
nor U1640 (N_1640,In_2637,In_1991);
nor U1641 (N_1641,In_385,In_2145);
or U1642 (N_1642,In_2669,In_2093);
xnor U1643 (N_1643,In_1729,In_2604);
or U1644 (N_1644,In_1498,In_2538);
nor U1645 (N_1645,In_1118,In_2182);
nor U1646 (N_1646,In_652,In_122);
and U1647 (N_1647,In_1961,In_2842);
nand U1648 (N_1648,In_494,In_1936);
or U1649 (N_1649,In_1765,In_864);
and U1650 (N_1650,In_1785,In_790);
nand U1651 (N_1651,In_185,In_1770);
and U1652 (N_1652,In_1827,In_2277);
nor U1653 (N_1653,In_2971,In_885);
or U1654 (N_1654,In_2787,In_144);
and U1655 (N_1655,In_1542,In_801);
nand U1656 (N_1656,In_1400,In_2407);
or U1657 (N_1657,In_482,In_2376);
or U1658 (N_1658,In_2644,In_827);
xnor U1659 (N_1659,In_67,In_1914);
nand U1660 (N_1660,In_1081,In_1052);
xor U1661 (N_1661,In_2011,In_929);
xor U1662 (N_1662,In_359,In_1064);
nand U1663 (N_1663,In_1139,In_1158);
nor U1664 (N_1664,In_2953,In_357);
or U1665 (N_1665,In_1191,In_863);
and U1666 (N_1666,In_2262,In_2314);
nand U1667 (N_1667,In_2036,In_2348);
nor U1668 (N_1668,In_1134,In_176);
and U1669 (N_1669,In_1629,In_1059);
nand U1670 (N_1670,In_2995,In_919);
or U1671 (N_1671,In_969,In_2630);
xnor U1672 (N_1672,In_1786,In_2947);
nand U1673 (N_1673,In_926,In_2656);
xor U1674 (N_1674,In_1649,In_729);
and U1675 (N_1675,In_648,In_2472);
or U1676 (N_1676,In_185,In_1207);
nor U1677 (N_1677,In_2691,In_868);
or U1678 (N_1678,In_2233,In_1007);
and U1679 (N_1679,In_1269,In_2615);
or U1680 (N_1680,In_1571,In_1068);
and U1681 (N_1681,In_21,In_2000);
or U1682 (N_1682,In_1221,In_2934);
or U1683 (N_1683,In_896,In_2841);
nor U1684 (N_1684,In_2100,In_2509);
and U1685 (N_1685,In_1946,In_506);
xor U1686 (N_1686,In_1445,In_1913);
nor U1687 (N_1687,In_172,In_1787);
xor U1688 (N_1688,In_1385,In_2596);
and U1689 (N_1689,In_79,In_1945);
nand U1690 (N_1690,In_1674,In_1);
nor U1691 (N_1691,In_2406,In_475);
nor U1692 (N_1692,In_1824,In_479);
nor U1693 (N_1693,In_2668,In_985);
or U1694 (N_1694,In_1983,In_1640);
nor U1695 (N_1695,In_932,In_1421);
nand U1696 (N_1696,In_95,In_2622);
nor U1697 (N_1697,In_243,In_530);
nand U1698 (N_1698,In_1594,In_1783);
nand U1699 (N_1699,In_1128,In_406);
and U1700 (N_1700,In_2166,In_1016);
and U1701 (N_1701,In_587,In_10);
nor U1702 (N_1702,In_2796,In_2284);
and U1703 (N_1703,In_2454,In_371);
xor U1704 (N_1704,In_2227,In_800);
nand U1705 (N_1705,In_2572,In_284);
and U1706 (N_1706,In_1725,In_2396);
or U1707 (N_1707,In_1226,In_2203);
and U1708 (N_1708,In_2884,In_1151);
xnor U1709 (N_1709,In_1372,In_944);
or U1710 (N_1710,In_1979,In_1510);
or U1711 (N_1711,In_1930,In_2035);
and U1712 (N_1712,In_44,In_1014);
nor U1713 (N_1713,In_1263,In_844);
nand U1714 (N_1714,In_2548,In_1095);
and U1715 (N_1715,In_1106,In_1081);
and U1716 (N_1716,In_236,In_1853);
nor U1717 (N_1717,In_239,In_1841);
or U1718 (N_1718,In_2494,In_1096);
nor U1719 (N_1719,In_647,In_2084);
or U1720 (N_1720,In_1519,In_800);
and U1721 (N_1721,In_687,In_1377);
or U1722 (N_1722,In_2513,In_559);
xnor U1723 (N_1723,In_1114,In_2590);
and U1724 (N_1724,In_392,In_1189);
nor U1725 (N_1725,In_2042,In_954);
nor U1726 (N_1726,In_1559,In_1452);
or U1727 (N_1727,In_2669,In_1749);
nand U1728 (N_1728,In_2113,In_2349);
or U1729 (N_1729,In_2208,In_1210);
or U1730 (N_1730,In_2568,In_452);
and U1731 (N_1731,In_1305,In_609);
xnor U1732 (N_1732,In_1963,In_2867);
and U1733 (N_1733,In_1920,In_336);
nor U1734 (N_1734,In_2355,In_2221);
xor U1735 (N_1735,In_2665,In_1862);
nand U1736 (N_1736,In_2330,In_932);
and U1737 (N_1737,In_711,In_1515);
nor U1738 (N_1738,In_603,In_445);
and U1739 (N_1739,In_1920,In_1244);
nor U1740 (N_1740,In_1618,In_1854);
and U1741 (N_1741,In_61,In_1702);
nor U1742 (N_1742,In_1733,In_1716);
and U1743 (N_1743,In_1564,In_2819);
nand U1744 (N_1744,In_989,In_33);
or U1745 (N_1745,In_1879,In_383);
and U1746 (N_1746,In_1624,In_1003);
or U1747 (N_1747,In_1009,In_2608);
xor U1748 (N_1748,In_363,In_404);
nand U1749 (N_1749,In_221,In_1201);
nor U1750 (N_1750,In_374,In_978);
nor U1751 (N_1751,In_1619,In_2872);
nor U1752 (N_1752,In_270,In_946);
xnor U1753 (N_1753,In_2944,In_1573);
nand U1754 (N_1754,In_1962,In_1856);
nor U1755 (N_1755,In_437,In_1383);
and U1756 (N_1756,In_2554,In_2103);
or U1757 (N_1757,In_542,In_2097);
or U1758 (N_1758,In_1190,In_1969);
xnor U1759 (N_1759,In_1317,In_2208);
nand U1760 (N_1760,In_2760,In_2669);
xnor U1761 (N_1761,In_1175,In_1092);
nor U1762 (N_1762,In_338,In_2159);
or U1763 (N_1763,In_592,In_589);
nor U1764 (N_1764,In_1024,In_1502);
nand U1765 (N_1765,In_2081,In_565);
nand U1766 (N_1766,In_491,In_2464);
nand U1767 (N_1767,In_2946,In_1701);
nand U1768 (N_1768,In_1329,In_387);
or U1769 (N_1769,In_1329,In_1486);
xnor U1770 (N_1770,In_383,In_997);
or U1771 (N_1771,In_1220,In_102);
and U1772 (N_1772,In_1290,In_138);
xor U1773 (N_1773,In_2854,In_2922);
nand U1774 (N_1774,In_104,In_1086);
nand U1775 (N_1775,In_2321,In_1893);
nor U1776 (N_1776,In_748,In_2651);
and U1777 (N_1777,In_1829,In_1317);
xnor U1778 (N_1778,In_382,In_1955);
or U1779 (N_1779,In_1504,In_692);
or U1780 (N_1780,In_702,In_2106);
nand U1781 (N_1781,In_1582,In_2800);
nand U1782 (N_1782,In_2388,In_2565);
nor U1783 (N_1783,In_2637,In_1393);
xnor U1784 (N_1784,In_492,In_48);
xnor U1785 (N_1785,In_794,In_31);
xnor U1786 (N_1786,In_1456,In_2898);
nor U1787 (N_1787,In_743,In_2500);
and U1788 (N_1788,In_1568,In_1185);
xor U1789 (N_1789,In_2056,In_2399);
or U1790 (N_1790,In_2014,In_1281);
xnor U1791 (N_1791,In_397,In_1349);
nand U1792 (N_1792,In_858,In_1380);
nand U1793 (N_1793,In_1476,In_416);
nand U1794 (N_1794,In_84,In_1638);
and U1795 (N_1795,In_2954,In_2017);
or U1796 (N_1796,In_247,In_1378);
xor U1797 (N_1797,In_1694,In_2598);
or U1798 (N_1798,In_581,In_457);
nand U1799 (N_1799,In_1641,In_1544);
nor U1800 (N_1800,In_1468,In_1690);
nand U1801 (N_1801,In_257,In_2197);
or U1802 (N_1802,In_2102,In_2397);
and U1803 (N_1803,In_472,In_2811);
or U1804 (N_1804,In_130,In_1519);
or U1805 (N_1805,In_973,In_1433);
xor U1806 (N_1806,In_789,In_1679);
and U1807 (N_1807,In_2906,In_2908);
and U1808 (N_1808,In_738,In_1031);
and U1809 (N_1809,In_1119,In_41);
and U1810 (N_1810,In_2742,In_1881);
and U1811 (N_1811,In_2346,In_2818);
or U1812 (N_1812,In_2799,In_1324);
nor U1813 (N_1813,In_1929,In_377);
xnor U1814 (N_1814,In_2257,In_2040);
or U1815 (N_1815,In_993,In_1697);
nor U1816 (N_1816,In_2650,In_660);
nor U1817 (N_1817,In_544,In_1731);
or U1818 (N_1818,In_2122,In_938);
and U1819 (N_1819,In_922,In_162);
and U1820 (N_1820,In_1871,In_1317);
nor U1821 (N_1821,In_1479,In_924);
nor U1822 (N_1822,In_2873,In_63);
and U1823 (N_1823,In_2726,In_1639);
nand U1824 (N_1824,In_2085,In_425);
or U1825 (N_1825,In_2280,In_1814);
or U1826 (N_1826,In_1770,In_1731);
nor U1827 (N_1827,In_918,In_2120);
nand U1828 (N_1828,In_2800,In_2382);
and U1829 (N_1829,In_2028,In_2951);
nor U1830 (N_1830,In_184,In_312);
nor U1831 (N_1831,In_702,In_885);
nor U1832 (N_1832,In_1588,In_2818);
or U1833 (N_1833,In_1788,In_2080);
nor U1834 (N_1834,In_2877,In_1972);
or U1835 (N_1835,In_966,In_583);
and U1836 (N_1836,In_1425,In_82);
xor U1837 (N_1837,In_2764,In_323);
and U1838 (N_1838,In_794,In_1809);
xnor U1839 (N_1839,In_197,In_287);
and U1840 (N_1840,In_1010,In_2418);
nand U1841 (N_1841,In_2232,In_122);
xnor U1842 (N_1842,In_2862,In_2656);
nand U1843 (N_1843,In_1540,In_1408);
and U1844 (N_1844,In_2502,In_1794);
nor U1845 (N_1845,In_1769,In_2144);
xnor U1846 (N_1846,In_135,In_332);
xnor U1847 (N_1847,In_1351,In_2004);
nand U1848 (N_1848,In_119,In_51);
nor U1849 (N_1849,In_1427,In_956);
nor U1850 (N_1850,In_1808,In_1994);
nand U1851 (N_1851,In_2965,In_710);
or U1852 (N_1852,In_2889,In_421);
nand U1853 (N_1853,In_621,In_70);
nor U1854 (N_1854,In_84,In_2910);
nor U1855 (N_1855,In_2290,In_1688);
and U1856 (N_1856,In_1697,In_2312);
or U1857 (N_1857,In_2525,In_1510);
nor U1858 (N_1858,In_203,In_232);
xor U1859 (N_1859,In_1713,In_2393);
or U1860 (N_1860,In_1653,In_2548);
and U1861 (N_1861,In_2924,In_2087);
nor U1862 (N_1862,In_1031,In_2169);
and U1863 (N_1863,In_99,In_882);
nand U1864 (N_1864,In_2961,In_882);
nand U1865 (N_1865,In_379,In_1775);
nor U1866 (N_1866,In_2807,In_2942);
nor U1867 (N_1867,In_835,In_587);
or U1868 (N_1868,In_898,In_836);
nand U1869 (N_1869,In_806,In_78);
xor U1870 (N_1870,In_1331,In_1281);
xnor U1871 (N_1871,In_511,In_1372);
xor U1872 (N_1872,In_1078,In_537);
xor U1873 (N_1873,In_2932,In_866);
and U1874 (N_1874,In_2239,In_163);
nand U1875 (N_1875,In_387,In_1547);
or U1876 (N_1876,In_995,In_873);
xnor U1877 (N_1877,In_2153,In_2083);
nand U1878 (N_1878,In_2109,In_1794);
and U1879 (N_1879,In_2423,In_678);
or U1880 (N_1880,In_1008,In_2873);
or U1881 (N_1881,In_1364,In_2382);
nor U1882 (N_1882,In_802,In_602);
xnor U1883 (N_1883,In_241,In_1808);
xor U1884 (N_1884,In_607,In_875);
and U1885 (N_1885,In_1794,In_254);
or U1886 (N_1886,In_819,In_2249);
and U1887 (N_1887,In_1979,In_549);
and U1888 (N_1888,In_2740,In_1015);
xor U1889 (N_1889,In_1610,In_2267);
xor U1890 (N_1890,In_1427,In_1638);
xor U1891 (N_1891,In_2281,In_963);
nor U1892 (N_1892,In_2405,In_1823);
nand U1893 (N_1893,In_2130,In_2219);
and U1894 (N_1894,In_2459,In_2014);
xor U1895 (N_1895,In_530,In_743);
nor U1896 (N_1896,In_2721,In_2221);
nor U1897 (N_1897,In_1894,In_2870);
nand U1898 (N_1898,In_2353,In_1829);
and U1899 (N_1899,In_888,In_884);
and U1900 (N_1900,In_2340,In_920);
nor U1901 (N_1901,In_1311,In_895);
nand U1902 (N_1902,In_1718,In_1737);
nand U1903 (N_1903,In_2822,In_1836);
or U1904 (N_1904,In_2350,In_1435);
nor U1905 (N_1905,In_2802,In_1060);
xor U1906 (N_1906,In_2928,In_629);
nor U1907 (N_1907,In_283,In_1567);
xnor U1908 (N_1908,In_1926,In_1505);
xor U1909 (N_1909,In_1109,In_451);
or U1910 (N_1910,In_1814,In_2072);
nor U1911 (N_1911,In_1455,In_229);
and U1912 (N_1912,In_611,In_1010);
nand U1913 (N_1913,In_208,In_2421);
nor U1914 (N_1914,In_804,In_774);
nand U1915 (N_1915,In_1741,In_1544);
and U1916 (N_1916,In_507,In_1248);
or U1917 (N_1917,In_2160,In_2269);
nor U1918 (N_1918,In_437,In_237);
or U1919 (N_1919,In_516,In_2728);
nor U1920 (N_1920,In_592,In_1245);
and U1921 (N_1921,In_1971,In_2828);
nor U1922 (N_1922,In_1158,In_465);
or U1923 (N_1923,In_1267,In_1712);
xnor U1924 (N_1924,In_1597,In_1853);
nand U1925 (N_1925,In_2750,In_1794);
xnor U1926 (N_1926,In_2937,In_70);
xor U1927 (N_1927,In_2446,In_942);
nand U1928 (N_1928,In_2154,In_709);
and U1929 (N_1929,In_2233,In_1933);
and U1930 (N_1930,In_378,In_851);
nor U1931 (N_1931,In_760,In_288);
nand U1932 (N_1932,In_337,In_1395);
or U1933 (N_1933,In_351,In_1317);
or U1934 (N_1934,In_819,In_968);
nor U1935 (N_1935,In_271,In_1345);
and U1936 (N_1936,In_1834,In_748);
xnor U1937 (N_1937,In_2442,In_2917);
or U1938 (N_1938,In_1459,In_1616);
and U1939 (N_1939,In_154,In_2948);
or U1940 (N_1940,In_2195,In_2119);
nor U1941 (N_1941,In_832,In_570);
nor U1942 (N_1942,In_362,In_2117);
and U1943 (N_1943,In_2329,In_2600);
or U1944 (N_1944,In_2255,In_916);
and U1945 (N_1945,In_1469,In_104);
xor U1946 (N_1946,In_596,In_296);
nand U1947 (N_1947,In_1747,In_1516);
nor U1948 (N_1948,In_1052,In_1145);
and U1949 (N_1949,In_2772,In_2998);
or U1950 (N_1950,In_1973,In_995);
and U1951 (N_1951,In_2179,In_1114);
and U1952 (N_1952,In_583,In_2288);
xor U1953 (N_1953,In_391,In_913);
nand U1954 (N_1954,In_839,In_2907);
and U1955 (N_1955,In_2891,In_1084);
xnor U1956 (N_1956,In_375,In_1906);
and U1957 (N_1957,In_2468,In_1279);
nand U1958 (N_1958,In_2612,In_760);
and U1959 (N_1959,In_1217,In_1970);
or U1960 (N_1960,In_1354,In_644);
xnor U1961 (N_1961,In_2171,In_1856);
nor U1962 (N_1962,In_837,In_843);
nand U1963 (N_1963,In_1884,In_2247);
nor U1964 (N_1964,In_775,In_1558);
and U1965 (N_1965,In_18,In_2988);
xnor U1966 (N_1966,In_291,In_2452);
nor U1967 (N_1967,In_816,In_2659);
nor U1968 (N_1968,In_2876,In_518);
or U1969 (N_1969,In_2861,In_2841);
or U1970 (N_1970,In_1556,In_1634);
or U1971 (N_1971,In_1743,In_0);
and U1972 (N_1972,In_2387,In_1831);
nand U1973 (N_1973,In_945,In_1759);
and U1974 (N_1974,In_639,In_334);
and U1975 (N_1975,In_1878,In_1434);
xor U1976 (N_1976,In_1137,In_2448);
or U1977 (N_1977,In_347,In_2225);
nor U1978 (N_1978,In_1776,In_1880);
or U1979 (N_1979,In_1699,In_1553);
xor U1980 (N_1980,In_1217,In_2465);
or U1981 (N_1981,In_2181,In_156);
xor U1982 (N_1982,In_297,In_1675);
nor U1983 (N_1983,In_2115,In_890);
or U1984 (N_1984,In_2126,In_786);
nor U1985 (N_1985,In_1697,In_1753);
and U1986 (N_1986,In_1153,In_1044);
and U1987 (N_1987,In_2144,In_2417);
or U1988 (N_1988,In_2953,In_775);
nor U1989 (N_1989,In_2234,In_506);
nand U1990 (N_1990,In_2268,In_2307);
nand U1991 (N_1991,In_1655,In_844);
nor U1992 (N_1992,In_2701,In_1049);
xnor U1993 (N_1993,In_641,In_599);
or U1994 (N_1994,In_2635,In_454);
and U1995 (N_1995,In_1106,In_1520);
nand U1996 (N_1996,In_1368,In_2619);
nor U1997 (N_1997,In_2096,In_773);
nor U1998 (N_1998,In_61,In_2516);
xor U1999 (N_1999,In_668,In_2158);
xor U2000 (N_2000,In_2627,In_202);
xnor U2001 (N_2001,In_2114,In_694);
nor U2002 (N_2002,In_2111,In_461);
nand U2003 (N_2003,In_1944,In_2025);
nor U2004 (N_2004,In_2883,In_1453);
xnor U2005 (N_2005,In_1126,In_602);
xnor U2006 (N_2006,In_2537,In_2195);
and U2007 (N_2007,In_1656,In_2283);
nand U2008 (N_2008,In_2622,In_1701);
xor U2009 (N_2009,In_1081,In_1643);
or U2010 (N_2010,In_1438,In_250);
xor U2011 (N_2011,In_1248,In_252);
nand U2012 (N_2012,In_1523,In_1001);
xnor U2013 (N_2013,In_252,In_1255);
xnor U2014 (N_2014,In_799,In_235);
or U2015 (N_2015,In_1598,In_1930);
nor U2016 (N_2016,In_2863,In_2658);
or U2017 (N_2017,In_1508,In_1157);
nor U2018 (N_2018,In_1942,In_2844);
or U2019 (N_2019,In_491,In_1260);
and U2020 (N_2020,In_2511,In_2146);
nor U2021 (N_2021,In_1758,In_1657);
nand U2022 (N_2022,In_1858,In_1608);
xnor U2023 (N_2023,In_2177,In_1712);
or U2024 (N_2024,In_2150,In_2480);
nand U2025 (N_2025,In_1183,In_2229);
xnor U2026 (N_2026,In_2981,In_2363);
xor U2027 (N_2027,In_2661,In_100);
or U2028 (N_2028,In_2291,In_1793);
xnor U2029 (N_2029,In_1884,In_149);
nor U2030 (N_2030,In_1437,In_1756);
nand U2031 (N_2031,In_2726,In_891);
nand U2032 (N_2032,In_1255,In_440);
nor U2033 (N_2033,In_754,In_2116);
xnor U2034 (N_2034,In_2311,In_1454);
and U2035 (N_2035,In_2996,In_2987);
and U2036 (N_2036,In_829,In_1159);
and U2037 (N_2037,In_855,In_1289);
or U2038 (N_2038,In_1654,In_122);
nand U2039 (N_2039,In_511,In_704);
or U2040 (N_2040,In_879,In_1780);
xor U2041 (N_2041,In_924,In_2153);
and U2042 (N_2042,In_208,In_1673);
and U2043 (N_2043,In_147,In_993);
nand U2044 (N_2044,In_2334,In_2109);
nand U2045 (N_2045,In_2766,In_621);
or U2046 (N_2046,In_964,In_2303);
or U2047 (N_2047,In_2482,In_232);
and U2048 (N_2048,In_394,In_2573);
and U2049 (N_2049,In_2337,In_2077);
or U2050 (N_2050,In_1051,In_1352);
xor U2051 (N_2051,In_687,In_547);
nand U2052 (N_2052,In_338,In_1857);
xor U2053 (N_2053,In_249,In_2317);
or U2054 (N_2054,In_2251,In_2565);
or U2055 (N_2055,In_1042,In_2127);
nor U2056 (N_2056,In_1247,In_439);
nand U2057 (N_2057,In_1470,In_1486);
xnor U2058 (N_2058,In_568,In_93);
and U2059 (N_2059,In_1778,In_294);
xor U2060 (N_2060,In_124,In_2833);
and U2061 (N_2061,In_1896,In_43);
nand U2062 (N_2062,In_48,In_2896);
nor U2063 (N_2063,In_728,In_614);
and U2064 (N_2064,In_1312,In_966);
nor U2065 (N_2065,In_1596,In_2354);
nor U2066 (N_2066,In_2070,In_2559);
nand U2067 (N_2067,In_2092,In_1640);
and U2068 (N_2068,In_2055,In_2306);
and U2069 (N_2069,In_97,In_2340);
and U2070 (N_2070,In_2405,In_2116);
and U2071 (N_2071,In_2841,In_1098);
and U2072 (N_2072,In_47,In_297);
or U2073 (N_2073,In_837,In_2781);
or U2074 (N_2074,In_461,In_349);
xnor U2075 (N_2075,In_2535,In_1403);
or U2076 (N_2076,In_2357,In_525);
and U2077 (N_2077,In_17,In_421);
and U2078 (N_2078,In_1752,In_1798);
and U2079 (N_2079,In_1374,In_2000);
nor U2080 (N_2080,In_1048,In_1157);
nand U2081 (N_2081,In_465,In_496);
and U2082 (N_2082,In_2296,In_720);
or U2083 (N_2083,In_2454,In_2479);
nand U2084 (N_2084,In_2791,In_1922);
xor U2085 (N_2085,In_2798,In_2278);
and U2086 (N_2086,In_1420,In_262);
xor U2087 (N_2087,In_950,In_870);
and U2088 (N_2088,In_2188,In_990);
and U2089 (N_2089,In_980,In_1261);
and U2090 (N_2090,In_1591,In_951);
or U2091 (N_2091,In_2613,In_2841);
nor U2092 (N_2092,In_546,In_2925);
xor U2093 (N_2093,In_2683,In_1649);
xor U2094 (N_2094,In_1710,In_1898);
and U2095 (N_2095,In_2376,In_521);
xnor U2096 (N_2096,In_338,In_1580);
and U2097 (N_2097,In_53,In_2520);
nor U2098 (N_2098,In_105,In_2815);
nand U2099 (N_2099,In_2901,In_1849);
nor U2100 (N_2100,In_1833,In_1407);
or U2101 (N_2101,In_1654,In_1697);
nand U2102 (N_2102,In_2570,In_406);
and U2103 (N_2103,In_761,In_2433);
or U2104 (N_2104,In_1189,In_999);
and U2105 (N_2105,In_1438,In_474);
or U2106 (N_2106,In_949,In_1719);
xor U2107 (N_2107,In_983,In_2595);
or U2108 (N_2108,In_794,In_67);
nor U2109 (N_2109,In_391,In_1713);
nor U2110 (N_2110,In_447,In_729);
or U2111 (N_2111,In_2715,In_1226);
nand U2112 (N_2112,In_2000,In_2981);
xor U2113 (N_2113,In_2243,In_2908);
xor U2114 (N_2114,In_261,In_104);
nor U2115 (N_2115,In_225,In_977);
or U2116 (N_2116,In_2149,In_1806);
xnor U2117 (N_2117,In_598,In_892);
or U2118 (N_2118,In_26,In_1492);
nand U2119 (N_2119,In_1843,In_576);
or U2120 (N_2120,In_924,In_547);
and U2121 (N_2121,In_133,In_1649);
and U2122 (N_2122,In_1761,In_1255);
xnor U2123 (N_2123,In_1867,In_2864);
or U2124 (N_2124,In_218,In_2338);
or U2125 (N_2125,In_602,In_2791);
or U2126 (N_2126,In_414,In_222);
or U2127 (N_2127,In_2689,In_1161);
and U2128 (N_2128,In_1711,In_2256);
or U2129 (N_2129,In_2147,In_363);
xnor U2130 (N_2130,In_2564,In_221);
and U2131 (N_2131,In_1295,In_1904);
and U2132 (N_2132,In_50,In_2744);
or U2133 (N_2133,In_2655,In_2329);
and U2134 (N_2134,In_2253,In_793);
and U2135 (N_2135,In_678,In_899);
nor U2136 (N_2136,In_2857,In_835);
and U2137 (N_2137,In_1884,In_1058);
and U2138 (N_2138,In_715,In_158);
xor U2139 (N_2139,In_209,In_2744);
or U2140 (N_2140,In_1752,In_828);
nand U2141 (N_2141,In_1751,In_2447);
xnor U2142 (N_2142,In_2837,In_2171);
and U2143 (N_2143,In_2883,In_292);
or U2144 (N_2144,In_1280,In_1392);
or U2145 (N_2145,In_1442,In_8);
and U2146 (N_2146,In_2765,In_1643);
and U2147 (N_2147,In_1750,In_1940);
xor U2148 (N_2148,In_210,In_764);
and U2149 (N_2149,In_2667,In_2198);
nor U2150 (N_2150,In_1995,In_592);
or U2151 (N_2151,In_2696,In_428);
or U2152 (N_2152,In_2712,In_2156);
and U2153 (N_2153,In_2435,In_2824);
nand U2154 (N_2154,In_1131,In_901);
nor U2155 (N_2155,In_1435,In_2934);
xnor U2156 (N_2156,In_2508,In_1777);
and U2157 (N_2157,In_666,In_500);
xor U2158 (N_2158,In_311,In_2741);
or U2159 (N_2159,In_1994,In_357);
nor U2160 (N_2160,In_683,In_757);
nor U2161 (N_2161,In_718,In_227);
or U2162 (N_2162,In_1972,In_2733);
nand U2163 (N_2163,In_1290,In_1979);
nand U2164 (N_2164,In_2449,In_1917);
xnor U2165 (N_2165,In_2857,In_2018);
nor U2166 (N_2166,In_2853,In_2899);
and U2167 (N_2167,In_1074,In_614);
and U2168 (N_2168,In_2146,In_2666);
nand U2169 (N_2169,In_2976,In_2721);
nand U2170 (N_2170,In_189,In_996);
nor U2171 (N_2171,In_439,In_2338);
nand U2172 (N_2172,In_2987,In_1093);
nor U2173 (N_2173,In_523,In_1962);
or U2174 (N_2174,In_2497,In_2165);
nor U2175 (N_2175,In_2191,In_2816);
xnor U2176 (N_2176,In_1025,In_738);
xor U2177 (N_2177,In_1480,In_2880);
or U2178 (N_2178,In_1065,In_1229);
xnor U2179 (N_2179,In_2905,In_1289);
nor U2180 (N_2180,In_754,In_2680);
nor U2181 (N_2181,In_2632,In_573);
or U2182 (N_2182,In_631,In_2435);
nor U2183 (N_2183,In_477,In_684);
nand U2184 (N_2184,In_2526,In_1813);
nor U2185 (N_2185,In_711,In_1112);
nor U2186 (N_2186,In_413,In_1134);
and U2187 (N_2187,In_2235,In_206);
nor U2188 (N_2188,In_2937,In_2075);
and U2189 (N_2189,In_537,In_1946);
or U2190 (N_2190,In_2907,In_1174);
and U2191 (N_2191,In_1545,In_2998);
nand U2192 (N_2192,In_1100,In_2696);
nor U2193 (N_2193,In_1201,In_434);
and U2194 (N_2194,In_1631,In_1491);
nor U2195 (N_2195,In_110,In_1587);
and U2196 (N_2196,In_1609,In_2533);
xnor U2197 (N_2197,In_2390,In_2241);
nand U2198 (N_2198,In_2233,In_1798);
xor U2199 (N_2199,In_2334,In_608);
and U2200 (N_2200,In_564,In_334);
nor U2201 (N_2201,In_1666,In_2865);
nand U2202 (N_2202,In_1828,In_1301);
nor U2203 (N_2203,In_2295,In_2046);
or U2204 (N_2204,In_2830,In_2824);
or U2205 (N_2205,In_1109,In_1355);
xor U2206 (N_2206,In_2770,In_660);
nand U2207 (N_2207,In_2999,In_2352);
nand U2208 (N_2208,In_1142,In_2589);
nor U2209 (N_2209,In_2749,In_2081);
nor U2210 (N_2210,In_1163,In_813);
xnor U2211 (N_2211,In_1221,In_264);
nor U2212 (N_2212,In_2794,In_1192);
xnor U2213 (N_2213,In_2766,In_2384);
xor U2214 (N_2214,In_1284,In_2579);
or U2215 (N_2215,In_843,In_2393);
and U2216 (N_2216,In_1373,In_2567);
nand U2217 (N_2217,In_2885,In_1338);
nor U2218 (N_2218,In_2764,In_476);
xnor U2219 (N_2219,In_1753,In_2909);
nand U2220 (N_2220,In_2120,In_1300);
xor U2221 (N_2221,In_1611,In_678);
xor U2222 (N_2222,In_892,In_2635);
nand U2223 (N_2223,In_1083,In_1338);
xor U2224 (N_2224,In_1264,In_26);
nor U2225 (N_2225,In_2446,In_646);
or U2226 (N_2226,In_2509,In_799);
nor U2227 (N_2227,In_339,In_110);
and U2228 (N_2228,In_142,In_2556);
nand U2229 (N_2229,In_484,In_78);
xnor U2230 (N_2230,In_1050,In_1125);
and U2231 (N_2231,In_2106,In_1064);
nand U2232 (N_2232,In_2266,In_817);
nor U2233 (N_2233,In_672,In_552);
or U2234 (N_2234,In_1311,In_553);
and U2235 (N_2235,In_509,In_356);
nor U2236 (N_2236,In_99,In_2614);
nand U2237 (N_2237,In_2276,In_1083);
nand U2238 (N_2238,In_2401,In_2071);
nor U2239 (N_2239,In_301,In_2002);
nand U2240 (N_2240,In_882,In_2029);
xor U2241 (N_2241,In_2590,In_536);
nand U2242 (N_2242,In_1767,In_2667);
nand U2243 (N_2243,In_2594,In_1837);
xnor U2244 (N_2244,In_2551,In_2268);
nor U2245 (N_2245,In_1185,In_220);
and U2246 (N_2246,In_853,In_884);
and U2247 (N_2247,In_832,In_463);
nor U2248 (N_2248,In_401,In_2727);
and U2249 (N_2249,In_2636,In_704);
and U2250 (N_2250,In_1726,In_819);
or U2251 (N_2251,In_1604,In_2597);
and U2252 (N_2252,In_2797,In_881);
and U2253 (N_2253,In_1456,In_1039);
nand U2254 (N_2254,In_2054,In_1286);
or U2255 (N_2255,In_2758,In_350);
nor U2256 (N_2256,In_1744,In_923);
and U2257 (N_2257,In_860,In_2979);
or U2258 (N_2258,In_223,In_2054);
nand U2259 (N_2259,In_1906,In_2381);
and U2260 (N_2260,In_929,In_2248);
xnor U2261 (N_2261,In_2548,In_2199);
xor U2262 (N_2262,In_2728,In_930);
xor U2263 (N_2263,In_1746,In_2110);
xnor U2264 (N_2264,In_1672,In_2980);
or U2265 (N_2265,In_722,In_2193);
or U2266 (N_2266,In_2354,In_613);
nand U2267 (N_2267,In_1328,In_2268);
or U2268 (N_2268,In_2223,In_1656);
and U2269 (N_2269,In_1502,In_2280);
nand U2270 (N_2270,In_633,In_2946);
nor U2271 (N_2271,In_2066,In_1825);
xor U2272 (N_2272,In_1138,In_1583);
nand U2273 (N_2273,In_326,In_868);
nand U2274 (N_2274,In_1792,In_2350);
or U2275 (N_2275,In_2362,In_2368);
or U2276 (N_2276,In_2138,In_2017);
xnor U2277 (N_2277,In_818,In_2851);
xor U2278 (N_2278,In_2109,In_523);
nor U2279 (N_2279,In_658,In_2013);
nor U2280 (N_2280,In_1023,In_1001);
and U2281 (N_2281,In_1818,In_609);
xor U2282 (N_2282,In_1518,In_608);
xnor U2283 (N_2283,In_2405,In_1818);
nor U2284 (N_2284,In_1519,In_1797);
nor U2285 (N_2285,In_2668,In_444);
or U2286 (N_2286,In_2168,In_865);
xor U2287 (N_2287,In_2319,In_2233);
xor U2288 (N_2288,In_2147,In_338);
nand U2289 (N_2289,In_914,In_2446);
nand U2290 (N_2290,In_839,In_198);
xnor U2291 (N_2291,In_2488,In_2886);
nand U2292 (N_2292,In_471,In_2876);
nand U2293 (N_2293,In_1563,In_998);
and U2294 (N_2294,In_2690,In_1664);
and U2295 (N_2295,In_966,In_2392);
and U2296 (N_2296,In_2772,In_2512);
xnor U2297 (N_2297,In_1059,In_2761);
xnor U2298 (N_2298,In_1727,In_323);
and U2299 (N_2299,In_1653,In_2346);
xor U2300 (N_2300,In_871,In_215);
and U2301 (N_2301,In_1589,In_1253);
nand U2302 (N_2302,In_2485,In_2646);
and U2303 (N_2303,In_2378,In_2592);
or U2304 (N_2304,In_2755,In_1819);
and U2305 (N_2305,In_1683,In_1697);
nand U2306 (N_2306,In_2427,In_603);
nor U2307 (N_2307,In_1745,In_2807);
nand U2308 (N_2308,In_1810,In_2023);
nor U2309 (N_2309,In_2394,In_1621);
and U2310 (N_2310,In_1664,In_1957);
nand U2311 (N_2311,In_2931,In_2418);
or U2312 (N_2312,In_78,In_232);
and U2313 (N_2313,In_1433,In_2990);
xnor U2314 (N_2314,In_686,In_451);
nand U2315 (N_2315,In_1932,In_1195);
nand U2316 (N_2316,In_2381,In_804);
or U2317 (N_2317,In_1616,In_549);
xnor U2318 (N_2318,In_217,In_954);
or U2319 (N_2319,In_2137,In_175);
or U2320 (N_2320,In_306,In_1164);
nor U2321 (N_2321,In_429,In_392);
or U2322 (N_2322,In_1543,In_1147);
or U2323 (N_2323,In_1349,In_2781);
xnor U2324 (N_2324,In_2182,In_2438);
nand U2325 (N_2325,In_332,In_2797);
and U2326 (N_2326,In_2374,In_1408);
nor U2327 (N_2327,In_742,In_1887);
nand U2328 (N_2328,In_2485,In_2860);
nor U2329 (N_2329,In_2568,In_354);
or U2330 (N_2330,In_417,In_387);
xnor U2331 (N_2331,In_1726,In_1748);
and U2332 (N_2332,In_128,In_148);
or U2333 (N_2333,In_2379,In_1289);
and U2334 (N_2334,In_786,In_1770);
and U2335 (N_2335,In_2344,In_1254);
and U2336 (N_2336,In_2992,In_329);
or U2337 (N_2337,In_2764,In_1111);
nor U2338 (N_2338,In_1988,In_894);
nand U2339 (N_2339,In_1111,In_2631);
nor U2340 (N_2340,In_1453,In_1510);
or U2341 (N_2341,In_2156,In_1413);
xor U2342 (N_2342,In_954,In_1539);
nand U2343 (N_2343,In_2234,In_1710);
nor U2344 (N_2344,In_2599,In_208);
xor U2345 (N_2345,In_2131,In_2755);
nor U2346 (N_2346,In_850,In_909);
nor U2347 (N_2347,In_1549,In_2114);
nand U2348 (N_2348,In_1706,In_1411);
nor U2349 (N_2349,In_1088,In_204);
or U2350 (N_2350,In_1402,In_32);
nor U2351 (N_2351,In_63,In_2058);
nor U2352 (N_2352,In_590,In_55);
nor U2353 (N_2353,In_2149,In_591);
nand U2354 (N_2354,In_2536,In_2187);
and U2355 (N_2355,In_2654,In_844);
and U2356 (N_2356,In_1656,In_848);
nand U2357 (N_2357,In_1984,In_2578);
xnor U2358 (N_2358,In_914,In_610);
nand U2359 (N_2359,In_1672,In_2892);
xnor U2360 (N_2360,In_819,In_2422);
or U2361 (N_2361,In_1134,In_2307);
xnor U2362 (N_2362,In_2641,In_2935);
or U2363 (N_2363,In_1168,In_1267);
xnor U2364 (N_2364,In_1381,In_980);
xor U2365 (N_2365,In_1902,In_1498);
and U2366 (N_2366,In_462,In_17);
nand U2367 (N_2367,In_932,In_1116);
xnor U2368 (N_2368,In_506,In_2456);
or U2369 (N_2369,In_2013,In_2009);
nor U2370 (N_2370,In_2553,In_327);
and U2371 (N_2371,In_904,In_2454);
xnor U2372 (N_2372,In_2094,In_87);
or U2373 (N_2373,In_83,In_174);
xnor U2374 (N_2374,In_1855,In_1980);
or U2375 (N_2375,In_129,In_2677);
or U2376 (N_2376,In_537,In_2215);
xnor U2377 (N_2377,In_2252,In_309);
and U2378 (N_2378,In_1414,In_9);
nor U2379 (N_2379,In_755,In_1789);
and U2380 (N_2380,In_2748,In_1108);
and U2381 (N_2381,In_2705,In_2090);
nand U2382 (N_2382,In_2061,In_1782);
and U2383 (N_2383,In_303,In_2670);
xor U2384 (N_2384,In_1694,In_2144);
nor U2385 (N_2385,In_2672,In_1930);
nor U2386 (N_2386,In_2573,In_2778);
and U2387 (N_2387,In_166,In_999);
or U2388 (N_2388,In_2677,In_1318);
xor U2389 (N_2389,In_128,In_2495);
xnor U2390 (N_2390,In_2033,In_708);
xnor U2391 (N_2391,In_2484,In_2349);
and U2392 (N_2392,In_850,In_1136);
or U2393 (N_2393,In_683,In_2580);
nand U2394 (N_2394,In_2128,In_50);
nor U2395 (N_2395,In_34,In_2123);
or U2396 (N_2396,In_1729,In_307);
or U2397 (N_2397,In_1227,In_879);
nand U2398 (N_2398,In_2915,In_227);
or U2399 (N_2399,In_1394,In_743);
xor U2400 (N_2400,In_2604,In_1548);
and U2401 (N_2401,In_252,In_2381);
nor U2402 (N_2402,In_2860,In_2704);
nand U2403 (N_2403,In_542,In_288);
or U2404 (N_2404,In_529,In_2518);
or U2405 (N_2405,In_2358,In_2541);
nand U2406 (N_2406,In_1552,In_121);
nor U2407 (N_2407,In_857,In_1678);
nand U2408 (N_2408,In_1155,In_881);
nand U2409 (N_2409,In_2276,In_439);
and U2410 (N_2410,In_1145,In_183);
nor U2411 (N_2411,In_638,In_1352);
or U2412 (N_2412,In_2739,In_2130);
or U2413 (N_2413,In_1863,In_2399);
or U2414 (N_2414,In_584,In_1780);
and U2415 (N_2415,In_1496,In_1801);
xor U2416 (N_2416,In_2208,In_911);
nand U2417 (N_2417,In_2028,In_144);
and U2418 (N_2418,In_2415,In_1817);
xnor U2419 (N_2419,In_451,In_844);
xnor U2420 (N_2420,In_2418,In_2400);
and U2421 (N_2421,In_390,In_898);
and U2422 (N_2422,In_388,In_2909);
nand U2423 (N_2423,In_1662,In_986);
and U2424 (N_2424,In_1488,In_946);
and U2425 (N_2425,In_2911,In_2570);
and U2426 (N_2426,In_1213,In_1772);
or U2427 (N_2427,In_1502,In_292);
nor U2428 (N_2428,In_16,In_2918);
and U2429 (N_2429,In_2685,In_2602);
xor U2430 (N_2430,In_2950,In_579);
nor U2431 (N_2431,In_1657,In_1508);
and U2432 (N_2432,In_2072,In_2140);
nand U2433 (N_2433,In_456,In_1124);
xnor U2434 (N_2434,In_1178,In_1046);
nand U2435 (N_2435,In_489,In_2914);
nand U2436 (N_2436,In_26,In_1102);
nand U2437 (N_2437,In_459,In_495);
and U2438 (N_2438,In_1651,In_130);
and U2439 (N_2439,In_1421,In_2316);
nor U2440 (N_2440,In_1298,In_2266);
xor U2441 (N_2441,In_1760,In_2473);
or U2442 (N_2442,In_957,In_2249);
and U2443 (N_2443,In_2279,In_2393);
nor U2444 (N_2444,In_1026,In_725);
and U2445 (N_2445,In_908,In_1240);
nor U2446 (N_2446,In_1108,In_2623);
nor U2447 (N_2447,In_1443,In_578);
nand U2448 (N_2448,In_1765,In_2493);
nor U2449 (N_2449,In_436,In_404);
xor U2450 (N_2450,In_138,In_1465);
nand U2451 (N_2451,In_625,In_1201);
or U2452 (N_2452,In_1132,In_670);
nand U2453 (N_2453,In_298,In_848);
or U2454 (N_2454,In_1526,In_1030);
xnor U2455 (N_2455,In_1195,In_2340);
nand U2456 (N_2456,In_363,In_2744);
or U2457 (N_2457,In_717,In_2624);
xnor U2458 (N_2458,In_598,In_281);
xor U2459 (N_2459,In_2987,In_2343);
nor U2460 (N_2460,In_437,In_288);
xnor U2461 (N_2461,In_2665,In_2137);
xnor U2462 (N_2462,In_1654,In_217);
nand U2463 (N_2463,In_859,In_2596);
or U2464 (N_2464,In_2321,In_2735);
or U2465 (N_2465,In_191,In_2540);
nor U2466 (N_2466,In_1277,In_1395);
and U2467 (N_2467,In_2911,In_970);
nor U2468 (N_2468,In_752,In_1888);
and U2469 (N_2469,In_261,In_1327);
nand U2470 (N_2470,In_518,In_1681);
and U2471 (N_2471,In_1874,In_2404);
nor U2472 (N_2472,In_2982,In_94);
xor U2473 (N_2473,In_1112,In_1921);
nand U2474 (N_2474,In_1725,In_2874);
nor U2475 (N_2475,In_2210,In_2434);
nand U2476 (N_2476,In_23,In_2577);
and U2477 (N_2477,In_468,In_2392);
nor U2478 (N_2478,In_824,In_383);
and U2479 (N_2479,In_1377,In_2423);
and U2480 (N_2480,In_915,In_1039);
nor U2481 (N_2481,In_2592,In_715);
nor U2482 (N_2482,In_1423,In_760);
nand U2483 (N_2483,In_574,In_1586);
or U2484 (N_2484,In_2047,In_811);
or U2485 (N_2485,In_2949,In_1479);
nor U2486 (N_2486,In_825,In_931);
and U2487 (N_2487,In_2062,In_1006);
and U2488 (N_2488,In_169,In_2360);
nor U2489 (N_2489,In_555,In_2946);
nor U2490 (N_2490,In_841,In_2533);
and U2491 (N_2491,In_2707,In_91);
and U2492 (N_2492,In_1408,In_1108);
nor U2493 (N_2493,In_2128,In_288);
and U2494 (N_2494,In_2235,In_1171);
xor U2495 (N_2495,In_847,In_1781);
and U2496 (N_2496,In_697,In_971);
xnor U2497 (N_2497,In_2108,In_2656);
or U2498 (N_2498,In_2143,In_1561);
nor U2499 (N_2499,In_377,In_1268);
nor U2500 (N_2500,In_2229,In_1091);
or U2501 (N_2501,In_668,In_1124);
nand U2502 (N_2502,In_2567,In_235);
xnor U2503 (N_2503,In_1858,In_46);
nand U2504 (N_2504,In_1740,In_1158);
or U2505 (N_2505,In_1872,In_425);
and U2506 (N_2506,In_1330,In_2136);
and U2507 (N_2507,In_2709,In_1934);
and U2508 (N_2508,In_1324,In_849);
xor U2509 (N_2509,In_293,In_259);
nor U2510 (N_2510,In_2642,In_2906);
xnor U2511 (N_2511,In_2462,In_2931);
and U2512 (N_2512,In_1933,In_463);
nor U2513 (N_2513,In_2125,In_137);
nor U2514 (N_2514,In_2139,In_2475);
and U2515 (N_2515,In_10,In_832);
xnor U2516 (N_2516,In_606,In_610);
nor U2517 (N_2517,In_1973,In_810);
nor U2518 (N_2518,In_2978,In_529);
nand U2519 (N_2519,In_826,In_1850);
and U2520 (N_2520,In_621,In_4);
or U2521 (N_2521,In_2768,In_1429);
and U2522 (N_2522,In_380,In_2862);
or U2523 (N_2523,In_811,In_2561);
nand U2524 (N_2524,In_1689,In_2973);
nor U2525 (N_2525,In_2872,In_2358);
xor U2526 (N_2526,In_237,In_1858);
xor U2527 (N_2527,In_28,In_1024);
nand U2528 (N_2528,In_2508,In_15);
or U2529 (N_2529,In_1320,In_1206);
nor U2530 (N_2530,In_2070,In_946);
or U2531 (N_2531,In_734,In_435);
or U2532 (N_2532,In_557,In_1418);
nor U2533 (N_2533,In_976,In_1257);
nand U2534 (N_2534,In_1938,In_2579);
nor U2535 (N_2535,In_2233,In_1556);
nand U2536 (N_2536,In_1766,In_1442);
nand U2537 (N_2537,In_1188,In_127);
nor U2538 (N_2538,In_567,In_2475);
nand U2539 (N_2539,In_2459,In_2262);
xnor U2540 (N_2540,In_137,In_332);
or U2541 (N_2541,In_2141,In_2608);
or U2542 (N_2542,In_1909,In_1528);
and U2543 (N_2543,In_564,In_2136);
xnor U2544 (N_2544,In_1936,In_1622);
nor U2545 (N_2545,In_2286,In_1709);
nor U2546 (N_2546,In_183,In_1745);
xor U2547 (N_2547,In_1129,In_248);
or U2548 (N_2548,In_810,In_1515);
xnor U2549 (N_2549,In_2376,In_1768);
xor U2550 (N_2550,In_1029,In_1756);
or U2551 (N_2551,In_1331,In_531);
nor U2552 (N_2552,In_1413,In_1469);
nand U2553 (N_2553,In_295,In_867);
and U2554 (N_2554,In_408,In_1546);
and U2555 (N_2555,In_284,In_2985);
and U2556 (N_2556,In_1358,In_597);
nand U2557 (N_2557,In_2280,In_1883);
nand U2558 (N_2558,In_2154,In_84);
xor U2559 (N_2559,In_770,In_1407);
nor U2560 (N_2560,In_308,In_2471);
xnor U2561 (N_2561,In_930,In_2032);
and U2562 (N_2562,In_461,In_726);
nand U2563 (N_2563,In_2652,In_2364);
xor U2564 (N_2564,In_1827,In_2285);
xor U2565 (N_2565,In_2118,In_860);
nor U2566 (N_2566,In_2985,In_1278);
nor U2567 (N_2567,In_1902,In_224);
xor U2568 (N_2568,In_25,In_942);
nand U2569 (N_2569,In_2690,In_749);
or U2570 (N_2570,In_2760,In_268);
xnor U2571 (N_2571,In_1903,In_1589);
nor U2572 (N_2572,In_1319,In_2510);
and U2573 (N_2573,In_2118,In_2504);
or U2574 (N_2574,In_2588,In_436);
and U2575 (N_2575,In_1617,In_2322);
xor U2576 (N_2576,In_21,In_951);
nand U2577 (N_2577,In_289,In_2300);
and U2578 (N_2578,In_2282,In_1796);
or U2579 (N_2579,In_1670,In_2025);
or U2580 (N_2580,In_2173,In_2346);
nor U2581 (N_2581,In_1405,In_731);
xor U2582 (N_2582,In_315,In_2807);
and U2583 (N_2583,In_1203,In_2010);
xnor U2584 (N_2584,In_2667,In_1970);
nand U2585 (N_2585,In_673,In_581);
and U2586 (N_2586,In_2196,In_2494);
or U2587 (N_2587,In_451,In_56);
or U2588 (N_2588,In_1052,In_1103);
and U2589 (N_2589,In_1475,In_2555);
and U2590 (N_2590,In_369,In_265);
nor U2591 (N_2591,In_1463,In_2483);
or U2592 (N_2592,In_572,In_2719);
and U2593 (N_2593,In_2749,In_919);
xor U2594 (N_2594,In_624,In_272);
and U2595 (N_2595,In_1699,In_2262);
nor U2596 (N_2596,In_1239,In_2244);
and U2597 (N_2597,In_1652,In_2392);
and U2598 (N_2598,In_576,In_1682);
or U2599 (N_2599,In_1672,In_2732);
or U2600 (N_2600,In_1518,In_2564);
or U2601 (N_2601,In_1333,In_1801);
and U2602 (N_2602,In_2162,In_1274);
or U2603 (N_2603,In_1745,In_514);
nor U2604 (N_2604,In_438,In_611);
and U2605 (N_2605,In_2827,In_1967);
nand U2606 (N_2606,In_522,In_1828);
xor U2607 (N_2607,In_2384,In_540);
or U2608 (N_2608,In_1286,In_1337);
nand U2609 (N_2609,In_2560,In_2756);
xnor U2610 (N_2610,In_1811,In_2727);
and U2611 (N_2611,In_435,In_2885);
xnor U2612 (N_2612,In_58,In_1363);
and U2613 (N_2613,In_175,In_408);
nor U2614 (N_2614,In_1813,In_2798);
and U2615 (N_2615,In_581,In_2112);
nand U2616 (N_2616,In_392,In_2669);
nand U2617 (N_2617,In_1955,In_1127);
or U2618 (N_2618,In_608,In_2783);
or U2619 (N_2619,In_1502,In_2394);
nor U2620 (N_2620,In_1810,In_2750);
or U2621 (N_2621,In_1881,In_1287);
nor U2622 (N_2622,In_1812,In_262);
nand U2623 (N_2623,In_2399,In_2653);
nand U2624 (N_2624,In_2113,In_700);
or U2625 (N_2625,In_858,In_2571);
and U2626 (N_2626,In_2709,In_1994);
nor U2627 (N_2627,In_1086,In_1209);
nand U2628 (N_2628,In_2752,In_305);
and U2629 (N_2629,In_1818,In_113);
and U2630 (N_2630,In_1365,In_647);
or U2631 (N_2631,In_1227,In_2817);
nor U2632 (N_2632,In_1617,In_315);
nor U2633 (N_2633,In_2766,In_348);
nor U2634 (N_2634,In_2886,In_136);
nor U2635 (N_2635,In_1757,In_2114);
and U2636 (N_2636,In_1303,In_945);
and U2637 (N_2637,In_1225,In_1778);
and U2638 (N_2638,In_1718,In_26);
nor U2639 (N_2639,In_1223,In_1988);
and U2640 (N_2640,In_857,In_937);
nand U2641 (N_2641,In_836,In_2866);
and U2642 (N_2642,In_1665,In_982);
nor U2643 (N_2643,In_847,In_397);
and U2644 (N_2644,In_521,In_1257);
and U2645 (N_2645,In_2619,In_1666);
nor U2646 (N_2646,In_676,In_706);
nor U2647 (N_2647,In_953,In_1700);
nor U2648 (N_2648,In_2053,In_1672);
xnor U2649 (N_2649,In_2239,In_1190);
or U2650 (N_2650,In_2103,In_1846);
nand U2651 (N_2651,In_1392,In_248);
nand U2652 (N_2652,In_28,In_680);
nand U2653 (N_2653,In_1858,In_1304);
nand U2654 (N_2654,In_410,In_2090);
and U2655 (N_2655,In_1848,In_477);
nor U2656 (N_2656,In_305,In_251);
nand U2657 (N_2657,In_1792,In_1871);
and U2658 (N_2658,In_2417,In_1777);
nand U2659 (N_2659,In_2895,In_789);
xnor U2660 (N_2660,In_1215,In_50);
and U2661 (N_2661,In_1208,In_2480);
nor U2662 (N_2662,In_2435,In_379);
nand U2663 (N_2663,In_1596,In_1029);
nor U2664 (N_2664,In_1869,In_530);
xor U2665 (N_2665,In_56,In_2563);
nor U2666 (N_2666,In_630,In_1871);
nor U2667 (N_2667,In_2892,In_2465);
nand U2668 (N_2668,In_657,In_2893);
nand U2669 (N_2669,In_90,In_1477);
or U2670 (N_2670,In_2012,In_505);
xor U2671 (N_2671,In_2725,In_699);
and U2672 (N_2672,In_2343,In_1277);
nand U2673 (N_2673,In_2406,In_671);
or U2674 (N_2674,In_2966,In_299);
nor U2675 (N_2675,In_2561,In_101);
xor U2676 (N_2676,In_2015,In_1178);
nand U2677 (N_2677,In_2771,In_1781);
and U2678 (N_2678,In_1074,In_2366);
nand U2679 (N_2679,In_1415,In_212);
and U2680 (N_2680,In_333,In_550);
and U2681 (N_2681,In_1776,In_1089);
nor U2682 (N_2682,In_356,In_2912);
and U2683 (N_2683,In_1115,In_1984);
and U2684 (N_2684,In_1157,In_91);
nor U2685 (N_2685,In_639,In_1348);
and U2686 (N_2686,In_1560,In_1692);
nor U2687 (N_2687,In_2595,In_1219);
nor U2688 (N_2688,In_653,In_2698);
and U2689 (N_2689,In_2510,In_1231);
or U2690 (N_2690,In_1877,In_2551);
nand U2691 (N_2691,In_2600,In_1307);
and U2692 (N_2692,In_2840,In_323);
or U2693 (N_2693,In_2230,In_1204);
or U2694 (N_2694,In_2514,In_686);
xnor U2695 (N_2695,In_406,In_810);
nand U2696 (N_2696,In_612,In_2960);
nand U2697 (N_2697,In_2885,In_80);
nor U2698 (N_2698,In_929,In_2962);
nor U2699 (N_2699,In_2846,In_1938);
nor U2700 (N_2700,In_349,In_402);
and U2701 (N_2701,In_1382,In_2);
nand U2702 (N_2702,In_1276,In_2478);
nand U2703 (N_2703,In_2578,In_2950);
or U2704 (N_2704,In_2,In_2101);
xnor U2705 (N_2705,In_843,In_1352);
or U2706 (N_2706,In_2193,In_2637);
and U2707 (N_2707,In_1719,In_2965);
nand U2708 (N_2708,In_1973,In_988);
nor U2709 (N_2709,In_2740,In_2207);
or U2710 (N_2710,In_1796,In_410);
xor U2711 (N_2711,In_274,In_1813);
nand U2712 (N_2712,In_2155,In_1934);
or U2713 (N_2713,In_942,In_512);
nand U2714 (N_2714,In_663,In_1713);
nor U2715 (N_2715,In_2817,In_1903);
and U2716 (N_2716,In_898,In_2430);
nor U2717 (N_2717,In_524,In_23);
and U2718 (N_2718,In_1470,In_1044);
xor U2719 (N_2719,In_1520,In_804);
xor U2720 (N_2720,In_382,In_946);
nor U2721 (N_2721,In_2488,In_1535);
or U2722 (N_2722,In_1633,In_2947);
xor U2723 (N_2723,In_1342,In_2734);
nor U2724 (N_2724,In_1944,In_660);
or U2725 (N_2725,In_743,In_1482);
xor U2726 (N_2726,In_428,In_1256);
nor U2727 (N_2727,In_614,In_632);
nor U2728 (N_2728,In_80,In_2163);
nand U2729 (N_2729,In_2236,In_508);
xnor U2730 (N_2730,In_2442,In_2862);
nand U2731 (N_2731,In_713,In_1733);
xnor U2732 (N_2732,In_652,In_1258);
or U2733 (N_2733,In_567,In_1692);
nand U2734 (N_2734,In_1400,In_1282);
and U2735 (N_2735,In_1091,In_1647);
and U2736 (N_2736,In_1669,In_255);
and U2737 (N_2737,In_232,In_1468);
nand U2738 (N_2738,In_740,In_2404);
xnor U2739 (N_2739,In_1534,In_586);
or U2740 (N_2740,In_1253,In_924);
nor U2741 (N_2741,In_2167,In_2019);
xnor U2742 (N_2742,In_499,In_46);
xnor U2743 (N_2743,In_703,In_1390);
nand U2744 (N_2744,In_490,In_55);
nor U2745 (N_2745,In_1068,In_2362);
nor U2746 (N_2746,In_2155,In_1422);
and U2747 (N_2747,In_1812,In_2355);
nor U2748 (N_2748,In_2771,In_390);
or U2749 (N_2749,In_2564,In_1485);
and U2750 (N_2750,In_83,In_970);
and U2751 (N_2751,In_2699,In_2908);
and U2752 (N_2752,In_2770,In_1745);
xnor U2753 (N_2753,In_2393,In_495);
and U2754 (N_2754,In_2414,In_1095);
xor U2755 (N_2755,In_2127,In_315);
and U2756 (N_2756,In_1977,In_164);
and U2757 (N_2757,In_269,In_620);
xor U2758 (N_2758,In_1278,In_511);
nor U2759 (N_2759,In_1406,In_681);
and U2760 (N_2760,In_1326,In_1852);
nand U2761 (N_2761,In_385,In_2664);
nand U2762 (N_2762,In_686,In_2885);
xnor U2763 (N_2763,In_2089,In_1851);
nand U2764 (N_2764,In_266,In_185);
nor U2765 (N_2765,In_800,In_2879);
xor U2766 (N_2766,In_548,In_1229);
xor U2767 (N_2767,In_2486,In_1343);
nor U2768 (N_2768,In_2802,In_2924);
nand U2769 (N_2769,In_718,In_2492);
or U2770 (N_2770,In_1174,In_2371);
nor U2771 (N_2771,In_1771,In_2248);
nor U2772 (N_2772,In_1470,In_1732);
xnor U2773 (N_2773,In_3,In_2863);
nand U2774 (N_2774,In_208,In_2849);
nand U2775 (N_2775,In_456,In_881);
nor U2776 (N_2776,In_1360,In_1793);
and U2777 (N_2777,In_1478,In_1603);
xor U2778 (N_2778,In_1151,In_883);
nand U2779 (N_2779,In_2158,In_2350);
or U2780 (N_2780,In_563,In_2884);
or U2781 (N_2781,In_2986,In_1840);
or U2782 (N_2782,In_1466,In_1450);
and U2783 (N_2783,In_912,In_980);
xor U2784 (N_2784,In_1912,In_1662);
and U2785 (N_2785,In_100,In_667);
or U2786 (N_2786,In_631,In_913);
and U2787 (N_2787,In_1898,In_2531);
and U2788 (N_2788,In_1840,In_740);
nor U2789 (N_2789,In_703,In_841);
or U2790 (N_2790,In_130,In_1676);
and U2791 (N_2791,In_2770,In_181);
and U2792 (N_2792,In_2663,In_432);
xor U2793 (N_2793,In_2825,In_2639);
nand U2794 (N_2794,In_804,In_486);
or U2795 (N_2795,In_261,In_476);
xor U2796 (N_2796,In_2485,In_1305);
nand U2797 (N_2797,In_1742,In_451);
or U2798 (N_2798,In_1060,In_2190);
or U2799 (N_2799,In_503,In_2631);
or U2800 (N_2800,In_835,In_1661);
and U2801 (N_2801,In_693,In_2739);
xnor U2802 (N_2802,In_1793,In_1767);
xnor U2803 (N_2803,In_1638,In_736);
xor U2804 (N_2804,In_1132,In_981);
and U2805 (N_2805,In_760,In_176);
and U2806 (N_2806,In_1014,In_503);
nand U2807 (N_2807,In_1772,In_1878);
nand U2808 (N_2808,In_2039,In_1189);
nor U2809 (N_2809,In_19,In_2976);
or U2810 (N_2810,In_1565,In_526);
nand U2811 (N_2811,In_456,In_301);
or U2812 (N_2812,In_2521,In_1301);
nand U2813 (N_2813,In_1343,In_2050);
nor U2814 (N_2814,In_2378,In_2093);
and U2815 (N_2815,In_692,In_2865);
xor U2816 (N_2816,In_1133,In_1171);
and U2817 (N_2817,In_725,In_1420);
or U2818 (N_2818,In_1560,In_2017);
nand U2819 (N_2819,In_2343,In_1444);
nand U2820 (N_2820,In_282,In_1847);
nor U2821 (N_2821,In_1815,In_521);
xnor U2822 (N_2822,In_2452,In_530);
and U2823 (N_2823,In_1320,In_2848);
and U2824 (N_2824,In_902,In_2502);
and U2825 (N_2825,In_158,In_1173);
and U2826 (N_2826,In_326,In_204);
xnor U2827 (N_2827,In_2579,In_67);
nand U2828 (N_2828,In_2990,In_951);
nand U2829 (N_2829,In_394,In_964);
or U2830 (N_2830,In_1321,In_2570);
nand U2831 (N_2831,In_663,In_1418);
nand U2832 (N_2832,In_134,In_1157);
and U2833 (N_2833,In_349,In_1129);
nor U2834 (N_2834,In_2606,In_602);
nand U2835 (N_2835,In_849,In_2062);
and U2836 (N_2836,In_86,In_2708);
or U2837 (N_2837,In_1620,In_2380);
and U2838 (N_2838,In_1898,In_1753);
xnor U2839 (N_2839,In_674,In_1112);
xnor U2840 (N_2840,In_901,In_2353);
xnor U2841 (N_2841,In_73,In_835);
and U2842 (N_2842,In_2138,In_2576);
or U2843 (N_2843,In_1549,In_1744);
and U2844 (N_2844,In_2066,In_1916);
nand U2845 (N_2845,In_2886,In_2547);
nor U2846 (N_2846,In_2621,In_1816);
or U2847 (N_2847,In_694,In_1059);
or U2848 (N_2848,In_2346,In_1336);
xor U2849 (N_2849,In_2288,In_632);
xnor U2850 (N_2850,In_1122,In_201);
nand U2851 (N_2851,In_1176,In_2378);
and U2852 (N_2852,In_2259,In_2842);
or U2853 (N_2853,In_2881,In_210);
xor U2854 (N_2854,In_2163,In_750);
nor U2855 (N_2855,In_2619,In_1560);
and U2856 (N_2856,In_181,In_2372);
or U2857 (N_2857,In_1745,In_647);
xor U2858 (N_2858,In_1383,In_1386);
xor U2859 (N_2859,In_1086,In_39);
nor U2860 (N_2860,In_1885,In_2142);
xor U2861 (N_2861,In_1031,In_327);
or U2862 (N_2862,In_2758,In_1729);
and U2863 (N_2863,In_2481,In_294);
nand U2864 (N_2864,In_2119,In_1856);
nand U2865 (N_2865,In_961,In_1892);
or U2866 (N_2866,In_2825,In_1830);
and U2867 (N_2867,In_2134,In_1856);
xor U2868 (N_2868,In_1806,In_1842);
xnor U2869 (N_2869,In_1082,In_2975);
or U2870 (N_2870,In_2669,In_2151);
nor U2871 (N_2871,In_2100,In_543);
xor U2872 (N_2872,In_2583,In_724);
nand U2873 (N_2873,In_462,In_1346);
and U2874 (N_2874,In_1219,In_127);
or U2875 (N_2875,In_2320,In_828);
or U2876 (N_2876,In_1976,In_1490);
xnor U2877 (N_2877,In_829,In_2299);
nor U2878 (N_2878,In_460,In_1938);
or U2879 (N_2879,In_107,In_2854);
and U2880 (N_2880,In_2730,In_2635);
xnor U2881 (N_2881,In_2690,In_2278);
nand U2882 (N_2882,In_1784,In_2092);
xor U2883 (N_2883,In_819,In_1585);
and U2884 (N_2884,In_758,In_477);
and U2885 (N_2885,In_1743,In_1768);
and U2886 (N_2886,In_399,In_277);
or U2887 (N_2887,In_2189,In_1762);
or U2888 (N_2888,In_652,In_1252);
or U2889 (N_2889,In_1127,In_645);
xor U2890 (N_2890,In_2309,In_2731);
or U2891 (N_2891,In_58,In_1600);
or U2892 (N_2892,In_1138,In_2051);
or U2893 (N_2893,In_565,In_2633);
nand U2894 (N_2894,In_2366,In_604);
and U2895 (N_2895,In_1528,In_1536);
and U2896 (N_2896,In_376,In_458);
xor U2897 (N_2897,In_81,In_1727);
or U2898 (N_2898,In_1888,In_2987);
nor U2899 (N_2899,In_2291,In_1181);
or U2900 (N_2900,In_2519,In_2082);
xor U2901 (N_2901,In_2597,In_2863);
or U2902 (N_2902,In_568,In_1028);
xor U2903 (N_2903,In_346,In_1234);
xnor U2904 (N_2904,In_492,In_1923);
or U2905 (N_2905,In_1144,In_1345);
nor U2906 (N_2906,In_1601,In_2237);
nand U2907 (N_2907,In_1368,In_515);
nor U2908 (N_2908,In_1930,In_1130);
and U2909 (N_2909,In_2284,In_2927);
nor U2910 (N_2910,In_2457,In_372);
nand U2911 (N_2911,In_2456,In_1731);
nand U2912 (N_2912,In_1254,In_370);
and U2913 (N_2913,In_1017,In_456);
or U2914 (N_2914,In_135,In_1608);
nor U2915 (N_2915,In_1137,In_1269);
nor U2916 (N_2916,In_2463,In_857);
and U2917 (N_2917,In_1933,In_732);
nor U2918 (N_2918,In_1935,In_2849);
or U2919 (N_2919,In_25,In_2245);
or U2920 (N_2920,In_742,In_1703);
and U2921 (N_2921,In_871,In_303);
xnor U2922 (N_2922,In_2795,In_1326);
nand U2923 (N_2923,In_1383,In_783);
nor U2924 (N_2924,In_2749,In_2099);
or U2925 (N_2925,In_2313,In_1692);
nor U2926 (N_2926,In_1177,In_788);
nand U2927 (N_2927,In_1697,In_1325);
and U2928 (N_2928,In_1123,In_726);
nand U2929 (N_2929,In_418,In_945);
and U2930 (N_2930,In_2921,In_2404);
nor U2931 (N_2931,In_2925,In_320);
or U2932 (N_2932,In_2584,In_866);
or U2933 (N_2933,In_180,In_2698);
or U2934 (N_2934,In_1063,In_2838);
nor U2935 (N_2935,In_1556,In_860);
nor U2936 (N_2936,In_378,In_741);
nor U2937 (N_2937,In_2151,In_1834);
and U2938 (N_2938,In_910,In_2328);
nand U2939 (N_2939,In_1105,In_2097);
nand U2940 (N_2940,In_1260,In_2629);
or U2941 (N_2941,In_371,In_2148);
nor U2942 (N_2942,In_2130,In_1780);
and U2943 (N_2943,In_1784,In_1616);
nor U2944 (N_2944,In_2231,In_1037);
nor U2945 (N_2945,In_2430,In_611);
and U2946 (N_2946,In_189,In_2877);
and U2947 (N_2947,In_2294,In_1206);
xnor U2948 (N_2948,In_1465,In_2150);
xnor U2949 (N_2949,In_1512,In_1898);
or U2950 (N_2950,In_2362,In_940);
nor U2951 (N_2951,In_772,In_2223);
nand U2952 (N_2952,In_2772,In_131);
nand U2953 (N_2953,In_2648,In_2876);
and U2954 (N_2954,In_66,In_862);
or U2955 (N_2955,In_1176,In_819);
and U2956 (N_2956,In_105,In_2672);
xor U2957 (N_2957,In_1674,In_2911);
and U2958 (N_2958,In_2189,In_2640);
nand U2959 (N_2959,In_2022,In_655);
nand U2960 (N_2960,In_2619,In_2325);
xor U2961 (N_2961,In_428,In_2104);
nand U2962 (N_2962,In_1272,In_1391);
nor U2963 (N_2963,In_2156,In_2765);
nor U2964 (N_2964,In_137,In_2849);
nor U2965 (N_2965,In_1288,In_20);
nor U2966 (N_2966,In_939,In_706);
nor U2967 (N_2967,In_481,In_1096);
nor U2968 (N_2968,In_1788,In_2156);
and U2969 (N_2969,In_1265,In_2525);
xnor U2970 (N_2970,In_209,In_693);
nand U2971 (N_2971,In_2966,In_2990);
and U2972 (N_2972,In_467,In_922);
xor U2973 (N_2973,In_989,In_2423);
or U2974 (N_2974,In_332,In_1205);
and U2975 (N_2975,In_1155,In_2840);
nor U2976 (N_2976,In_546,In_1008);
xnor U2977 (N_2977,In_2226,In_2815);
nor U2978 (N_2978,In_1287,In_2861);
xnor U2979 (N_2979,In_2755,In_583);
and U2980 (N_2980,In_1387,In_1630);
xnor U2981 (N_2981,In_1227,In_2487);
and U2982 (N_2982,In_1992,In_1285);
and U2983 (N_2983,In_2672,In_1568);
or U2984 (N_2984,In_2685,In_2735);
or U2985 (N_2985,In_1834,In_517);
and U2986 (N_2986,In_2503,In_430);
xnor U2987 (N_2987,In_529,In_469);
nand U2988 (N_2988,In_816,In_2918);
nand U2989 (N_2989,In_1,In_1951);
nand U2990 (N_2990,In_2519,In_585);
and U2991 (N_2991,In_2961,In_522);
nor U2992 (N_2992,In_2000,In_2001);
xnor U2993 (N_2993,In_242,In_569);
xor U2994 (N_2994,In_2726,In_677);
and U2995 (N_2995,In_2010,In_2704);
or U2996 (N_2996,In_2770,In_1856);
or U2997 (N_2997,In_1520,In_2879);
nor U2998 (N_2998,In_2057,In_1149);
and U2999 (N_2999,In_585,In_2602);
xnor U3000 (N_3000,In_1446,In_146);
or U3001 (N_3001,In_1143,In_1094);
and U3002 (N_3002,In_307,In_2720);
nand U3003 (N_3003,In_2980,In_2071);
nand U3004 (N_3004,In_2511,In_143);
xnor U3005 (N_3005,In_55,In_2152);
or U3006 (N_3006,In_568,In_1405);
nor U3007 (N_3007,In_1594,In_783);
nor U3008 (N_3008,In_332,In_2691);
and U3009 (N_3009,In_102,In_466);
xnor U3010 (N_3010,In_73,In_2496);
or U3011 (N_3011,In_392,In_268);
nor U3012 (N_3012,In_286,In_754);
and U3013 (N_3013,In_1012,In_2944);
or U3014 (N_3014,In_947,In_2352);
nor U3015 (N_3015,In_2570,In_1693);
and U3016 (N_3016,In_854,In_822);
or U3017 (N_3017,In_1916,In_424);
nand U3018 (N_3018,In_561,In_1175);
nand U3019 (N_3019,In_2057,In_2204);
or U3020 (N_3020,In_653,In_872);
or U3021 (N_3021,In_417,In_2822);
and U3022 (N_3022,In_2152,In_1701);
nand U3023 (N_3023,In_1644,In_275);
xor U3024 (N_3024,In_2472,In_174);
or U3025 (N_3025,In_2954,In_2923);
nor U3026 (N_3026,In_1881,In_2097);
and U3027 (N_3027,In_2957,In_131);
and U3028 (N_3028,In_1975,In_1427);
and U3029 (N_3029,In_2108,In_1519);
or U3030 (N_3030,In_2503,In_298);
nor U3031 (N_3031,In_2696,In_2392);
nor U3032 (N_3032,In_2551,In_563);
nand U3033 (N_3033,In_823,In_2082);
nor U3034 (N_3034,In_1410,In_1267);
and U3035 (N_3035,In_2225,In_958);
nor U3036 (N_3036,In_2474,In_2464);
xor U3037 (N_3037,In_981,In_807);
and U3038 (N_3038,In_207,In_2988);
and U3039 (N_3039,In_1951,In_398);
nand U3040 (N_3040,In_1246,In_978);
xnor U3041 (N_3041,In_2989,In_2620);
xnor U3042 (N_3042,In_2297,In_2484);
nor U3043 (N_3043,In_931,In_1764);
or U3044 (N_3044,In_283,In_1518);
nand U3045 (N_3045,In_2628,In_1496);
nand U3046 (N_3046,In_988,In_2408);
nor U3047 (N_3047,In_1627,In_317);
or U3048 (N_3048,In_1454,In_1457);
nand U3049 (N_3049,In_2108,In_737);
or U3050 (N_3050,In_2798,In_1940);
and U3051 (N_3051,In_787,In_371);
nand U3052 (N_3052,In_2666,In_912);
nand U3053 (N_3053,In_1848,In_281);
or U3054 (N_3054,In_2809,In_705);
or U3055 (N_3055,In_1352,In_109);
or U3056 (N_3056,In_132,In_1493);
nand U3057 (N_3057,In_564,In_1627);
nand U3058 (N_3058,In_1814,In_639);
nand U3059 (N_3059,In_1438,In_2484);
or U3060 (N_3060,In_418,In_75);
nand U3061 (N_3061,In_2390,In_2318);
or U3062 (N_3062,In_1669,In_2083);
or U3063 (N_3063,In_2076,In_1735);
nor U3064 (N_3064,In_707,In_499);
nor U3065 (N_3065,In_1107,In_2104);
and U3066 (N_3066,In_2226,In_909);
and U3067 (N_3067,In_2757,In_1261);
and U3068 (N_3068,In_2434,In_2490);
nand U3069 (N_3069,In_2536,In_2334);
xnor U3070 (N_3070,In_2142,In_833);
nand U3071 (N_3071,In_2847,In_1064);
nor U3072 (N_3072,In_843,In_1448);
nor U3073 (N_3073,In_1135,In_1203);
nor U3074 (N_3074,In_1410,In_1245);
and U3075 (N_3075,In_2677,In_2793);
nor U3076 (N_3076,In_1490,In_617);
and U3077 (N_3077,In_2208,In_2218);
and U3078 (N_3078,In_2036,In_94);
and U3079 (N_3079,In_2299,In_438);
or U3080 (N_3080,In_147,In_2341);
nor U3081 (N_3081,In_91,In_575);
or U3082 (N_3082,In_1717,In_2455);
or U3083 (N_3083,In_882,In_678);
xor U3084 (N_3084,In_508,In_2690);
and U3085 (N_3085,In_1146,In_993);
or U3086 (N_3086,In_2122,In_1661);
and U3087 (N_3087,In_1893,In_1170);
and U3088 (N_3088,In_1853,In_1494);
nand U3089 (N_3089,In_715,In_2404);
nor U3090 (N_3090,In_299,In_71);
or U3091 (N_3091,In_1128,In_1275);
or U3092 (N_3092,In_573,In_2315);
xor U3093 (N_3093,In_841,In_593);
nor U3094 (N_3094,In_672,In_1017);
or U3095 (N_3095,In_2216,In_2486);
and U3096 (N_3096,In_1952,In_1513);
or U3097 (N_3097,In_945,In_1497);
nor U3098 (N_3098,In_1719,In_351);
xnor U3099 (N_3099,In_1604,In_521);
or U3100 (N_3100,In_1375,In_12);
xnor U3101 (N_3101,In_2515,In_2924);
and U3102 (N_3102,In_2001,In_215);
nor U3103 (N_3103,In_1151,In_39);
or U3104 (N_3104,In_506,In_577);
nor U3105 (N_3105,In_1029,In_2872);
nor U3106 (N_3106,In_712,In_2172);
or U3107 (N_3107,In_245,In_2483);
and U3108 (N_3108,In_1658,In_1699);
nand U3109 (N_3109,In_1196,In_1707);
or U3110 (N_3110,In_1163,In_1040);
and U3111 (N_3111,In_2,In_1006);
nor U3112 (N_3112,In_2399,In_216);
and U3113 (N_3113,In_2556,In_2906);
nor U3114 (N_3114,In_2336,In_1981);
and U3115 (N_3115,In_1875,In_836);
nand U3116 (N_3116,In_2862,In_387);
xnor U3117 (N_3117,In_2231,In_2127);
xnor U3118 (N_3118,In_1915,In_2067);
xor U3119 (N_3119,In_1183,In_2856);
nand U3120 (N_3120,In_1385,In_898);
xor U3121 (N_3121,In_2437,In_2493);
xnor U3122 (N_3122,In_388,In_958);
xor U3123 (N_3123,In_605,In_2163);
nor U3124 (N_3124,In_1081,In_2405);
nand U3125 (N_3125,In_2681,In_522);
nand U3126 (N_3126,In_1454,In_586);
or U3127 (N_3127,In_1709,In_548);
xnor U3128 (N_3128,In_326,In_1355);
xor U3129 (N_3129,In_899,In_319);
or U3130 (N_3130,In_2181,In_1201);
nand U3131 (N_3131,In_1075,In_2445);
nand U3132 (N_3132,In_1715,In_2713);
and U3133 (N_3133,In_1847,In_2390);
and U3134 (N_3134,In_588,In_1162);
xnor U3135 (N_3135,In_45,In_392);
nand U3136 (N_3136,In_1531,In_2064);
nand U3137 (N_3137,In_2531,In_2160);
and U3138 (N_3138,In_2793,In_858);
or U3139 (N_3139,In_201,In_2672);
nor U3140 (N_3140,In_286,In_1133);
nand U3141 (N_3141,In_2654,In_1090);
or U3142 (N_3142,In_2412,In_1590);
nand U3143 (N_3143,In_1158,In_1354);
nand U3144 (N_3144,In_450,In_1236);
xor U3145 (N_3145,In_2662,In_593);
and U3146 (N_3146,In_1419,In_1092);
nor U3147 (N_3147,In_281,In_1702);
nand U3148 (N_3148,In_958,In_435);
nand U3149 (N_3149,In_2429,In_1900);
nand U3150 (N_3150,In_262,In_1021);
xnor U3151 (N_3151,In_624,In_2718);
nor U3152 (N_3152,In_1758,In_2578);
and U3153 (N_3153,In_1242,In_1183);
or U3154 (N_3154,In_1070,In_1569);
nor U3155 (N_3155,In_1418,In_793);
nor U3156 (N_3156,In_611,In_2404);
nand U3157 (N_3157,In_831,In_2966);
xnor U3158 (N_3158,In_2915,In_747);
xnor U3159 (N_3159,In_2037,In_893);
and U3160 (N_3160,In_2936,In_1861);
nand U3161 (N_3161,In_1417,In_309);
and U3162 (N_3162,In_2104,In_1027);
nand U3163 (N_3163,In_2478,In_2612);
xor U3164 (N_3164,In_1144,In_194);
nand U3165 (N_3165,In_836,In_2096);
or U3166 (N_3166,In_1028,In_2266);
nand U3167 (N_3167,In_2768,In_392);
xnor U3168 (N_3168,In_2953,In_620);
nand U3169 (N_3169,In_1167,In_2697);
xnor U3170 (N_3170,In_689,In_1964);
nand U3171 (N_3171,In_585,In_2444);
nor U3172 (N_3172,In_497,In_384);
nand U3173 (N_3173,In_1843,In_1237);
nor U3174 (N_3174,In_2489,In_738);
or U3175 (N_3175,In_481,In_315);
xor U3176 (N_3176,In_1791,In_1331);
xnor U3177 (N_3177,In_1471,In_229);
nand U3178 (N_3178,In_119,In_1819);
nor U3179 (N_3179,In_1805,In_515);
xor U3180 (N_3180,In_138,In_2591);
or U3181 (N_3181,In_180,In_1974);
xor U3182 (N_3182,In_798,In_2186);
xnor U3183 (N_3183,In_967,In_2211);
xor U3184 (N_3184,In_2135,In_907);
and U3185 (N_3185,In_539,In_205);
nand U3186 (N_3186,In_2300,In_986);
nand U3187 (N_3187,In_1057,In_1383);
nor U3188 (N_3188,In_1098,In_2337);
xnor U3189 (N_3189,In_189,In_141);
or U3190 (N_3190,In_329,In_2723);
xor U3191 (N_3191,In_1917,In_1981);
or U3192 (N_3192,In_540,In_1759);
nand U3193 (N_3193,In_2772,In_2775);
nor U3194 (N_3194,In_2916,In_1308);
xor U3195 (N_3195,In_2441,In_1914);
or U3196 (N_3196,In_1921,In_1697);
nand U3197 (N_3197,In_2595,In_1631);
or U3198 (N_3198,In_1642,In_2842);
or U3199 (N_3199,In_1692,In_2557);
xnor U3200 (N_3200,In_1153,In_2089);
and U3201 (N_3201,In_1430,In_523);
nor U3202 (N_3202,In_459,In_946);
xor U3203 (N_3203,In_1187,In_2778);
and U3204 (N_3204,In_1263,In_2947);
and U3205 (N_3205,In_1605,In_2845);
nand U3206 (N_3206,In_2501,In_22);
xnor U3207 (N_3207,In_47,In_2326);
or U3208 (N_3208,In_1808,In_625);
and U3209 (N_3209,In_1530,In_1299);
or U3210 (N_3210,In_2151,In_2327);
nor U3211 (N_3211,In_1939,In_611);
or U3212 (N_3212,In_1344,In_2214);
xnor U3213 (N_3213,In_1523,In_1475);
xor U3214 (N_3214,In_697,In_818);
and U3215 (N_3215,In_540,In_1647);
and U3216 (N_3216,In_1619,In_601);
or U3217 (N_3217,In_1821,In_1964);
nand U3218 (N_3218,In_917,In_1258);
nand U3219 (N_3219,In_903,In_2500);
nand U3220 (N_3220,In_2710,In_431);
nand U3221 (N_3221,In_2775,In_326);
and U3222 (N_3222,In_392,In_892);
nor U3223 (N_3223,In_1397,In_2343);
or U3224 (N_3224,In_2981,In_2970);
xor U3225 (N_3225,In_1576,In_2527);
or U3226 (N_3226,In_927,In_2572);
or U3227 (N_3227,In_97,In_233);
nor U3228 (N_3228,In_639,In_1472);
nand U3229 (N_3229,In_1630,In_1854);
nand U3230 (N_3230,In_450,In_1487);
xnor U3231 (N_3231,In_602,In_1855);
nor U3232 (N_3232,In_1332,In_424);
and U3233 (N_3233,In_1834,In_586);
or U3234 (N_3234,In_559,In_745);
xnor U3235 (N_3235,In_2035,In_935);
nor U3236 (N_3236,In_1159,In_831);
xnor U3237 (N_3237,In_818,In_1446);
xnor U3238 (N_3238,In_13,In_1552);
nand U3239 (N_3239,In_1800,In_1510);
or U3240 (N_3240,In_141,In_358);
nor U3241 (N_3241,In_2176,In_737);
nand U3242 (N_3242,In_845,In_696);
nor U3243 (N_3243,In_2466,In_2986);
and U3244 (N_3244,In_1820,In_181);
xor U3245 (N_3245,In_830,In_1278);
or U3246 (N_3246,In_93,In_95);
xnor U3247 (N_3247,In_987,In_1041);
or U3248 (N_3248,In_2431,In_1345);
nor U3249 (N_3249,In_2523,In_1100);
and U3250 (N_3250,In_865,In_895);
nand U3251 (N_3251,In_1965,In_1414);
or U3252 (N_3252,In_1250,In_1612);
or U3253 (N_3253,In_1476,In_2402);
nor U3254 (N_3254,In_1026,In_2335);
nor U3255 (N_3255,In_55,In_2217);
xor U3256 (N_3256,In_2989,In_1934);
and U3257 (N_3257,In_2331,In_172);
and U3258 (N_3258,In_285,In_425);
nand U3259 (N_3259,In_1354,In_558);
and U3260 (N_3260,In_2164,In_2410);
xnor U3261 (N_3261,In_1168,In_2981);
xor U3262 (N_3262,In_1199,In_1968);
nor U3263 (N_3263,In_2686,In_1886);
nand U3264 (N_3264,In_1660,In_1845);
or U3265 (N_3265,In_1147,In_1135);
and U3266 (N_3266,In_927,In_2768);
or U3267 (N_3267,In_223,In_1209);
nand U3268 (N_3268,In_3,In_547);
or U3269 (N_3269,In_2691,In_2245);
nor U3270 (N_3270,In_1163,In_1319);
nand U3271 (N_3271,In_230,In_1300);
xnor U3272 (N_3272,In_2366,In_1855);
nor U3273 (N_3273,In_2351,In_2598);
or U3274 (N_3274,In_2046,In_1843);
or U3275 (N_3275,In_890,In_1090);
nor U3276 (N_3276,In_2305,In_1581);
nor U3277 (N_3277,In_363,In_2351);
or U3278 (N_3278,In_2192,In_2024);
and U3279 (N_3279,In_2789,In_2464);
or U3280 (N_3280,In_411,In_1880);
xor U3281 (N_3281,In_74,In_926);
nor U3282 (N_3282,In_485,In_2512);
xor U3283 (N_3283,In_997,In_2794);
or U3284 (N_3284,In_1679,In_1113);
nor U3285 (N_3285,In_1891,In_1601);
nor U3286 (N_3286,In_1453,In_2742);
xnor U3287 (N_3287,In_1971,In_1128);
nand U3288 (N_3288,In_1283,In_1906);
nor U3289 (N_3289,In_1473,In_2552);
nor U3290 (N_3290,In_478,In_1253);
nor U3291 (N_3291,In_1492,In_2169);
nor U3292 (N_3292,In_1152,In_2470);
and U3293 (N_3293,In_649,In_853);
or U3294 (N_3294,In_1133,In_2213);
and U3295 (N_3295,In_1164,In_1918);
nand U3296 (N_3296,In_166,In_2267);
or U3297 (N_3297,In_864,In_228);
nand U3298 (N_3298,In_2185,In_1578);
nand U3299 (N_3299,In_1459,In_1715);
nand U3300 (N_3300,In_2945,In_996);
and U3301 (N_3301,In_1820,In_479);
or U3302 (N_3302,In_2758,In_2900);
and U3303 (N_3303,In_2749,In_2510);
xor U3304 (N_3304,In_2067,In_1693);
nor U3305 (N_3305,In_2114,In_1900);
nor U3306 (N_3306,In_1534,In_1779);
xor U3307 (N_3307,In_523,In_1611);
or U3308 (N_3308,In_2477,In_2103);
and U3309 (N_3309,In_2848,In_1287);
nor U3310 (N_3310,In_1832,In_286);
or U3311 (N_3311,In_1117,In_2148);
nor U3312 (N_3312,In_223,In_270);
nand U3313 (N_3313,In_1240,In_1202);
xor U3314 (N_3314,In_1300,In_2610);
or U3315 (N_3315,In_447,In_202);
and U3316 (N_3316,In_2933,In_2527);
xnor U3317 (N_3317,In_1310,In_1120);
nand U3318 (N_3318,In_75,In_1540);
and U3319 (N_3319,In_353,In_1724);
xnor U3320 (N_3320,In_2616,In_1678);
nor U3321 (N_3321,In_2017,In_783);
xor U3322 (N_3322,In_476,In_1273);
nor U3323 (N_3323,In_936,In_2044);
xnor U3324 (N_3324,In_1634,In_2773);
nor U3325 (N_3325,In_1157,In_400);
xnor U3326 (N_3326,In_2527,In_949);
and U3327 (N_3327,In_1190,In_596);
and U3328 (N_3328,In_2009,In_929);
and U3329 (N_3329,In_1132,In_2446);
and U3330 (N_3330,In_1688,In_2197);
nor U3331 (N_3331,In_1093,In_2138);
nor U3332 (N_3332,In_891,In_2755);
and U3333 (N_3333,In_1347,In_986);
xnor U3334 (N_3334,In_2081,In_240);
xor U3335 (N_3335,In_2112,In_1049);
nor U3336 (N_3336,In_1565,In_861);
nor U3337 (N_3337,In_187,In_2075);
xor U3338 (N_3338,In_2736,In_1672);
and U3339 (N_3339,In_120,In_2685);
nand U3340 (N_3340,In_2336,In_579);
and U3341 (N_3341,In_348,In_915);
and U3342 (N_3342,In_2001,In_2612);
xor U3343 (N_3343,In_2152,In_2927);
nor U3344 (N_3344,In_2070,In_111);
xor U3345 (N_3345,In_2931,In_2452);
or U3346 (N_3346,In_519,In_436);
xnor U3347 (N_3347,In_1329,In_66);
and U3348 (N_3348,In_781,In_1193);
and U3349 (N_3349,In_2562,In_1961);
or U3350 (N_3350,In_801,In_732);
and U3351 (N_3351,In_2379,In_2487);
or U3352 (N_3352,In_1616,In_2242);
nand U3353 (N_3353,In_2407,In_540);
nor U3354 (N_3354,In_2694,In_371);
and U3355 (N_3355,In_1535,In_63);
xnor U3356 (N_3356,In_2315,In_996);
or U3357 (N_3357,In_1717,In_2887);
nand U3358 (N_3358,In_1510,In_1061);
and U3359 (N_3359,In_1927,In_2254);
xnor U3360 (N_3360,In_1575,In_1056);
and U3361 (N_3361,In_2221,In_2124);
or U3362 (N_3362,In_2541,In_210);
or U3363 (N_3363,In_938,In_2874);
and U3364 (N_3364,In_2052,In_59);
xnor U3365 (N_3365,In_1641,In_2300);
or U3366 (N_3366,In_1550,In_1005);
nor U3367 (N_3367,In_2587,In_2858);
nand U3368 (N_3368,In_721,In_558);
xor U3369 (N_3369,In_954,In_2980);
nand U3370 (N_3370,In_478,In_2885);
and U3371 (N_3371,In_1625,In_1009);
xor U3372 (N_3372,In_2845,In_118);
nor U3373 (N_3373,In_641,In_683);
nand U3374 (N_3374,In_1185,In_13);
nand U3375 (N_3375,In_2368,In_2853);
or U3376 (N_3376,In_1469,In_1501);
or U3377 (N_3377,In_827,In_837);
xor U3378 (N_3378,In_757,In_2876);
or U3379 (N_3379,In_2197,In_1338);
nand U3380 (N_3380,In_1566,In_1835);
nor U3381 (N_3381,In_2795,In_1279);
xor U3382 (N_3382,In_618,In_2592);
and U3383 (N_3383,In_220,In_2556);
and U3384 (N_3384,In_1044,In_1014);
or U3385 (N_3385,In_670,In_1661);
nor U3386 (N_3386,In_196,In_619);
and U3387 (N_3387,In_2815,In_1341);
or U3388 (N_3388,In_1194,In_426);
nor U3389 (N_3389,In_1358,In_1948);
nand U3390 (N_3390,In_1609,In_1543);
nand U3391 (N_3391,In_2527,In_1642);
nand U3392 (N_3392,In_1820,In_224);
nor U3393 (N_3393,In_2772,In_123);
or U3394 (N_3394,In_2117,In_2101);
or U3395 (N_3395,In_2080,In_706);
and U3396 (N_3396,In_1852,In_429);
xnor U3397 (N_3397,In_2684,In_718);
or U3398 (N_3398,In_1094,In_1274);
or U3399 (N_3399,In_2090,In_2543);
nor U3400 (N_3400,In_950,In_270);
nand U3401 (N_3401,In_405,In_594);
and U3402 (N_3402,In_2455,In_2972);
or U3403 (N_3403,In_2005,In_2061);
and U3404 (N_3404,In_610,In_1292);
nand U3405 (N_3405,In_732,In_717);
nor U3406 (N_3406,In_2322,In_713);
xnor U3407 (N_3407,In_2766,In_233);
nand U3408 (N_3408,In_1229,In_2735);
xor U3409 (N_3409,In_865,In_2924);
nand U3410 (N_3410,In_2234,In_377);
nor U3411 (N_3411,In_1721,In_491);
and U3412 (N_3412,In_195,In_614);
and U3413 (N_3413,In_1411,In_2566);
nand U3414 (N_3414,In_1897,In_1285);
xor U3415 (N_3415,In_510,In_865);
and U3416 (N_3416,In_1167,In_1261);
nor U3417 (N_3417,In_2251,In_749);
nor U3418 (N_3418,In_531,In_1469);
xnor U3419 (N_3419,In_1020,In_661);
nand U3420 (N_3420,In_182,In_2355);
and U3421 (N_3421,In_1972,In_2317);
and U3422 (N_3422,In_2568,In_2236);
xnor U3423 (N_3423,In_2299,In_1961);
nand U3424 (N_3424,In_1774,In_1234);
xor U3425 (N_3425,In_2696,In_1818);
and U3426 (N_3426,In_1375,In_883);
nand U3427 (N_3427,In_291,In_13);
and U3428 (N_3428,In_619,In_1478);
nand U3429 (N_3429,In_2543,In_31);
nand U3430 (N_3430,In_2920,In_717);
nand U3431 (N_3431,In_290,In_1488);
nor U3432 (N_3432,In_2562,In_983);
nand U3433 (N_3433,In_0,In_2422);
nor U3434 (N_3434,In_359,In_2510);
and U3435 (N_3435,In_1800,In_2943);
nand U3436 (N_3436,In_185,In_472);
xnor U3437 (N_3437,In_2422,In_1873);
nor U3438 (N_3438,In_254,In_1224);
xor U3439 (N_3439,In_300,In_2469);
or U3440 (N_3440,In_2313,In_1403);
nor U3441 (N_3441,In_1468,In_2850);
xnor U3442 (N_3442,In_494,In_93);
xnor U3443 (N_3443,In_2959,In_1438);
nor U3444 (N_3444,In_1840,In_170);
nand U3445 (N_3445,In_568,In_485);
nand U3446 (N_3446,In_2211,In_1888);
or U3447 (N_3447,In_2238,In_1498);
nor U3448 (N_3448,In_742,In_1838);
nand U3449 (N_3449,In_2198,In_2086);
and U3450 (N_3450,In_1437,In_2774);
and U3451 (N_3451,In_2652,In_1442);
nand U3452 (N_3452,In_1980,In_713);
or U3453 (N_3453,In_391,In_1230);
nor U3454 (N_3454,In_1067,In_2807);
and U3455 (N_3455,In_966,In_2023);
and U3456 (N_3456,In_666,In_2687);
nand U3457 (N_3457,In_1802,In_2166);
xnor U3458 (N_3458,In_454,In_1890);
and U3459 (N_3459,In_1474,In_1508);
xnor U3460 (N_3460,In_192,In_2982);
or U3461 (N_3461,In_2177,In_1361);
nand U3462 (N_3462,In_574,In_2473);
nand U3463 (N_3463,In_2448,In_2352);
xnor U3464 (N_3464,In_1802,In_2145);
or U3465 (N_3465,In_412,In_806);
nor U3466 (N_3466,In_2884,In_222);
nor U3467 (N_3467,In_2693,In_259);
xnor U3468 (N_3468,In_1108,In_356);
xnor U3469 (N_3469,In_1748,In_2508);
and U3470 (N_3470,In_2714,In_143);
and U3471 (N_3471,In_493,In_2775);
xor U3472 (N_3472,In_1648,In_1280);
and U3473 (N_3473,In_662,In_2273);
and U3474 (N_3474,In_695,In_1440);
nand U3475 (N_3475,In_142,In_2811);
and U3476 (N_3476,In_2870,In_1897);
nand U3477 (N_3477,In_936,In_186);
xor U3478 (N_3478,In_2211,In_70);
nor U3479 (N_3479,In_959,In_1194);
or U3480 (N_3480,In_760,In_2851);
xor U3481 (N_3481,In_492,In_1618);
or U3482 (N_3482,In_2897,In_2629);
nor U3483 (N_3483,In_1554,In_52);
xor U3484 (N_3484,In_2761,In_2419);
or U3485 (N_3485,In_1005,In_638);
or U3486 (N_3486,In_145,In_233);
nand U3487 (N_3487,In_506,In_518);
xnor U3488 (N_3488,In_1748,In_2671);
nand U3489 (N_3489,In_1109,In_863);
or U3490 (N_3490,In_426,In_2340);
or U3491 (N_3491,In_1243,In_464);
and U3492 (N_3492,In_163,In_114);
nor U3493 (N_3493,In_974,In_1879);
and U3494 (N_3494,In_124,In_1037);
nand U3495 (N_3495,In_1792,In_178);
xor U3496 (N_3496,In_2895,In_1855);
and U3497 (N_3497,In_2120,In_213);
xor U3498 (N_3498,In_467,In_2845);
xor U3499 (N_3499,In_2791,In_1680);
and U3500 (N_3500,In_2316,In_708);
xor U3501 (N_3501,In_335,In_1773);
xor U3502 (N_3502,In_557,In_357);
nor U3503 (N_3503,In_2491,In_1547);
and U3504 (N_3504,In_2871,In_2956);
and U3505 (N_3505,In_1348,In_1159);
and U3506 (N_3506,In_1386,In_1273);
and U3507 (N_3507,In_470,In_2020);
and U3508 (N_3508,In_1546,In_430);
nand U3509 (N_3509,In_27,In_420);
and U3510 (N_3510,In_2829,In_944);
and U3511 (N_3511,In_1160,In_1914);
xor U3512 (N_3512,In_2500,In_1148);
nor U3513 (N_3513,In_2590,In_2411);
nor U3514 (N_3514,In_1785,In_75);
and U3515 (N_3515,In_7,In_1799);
or U3516 (N_3516,In_2789,In_1030);
nor U3517 (N_3517,In_1269,In_644);
nor U3518 (N_3518,In_1042,In_1579);
or U3519 (N_3519,In_95,In_2514);
xor U3520 (N_3520,In_354,In_469);
nand U3521 (N_3521,In_1586,In_1711);
nor U3522 (N_3522,In_1478,In_74);
and U3523 (N_3523,In_2670,In_517);
xor U3524 (N_3524,In_265,In_2176);
and U3525 (N_3525,In_327,In_2663);
nand U3526 (N_3526,In_2278,In_1475);
and U3527 (N_3527,In_2242,In_2663);
xor U3528 (N_3528,In_909,In_1866);
xnor U3529 (N_3529,In_2707,In_1808);
nand U3530 (N_3530,In_2997,In_1626);
xor U3531 (N_3531,In_1491,In_17);
xnor U3532 (N_3532,In_1253,In_1377);
nand U3533 (N_3533,In_1375,In_1110);
and U3534 (N_3534,In_860,In_308);
xor U3535 (N_3535,In_1786,In_911);
and U3536 (N_3536,In_1615,In_1088);
nand U3537 (N_3537,In_2757,In_1172);
and U3538 (N_3538,In_1291,In_2661);
or U3539 (N_3539,In_559,In_1995);
nor U3540 (N_3540,In_1239,In_2978);
xnor U3541 (N_3541,In_1782,In_2949);
or U3542 (N_3542,In_1245,In_2774);
or U3543 (N_3543,In_388,In_346);
or U3544 (N_3544,In_567,In_2271);
nor U3545 (N_3545,In_2059,In_2102);
or U3546 (N_3546,In_1088,In_2443);
or U3547 (N_3547,In_2456,In_65);
and U3548 (N_3548,In_1545,In_2850);
or U3549 (N_3549,In_2863,In_2726);
nand U3550 (N_3550,In_680,In_1020);
or U3551 (N_3551,In_341,In_603);
nand U3552 (N_3552,In_498,In_905);
and U3553 (N_3553,In_322,In_2260);
nand U3554 (N_3554,In_960,In_918);
nand U3555 (N_3555,In_1065,In_2397);
xor U3556 (N_3556,In_2628,In_1229);
nor U3557 (N_3557,In_2338,In_329);
or U3558 (N_3558,In_1835,In_2901);
xnor U3559 (N_3559,In_2046,In_419);
and U3560 (N_3560,In_1889,In_260);
and U3561 (N_3561,In_491,In_359);
xnor U3562 (N_3562,In_376,In_2305);
nor U3563 (N_3563,In_16,In_2150);
xnor U3564 (N_3564,In_1468,In_2112);
nor U3565 (N_3565,In_2232,In_2475);
or U3566 (N_3566,In_1803,In_1189);
and U3567 (N_3567,In_369,In_823);
xnor U3568 (N_3568,In_541,In_2924);
and U3569 (N_3569,In_422,In_154);
and U3570 (N_3570,In_2456,In_2144);
or U3571 (N_3571,In_621,In_677);
nor U3572 (N_3572,In_169,In_419);
or U3573 (N_3573,In_235,In_1733);
nor U3574 (N_3574,In_729,In_2173);
or U3575 (N_3575,In_2391,In_607);
nor U3576 (N_3576,In_121,In_852);
nor U3577 (N_3577,In_1239,In_63);
or U3578 (N_3578,In_2213,In_2774);
xnor U3579 (N_3579,In_371,In_812);
and U3580 (N_3580,In_747,In_2015);
xor U3581 (N_3581,In_2638,In_2953);
nand U3582 (N_3582,In_515,In_1737);
nand U3583 (N_3583,In_2816,In_1152);
and U3584 (N_3584,In_1477,In_427);
xor U3585 (N_3585,In_1982,In_508);
nand U3586 (N_3586,In_2338,In_2861);
nor U3587 (N_3587,In_2824,In_1186);
xor U3588 (N_3588,In_2133,In_1815);
or U3589 (N_3589,In_345,In_117);
nor U3590 (N_3590,In_1112,In_2459);
nand U3591 (N_3591,In_588,In_955);
or U3592 (N_3592,In_2678,In_2619);
xnor U3593 (N_3593,In_879,In_1754);
nor U3594 (N_3594,In_2114,In_1123);
nand U3595 (N_3595,In_341,In_1438);
xor U3596 (N_3596,In_2849,In_942);
nand U3597 (N_3597,In_58,In_1714);
nor U3598 (N_3598,In_2959,In_2900);
nand U3599 (N_3599,In_2282,In_1720);
xor U3600 (N_3600,In_2553,In_45);
or U3601 (N_3601,In_2549,In_1399);
or U3602 (N_3602,In_2389,In_1867);
or U3603 (N_3603,In_1654,In_1026);
nor U3604 (N_3604,In_2490,In_547);
xnor U3605 (N_3605,In_1474,In_2703);
nand U3606 (N_3606,In_1936,In_1152);
and U3607 (N_3607,In_392,In_42);
nor U3608 (N_3608,In_1825,In_1683);
or U3609 (N_3609,In_2513,In_2300);
or U3610 (N_3610,In_1602,In_610);
and U3611 (N_3611,In_2552,In_2928);
xor U3612 (N_3612,In_1143,In_1999);
or U3613 (N_3613,In_2105,In_759);
or U3614 (N_3614,In_1556,In_2079);
or U3615 (N_3615,In_1727,In_1224);
xnor U3616 (N_3616,In_382,In_1178);
nand U3617 (N_3617,In_1996,In_411);
or U3618 (N_3618,In_525,In_1836);
nand U3619 (N_3619,In_2525,In_2906);
or U3620 (N_3620,In_2056,In_1652);
and U3621 (N_3621,In_2718,In_1682);
nand U3622 (N_3622,In_2381,In_345);
nor U3623 (N_3623,In_1633,In_1274);
nand U3624 (N_3624,In_2340,In_264);
or U3625 (N_3625,In_2945,In_619);
or U3626 (N_3626,In_1893,In_2229);
or U3627 (N_3627,In_402,In_2925);
nand U3628 (N_3628,In_778,In_2190);
and U3629 (N_3629,In_823,In_229);
xnor U3630 (N_3630,In_127,In_1651);
nand U3631 (N_3631,In_1883,In_2451);
nor U3632 (N_3632,In_2522,In_832);
nor U3633 (N_3633,In_750,In_736);
nand U3634 (N_3634,In_2556,In_483);
and U3635 (N_3635,In_1104,In_2876);
and U3636 (N_3636,In_2100,In_2083);
or U3637 (N_3637,In_2662,In_672);
or U3638 (N_3638,In_277,In_861);
xnor U3639 (N_3639,In_2071,In_355);
or U3640 (N_3640,In_465,In_1294);
and U3641 (N_3641,In_908,In_187);
nand U3642 (N_3642,In_1543,In_906);
nand U3643 (N_3643,In_1600,In_1242);
xnor U3644 (N_3644,In_362,In_324);
or U3645 (N_3645,In_2015,In_733);
nor U3646 (N_3646,In_397,In_1428);
nor U3647 (N_3647,In_2191,In_1822);
nor U3648 (N_3648,In_1622,In_470);
and U3649 (N_3649,In_1796,In_2405);
xnor U3650 (N_3650,In_1026,In_832);
nor U3651 (N_3651,In_1405,In_1619);
nand U3652 (N_3652,In_134,In_2923);
nand U3653 (N_3653,In_1217,In_2418);
xnor U3654 (N_3654,In_2988,In_688);
xnor U3655 (N_3655,In_560,In_398);
or U3656 (N_3656,In_2676,In_2366);
or U3657 (N_3657,In_2295,In_973);
and U3658 (N_3658,In_80,In_2355);
or U3659 (N_3659,In_354,In_2753);
nor U3660 (N_3660,In_2106,In_2552);
nand U3661 (N_3661,In_1743,In_2501);
and U3662 (N_3662,In_1629,In_597);
or U3663 (N_3663,In_1990,In_1364);
nor U3664 (N_3664,In_2287,In_740);
nor U3665 (N_3665,In_1938,In_425);
and U3666 (N_3666,In_432,In_248);
xnor U3667 (N_3667,In_2846,In_283);
nand U3668 (N_3668,In_1537,In_954);
or U3669 (N_3669,In_670,In_2000);
xor U3670 (N_3670,In_2314,In_1291);
nand U3671 (N_3671,In_2558,In_1314);
and U3672 (N_3672,In_990,In_172);
nor U3673 (N_3673,In_1469,In_1836);
or U3674 (N_3674,In_245,In_471);
and U3675 (N_3675,In_2641,In_421);
xor U3676 (N_3676,In_886,In_249);
or U3677 (N_3677,In_2403,In_845);
nor U3678 (N_3678,In_129,In_2127);
or U3679 (N_3679,In_2292,In_2148);
nand U3680 (N_3680,In_524,In_63);
nor U3681 (N_3681,In_2300,In_358);
nand U3682 (N_3682,In_496,In_174);
or U3683 (N_3683,In_1967,In_2012);
xor U3684 (N_3684,In_1777,In_837);
nor U3685 (N_3685,In_1844,In_2038);
and U3686 (N_3686,In_2459,In_823);
and U3687 (N_3687,In_140,In_2520);
xnor U3688 (N_3688,In_2071,In_1304);
nand U3689 (N_3689,In_1125,In_447);
nand U3690 (N_3690,In_2637,In_654);
xnor U3691 (N_3691,In_111,In_454);
or U3692 (N_3692,In_228,In_2121);
and U3693 (N_3693,In_246,In_1367);
nor U3694 (N_3694,In_2006,In_2338);
nand U3695 (N_3695,In_1604,In_390);
nor U3696 (N_3696,In_1841,In_220);
and U3697 (N_3697,In_602,In_2858);
xor U3698 (N_3698,In_54,In_2429);
nor U3699 (N_3699,In_2493,In_884);
nand U3700 (N_3700,In_779,In_1646);
xor U3701 (N_3701,In_2131,In_1274);
nand U3702 (N_3702,In_1336,In_1851);
or U3703 (N_3703,In_1614,In_2335);
or U3704 (N_3704,In_688,In_1065);
xnor U3705 (N_3705,In_1514,In_2367);
or U3706 (N_3706,In_2818,In_210);
and U3707 (N_3707,In_2819,In_1806);
and U3708 (N_3708,In_2651,In_974);
nand U3709 (N_3709,In_1139,In_519);
xor U3710 (N_3710,In_61,In_734);
or U3711 (N_3711,In_903,In_2869);
or U3712 (N_3712,In_1412,In_1035);
nand U3713 (N_3713,In_2564,In_2800);
nand U3714 (N_3714,In_1257,In_1342);
nand U3715 (N_3715,In_2222,In_2894);
xnor U3716 (N_3716,In_1472,In_944);
and U3717 (N_3717,In_671,In_1124);
nor U3718 (N_3718,In_702,In_41);
nor U3719 (N_3719,In_382,In_1511);
nand U3720 (N_3720,In_1778,In_400);
nor U3721 (N_3721,In_857,In_2214);
or U3722 (N_3722,In_2848,In_771);
nand U3723 (N_3723,In_1984,In_1702);
xor U3724 (N_3724,In_393,In_2202);
or U3725 (N_3725,In_1840,In_1375);
nand U3726 (N_3726,In_654,In_2880);
or U3727 (N_3727,In_2094,In_2276);
and U3728 (N_3728,In_2998,In_2909);
nor U3729 (N_3729,In_619,In_690);
xor U3730 (N_3730,In_1477,In_270);
and U3731 (N_3731,In_1715,In_2375);
or U3732 (N_3732,In_1839,In_1541);
and U3733 (N_3733,In_937,In_1709);
nor U3734 (N_3734,In_1772,In_1220);
nor U3735 (N_3735,In_2898,In_763);
nand U3736 (N_3736,In_1724,In_94);
xnor U3737 (N_3737,In_1745,In_1096);
and U3738 (N_3738,In_2536,In_2680);
nor U3739 (N_3739,In_1384,In_444);
nand U3740 (N_3740,In_1526,In_2788);
and U3741 (N_3741,In_2488,In_1134);
xnor U3742 (N_3742,In_112,In_2191);
or U3743 (N_3743,In_1248,In_2519);
and U3744 (N_3744,In_1362,In_2514);
nand U3745 (N_3745,In_153,In_376);
and U3746 (N_3746,In_1200,In_1845);
nor U3747 (N_3747,In_587,In_2755);
nand U3748 (N_3748,In_2357,In_1960);
xnor U3749 (N_3749,In_841,In_2479);
nand U3750 (N_3750,In_2881,In_781);
and U3751 (N_3751,In_2991,In_1905);
nand U3752 (N_3752,In_2521,In_230);
nor U3753 (N_3753,In_2691,In_1032);
xnor U3754 (N_3754,In_888,In_2064);
and U3755 (N_3755,In_2086,In_815);
xnor U3756 (N_3756,In_613,In_1131);
nor U3757 (N_3757,In_999,In_1428);
xnor U3758 (N_3758,In_2681,In_2221);
and U3759 (N_3759,In_1468,In_1520);
and U3760 (N_3760,In_658,In_277);
and U3761 (N_3761,In_1782,In_1394);
and U3762 (N_3762,In_1734,In_2418);
or U3763 (N_3763,In_1247,In_1751);
nor U3764 (N_3764,In_1223,In_36);
nand U3765 (N_3765,In_840,In_1959);
or U3766 (N_3766,In_2860,In_777);
nor U3767 (N_3767,In_343,In_2190);
or U3768 (N_3768,In_1601,In_290);
or U3769 (N_3769,In_1731,In_2844);
xor U3770 (N_3770,In_78,In_2471);
or U3771 (N_3771,In_2942,In_1132);
nor U3772 (N_3772,In_780,In_458);
or U3773 (N_3773,In_1772,In_2555);
xor U3774 (N_3774,In_1315,In_419);
nor U3775 (N_3775,In_90,In_893);
nand U3776 (N_3776,In_1990,In_264);
or U3777 (N_3777,In_1250,In_909);
nor U3778 (N_3778,In_2790,In_1696);
nand U3779 (N_3779,In_1694,In_211);
nand U3780 (N_3780,In_91,In_2438);
and U3781 (N_3781,In_201,In_650);
nand U3782 (N_3782,In_2087,In_620);
nand U3783 (N_3783,In_499,In_924);
nor U3784 (N_3784,In_2825,In_2770);
or U3785 (N_3785,In_2910,In_247);
xnor U3786 (N_3786,In_2217,In_1388);
or U3787 (N_3787,In_376,In_1290);
and U3788 (N_3788,In_977,In_2816);
nand U3789 (N_3789,In_1345,In_2943);
and U3790 (N_3790,In_2872,In_2858);
nand U3791 (N_3791,In_498,In_2967);
or U3792 (N_3792,In_951,In_2995);
xnor U3793 (N_3793,In_465,In_1425);
nand U3794 (N_3794,In_2506,In_1795);
nand U3795 (N_3795,In_2625,In_1060);
xor U3796 (N_3796,In_168,In_2201);
or U3797 (N_3797,In_1117,In_2656);
nor U3798 (N_3798,In_2882,In_2689);
nand U3799 (N_3799,In_1774,In_2159);
or U3800 (N_3800,In_23,In_17);
or U3801 (N_3801,In_1868,In_2381);
nor U3802 (N_3802,In_633,In_138);
xor U3803 (N_3803,In_2201,In_792);
or U3804 (N_3804,In_2099,In_2642);
and U3805 (N_3805,In_399,In_1733);
nor U3806 (N_3806,In_127,In_2535);
or U3807 (N_3807,In_2903,In_1939);
nor U3808 (N_3808,In_2284,In_2997);
nand U3809 (N_3809,In_1152,In_2611);
and U3810 (N_3810,In_2714,In_168);
xnor U3811 (N_3811,In_2503,In_1782);
nor U3812 (N_3812,In_1330,In_533);
nand U3813 (N_3813,In_1000,In_2173);
or U3814 (N_3814,In_10,In_2597);
nor U3815 (N_3815,In_1882,In_640);
nor U3816 (N_3816,In_2090,In_2874);
and U3817 (N_3817,In_2563,In_680);
nor U3818 (N_3818,In_1445,In_1565);
nand U3819 (N_3819,In_1300,In_1055);
and U3820 (N_3820,In_2642,In_472);
or U3821 (N_3821,In_1781,In_2866);
or U3822 (N_3822,In_1320,In_2304);
nand U3823 (N_3823,In_189,In_464);
nand U3824 (N_3824,In_39,In_1387);
and U3825 (N_3825,In_2689,In_621);
nand U3826 (N_3826,In_1138,In_2079);
nand U3827 (N_3827,In_2951,In_483);
nand U3828 (N_3828,In_2319,In_9);
and U3829 (N_3829,In_1403,In_2438);
nand U3830 (N_3830,In_808,In_653);
xor U3831 (N_3831,In_1839,In_1594);
or U3832 (N_3832,In_295,In_2171);
or U3833 (N_3833,In_2886,In_736);
nor U3834 (N_3834,In_1870,In_1119);
nor U3835 (N_3835,In_169,In_825);
nand U3836 (N_3836,In_1233,In_2903);
or U3837 (N_3837,In_2328,In_1076);
nand U3838 (N_3838,In_1953,In_791);
xor U3839 (N_3839,In_2482,In_584);
nand U3840 (N_3840,In_1029,In_2180);
and U3841 (N_3841,In_1788,In_1892);
xnor U3842 (N_3842,In_1966,In_2406);
or U3843 (N_3843,In_1260,In_691);
or U3844 (N_3844,In_1660,In_1126);
and U3845 (N_3845,In_309,In_833);
xnor U3846 (N_3846,In_2798,In_2950);
nor U3847 (N_3847,In_1786,In_150);
nand U3848 (N_3848,In_2912,In_1241);
nand U3849 (N_3849,In_1943,In_1112);
or U3850 (N_3850,In_955,In_2915);
nand U3851 (N_3851,In_2741,In_1643);
and U3852 (N_3852,In_781,In_2412);
nor U3853 (N_3853,In_96,In_357);
or U3854 (N_3854,In_1343,In_2352);
nor U3855 (N_3855,In_954,In_1914);
xor U3856 (N_3856,In_1988,In_1093);
nor U3857 (N_3857,In_630,In_1719);
nand U3858 (N_3858,In_1667,In_976);
and U3859 (N_3859,In_144,In_279);
or U3860 (N_3860,In_135,In_1911);
nor U3861 (N_3861,In_2576,In_1063);
nand U3862 (N_3862,In_2018,In_2967);
nand U3863 (N_3863,In_100,In_1771);
nor U3864 (N_3864,In_2727,In_1384);
and U3865 (N_3865,In_1810,In_2734);
xnor U3866 (N_3866,In_2907,In_2884);
and U3867 (N_3867,In_2189,In_653);
xor U3868 (N_3868,In_1610,In_2445);
or U3869 (N_3869,In_2844,In_1459);
xor U3870 (N_3870,In_2159,In_1803);
nor U3871 (N_3871,In_1352,In_1719);
nand U3872 (N_3872,In_503,In_1429);
nand U3873 (N_3873,In_1650,In_2479);
and U3874 (N_3874,In_2532,In_2864);
xor U3875 (N_3875,In_739,In_1050);
xnor U3876 (N_3876,In_1362,In_1706);
nand U3877 (N_3877,In_2496,In_1263);
or U3878 (N_3878,In_2748,In_2108);
xor U3879 (N_3879,In_623,In_2480);
xnor U3880 (N_3880,In_881,In_1231);
or U3881 (N_3881,In_133,In_761);
nor U3882 (N_3882,In_291,In_1261);
and U3883 (N_3883,In_593,In_1549);
or U3884 (N_3884,In_127,In_522);
or U3885 (N_3885,In_2734,In_383);
xor U3886 (N_3886,In_327,In_1140);
nor U3887 (N_3887,In_2191,In_1976);
and U3888 (N_3888,In_115,In_1424);
and U3889 (N_3889,In_584,In_1985);
or U3890 (N_3890,In_1082,In_1881);
or U3891 (N_3891,In_1680,In_1829);
or U3892 (N_3892,In_1359,In_2958);
nor U3893 (N_3893,In_2244,In_1647);
nor U3894 (N_3894,In_1465,In_288);
and U3895 (N_3895,In_1908,In_635);
or U3896 (N_3896,In_194,In_255);
and U3897 (N_3897,In_2125,In_2606);
xor U3898 (N_3898,In_877,In_173);
or U3899 (N_3899,In_2119,In_796);
nor U3900 (N_3900,In_2621,In_1285);
xor U3901 (N_3901,In_2685,In_1499);
and U3902 (N_3902,In_2880,In_2720);
nand U3903 (N_3903,In_2156,In_546);
nand U3904 (N_3904,In_512,In_19);
nor U3905 (N_3905,In_1456,In_1444);
xor U3906 (N_3906,In_1104,In_2295);
nand U3907 (N_3907,In_1625,In_287);
nand U3908 (N_3908,In_122,In_1690);
xor U3909 (N_3909,In_535,In_719);
nor U3910 (N_3910,In_330,In_772);
nor U3911 (N_3911,In_1314,In_44);
and U3912 (N_3912,In_2704,In_422);
nand U3913 (N_3913,In_2197,In_2878);
and U3914 (N_3914,In_770,In_963);
xor U3915 (N_3915,In_1464,In_387);
nor U3916 (N_3916,In_1827,In_845);
nor U3917 (N_3917,In_2806,In_55);
and U3918 (N_3918,In_2266,In_1244);
or U3919 (N_3919,In_2840,In_2650);
nor U3920 (N_3920,In_126,In_1584);
nor U3921 (N_3921,In_300,In_961);
xnor U3922 (N_3922,In_916,In_2280);
or U3923 (N_3923,In_287,In_268);
nand U3924 (N_3924,In_743,In_604);
xnor U3925 (N_3925,In_2298,In_381);
and U3926 (N_3926,In_1455,In_2335);
nand U3927 (N_3927,In_908,In_2601);
or U3928 (N_3928,In_2037,In_1216);
nand U3929 (N_3929,In_537,In_2153);
and U3930 (N_3930,In_2948,In_2357);
or U3931 (N_3931,In_1485,In_1807);
nor U3932 (N_3932,In_548,In_1223);
nor U3933 (N_3933,In_1507,In_2221);
nor U3934 (N_3934,In_2039,In_873);
nor U3935 (N_3935,In_2227,In_1609);
nand U3936 (N_3936,In_2259,In_1043);
xor U3937 (N_3937,In_563,In_1684);
xor U3938 (N_3938,In_2822,In_630);
nand U3939 (N_3939,In_2508,In_232);
nor U3940 (N_3940,In_1548,In_1124);
nor U3941 (N_3941,In_2032,In_1698);
nor U3942 (N_3942,In_1504,In_967);
or U3943 (N_3943,In_1781,In_145);
nand U3944 (N_3944,In_1785,In_282);
and U3945 (N_3945,In_2440,In_1494);
nor U3946 (N_3946,In_2362,In_1209);
and U3947 (N_3947,In_2411,In_1771);
nand U3948 (N_3948,In_1730,In_2784);
nand U3949 (N_3949,In_510,In_2421);
or U3950 (N_3950,In_959,In_2522);
xor U3951 (N_3951,In_1528,In_112);
and U3952 (N_3952,In_212,In_2198);
xnor U3953 (N_3953,In_2097,In_1717);
xnor U3954 (N_3954,In_2304,In_1257);
nand U3955 (N_3955,In_1632,In_980);
or U3956 (N_3956,In_1692,In_884);
or U3957 (N_3957,In_2430,In_2036);
nand U3958 (N_3958,In_956,In_1088);
nand U3959 (N_3959,In_506,In_1641);
nor U3960 (N_3960,In_1655,In_1388);
or U3961 (N_3961,In_1344,In_2755);
and U3962 (N_3962,In_2766,In_2375);
and U3963 (N_3963,In_1525,In_671);
xnor U3964 (N_3964,In_1487,In_1937);
xnor U3965 (N_3965,In_2606,In_2447);
nor U3966 (N_3966,In_610,In_322);
and U3967 (N_3967,In_2217,In_1123);
xnor U3968 (N_3968,In_627,In_587);
xnor U3969 (N_3969,In_638,In_2222);
and U3970 (N_3970,In_946,In_1393);
and U3971 (N_3971,In_2306,In_1099);
xnor U3972 (N_3972,In_402,In_715);
or U3973 (N_3973,In_1737,In_2696);
and U3974 (N_3974,In_1822,In_2284);
or U3975 (N_3975,In_2718,In_89);
or U3976 (N_3976,In_1239,In_1411);
xor U3977 (N_3977,In_1671,In_262);
nor U3978 (N_3978,In_1884,In_2472);
nand U3979 (N_3979,In_418,In_2410);
xnor U3980 (N_3980,In_1815,In_316);
or U3981 (N_3981,In_758,In_1568);
xnor U3982 (N_3982,In_1225,In_2662);
and U3983 (N_3983,In_1183,In_175);
xor U3984 (N_3984,In_205,In_2398);
nand U3985 (N_3985,In_2558,In_1611);
nand U3986 (N_3986,In_446,In_817);
xnor U3987 (N_3987,In_534,In_278);
nand U3988 (N_3988,In_432,In_696);
nor U3989 (N_3989,In_779,In_382);
or U3990 (N_3990,In_1611,In_1734);
or U3991 (N_3991,In_495,In_1711);
nand U3992 (N_3992,In_615,In_2630);
or U3993 (N_3993,In_2254,In_201);
and U3994 (N_3994,In_2670,In_1118);
xnor U3995 (N_3995,In_529,In_1754);
nor U3996 (N_3996,In_891,In_1320);
nor U3997 (N_3997,In_2053,In_79);
nand U3998 (N_3998,In_1782,In_1400);
xnor U3999 (N_3999,In_1918,In_2243);
or U4000 (N_4000,In_55,In_194);
nand U4001 (N_4001,In_2701,In_2515);
nor U4002 (N_4002,In_186,In_197);
nor U4003 (N_4003,In_229,In_175);
xnor U4004 (N_4004,In_428,In_1241);
and U4005 (N_4005,In_548,In_951);
and U4006 (N_4006,In_2047,In_2528);
nand U4007 (N_4007,In_1385,In_2851);
nor U4008 (N_4008,In_2120,In_1306);
nor U4009 (N_4009,In_2449,In_2865);
and U4010 (N_4010,In_1619,In_236);
or U4011 (N_4011,In_1291,In_1941);
nand U4012 (N_4012,In_1943,In_1214);
nor U4013 (N_4013,In_783,In_616);
xnor U4014 (N_4014,In_1535,In_1167);
or U4015 (N_4015,In_2890,In_2769);
xnor U4016 (N_4016,In_1588,In_1805);
nand U4017 (N_4017,In_2887,In_1895);
and U4018 (N_4018,In_2951,In_302);
or U4019 (N_4019,In_2441,In_867);
or U4020 (N_4020,In_1462,In_1926);
nand U4021 (N_4021,In_1117,In_2009);
nand U4022 (N_4022,In_1819,In_724);
nor U4023 (N_4023,In_887,In_779);
nor U4024 (N_4024,In_746,In_2676);
and U4025 (N_4025,In_1452,In_2205);
or U4026 (N_4026,In_741,In_1435);
or U4027 (N_4027,In_1851,In_437);
xor U4028 (N_4028,In_2760,In_1834);
and U4029 (N_4029,In_2738,In_1895);
or U4030 (N_4030,In_1422,In_1786);
nor U4031 (N_4031,In_430,In_862);
nor U4032 (N_4032,In_1636,In_1312);
or U4033 (N_4033,In_239,In_123);
or U4034 (N_4034,In_1519,In_2353);
nor U4035 (N_4035,In_640,In_2941);
or U4036 (N_4036,In_1285,In_1488);
xor U4037 (N_4037,In_2338,In_1587);
nor U4038 (N_4038,In_1111,In_194);
nand U4039 (N_4039,In_1197,In_2076);
xor U4040 (N_4040,In_1193,In_1208);
and U4041 (N_4041,In_741,In_1360);
xnor U4042 (N_4042,In_1039,In_1257);
and U4043 (N_4043,In_2804,In_832);
nand U4044 (N_4044,In_2231,In_114);
nor U4045 (N_4045,In_1218,In_1299);
and U4046 (N_4046,In_1269,In_226);
and U4047 (N_4047,In_2365,In_2685);
or U4048 (N_4048,In_134,In_1323);
nor U4049 (N_4049,In_2710,In_442);
nor U4050 (N_4050,In_1878,In_1098);
xnor U4051 (N_4051,In_171,In_669);
or U4052 (N_4052,In_1234,In_2752);
nor U4053 (N_4053,In_2556,In_410);
nand U4054 (N_4054,In_1738,In_1331);
nor U4055 (N_4055,In_2739,In_2127);
nor U4056 (N_4056,In_954,In_2497);
nand U4057 (N_4057,In_1909,In_191);
or U4058 (N_4058,In_2600,In_1504);
or U4059 (N_4059,In_282,In_2502);
and U4060 (N_4060,In_506,In_1950);
or U4061 (N_4061,In_2747,In_1059);
xnor U4062 (N_4062,In_308,In_1267);
and U4063 (N_4063,In_1043,In_1231);
xnor U4064 (N_4064,In_2654,In_1020);
or U4065 (N_4065,In_1237,In_2723);
or U4066 (N_4066,In_1661,In_700);
xnor U4067 (N_4067,In_672,In_1612);
and U4068 (N_4068,In_1367,In_1941);
and U4069 (N_4069,In_181,In_1437);
nor U4070 (N_4070,In_2191,In_25);
nand U4071 (N_4071,In_2115,In_594);
nand U4072 (N_4072,In_932,In_584);
nand U4073 (N_4073,In_2809,In_2513);
nand U4074 (N_4074,In_1844,In_1022);
xnor U4075 (N_4075,In_1850,In_381);
nor U4076 (N_4076,In_586,In_2539);
xor U4077 (N_4077,In_512,In_1199);
nand U4078 (N_4078,In_2802,In_587);
xor U4079 (N_4079,In_570,In_1664);
or U4080 (N_4080,In_291,In_1915);
or U4081 (N_4081,In_2472,In_1833);
xor U4082 (N_4082,In_1870,In_653);
nor U4083 (N_4083,In_1635,In_553);
nor U4084 (N_4084,In_1054,In_2567);
and U4085 (N_4085,In_1650,In_2576);
xnor U4086 (N_4086,In_705,In_473);
or U4087 (N_4087,In_98,In_1300);
nand U4088 (N_4088,In_2127,In_2012);
or U4089 (N_4089,In_2386,In_2802);
nor U4090 (N_4090,In_1638,In_837);
nor U4091 (N_4091,In_2709,In_1740);
nand U4092 (N_4092,In_63,In_1707);
nor U4093 (N_4093,In_494,In_2265);
xnor U4094 (N_4094,In_673,In_2338);
nand U4095 (N_4095,In_2571,In_723);
and U4096 (N_4096,In_11,In_1372);
nor U4097 (N_4097,In_2402,In_1208);
and U4098 (N_4098,In_1846,In_1424);
nand U4099 (N_4099,In_727,In_901);
xnor U4100 (N_4100,In_975,In_1357);
and U4101 (N_4101,In_2610,In_60);
nand U4102 (N_4102,In_2506,In_2386);
and U4103 (N_4103,In_957,In_394);
and U4104 (N_4104,In_800,In_450);
nor U4105 (N_4105,In_2136,In_2415);
xnor U4106 (N_4106,In_166,In_2244);
xor U4107 (N_4107,In_2208,In_489);
or U4108 (N_4108,In_500,In_2399);
or U4109 (N_4109,In_309,In_2928);
nand U4110 (N_4110,In_2317,In_2293);
or U4111 (N_4111,In_1134,In_2661);
nand U4112 (N_4112,In_487,In_1751);
or U4113 (N_4113,In_2421,In_2687);
xnor U4114 (N_4114,In_1998,In_1037);
or U4115 (N_4115,In_1599,In_121);
and U4116 (N_4116,In_553,In_2110);
xor U4117 (N_4117,In_2990,In_190);
and U4118 (N_4118,In_2879,In_2153);
nor U4119 (N_4119,In_121,In_2366);
nor U4120 (N_4120,In_823,In_2909);
or U4121 (N_4121,In_1436,In_2189);
nand U4122 (N_4122,In_2375,In_84);
xor U4123 (N_4123,In_2609,In_543);
and U4124 (N_4124,In_2516,In_16);
or U4125 (N_4125,In_1164,In_2796);
nand U4126 (N_4126,In_2686,In_2175);
nor U4127 (N_4127,In_466,In_590);
and U4128 (N_4128,In_934,In_2797);
or U4129 (N_4129,In_2048,In_1021);
or U4130 (N_4130,In_1463,In_806);
and U4131 (N_4131,In_1002,In_2495);
and U4132 (N_4132,In_754,In_1809);
nor U4133 (N_4133,In_2758,In_2578);
nor U4134 (N_4134,In_2501,In_769);
nand U4135 (N_4135,In_2678,In_2874);
and U4136 (N_4136,In_1319,In_2321);
and U4137 (N_4137,In_1378,In_2165);
and U4138 (N_4138,In_227,In_2979);
xor U4139 (N_4139,In_1848,In_2923);
or U4140 (N_4140,In_2819,In_705);
and U4141 (N_4141,In_1975,In_784);
nand U4142 (N_4142,In_2884,In_2401);
nand U4143 (N_4143,In_2442,In_283);
nand U4144 (N_4144,In_2534,In_2562);
nand U4145 (N_4145,In_2417,In_37);
or U4146 (N_4146,In_2372,In_2625);
nor U4147 (N_4147,In_1797,In_78);
xnor U4148 (N_4148,In_180,In_1639);
or U4149 (N_4149,In_2209,In_1479);
xor U4150 (N_4150,In_2367,In_2759);
nand U4151 (N_4151,In_437,In_2227);
nand U4152 (N_4152,In_1105,In_1289);
nand U4153 (N_4153,In_1869,In_2342);
xor U4154 (N_4154,In_2541,In_2802);
or U4155 (N_4155,In_789,In_2813);
nor U4156 (N_4156,In_237,In_1411);
or U4157 (N_4157,In_286,In_147);
xnor U4158 (N_4158,In_2524,In_2570);
nand U4159 (N_4159,In_768,In_2923);
xnor U4160 (N_4160,In_67,In_1081);
nand U4161 (N_4161,In_154,In_551);
nand U4162 (N_4162,In_2992,In_914);
nand U4163 (N_4163,In_1903,In_2518);
nand U4164 (N_4164,In_637,In_1769);
and U4165 (N_4165,In_306,In_2989);
xor U4166 (N_4166,In_2129,In_2500);
nor U4167 (N_4167,In_142,In_2346);
nor U4168 (N_4168,In_1134,In_5);
nor U4169 (N_4169,In_2761,In_2153);
xnor U4170 (N_4170,In_2494,In_1690);
and U4171 (N_4171,In_1292,In_1811);
and U4172 (N_4172,In_2268,In_1901);
and U4173 (N_4173,In_1789,In_500);
and U4174 (N_4174,In_1159,In_2643);
or U4175 (N_4175,In_46,In_230);
nand U4176 (N_4176,In_449,In_915);
xnor U4177 (N_4177,In_578,In_2540);
xnor U4178 (N_4178,In_1625,In_1032);
or U4179 (N_4179,In_1326,In_2776);
and U4180 (N_4180,In_2024,In_2380);
and U4181 (N_4181,In_163,In_1251);
nor U4182 (N_4182,In_688,In_2354);
nand U4183 (N_4183,In_2613,In_2152);
and U4184 (N_4184,In_1620,In_632);
and U4185 (N_4185,In_2795,In_918);
or U4186 (N_4186,In_1220,In_410);
and U4187 (N_4187,In_2560,In_956);
nand U4188 (N_4188,In_659,In_2317);
nand U4189 (N_4189,In_1492,In_2638);
nor U4190 (N_4190,In_1303,In_24);
and U4191 (N_4191,In_627,In_2106);
nor U4192 (N_4192,In_1553,In_488);
nor U4193 (N_4193,In_2410,In_2048);
nor U4194 (N_4194,In_2110,In_2400);
nor U4195 (N_4195,In_1340,In_477);
or U4196 (N_4196,In_2588,In_36);
nor U4197 (N_4197,In_1177,In_1820);
nand U4198 (N_4198,In_1601,In_2366);
xnor U4199 (N_4199,In_2040,In_1843);
and U4200 (N_4200,In_2064,In_788);
and U4201 (N_4201,In_1393,In_1207);
or U4202 (N_4202,In_1584,In_2317);
nor U4203 (N_4203,In_353,In_2874);
nor U4204 (N_4204,In_2463,In_2704);
or U4205 (N_4205,In_1963,In_424);
xnor U4206 (N_4206,In_2390,In_598);
nor U4207 (N_4207,In_1429,In_220);
and U4208 (N_4208,In_2015,In_1618);
or U4209 (N_4209,In_2071,In_1658);
and U4210 (N_4210,In_2265,In_1972);
nand U4211 (N_4211,In_4,In_2362);
or U4212 (N_4212,In_826,In_1217);
xnor U4213 (N_4213,In_893,In_1070);
xnor U4214 (N_4214,In_142,In_2937);
nor U4215 (N_4215,In_1231,In_1915);
nand U4216 (N_4216,In_838,In_2734);
and U4217 (N_4217,In_99,In_1271);
xnor U4218 (N_4218,In_1258,In_2597);
or U4219 (N_4219,In_2327,In_2107);
nand U4220 (N_4220,In_1060,In_954);
nand U4221 (N_4221,In_2925,In_2366);
nand U4222 (N_4222,In_1212,In_175);
or U4223 (N_4223,In_2470,In_791);
nand U4224 (N_4224,In_79,In_170);
xor U4225 (N_4225,In_1270,In_1128);
or U4226 (N_4226,In_398,In_1945);
or U4227 (N_4227,In_917,In_2165);
or U4228 (N_4228,In_564,In_1558);
or U4229 (N_4229,In_2248,In_724);
and U4230 (N_4230,In_1745,In_1428);
xor U4231 (N_4231,In_1446,In_2629);
and U4232 (N_4232,In_2949,In_743);
and U4233 (N_4233,In_1544,In_2604);
or U4234 (N_4234,In_207,In_1703);
xnor U4235 (N_4235,In_312,In_825);
or U4236 (N_4236,In_2675,In_2732);
xor U4237 (N_4237,In_2341,In_1467);
nor U4238 (N_4238,In_992,In_2112);
xor U4239 (N_4239,In_96,In_801);
or U4240 (N_4240,In_1990,In_1210);
nand U4241 (N_4241,In_679,In_2938);
xor U4242 (N_4242,In_2577,In_1262);
xor U4243 (N_4243,In_1126,In_2158);
nor U4244 (N_4244,In_2957,In_538);
xnor U4245 (N_4245,In_2871,In_421);
and U4246 (N_4246,In_1547,In_2764);
xor U4247 (N_4247,In_1376,In_2856);
or U4248 (N_4248,In_176,In_680);
xor U4249 (N_4249,In_1502,In_2922);
or U4250 (N_4250,In_1658,In_453);
nor U4251 (N_4251,In_251,In_1206);
nor U4252 (N_4252,In_1695,In_2777);
or U4253 (N_4253,In_2840,In_1635);
and U4254 (N_4254,In_1969,In_1055);
nor U4255 (N_4255,In_1152,In_1905);
or U4256 (N_4256,In_105,In_1683);
or U4257 (N_4257,In_1768,In_2944);
xnor U4258 (N_4258,In_1202,In_1699);
and U4259 (N_4259,In_1928,In_1904);
and U4260 (N_4260,In_2998,In_2942);
xor U4261 (N_4261,In_630,In_582);
nor U4262 (N_4262,In_1062,In_1534);
or U4263 (N_4263,In_1488,In_173);
and U4264 (N_4264,In_819,In_1127);
xnor U4265 (N_4265,In_31,In_1650);
or U4266 (N_4266,In_1335,In_2974);
and U4267 (N_4267,In_493,In_1669);
xnor U4268 (N_4268,In_774,In_1619);
nand U4269 (N_4269,In_2320,In_2839);
or U4270 (N_4270,In_2919,In_2169);
and U4271 (N_4271,In_2573,In_453);
and U4272 (N_4272,In_939,In_508);
nand U4273 (N_4273,In_1799,In_1379);
xnor U4274 (N_4274,In_1209,In_2156);
nand U4275 (N_4275,In_2881,In_1220);
and U4276 (N_4276,In_1167,In_1902);
nand U4277 (N_4277,In_428,In_462);
or U4278 (N_4278,In_801,In_425);
nand U4279 (N_4279,In_357,In_244);
xor U4280 (N_4280,In_2441,In_849);
and U4281 (N_4281,In_2306,In_2407);
and U4282 (N_4282,In_306,In_150);
xnor U4283 (N_4283,In_1206,In_456);
xnor U4284 (N_4284,In_2961,In_1497);
nor U4285 (N_4285,In_1858,In_2557);
or U4286 (N_4286,In_590,In_123);
and U4287 (N_4287,In_2132,In_276);
or U4288 (N_4288,In_2505,In_1103);
and U4289 (N_4289,In_1536,In_1684);
and U4290 (N_4290,In_1154,In_2591);
and U4291 (N_4291,In_1366,In_1850);
xnor U4292 (N_4292,In_443,In_1361);
and U4293 (N_4293,In_2688,In_1088);
nor U4294 (N_4294,In_441,In_1893);
nor U4295 (N_4295,In_1448,In_2703);
xor U4296 (N_4296,In_1507,In_2469);
or U4297 (N_4297,In_673,In_2763);
nand U4298 (N_4298,In_632,In_400);
or U4299 (N_4299,In_1317,In_1509);
xor U4300 (N_4300,In_1498,In_2075);
or U4301 (N_4301,In_1576,In_2393);
nor U4302 (N_4302,In_2843,In_1683);
xnor U4303 (N_4303,In_112,In_957);
xor U4304 (N_4304,In_2208,In_2054);
nor U4305 (N_4305,In_2242,In_154);
or U4306 (N_4306,In_2966,In_28);
xnor U4307 (N_4307,In_1623,In_1266);
nand U4308 (N_4308,In_879,In_269);
xor U4309 (N_4309,In_787,In_2217);
nor U4310 (N_4310,In_2912,In_2428);
nand U4311 (N_4311,In_1309,In_2672);
nand U4312 (N_4312,In_1437,In_1241);
and U4313 (N_4313,In_643,In_965);
or U4314 (N_4314,In_2326,In_219);
nand U4315 (N_4315,In_1524,In_256);
and U4316 (N_4316,In_736,In_312);
xnor U4317 (N_4317,In_2992,In_2289);
nand U4318 (N_4318,In_1270,In_980);
and U4319 (N_4319,In_1628,In_643);
xnor U4320 (N_4320,In_2399,In_932);
or U4321 (N_4321,In_920,In_2737);
and U4322 (N_4322,In_1754,In_985);
or U4323 (N_4323,In_1527,In_1390);
xor U4324 (N_4324,In_2140,In_749);
and U4325 (N_4325,In_1018,In_1370);
nand U4326 (N_4326,In_1925,In_1088);
nand U4327 (N_4327,In_1391,In_1654);
and U4328 (N_4328,In_2286,In_477);
or U4329 (N_4329,In_2330,In_1799);
nand U4330 (N_4330,In_2205,In_2913);
or U4331 (N_4331,In_1898,In_2309);
or U4332 (N_4332,In_1823,In_2925);
nor U4333 (N_4333,In_2532,In_2860);
xor U4334 (N_4334,In_1676,In_1373);
xnor U4335 (N_4335,In_741,In_989);
nor U4336 (N_4336,In_1607,In_2915);
and U4337 (N_4337,In_675,In_385);
nor U4338 (N_4338,In_1825,In_2863);
nand U4339 (N_4339,In_933,In_2747);
xor U4340 (N_4340,In_2833,In_2254);
nand U4341 (N_4341,In_298,In_989);
or U4342 (N_4342,In_1231,In_671);
xnor U4343 (N_4343,In_1531,In_2722);
nor U4344 (N_4344,In_1439,In_1351);
xor U4345 (N_4345,In_159,In_2120);
and U4346 (N_4346,In_506,In_141);
and U4347 (N_4347,In_2184,In_1482);
nand U4348 (N_4348,In_1204,In_1515);
nand U4349 (N_4349,In_2336,In_988);
and U4350 (N_4350,In_190,In_2106);
xor U4351 (N_4351,In_1438,In_1699);
xor U4352 (N_4352,In_1742,In_183);
and U4353 (N_4353,In_280,In_2405);
nor U4354 (N_4354,In_1622,In_565);
xor U4355 (N_4355,In_2298,In_2835);
xor U4356 (N_4356,In_1904,In_2006);
xnor U4357 (N_4357,In_1505,In_2870);
and U4358 (N_4358,In_944,In_439);
xnor U4359 (N_4359,In_1996,In_2748);
nor U4360 (N_4360,In_1672,In_364);
nor U4361 (N_4361,In_1585,In_982);
and U4362 (N_4362,In_2931,In_2248);
and U4363 (N_4363,In_1553,In_1586);
nor U4364 (N_4364,In_2639,In_1641);
nor U4365 (N_4365,In_2734,In_1174);
or U4366 (N_4366,In_262,In_2475);
nor U4367 (N_4367,In_2970,In_645);
or U4368 (N_4368,In_546,In_2643);
and U4369 (N_4369,In_642,In_1072);
or U4370 (N_4370,In_940,In_2912);
nor U4371 (N_4371,In_1283,In_939);
or U4372 (N_4372,In_1942,In_291);
nor U4373 (N_4373,In_745,In_2235);
xnor U4374 (N_4374,In_2737,In_1952);
nor U4375 (N_4375,In_2207,In_2041);
nor U4376 (N_4376,In_2725,In_103);
or U4377 (N_4377,In_2595,In_728);
and U4378 (N_4378,In_2322,In_77);
nand U4379 (N_4379,In_1592,In_2432);
and U4380 (N_4380,In_280,In_27);
and U4381 (N_4381,In_1616,In_1451);
and U4382 (N_4382,In_2482,In_2224);
nor U4383 (N_4383,In_2975,In_2520);
nor U4384 (N_4384,In_983,In_812);
nand U4385 (N_4385,In_2756,In_888);
or U4386 (N_4386,In_2320,In_871);
nand U4387 (N_4387,In_2198,In_1703);
xor U4388 (N_4388,In_662,In_2161);
and U4389 (N_4389,In_1990,In_541);
nand U4390 (N_4390,In_607,In_2319);
or U4391 (N_4391,In_2530,In_1638);
or U4392 (N_4392,In_2431,In_395);
and U4393 (N_4393,In_805,In_113);
or U4394 (N_4394,In_335,In_706);
or U4395 (N_4395,In_19,In_149);
and U4396 (N_4396,In_1545,In_343);
nor U4397 (N_4397,In_2834,In_2409);
xor U4398 (N_4398,In_1875,In_1647);
or U4399 (N_4399,In_13,In_1347);
or U4400 (N_4400,In_1276,In_93);
and U4401 (N_4401,In_1063,In_817);
and U4402 (N_4402,In_468,In_1842);
or U4403 (N_4403,In_422,In_2575);
xor U4404 (N_4404,In_1339,In_1465);
nand U4405 (N_4405,In_2663,In_2761);
and U4406 (N_4406,In_332,In_992);
and U4407 (N_4407,In_2082,In_2270);
or U4408 (N_4408,In_287,In_578);
xor U4409 (N_4409,In_1547,In_2890);
and U4410 (N_4410,In_2170,In_1366);
nor U4411 (N_4411,In_931,In_898);
nor U4412 (N_4412,In_1053,In_250);
and U4413 (N_4413,In_536,In_938);
and U4414 (N_4414,In_2378,In_1425);
nand U4415 (N_4415,In_1139,In_2034);
nor U4416 (N_4416,In_216,In_2824);
or U4417 (N_4417,In_396,In_673);
or U4418 (N_4418,In_2435,In_2751);
nor U4419 (N_4419,In_4,In_2733);
or U4420 (N_4420,In_676,In_991);
xor U4421 (N_4421,In_2372,In_1197);
nand U4422 (N_4422,In_2397,In_2232);
and U4423 (N_4423,In_16,In_2468);
xor U4424 (N_4424,In_1008,In_1949);
or U4425 (N_4425,In_2524,In_819);
and U4426 (N_4426,In_1429,In_1161);
nor U4427 (N_4427,In_2374,In_1223);
nor U4428 (N_4428,In_2419,In_1964);
nor U4429 (N_4429,In_998,In_1006);
xor U4430 (N_4430,In_2695,In_2229);
nand U4431 (N_4431,In_447,In_2607);
nor U4432 (N_4432,In_1292,In_2145);
and U4433 (N_4433,In_842,In_2417);
and U4434 (N_4434,In_2490,In_1590);
or U4435 (N_4435,In_2896,In_2326);
xor U4436 (N_4436,In_1659,In_652);
nand U4437 (N_4437,In_779,In_616);
nand U4438 (N_4438,In_890,In_1101);
and U4439 (N_4439,In_1566,In_569);
nor U4440 (N_4440,In_2265,In_2862);
or U4441 (N_4441,In_739,In_2582);
xnor U4442 (N_4442,In_453,In_369);
nand U4443 (N_4443,In_1892,In_1699);
nor U4444 (N_4444,In_1842,In_1665);
and U4445 (N_4445,In_1894,In_1141);
nand U4446 (N_4446,In_2972,In_2679);
or U4447 (N_4447,In_686,In_1005);
nor U4448 (N_4448,In_114,In_1231);
nand U4449 (N_4449,In_2109,In_2225);
nor U4450 (N_4450,In_2191,In_27);
xor U4451 (N_4451,In_2151,In_1100);
or U4452 (N_4452,In_1011,In_2103);
nor U4453 (N_4453,In_2960,In_1586);
or U4454 (N_4454,In_831,In_2557);
nor U4455 (N_4455,In_1726,In_649);
nor U4456 (N_4456,In_72,In_582);
or U4457 (N_4457,In_2033,In_168);
and U4458 (N_4458,In_446,In_1632);
and U4459 (N_4459,In_913,In_1753);
xnor U4460 (N_4460,In_2742,In_1542);
nand U4461 (N_4461,In_2879,In_1339);
and U4462 (N_4462,In_1609,In_2730);
xor U4463 (N_4463,In_41,In_123);
xor U4464 (N_4464,In_1410,In_2223);
xnor U4465 (N_4465,In_888,In_1831);
or U4466 (N_4466,In_268,In_1216);
nor U4467 (N_4467,In_1568,In_2929);
nand U4468 (N_4468,In_2924,In_270);
nor U4469 (N_4469,In_982,In_2319);
nand U4470 (N_4470,In_870,In_1415);
nor U4471 (N_4471,In_649,In_2643);
and U4472 (N_4472,In_1501,In_2830);
xnor U4473 (N_4473,In_997,In_710);
nand U4474 (N_4474,In_100,In_756);
xor U4475 (N_4475,In_833,In_652);
and U4476 (N_4476,In_191,In_2155);
nor U4477 (N_4477,In_2548,In_644);
and U4478 (N_4478,In_2277,In_778);
or U4479 (N_4479,In_1048,In_1745);
xnor U4480 (N_4480,In_576,In_1933);
xnor U4481 (N_4481,In_1531,In_2332);
xor U4482 (N_4482,In_1093,In_2421);
and U4483 (N_4483,In_2851,In_449);
xnor U4484 (N_4484,In_594,In_2743);
nand U4485 (N_4485,In_2194,In_1085);
and U4486 (N_4486,In_1712,In_1840);
nand U4487 (N_4487,In_1046,In_1969);
and U4488 (N_4488,In_362,In_2487);
and U4489 (N_4489,In_1544,In_1754);
nor U4490 (N_4490,In_1351,In_2610);
or U4491 (N_4491,In_1245,In_2610);
nand U4492 (N_4492,In_584,In_1678);
and U4493 (N_4493,In_617,In_2434);
or U4494 (N_4494,In_2905,In_908);
or U4495 (N_4495,In_1899,In_1464);
nand U4496 (N_4496,In_1583,In_235);
nor U4497 (N_4497,In_2636,In_1811);
xnor U4498 (N_4498,In_2083,In_1509);
nand U4499 (N_4499,In_370,In_621);
or U4500 (N_4500,In_2666,In_739);
xor U4501 (N_4501,In_755,In_2412);
or U4502 (N_4502,In_1799,In_1125);
nor U4503 (N_4503,In_1370,In_2907);
or U4504 (N_4504,In_593,In_874);
nand U4505 (N_4505,In_2661,In_193);
and U4506 (N_4506,In_792,In_2757);
or U4507 (N_4507,In_2560,In_2381);
nand U4508 (N_4508,In_2429,In_493);
nand U4509 (N_4509,In_1849,In_2549);
xor U4510 (N_4510,In_2084,In_1849);
or U4511 (N_4511,In_190,In_2566);
nor U4512 (N_4512,In_1484,In_167);
xor U4513 (N_4513,In_699,In_445);
and U4514 (N_4514,In_2951,In_1799);
nor U4515 (N_4515,In_2577,In_191);
nor U4516 (N_4516,In_1541,In_2800);
nor U4517 (N_4517,In_1325,In_736);
nand U4518 (N_4518,In_810,In_579);
or U4519 (N_4519,In_646,In_383);
or U4520 (N_4520,In_2063,In_2297);
and U4521 (N_4521,In_2308,In_1678);
nand U4522 (N_4522,In_2692,In_1470);
and U4523 (N_4523,In_668,In_1135);
or U4524 (N_4524,In_129,In_231);
xnor U4525 (N_4525,In_1942,In_2291);
or U4526 (N_4526,In_537,In_2527);
and U4527 (N_4527,In_2338,In_974);
and U4528 (N_4528,In_2677,In_1259);
or U4529 (N_4529,In_701,In_741);
or U4530 (N_4530,In_276,In_1825);
nand U4531 (N_4531,In_1363,In_2246);
nand U4532 (N_4532,In_311,In_1569);
nand U4533 (N_4533,In_2824,In_2879);
xnor U4534 (N_4534,In_982,In_590);
nand U4535 (N_4535,In_2345,In_591);
xor U4536 (N_4536,In_1075,In_167);
and U4537 (N_4537,In_1630,In_999);
nor U4538 (N_4538,In_2896,In_2804);
and U4539 (N_4539,In_582,In_1392);
nor U4540 (N_4540,In_2255,In_715);
nand U4541 (N_4541,In_1017,In_781);
xor U4542 (N_4542,In_68,In_2232);
or U4543 (N_4543,In_1648,In_1769);
and U4544 (N_4544,In_566,In_96);
nor U4545 (N_4545,In_1915,In_155);
nor U4546 (N_4546,In_2581,In_1880);
nor U4547 (N_4547,In_791,In_2669);
xor U4548 (N_4548,In_1240,In_806);
xnor U4549 (N_4549,In_716,In_148);
nand U4550 (N_4550,In_1326,In_1491);
nand U4551 (N_4551,In_1392,In_2064);
and U4552 (N_4552,In_2811,In_1204);
xor U4553 (N_4553,In_1957,In_2732);
xor U4554 (N_4554,In_2770,In_270);
or U4555 (N_4555,In_2675,In_2596);
nor U4556 (N_4556,In_470,In_165);
nand U4557 (N_4557,In_2252,In_369);
nand U4558 (N_4558,In_2379,In_65);
nand U4559 (N_4559,In_941,In_1743);
nand U4560 (N_4560,In_2724,In_814);
or U4561 (N_4561,In_925,In_2822);
and U4562 (N_4562,In_1973,In_2943);
nor U4563 (N_4563,In_2496,In_2338);
xor U4564 (N_4564,In_1179,In_426);
or U4565 (N_4565,In_786,In_2181);
or U4566 (N_4566,In_1818,In_1406);
and U4567 (N_4567,In_1898,In_2574);
nand U4568 (N_4568,In_141,In_442);
nand U4569 (N_4569,In_2206,In_1276);
nand U4570 (N_4570,In_785,In_2235);
nor U4571 (N_4571,In_402,In_1621);
and U4572 (N_4572,In_2291,In_1258);
or U4573 (N_4573,In_630,In_888);
or U4574 (N_4574,In_2762,In_1258);
nand U4575 (N_4575,In_1208,In_131);
nor U4576 (N_4576,In_2345,In_2522);
or U4577 (N_4577,In_1046,In_776);
and U4578 (N_4578,In_792,In_2344);
or U4579 (N_4579,In_2020,In_1543);
nand U4580 (N_4580,In_1496,In_1969);
xnor U4581 (N_4581,In_1471,In_2554);
and U4582 (N_4582,In_683,In_1992);
nand U4583 (N_4583,In_1715,In_484);
and U4584 (N_4584,In_2168,In_2170);
nand U4585 (N_4585,In_1272,In_1781);
nor U4586 (N_4586,In_542,In_1648);
xor U4587 (N_4587,In_2582,In_1738);
nand U4588 (N_4588,In_951,In_2250);
xnor U4589 (N_4589,In_33,In_756);
xor U4590 (N_4590,In_1596,In_2084);
nand U4591 (N_4591,In_1883,In_2596);
xnor U4592 (N_4592,In_2596,In_172);
nor U4593 (N_4593,In_1705,In_432);
or U4594 (N_4594,In_1287,In_181);
and U4595 (N_4595,In_2389,In_2465);
xnor U4596 (N_4596,In_571,In_2271);
or U4597 (N_4597,In_57,In_2595);
nand U4598 (N_4598,In_848,In_740);
xor U4599 (N_4599,In_1047,In_2451);
or U4600 (N_4600,In_422,In_822);
and U4601 (N_4601,In_993,In_1093);
nand U4602 (N_4602,In_1531,In_480);
and U4603 (N_4603,In_1656,In_146);
nor U4604 (N_4604,In_1551,In_408);
nand U4605 (N_4605,In_2111,In_72);
nor U4606 (N_4606,In_2630,In_1297);
and U4607 (N_4607,In_1769,In_2686);
or U4608 (N_4608,In_1338,In_884);
xnor U4609 (N_4609,In_261,In_446);
and U4610 (N_4610,In_2785,In_991);
xnor U4611 (N_4611,In_171,In_18);
xnor U4612 (N_4612,In_1149,In_2016);
nor U4613 (N_4613,In_1925,In_2741);
or U4614 (N_4614,In_1296,In_1351);
nand U4615 (N_4615,In_922,In_742);
xor U4616 (N_4616,In_986,In_2821);
nand U4617 (N_4617,In_2455,In_592);
xnor U4618 (N_4618,In_666,In_683);
xor U4619 (N_4619,In_461,In_434);
or U4620 (N_4620,In_130,In_2155);
nor U4621 (N_4621,In_391,In_2291);
nor U4622 (N_4622,In_933,In_633);
xnor U4623 (N_4623,In_461,In_2821);
nand U4624 (N_4624,In_1321,In_2727);
nor U4625 (N_4625,In_2122,In_283);
nand U4626 (N_4626,In_324,In_566);
nand U4627 (N_4627,In_2043,In_789);
nand U4628 (N_4628,In_118,In_464);
or U4629 (N_4629,In_2286,In_838);
nand U4630 (N_4630,In_2812,In_1401);
and U4631 (N_4631,In_345,In_656);
nor U4632 (N_4632,In_553,In_2246);
xor U4633 (N_4633,In_1504,In_882);
or U4634 (N_4634,In_747,In_294);
and U4635 (N_4635,In_2075,In_1675);
or U4636 (N_4636,In_1229,In_601);
xnor U4637 (N_4637,In_1625,In_2343);
xor U4638 (N_4638,In_2210,In_303);
or U4639 (N_4639,In_1409,In_143);
or U4640 (N_4640,In_981,In_2307);
nor U4641 (N_4641,In_134,In_118);
or U4642 (N_4642,In_1762,In_2150);
nor U4643 (N_4643,In_2668,In_187);
xor U4644 (N_4644,In_1309,In_604);
xor U4645 (N_4645,In_1869,In_337);
and U4646 (N_4646,In_1062,In_168);
and U4647 (N_4647,In_719,In_1891);
nor U4648 (N_4648,In_1179,In_2249);
xor U4649 (N_4649,In_221,In_2874);
and U4650 (N_4650,In_1864,In_842);
nor U4651 (N_4651,In_2970,In_1642);
and U4652 (N_4652,In_500,In_2705);
and U4653 (N_4653,In_1635,In_2131);
nor U4654 (N_4654,In_2356,In_2177);
nor U4655 (N_4655,In_133,In_1490);
xnor U4656 (N_4656,In_997,In_1975);
nor U4657 (N_4657,In_1430,In_1285);
and U4658 (N_4658,In_2673,In_2812);
and U4659 (N_4659,In_2013,In_1483);
or U4660 (N_4660,In_571,In_329);
xor U4661 (N_4661,In_278,In_2230);
nand U4662 (N_4662,In_2681,In_2486);
and U4663 (N_4663,In_188,In_2533);
and U4664 (N_4664,In_343,In_1680);
or U4665 (N_4665,In_289,In_927);
or U4666 (N_4666,In_481,In_2817);
or U4667 (N_4667,In_2436,In_960);
or U4668 (N_4668,In_1544,In_17);
nor U4669 (N_4669,In_1998,In_1667);
nand U4670 (N_4670,In_1848,In_1977);
nand U4671 (N_4671,In_2185,In_981);
xnor U4672 (N_4672,In_542,In_505);
xor U4673 (N_4673,In_2711,In_1008);
or U4674 (N_4674,In_169,In_1516);
xnor U4675 (N_4675,In_2805,In_20);
xnor U4676 (N_4676,In_463,In_346);
nand U4677 (N_4677,In_2873,In_1629);
or U4678 (N_4678,In_1659,In_1534);
or U4679 (N_4679,In_981,In_467);
or U4680 (N_4680,In_1972,In_1479);
and U4681 (N_4681,In_1297,In_1544);
nor U4682 (N_4682,In_2786,In_103);
and U4683 (N_4683,In_982,In_2542);
or U4684 (N_4684,In_206,In_249);
nand U4685 (N_4685,In_2148,In_239);
and U4686 (N_4686,In_677,In_2216);
and U4687 (N_4687,In_2192,In_775);
or U4688 (N_4688,In_1826,In_2754);
nand U4689 (N_4689,In_1003,In_1551);
nand U4690 (N_4690,In_2788,In_2457);
nand U4691 (N_4691,In_2506,In_1651);
nand U4692 (N_4692,In_960,In_686);
or U4693 (N_4693,In_819,In_2003);
nor U4694 (N_4694,In_756,In_1032);
nor U4695 (N_4695,In_1124,In_2742);
nand U4696 (N_4696,In_318,In_1617);
nand U4697 (N_4697,In_2521,In_2800);
and U4698 (N_4698,In_59,In_1172);
xnor U4699 (N_4699,In_820,In_571);
nor U4700 (N_4700,In_624,In_2129);
nand U4701 (N_4701,In_949,In_1671);
nor U4702 (N_4702,In_2750,In_1748);
nand U4703 (N_4703,In_2582,In_153);
nand U4704 (N_4704,In_1965,In_784);
nor U4705 (N_4705,In_1945,In_73);
and U4706 (N_4706,In_2235,In_196);
or U4707 (N_4707,In_1053,In_2637);
and U4708 (N_4708,In_1805,In_1727);
nand U4709 (N_4709,In_2262,In_2999);
nor U4710 (N_4710,In_1113,In_1819);
and U4711 (N_4711,In_999,In_2533);
or U4712 (N_4712,In_2144,In_2063);
xor U4713 (N_4713,In_2049,In_144);
nand U4714 (N_4714,In_46,In_1019);
nand U4715 (N_4715,In_486,In_510);
xor U4716 (N_4716,In_989,In_1535);
and U4717 (N_4717,In_456,In_1240);
xor U4718 (N_4718,In_2122,In_2330);
or U4719 (N_4719,In_2699,In_2799);
and U4720 (N_4720,In_1037,In_2232);
nand U4721 (N_4721,In_680,In_1546);
xnor U4722 (N_4722,In_2290,In_1765);
nor U4723 (N_4723,In_2405,In_1376);
nand U4724 (N_4724,In_2527,In_1889);
nand U4725 (N_4725,In_2607,In_297);
nor U4726 (N_4726,In_39,In_818);
and U4727 (N_4727,In_159,In_2089);
and U4728 (N_4728,In_2172,In_561);
nor U4729 (N_4729,In_657,In_2122);
and U4730 (N_4730,In_1396,In_1564);
or U4731 (N_4731,In_844,In_2266);
nand U4732 (N_4732,In_19,In_2578);
xor U4733 (N_4733,In_2124,In_195);
nor U4734 (N_4734,In_2894,In_2662);
or U4735 (N_4735,In_2667,In_126);
or U4736 (N_4736,In_916,In_2081);
and U4737 (N_4737,In_531,In_1856);
and U4738 (N_4738,In_796,In_1036);
nor U4739 (N_4739,In_1260,In_1005);
xor U4740 (N_4740,In_1845,In_2198);
nand U4741 (N_4741,In_1366,In_2798);
xor U4742 (N_4742,In_1467,In_560);
xnor U4743 (N_4743,In_2788,In_2442);
nor U4744 (N_4744,In_1510,In_1931);
and U4745 (N_4745,In_1472,In_604);
nand U4746 (N_4746,In_1752,In_2547);
and U4747 (N_4747,In_814,In_1540);
nand U4748 (N_4748,In_877,In_2918);
xor U4749 (N_4749,In_2950,In_565);
nand U4750 (N_4750,In_1751,In_2249);
or U4751 (N_4751,In_1051,In_711);
or U4752 (N_4752,In_2853,In_984);
nor U4753 (N_4753,In_2958,In_648);
and U4754 (N_4754,In_1326,In_1599);
and U4755 (N_4755,In_1467,In_1636);
xnor U4756 (N_4756,In_1239,In_2187);
nand U4757 (N_4757,In_2574,In_1258);
or U4758 (N_4758,In_2500,In_2302);
and U4759 (N_4759,In_545,In_1962);
nor U4760 (N_4760,In_775,In_1948);
nor U4761 (N_4761,In_2890,In_2200);
xnor U4762 (N_4762,In_2377,In_619);
nand U4763 (N_4763,In_1507,In_2269);
nand U4764 (N_4764,In_439,In_2141);
nor U4765 (N_4765,In_2049,In_2647);
nand U4766 (N_4766,In_1133,In_1303);
or U4767 (N_4767,In_549,In_956);
or U4768 (N_4768,In_106,In_1919);
nor U4769 (N_4769,In_1117,In_2469);
and U4770 (N_4770,In_970,In_886);
xor U4771 (N_4771,In_2180,In_320);
nor U4772 (N_4772,In_586,In_317);
nor U4773 (N_4773,In_2388,In_1010);
nand U4774 (N_4774,In_2566,In_641);
nand U4775 (N_4775,In_2515,In_2834);
and U4776 (N_4776,In_2686,In_1795);
xor U4777 (N_4777,In_2311,In_760);
nor U4778 (N_4778,In_2913,In_1474);
nand U4779 (N_4779,In_912,In_280);
nand U4780 (N_4780,In_1934,In_1773);
or U4781 (N_4781,In_2316,In_1599);
nand U4782 (N_4782,In_2124,In_1244);
xor U4783 (N_4783,In_2377,In_2822);
xor U4784 (N_4784,In_1104,In_1500);
and U4785 (N_4785,In_2897,In_1721);
and U4786 (N_4786,In_1772,In_235);
xnor U4787 (N_4787,In_2984,In_2697);
nor U4788 (N_4788,In_2422,In_2454);
or U4789 (N_4789,In_684,In_1373);
xnor U4790 (N_4790,In_1357,In_2365);
and U4791 (N_4791,In_662,In_938);
or U4792 (N_4792,In_273,In_1302);
or U4793 (N_4793,In_714,In_800);
nand U4794 (N_4794,In_1329,In_242);
or U4795 (N_4795,In_406,In_22);
and U4796 (N_4796,In_430,In_180);
or U4797 (N_4797,In_211,In_1147);
or U4798 (N_4798,In_655,In_504);
nor U4799 (N_4799,In_1059,In_1775);
or U4800 (N_4800,In_1973,In_2120);
and U4801 (N_4801,In_2398,In_10);
nor U4802 (N_4802,In_2270,In_2244);
or U4803 (N_4803,In_1697,In_1118);
and U4804 (N_4804,In_1685,In_2972);
or U4805 (N_4805,In_1077,In_1791);
or U4806 (N_4806,In_1492,In_2997);
or U4807 (N_4807,In_2544,In_1305);
or U4808 (N_4808,In_2450,In_2928);
nor U4809 (N_4809,In_398,In_2002);
or U4810 (N_4810,In_2777,In_1496);
nor U4811 (N_4811,In_2649,In_1035);
nand U4812 (N_4812,In_1256,In_449);
nand U4813 (N_4813,In_1571,In_1130);
or U4814 (N_4814,In_1359,In_237);
nor U4815 (N_4815,In_2708,In_2112);
nor U4816 (N_4816,In_1189,In_2843);
xnor U4817 (N_4817,In_1024,In_2656);
xnor U4818 (N_4818,In_1060,In_2249);
xor U4819 (N_4819,In_782,In_1157);
or U4820 (N_4820,In_696,In_975);
xor U4821 (N_4821,In_674,In_1053);
xnor U4822 (N_4822,In_811,In_2267);
or U4823 (N_4823,In_115,In_13);
xnor U4824 (N_4824,In_2636,In_386);
and U4825 (N_4825,In_287,In_665);
nand U4826 (N_4826,In_2950,In_1816);
and U4827 (N_4827,In_2481,In_1090);
and U4828 (N_4828,In_2833,In_1382);
nor U4829 (N_4829,In_84,In_1243);
nor U4830 (N_4830,In_2746,In_1576);
or U4831 (N_4831,In_2165,In_1595);
xnor U4832 (N_4832,In_1016,In_1714);
and U4833 (N_4833,In_2891,In_1823);
or U4834 (N_4834,In_140,In_2594);
nand U4835 (N_4835,In_52,In_1965);
and U4836 (N_4836,In_2373,In_1194);
nor U4837 (N_4837,In_1631,In_1142);
or U4838 (N_4838,In_1938,In_377);
nand U4839 (N_4839,In_2954,In_1400);
nand U4840 (N_4840,In_2341,In_357);
xnor U4841 (N_4841,In_1169,In_1350);
or U4842 (N_4842,In_2081,In_2992);
or U4843 (N_4843,In_1482,In_1579);
nand U4844 (N_4844,In_800,In_2849);
xor U4845 (N_4845,In_1661,In_1881);
nor U4846 (N_4846,In_673,In_2167);
xor U4847 (N_4847,In_1788,In_589);
xnor U4848 (N_4848,In_48,In_1110);
and U4849 (N_4849,In_1404,In_1368);
xor U4850 (N_4850,In_1124,In_830);
or U4851 (N_4851,In_704,In_2560);
or U4852 (N_4852,In_2651,In_231);
nand U4853 (N_4853,In_2203,In_248);
or U4854 (N_4854,In_585,In_849);
nor U4855 (N_4855,In_1441,In_564);
or U4856 (N_4856,In_1634,In_2803);
nand U4857 (N_4857,In_1883,In_471);
xor U4858 (N_4858,In_2625,In_2292);
nand U4859 (N_4859,In_1786,In_2052);
or U4860 (N_4860,In_1906,In_1290);
xnor U4861 (N_4861,In_2977,In_2165);
nor U4862 (N_4862,In_2536,In_2362);
nand U4863 (N_4863,In_836,In_58);
nor U4864 (N_4864,In_2903,In_49);
or U4865 (N_4865,In_2197,In_1670);
xnor U4866 (N_4866,In_2214,In_2581);
xor U4867 (N_4867,In_325,In_1166);
and U4868 (N_4868,In_450,In_255);
nand U4869 (N_4869,In_2009,In_2955);
xnor U4870 (N_4870,In_1198,In_15);
nor U4871 (N_4871,In_2962,In_2681);
nand U4872 (N_4872,In_2672,In_1307);
and U4873 (N_4873,In_2616,In_803);
or U4874 (N_4874,In_1838,In_581);
or U4875 (N_4875,In_968,In_2873);
or U4876 (N_4876,In_1537,In_2563);
and U4877 (N_4877,In_2184,In_2510);
or U4878 (N_4878,In_1246,In_2185);
nand U4879 (N_4879,In_2843,In_818);
xnor U4880 (N_4880,In_1766,In_400);
and U4881 (N_4881,In_2914,In_281);
nor U4882 (N_4882,In_2733,In_1883);
nand U4883 (N_4883,In_721,In_613);
nor U4884 (N_4884,In_2774,In_1565);
nor U4885 (N_4885,In_395,In_2299);
and U4886 (N_4886,In_1507,In_51);
xnor U4887 (N_4887,In_2588,In_333);
or U4888 (N_4888,In_2038,In_1606);
xnor U4889 (N_4889,In_1658,In_231);
xor U4890 (N_4890,In_2733,In_2296);
nor U4891 (N_4891,In_1078,In_552);
or U4892 (N_4892,In_414,In_201);
xor U4893 (N_4893,In_261,In_2799);
nand U4894 (N_4894,In_769,In_1871);
nor U4895 (N_4895,In_1902,In_1400);
nor U4896 (N_4896,In_1162,In_2284);
nor U4897 (N_4897,In_1975,In_652);
or U4898 (N_4898,In_1485,In_400);
and U4899 (N_4899,In_2610,In_1347);
xor U4900 (N_4900,In_173,In_904);
nor U4901 (N_4901,In_459,In_1574);
nand U4902 (N_4902,In_2223,In_1200);
and U4903 (N_4903,In_2804,In_2705);
nor U4904 (N_4904,In_596,In_2179);
xor U4905 (N_4905,In_1790,In_31);
or U4906 (N_4906,In_1313,In_1608);
or U4907 (N_4907,In_2684,In_2161);
nor U4908 (N_4908,In_1924,In_1446);
or U4909 (N_4909,In_2323,In_1430);
and U4910 (N_4910,In_841,In_2544);
nand U4911 (N_4911,In_1860,In_955);
or U4912 (N_4912,In_2550,In_1627);
nor U4913 (N_4913,In_600,In_1199);
nor U4914 (N_4914,In_2437,In_2466);
or U4915 (N_4915,In_1392,In_2747);
xnor U4916 (N_4916,In_2237,In_1146);
and U4917 (N_4917,In_2437,In_763);
nand U4918 (N_4918,In_678,In_726);
xor U4919 (N_4919,In_2456,In_1409);
xor U4920 (N_4920,In_2499,In_1416);
nand U4921 (N_4921,In_2052,In_2692);
xnor U4922 (N_4922,In_156,In_2638);
and U4923 (N_4923,In_1232,In_2442);
nand U4924 (N_4924,In_2086,In_2364);
nand U4925 (N_4925,In_2830,In_633);
or U4926 (N_4926,In_1988,In_2044);
xor U4927 (N_4927,In_2605,In_727);
nand U4928 (N_4928,In_1040,In_1195);
nand U4929 (N_4929,In_2479,In_910);
or U4930 (N_4930,In_1237,In_1034);
xnor U4931 (N_4931,In_292,In_1490);
nor U4932 (N_4932,In_2143,In_344);
xnor U4933 (N_4933,In_910,In_358);
or U4934 (N_4934,In_2701,In_546);
xnor U4935 (N_4935,In_2828,In_2055);
or U4936 (N_4936,In_2475,In_1257);
or U4937 (N_4937,In_2322,In_1026);
xnor U4938 (N_4938,In_1336,In_1185);
nor U4939 (N_4939,In_1303,In_332);
nand U4940 (N_4940,In_2912,In_1158);
xnor U4941 (N_4941,In_3,In_953);
nor U4942 (N_4942,In_177,In_2109);
nand U4943 (N_4943,In_643,In_73);
and U4944 (N_4944,In_2968,In_1619);
and U4945 (N_4945,In_1931,In_749);
xor U4946 (N_4946,In_782,In_651);
nor U4947 (N_4947,In_2801,In_2606);
nor U4948 (N_4948,In_105,In_464);
or U4949 (N_4949,In_2175,In_680);
nand U4950 (N_4950,In_2215,In_349);
xnor U4951 (N_4951,In_2341,In_1590);
or U4952 (N_4952,In_127,In_837);
nand U4953 (N_4953,In_714,In_1447);
and U4954 (N_4954,In_1329,In_2673);
xor U4955 (N_4955,In_1643,In_1906);
and U4956 (N_4956,In_2931,In_1610);
or U4957 (N_4957,In_1233,In_1559);
xnor U4958 (N_4958,In_2506,In_1284);
nor U4959 (N_4959,In_715,In_2037);
xor U4960 (N_4960,In_97,In_557);
and U4961 (N_4961,In_1499,In_548);
nor U4962 (N_4962,In_531,In_656);
or U4963 (N_4963,In_1699,In_1420);
or U4964 (N_4964,In_2337,In_1580);
nor U4965 (N_4965,In_1014,In_861);
nand U4966 (N_4966,In_519,In_1510);
or U4967 (N_4967,In_1233,In_2941);
nand U4968 (N_4968,In_1845,In_1475);
and U4969 (N_4969,In_1069,In_2772);
nand U4970 (N_4970,In_1930,In_1663);
and U4971 (N_4971,In_2585,In_1224);
nor U4972 (N_4972,In_726,In_365);
or U4973 (N_4973,In_1279,In_2249);
xnor U4974 (N_4974,In_591,In_2629);
or U4975 (N_4975,In_2468,In_2697);
nand U4976 (N_4976,In_2455,In_2534);
or U4977 (N_4977,In_2530,In_1235);
or U4978 (N_4978,In_2101,In_1687);
and U4979 (N_4979,In_738,In_2381);
nand U4980 (N_4980,In_2691,In_330);
or U4981 (N_4981,In_1240,In_825);
nor U4982 (N_4982,In_515,In_74);
or U4983 (N_4983,In_1272,In_159);
and U4984 (N_4984,In_2591,In_805);
or U4985 (N_4985,In_44,In_2811);
and U4986 (N_4986,In_89,In_1462);
or U4987 (N_4987,In_1262,In_787);
and U4988 (N_4988,In_594,In_1343);
nand U4989 (N_4989,In_42,In_440);
or U4990 (N_4990,In_1861,In_38);
xnor U4991 (N_4991,In_50,In_2508);
xor U4992 (N_4992,In_1751,In_2209);
or U4993 (N_4993,In_1584,In_2263);
and U4994 (N_4994,In_1219,In_1850);
and U4995 (N_4995,In_681,In_1523);
nand U4996 (N_4996,In_201,In_1890);
nor U4997 (N_4997,In_801,In_2447);
and U4998 (N_4998,In_2552,In_201);
or U4999 (N_4999,In_1301,In_381);
or U5000 (N_5000,N_716,N_1512);
xor U5001 (N_5001,N_3401,N_37);
nor U5002 (N_5002,N_2411,N_3329);
and U5003 (N_5003,N_20,N_2601);
and U5004 (N_5004,N_83,N_460);
or U5005 (N_5005,N_3480,N_3288);
xnor U5006 (N_5006,N_53,N_1931);
nor U5007 (N_5007,N_1952,N_4616);
nor U5008 (N_5008,N_682,N_2707);
xnor U5009 (N_5009,N_2805,N_1711);
or U5010 (N_5010,N_2547,N_3506);
xor U5011 (N_5011,N_3019,N_1483);
xor U5012 (N_5012,N_4902,N_362);
and U5013 (N_5013,N_3039,N_527);
and U5014 (N_5014,N_3676,N_1649);
nor U5015 (N_5015,N_4236,N_2982);
or U5016 (N_5016,N_1358,N_1607);
xnor U5017 (N_5017,N_3146,N_2834);
or U5018 (N_5018,N_2676,N_1984);
nor U5019 (N_5019,N_3699,N_3698);
nor U5020 (N_5020,N_2893,N_3445);
xor U5021 (N_5021,N_652,N_4939);
xnor U5022 (N_5022,N_244,N_3788);
or U5023 (N_5023,N_912,N_4361);
or U5024 (N_5024,N_3047,N_4183);
nor U5025 (N_5025,N_4261,N_1489);
nand U5026 (N_5026,N_1290,N_141);
nand U5027 (N_5027,N_3556,N_1862);
xnor U5028 (N_5028,N_591,N_2145);
or U5029 (N_5029,N_11,N_1153);
or U5030 (N_5030,N_2136,N_2196);
nor U5031 (N_5031,N_96,N_2387);
xor U5032 (N_5032,N_1331,N_3978);
xor U5033 (N_5033,N_3755,N_1226);
nor U5034 (N_5034,N_3490,N_304);
or U5035 (N_5035,N_4719,N_2261);
xnor U5036 (N_5036,N_928,N_351);
and U5037 (N_5037,N_4079,N_1492);
nor U5038 (N_5038,N_1547,N_4135);
or U5039 (N_5039,N_1637,N_4366);
or U5040 (N_5040,N_1556,N_2554);
xor U5041 (N_5041,N_4857,N_243);
nand U5042 (N_5042,N_2067,N_369);
or U5043 (N_5043,N_3128,N_338);
nand U5044 (N_5044,N_1840,N_182);
or U5045 (N_5045,N_3374,N_3562);
nand U5046 (N_5046,N_105,N_2356);
or U5047 (N_5047,N_117,N_486);
and U5048 (N_5048,N_300,N_1966);
nand U5049 (N_5049,N_1872,N_3271);
nand U5050 (N_5050,N_885,N_4766);
nor U5051 (N_5051,N_2665,N_505);
nor U5052 (N_5052,N_4259,N_4075);
nor U5053 (N_5053,N_29,N_1465);
nor U5054 (N_5054,N_3859,N_2321);
and U5055 (N_5055,N_1687,N_4073);
nor U5056 (N_5056,N_2303,N_4955);
nor U5057 (N_5057,N_26,N_3874);
nor U5058 (N_5058,N_70,N_3162);
xnor U5059 (N_5059,N_2590,N_2209);
nor U5060 (N_5060,N_4953,N_3649);
and U5061 (N_5061,N_3763,N_3514);
or U5062 (N_5062,N_2853,N_2637);
and U5063 (N_5063,N_2456,N_623);
nand U5064 (N_5064,N_2365,N_2406);
nand U5065 (N_5065,N_1460,N_1113);
xor U5066 (N_5066,N_2482,N_1395);
nand U5067 (N_5067,N_2685,N_4928);
nand U5068 (N_5068,N_3504,N_2239);
nand U5069 (N_5069,N_4301,N_414);
and U5070 (N_5070,N_2632,N_1798);
xor U5071 (N_5071,N_4578,N_719);
and U5072 (N_5072,N_3622,N_17);
xnor U5073 (N_5073,N_4168,N_2920);
xor U5074 (N_5074,N_4281,N_1316);
or U5075 (N_5075,N_1625,N_1454);
and U5076 (N_5076,N_1415,N_1030);
and U5077 (N_5077,N_3416,N_3775);
nand U5078 (N_5078,N_4609,N_219);
xor U5079 (N_5079,N_2249,N_3468);
nor U5080 (N_5080,N_2922,N_2030);
or U5081 (N_5081,N_4039,N_173);
or U5082 (N_5082,N_1232,N_3345);
and U5083 (N_5083,N_2263,N_1342);
nor U5084 (N_5084,N_3992,N_1664);
xor U5085 (N_5085,N_554,N_1171);
nand U5086 (N_5086,N_461,N_3609);
nand U5087 (N_5087,N_4990,N_312);
xnor U5088 (N_5088,N_854,N_3509);
and U5089 (N_5089,N_1472,N_4276);
or U5090 (N_5090,N_2400,N_762);
nor U5091 (N_5091,N_4147,N_245);
and U5092 (N_5092,N_1764,N_979);
nand U5093 (N_5093,N_4100,N_2772);
nand U5094 (N_5094,N_344,N_4241);
xnor U5095 (N_5095,N_4492,N_3139);
xnor U5096 (N_5096,N_124,N_697);
nand U5097 (N_5097,N_779,N_2069);
nor U5098 (N_5098,N_4243,N_1621);
xnor U5099 (N_5099,N_2536,N_2592);
or U5100 (N_5100,N_1533,N_4153);
and U5101 (N_5101,N_4128,N_597);
nor U5102 (N_5102,N_1384,N_1849);
or U5103 (N_5103,N_1792,N_2522);
and U5104 (N_5104,N_1105,N_3053);
and U5105 (N_5105,N_1932,N_4513);
or U5106 (N_5106,N_2240,N_3063);
nand U5107 (N_5107,N_4893,N_307);
and U5108 (N_5108,N_1005,N_4845);
nor U5109 (N_5109,N_3415,N_996);
and U5110 (N_5110,N_2755,N_2120);
nand U5111 (N_5111,N_3021,N_94);
xnor U5112 (N_5112,N_3145,N_2103);
and U5113 (N_5113,N_2430,N_568);
and U5114 (N_5114,N_1161,N_1726);
nand U5115 (N_5115,N_1401,N_3362);
nor U5116 (N_5116,N_1995,N_2107);
or U5117 (N_5117,N_1674,N_4657);
and U5118 (N_5118,N_2508,N_16);
or U5119 (N_5119,N_1513,N_2135);
and U5120 (N_5120,N_4993,N_614);
or U5121 (N_5121,N_2088,N_749);
or U5122 (N_5122,N_4035,N_2859);
or U5123 (N_5123,N_2917,N_2998);
or U5124 (N_5124,N_2594,N_4982);
nand U5125 (N_5125,N_1616,N_3618);
nand U5126 (N_5126,N_3024,N_2811);
and U5127 (N_5127,N_2899,N_4500);
nand U5128 (N_5128,N_3120,N_4806);
or U5129 (N_5129,N_3780,N_3955);
nand U5130 (N_5130,N_1469,N_3140);
nand U5131 (N_5131,N_3267,N_4758);
nand U5132 (N_5132,N_4519,N_1581);
nor U5133 (N_5133,N_33,N_1532);
xnor U5134 (N_5134,N_883,N_1385);
xor U5135 (N_5135,N_441,N_2642);
nand U5136 (N_5136,N_3430,N_2229);
xor U5137 (N_5137,N_2598,N_2775);
or U5138 (N_5138,N_1519,N_2394);
and U5139 (N_5139,N_274,N_4099);
xnor U5140 (N_5140,N_2606,N_163);
nor U5141 (N_5141,N_4569,N_831);
or U5142 (N_5142,N_292,N_255);
nor U5143 (N_5143,N_4499,N_4891);
xor U5144 (N_5144,N_4687,N_4828);
xnor U5145 (N_5145,N_1693,N_3383);
nand U5146 (N_5146,N_113,N_2050);
nand U5147 (N_5147,N_1334,N_343);
and U5148 (N_5148,N_1143,N_25);
nand U5149 (N_5149,N_1987,N_1955);
nand U5150 (N_5150,N_2327,N_651);
and U5151 (N_5151,N_299,N_2906);
nor U5152 (N_5152,N_4143,N_2876);
or U5153 (N_5153,N_477,N_994);
nand U5154 (N_5154,N_4584,N_3920);
and U5155 (N_5155,N_1748,N_176);
nor U5156 (N_5156,N_4068,N_2228);
or U5157 (N_5157,N_1322,N_3570);
nor U5158 (N_5158,N_3131,N_4413);
nor U5159 (N_5159,N_3358,N_780);
or U5160 (N_5160,N_1388,N_2934);
xnor U5161 (N_5161,N_4898,N_3183);
nand U5162 (N_5162,N_2346,N_1837);
or U5163 (N_5163,N_4506,N_3890);
nand U5164 (N_5164,N_4400,N_2881);
and U5165 (N_5165,N_4539,N_1942);
or U5166 (N_5166,N_2518,N_4227);
and U5167 (N_5167,N_214,N_2612);
or U5168 (N_5168,N_646,N_2910);
or U5169 (N_5169,N_2187,N_657);
or U5170 (N_5170,N_3898,N_2947);
or U5171 (N_5171,N_1058,N_2155);
nor U5172 (N_5172,N_4226,N_1700);
xnor U5173 (N_5173,N_3850,N_1651);
nand U5174 (N_5174,N_3248,N_3298);
or U5175 (N_5175,N_1079,N_3369);
nand U5176 (N_5176,N_2210,N_1000);
nand U5177 (N_5177,N_3793,N_7);
or U5178 (N_5178,N_4387,N_2316);
nand U5179 (N_5179,N_381,N_4603);
xnor U5180 (N_5180,N_2757,N_3541);
and U5181 (N_5181,N_259,N_1173);
and U5182 (N_5182,N_86,N_3175);
nor U5183 (N_5183,N_3089,N_639);
xnor U5184 (N_5184,N_1676,N_4007);
nand U5185 (N_5185,N_3070,N_3238);
and U5186 (N_5186,N_3719,N_2528);
or U5187 (N_5187,N_3442,N_2515);
and U5188 (N_5188,N_4551,N_3255);
xnor U5189 (N_5189,N_901,N_1588);
or U5190 (N_5190,N_1704,N_549);
xor U5191 (N_5191,N_2911,N_58);
xnor U5192 (N_5192,N_1220,N_3451);
or U5193 (N_5193,N_1425,N_4477);
nor U5194 (N_5194,N_1963,N_1575);
and U5195 (N_5195,N_3821,N_2014);
or U5196 (N_5196,N_4054,N_162);
nand U5197 (N_5197,N_2330,N_4736);
and U5198 (N_5198,N_701,N_856);
and U5199 (N_5199,N_4977,N_1245);
nand U5200 (N_5200,N_4171,N_1537);
nor U5201 (N_5201,N_1056,N_221);
nor U5202 (N_5202,N_1082,N_4232);
nand U5203 (N_5203,N_1249,N_638);
or U5204 (N_5204,N_3737,N_1543);
nand U5205 (N_5205,N_3249,N_2868);
nand U5206 (N_5206,N_1059,N_4187);
nor U5207 (N_5207,N_1284,N_1852);
and U5208 (N_5208,N_1025,N_4764);
nand U5209 (N_5209,N_2354,N_758);
and U5210 (N_5210,N_4055,N_795);
xnor U5211 (N_5211,N_4123,N_1808);
or U5212 (N_5212,N_1634,N_2506);
nor U5213 (N_5213,N_4694,N_4072);
and U5214 (N_5214,N_409,N_3185);
and U5215 (N_5215,N_4331,N_3022);
xnor U5216 (N_5216,N_2977,N_796);
xor U5217 (N_5217,N_843,N_770);
xnor U5218 (N_5218,N_3372,N_3321);
or U5219 (N_5219,N_3899,N_2909);
nand U5220 (N_5220,N_2305,N_3466);
or U5221 (N_5221,N_2426,N_4683);
nand U5222 (N_5222,N_281,N_2855);
or U5223 (N_5223,N_3460,N_2903);
nor U5224 (N_5224,N_3380,N_662);
nor U5225 (N_5225,N_422,N_846);
and U5226 (N_5226,N_2376,N_1742);
or U5227 (N_5227,N_1372,N_2753);
nor U5228 (N_5228,N_1571,N_1526);
xnor U5229 (N_5229,N_4860,N_1629);
xor U5230 (N_5230,N_3328,N_4163);
nor U5231 (N_5231,N_1751,N_2268);
and U5232 (N_5232,N_989,N_1004);
and U5233 (N_5233,N_1906,N_1179);
or U5234 (N_5234,N_2125,N_2495);
xor U5235 (N_5235,N_797,N_3130);
nor U5236 (N_5236,N_4254,N_3244);
or U5237 (N_5237,N_3276,N_570);
and U5238 (N_5238,N_4959,N_415);
or U5239 (N_5239,N_2488,N_2271);
and U5240 (N_5240,N_2016,N_1160);
xor U5241 (N_5241,N_1788,N_4491);
or U5242 (N_5242,N_3572,N_4752);
nor U5243 (N_5243,N_2060,N_2057);
or U5244 (N_5244,N_2778,N_2238);
and U5245 (N_5245,N_3212,N_4435);
nor U5246 (N_5246,N_4204,N_756);
xor U5247 (N_5247,N_4775,N_2458);
and U5248 (N_5248,N_4782,N_3475);
xnor U5249 (N_5249,N_155,N_3494);
or U5250 (N_5250,N_2424,N_1757);
or U5251 (N_5251,N_2819,N_863);
xor U5252 (N_5252,N_3915,N_3510);
xnor U5253 (N_5253,N_323,N_2277);
xor U5254 (N_5254,N_2258,N_3027);
and U5255 (N_5255,N_2956,N_4900);
and U5256 (N_5256,N_870,N_3364);
xnor U5257 (N_5257,N_1071,N_4394);
xor U5258 (N_5258,N_3958,N_4947);
and U5259 (N_5259,N_1531,N_1003);
or U5260 (N_5260,N_4695,N_669);
or U5261 (N_5261,N_2065,N_4798);
xor U5262 (N_5262,N_2608,N_1680);
or U5263 (N_5263,N_1124,N_419);
and U5264 (N_5264,N_2595,N_3660);
or U5265 (N_5265,N_3394,N_19);
or U5266 (N_5266,N_2555,N_1254);
and U5267 (N_5267,N_4293,N_4269);
nand U5268 (N_5268,N_4644,N_2625);
nand U5269 (N_5269,N_907,N_4377);
xnor U5270 (N_5270,N_1690,N_4345);
nand U5271 (N_5271,N_1560,N_4576);
and U5272 (N_5272,N_3492,N_2573);
nand U5273 (N_5273,N_87,N_151);
nor U5274 (N_5274,N_1424,N_2317);
xor U5275 (N_5275,N_8,N_4048);
nand U5276 (N_5276,N_1362,N_4997);
xnor U5277 (N_5277,N_2797,N_2599);
or U5278 (N_5278,N_2435,N_1294);
nand U5279 (N_5279,N_1278,N_1253);
or U5280 (N_5280,N_4218,N_2686);
nand U5281 (N_5281,N_3231,N_181);
xor U5282 (N_5282,N_3789,N_1248);
nor U5283 (N_5283,N_4749,N_4399);
or U5284 (N_5284,N_2979,N_3371);
xor U5285 (N_5285,N_3631,N_4188);
and U5286 (N_5286,N_4050,N_2022);
nand U5287 (N_5287,N_2476,N_1427);
nor U5288 (N_5288,N_4654,N_4800);
nand U5289 (N_5289,N_1701,N_3685);
xnor U5290 (N_5290,N_376,N_339);
xor U5291 (N_5291,N_2393,N_2201);
nor U5292 (N_5292,N_4840,N_4363);
and U5293 (N_5293,N_4235,N_2513);
nand U5294 (N_5294,N_872,N_518);
and U5295 (N_5295,N_4486,N_3455);
xnor U5296 (N_5296,N_4896,N_648);
and U5297 (N_5297,N_3686,N_1018);
nor U5298 (N_5298,N_3962,N_508);
or U5299 (N_5299,N_464,N_1091);
and U5300 (N_5300,N_4270,N_2688);
and U5301 (N_5301,N_4078,N_4027);
nor U5302 (N_5302,N_4481,N_2254);
or U5303 (N_5303,N_1477,N_190);
and U5304 (N_5304,N_297,N_2138);
xnor U5305 (N_5305,N_13,N_4961);
xor U5306 (N_5306,N_67,N_4323);
or U5307 (N_5307,N_4927,N_2081);
and U5308 (N_5308,N_3703,N_3757);
xnor U5309 (N_5309,N_2664,N_2603);
nand U5310 (N_5310,N_315,N_3613);
nand U5311 (N_5311,N_1732,N_3310);
or U5312 (N_5312,N_3161,N_3814);
and U5313 (N_5313,N_92,N_1406);
or U5314 (N_5314,N_4464,N_1020);
xor U5315 (N_5315,N_1439,N_3155);
nand U5316 (N_5316,N_1193,N_4597);
xnor U5317 (N_5317,N_1628,N_23);
xnor U5318 (N_5318,N_3597,N_193);
and U5319 (N_5319,N_4937,N_2337);
and U5320 (N_5320,N_2174,N_2163);
or U5321 (N_5321,N_4637,N_1196);
xnor U5322 (N_5322,N_1974,N_1936);
nand U5323 (N_5323,N_1389,N_2236);
nand U5324 (N_5324,N_4508,N_2856);
nand U5325 (N_5325,N_4441,N_480);
nor U5326 (N_5326,N_144,N_2894);
and U5327 (N_5327,N_4647,N_670);
or U5328 (N_5328,N_41,N_2214);
nor U5329 (N_5329,N_1501,N_1157);
xor U5330 (N_5330,N_2211,N_384);
and U5331 (N_5331,N_4643,N_3786);
nor U5332 (N_5332,N_1149,N_3528);
and U5333 (N_5333,N_2809,N_4032);
and U5334 (N_5334,N_4520,N_3457);
nand U5335 (N_5335,N_1373,N_1898);
xor U5336 (N_5336,N_1159,N_3444);
or U5337 (N_5337,N_4386,N_3359);
or U5338 (N_5338,N_4192,N_2777);
nand U5339 (N_5339,N_1654,N_246);
xor U5340 (N_5340,N_371,N_256);
xor U5341 (N_5341,N_1304,N_3315);
nor U5342 (N_5342,N_4976,N_4557);
and U5343 (N_5343,N_161,N_4839);
xnor U5344 (N_5344,N_3137,N_2764);
xnor U5345 (N_5345,N_2056,N_3171);
nor U5346 (N_5346,N_2441,N_3654);
nand U5347 (N_5347,N_1536,N_2086);
nand U5348 (N_5348,N_1781,N_926);
or U5349 (N_5349,N_4869,N_588);
xor U5350 (N_5350,N_3102,N_2250);
nand U5351 (N_5351,N_4599,N_2102);
xor U5352 (N_5352,N_2567,N_1414);
xor U5353 (N_5353,N_604,N_3530);
or U5354 (N_5354,N_3715,N_3797);
nand U5355 (N_5355,N_909,N_3254);
xnor U5356 (N_5356,N_2929,N_3050);
or U5357 (N_5357,N_822,N_4951);
nand U5358 (N_5358,N_2167,N_1793);
nor U5359 (N_5359,N_737,N_2212);
or U5360 (N_5360,N_2436,N_2864);
nor U5361 (N_5361,N_1260,N_4447);
and U5362 (N_5362,N_4468,N_1309);
nor U5363 (N_5363,N_3524,N_4022);
and U5364 (N_5364,N_1431,N_730);
nor U5365 (N_5365,N_1262,N_1842);
or U5366 (N_5366,N_2063,N_2298);
xor U5367 (N_5367,N_4240,N_411);
or U5368 (N_5368,N_3900,N_2615);
xor U5369 (N_5369,N_2110,N_1943);
xnor U5370 (N_5370,N_3341,N_2862);
or U5371 (N_5371,N_4859,N_4575);
nand U5372 (N_5372,N_3972,N_1247);
or U5373 (N_5373,N_3028,N_4601);
nor U5374 (N_5374,N_722,N_1933);
and U5375 (N_5375,N_4691,N_283);
nand U5376 (N_5376,N_2620,N_2530);
xor U5377 (N_5377,N_4784,N_1259);
xor U5378 (N_5378,N_2459,N_1463);
xnor U5379 (N_5379,N_956,N_3602);
or U5380 (N_5380,N_1484,N_1026);
or U5381 (N_5381,N_429,N_4586);
nor U5382 (N_5382,N_4822,N_3302);
or U5383 (N_5383,N_1035,N_985);
and U5384 (N_5384,N_1721,N_110);
nand U5385 (N_5385,N_4266,N_4850);
nor U5386 (N_5386,N_4428,N_4638);
nor U5387 (N_5387,N_2200,N_3262);
xor U5388 (N_5388,N_4527,N_1102);
nor U5389 (N_5389,N_3710,N_2494);
xor U5390 (N_5390,N_2472,N_4640);
and U5391 (N_5391,N_2915,N_1111);
nor U5392 (N_5392,N_4669,N_4214);
nand U5393 (N_5393,N_3834,N_4871);
or U5394 (N_5394,N_2546,N_3097);
nand U5395 (N_5395,N_1990,N_3658);
xnor U5396 (N_5396,N_3179,N_2444);
xnor U5397 (N_5397,N_2372,N_1008);
xor U5398 (N_5398,N_550,N_3208);
nand U5399 (N_5399,N_3656,N_1166);
xnor U5400 (N_5400,N_3877,N_3104);
or U5401 (N_5401,N_850,N_1587);
xnor U5402 (N_5402,N_4618,N_3352);
xnor U5403 (N_5403,N_4625,N_2111);
nand U5404 (N_5404,N_4696,N_3396);
nand U5405 (N_5405,N_472,N_3800);
nor U5406 (N_5406,N_1135,N_2692);
and U5407 (N_5407,N_2351,N_2213);
xor U5408 (N_5408,N_1522,N_4745);
nor U5409 (N_5409,N_1662,N_2429);
or U5410 (N_5410,N_4761,N_2533);
nor U5411 (N_5411,N_2044,N_1214);
nand U5412 (N_5412,N_2269,N_1601);
nor U5413 (N_5413,N_2829,N_3088);
xor U5414 (N_5414,N_814,N_2743);
nor U5415 (N_5415,N_4979,N_126);
and U5416 (N_5416,N_602,N_1636);
or U5417 (N_5417,N_2175,N_4167);
nor U5418 (N_5418,N_818,N_3426);
or U5419 (N_5419,N_3984,N_427);
nand U5420 (N_5420,N_4368,N_2410);
or U5421 (N_5421,N_3343,N_1724);
xor U5422 (N_5422,N_4327,N_813);
and U5423 (N_5423,N_3356,N_3989);
nor U5424 (N_5424,N_4910,N_4907);
and U5425 (N_5425,N_1529,N_322);
nor U5426 (N_5426,N_3599,N_102);
nand U5427 (N_5427,N_839,N_3496);
nand U5428 (N_5428,N_3393,N_1848);
nor U5429 (N_5429,N_4579,N_3785);
and U5430 (N_5430,N_3577,N_1789);
nand U5431 (N_5431,N_4524,N_922);
and U5432 (N_5432,N_3291,N_2725);
and U5433 (N_5433,N_906,N_1712);
or U5434 (N_5434,N_1502,N_1189);
nor U5435 (N_5435,N_3092,N_4941);
or U5436 (N_5436,N_327,N_1274);
or U5437 (N_5437,N_3354,N_3589);
or U5438 (N_5438,N_4103,N_1491);
and U5439 (N_5439,N_4556,N_2966);
or U5440 (N_5440,N_1224,N_2651);
and U5441 (N_5441,N_373,N_202);
and U5442 (N_5442,N_1807,N_1381);
xnor U5443 (N_5443,N_4217,N_3118);
and U5444 (N_5444,N_2468,N_2011);
xnor U5445 (N_5445,N_447,N_1811);
xor U5446 (N_5446,N_2641,N_417);
or U5447 (N_5447,N_2395,N_3742);
or U5448 (N_5448,N_675,N_2521);
xor U5449 (N_5449,N_2153,N_1517);
nor U5450 (N_5450,N_3760,N_3497);
xnor U5451 (N_5451,N_936,N_2611);
or U5452 (N_5452,N_2680,N_2313);
xor U5453 (N_5453,N_984,N_1663);
nand U5454 (N_5454,N_1813,N_3236);
xnor U5455 (N_5455,N_1100,N_4440);
xnor U5456 (N_5456,N_1313,N_308);
and U5457 (N_5457,N_3191,N_3441);
and U5458 (N_5458,N_2283,N_700);
or U5459 (N_5459,N_1720,N_4472);
or U5460 (N_5460,N_150,N_4746);
xnor U5461 (N_5461,N_3007,N_1735);
nand U5462 (N_5462,N_690,N_3848);
nand U5463 (N_5463,N_4182,N_1233);
nor U5464 (N_5464,N_4023,N_2689);
or U5465 (N_5465,N_2556,N_2134);
or U5466 (N_5466,N_1800,N_1882);
nor U5467 (N_5467,N_3193,N_3199);
nor U5468 (N_5468,N_2477,N_4157);
nand U5469 (N_5469,N_1349,N_4229);
xnor U5470 (N_5470,N_3127,N_2945);
nor U5471 (N_5471,N_745,N_4414);
xor U5472 (N_5472,N_346,N_1235);
nor U5473 (N_5473,N_627,N_3844);
nor U5474 (N_5474,N_887,N_3368);
or U5475 (N_5475,N_4203,N_1413);
nand U5476 (N_5476,N_3096,N_4335);
nor U5477 (N_5477,N_1877,N_4936);
or U5478 (N_5478,N_621,N_2918);
nor U5479 (N_5479,N_3339,N_2364);
and U5480 (N_5480,N_1473,N_1550);
xnor U5481 (N_5481,N_2259,N_444);
nand U5482 (N_5482,N_2027,N_628);
nor U5483 (N_5483,N_4783,N_1398);
nor U5484 (N_5484,N_4705,N_247);
or U5485 (N_5485,N_2813,N_4626);
nand U5486 (N_5486,N_548,N_1935);
nor U5487 (N_5487,N_4821,N_1243);
and U5488 (N_5488,N_4968,N_747);
nor U5489 (N_5489,N_3195,N_402);
and U5490 (N_5490,N_1780,N_2405);
and U5491 (N_5491,N_2880,N_4915);
nor U5492 (N_5492,N_1039,N_3033);
xor U5493 (N_5493,N_1604,N_492);
nand U5494 (N_5494,N_4081,N_1350);
nor U5495 (N_5495,N_2784,N_3031);
xor U5496 (N_5496,N_2671,N_2090);
nand U5497 (N_5497,N_2098,N_1044);
or U5498 (N_5498,N_3873,N_3370);
and U5499 (N_5499,N_2795,N_4089);
and U5500 (N_5500,N_4887,N_2350);
nand U5501 (N_5501,N_112,N_692);
and U5502 (N_5502,N_3057,N_4260);
xor U5503 (N_5503,N_4501,N_1535);
and U5504 (N_5504,N_4053,N_3068);
or U5505 (N_5505,N_434,N_4033);
xnor U5506 (N_5506,N_3881,N_1154);
nor U5507 (N_5507,N_3474,N_4837);
xor U5508 (N_5508,N_595,N_2024);
or U5509 (N_5509,N_4518,N_4256);
xnor U5510 (N_5510,N_4562,N_1846);
or U5511 (N_5511,N_3489,N_3075);
or U5512 (N_5512,N_2936,N_2541);
and U5513 (N_5513,N_3857,N_2362);
or U5514 (N_5514,N_2485,N_1038);
xor U5515 (N_5515,N_4734,N_869);
or U5516 (N_5516,N_2055,N_2121);
xnor U5517 (N_5517,N_2370,N_4791);
xor U5518 (N_5518,N_2991,N_4397);
xnor U5519 (N_5519,N_342,N_4410);
nor U5520 (N_5520,N_4372,N_1023);
nand U5521 (N_5521,N_2663,N_1212);
and U5522 (N_5522,N_4854,N_4946);
or U5523 (N_5523,N_2916,N_1392);
and U5524 (N_5524,N_900,N_90);
or U5525 (N_5525,N_1619,N_2366);
nor U5526 (N_5526,N_3280,N_4322);
or U5527 (N_5527,N_340,N_3389);
or U5528 (N_5528,N_3619,N_2445);
nor U5529 (N_5529,N_1868,N_3993);
and U5530 (N_5530,N_206,N_2073);
or U5531 (N_5531,N_3750,N_1779);
xnor U5532 (N_5532,N_4747,N_4344);
nor U5533 (N_5533,N_753,N_3713);
or U5534 (N_5534,N_2748,N_4658);
nand U5535 (N_5535,N_204,N_85);
nor U5536 (N_5536,N_966,N_3614);
or U5537 (N_5537,N_3729,N_3052);
nor U5538 (N_5538,N_3573,N_1246);
xnor U5539 (N_5539,N_4834,N_899);
and U5540 (N_5540,N_3943,N_4268);
nor U5541 (N_5541,N_230,N_1773);
and U5542 (N_5542,N_1266,N_693);
and U5543 (N_5543,N_1325,N_3592);
xnor U5544 (N_5544,N_4351,N_1272);
nand U5545 (N_5545,N_4442,N_1617);
nor U5546 (N_5546,N_2950,N_104);
nand U5547 (N_5547,N_1308,N_2028);
and U5548 (N_5548,N_2818,N_2766);
or U5549 (N_5549,N_1699,N_3644);
nor U5550 (N_5550,N_2177,N_3628);
and U5551 (N_5551,N_1640,N_1754);
nor U5552 (N_5552,N_1648,N_228);
nand U5553 (N_5553,N_4245,N_3260);
or U5554 (N_5554,N_3519,N_809);
xnor U5555 (N_5555,N_2836,N_3471);
xnor U5556 (N_5556,N_4052,N_205);
nor U5557 (N_5557,N_4130,N_2768);
or U5558 (N_5558,N_2800,N_399);
nand U5559 (N_5559,N_1734,N_4096);
nand U5560 (N_5560,N_2463,N_4911);
nand U5561 (N_5561,N_4801,N_2493);
xnor U5562 (N_5562,N_988,N_309);
and U5563 (N_5563,N_2363,N_4743);
nand U5564 (N_5564,N_2181,N_2981);
xor U5565 (N_5565,N_2581,N_2418);
or U5566 (N_5566,N_1727,N_433);
and U5567 (N_5567,N_4006,N_4057);
nand U5568 (N_5568,N_24,N_4333);
or U5569 (N_5569,N_4403,N_3428);
nor U5570 (N_5570,N_2785,N_4537);
xor U5571 (N_5571,N_2803,N_4570);
or U5572 (N_5572,N_4697,N_3287);
and U5573 (N_5573,N_1505,N_3624);
xor U5574 (N_5574,N_4086,N_4150);
and U5575 (N_5575,N_4304,N_4367);
nor U5576 (N_5576,N_4855,N_2532);
nor U5577 (N_5577,N_2782,N_4984);
nand U5578 (N_5578,N_2794,N_1099);
or U5579 (N_5579,N_1585,N_535);
nor U5580 (N_5580,N_2507,N_3126);
and U5581 (N_5581,N_4176,N_4267);
xnor U5582 (N_5582,N_3674,N_3136);
and U5583 (N_5583,N_4141,N_135);
and U5584 (N_5584,N_547,N_3187);
nor U5585 (N_5585,N_3904,N_3913);
xor U5586 (N_5586,N_3952,N_1694);
nand U5587 (N_5587,N_4185,N_445);
nand U5588 (N_5588,N_1775,N_2217);
nor U5589 (N_5589,N_3764,N_650);
nor U5590 (N_5590,N_4220,N_3274);
nor U5591 (N_5591,N_3080,N_2810);
or U5592 (N_5592,N_325,N_2161);
nand U5593 (N_5593,N_4149,N_4865);
nor U5594 (N_5594,N_2720,N_1191);
or U5595 (N_5595,N_1772,N_1192);
xnor U5596 (N_5596,N_864,N_1633);
xor U5597 (N_5597,N_2043,N_537);
nor U5598 (N_5598,N_3446,N_2993);
xor U5599 (N_5599,N_4152,N_2425);
nor U5600 (N_5600,N_3590,N_3991);
nor U5601 (N_5601,N_288,N_649);
xnor U5602 (N_5602,N_4380,N_3584);
xor U5603 (N_5603,N_2002,N_3880);
or U5604 (N_5604,N_3122,N_3935);
nor U5605 (N_5605,N_3828,N_4862);
and U5606 (N_5606,N_1538,N_787);
or U5607 (N_5607,N_2064,N_3555);
or U5608 (N_5608,N_4666,N_1610);
nor U5609 (N_5609,N_4036,N_1273);
nor U5610 (N_5610,N_316,N_4938);
nor U5611 (N_5611,N_1816,N_4317);
or U5612 (N_5612,N_3776,N_534);
nand U5613 (N_5613,N_1624,N_1796);
nor U5614 (N_5614,N_1746,N_4650);
xor U5615 (N_5615,N_2806,N_4355);
or U5616 (N_5616,N_107,N_421);
nand U5617 (N_5617,N_1032,N_4738);
xor U5618 (N_5618,N_1835,N_4411);
xnor U5619 (N_5619,N_2652,N_1886);
nor U5620 (N_5620,N_3652,N_2007);
nor U5621 (N_5621,N_2108,N_4934);
nand U5622 (N_5622,N_4574,N_4682);
or U5623 (N_5623,N_4932,N_2178);
nor U5624 (N_5624,N_2257,N_1561);
and U5625 (N_5625,N_504,N_2558);
or U5626 (N_5626,N_585,N_3748);
or U5627 (N_5627,N_1125,N_1051);
xnor U5628 (N_5628,N_4525,N_1857);
or U5629 (N_5629,N_4581,N_905);
nand U5630 (N_5630,N_147,N_3182);
or U5631 (N_5631,N_618,N_2075);
and U5632 (N_5632,N_1762,N_2774);
and U5633 (N_5633,N_2634,N_3564);
or U5634 (N_5634,N_234,N_4393);
and U5635 (N_5635,N_4450,N_1267);
or U5636 (N_5636,N_375,N_4895);
xor U5637 (N_5637,N_4299,N_3400);
xor U5638 (N_5638,N_4794,N_3493);
xor U5639 (N_5639,N_4550,N_1016);
nor U5640 (N_5640,N_4140,N_4431);
nor U5641 (N_5641,N_2889,N_1393);
nor U5642 (N_5642,N_2552,N_4876);
and U5643 (N_5643,N_4656,N_3808);
xnor U5644 (N_5644,N_1681,N_728);
and U5645 (N_5645,N_2419,N_4545);
nor U5646 (N_5646,N_3896,N_2923);
nor U5647 (N_5647,N_4202,N_3743);
and U5648 (N_5648,N_4222,N_1172);
or U5649 (N_5649,N_2962,N_1507);
or U5650 (N_5650,N_2718,N_318);
nor U5651 (N_5651,N_233,N_727);
xor U5652 (N_5652,N_2001,N_2559);
xnor U5653 (N_5653,N_2708,N_4016);
and U5654 (N_5654,N_629,N_1217);
or U5655 (N_5655,N_4899,N_3125);
or U5656 (N_5656,N_239,N_1911);
nand U5657 (N_5657,N_3970,N_946);
nand U5658 (N_5658,N_507,N_1622);
xor U5659 (N_5659,N_2094,N_999);
nor U5660 (N_5660,N_2566,N_3895);
and U5661 (N_5661,N_696,N_1289);
and U5662 (N_5662,N_1874,N_4114);
and U5663 (N_5663,N_1437,N_2159);
nor U5664 (N_5664,N_3771,N_4164);
or U5665 (N_5665,N_4874,N_2189);
or U5666 (N_5666,N_1239,N_357);
or U5667 (N_5667,N_1763,N_1364);
or U5668 (N_5668,N_541,N_295);
or U5669 (N_5669,N_4838,N_1630);
and U5670 (N_5670,N_3988,N_3085);
or U5671 (N_5671,N_545,N_437);
nand U5672 (N_5672,N_2504,N_521);
xor U5673 (N_5673,N_4158,N_2246);
xnor U5674 (N_5674,N_2801,N_3111);
xnor U5675 (N_5675,N_4565,N_3035);
nor U5676 (N_5676,N_287,N_4077);
nand U5677 (N_5677,N_1148,N_1185);
xor U5678 (N_5678,N_792,N_2194);
and U5679 (N_5679,N_1758,N_3670);
nand U5680 (N_5680,N_254,N_4004);
nand U5681 (N_5681,N_2384,N_3999);
or U5682 (N_5682,N_2483,N_4487);
and U5683 (N_5683,N_1947,N_3218);
xnor U5684 (N_5684,N_499,N_1132);
nand U5685 (N_5685,N_2600,N_4890);
xnor U5686 (N_5686,N_3629,N_2804);
nor U5687 (N_5687,N_3672,N_2902);
nor U5688 (N_5688,N_330,N_4233);
xnor U5689 (N_5689,N_4420,N_1487);
nand U5690 (N_5690,N_4593,N_4739);
and U5691 (N_5691,N_4415,N_741);
nand U5692 (N_5692,N_2068,N_2735);
nand U5693 (N_5693,N_4230,N_708);
and U5694 (N_5694,N_524,N_3617);
xnor U5695 (N_5695,N_666,N_3856);
and U5696 (N_5696,N_3661,N_4948);
nor U5697 (N_5697,N_2180,N_109);
xnor U5698 (N_5698,N_1285,N_4422);
or U5699 (N_5699,N_3294,N_4146);
and U5700 (N_5700,N_765,N_1671);
and U5701 (N_5701,N_2828,N_4608);
xor U5702 (N_5702,N_4605,N_260);
xnor U5703 (N_5703,N_526,N_4272);
or U5704 (N_5704,N_3998,N_3807);
or U5705 (N_5705,N_4309,N_275);
xnor U5706 (N_5706,N_2883,N_4978);
and U5707 (N_5707,N_4848,N_396);
xnor U5708 (N_5708,N_4255,N_1900);
xor U5709 (N_5709,N_2563,N_4832);
xnor U5710 (N_5710,N_18,N_4962);
and U5711 (N_5711,N_4846,N_185);
xor U5712 (N_5712,N_1174,N_2397);
nand U5713 (N_5713,N_424,N_3135);
nor U5714 (N_5714,N_3862,N_4124);
and U5715 (N_5715,N_3210,N_2438);
nor U5716 (N_5716,N_3911,N_3011);
and U5717 (N_5717,N_4195,N_4595);
and U5718 (N_5718,N_271,N_3861);
or U5719 (N_5719,N_183,N_790);
xnor U5720 (N_5720,N_4750,N_2550);
and U5721 (N_5721,N_82,N_4189);
nand U5722 (N_5722,N_1404,N_2484);
and U5723 (N_5723,N_4318,N_1187);
or U5724 (N_5724,N_3232,N_103);
and U5725 (N_5725,N_2047,N_2339);
xor U5726 (N_5726,N_4776,N_4831);
or U5727 (N_5727,N_1047,N_1844);
nor U5728 (N_5728,N_967,N_743);
nand U5729 (N_5729,N_4681,N_4329);
and U5730 (N_5730,N_3105,N_4731);
nand U5731 (N_5731,N_2815,N_3066);
and U5732 (N_5732,N_226,N_586);
nand U5733 (N_5733,N_3740,N_1922);
nor U5734 (N_5734,N_4265,N_3885);
nor U5735 (N_5735,N_1964,N_1678);
nor U5736 (N_5736,N_4505,N_4526);
and U5737 (N_5737,N_3361,N_3237);
xnor U5738 (N_5738,N_2690,N_408);
or U5739 (N_5739,N_1055,N_413);
xnor U5740 (N_5740,N_3995,N_4066);
or U5741 (N_5741,N_2799,N_3693);
xor U5742 (N_5742,N_3684,N_156);
nor U5743 (N_5743,N_69,N_3042);
xnor U5744 (N_5744,N_4352,N_1444);
xnor U5745 (N_5745,N_1967,N_1710);
and U5746 (N_5746,N_2165,N_1658);
and U5747 (N_5747,N_3870,N_3002);
xnor U5748 (N_5748,N_3914,N_4824);
xor U5749 (N_5749,N_3974,N_4805);
or U5750 (N_5750,N_3392,N_4137);
xnor U5751 (N_5751,N_2374,N_3367);
nand U5752 (N_5752,N_2322,N_4760);
or U5753 (N_5753,N_2695,N_290);
and U5754 (N_5754,N_1104,N_332);
nand U5755 (N_5755,N_3041,N_2008);
and U5756 (N_5756,N_1921,N_91);
or U5757 (N_5757,N_1048,N_2733);
nand U5758 (N_5758,N_1797,N_1767);
or U5759 (N_5759,N_4702,N_3600);
and U5760 (N_5760,N_2404,N_4634);
and U5761 (N_5761,N_724,N_2630);
nand U5762 (N_5762,N_2389,N_2169);
or U5763 (N_5763,N_4533,N_1064);
and U5764 (N_5764,N_2691,N_4727);
xor U5765 (N_5765,N_377,N_1061);
and U5766 (N_5766,N_4778,N_1608);
xnor U5767 (N_5767,N_3346,N_1287);
or U5768 (N_5768,N_2119,N_232);
or U5769 (N_5769,N_785,N_1277);
or U5770 (N_5770,N_3012,N_9);
xnor U5771 (N_5771,N_998,N_731);
xnor U5772 (N_5772,N_1706,N_884);
or U5773 (N_5773,N_3116,N_920);
nand U5774 (N_5774,N_3583,N_2202);
xor U5775 (N_5775,N_2670,N_2887);
and U5776 (N_5776,N_3901,N_4105);
and U5777 (N_5777,N_3424,N_3323);
and U5778 (N_5778,N_2564,N_1542);
nor U5779 (N_5779,N_4585,N_1354);
or U5780 (N_5780,N_590,N_3003);
and U5781 (N_5781,N_620,N_1810);
nand U5782 (N_5782,N_2844,N_3351);
xnor U5783 (N_5783,N_4257,N_3735);
nor U5784 (N_5784,N_4802,N_1635);
nor U5785 (N_5785,N_2792,N_2839);
and U5786 (N_5786,N_210,N_617);
or U5787 (N_5787,N_973,N_317);
nand U5788 (N_5788,N_4478,N_4720);
and U5789 (N_5789,N_356,N_1769);
or U5790 (N_5790,N_1918,N_4253);
and U5791 (N_5791,N_1518,N_2199);
nor U5792 (N_5792,N_1697,N_1885);
or U5793 (N_5793,N_1818,N_3049);
xor U5794 (N_5794,N_4918,N_3997);
and U5795 (N_5795,N_1723,N_3726);
and U5796 (N_5796,N_3853,N_2681);
nor U5797 (N_5797,N_1386,N_3687);
nor U5798 (N_5798,N_21,N_191);
and U5799 (N_5799,N_3337,N_3511);
nor U5800 (N_5800,N_4972,N_1458);
xor U5801 (N_5801,N_4944,N_3447);
nor U5802 (N_5802,N_2373,N_3957);
nor U5803 (N_5803,N_2193,N_4986);
nand U5804 (N_5804,N_695,N_1623);
and U5805 (N_5805,N_1409,N_845);
and U5806 (N_5806,N_1859,N_1396);
nand U5807 (N_5807,N_2020,N_4374);
nor U5808 (N_5808,N_2683,N_4373);
nor U5809 (N_5809,N_2647,N_2332);
xor U5810 (N_5810,N_3407,N_3173);
or U5811 (N_5811,N_3350,N_3168);
and U5812 (N_5812,N_400,N_1092);
or U5813 (N_5813,N_89,N_3831);
or U5814 (N_5814,N_1783,N_2816);
xor U5815 (N_5815,N_4945,N_3539);
and U5816 (N_5816,N_1530,N_133);
and U5817 (N_5817,N_4851,N_1820);
nor U5818 (N_5818,N_501,N_3094);
nand U5819 (N_5819,N_4957,N_483);
xor U5820 (N_5820,N_2266,N_4692);
nor U5821 (N_5821,N_1665,N_663);
or U5822 (N_5822,N_2988,N_2052);
nor U5823 (N_5823,N_587,N_4336);
or U5824 (N_5824,N_2739,N_3603);
nor U5825 (N_5825,N_3700,N_788);
xor U5826 (N_5826,N_1641,N_1545);
and U5827 (N_5827,N_3263,N_370);
xor U5828 (N_5828,N_1108,N_2371);
or U5829 (N_5829,N_576,N_4091);
and U5830 (N_5830,N_1855,N_1209);
nor U5831 (N_5831,N_1562,N_3087);
nor U5832 (N_5832,N_1255,N_2745);
nor U5833 (N_5833,N_3463,N_871);
or U5834 (N_5834,N_3933,N_298);
or U5835 (N_5835,N_3178,N_1040);
xor U5836 (N_5836,N_2227,N_704);
xnor U5837 (N_5837,N_137,N_3349);
nor U5838 (N_5838,N_1856,N_301);
and U5839 (N_5839,N_2005,N_1864);
or U5840 (N_5840,N_1027,N_2593);
nand U5841 (N_5841,N_3072,N_3659);
xnor U5842 (N_5842,N_622,N_4950);
and U5843 (N_5843,N_2455,N_2385);
and U5844 (N_5844,N_4277,N_3837);
nor U5845 (N_5845,N_2841,N_3538);
and U5846 (N_5846,N_644,N_2953);
xnor U5847 (N_5847,N_3100,N_3452);
nand U5848 (N_5848,N_4291,N_1657);
xor U5849 (N_5849,N_51,N_3293);
and U5850 (N_5850,N_1743,N_4648);
nand U5851 (N_5851,N_1017,N_3286);
and U5852 (N_5852,N_4635,N_3611);
xnor U5853 (N_5853,N_3241,N_510);
or U5854 (N_5854,N_4328,N_1832);
nand U5855 (N_5855,N_2721,N_3230);
nor U5856 (N_5856,N_929,N_821);
or U5857 (N_5857,N_3414,N_4402);
or U5858 (N_5858,N_4456,N_2264);
xnor U5859 (N_5859,N_4223,N_97);
or U5860 (N_5860,N_4612,N_4194);
nand U5861 (N_5861,N_1452,N_4920);
and U5862 (N_5862,N_3815,N_3151);
and U5863 (N_5863,N_2017,N_2763);
nor U5864 (N_5864,N_2497,N_566);
nand U5865 (N_5865,N_2038,N_3633);
or U5866 (N_5866,N_4878,N_4885);
nand U5867 (N_5867,N_159,N_4237);
or U5868 (N_5868,N_1838,N_4443);
and U5869 (N_5869,N_100,N_1347);
xor U5870 (N_5870,N_3515,N_2571);
xnor U5871 (N_5871,N_2904,N_4170);
nor U5872 (N_5872,N_4958,N_2627);
xor U5873 (N_5873,N_1756,N_4512);
nor U5874 (N_5874,N_1824,N_551);
nand U5875 (N_5875,N_3229,N_3038);
and U5876 (N_5876,N_671,N_3947);
xor U5877 (N_5877,N_2890,N_207);
xor U5878 (N_5878,N_3439,N_390);
nand U5879 (N_5879,N_951,N_4725);
xnor U5880 (N_5880,N_157,N_2139);
and U5881 (N_5881,N_4534,N_2919);
xnor U5882 (N_5882,N_3078,N_810);
or U5883 (N_5883,N_1825,N_3707);
nand U5884 (N_5884,N_1435,N_710);
or U5885 (N_5885,N_3811,N_1479);
and U5886 (N_5886,N_1854,N_1656);
and U5887 (N_5887,N_4289,N_2851);
nor U5888 (N_5888,N_2891,N_2983);
xnor U5889 (N_5889,N_4113,N_418);
and U5890 (N_5890,N_2010,N_3925);
nand U5891 (N_5891,N_3077,N_3454);
xor U5892 (N_5892,N_3657,N_1905);
nand U5893 (N_5893,N_4286,N_1867);
nor U5894 (N_5894,N_897,N_454);
nor U5895 (N_5895,N_1296,N_2012);
nand U5896 (N_5896,N_2415,N_517);
xnor U5897 (N_5897,N_592,N_1890);
nand U5898 (N_5898,N_4,N_3313);
nor U5899 (N_5899,N_4715,N_22);
nor U5900 (N_5900,N_2253,N_3180);
or U5901 (N_5901,N_3117,N_619);
nand U5902 (N_5902,N_1011,N_1552);
nand U5903 (N_5903,N_4923,N_2326);
xor U5904 (N_5904,N_2359,N_3745);
nor U5905 (N_5905,N_4302,N_4426);
nand U5906 (N_5906,N_2744,N_4315);
nor U5907 (N_5907,N_2543,N_3876);
xor U5908 (N_5908,N_3731,N_3079);
or U5909 (N_5909,N_4732,N_2783);
or U5910 (N_5910,N_2531,N_4541);
nand U5911 (N_5911,N_2255,N_1652);
and U5912 (N_5912,N_1627,N_3845);
nor U5913 (N_5913,N_1576,N_4566);
nor U5914 (N_5914,N_3960,N_277);
or U5915 (N_5915,N_4308,N_2137);
or U5916 (N_5916,N_3948,N_240);
and U5917 (N_5917,N_175,N_3551);
nor U5918 (N_5918,N_1985,N_4412);
or U5919 (N_5919,N_3867,N_241);
or U5920 (N_5920,N_2931,N_3824);
and U5921 (N_5921,N_4358,N_1805);
nand U5922 (N_5922,N_1930,N_2095);
or U5923 (N_5923,N_3219,N_1821);
or U5924 (N_5924,N_4906,N_160);
xor U5925 (N_5925,N_514,N_1298);
xnor U5926 (N_5926,N_2607,N_2793);
nand U5927 (N_5927,N_891,N_4742);
and U5928 (N_5928,N_1050,N_1999);
or U5929 (N_5929,N_2147,N_3324);
or U5930 (N_5930,N_2117,N_1407);
nor U5931 (N_5931,N_1814,N_1083);
nand U5932 (N_5932,N_4295,N_257);
nand U5933 (N_5933,N_1696,N_4076);
or U5934 (N_5934,N_1208,N_820);
nand U5935 (N_5935,N_3711,N_4065);
and U5936 (N_5936,N_4488,N_2375);
nor U5937 (N_5937,N_4868,N_153);
or U5938 (N_5938,N_630,N_4396);
nor U5939 (N_5939,N_3521,N_886);
xnor U5940 (N_5940,N_2072,N_293);
or U5941 (N_5941,N_865,N_2281);
nor U5942 (N_5942,N_2006,N_4810);
nor U5943 (N_5943,N_733,N_2114);
or U5944 (N_5944,N_711,N_3440);
and U5945 (N_5945,N_3918,N_520);
nand U5946 (N_5946,N_3001,N_1753);
nand U5947 (N_5947,N_610,N_702);
xnor U5948 (N_5948,N_3335,N_3545);
and U5949 (N_5949,N_2677,N_1851);
or U5950 (N_5950,N_958,N_2469);
or U5951 (N_5951,N_1714,N_677);
or U5952 (N_5952,N_596,N_4594);
and U5953 (N_5953,N_4013,N_2519);
or U5954 (N_5954,N_2208,N_2335);
xnor U5955 (N_5955,N_4528,N_3469);
and U5956 (N_5956,N_4173,N_1033);
nor U5957 (N_5957,N_4744,N_1200);
and U5958 (N_5958,N_1466,N_2401);
xor U5959 (N_5959,N_1679,N_450);
nor U5960 (N_5960,N_2617,N_2130);
xnor U5961 (N_5961,N_4332,N_1357);
nor U5962 (N_5962,N_4975,N_4816);
nand U5963 (N_5963,N_363,N_3692);
nor U5964 (N_5964,N_2183,N_2341);
xnor U5965 (N_5965,N_2802,N_4339);
or U5966 (N_5966,N_2523,N_1408);
and U5967 (N_5967,N_3121,N_4132);
xnor U5968 (N_5968,N_685,N_2413);
and U5969 (N_5969,N_1380,N_528);
nand U5970 (N_5970,N_2379,N_1703);
xor U5971 (N_5971,N_2383,N_3812);
and U5972 (N_5972,N_1613,N_2656);
xor U5973 (N_5973,N_129,N_188);
nand U5974 (N_5974,N_3987,N_491);
or U5975 (N_5975,N_331,N_1355);
nand U5976 (N_5976,N_761,N_3409);
nor U5977 (N_5977,N_1959,N_4571);
nor U5978 (N_5978,N_3841,N_324);
and U5979 (N_5979,N_3549,N_2940);
nor U5980 (N_5980,N_3157,N_237);
nor U5981 (N_5981,N_3266,N_766);
nor U5982 (N_5982,N_713,N_2319);
nor U5983 (N_5983,N_2233,N_4909);
and U5984 (N_5984,N_395,N_2935);
and U5985 (N_5985,N_715,N_2478);
and U5986 (N_5986,N_4721,N_1572);
or U5987 (N_5987,N_771,N_3535);
nand U5988 (N_5988,N_2752,N_1010);
nand U5989 (N_5989,N_3170,N_4903);
and U5990 (N_5990,N_3176,N_451);
nand U5991 (N_5991,N_3290,N_3638);
and U5992 (N_5992,N_2616,N_273);
nand U5993 (N_5993,N_3769,N_4552);
xor U5994 (N_5994,N_378,N_1118);
nor U5995 (N_5995,N_2830,N_2654);
and U5996 (N_5996,N_2732,N_2585);
or U5997 (N_5997,N_4572,N_2992);
xor U5998 (N_5998,N_2128,N_3423);
xor U5999 (N_5999,N_1916,N_1338);
nand U6000 (N_6000,N_360,N_3980);
xnor U6001 (N_6001,N_52,N_1553);
xnor U6002 (N_6002,N_653,N_2781);
nand U6003 (N_6003,N_1929,N_740);
and U6004 (N_6004,N_862,N_2026);
nand U6005 (N_6005,N_2900,N_1078);
or U6006 (N_6006,N_1770,N_2572);
xor U6007 (N_6007,N_1115,N_995);
nand U6008 (N_6008,N_718,N_3975);
nand U6009 (N_6009,N_4762,N_4406);
and U6010 (N_6010,N_2674,N_645);
xnor U6011 (N_6011,N_881,N_1194);
xor U6012 (N_6012,N_2925,N_990);
or U6013 (N_6013,N_4685,N_2031);
nor U6014 (N_6014,N_563,N_3278);
and U6015 (N_6015,N_3464,N_1826);
nand U6016 (N_6016,N_1937,N_348);
and U6017 (N_6017,N_3384,N_705);
nor U6018 (N_6018,N_3247,N_78);
nor U6019 (N_6019,N_565,N_1197);
or U6020 (N_6020,N_1410,N_1403);
nor U6021 (N_6021,N_252,N_225);
nor U6022 (N_6022,N_2588,N_4401);
xor U6023 (N_6023,N_1884,N_4913);
xnor U6024 (N_6024,N_223,N_2845);
xnor U6025 (N_6025,N_1829,N_698);
xnor U6026 (N_6026,N_2053,N_889);
nor U6027 (N_6027,N_1686,N_511);
nor U6028 (N_6028,N_265,N_4511);
and U6029 (N_6029,N_1755,N_3025);
nand U6030 (N_6030,N_4954,N_1819);
nor U6031 (N_6031,N_1280,N_2758);
nand U6032 (N_6032,N_672,N_4676);
and U6033 (N_6033,N_3054,N_3376);
nor U6034 (N_6034,N_3953,N_2083);
and U6035 (N_6035,N_3796,N_552);
nand U6036 (N_6036,N_1002,N_1598);
xor U6037 (N_6037,N_1761,N_4273);
nand U6038 (N_6038,N_4228,N_2);
nor U6039 (N_6039,N_2129,N_1899);
nor U6040 (N_6040,N_2990,N_1069);
nand U6041 (N_6041,N_3529,N_3486);
or U6042 (N_6042,N_4088,N_2396);
nand U6043 (N_6043,N_4825,N_2629);
xor U6044 (N_6044,N_341,N_1109);
and U6045 (N_6045,N_4779,N_3108);
nor U6046 (N_6046,N_4129,N_4879);
or U6047 (N_6047,N_561,N_1087);
and U6048 (N_6048,N_2096,N_2714);
xor U6049 (N_6049,N_2242,N_4430);
and U6050 (N_6050,N_970,N_1448);
xnor U6051 (N_6051,N_4433,N_4974);
or U6052 (N_6052,N_1299,N_4310);
nor U6053 (N_6053,N_1374,N_4193);
and U6054 (N_6054,N_2289,N_4614);
and U6055 (N_6055,N_1333,N_1049);
or U6056 (N_6056,N_2959,N_3781);
nand U6057 (N_6057,N_3836,N_2823);
nand U6058 (N_6058,N_2957,N_114);
nand U6059 (N_6059,N_4059,N_3517);
xnor U6060 (N_6060,N_3242,N_3653);
nand U6061 (N_6061,N_2675,N_764);
nor U6062 (N_6062,N_2773,N_4684);
and U6063 (N_6063,N_799,N_4922);
or U6064 (N_6064,N_2822,N_3630);
or U6065 (N_6065,N_1673,N_1989);
and U6066 (N_6066,N_3214,N_1244);
nand U6067 (N_6067,N_1321,N_218);
or U6068 (N_6068,N_2892,N_4707);
xor U6069 (N_6069,N_1897,N_1141);
nor U6070 (N_6070,N_2314,N_3727);
and U6071 (N_6071,N_2986,N_503);
xor U6072 (N_6072,N_3759,N_1168);
nand U6073 (N_6073,N_4476,N_888);
nand U6074 (N_6074,N_2358,N_3405);
nor U6075 (N_6075,N_519,N_1488);
and U6076 (N_6076,N_189,N_2160);
nor U6077 (N_6077,N_1297,N_2798);
nor U6078 (N_6078,N_833,N_4021);
nor U6079 (N_6079,N_1258,N_1709);
xnor U6080 (N_6080,N_2529,N_1730);
and U6081 (N_6081,N_3273,N_2655);
or U6082 (N_6082,N_532,N_838);
nand U6083 (N_6083,N_496,N_1737);
or U6084 (N_6084,N_608,N_4092);
and U6085 (N_6085,N_35,N_3910);
or U6086 (N_6086,N_1997,N_3375);
nand U6087 (N_6087,N_4629,N_4063);
or U6088 (N_6088,N_3635,N_4250);
nand U6089 (N_6089,N_478,N_506);
or U6090 (N_6090,N_546,N_4737);
xnor U6091 (N_6091,N_1493,N_3994);
xnor U6092 (N_6092,N_939,N_957);
nor U6093 (N_6093,N_4722,N_4602);
and U6094 (N_6094,N_1731,N_1759);
xnor U6095 (N_6095,N_1803,N_4015);
xnor U6096 (N_6096,N_425,N_4342);
nor U6097 (N_6097,N_46,N_2914);
and U6098 (N_6098,N_1068,N_4884);
or U6099 (N_6099,N_2579,N_580);
and U6100 (N_6100,N_4949,N_3154);
or U6101 (N_6101,N_1015,N_3640);
nand U6102 (N_6102,N_736,N_116);
and U6103 (N_6103,N_2308,N_3091);
nand U6104 (N_6104,N_1382,N_1747);
nor U6105 (N_6105,N_2628,N_2369);
nor U6106 (N_6106,N_3158,N_3340);
nor U6107 (N_6107,N_840,N_1698);
and U6108 (N_6108,N_4861,N_61);
nand U6109 (N_6109,N_4880,N_1441);
or U6110 (N_6110,N_3336,N_3767);
or U6111 (N_6111,N_2817,N_4796);
and U6112 (N_6112,N_3344,N_282);
xor U6113 (N_6113,N_2877,N_4596);
nor U6114 (N_6114,N_658,N_1270);
xnor U6115 (N_6115,N_2932,N_4894);
nand U6116 (N_6116,N_1595,N_1306);
nand U6117 (N_6117,N_3332,N_2553);
or U6118 (N_6118,N_3929,N_2924);
and U6119 (N_6119,N_2980,N_3714);
xnor U6120 (N_6120,N_1570,N_3397);
nand U6121 (N_6121,N_1170,N_3596);
xnor U6122 (N_6122,N_876,N_4418);
or U6123 (N_6123,N_1136,N_1817);
or U6124 (N_6124,N_2460,N_2320);
nor U6125 (N_6125,N_2847,N_4383);
or U6126 (N_6126,N_4098,N_2051);
and U6127 (N_6127,N_789,N_4371);
and U6128 (N_6128,N_1429,N_4701);
nor U6129 (N_6129,N_3801,N_2192);
xor U6130 (N_6130,N_4404,N_703);
or U6131 (N_6131,N_2152,N_4769);
nand U6132 (N_6132,N_1904,N_4664);
nor U6133 (N_6133,N_2843,N_1447);
xor U6134 (N_6134,N_1310,N_3894);
nand U6135 (N_6135,N_4833,N_2204);
and U6136 (N_6136,N_3269,N_3207);
or U6137 (N_6137,N_136,N_3946);
nand U6138 (N_6138,N_264,N_867);
nor U6139 (N_6139,N_3724,N_3300);
xor U6140 (N_6140,N_267,N_1958);
nand U6141 (N_6141,N_1305,N_3220);
xor U6142 (N_6142,N_3036,N_987);
nor U6143 (N_6143,N_4416,N_2560);
nand U6144 (N_6144,N_3942,N_372);
and U6145 (N_6145,N_1923,N_2226);
nand U6146 (N_6146,N_2944,N_2509);
nor U6147 (N_6147,N_56,N_4600);
nand U6148 (N_6148,N_2092,N_4607);
and U6149 (N_6149,N_1972,N_1379);
nand U6150 (N_6150,N_3770,N_1024);
or U6151 (N_6151,N_3679,N_538);
or U6152 (N_6152,N_3982,N_2973);
xor U6153 (N_6153,N_3044,N_1138);
xor U6154 (N_6154,N_2078,N_1461);
or U6155 (N_6155,N_4795,N_2937);
and U6156 (N_6156,N_3637,N_3223);
or U6157 (N_6157,N_2473,N_1146);
or U6158 (N_6158,N_2336,N_2669);
or U6159 (N_6159,N_1584,N_3736);
nor U6160 (N_6160,N_1365,N_2650);
and U6161 (N_6161,N_2907,N_213);
nor U6162 (N_6162,N_1961,N_3478);
nand U6163 (N_6163,N_684,N_2604);
nand U6164 (N_6164,N_3959,N_594);
xor U6165 (N_6165,N_4807,N_391);
and U6166 (N_6166,N_4754,N_1944);
and U6167 (N_6167,N_2635,N_2085);
nand U6168 (N_6168,N_1144,N_4151);
xor U6169 (N_6169,N_4246,N_556);
nor U6170 (N_6170,N_1028,N_4012);
or U6171 (N_6171,N_3662,N_2417);
and U6172 (N_6172,N_68,N_2870);
xnor U6173 (N_6173,N_2633,N_4005);
and U6174 (N_6174,N_3608,N_3531);
nor U6175 (N_6175,N_2076,N_2176);
and U6176 (N_6176,N_2510,N_1234);
nand U6177 (N_6177,N_935,N_2838);
nor U6178 (N_6178,N_2474,N_3554);
nand U6179 (N_6179,N_1317,N_3482);
nor U6180 (N_6180,N_2984,N_2827);
nand U6181 (N_6181,N_1126,N_4988);
nor U6182 (N_6182,N_3233,N_964);
or U6183 (N_6183,N_74,N_2850);
and U6184 (N_6184,N_2353,N_4489);
xnor U6185 (N_6185,N_1812,N_4710);
nand U6186 (N_6186,N_4924,N_2272);
nand U6187 (N_6187,N_1348,N_3986);
nor U6188 (N_6188,N_359,N_98);
nand U6189 (N_6189,N_3093,N_3);
xnor U6190 (N_6190,N_4097,N_2037);
or U6191 (N_6191,N_1151,N_2462);
nor U6192 (N_6192,N_4933,N_3683);
xor U6193 (N_6193,N_4494,N_2742);
or U6194 (N_6194,N_2605,N_2535);
and U6195 (N_6195,N_647,N_4991);
or U6196 (N_6196,N_4208,N_1554);
and U6197 (N_6197,N_3502,N_2751);
and U6198 (N_6198,N_95,N_4207);
and U6199 (N_6199,N_3641,N_673);
nor U6200 (N_6200,N_2539,N_949);
xor U6201 (N_6201,N_1892,N_2168);
nor U6202 (N_6202,N_3536,N_2154);
nor U6203 (N_6203,N_3949,N_4001);
nand U6204 (N_6204,N_1546,N_1893);
and U6205 (N_6205,N_286,N_757);
and U6206 (N_6206,N_4835,N_3123);
nand U6207 (N_6207,N_3547,N_2162);
nand U6208 (N_6208,N_2171,N_1103);
or U6209 (N_6209,N_2825,N_2736);
and U6210 (N_6210,N_2032,N_4630);
nand U6211 (N_6211,N_3766,N_249);
nand U6212 (N_6212,N_4804,N_3473);
and U6213 (N_6213,N_2077,N_3030);
nor U6214 (N_6214,N_3546,N_3381);
or U6215 (N_6215,N_99,N_3270);
or U6216 (N_6216,N_2015,N_1096);
or U6217 (N_6217,N_2860,N_1873);
xor U6218 (N_6218,N_3802,N_2858);
and U6219 (N_6219,N_2480,N_4641);
nor U6220 (N_6220,N_3650,N_4138);
nand U6221 (N_6221,N_976,N_1907);
nand U6222 (N_6222,N_4324,N_3931);
nand U6223 (N_6223,N_1006,N_1926);
or U6224 (N_6224,N_1063,N_3309);
nand U6225 (N_6225,N_386,N_4264);
nand U6226 (N_6226,N_3926,N_481);
or U6227 (N_6227,N_2747,N_1075);
xor U6228 (N_6228,N_4590,N_4536);
and U6229 (N_6229,N_2807,N_4364);
xnor U6230 (N_6230,N_969,N_2421);
or U6231 (N_6231,N_3612,N_654);
xnor U6232 (N_6232,N_1293,N_3930);
xor U6233 (N_6233,N_192,N_1074);
xor U6234 (N_6234,N_1195,N_3192);
or U6235 (N_6235,N_4405,N_2270);
and U6236 (N_6236,N_755,N_1950);
nand U6237 (N_6237,N_1088,N_2282);
and U6238 (N_6238,N_235,N_3606);
and U6239 (N_6239,N_180,N_38);
nor U6240 (N_6240,N_530,N_959);
or U6241 (N_6241,N_15,N_2867);
or U6242 (N_6242,N_4709,N_3668);
nand U6243 (N_6243,N_4118,N_4662);
and U6244 (N_6244,N_3523,N_1618);
xnor U6245 (N_6245,N_3580,N_4646);
and U6246 (N_6246,N_750,N_314);
xor U6247 (N_6247,N_3284,N_138);
xnor U6248 (N_6248,N_825,N_2450);
xor U6249 (N_6249,N_904,N_4115);
nand U6250 (N_6250,N_1169,N_4863);
or U6251 (N_6251,N_2399,N_2329);
nand U6252 (N_6252,N_4803,N_2659);
or U6253 (N_6253,N_1981,N_1351);
xnor U6254 (N_6254,N_960,N_4671);
nand U6255 (N_6255,N_1106,N_2443);
nand U6256 (N_6256,N_4622,N_4298);
xor U6257 (N_6257,N_1549,N_4591);
xnor U6258 (N_6258,N_2118,N_4307);
and U6259 (N_6259,N_3782,N_3425);
and U6260 (N_6260,N_2886,N_178);
nor U6261 (N_6261,N_3525,N_4966);
nand U6262 (N_6262,N_4716,N_4300);
and U6263 (N_6263,N_1256,N_4587);
or U6264 (N_6264,N_2235,N_533);
nand U6265 (N_6265,N_2580,N_3576);
and U6266 (N_6266,N_4028,N_3379);
nand U6267 (N_6267,N_801,N_3561);
or U6268 (N_6268,N_394,N_446);
or U6269 (N_6269,N_1471,N_4159);
nand U6270 (N_6270,N_2386,N_63);
and U6271 (N_6271,N_1344,N_1468);
or U6272 (N_6272,N_2079,N_405);
nand U6273 (N_6273,N_1996,N_1928);
xnor U6274 (N_6274,N_4375,N_3594);
and U6275 (N_6275,N_1510,N_1279);
xor U6276 (N_6276,N_59,N_4206);
nand U6277 (N_6277,N_860,N_2109);
and U6278 (N_6278,N_3718,N_4060);
xor U6279 (N_6279,N_3304,N_3543);
nand U6280 (N_6280,N_3421,N_1593);
and U6281 (N_6281,N_1391,N_3941);
or U6282 (N_6282,N_1728,N_516);
xor U6283 (N_6283,N_751,N_4613);
nor U6284 (N_6284,N_2439,N_3373);
and U6285 (N_6285,N_4983,N_641);
or U6286 (N_6286,N_3338,N_2331);
xnor U6287 (N_6287,N_4530,N_365);
and U6288 (N_6288,N_3476,N_1992);
and U6289 (N_6289,N_3282,N_2046);
nand U6290 (N_6290,N_3533,N_3132);
xor U6291 (N_6291,N_3851,N_4212);
nand U6292 (N_6292,N_1568,N_2517);
and U6293 (N_6293,N_1,N_4770);
or U6294 (N_6294,N_955,N_1919);
and U6295 (N_6295,N_4120,N_199);
nand U6296 (N_6296,N_572,N_3795);
xnor U6297 (N_6297,N_2698,N_3422);
xnor U6298 (N_6298,N_3557,N_4209);
or U6299 (N_6299,N_1320,N_1741);
or U6300 (N_6300,N_2526,N_3932);
or U6301 (N_6301,N_3565,N_4480);
nor U6302 (N_6302,N_3639,N_4713);
nor U6303 (N_6303,N_4142,N_3588);
xor U6304 (N_6304,N_857,N_1760);
nand U6305 (N_6305,N_943,N_1301);
and U6306 (N_6306,N_4330,N_2643);
and U6307 (N_6307,N_3308,N_2280);
nor U6308 (N_6308,N_4919,N_4882);
xnor U6309 (N_6309,N_2437,N_148);
or U6310 (N_6310,N_2195,N_4532);
xor U6311 (N_6311,N_1567,N_2657);
and U6312 (N_6312,N_2230,N_3048);
nor U6313 (N_6313,N_2626,N_3240);
nor U6314 (N_6314,N_2874,N_1140);
or U6315 (N_6315,N_2848,N_829);
or U6316 (N_6316,N_1131,N_4216);
nand U6317 (N_6317,N_4856,N_3749);
nand U6318 (N_6318,N_1573,N_231);
or U6319 (N_6319,N_4359,N_3704);
nor U6320 (N_6320,N_837,N_393);
nor U6321 (N_6321,N_3883,N_2700);
nor U6322 (N_6322,N_4009,N_2997);
xor U6323 (N_6323,N_3682,N_3342);
xor U6324 (N_6324,N_3758,N_2878);
and U6325 (N_6325,N_1119,N_3581);
nor U6326 (N_6326,N_931,N_4980);
nand U6327 (N_6327,N_4389,N_2965);
nor U6328 (N_6328,N_3205,N_4886);
nand U6329 (N_6329,N_1375,N_1895);
nand U6330 (N_6330,N_4424,N_3073);
or U6331 (N_6331,N_2908,N_2779);
nand U6332 (N_6332,N_631,N_4793);
and U6333 (N_6333,N_358,N_266);
and U6334 (N_6334,N_2964,N_442);
or U6335 (N_6335,N_1896,N_1689);
and U6336 (N_6336,N_2301,N_1328);
and U6337 (N_6337,N_4340,N_269);
and U6338 (N_6338,N_3981,N_938);
nand U6339 (N_6339,N_4780,N_3264);
or U6340 (N_6340,N_374,N_1426);
nand U6341 (N_6341,N_2976,N_2170);
xor U6342 (N_6342,N_3465,N_4454);
or U6343 (N_6343,N_2021,N_4003);
xor U6344 (N_6344,N_1467,N_2112);
nor U6345 (N_6345,N_1021,N_3017);
nand U6346 (N_6346,N_640,N_3887);
and U6347 (N_6347,N_3889,N_2837);
xor U6348 (N_6348,N_633,N_1152);
xnor U6349 (N_6349,N_272,N_1053);
nand U6350 (N_6350,N_2248,N_2278);
and U6351 (N_6351,N_4733,N_2538);
nor U6352 (N_6352,N_2716,N_1302);
or U6353 (N_6353,N_879,N_2380);
and U6354 (N_6354,N_2464,N_2568);
and U6355 (N_6355,N_739,N_127);
or U6356 (N_6356,N_2453,N_1001);
nor U6357 (N_6357,N_738,N_1791);
or U6358 (N_6358,N_806,N_389);
xor U6359 (N_6359,N_1677,N_1909);
xnor U6360 (N_6360,N_1776,N_4470);
nor U6361 (N_6361,N_2059,N_4313);
nand U6362 (N_6362,N_4398,N_3882);
nand U6363 (N_6363,N_426,N_4172);
nor U6364 (N_6364,N_573,N_983);
or U6365 (N_6365,N_2035,N_3275);
nor U6366 (N_6366,N_1660,N_170);
xnor U6367 (N_6367,N_1295,N_683);
xnor U6368 (N_6368,N_3153,N_1066);
xnor U6369 (N_6369,N_248,N_3761);
or U6370 (N_6370,N_1336,N_3062);
nor U6371 (N_6371,N_699,N_1353);
nand U6372 (N_6372,N_4179,N_4753);
or U6373 (N_6373,N_4844,N_1548);
nor U6374 (N_6374,N_1163,N_4378);
and U6375 (N_6375,N_4853,N_4708);
xor U6376 (N_6376,N_3762,N_3325);
xnor U6377 (N_6377,N_667,N_186);
xor U6378 (N_6378,N_2207,N_3164);
nor U6379 (N_6379,N_2776,N_1416);
nor U6380 (N_6380,N_3847,N_1982);
xnor U6381 (N_6381,N_3799,N_878);
nand U6382 (N_6382,N_2661,N_4952);
nor U6383 (N_6383,N_2912,N_2244);
or U6384 (N_6384,N_1114,N_4279);
nor U6385 (N_6385,N_2311,N_3921);
xnor U6386 (N_6386,N_1402,N_3043);
and U6387 (N_6387,N_4921,N_3000);
or U6388 (N_6388,N_328,N_3884);
and U6389 (N_6389,N_3259,N_3712);
and U6390 (N_6390,N_3809,N_132);
or U6391 (N_6391,N_1417,N_216);
nor U6392 (N_6392,N_2653,N_172);
nor U6393 (N_6393,N_2987,N_4275);
nand U6394 (N_6394,N_986,N_569);
and U6395 (N_6395,N_3306,N_1184);
nand U6396 (N_6396,N_2668,N_3228);
nand U6397 (N_6397,N_3353,N_0);
xnor U6398 (N_6398,N_2061,N_1230);
nor U6399 (N_6399,N_2702,N_3292);
nand U6400 (N_6400,N_720,N_2066);
nand U6401 (N_6401,N_3723,N_2699);
and U6402 (N_6402,N_2542,N_544);
xnor U6403 (N_6403,N_3503,N_1263);
nor U6404 (N_6404,N_2312,N_1516);
xnor U6405 (N_6405,N_1881,N_2791);
nand U6406 (N_6406,N_977,N_1675);
and U6407 (N_6407,N_2713,N_31);
nand U6408 (N_6408,N_3213,N_3305);
xor U6409 (N_6409,N_1445,N_55);
and U6410 (N_6410,N_4925,N_557);
xor U6411 (N_6411,N_4881,N_4017);
or U6412 (N_6412,N_313,N_4632);
xnor U6413 (N_6413,N_1371,N_333);
xnor U6414 (N_6414,N_1611,N_4384);
nor U6415 (N_6415,N_4107,N_81);
xnor U6416 (N_6416,N_3250,N_1360);
and U6417 (N_6417,N_3648,N_567);
nor U6418 (N_6418,N_2496,N_3436);
xor U6419 (N_6419,N_2151,N_2710);
and U6420 (N_6420,N_3507,N_3488);
or U6421 (N_6421,N_933,N_1329);
nand U6422 (N_6422,N_2896,N_1073);
xor U6423 (N_6423,N_3006,N_3160);
nand U6424 (N_6424,N_4969,N_1022);
or U6425 (N_6425,N_1067,N_3156);
nor U6426 (N_6426,N_311,N_3976);
nor U6427 (N_6427,N_4436,N_195);
or U6428 (N_6428,N_4407,N_1861);
and U6429 (N_6429,N_4956,N_3265);
and U6430 (N_6430,N_3234,N_187);
or U6431 (N_6431,N_1596,N_1377);
nor U6432 (N_6432,N_3427,N_1080);
and U6433 (N_6433,N_4703,N_3165);
nand U6434 (N_6434,N_3741,N_2969);
or U6435 (N_6435,N_1902,N_4503);
or U6436 (N_6436,N_1682,N_1250);
xor U6437 (N_6437,N_3103,N_4064);
or U6438 (N_6438,N_439,N_3076);
nor U6439 (N_6439,N_432,N_2682);
xor U6440 (N_6440,N_3756,N_2622);
nor U6441 (N_6441,N_940,N_4238);
xnor U6442 (N_6442,N_4234,N_4704);
xnor U6443 (N_6443,N_1993,N_4889);
or U6444 (N_6444,N_3483,N_4287);
nand U6445 (N_6445,N_72,N_2871);
nor U6446 (N_6446,N_1828,N_2949);
or U6447 (N_6447,N_2884,N_4388);
and U6448 (N_6448,N_1786,N_3296);
nand U6449 (N_6449,N_1705,N_3485);
or U6450 (N_6450,N_3403,N_1060);
nand U6451 (N_6451,N_2318,N_3587);
nor U6452 (N_6452,N_2951,N_4166);
or U6453 (N_6453,N_4449,N_1261);
and U6454 (N_6454,N_4777,N_3484);
and U6455 (N_6455,N_43,N_4154);
xor U6456 (N_6456,N_2557,N_1715);
xnor U6457 (N_6457,N_4904,N_489);
nand U6458 (N_6458,N_3558,N_2583);
nor U6459 (N_6459,N_2756,N_1276);
xnor U6460 (N_6460,N_3026,N_1478);
or U6461 (N_6461,N_3470,N_4349);
nor U6462 (N_6462,N_3172,N_2824);
nand U6463 (N_6463,N_4767,N_1733);
or U6464 (N_6464,N_848,N_4199);
or U6465 (N_6465,N_849,N_1566);
or U6466 (N_6466,N_3023,N_1503);
and U6467 (N_6467,N_853,N_349);
nand U6468 (N_6468,N_2433,N_2442);
nand U6469 (N_6469,N_609,N_4852);
nor U6470 (N_6470,N_3477,N_4989);
and U6471 (N_6471,N_1915,N_2403);
or U6472 (N_6472,N_4771,N_142);
xor U6473 (N_6473,N_4543,N_4231);
and U6474 (N_6474,N_3560,N_3391);
nand U6475 (N_6475,N_4423,N_1070);
nand U6476 (N_6476,N_2262,N_2294);
nor U6477 (N_6477,N_1134,N_3827);
nand U6478 (N_6478,N_4432,N_30);
nand U6479 (N_6479,N_3090,N_353);
nand U6480 (N_6480,N_3716,N_4044);
nand U6481 (N_6481,N_3434,N_2544);
nor U6482 (N_6482,N_3968,N_1605);
nand U6483 (N_6483,N_3491,N_4200);
xor U6484 (N_6484,N_1227,N_1490);
and U6485 (N_6485,N_636,N_475);
nand U6486 (N_6486,N_1121,N_717);
nand U6487 (N_6487,N_3671,N_4724);
nand U6488 (N_6488,N_4826,N_1013);
xnor U6489 (N_6489,N_236,N_3217);
and U6490 (N_6490,N_423,N_1345);
and U6491 (N_6491,N_4917,N_2412);
nor U6492 (N_6492,N_3225,N_1356);
nand U6493 (N_6493,N_4774,N_4357);
or U6494 (N_6494,N_941,N_4139);
nand U6495 (N_6495,N_2660,N_2198);
nand U6496 (N_6496,N_412,N_4280);
xnor U6497 (N_6497,N_2684,N_2124);
and U6498 (N_6498,N_3209,N_2449);
and U6499 (N_6499,N_1210,N_2324);
and U6500 (N_6500,N_1218,N_971);
nand U6501 (N_6501,N_2042,N_4062);
xnor U6502 (N_6502,N_1752,N_4274);
nor U6503 (N_6503,N_2084,N_4211);
xnor U6504 (N_6504,N_4522,N_2577);
or U6505 (N_6505,N_4971,N_321);
and U6506 (N_6506,N_3508,N_2422);
or U6507 (N_6507,N_1590,N_4509);
xor U6508 (N_6508,N_1089,N_3956);
and U6509 (N_6509,N_122,N_1042);
and U6510 (N_6510,N_2948,N_1653);
nor U6511 (N_6511,N_1352,N_4316);
nand U6512 (N_6512,N_1969,N_2952);
or U6513 (N_6513,N_2644,N_1998);
nand U6514 (N_6514,N_3479,N_2185);
nor U6515 (N_6515,N_196,N_1831);
nand U6516 (N_6516,N_1768,N_786);
nand U6517 (N_6517,N_335,N_4812);
nor U6518 (N_6518,N_1130,N_4196);
nand U6519 (N_6519,N_3505,N_465);
or U6520 (N_6520,N_577,N_2338);
xor U6521 (N_6521,N_681,N_1421);
xnor U6522 (N_6522,N_1167,N_3522);
or U6523 (N_6523,N_3449,N_2901);
and U6524 (N_6524,N_4498,N_844);
or U6525 (N_6525,N_665,N_599);
or U6526 (N_6526,N_1150,N_1765);
nor U6527 (N_6527,N_462,N_2975);
xnor U6528 (N_6528,N_1968,N_1991);
nor U6529 (N_6529,N_1612,N_3281);
xnor U6530 (N_6530,N_613,N_3865);
xor U6531 (N_6531,N_4444,N_1514);
nor U6532 (N_6532,N_3410,N_3334);
nor U6533 (N_6533,N_1434,N_1565);
nor U6534 (N_6534,N_1181,N_4144);
nand U6535 (N_6535,N_1065,N_3051);
and U6536 (N_6536,N_4620,N_2849);
nor U6537 (N_6537,N_558,N_211);
and U6538 (N_6538,N_914,N_2489);
xor U6539 (N_6539,N_1749,N_1544);
nand U6540 (N_6540,N_428,N_4483);
xor U6541 (N_6541,N_4799,N_2726);
xor U6542 (N_6542,N_1303,N_2502);
nor U6543 (N_6543,N_2645,N_1085);
nand U6544 (N_6544,N_2431,N_1866);
nor U6545 (N_6545,N_744,N_910);
nand U6546 (N_6546,N_3169,N_3790);
or U6547 (N_6547,N_3902,N_4419);
xnor U6548 (N_6548,N_3593,N_4175);
nor U6549 (N_6549,N_3681,N_3472);
nand U6550 (N_6550,N_3261,N_1564);
and U6551 (N_6551,N_2514,N_4680);
nor U6552 (N_6552,N_815,N_1589);
or U6553 (N_6553,N_1318,N_1736);
xnor U6554 (N_6554,N_4987,N_2821);
and U6555 (N_6555,N_4467,N_3016);
and U6556 (N_6556,N_3983,N_3860);
and U6557 (N_6557,N_1485,N_3115);
and U6558 (N_6558,N_2760,N_1912);
nand U6559 (N_6559,N_2487,N_4516);
nor U6560 (N_6560,N_584,N_4133);
and U6561 (N_6561,N_2978,N_3272);
nand U6562 (N_6562,N_748,N_2759);
xnor U6563 (N_6563,N_3395,N_3916);
or U6564 (N_6564,N_3872,N_1850);
or U6565 (N_6565,N_800,N_329);
nand U6566 (N_6566,N_401,N_3825);
xnor U6567 (N_6567,N_3082,N_2995);
nand U6568 (N_6568,N_179,N_1498);
and U6569 (N_6569,N_4485,N_4759);
nand U6570 (N_6570,N_4819,N_4125);
nand U6571 (N_6571,N_1326,N_3418);
and U6572 (N_6572,N_4069,N_4529);
or U6573 (N_6573,N_4024,N_2955);
xor U6574 (N_6574,N_469,N_937);
xor U6575 (N_6575,N_512,N_2584);
or U6576 (N_6576,N_3119,N_2267);
or U6577 (N_6577,N_4943,N_4385);
xnor U6578 (N_6578,N_2938,N_2471);
or U6579 (N_6579,N_3765,N_1750);
or U6580 (N_6580,N_626,N_2273);
and U6581 (N_6581,N_1231,N_3697);
and U6582 (N_6582,N_1097,N_1432);
or U6583 (N_6583,N_2127,N_3922);
or U6584 (N_6584,N_3064,N_3973);
and U6585 (N_6585,N_637,N_2888);
or U6586 (N_6586,N_2223,N_84);
or U6587 (N_6587,N_1341,N_319);
or U6588 (N_6588,N_1716,N_589);
xor U6589 (N_6589,N_1052,N_2285);
nor U6590 (N_6590,N_2741,N_4700);
and U6591 (N_6591,N_2286,N_436);
nand U6592 (N_6592,N_1994,N_759);
nand U6593 (N_6593,N_3167,N_913);
nor U6594 (N_6594,N_944,N_3537);
xor U6595 (N_6595,N_1541,N_2029);
nand U6596 (N_6596,N_1165,N_3601);
nand U6597 (N_6597,N_305,N_2942);
nor U6598 (N_6598,N_1419,N_1446);
and U6599 (N_6599,N_4843,N_3243);
and U6600 (N_6600,N_4303,N_3387);
xnor U6601 (N_6601,N_3966,N_2565);
and U6602 (N_6602,N_4540,N_714);
nor U6603 (N_6603,N_222,N_482);
xnor U6604 (N_6604,N_942,N_3411);
and U6605 (N_6605,N_893,N_488);
nor U6606 (N_6606,N_1685,N_2728);
or U6607 (N_6607,N_1938,N_1094);
xnor U6608 (N_6608,N_420,N_2921);
and U6609 (N_6609,N_3045,N_347);
nor U6610 (N_6610,N_1948,N_2927);
nand U6611 (N_6611,N_34,N_4755);
nand U6612 (N_6612,N_471,N_2287);
or U6613 (N_6613,N_1470,N_3360);
and U6614 (N_6614,N_4674,N_3907);
nor U6615 (N_6615,N_1586,N_3412);
nor U6616 (N_6616,N_1430,N_440);
and U6617 (N_6617,N_3113,N_1147);
nand U6618 (N_6618,N_4338,N_3382);
nand U6619 (N_6619,N_811,N_1221);
xor U6620 (N_6620,N_36,N_1497);
and U6621 (N_6621,N_3198,N_3347);
and U6622 (N_6622,N_895,N_917);
or U6623 (N_6623,N_911,N_4284);
nor U6624 (N_6624,N_320,N_366);
or U6625 (N_6625,N_807,N_3194);
nand U6626 (N_6626,N_2304,N_3832);
and U6627 (N_6627,N_2048,N_832);
nand U6628 (N_6628,N_4242,N_1888);
and U6629 (N_6629,N_270,N_4051);
or U6630 (N_6630,N_1186,N_1740);
nand U6631 (N_6631,N_2100,N_3467);
xnor U6632 (N_6632,N_3620,N_4337);
nor U6633 (N_6633,N_2144,N_3283);
nand U6634 (N_6634,N_1314,N_3945);
or U6635 (N_6635,N_4311,N_2505);
nor U6636 (N_6636,N_291,N_212);
and U6637 (N_6637,N_3721,N_1833);
and U6638 (N_6638,N_2578,N_4663);
or U6639 (N_6639,N_4649,N_963);
and U6640 (N_6640,N_760,N_4633);
and U6641 (N_6641,N_3513,N_4967);
xnor U6642 (N_6642,N_2694,N_303);
xor U6643 (N_6643,N_2292,N_2036);
nor U6644 (N_6644,N_3174,N_2381);
nand U6645 (N_6645,N_732,N_2666);
and U6646 (N_6646,N_2423,N_1574);
or U6647 (N_6647,N_1847,N_1137);
xor U6648 (N_6648,N_4109,N_3954);
or U6649 (N_6649,N_2003,N_4463);
or U6650 (N_6650,N_4908,N_2491);
nand U6651 (N_6651,N_1863,N_2392);
nor U6652 (N_6652,N_4180,N_3886);
or U6653 (N_6653,N_529,N_4451);
and U6654 (N_6654,N_3099,N_2750);
nand U6655 (N_6655,N_746,N_3326);
nor U6656 (N_6656,N_1286,N_2288);
nor U6657 (N_6657,N_2895,N_3227);
xor U6658 (N_6658,N_678,N_4535);
nand U6659 (N_6659,N_302,N_1205);
nand U6660 (N_6660,N_1729,N_4479);
and U6661 (N_6661,N_1440,N_3404);
or U6662 (N_6662,N_2971,N_817);
nor U6663 (N_6663,N_898,N_827);
or U6664 (N_6664,N_1597,N_1946);
nand U6665 (N_6665,N_2930,N_3830);
nand U6666 (N_6666,N_1190,N_947);
xor U6667 (N_6667,N_1878,N_4763);
nand U6668 (N_6668,N_908,N_4395);
and U6669 (N_6669,N_3516,N_624);
xnor U6670 (N_6670,N_3544,N_1036);
nand U6671 (N_6671,N_3626,N_1223);
nor U6672 (N_6672,N_4178,N_4815);
nand U6673 (N_6673,N_3226,N_3316);
nand U6674 (N_6674,N_2342,N_164);
or U6675 (N_6675,N_118,N_2113);
xnor U6676 (N_6676,N_2146,N_2141);
nand U6677 (N_6677,N_2355,N_4429);
nor U6678 (N_6678,N_134,N_3647);
xor U6679 (N_6679,N_1925,N_1481);
and U6680 (N_6680,N_4789,N_4136);
nand U6681 (N_6681,N_3928,N_2345);
and U6682 (N_6682,N_4583,N_1264);
or U6683 (N_6683,N_215,N_1953);
or U6684 (N_6684,N_1443,N_3645);
nand U6685 (N_6685,N_6,N_2179);
nand U6686 (N_6686,N_4071,N_1451);
nor U6687 (N_6687,N_3141,N_3891);
or U6688 (N_6688,N_3432,N_1971);
nand U6689 (N_6689,N_2231,N_3289);
xnor U6690 (N_6690,N_4790,N_1459);
nor U6691 (N_6691,N_2274,N_2780);
nand U6692 (N_6692,N_4521,N_50);
and U6693 (N_6693,N_2402,N_992);
and U6694 (N_6694,N_2602,N_2582);
xor U6695 (N_6695,N_4047,N_1806);
nand U6696 (N_6696,N_3846,N_687);
nand U6697 (N_6697,N_3852,N_495);
xnor U6698 (N_6698,N_3203,N_1528);
nand U6699 (N_6699,N_32,N_3059);
or U6700 (N_6700,N_1155,N_2648);
xnor U6701 (N_6701,N_4190,N_2265);
or U6702 (N_6702,N_4542,N_3277);
and U6703 (N_6703,N_615,N_4473);
nor U6704 (N_6704,N_2738,N_1809);
and U6705 (N_6705,N_2307,N_4445);
nor U6706 (N_6706,N_3854,N_3196);
nor U6707 (N_6707,N_2596,N_819);
xnor U6708 (N_6708,N_1976,N_258);
and U6709 (N_6709,N_1785,N_4714);
or U6710 (N_6710,N_3406,N_868);
and U6711 (N_6711,N_873,N_2377);
nand U6712 (N_6712,N_4849,N_3939);
nor U6713 (N_6713,N_1606,N_1162);
xnor U6714 (N_6714,N_2440,N_4627);
and U6715 (N_6715,N_2788,N_3500);
nor U6716 (N_6716,N_3694,N_1269);
xor U6717 (N_6717,N_3224,N_1282);
and U6718 (N_6718,N_993,N_3061);
nor U6719 (N_6719,N_3067,N_4652);
and U6720 (N_6720,N_3046,N_4446);
nand U6721 (N_6721,N_2500,N_3610);
nand U6722 (N_6722,N_397,N_2840);
and U6723 (N_6723,N_2220,N_3110);
or U6724 (N_6724,N_4131,N_781);
nand U6725 (N_6725,N_1178,N_4156);
xnor U6726 (N_6726,N_1175,N_4294);
nand U6727 (N_6727,N_119,N_4184);
xnor U6728 (N_6728,N_47,N_4560);
xnor U6729 (N_6729,N_2143,N_4177);
xnor U6730 (N_6730,N_2221,N_3301);
or U6731 (N_6731,N_2761,N_1019);
nand U6732 (N_6732,N_3159,N_171);
nor U6733 (N_6733,N_1901,N_4610);
nand U6734 (N_6734,N_816,N_2672);
or U6735 (N_6735,N_3004,N_1422);
nor U6736 (N_6736,N_1661,N_1225);
nand U6737 (N_6737,N_452,N_2928);
xnor U6738 (N_6738,N_3148,N_1288);
nand U6739 (N_6739,N_4126,N_3738);
or U6740 (N_6740,N_1133,N_27);
nand U6741 (N_6741,N_2157,N_1271);
or U6742 (N_6742,N_2873,N_4290);
nand U6743 (N_6743,N_777,N_487);
xor U6744 (N_6744,N_2591,N_2451);
and U6745 (N_6745,N_1815,N_3744);
xor U6746 (N_6746,N_2970,N_1215);
nand U6747 (N_6747,N_1405,N_3734);
and U6748 (N_6748,N_981,N_688);
nand U6749 (N_6749,N_3623,N_3083);
nand U6750 (N_6750,N_3855,N_2730);
xnor U6751 (N_6751,N_2861,N_4067);
and U6752 (N_6752,N_783,N_1869);
or U6753 (N_6753,N_4262,N_2275);
and U6754 (N_6754,N_4043,N_600);
nand U6755 (N_6755,N_3869,N_4740);
or U6756 (N_6756,N_828,N_457);
nand U6757 (N_6757,N_3420,N_4210);
nand U6758 (N_6758,N_4841,N_1774);
nand U6759 (N_6759,N_1858,N_3739);
xor U6760 (N_6760,N_1551,N_2749);
and U6761 (N_6761,N_3582,N_4698);
xnor U6762 (N_6762,N_4121,N_4653);
nand U6763 (N_6763,N_280,N_1346);
and U6764 (N_6764,N_4134,N_3675);
or U6765 (N_6765,N_4014,N_4160);
and U6766 (N_6766,N_1695,N_4502);
or U6767 (N_6767,N_1853,N_4360);
and U6768 (N_6768,N_1242,N_4462);
xor U6769 (N_6769,N_4046,N_1917);
nor U6770 (N_6770,N_2013,N_1330);
or U6771 (N_6771,N_4495,N_3833);
and U6772 (N_6772,N_1744,N_2717);
nand U6773 (N_6773,N_2631,N_2897);
nand U6774 (N_6774,N_3235,N_2352);
nor U6775 (N_6775,N_2609,N_826);
and U6776 (N_6776,N_4507,N_3621);
or U6777 (N_6777,N_1647,N_4730);
nand U6778 (N_6778,N_4117,N_1436);
xor U6779 (N_6779,N_1580,N_1177);
or U6780 (N_6780,N_3909,N_4408);
and U6781 (N_6781,N_1204,N_3029);
and U6782 (N_6782,N_2357,N_2820);
xnor U6783 (N_6783,N_1975,N_4547);
nor U6784 (N_6784,N_2658,N_3520);
nand U6785 (N_6785,N_2252,N_1646);
nand U6786 (N_6786,N_4809,N_3071);
or U6787 (N_6787,N_2943,N_1883);
or U6788 (N_6788,N_3804,N_217);
and U6789 (N_6789,N_3307,N_774);
or U6790 (N_6790,N_2309,N_2846);
nand U6791 (N_6791,N_1499,N_1268);
and U6792 (N_6792,N_841,N_3908);
nor U6793 (N_6793,N_3032,N_1120);
or U6794 (N_6794,N_4343,N_3348);
nor U6795 (N_6795,N_2587,N_2512);
or U6796 (N_6796,N_1476,N_1062);
nor U6797 (N_6797,N_1927,N_4588);
or U6798 (N_6798,N_1632,N_2466);
nand U6799 (N_6799,N_1965,N_1738);
xor U6800 (N_6800,N_3365,N_3060);
nand U6801 (N_6801,N_686,N_1876);
nand U6802 (N_6802,N_4897,N_289);
and U6803 (N_6803,N_3438,N_1794);
or U6804 (N_6804,N_2234,N_169);
nand U6805 (N_6805,N_3134,N_2388);
nand U6806 (N_6806,N_4867,N_3331);
and U6807 (N_6807,N_805,N_894);
nand U6808 (N_6808,N_4555,N_263);
and U6809 (N_6809,N_4101,N_2787);
and U6810 (N_6810,N_3937,N_1222);
and U6811 (N_6811,N_3138,N_2247);
nor U6812 (N_6812,N_767,N_2933);
and U6813 (N_6813,N_2300,N_2340);
xnor U6814 (N_6814,N_4482,N_4621);
and U6815 (N_6815,N_4326,N_2624);
or U6816 (N_6816,N_1827,N_2679);
nor U6817 (N_6817,N_3133,N_2297);
and U6818 (N_6818,N_3069,N_655);
xor U6819 (N_6819,N_4111,N_2039);
xnor U6820 (N_6820,N_2866,N_1521);
nand U6821 (N_6821,N_3905,N_1399);
and U6822 (N_6822,N_3318,N_1908);
nor U6823 (N_6823,N_2996,N_4041);
nand U6824 (N_6824,N_3607,N_166);
nand U6825 (N_6825,N_2946,N_707);
and U6826 (N_6826,N_4773,N_3823);
xor U6827 (N_6827,N_4425,N_4434);
xor U6828 (N_6828,N_4781,N_1335);
nor U6829 (N_6829,N_1464,N_229);
and U6830 (N_6830,N_4094,N_3563);
or U6831 (N_6831,N_3936,N_1626);
nand U6832 (N_6832,N_3462,N_2869);
and U6833 (N_6833,N_2724,N_1095);
or U6834 (N_6834,N_4174,N_866);
nand U6835 (N_6835,N_542,N_3632);
or U6836 (N_6836,N_284,N_3550);
nand U6837 (N_6837,N_2150,N_336);
or U6838 (N_6838,N_2667,N_616);
and U6839 (N_6839,N_470,N_3977);
xnor U6840 (N_6840,N_1359,N_5);
and U6841 (N_6841,N_4858,N_769);
xnor U6842 (N_6842,N_2295,N_3733);
nor U6843 (N_6843,N_1639,N_3005);
nand U6844 (N_6844,N_3879,N_3390);
nand U6845 (N_6845,N_2790,N_4037);
nor U6846 (N_6846,N_449,N_4931);
or U6847 (N_6847,N_2525,N_1891);
nor U6848 (N_6848,N_4690,N_3709);
xor U6849 (N_6849,N_4008,N_125);
nor U6850 (N_6850,N_2729,N_64);
or U6851 (N_6851,N_484,N_220);
xnor U6852 (N_6852,N_3429,N_2082);
nor U6853 (N_6853,N_392,N_4119);
nor U6854 (N_6854,N_3798,N_1822);
nor U6855 (N_6855,N_2649,N_4792);
xor U6856 (N_6856,N_4320,N_2106);
or U6857 (N_6857,N_4465,N_4592);
nor U6858 (N_6858,N_4531,N_2245);
xor U6859 (N_6859,N_3527,N_1251);
or U6860 (N_6860,N_3893,N_2409);
xor U6861 (N_6861,N_1702,N_3319);
and U6862 (N_6862,N_3567,N_4992);
and U6863 (N_6863,N_44,N_4082);
xor U6864 (N_6864,N_4788,N_238);
or U6865 (N_6865,N_4490,N_120);
and U6866 (N_6866,N_1631,N_1823);
nand U6867 (N_6867,N_2454,N_42);
nand U6868 (N_6868,N_4427,N_4717);
or U6869 (N_6869,N_4116,N_2974);
nor U6870 (N_6870,N_2576,N_3615);
xnor U6871 (N_6871,N_4675,N_4191);
or U6872 (N_6872,N_4475,N_2333);
nor U6873 (N_6873,N_1782,N_661);
nor U6874 (N_6874,N_4875,N_2941);
nand U6875 (N_6875,N_4811,N_2131);
nand U6876 (N_6876,N_143,N_3450);
xor U6877 (N_6877,N_60,N_4823);
or U6878 (N_6878,N_3211,N_2323);
nor U6879 (N_6879,N_3690,N_2549);
nor U6880 (N_6880,N_706,N_497);
xor U6881 (N_6881,N_861,N_1887);
or U6882 (N_6882,N_4559,N_4285);
xnor U6883 (N_6883,N_3322,N_1659);
and U6884 (N_6884,N_145,N_2461);
nor U6885 (N_6885,N_3747,N_2872);
xnor U6886 (N_6886,N_1951,N_1784);
xor U6887 (N_6887,N_4929,N_1557);
nand U6888 (N_6888,N_4661,N_276);
xor U6889 (N_6889,N_2009,N_337);
xnor U6890 (N_6890,N_158,N_754);
nand U6891 (N_6891,N_4619,N_4466);
xnor U6892 (N_6892,N_4827,N_93);
and U6893 (N_6893,N_1009,N_407);
xnor U6894 (N_6894,N_3355,N_522);
nor U6895 (N_6895,N_3702,N_4864);
or U6896 (N_6896,N_4106,N_3871);
xnor U6897 (N_6897,N_3239,N_1428);
xnor U6898 (N_6898,N_2696,N_3625);
and U6899 (N_6899,N_4321,N_4148);
and U6900 (N_6900,N_3863,N_668);
and U6901 (N_6901,N_2398,N_2673);
nor U6902 (N_6902,N_1523,N_4455);
nand U6903 (N_6903,N_2826,N_4080);
xor U6904 (N_6904,N_4201,N_954);
or U6905 (N_6905,N_1041,N_2041);
xor U6906 (N_6906,N_2586,N_4741);
and U6907 (N_6907,N_1307,N_798);
nand U6908 (N_6908,N_1666,N_1960);
xnor U6909 (N_6909,N_3084,N_2132);
nand U6910 (N_6910,N_2835,N_350);
nand U6911 (N_6911,N_1453,N_1645);
nor U6912 (N_6912,N_2360,N_1739);
nand U6913 (N_6913,N_930,N_4517);
nor U6914 (N_6914,N_3256,N_2831);
nand U6915 (N_6915,N_3696,N_3779);
xnor U6916 (N_6916,N_4998,N_2428);
or U6917 (N_6917,N_1449,N_3202);
and U6918 (N_6918,N_4085,N_4999);
nand U6919 (N_6919,N_3705,N_3813);
nor U6920 (N_6920,N_242,N_1054);
and U6921 (N_6921,N_1692,N_3253);
or U6922 (N_6922,N_2769,N_3559);
nor U6923 (N_6923,N_3297,N_364);
xor U6924 (N_6924,N_3816,N_4883);
or U6925 (N_6925,N_3829,N_2296);
nand U6926 (N_6926,N_734,N_1495);
xor U6927 (N_6927,N_1845,N_4665);
or U6928 (N_6928,N_2122,N_1007);
nand U6929 (N_6929,N_606,N_403);
nand U6930 (N_6930,N_268,N_3419);
and U6931 (N_6931,N_285,N_4353);
xnor U6932 (N_6932,N_1843,N_2498);
nand U6933 (N_6933,N_4995,N_4660);
nor U6934 (N_6934,N_253,N_2123);
or U6935 (N_6935,N_4728,N_354);
nand U6936 (N_6936,N_4409,N_1875);
nor U6937 (N_6937,N_2062,N_3673);
and U6938 (N_6938,N_4820,N_3378);
and U6939 (N_6939,N_2347,N_882);
xnor U6940 (N_6940,N_4589,N_2687);
nand U6941 (N_6941,N_3578,N_3591);
and U6942 (N_6942,N_1182,N_2216);
nor U6943 (N_6943,N_131,N_834);
nand U6944 (N_6944,N_3938,N_4390);
nor U6945 (N_6945,N_1394,N_66);
xor U6946 (N_6946,N_2306,N_991);
nor U6947 (N_6947,N_2875,N_4631);
nand U6948 (N_6948,N_1127,N_165);
or U6949 (N_6949,N_1836,N_4598);
or U6950 (N_6950,N_1524,N_1238);
nand U6951 (N_6951,N_4772,N_2693);
or U6952 (N_6952,N_2054,N_1683);
xnor U6953 (N_6953,N_605,N_468);
nand U6954 (N_6954,N_3216,N_203);
and U6955 (N_6955,N_2328,N_1311);
nor U6956 (N_6956,N_4564,N_4288);
and U6957 (N_6957,N_3616,N_3201);
nor U6958 (N_6958,N_968,N_4484);
nand U6959 (N_6959,N_3826,N_4110);
xnor U6960 (N_6960,N_782,N_453);
xor U6961 (N_6961,N_4093,N_3257);
nand U6962 (N_6962,N_3532,N_2808);
nor U6963 (N_6963,N_723,N_634);
xor U6964 (N_6964,N_3453,N_4474);
nor U6965 (N_6965,N_2737,N_3311);
nand U6966 (N_6966,N_4785,N_2814);
xnor U6967 (N_6967,N_3413,N_1340);
nor U6968 (N_6968,N_4673,N_2142);
and U6969 (N_6969,N_3646,N_4813);
nor U6970 (N_6970,N_4877,N_997);
xor U6971 (N_6971,N_1980,N_2562);
nand U6972 (N_6972,N_2467,N_3566);
nor U6973 (N_6973,N_3688,N_564);
and U6974 (N_6974,N_3774,N_4723);
xor U6975 (N_6975,N_1970,N_250);
nor U6976 (N_6976,N_784,N_4030);
and U6977 (N_6977,N_3571,N_1363);
nand U6978 (N_6978,N_383,N_2678);
nor U6979 (N_6979,N_4108,N_3086);
xor U6980 (N_6980,N_4049,N_2771);
xor U6981 (N_6981,N_3222,N_3820);
or U6982 (N_6982,N_980,N_1319);
xnor U6983 (N_6983,N_4459,N_1370);
nand U6984 (N_6984,N_3540,N_659);
and U6985 (N_6985,N_3919,N_2222);
nand U6986 (N_6986,N_197,N_1719);
xnor U6987 (N_6987,N_531,N_111);
and U6988 (N_6988,N_279,N_2025);
or U6989 (N_6989,N_855,N_3189);
nor U6990 (N_6990,N_1275,N_2251);
nand U6991 (N_6991,N_1400,N_1480);
and U6992 (N_6992,N_2722,N_3461);
or U6993 (N_6993,N_3598,N_3752);
nand U6994 (N_6994,N_4964,N_2172);
nand U6995 (N_6995,N_804,N_108);
and U6996 (N_6996,N_4213,N_593);
nand U6997 (N_6997,N_1281,N_3399);
xnor U6998 (N_6998,N_4624,N_3768);
or U6999 (N_6999,N_1506,N_802);
and U7000 (N_7000,N_177,N_4659);
and U7001 (N_7001,N_2520,N_2070);
xnor U7002 (N_7002,N_1123,N_875);
xor U7003 (N_7003,N_934,N_2613);
or U7004 (N_7004,N_3822,N_4563);
xor U7005 (N_7005,N_1940,N_1486);
or U7006 (N_7006,N_4636,N_4042);
or U7007 (N_7007,N_198,N_4814);
nor U7008 (N_7008,N_1986,N_3552);
xor U7009 (N_7009,N_2243,N_4306);
or U7010 (N_7010,N_2697,N_2215);
or U7011 (N_7011,N_2284,N_4642);
or U7012 (N_7012,N_3197,N_184);
and U7013 (N_7013,N_2501,N_1327);
or U7014 (N_7014,N_4818,N_2852);
or U7015 (N_7015,N_4582,N_1841);
nor U7016 (N_7016,N_2448,N_3124);
and U7017 (N_7017,N_4421,N_4935);
nor U7018 (N_7018,N_2985,N_1879);
nand U7019 (N_7019,N_1508,N_2104);
nand U7020 (N_7020,N_2097,N_3951);
xnor U7021 (N_7021,N_398,N_823);
or U7022 (N_7022,N_3015,N_1117);
xnor U7023 (N_7023,N_1323,N_3144);
xor U7024 (N_7024,N_3875,N_2704);
nand U7025 (N_7025,N_4493,N_500);
xor U7026 (N_7026,N_1236,N_1830);
nor U7027 (N_7027,N_1977,N_1450);
nand U7028 (N_7028,N_4122,N_4729);
or U7029 (N_7029,N_1962,N_4382);
or U7030 (N_7030,N_1594,N_1672);
or U7031 (N_7031,N_2219,N_4751);
or U7032 (N_7032,N_4756,N_3186);
and U7033 (N_7033,N_2619,N_4282);
nand U7034 (N_7034,N_3858,N_4561);
and U7035 (N_7035,N_2638,N_4617);
and U7036 (N_7036,N_3730,N_4787);
nor U7037 (N_7037,N_3574,N_3435);
nor U7038 (N_7038,N_4538,N_2863);
nor U7039 (N_7039,N_852,N_3034);
and U7040 (N_7040,N_2058,N_368);
and U7041 (N_7041,N_2099,N_961);
or U7042 (N_7042,N_4808,N_4102);
nand U7043 (N_7043,N_1129,N_352);
and U7044 (N_7044,N_3320,N_1525);
nor U7045 (N_7045,N_1920,N_2786);
nand U7046 (N_7046,N_2166,N_294);
or U7047 (N_7047,N_4639,N_10);
and U7048 (N_7048,N_632,N_2481);
nor U7049 (N_7049,N_1620,N_2479);
nor U7050 (N_7050,N_1228,N_923);
nand U7051 (N_7051,N_808,N_494);
nand U7052 (N_7052,N_874,N_1949);
xor U7053 (N_7053,N_466,N_1252);
xnor U7054 (N_7054,N_4045,N_1369);
or U7055 (N_7055,N_3377,N_1509);
or U7056 (N_7056,N_388,N_3575);
or U7057 (N_7057,N_3979,N_474);
and U7058 (N_7058,N_4258,N_2206);
and U7059 (N_7059,N_1142,N_1650);
nor U7060 (N_7060,N_4829,N_3548);
nand U7061 (N_7061,N_612,N_1034);
and U7062 (N_7062,N_1098,N_4981);
nor U7063 (N_7063,N_4628,N_3818);
nand U7064 (N_7064,N_1804,N_4283);
nor U7065 (N_7065,N_4034,N_709);
or U7066 (N_7066,N_3534,N_2960);
xnor U7067 (N_7067,N_3398,N_1072);
and U7068 (N_7068,N_2503,N_3245);
or U7069 (N_7069,N_2961,N_2765);
or U7070 (N_7070,N_2636,N_4219);
xnor U7071 (N_7071,N_4225,N_1418);
or U7072 (N_7072,N_2723,N_4438);
nand U7073 (N_7073,N_3385,N_583);
nor U7074 (N_7074,N_2205,N_410);
nor U7075 (N_7075,N_3433,N_3751);
nand U7076 (N_7076,N_3258,N_2348);
xnor U7077 (N_7077,N_1578,N_3285);
or U7078 (N_7078,N_4354,N_3695);
xor U7079 (N_7079,N_598,N_1332);
xor U7080 (N_7080,N_1312,N_950);
or U7081 (N_7081,N_3934,N_4558);
xor U7082 (N_7082,N_4786,N_3366);
or U7083 (N_7083,N_3177,N_842);
or U7084 (N_7084,N_676,N_2310);
xnor U7085 (N_7085,N_919,N_3669);
nand U7086 (N_7086,N_77,N_2551);
nor U7087 (N_7087,N_2040,N_2133);
xor U7088 (N_7088,N_1778,N_1093);
or U7089 (N_7089,N_581,N_4942);
and U7090 (N_7090,N_3166,N_3106);
or U7091 (N_7091,N_167,N_3940);
nand U7092 (N_7092,N_3805,N_1455);
nand U7093 (N_7093,N_4341,N_40);
nor U7094 (N_7094,N_656,N_2004);
nand U7095 (N_7095,N_4169,N_2715);
or U7096 (N_7096,N_1164,N_4615);
xnor U7097 (N_7097,N_2279,N_1722);
or U7098 (N_7098,N_3634,N_4000);
and U7099 (N_7099,N_4905,N_2191);
nand U7100 (N_7100,N_2116,N_79);
xor U7101 (N_7101,N_334,N_1475);
nor U7102 (N_7102,N_387,N_965);
nor U7103 (N_7103,N_438,N_3569);
nor U7104 (N_7104,N_4458,N_2712);
and U7105 (N_7105,N_3279,N_4348);
nand U7106 (N_7106,N_3912,N_3636);
nor U7107 (N_7107,N_4523,N_3868);
xor U7108 (N_7108,N_139,N_553);
or U7109 (N_7109,N_430,N_224);
and U7110 (N_7110,N_513,N_2499);
xnor U7111 (N_7111,N_4010,N_2865);
nand U7112 (N_7112,N_2148,N_2344);
xnor U7113 (N_7113,N_4985,N_2465);
nor U7114 (N_7114,N_2994,N_2646);
nand U7115 (N_7115,N_4070,N_3443);
and U7116 (N_7116,N_3838,N_1229);
or U7117 (N_7117,N_4247,N_4038);
nand U7118 (N_7118,N_3664,N_1691);
xnor U7119 (N_7119,N_2457,N_2368);
and U7120 (N_7120,N_689,N_642);
and U7121 (N_7121,N_2224,N_691);
and U7122 (N_7122,N_3152,N_4711);
and U7123 (N_7123,N_1870,N_1941);
or U7124 (N_7124,N_2091,N_1324);
nand U7125 (N_7125,N_435,N_2334);
xnor U7126 (N_7126,N_2705,N_4155);
nor U7127 (N_7127,N_3074,N_2447);
xnor U7128 (N_7128,N_1112,N_101);
nor U7129 (N_7129,N_1555,N_4679);
and U7130 (N_7130,N_2833,N_1014);
or U7131 (N_7131,N_1122,N_1591);
nand U7132 (N_7132,N_1207,N_1339);
nand U7133 (N_7133,N_296,N_2999);
xnor U7134 (N_7134,N_1642,N_4252);
nor U7135 (N_7135,N_4765,N_1910);
and U7136 (N_7136,N_463,N_3965);
nor U7137 (N_7137,N_88,N_2049);
nand U7138 (N_7138,N_2524,N_540);
xnor U7139 (N_7139,N_932,N_2711);
nand U7140 (N_7140,N_1128,N_1504);
and U7141 (N_7141,N_73,N_3586);
nor U7142 (N_7142,N_877,N_3971);
or U7143 (N_7143,N_523,N_1614);
nand U7144 (N_7144,N_4546,N_4672);
nand U7145 (N_7145,N_974,N_975);
or U7146 (N_7146,N_4549,N_3680);
or U7147 (N_7147,N_2173,N_4278);
or U7148 (N_7148,N_2623,N_2703);
xnor U7149 (N_7149,N_4347,N_3722);
xor U7150 (N_7150,N_2701,N_560);
or U7151 (N_7151,N_1202,N_2548);
or U7152 (N_7152,N_2378,N_458);
xnor U7153 (N_7153,N_2734,N_1076);
and U7154 (N_7154,N_2470,N_1718);
and U7155 (N_7155,N_1199,N_14);
nor U7156 (N_7156,N_2302,N_1216);
or U7157 (N_7157,N_1802,N_4031);
xnor U7158 (N_7158,N_455,N_65);
nand U7159 (N_7159,N_1939,N_725);
and U7160 (N_7160,N_555,N_2390);
xnor U7161 (N_7161,N_1456,N_1420);
nor U7162 (N_7162,N_3459,N_1956);
xor U7163 (N_7163,N_1913,N_3585);
and U7164 (N_7164,N_4346,N_1457);
xor U7165 (N_7165,N_4514,N_1599);
nand U7166 (N_7166,N_2972,N_2432);
or U7167 (N_7167,N_3498,N_1084);
or U7168 (N_7168,N_4392,N_1188);
and U7169 (N_7169,N_479,N_978);
and U7170 (N_7170,N_168,N_4901);
or U7171 (N_7171,N_3055,N_57);
nor U7172 (N_7172,N_3842,N_201);
or U7173 (N_7173,N_3990,N_1534);
xnor U7174 (N_7174,N_972,N_130);
nor U7175 (N_7175,N_3806,N_4249);
nor U7176 (N_7176,N_4362,N_1219);
nand U7177 (N_7177,N_1412,N_3215);
nand U7178 (N_7178,N_3417,N_1265);
nand U7179 (N_7179,N_12,N_2812);
or U7180 (N_7180,N_498,N_115);
nor U7181 (N_7181,N_3388,N_1577);
nand U7182 (N_7182,N_3333,N_611);
or U7183 (N_7183,N_4019,N_880);
nand U7184 (N_7184,N_4914,N_1880);
nor U7185 (N_7185,N_3142,N_4994);
nand U7186 (N_7186,N_3817,N_3013);
nor U7187 (N_7187,N_1203,N_3903);
xnor U7188 (N_7188,N_4892,N_1988);
nor U7189 (N_7189,N_607,N_3667);
xor U7190 (N_7190,N_3717,N_1201);
xor U7191 (N_7191,N_1496,N_3792);
and U7192 (N_7192,N_3927,N_2662);
nand U7193 (N_7193,N_1361,N_1978);
or U7194 (N_7194,N_4678,N_71);
nand U7195 (N_7195,N_1211,N_1383);
and U7196 (N_7196,N_4830,N_4960);
nor U7197 (N_7197,N_1237,N_1934);
xnor U7198 (N_7198,N_3481,N_1644);
and U7199 (N_7199,N_3081,N_4912);
xor U7200 (N_7200,N_3605,N_2071);
nand U7201 (N_7201,N_1592,N_3018);
nor U7202 (N_7202,N_3458,N_278);
or U7203 (N_7203,N_4965,N_3008);
and U7204 (N_7204,N_2033,N_1603);
xor U7205 (N_7205,N_916,N_4251);
nor U7206 (N_7206,N_2486,N_3014);
or U7207 (N_7207,N_4668,N_4748);
and U7208 (N_7208,N_361,N_106);
nand U7209 (N_7209,N_1077,N_443);
xnor U7210 (N_7210,N_4873,N_1559);
nor U7211 (N_7211,N_3728,N_794);
xnor U7212 (N_7212,N_2115,N_1474);
nor U7213 (N_7213,N_2537,N_830);
xor U7214 (N_7214,N_2898,N_2188);
nor U7215 (N_7215,N_2184,N_4667);
nor U7216 (N_7216,N_4651,N_3754);
and U7217 (N_7217,N_509,N_1390);
xnor U7218 (N_7218,N_3655,N_3964);
nor U7219 (N_7219,N_3924,N_1511);
or U7220 (N_7220,N_4757,N_2796);
and U7221 (N_7221,N_355,N_49);
xor U7222 (N_7222,N_2905,N_1029);
or U7223 (N_7223,N_1043,N_208);
and U7224 (N_7224,N_902,N_385);
and U7225 (N_7225,N_1343,N_4127);
and U7226 (N_7226,N_1315,N_48);
or U7227 (N_7227,N_3327,N_4198);
and U7228 (N_7228,N_2967,N_4056);
nand U7229 (N_7229,N_2963,N_149);
nand U7230 (N_7230,N_674,N_1569);
and U7231 (N_7231,N_2434,N_4888);
nor U7232 (N_7232,N_4145,N_847);
or U7233 (N_7233,N_625,N_603);
nor U7234 (N_7234,N_763,N_3101);
and U7235 (N_7235,N_3065,N_2545);
xnor U7236 (N_7236,N_1046,N_525);
or U7237 (N_7237,N_726,N_1494);
nor U7238 (N_7238,N_1438,N_1643);
and U7239 (N_7239,N_1411,N_1834);
nand U7240 (N_7240,N_4350,N_2000);
xnor U7241 (N_7241,N_4689,N_1442);
nand U7242 (N_7242,N_3791,N_3678);
or U7243 (N_7243,N_2789,N_948);
xor U7244 (N_7244,N_735,N_3431);
nor U7245 (N_7245,N_775,N_3268);
and U7246 (N_7246,N_345,N_2367);
and U7247 (N_7247,N_3689,N_262);
xor U7248 (N_7248,N_2186,N_1582);
nor U7249 (N_7249,N_4836,N_456);
xor U7250 (N_7250,N_4504,N_1563);
xor U7251 (N_7251,N_4645,N_4580);
nor U7252 (N_7252,N_721,N_2087);
and U7253 (N_7253,N_4334,N_4161);
nor U7254 (N_7254,N_2842,N_2857);
and U7255 (N_7255,N_2414,N_921);
and U7256 (N_7256,N_4611,N_836);
xor U7257 (N_7257,N_1462,N_1766);
or U7258 (N_7258,N_2349,N_918);
xor U7259 (N_7259,N_2427,N_1180);
nor U7260 (N_7260,N_574,N_1558);
xor U7261 (N_7261,N_4197,N_3363);
xor U7262 (N_7262,N_1086,N_664);
or U7263 (N_7263,N_4515,N_3677);
and U7264 (N_7264,N_2885,N_2325);
and U7265 (N_7265,N_2614,N_3892);
or U7266 (N_7266,N_2276,N_4726);
and U7267 (N_7267,N_1366,N_4112);
and U7268 (N_7268,N_1777,N_4872);
nand U7269 (N_7269,N_915,N_3184);
nand U7270 (N_7270,N_2492,N_575);
nor U7271 (N_7271,N_1156,N_1337);
nor U7272 (N_7272,N_152,N_2570);
and U7273 (N_7273,N_3181,N_3773);
nand U7274 (N_7274,N_1482,N_803);
or U7275 (N_7275,N_2589,N_2719);
xnor U7276 (N_7276,N_2511,N_4577);
nor U7277 (N_7277,N_543,N_2237);
or U7278 (N_7278,N_3772,N_379);
nor U7279 (N_7279,N_4248,N_4002);
xor U7280 (N_7280,N_3056,N_4567);
xor U7281 (N_7281,N_4686,N_3706);
xor U7282 (N_7282,N_742,N_1954);
xor U7283 (N_7283,N_571,N_459);
xor U7284 (N_7284,N_4305,N_903);
or U7285 (N_7285,N_1600,N_4356);
nor U7286 (N_7286,N_4074,N_62);
nor U7287 (N_7287,N_1894,N_3810);
or U7288 (N_7288,N_4496,N_4963);
xnor U7289 (N_7289,N_4842,N_4469);
nand U7290 (N_7290,N_778,N_2475);
and U7291 (N_7291,N_3303,N_3010);
and U7292 (N_7292,N_729,N_2926);
nand U7293 (N_7293,N_679,N_1515);
nand U7294 (N_7294,N_3666,N_3037);
xor U7295 (N_7295,N_4018,N_2256);
nand U7296 (N_7296,N_2074,N_3866);
nand U7297 (N_7297,N_4040,N_1914);
or U7298 (N_7298,N_1540,N_1655);
or U7299 (N_7299,N_2018,N_962);
nor U7300 (N_7300,N_4026,N_3985);
or U7301 (N_7301,N_502,N_2731);
xor U7302 (N_7302,N_2527,N_1158);
xor U7303 (N_7303,N_4215,N_2618);
xnor U7304 (N_7304,N_4688,N_4670);
and U7305 (N_7305,N_2093,N_924);
xor U7306 (N_7306,N_4655,N_4365);
nor U7307 (N_7307,N_174,N_4996);
and U7308 (N_7308,N_1745,N_890);
and U7309 (N_7309,N_4604,N_2446);
or U7310 (N_7310,N_1527,N_367);
xor U7311 (N_7311,N_4029,N_635);
nor U7312 (N_7312,N_1609,N_4768);
nor U7313 (N_7313,N_1198,N_1684);
or U7314 (N_7314,N_2621,N_896);
nand U7315 (N_7315,N_1903,N_773);
xnor U7316 (N_7316,N_3317,N_953);
xnor U7317 (N_7317,N_3701,N_3843);
or U7318 (N_7318,N_3950,N_326);
xor U7319 (N_7319,N_2610,N_3456);
nor U7320 (N_7320,N_4437,N_2640);
and U7321 (N_7321,N_2913,N_2290);
xor U7322 (N_7322,N_4011,N_1670);
xor U7323 (N_7323,N_2089,N_4866);
xnor U7324 (N_7324,N_4292,N_559);
xnor U7325 (N_7325,N_2182,N_1539);
nand U7326 (N_7326,N_3835,N_3246);
and U7327 (N_7327,N_4319,N_406);
nand U7328 (N_7328,N_2158,N_4020);
xor U7329 (N_7329,N_1376,N_1012);
nor U7330 (N_7330,N_146,N_1667);
nand U7331 (N_7331,N_3595,N_4916);
and U7332 (N_7332,N_4090,N_1979);
and U7333 (N_7333,N_76,N_1839);
nor U7334 (N_7334,N_2293,N_3864);
or U7335 (N_7335,N_4381,N_3437);
nand U7336 (N_7336,N_3753,N_4706);
nand U7337 (N_7337,N_1081,N_154);
nor U7338 (N_7338,N_3923,N_1707);
xor U7339 (N_7339,N_945,N_467);
nor U7340 (N_7340,N_4025,N_3819);
xnor U7341 (N_7341,N_694,N_4083);
or U7342 (N_7342,N_3663,N_562);
xor U7343 (N_7343,N_1107,N_4439);
and U7344 (N_7344,N_2156,N_3040);
xnor U7345 (N_7345,N_4244,N_927);
and U7346 (N_7346,N_1717,N_2540);
xor U7347 (N_7347,N_3803,N_3357);
nor U7348 (N_7348,N_1795,N_1045);
and U7349 (N_7349,N_2516,N_1176);
or U7350 (N_7350,N_539,N_3150);
xor U7351 (N_7351,N_200,N_1668);
or U7352 (N_7352,N_3312,N_3627);
nand U7353 (N_7353,N_3518,N_3778);
nor U7354 (N_7354,N_306,N_3501);
nand U7355 (N_7355,N_601,N_2762);
nor U7356 (N_7356,N_3109,N_3651);
nor U7357 (N_7357,N_2218,N_4417);
and U7358 (N_7358,N_2452,N_261);
nor U7359 (N_7359,N_3969,N_3725);
nor U7360 (N_7360,N_2019,N_1139);
nor U7361 (N_7361,N_4391,N_2126);
and U7362 (N_7362,N_3252,N_3732);
xor U7363 (N_7363,N_3149,N_2746);
xnor U7364 (N_7364,N_4940,N_776);
nand U7365 (N_7365,N_3114,N_3188);
xnor U7366 (N_7366,N_2361,N_3314);
nor U7367 (N_7367,N_2968,N_4095);
xor U7368 (N_7368,N_4973,N_75);
nand U7369 (N_7369,N_3098,N_382);
xnor U7370 (N_7370,N_4548,N_1945);
nor U7371 (N_7371,N_2770,N_2989);
or U7372 (N_7372,N_1583,N_3691);
nand U7373 (N_7373,N_1397,N_3783);
or U7374 (N_7374,N_2149,N_2299);
and U7375 (N_7375,N_3777,N_4461);
xnor U7376 (N_7376,N_2382,N_3849);
nor U7377 (N_7377,N_4460,N_1871);
nand U7378 (N_7378,N_4970,N_4712);
nand U7379 (N_7379,N_680,N_3206);
nand U7380 (N_7380,N_851,N_4606);
nor U7381 (N_7381,N_2241,N_793);
nor U7382 (N_7382,N_4568,N_2561);
xor U7383 (N_7383,N_2854,N_2080);
xnor U7384 (N_7384,N_2882,N_3163);
nand U7385 (N_7385,N_835,N_1368);
xnor U7386 (N_7386,N_1865,N_2343);
nand U7387 (N_7387,N_3058,N_4379);
nand U7388 (N_7388,N_1638,N_54);
nor U7389 (N_7389,N_1801,N_3542);
nor U7390 (N_7390,N_4263,N_4847);
nand U7391 (N_7391,N_3190,N_4554);
xor U7392 (N_7392,N_128,N_4926);
nand U7393 (N_7393,N_4165,N_3112);
and U7394 (N_7394,N_952,N_4693);
xor U7395 (N_7395,N_4087,N_3402);
nand U7396 (N_7396,N_1116,N_1037);
nor U7397 (N_7397,N_2203,N_3784);
xnor U7398 (N_7398,N_3961,N_1090);
nand U7399 (N_7399,N_4370,N_473);
nor U7400 (N_7400,N_1145,N_3579);
and U7401 (N_7401,N_3917,N_752);
xnor U7402 (N_7402,N_2706,N_3495);
nor U7403 (N_7403,N_2232,N_1520);
or U7404 (N_7404,N_4471,N_3143);
nand U7405 (N_7405,N_2140,N_925);
nand U7406 (N_7406,N_4817,N_791);
nand U7407 (N_7407,N_1669,N_1579);
nor U7408 (N_7408,N_4314,N_3251);
xor U7409 (N_7409,N_4205,N_1713);
xnor U7410 (N_7410,N_4510,N_4457);
or U7411 (N_7411,N_3200,N_1057);
and U7412 (N_7412,N_4061,N_2023);
xnor U7413 (N_7413,N_3408,N_643);
and U7414 (N_7414,N_3107,N_2391);
and U7415 (N_7415,N_3720,N_1213);
nor U7416 (N_7416,N_4573,N_768);
nand U7417 (N_7417,N_2754,N_824);
xor U7418 (N_7418,N_4544,N_3295);
nor U7419 (N_7419,N_3568,N_3020);
or U7420 (N_7420,N_4221,N_4369);
or U7421 (N_7421,N_3512,N_4271);
or U7422 (N_7422,N_3299,N_1771);
nor U7423 (N_7423,N_2190,N_4104);
nor U7424 (N_7424,N_536,N_4735);
or U7425 (N_7425,N_28,N_3708);
and U7426 (N_7426,N_712,N_3746);
or U7427 (N_7427,N_485,N_1257);
nor U7428 (N_7428,N_2597,N_4325);
nand U7429 (N_7429,N_2490,N_1433);
xor U7430 (N_7430,N_3526,N_4181);
xnor U7431 (N_7431,N_578,N_2639);
nand U7432 (N_7432,N_859,N_1101);
nand U7433 (N_7433,N_3794,N_1387);
xor U7434 (N_7434,N_4376,N_1367);
and U7435 (N_7435,N_2034,N_1602);
nand U7436 (N_7436,N_2101,N_982);
xnor U7437 (N_7437,N_3840,N_1787);
and U7438 (N_7438,N_1500,N_1206);
nand U7439 (N_7439,N_3888,N_45);
nand U7440 (N_7440,N_1799,N_1110);
nor U7441 (N_7441,N_2045,N_2954);
nand U7442 (N_7442,N_4623,N_4312);
or U7443 (N_7443,N_4224,N_2575);
or U7444 (N_7444,N_2407,N_1283);
nor U7445 (N_7445,N_4497,N_1860);
or U7446 (N_7446,N_123,N_194);
nor U7447 (N_7447,N_1240,N_140);
nand U7448 (N_7448,N_4797,N_476);
nand U7449 (N_7449,N_2416,N_1725);
or U7450 (N_7450,N_3996,N_2958);
or U7451 (N_7451,N_3487,N_582);
or U7452 (N_7452,N_448,N_1291);
or U7453 (N_7453,N_2197,N_4870);
and U7454 (N_7454,N_2260,N_1292);
nand U7455 (N_7455,N_2767,N_2569);
and U7456 (N_7456,N_310,N_3221);
nor U7457 (N_7457,N_121,N_3386);
xnor U7458 (N_7458,N_1790,N_251);
and U7459 (N_7459,N_3499,N_1423);
or U7460 (N_7460,N_2315,N_493);
or U7461 (N_7461,N_3787,N_1924);
or U7462 (N_7462,N_2709,N_4718);
nor U7463 (N_7463,N_4553,N_4297);
nand U7464 (N_7464,N_2879,N_2727);
xnor U7465 (N_7465,N_3129,N_1615);
nand U7466 (N_7466,N_858,N_3095);
nand U7467 (N_7467,N_1183,N_1957);
nor U7468 (N_7468,N_772,N_380);
and U7469 (N_7469,N_209,N_4448);
xnor U7470 (N_7470,N_4930,N_515);
or U7471 (N_7471,N_3963,N_2291);
xnor U7472 (N_7472,N_80,N_39);
nand U7473 (N_7473,N_490,N_4084);
nand U7474 (N_7474,N_2740,N_1889);
nor U7475 (N_7475,N_4162,N_2408);
xnor U7476 (N_7476,N_3009,N_404);
nor U7477 (N_7477,N_1241,N_3330);
nor U7478 (N_7478,N_1031,N_3604);
and U7479 (N_7479,N_1300,N_3897);
xor U7480 (N_7480,N_3553,N_4677);
nand U7481 (N_7481,N_2534,N_4296);
or U7482 (N_7482,N_892,N_2420);
and U7483 (N_7483,N_2164,N_431);
xor U7484 (N_7484,N_4699,N_3642);
nand U7485 (N_7485,N_1983,N_2574);
nor U7486 (N_7486,N_579,N_812);
nand U7487 (N_7487,N_3906,N_3839);
nand U7488 (N_7488,N_2939,N_3878);
and U7489 (N_7489,N_3967,N_4058);
nand U7490 (N_7490,N_4453,N_660);
nor U7491 (N_7491,N_3643,N_4239);
or U7492 (N_7492,N_227,N_1973);
nor U7493 (N_7493,N_3944,N_4186);
nor U7494 (N_7494,N_3665,N_416);
nand U7495 (N_7495,N_3204,N_1378);
or U7496 (N_7496,N_4452,N_2832);
or U7497 (N_7497,N_1688,N_3147);
nand U7498 (N_7498,N_2105,N_2225);
nor U7499 (N_7499,N_1708,N_3448);
nand U7500 (N_7500,N_152,N_992);
or U7501 (N_7501,N_3056,N_2861);
and U7502 (N_7502,N_2978,N_3347);
nor U7503 (N_7503,N_624,N_3657);
or U7504 (N_7504,N_292,N_2258);
nor U7505 (N_7505,N_1481,N_1536);
or U7506 (N_7506,N_4976,N_1807);
nor U7507 (N_7507,N_1798,N_3153);
nand U7508 (N_7508,N_3281,N_4409);
and U7509 (N_7509,N_3343,N_3496);
or U7510 (N_7510,N_884,N_40);
nor U7511 (N_7511,N_1103,N_1979);
nor U7512 (N_7512,N_4361,N_2115);
and U7513 (N_7513,N_3786,N_2471);
nand U7514 (N_7514,N_4648,N_4571);
nand U7515 (N_7515,N_2086,N_2663);
xor U7516 (N_7516,N_1202,N_3752);
and U7517 (N_7517,N_2539,N_3067);
nand U7518 (N_7518,N_1721,N_846);
and U7519 (N_7519,N_4238,N_4545);
xnor U7520 (N_7520,N_3244,N_795);
xnor U7521 (N_7521,N_643,N_4457);
xnor U7522 (N_7522,N_2718,N_406);
nor U7523 (N_7523,N_2684,N_3468);
nand U7524 (N_7524,N_2784,N_2134);
nand U7525 (N_7525,N_782,N_1894);
and U7526 (N_7526,N_4863,N_2943);
and U7527 (N_7527,N_3131,N_2000);
nor U7528 (N_7528,N_2236,N_2515);
and U7529 (N_7529,N_1953,N_3337);
xor U7530 (N_7530,N_34,N_4154);
nor U7531 (N_7531,N_4466,N_4877);
nand U7532 (N_7532,N_3135,N_2500);
nor U7533 (N_7533,N_2907,N_1683);
and U7534 (N_7534,N_4355,N_4977);
nor U7535 (N_7535,N_2360,N_159);
nor U7536 (N_7536,N_483,N_2509);
and U7537 (N_7537,N_355,N_4586);
or U7538 (N_7538,N_4878,N_679);
xor U7539 (N_7539,N_4289,N_2879);
xor U7540 (N_7540,N_235,N_2166);
and U7541 (N_7541,N_2119,N_2337);
and U7542 (N_7542,N_1910,N_2134);
nor U7543 (N_7543,N_1035,N_3538);
nand U7544 (N_7544,N_4558,N_2566);
nor U7545 (N_7545,N_4634,N_4963);
and U7546 (N_7546,N_4522,N_3649);
nor U7547 (N_7547,N_2938,N_1406);
and U7548 (N_7548,N_1727,N_3558);
and U7549 (N_7549,N_385,N_4744);
or U7550 (N_7550,N_4716,N_3144);
nor U7551 (N_7551,N_501,N_1653);
nor U7552 (N_7552,N_4390,N_409);
xor U7553 (N_7553,N_4147,N_1266);
xor U7554 (N_7554,N_2547,N_2797);
nand U7555 (N_7555,N_4904,N_3108);
xor U7556 (N_7556,N_4728,N_1985);
or U7557 (N_7557,N_1345,N_4508);
or U7558 (N_7558,N_2552,N_3809);
and U7559 (N_7559,N_4725,N_3197);
or U7560 (N_7560,N_863,N_2913);
xor U7561 (N_7561,N_1884,N_3421);
nor U7562 (N_7562,N_3983,N_2104);
nand U7563 (N_7563,N_3858,N_3533);
and U7564 (N_7564,N_4179,N_606);
xor U7565 (N_7565,N_1689,N_1285);
nor U7566 (N_7566,N_4151,N_2848);
nand U7567 (N_7567,N_3028,N_4780);
and U7568 (N_7568,N_2117,N_1215);
nor U7569 (N_7569,N_3658,N_4025);
nand U7570 (N_7570,N_947,N_4611);
xnor U7571 (N_7571,N_2677,N_1854);
and U7572 (N_7572,N_1870,N_4906);
and U7573 (N_7573,N_393,N_184);
and U7574 (N_7574,N_2353,N_1498);
nand U7575 (N_7575,N_2052,N_3114);
and U7576 (N_7576,N_1627,N_3777);
xnor U7577 (N_7577,N_1808,N_938);
nand U7578 (N_7578,N_4596,N_1791);
xnor U7579 (N_7579,N_3577,N_1004);
and U7580 (N_7580,N_3450,N_178);
and U7581 (N_7581,N_4488,N_592);
nand U7582 (N_7582,N_76,N_3121);
and U7583 (N_7583,N_2571,N_2660);
or U7584 (N_7584,N_4334,N_2909);
or U7585 (N_7585,N_721,N_1025);
and U7586 (N_7586,N_3071,N_1393);
xnor U7587 (N_7587,N_1538,N_1098);
nor U7588 (N_7588,N_463,N_4475);
or U7589 (N_7589,N_1260,N_2005);
nor U7590 (N_7590,N_3749,N_542);
nand U7591 (N_7591,N_18,N_253);
nand U7592 (N_7592,N_3301,N_115);
nor U7593 (N_7593,N_4205,N_925);
nand U7594 (N_7594,N_3910,N_3504);
or U7595 (N_7595,N_4439,N_1595);
nand U7596 (N_7596,N_4591,N_1779);
nor U7597 (N_7597,N_1061,N_2643);
or U7598 (N_7598,N_3067,N_4667);
or U7599 (N_7599,N_1874,N_2516);
xnor U7600 (N_7600,N_1084,N_3139);
or U7601 (N_7601,N_2234,N_3487);
or U7602 (N_7602,N_2600,N_3984);
and U7603 (N_7603,N_1020,N_4160);
nand U7604 (N_7604,N_1237,N_3242);
or U7605 (N_7605,N_1554,N_4225);
or U7606 (N_7606,N_3620,N_1049);
xnor U7607 (N_7607,N_3243,N_4091);
nand U7608 (N_7608,N_2841,N_779);
xnor U7609 (N_7609,N_578,N_4462);
xnor U7610 (N_7610,N_4445,N_3840);
or U7611 (N_7611,N_2260,N_2727);
xnor U7612 (N_7612,N_3467,N_90);
xnor U7613 (N_7613,N_4177,N_3465);
nand U7614 (N_7614,N_3831,N_1921);
or U7615 (N_7615,N_768,N_1461);
and U7616 (N_7616,N_1503,N_420);
or U7617 (N_7617,N_4353,N_3845);
nor U7618 (N_7618,N_4599,N_1893);
nand U7619 (N_7619,N_2204,N_1472);
xor U7620 (N_7620,N_4291,N_999);
nand U7621 (N_7621,N_2220,N_3160);
or U7622 (N_7622,N_4126,N_1283);
and U7623 (N_7623,N_1006,N_1283);
nand U7624 (N_7624,N_4375,N_2535);
nor U7625 (N_7625,N_3029,N_2053);
nor U7626 (N_7626,N_3683,N_3087);
nand U7627 (N_7627,N_1758,N_1613);
nor U7628 (N_7628,N_961,N_4233);
or U7629 (N_7629,N_203,N_4398);
xnor U7630 (N_7630,N_2356,N_2168);
and U7631 (N_7631,N_1811,N_923);
xnor U7632 (N_7632,N_1543,N_2053);
and U7633 (N_7633,N_4032,N_3635);
xor U7634 (N_7634,N_1348,N_873);
and U7635 (N_7635,N_1712,N_2929);
and U7636 (N_7636,N_3725,N_2070);
and U7637 (N_7637,N_3442,N_1337);
or U7638 (N_7638,N_3483,N_4429);
nand U7639 (N_7639,N_1179,N_3318);
or U7640 (N_7640,N_2067,N_4614);
xor U7641 (N_7641,N_2989,N_3225);
or U7642 (N_7642,N_2302,N_1733);
nor U7643 (N_7643,N_1881,N_2404);
nor U7644 (N_7644,N_2867,N_760);
xnor U7645 (N_7645,N_1410,N_2383);
xnor U7646 (N_7646,N_4705,N_1906);
nand U7647 (N_7647,N_3225,N_2959);
nor U7648 (N_7648,N_1817,N_2794);
nor U7649 (N_7649,N_969,N_4021);
or U7650 (N_7650,N_1354,N_2007);
or U7651 (N_7651,N_4048,N_159);
nand U7652 (N_7652,N_3375,N_2862);
nand U7653 (N_7653,N_203,N_1420);
and U7654 (N_7654,N_3777,N_1703);
xnor U7655 (N_7655,N_1585,N_1121);
and U7656 (N_7656,N_2478,N_4597);
nor U7657 (N_7657,N_3010,N_1672);
or U7658 (N_7658,N_4204,N_2997);
or U7659 (N_7659,N_130,N_3306);
or U7660 (N_7660,N_465,N_2734);
xnor U7661 (N_7661,N_1191,N_2559);
or U7662 (N_7662,N_1483,N_2030);
xor U7663 (N_7663,N_3131,N_2773);
nand U7664 (N_7664,N_502,N_546);
or U7665 (N_7665,N_2071,N_1654);
xnor U7666 (N_7666,N_855,N_3696);
xor U7667 (N_7667,N_3211,N_2929);
nor U7668 (N_7668,N_3099,N_4755);
xor U7669 (N_7669,N_3138,N_3504);
nor U7670 (N_7670,N_181,N_4356);
xnor U7671 (N_7671,N_533,N_4549);
nor U7672 (N_7672,N_364,N_2498);
or U7673 (N_7673,N_4873,N_1870);
nor U7674 (N_7674,N_2949,N_4878);
nor U7675 (N_7675,N_2791,N_3908);
and U7676 (N_7676,N_2191,N_2591);
and U7677 (N_7677,N_4775,N_1148);
and U7678 (N_7678,N_668,N_451);
nand U7679 (N_7679,N_1101,N_3081);
and U7680 (N_7680,N_442,N_161);
or U7681 (N_7681,N_4065,N_3829);
nor U7682 (N_7682,N_1491,N_4116);
nor U7683 (N_7683,N_3265,N_4415);
or U7684 (N_7684,N_2376,N_1315);
nand U7685 (N_7685,N_1127,N_1289);
and U7686 (N_7686,N_2258,N_338);
xnor U7687 (N_7687,N_2599,N_4186);
xor U7688 (N_7688,N_4968,N_4410);
or U7689 (N_7689,N_129,N_1567);
nor U7690 (N_7690,N_591,N_1501);
and U7691 (N_7691,N_63,N_3715);
xor U7692 (N_7692,N_3471,N_4305);
nand U7693 (N_7693,N_3043,N_3674);
nor U7694 (N_7694,N_1849,N_3387);
nor U7695 (N_7695,N_866,N_206);
nor U7696 (N_7696,N_3819,N_3241);
xor U7697 (N_7697,N_471,N_318);
nor U7698 (N_7698,N_2770,N_3097);
xnor U7699 (N_7699,N_2053,N_1386);
and U7700 (N_7700,N_11,N_969);
or U7701 (N_7701,N_4489,N_40);
nand U7702 (N_7702,N_4782,N_1950);
nand U7703 (N_7703,N_4200,N_4163);
xor U7704 (N_7704,N_1892,N_882);
nand U7705 (N_7705,N_2342,N_1889);
and U7706 (N_7706,N_4977,N_876);
xnor U7707 (N_7707,N_2076,N_2407);
nor U7708 (N_7708,N_1666,N_1278);
or U7709 (N_7709,N_1281,N_4249);
nor U7710 (N_7710,N_33,N_2918);
and U7711 (N_7711,N_1822,N_91);
and U7712 (N_7712,N_2360,N_1863);
or U7713 (N_7713,N_1278,N_4535);
and U7714 (N_7714,N_527,N_628);
xnor U7715 (N_7715,N_2912,N_992);
or U7716 (N_7716,N_3368,N_3994);
nand U7717 (N_7717,N_1443,N_572);
and U7718 (N_7718,N_2772,N_281);
and U7719 (N_7719,N_2700,N_2789);
and U7720 (N_7720,N_3307,N_2826);
nor U7721 (N_7721,N_4612,N_70);
xnor U7722 (N_7722,N_1695,N_2636);
or U7723 (N_7723,N_1701,N_1352);
nand U7724 (N_7724,N_1317,N_2736);
xnor U7725 (N_7725,N_2752,N_4038);
and U7726 (N_7726,N_4866,N_686);
nor U7727 (N_7727,N_3402,N_1290);
xnor U7728 (N_7728,N_2430,N_2195);
xor U7729 (N_7729,N_4835,N_2805);
xor U7730 (N_7730,N_795,N_1250);
and U7731 (N_7731,N_3611,N_3932);
and U7732 (N_7732,N_4764,N_3909);
and U7733 (N_7733,N_1300,N_4061);
nor U7734 (N_7734,N_4605,N_2484);
nor U7735 (N_7735,N_656,N_3337);
and U7736 (N_7736,N_3654,N_279);
or U7737 (N_7737,N_520,N_212);
nor U7738 (N_7738,N_2947,N_520);
or U7739 (N_7739,N_1357,N_1912);
nand U7740 (N_7740,N_1252,N_3524);
xnor U7741 (N_7741,N_9,N_4187);
nand U7742 (N_7742,N_904,N_2996);
or U7743 (N_7743,N_1422,N_356);
and U7744 (N_7744,N_2047,N_3472);
nor U7745 (N_7745,N_4573,N_137);
xor U7746 (N_7746,N_2957,N_1000);
or U7747 (N_7747,N_577,N_4537);
and U7748 (N_7748,N_4329,N_3186);
nor U7749 (N_7749,N_985,N_1053);
and U7750 (N_7750,N_1726,N_3964);
and U7751 (N_7751,N_3318,N_3197);
nand U7752 (N_7752,N_4987,N_2277);
xnor U7753 (N_7753,N_1459,N_139);
nor U7754 (N_7754,N_3713,N_540);
and U7755 (N_7755,N_438,N_3535);
nor U7756 (N_7756,N_4644,N_3700);
nor U7757 (N_7757,N_256,N_359);
or U7758 (N_7758,N_1104,N_778);
and U7759 (N_7759,N_1900,N_1506);
nand U7760 (N_7760,N_3785,N_4935);
or U7761 (N_7761,N_4815,N_4370);
or U7762 (N_7762,N_1313,N_3211);
or U7763 (N_7763,N_1058,N_2314);
and U7764 (N_7764,N_4704,N_2692);
and U7765 (N_7765,N_2997,N_123);
and U7766 (N_7766,N_4578,N_1709);
and U7767 (N_7767,N_3569,N_2059);
nand U7768 (N_7768,N_3459,N_2513);
and U7769 (N_7769,N_3374,N_734);
nor U7770 (N_7770,N_525,N_3767);
and U7771 (N_7771,N_1363,N_2080);
xnor U7772 (N_7772,N_3487,N_1431);
nor U7773 (N_7773,N_3687,N_1407);
nor U7774 (N_7774,N_3033,N_1569);
nand U7775 (N_7775,N_4328,N_2595);
or U7776 (N_7776,N_2329,N_2727);
and U7777 (N_7777,N_3104,N_1298);
and U7778 (N_7778,N_2090,N_4020);
and U7779 (N_7779,N_1967,N_1000);
or U7780 (N_7780,N_17,N_2363);
xnor U7781 (N_7781,N_300,N_2666);
and U7782 (N_7782,N_202,N_3483);
or U7783 (N_7783,N_2429,N_102);
nand U7784 (N_7784,N_3334,N_116);
or U7785 (N_7785,N_2617,N_238);
nor U7786 (N_7786,N_4233,N_3198);
xnor U7787 (N_7787,N_531,N_86);
nor U7788 (N_7788,N_4220,N_2719);
xnor U7789 (N_7789,N_1634,N_568);
and U7790 (N_7790,N_4526,N_3354);
xnor U7791 (N_7791,N_3761,N_4829);
nor U7792 (N_7792,N_4403,N_2903);
xnor U7793 (N_7793,N_4818,N_2998);
and U7794 (N_7794,N_4826,N_4567);
and U7795 (N_7795,N_524,N_133);
xnor U7796 (N_7796,N_2618,N_1656);
nand U7797 (N_7797,N_3883,N_1720);
and U7798 (N_7798,N_3434,N_2235);
or U7799 (N_7799,N_4193,N_129);
nor U7800 (N_7800,N_2585,N_4293);
nand U7801 (N_7801,N_510,N_4147);
xnor U7802 (N_7802,N_4238,N_948);
or U7803 (N_7803,N_185,N_3762);
nor U7804 (N_7804,N_1998,N_3122);
xor U7805 (N_7805,N_548,N_2706);
or U7806 (N_7806,N_4543,N_394);
nand U7807 (N_7807,N_1701,N_2602);
nor U7808 (N_7808,N_4222,N_1064);
nand U7809 (N_7809,N_2062,N_3227);
xor U7810 (N_7810,N_1855,N_4437);
xor U7811 (N_7811,N_2740,N_2949);
and U7812 (N_7812,N_25,N_1722);
nor U7813 (N_7813,N_4913,N_2676);
xnor U7814 (N_7814,N_2259,N_3781);
or U7815 (N_7815,N_4537,N_3364);
and U7816 (N_7816,N_2911,N_2493);
nor U7817 (N_7817,N_795,N_4427);
nand U7818 (N_7818,N_687,N_4254);
xnor U7819 (N_7819,N_3315,N_4196);
nor U7820 (N_7820,N_4620,N_1047);
xor U7821 (N_7821,N_1219,N_1650);
or U7822 (N_7822,N_4066,N_2205);
or U7823 (N_7823,N_1018,N_3512);
nand U7824 (N_7824,N_4598,N_2886);
and U7825 (N_7825,N_2473,N_3197);
xor U7826 (N_7826,N_3033,N_1772);
nand U7827 (N_7827,N_2975,N_1782);
or U7828 (N_7828,N_2280,N_1161);
nand U7829 (N_7829,N_1584,N_979);
or U7830 (N_7830,N_4274,N_3925);
or U7831 (N_7831,N_1356,N_3268);
nand U7832 (N_7832,N_3085,N_1243);
nand U7833 (N_7833,N_230,N_3429);
xor U7834 (N_7834,N_2406,N_4939);
xnor U7835 (N_7835,N_2314,N_3374);
nor U7836 (N_7836,N_2248,N_1157);
nor U7837 (N_7837,N_4737,N_3629);
nor U7838 (N_7838,N_1510,N_669);
or U7839 (N_7839,N_1351,N_637);
xor U7840 (N_7840,N_1312,N_898);
xnor U7841 (N_7841,N_4578,N_4025);
nand U7842 (N_7842,N_3272,N_3921);
and U7843 (N_7843,N_324,N_2778);
nand U7844 (N_7844,N_2939,N_847);
xnor U7845 (N_7845,N_975,N_4731);
nand U7846 (N_7846,N_3730,N_4241);
and U7847 (N_7847,N_609,N_4102);
nor U7848 (N_7848,N_2504,N_1311);
and U7849 (N_7849,N_1402,N_4473);
xor U7850 (N_7850,N_1357,N_178);
or U7851 (N_7851,N_1909,N_2441);
xnor U7852 (N_7852,N_2845,N_1357);
and U7853 (N_7853,N_220,N_1245);
nand U7854 (N_7854,N_165,N_1050);
and U7855 (N_7855,N_526,N_551);
xor U7856 (N_7856,N_4953,N_411);
and U7857 (N_7857,N_3270,N_1985);
and U7858 (N_7858,N_942,N_396);
or U7859 (N_7859,N_443,N_2210);
or U7860 (N_7860,N_1711,N_2699);
or U7861 (N_7861,N_2230,N_792);
and U7862 (N_7862,N_783,N_3685);
and U7863 (N_7863,N_627,N_3442);
nor U7864 (N_7864,N_3109,N_2650);
nor U7865 (N_7865,N_3761,N_469);
xnor U7866 (N_7866,N_2437,N_2780);
and U7867 (N_7867,N_4520,N_2703);
or U7868 (N_7868,N_190,N_2060);
xnor U7869 (N_7869,N_3317,N_895);
and U7870 (N_7870,N_2868,N_2259);
and U7871 (N_7871,N_1348,N_4834);
xnor U7872 (N_7872,N_463,N_3582);
and U7873 (N_7873,N_942,N_2844);
nor U7874 (N_7874,N_501,N_4359);
and U7875 (N_7875,N_3007,N_3585);
xor U7876 (N_7876,N_3734,N_2873);
or U7877 (N_7877,N_2244,N_251);
nor U7878 (N_7878,N_2833,N_229);
nand U7879 (N_7879,N_3318,N_4465);
nand U7880 (N_7880,N_4984,N_1477);
nor U7881 (N_7881,N_2194,N_1073);
xnor U7882 (N_7882,N_2816,N_1331);
or U7883 (N_7883,N_3498,N_4927);
nand U7884 (N_7884,N_785,N_4437);
nor U7885 (N_7885,N_2960,N_235);
nand U7886 (N_7886,N_279,N_53);
and U7887 (N_7887,N_4592,N_2276);
xor U7888 (N_7888,N_1995,N_4933);
and U7889 (N_7889,N_1988,N_2343);
and U7890 (N_7890,N_500,N_804);
nor U7891 (N_7891,N_2039,N_4262);
xnor U7892 (N_7892,N_529,N_2869);
nand U7893 (N_7893,N_3411,N_1791);
nand U7894 (N_7894,N_1012,N_976);
nand U7895 (N_7895,N_1821,N_1933);
xor U7896 (N_7896,N_2290,N_1536);
xor U7897 (N_7897,N_1252,N_2320);
xnor U7898 (N_7898,N_505,N_4712);
or U7899 (N_7899,N_854,N_2064);
or U7900 (N_7900,N_2003,N_244);
nand U7901 (N_7901,N_1175,N_3412);
nand U7902 (N_7902,N_3589,N_1951);
or U7903 (N_7903,N_2487,N_235);
xor U7904 (N_7904,N_2839,N_4178);
nor U7905 (N_7905,N_1922,N_1127);
and U7906 (N_7906,N_2539,N_4635);
nand U7907 (N_7907,N_3352,N_241);
xnor U7908 (N_7908,N_2600,N_278);
or U7909 (N_7909,N_2445,N_1083);
nor U7910 (N_7910,N_4677,N_2310);
xor U7911 (N_7911,N_2036,N_2786);
or U7912 (N_7912,N_2557,N_1111);
nand U7913 (N_7913,N_4502,N_1375);
nand U7914 (N_7914,N_396,N_1984);
or U7915 (N_7915,N_4500,N_1223);
xnor U7916 (N_7916,N_4410,N_767);
and U7917 (N_7917,N_2776,N_81);
nor U7918 (N_7918,N_4103,N_2942);
nor U7919 (N_7919,N_1958,N_1450);
nor U7920 (N_7920,N_2660,N_2977);
and U7921 (N_7921,N_2331,N_3706);
xor U7922 (N_7922,N_505,N_1741);
xnor U7923 (N_7923,N_3167,N_676);
xnor U7924 (N_7924,N_4428,N_1781);
nand U7925 (N_7925,N_2693,N_1775);
and U7926 (N_7926,N_3327,N_1437);
xnor U7927 (N_7927,N_1288,N_2016);
and U7928 (N_7928,N_298,N_3367);
nand U7929 (N_7929,N_3123,N_2507);
xnor U7930 (N_7930,N_595,N_1880);
or U7931 (N_7931,N_4808,N_4342);
nand U7932 (N_7932,N_3352,N_2618);
nand U7933 (N_7933,N_2208,N_553);
nand U7934 (N_7934,N_1835,N_2784);
and U7935 (N_7935,N_3930,N_628);
nor U7936 (N_7936,N_1837,N_4496);
or U7937 (N_7937,N_2189,N_3302);
nand U7938 (N_7938,N_3232,N_972);
and U7939 (N_7939,N_2289,N_3251);
and U7940 (N_7940,N_1187,N_960);
or U7941 (N_7941,N_838,N_4200);
or U7942 (N_7942,N_4093,N_278);
or U7943 (N_7943,N_891,N_4255);
and U7944 (N_7944,N_1280,N_2901);
or U7945 (N_7945,N_222,N_3371);
nand U7946 (N_7946,N_2092,N_3000);
xnor U7947 (N_7947,N_2205,N_1047);
nand U7948 (N_7948,N_4717,N_2931);
nand U7949 (N_7949,N_3122,N_3771);
nand U7950 (N_7950,N_3382,N_2346);
nand U7951 (N_7951,N_3343,N_4668);
xor U7952 (N_7952,N_879,N_4294);
or U7953 (N_7953,N_1838,N_3067);
xor U7954 (N_7954,N_3394,N_638);
nand U7955 (N_7955,N_4110,N_681);
and U7956 (N_7956,N_2772,N_36);
or U7957 (N_7957,N_4500,N_387);
and U7958 (N_7958,N_3140,N_1840);
or U7959 (N_7959,N_3681,N_1319);
nand U7960 (N_7960,N_4417,N_23);
and U7961 (N_7961,N_3795,N_306);
nor U7962 (N_7962,N_618,N_2708);
and U7963 (N_7963,N_1132,N_4707);
nand U7964 (N_7964,N_4578,N_422);
nor U7965 (N_7965,N_3964,N_3346);
and U7966 (N_7966,N_665,N_973);
and U7967 (N_7967,N_3065,N_2199);
or U7968 (N_7968,N_741,N_122);
or U7969 (N_7969,N_2224,N_4475);
or U7970 (N_7970,N_946,N_217);
nand U7971 (N_7971,N_3930,N_4431);
xnor U7972 (N_7972,N_3192,N_2876);
nand U7973 (N_7973,N_240,N_49);
nor U7974 (N_7974,N_845,N_4775);
nor U7975 (N_7975,N_4172,N_2281);
or U7976 (N_7976,N_1072,N_4451);
or U7977 (N_7977,N_2645,N_1866);
xnor U7978 (N_7978,N_849,N_2565);
and U7979 (N_7979,N_690,N_847);
nand U7980 (N_7980,N_2806,N_894);
or U7981 (N_7981,N_2721,N_4202);
or U7982 (N_7982,N_4413,N_1203);
xor U7983 (N_7983,N_1373,N_181);
xnor U7984 (N_7984,N_4637,N_3146);
and U7985 (N_7985,N_2120,N_1278);
nand U7986 (N_7986,N_4873,N_2894);
nor U7987 (N_7987,N_2026,N_2522);
nor U7988 (N_7988,N_4790,N_2048);
nor U7989 (N_7989,N_4625,N_2409);
nand U7990 (N_7990,N_2897,N_2843);
and U7991 (N_7991,N_1276,N_3446);
and U7992 (N_7992,N_813,N_4248);
nand U7993 (N_7993,N_3949,N_480);
or U7994 (N_7994,N_756,N_722);
nor U7995 (N_7995,N_2404,N_1875);
xor U7996 (N_7996,N_33,N_4464);
and U7997 (N_7997,N_135,N_1964);
xnor U7998 (N_7998,N_4094,N_4702);
and U7999 (N_7999,N_1763,N_4958);
nor U8000 (N_8000,N_140,N_3616);
xor U8001 (N_8001,N_2799,N_2942);
or U8002 (N_8002,N_947,N_3088);
and U8003 (N_8003,N_1585,N_1312);
nand U8004 (N_8004,N_3429,N_2676);
nor U8005 (N_8005,N_1573,N_4679);
xnor U8006 (N_8006,N_3235,N_1786);
or U8007 (N_8007,N_2455,N_3392);
nor U8008 (N_8008,N_2199,N_424);
xor U8009 (N_8009,N_3927,N_4897);
nor U8010 (N_8010,N_2786,N_3087);
nor U8011 (N_8011,N_1156,N_1755);
nand U8012 (N_8012,N_3030,N_3174);
xnor U8013 (N_8013,N_3169,N_1531);
nor U8014 (N_8014,N_3072,N_2467);
xnor U8015 (N_8015,N_4497,N_4493);
nor U8016 (N_8016,N_3955,N_1409);
nor U8017 (N_8017,N_3779,N_1964);
nor U8018 (N_8018,N_2675,N_1404);
or U8019 (N_8019,N_4437,N_2327);
nand U8020 (N_8020,N_3957,N_4181);
or U8021 (N_8021,N_505,N_1191);
xor U8022 (N_8022,N_190,N_383);
and U8023 (N_8023,N_2325,N_1988);
or U8024 (N_8024,N_1268,N_1425);
and U8025 (N_8025,N_1045,N_2924);
or U8026 (N_8026,N_219,N_1200);
nand U8027 (N_8027,N_3384,N_1022);
and U8028 (N_8028,N_1199,N_1818);
nand U8029 (N_8029,N_4764,N_978);
or U8030 (N_8030,N_893,N_2946);
or U8031 (N_8031,N_3098,N_3558);
xnor U8032 (N_8032,N_2194,N_1455);
and U8033 (N_8033,N_3867,N_910);
or U8034 (N_8034,N_1640,N_1334);
nand U8035 (N_8035,N_4978,N_2705);
nor U8036 (N_8036,N_3465,N_759);
nor U8037 (N_8037,N_3490,N_1571);
nor U8038 (N_8038,N_2122,N_4475);
nand U8039 (N_8039,N_3389,N_1161);
or U8040 (N_8040,N_1057,N_2581);
and U8041 (N_8041,N_1110,N_612);
xnor U8042 (N_8042,N_2659,N_3936);
or U8043 (N_8043,N_3959,N_4800);
nor U8044 (N_8044,N_3818,N_2617);
nor U8045 (N_8045,N_376,N_3331);
nor U8046 (N_8046,N_2015,N_95);
nand U8047 (N_8047,N_458,N_4993);
nand U8048 (N_8048,N_4943,N_3240);
and U8049 (N_8049,N_4874,N_1781);
nand U8050 (N_8050,N_3974,N_1063);
and U8051 (N_8051,N_1681,N_1062);
nand U8052 (N_8052,N_3408,N_2046);
and U8053 (N_8053,N_791,N_2098);
and U8054 (N_8054,N_4136,N_989);
nand U8055 (N_8055,N_1149,N_4056);
or U8056 (N_8056,N_524,N_982);
nor U8057 (N_8057,N_3892,N_820);
nor U8058 (N_8058,N_2094,N_1741);
nor U8059 (N_8059,N_2663,N_3354);
or U8060 (N_8060,N_4923,N_3881);
and U8061 (N_8061,N_2205,N_165);
xnor U8062 (N_8062,N_1771,N_2426);
xor U8063 (N_8063,N_2795,N_2000);
nand U8064 (N_8064,N_2761,N_58);
nand U8065 (N_8065,N_3832,N_202);
nor U8066 (N_8066,N_956,N_4267);
xnor U8067 (N_8067,N_773,N_3791);
nor U8068 (N_8068,N_3544,N_4763);
xor U8069 (N_8069,N_2410,N_3357);
nor U8070 (N_8070,N_3894,N_1973);
xnor U8071 (N_8071,N_1647,N_206);
and U8072 (N_8072,N_3980,N_2021);
nand U8073 (N_8073,N_4983,N_227);
and U8074 (N_8074,N_4285,N_895);
or U8075 (N_8075,N_2641,N_362);
nand U8076 (N_8076,N_3098,N_3145);
nor U8077 (N_8077,N_2849,N_1825);
nand U8078 (N_8078,N_4771,N_1309);
nor U8079 (N_8079,N_171,N_444);
or U8080 (N_8080,N_2946,N_1841);
xnor U8081 (N_8081,N_2047,N_4880);
nand U8082 (N_8082,N_3355,N_848);
nor U8083 (N_8083,N_121,N_2787);
nand U8084 (N_8084,N_3783,N_4812);
xor U8085 (N_8085,N_2731,N_33);
xnor U8086 (N_8086,N_2595,N_999);
nand U8087 (N_8087,N_4693,N_3376);
or U8088 (N_8088,N_2096,N_1212);
xor U8089 (N_8089,N_1528,N_4686);
xor U8090 (N_8090,N_4056,N_4920);
nand U8091 (N_8091,N_4409,N_4446);
and U8092 (N_8092,N_1274,N_2395);
xor U8093 (N_8093,N_1705,N_2768);
or U8094 (N_8094,N_3291,N_997);
xnor U8095 (N_8095,N_769,N_1527);
and U8096 (N_8096,N_3893,N_166);
nand U8097 (N_8097,N_668,N_180);
or U8098 (N_8098,N_3506,N_1124);
nor U8099 (N_8099,N_3891,N_3869);
nor U8100 (N_8100,N_1108,N_2022);
or U8101 (N_8101,N_4567,N_3330);
nor U8102 (N_8102,N_940,N_3075);
nor U8103 (N_8103,N_1570,N_4925);
nand U8104 (N_8104,N_1718,N_1340);
or U8105 (N_8105,N_673,N_1652);
nor U8106 (N_8106,N_732,N_3547);
nand U8107 (N_8107,N_1214,N_321);
nand U8108 (N_8108,N_4820,N_3196);
or U8109 (N_8109,N_393,N_1822);
nor U8110 (N_8110,N_4502,N_4302);
nand U8111 (N_8111,N_2676,N_4294);
nor U8112 (N_8112,N_3515,N_4452);
nor U8113 (N_8113,N_3010,N_791);
nor U8114 (N_8114,N_1808,N_4792);
nor U8115 (N_8115,N_2541,N_89);
nand U8116 (N_8116,N_4713,N_4177);
xnor U8117 (N_8117,N_1007,N_2572);
or U8118 (N_8118,N_1967,N_159);
and U8119 (N_8119,N_2392,N_2322);
nand U8120 (N_8120,N_1850,N_3411);
or U8121 (N_8121,N_3717,N_663);
nor U8122 (N_8122,N_3319,N_1570);
xor U8123 (N_8123,N_863,N_4492);
or U8124 (N_8124,N_3350,N_3597);
or U8125 (N_8125,N_1798,N_1567);
xnor U8126 (N_8126,N_1857,N_4868);
or U8127 (N_8127,N_1860,N_4837);
and U8128 (N_8128,N_2495,N_770);
or U8129 (N_8129,N_2094,N_1557);
or U8130 (N_8130,N_3220,N_953);
or U8131 (N_8131,N_1293,N_3236);
and U8132 (N_8132,N_3680,N_4468);
nand U8133 (N_8133,N_2312,N_4913);
or U8134 (N_8134,N_1885,N_3256);
nor U8135 (N_8135,N_4656,N_2962);
nor U8136 (N_8136,N_1033,N_3886);
nor U8137 (N_8137,N_558,N_2285);
or U8138 (N_8138,N_1821,N_2847);
and U8139 (N_8139,N_1411,N_1254);
nand U8140 (N_8140,N_2370,N_3953);
nor U8141 (N_8141,N_3634,N_2974);
nor U8142 (N_8142,N_1280,N_3129);
or U8143 (N_8143,N_315,N_1714);
nor U8144 (N_8144,N_35,N_4452);
xnor U8145 (N_8145,N_3452,N_1136);
nor U8146 (N_8146,N_362,N_746);
xnor U8147 (N_8147,N_1098,N_3593);
xnor U8148 (N_8148,N_3656,N_3167);
nor U8149 (N_8149,N_333,N_1517);
nand U8150 (N_8150,N_4670,N_2591);
xnor U8151 (N_8151,N_3407,N_3987);
xnor U8152 (N_8152,N_3539,N_509);
nand U8153 (N_8153,N_103,N_442);
nor U8154 (N_8154,N_2925,N_2310);
or U8155 (N_8155,N_3182,N_4990);
nor U8156 (N_8156,N_4406,N_2724);
nor U8157 (N_8157,N_1632,N_803);
or U8158 (N_8158,N_845,N_747);
or U8159 (N_8159,N_199,N_135);
xnor U8160 (N_8160,N_4785,N_4583);
and U8161 (N_8161,N_3729,N_3777);
and U8162 (N_8162,N_1089,N_256);
nor U8163 (N_8163,N_1106,N_3384);
or U8164 (N_8164,N_3982,N_4437);
nand U8165 (N_8165,N_77,N_491);
nor U8166 (N_8166,N_1744,N_557);
and U8167 (N_8167,N_989,N_807);
xnor U8168 (N_8168,N_3095,N_1988);
nand U8169 (N_8169,N_803,N_2552);
xor U8170 (N_8170,N_2915,N_2847);
xnor U8171 (N_8171,N_3422,N_1919);
nor U8172 (N_8172,N_4481,N_4564);
and U8173 (N_8173,N_303,N_4467);
or U8174 (N_8174,N_953,N_1470);
nor U8175 (N_8175,N_1485,N_1698);
nor U8176 (N_8176,N_4180,N_954);
nor U8177 (N_8177,N_3615,N_3717);
or U8178 (N_8178,N_3918,N_1036);
and U8179 (N_8179,N_2670,N_151);
or U8180 (N_8180,N_3879,N_1218);
or U8181 (N_8181,N_1242,N_3876);
xor U8182 (N_8182,N_4725,N_2250);
xor U8183 (N_8183,N_3184,N_4121);
nand U8184 (N_8184,N_3728,N_819);
nor U8185 (N_8185,N_2278,N_3076);
and U8186 (N_8186,N_1274,N_3504);
and U8187 (N_8187,N_2545,N_2124);
xnor U8188 (N_8188,N_2625,N_1873);
and U8189 (N_8189,N_2910,N_3207);
and U8190 (N_8190,N_3540,N_1637);
nand U8191 (N_8191,N_1266,N_3800);
or U8192 (N_8192,N_2106,N_3952);
and U8193 (N_8193,N_2165,N_2272);
nand U8194 (N_8194,N_3929,N_3168);
nor U8195 (N_8195,N_2142,N_3275);
and U8196 (N_8196,N_3736,N_4093);
nand U8197 (N_8197,N_2431,N_1959);
and U8198 (N_8198,N_3213,N_798);
xnor U8199 (N_8199,N_861,N_1242);
nor U8200 (N_8200,N_2366,N_1927);
nand U8201 (N_8201,N_2754,N_1082);
xnor U8202 (N_8202,N_4480,N_3502);
nor U8203 (N_8203,N_3436,N_172);
xor U8204 (N_8204,N_4645,N_1578);
nand U8205 (N_8205,N_3885,N_3777);
xnor U8206 (N_8206,N_3942,N_2703);
and U8207 (N_8207,N_3681,N_417);
nor U8208 (N_8208,N_993,N_1825);
xnor U8209 (N_8209,N_2011,N_2360);
nor U8210 (N_8210,N_2052,N_2092);
and U8211 (N_8211,N_2379,N_2712);
and U8212 (N_8212,N_2232,N_416);
or U8213 (N_8213,N_1599,N_2671);
xnor U8214 (N_8214,N_4295,N_14);
nand U8215 (N_8215,N_1640,N_354);
nor U8216 (N_8216,N_2837,N_2247);
or U8217 (N_8217,N_4856,N_3733);
nor U8218 (N_8218,N_2458,N_430);
nand U8219 (N_8219,N_1084,N_885);
nand U8220 (N_8220,N_1410,N_637);
or U8221 (N_8221,N_4700,N_4983);
nand U8222 (N_8222,N_2609,N_903);
or U8223 (N_8223,N_2423,N_3710);
xor U8224 (N_8224,N_4281,N_1984);
xnor U8225 (N_8225,N_2945,N_4149);
or U8226 (N_8226,N_529,N_884);
or U8227 (N_8227,N_1362,N_1899);
nand U8228 (N_8228,N_1560,N_4827);
xor U8229 (N_8229,N_3636,N_3282);
and U8230 (N_8230,N_2530,N_2551);
nand U8231 (N_8231,N_4452,N_1226);
xor U8232 (N_8232,N_3359,N_3116);
and U8233 (N_8233,N_2269,N_2196);
xnor U8234 (N_8234,N_4113,N_4430);
or U8235 (N_8235,N_4967,N_1966);
nor U8236 (N_8236,N_1833,N_809);
nor U8237 (N_8237,N_1698,N_3322);
and U8238 (N_8238,N_1618,N_1607);
nand U8239 (N_8239,N_2250,N_4240);
and U8240 (N_8240,N_764,N_3194);
or U8241 (N_8241,N_1081,N_2688);
or U8242 (N_8242,N_943,N_1230);
xnor U8243 (N_8243,N_704,N_4592);
and U8244 (N_8244,N_1223,N_4242);
xor U8245 (N_8245,N_1499,N_228);
or U8246 (N_8246,N_3826,N_2813);
nand U8247 (N_8247,N_4238,N_912);
nand U8248 (N_8248,N_2800,N_3065);
or U8249 (N_8249,N_3862,N_4085);
nor U8250 (N_8250,N_4615,N_4467);
and U8251 (N_8251,N_3869,N_258);
nor U8252 (N_8252,N_4765,N_4516);
xor U8253 (N_8253,N_2916,N_4538);
and U8254 (N_8254,N_334,N_4392);
nand U8255 (N_8255,N_3289,N_4483);
nor U8256 (N_8256,N_2921,N_4819);
nor U8257 (N_8257,N_4482,N_3389);
or U8258 (N_8258,N_3991,N_3966);
nand U8259 (N_8259,N_3852,N_3315);
xor U8260 (N_8260,N_1465,N_1753);
nor U8261 (N_8261,N_4253,N_4464);
and U8262 (N_8262,N_3517,N_3528);
nor U8263 (N_8263,N_4829,N_4906);
nand U8264 (N_8264,N_886,N_3619);
xor U8265 (N_8265,N_2009,N_19);
nand U8266 (N_8266,N_4287,N_1114);
xor U8267 (N_8267,N_2319,N_1794);
or U8268 (N_8268,N_4516,N_4413);
xor U8269 (N_8269,N_256,N_3255);
nor U8270 (N_8270,N_2368,N_1796);
or U8271 (N_8271,N_552,N_34);
or U8272 (N_8272,N_373,N_91);
xor U8273 (N_8273,N_2267,N_4824);
nor U8274 (N_8274,N_1718,N_153);
or U8275 (N_8275,N_695,N_1581);
nor U8276 (N_8276,N_3192,N_2829);
nor U8277 (N_8277,N_4105,N_1604);
nor U8278 (N_8278,N_4490,N_2897);
nand U8279 (N_8279,N_834,N_2051);
xnor U8280 (N_8280,N_923,N_2051);
nor U8281 (N_8281,N_2427,N_3442);
or U8282 (N_8282,N_2895,N_168);
nand U8283 (N_8283,N_2460,N_3497);
and U8284 (N_8284,N_4645,N_20);
or U8285 (N_8285,N_3629,N_381);
nand U8286 (N_8286,N_3564,N_4083);
nor U8287 (N_8287,N_2497,N_1579);
nand U8288 (N_8288,N_2012,N_864);
or U8289 (N_8289,N_1204,N_2333);
nand U8290 (N_8290,N_114,N_4227);
xor U8291 (N_8291,N_4732,N_4983);
and U8292 (N_8292,N_2885,N_2472);
or U8293 (N_8293,N_3101,N_43);
or U8294 (N_8294,N_3906,N_2360);
nor U8295 (N_8295,N_3250,N_3057);
and U8296 (N_8296,N_1180,N_3406);
nor U8297 (N_8297,N_3622,N_4857);
nand U8298 (N_8298,N_1594,N_1698);
nand U8299 (N_8299,N_4103,N_2718);
nand U8300 (N_8300,N_2377,N_3202);
and U8301 (N_8301,N_364,N_910);
xnor U8302 (N_8302,N_1623,N_863);
nor U8303 (N_8303,N_2632,N_1052);
nor U8304 (N_8304,N_284,N_2936);
and U8305 (N_8305,N_3618,N_3670);
or U8306 (N_8306,N_1976,N_4217);
or U8307 (N_8307,N_135,N_2078);
nand U8308 (N_8308,N_2915,N_1176);
or U8309 (N_8309,N_1490,N_4432);
xor U8310 (N_8310,N_371,N_3858);
nor U8311 (N_8311,N_2026,N_4831);
nand U8312 (N_8312,N_1518,N_1306);
and U8313 (N_8313,N_2398,N_878);
or U8314 (N_8314,N_3367,N_583);
nand U8315 (N_8315,N_3862,N_3585);
nand U8316 (N_8316,N_4019,N_36);
or U8317 (N_8317,N_4934,N_2773);
xnor U8318 (N_8318,N_4120,N_1191);
nor U8319 (N_8319,N_2671,N_4797);
nor U8320 (N_8320,N_2328,N_1620);
nand U8321 (N_8321,N_751,N_4250);
and U8322 (N_8322,N_986,N_1975);
nand U8323 (N_8323,N_2648,N_4808);
nand U8324 (N_8324,N_2104,N_929);
and U8325 (N_8325,N_4851,N_2494);
and U8326 (N_8326,N_4319,N_1419);
nor U8327 (N_8327,N_1762,N_4415);
xnor U8328 (N_8328,N_145,N_1044);
xnor U8329 (N_8329,N_4416,N_1609);
and U8330 (N_8330,N_4508,N_425);
nor U8331 (N_8331,N_3959,N_2519);
xor U8332 (N_8332,N_61,N_1350);
nor U8333 (N_8333,N_458,N_3915);
nand U8334 (N_8334,N_1923,N_1981);
and U8335 (N_8335,N_1791,N_3814);
nand U8336 (N_8336,N_365,N_2972);
or U8337 (N_8337,N_1835,N_1062);
and U8338 (N_8338,N_930,N_463);
and U8339 (N_8339,N_3600,N_2109);
and U8340 (N_8340,N_3776,N_1575);
and U8341 (N_8341,N_580,N_3615);
or U8342 (N_8342,N_3910,N_2496);
and U8343 (N_8343,N_1560,N_2054);
xor U8344 (N_8344,N_2644,N_164);
nor U8345 (N_8345,N_2888,N_1767);
or U8346 (N_8346,N_4571,N_4564);
nand U8347 (N_8347,N_1632,N_2556);
nand U8348 (N_8348,N_1001,N_4398);
and U8349 (N_8349,N_2112,N_3468);
nor U8350 (N_8350,N_1116,N_538);
xor U8351 (N_8351,N_4260,N_3727);
xnor U8352 (N_8352,N_3656,N_243);
nand U8353 (N_8353,N_2879,N_2888);
xor U8354 (N_8354,N_2186,N_1338);
and U8355 (N_8355,N_4547,N_3814);
nor U8356 (N_8356,N_515,N_3600);
nand U8357 (N_8357,N_3635,N_2280);
nand U8358 (N_8358,N_76,N_4176);
xnor U8359 (N_8359,N_3051,N_1228);
or U8360 (N_8360,N_348,N_216);
nand U8361 (N_8361,N_3823,N_4909);
and U8362 (N_8362,N_3416,N_1294);
xor U8363 (N_8363,N_2487,N_4758);
and U8364 (N_8364,N_4938,N_2930);
and U8365 (N_8365,N_1283,N_4772);
xor U8366 (N_8366,N_4306,N_3872);
nand U8367 (N_8367,N_2635,N_2141);
and U8368 (N_8368,N_1840,N_4341);
nand U8369 (N_8369,N_2754,N_3555);
nor U8370 (N_8370,N_2242,N_3156);
nor U8371 (N_8371,N_277,N_2327);
nand U8372 (N_8372,N_671,N_2989);
and U8373 (N_8373,N_1841,N_1967);
nor U8374 (N_8374,N_32,N_547);
or U8375 (N_8375,N_2689,N_2449);
nand U8376 (N_8376,N_2054,N_1047);
and U8377 (N_8377,N_4177,N_1258);
and U8378 (N_8378,N_4276,N_2507);
xor U8379 (N_8379,N_2108,N_605);
and U8380 (N_8380,N_2073,N_2402);
and U8381 (N_8381,N_4809,N_1095);
nor U8382 (N_8382,N_2172,N_3624);
or U8383 (N_8383,N_567,N_3563);
or U8384 (N_8384,N_225,N_2126);
nand U8385 (N_8385,N_4034,N_3261);
nand U8386 (N_8386,N_1836,N_777);
nand U8387 (N_8387,N_1345,N_715);
or U8388 (N_8388,N_3567,N_4164);
and U8389 (N_8389,N_4723,N_2438);
xor U8390 (N_8390,N_3003,N_3045);
and U8391 (N_8391,N_209,N_4105);
and U8392 (N_8392,N_370,N_4258);
nor U8393 (N_8393,N_3085,N_3366);
or U8394 (N_8394,N_2396,N_104);
or U8395 (N_8395,N_50,N_1256);
nand U8396 (N_8396,N_377,N_4107);
nand U8397 (N_8397,N_1732,N_4267);
xnor U8398 (N_8398,N_2468,N_1049);
and U8399 (N_8399,N_1688,N_245);
and U8400 (N_8400,N_755,N_3230);
nand U8401 (N_8401,N_2049,N_81);
and U8402 (N_8402,N_24,N_1627);
xor U8403 (N_8403,N_3801,N_4955);
nor U8404 (N_8404,N_1184,N_3358);
nor U8405 (N_8405,N_3153,N_3724);
or U8406 (N_8406,N_2974,N_715);
nand U8407 (N_8407,N_2813,N_1999);
xnor U8408 (N_8408,N_2809,N_243);
nand U8409 (N_8409,N_2916,N_3504);
xnor U8410 (N_8410,N_1944,N_827);
or U8411 (N_8411,N_1346,N_4617);
xnor U8412 (N_8412,N_2687,N_2465);
xor U8413 (N_8413,N_3995,N_4869);
nand U8414 (N_8414,N_2030,N_4608);
nor U8415 (N_8415,N_3347,N_1258);
and U8416 (N_8416,N_1656,N_4307);
nand U8417 (N_8417,N_3117,N_2520);
xor U8418 (N_8418,N_1205,N_241);
and U8419 (N_8419,N_3886,N_423);
xor U8420 (N_8420,N_439,N_1951);
nor U8421 (N_8421,N_4908,N_1848);
nor U8422 (N_8422,N_2797,N_1784);
xnor U8423 (N_8423,N_2041,N_3453);
and U8424 (N_8424,N_659,N_3684);
xor U8425 (N_8425,N_1977,N_4884);
and U8426 (N_8426,N_2732,N_1986);
or U8427 (N_8427,N_1944,N_1570);
or U8428 (N_8428,N_4425,N_4486);
xor U8429 (N_8429,N_3476,N_3555);
and U8430 (N_8430,N_465,N_3167);
and U8431 (N_8431,N_1442,N_328);
and U8432 (N_8432,N_4069,N_4193);
and U8433 (N_8433,N_2132,N_2751);
or U8434 (N_8434,N_373,N_529);
nand U8435 (N_8435,N_3591,N_4531);
nor U8436 (N_8436,N_3,N_987);
xnor U8437 (N_8437,N_1594,N_3273);
nand U8438 (N_8438,N_2117,N_777);
xor U8439 (N_8439,N_25,N_1547);
nand U8440 (N_8440,N_287,N_2304);
and U8441 (N_8441,N_4575,N_2813);
and U8442 (N_8442,N_725,N_3485);
or U8443 (N_8443,N_1443,N_2920);
nand U8444 (N_8444,N_4642,N_2835);
or U8445 (N_8445,N_4190,N_1939);
xor U8446 (N_8446,N_1551,N_1670);
nand U8447 (N_8447,N_3630,N_4439);
or U8448 (N_8448,N_2896,N_1324);
or U8449 (N_8449,N_2603,N_2810);
nand U8450 (N_8450,N_397,N_3736);
or U8451 (N_8451,N_2525,N_4454);
xnor U8452 (N_8452,N_307,N_2720);
or U8453 (N_8453,N_1413,N_4558);
or U8454 (N_8454,N_3527,N_167);
xnor U8455 (N_8455,N_2358,N_767);
or U8456 (N_8456,N_4417,N_2907);
nand U8457 (N_8457,N_732,N_2302);
nor U8458 (N_8458,N_1333,N_2468);
nor U8459 (N_8459,N_3216,N_4857);
nand U8460 (N_8460,N_1400,N_4483);
and U8461 (N_8461,N_175,N_867);
nand U8462 (N_8462,N_1017,N_3535);
nor U8463 (N_8463,N_4169,N_4566);
and U8464 (N_8464,N_4705,N_1952);
or U8465 (N_8465,N_3016,N_4591);
nand U8466 (N_8466,N_2982,N_3653);
nor U8467 (N_8467,N_4944,N_4207);
nand U8468 (N_8468,N_320,N_2502);
nand U8469 (N_8469,N_3933,N_3479);
or U8470 (N_8470,N_4103,N_4765);
xor U8471 (N_8471,N_2159,N_1903);
xor U8472 (N_8472,N_4705,N_94);
xor U8473 (N_8473,N_4243,N_3767);
xor U8474 (N_8474,N_2748,N_4615);
nand U8475 (N_8475,N_2304,N_448);
or U8476 (N_8476,N_3538,N_44);
nor U8477 (N_8477,N_2142,N_1379);
and U8478 (N_8478,N_1494,N_1562);
nor U8479 (N_8479,N_4756,N_968);
xnor U8480 (N_8480,N_1175,N_108);
nand U8481 (N_8481,N_4173,N_627);
nand U8482 (N_8482,N_1379,N_4719);
xor U8483 (N_8483,N_2766,N_4629);
nor U8484 (N_8484,N_4753,N_1739);
nor U8485 (N_8485,N_2036,N_4255);
xor U8486 (N_8486,N_2771,N_3861);
and U8487 (N_8487,N_2688,N_4884);
xnor U8488 (N_8488,N_2684,N_3382);
or U8489 (N_8489,N_4042,N_639);
nand U8490 (N_8490,N_213,N_2999);
nor U8491 (N_8491,N_3266,N_2678);
nor U8492 (N_8492,N_4935,N_2945);
or U8493 (N_8493,N_3570,N_1122);
xnor U8494 (N_8494,N_3468,N_3988);
xor U8495 (N_8495,N_2500,N_3000);
xnor U8496 (N_8496,N_2527,N_1412);
and U8497 (N_8497,N_1336,N_3588);
xor U8498 (N_8498,N_859,N_4669);
or U8499 (N_8499,N_3512,N_813);
nand U8500 (N_8500,N_1327,N_3140);
and U8501 (N_8501,N_570,N_4875);
xnor U8502 (N_8502,N_484,N_4088);
or U8503 (N_8503,N_76,N_318);
nand U8504 (N_8504,N_3620,N_4298);
or U8505 (N_8505,N_3689,N_4602);
and U8506 (N_8506,N_4923,N_4111);
or U8507 (N_8507,N_4767,N_4215);
nand U8508 (N_8508,N_4447,N_961);
or U8509 (N_8509,N_3464,N_4549);
nand U8510 (N_8510,N_350,N_1323);
nor U8511 (N_8511,N_2216,N_4345);
and U8512 (N_8512,N_3724,N_2070);
xor U8513 (N_8513,N_1374,N_2688);
nand U8514 (N_8514,N_1915,N_1266);
nand U8515 (N_8515,N_3803,N_1581);
xor U8516 (N_8516,N_3997,N_2678);
nor U8517 (N_8517,N_3326,N_2485);
nor U8518 (N_8518,N_4494,N_2214);
nor U8519 (N_8519,N_2451,N_666);
xnor U8520 (N_8520,N_4423,N_4315);
and U8521 (N_8521,N_381,N_242);
nand U8522 (N_8522,N_3757,N_2970);
xor U8523 (N_8523,N_82,N_4890);
and U8524 (N_8524,N_715,N_1687);
or U8525 (N_8525,N_1150,N_3704);
or U8526 (N_8526,N_1757,N_2855);
and U8527 (N_8527,N_4876,N_3871);
nand U8528 (N_8528,N_3679,N_3823);
or U8529 (N_8529,N_4383,N_3691);
nor U8530 (N_8530,N_2143,N_44);
or U8531 (N_8531,N_909,N_1207);
and U8532 (N_8532,N_443,N_4938);
nor U8533 (N_8533,N_107,N_640);
xor U8534 (N_8534,N_2761,N_2080);
nand U8535 (N_8535,N_4995,N_4312);
nand U8536 (N_8536,N_2725,N_1647);
nor U8537 (N_8537,N_271,N_1923);
or U8538 (N_8538,N_946,N_3593);
xnor U8539 (N_8539,N_1967,N_1310);
or U8540 (N_8540,N_3307,N_2232);
xor U8541 (N_8541,N_113,N_3062);
xor U8542 (N_8542,N_1979,N_3173);
nor U8543 (N_8543,N_435,N_3964);
or U8544 (N_8544,N_2813,N_2994);
and U8545 (N_8545,N_408,N_4662);
and U8546 (N_8546,N_1600,N_4086);
xnor U8547 (N_8547,N_3745,N_2779);
and U8548 (N_8548,N_569,N_1287);
or U8549 (N_8549,N_337,N_1019);
and U8550 (N_8550,N_4661,N_1032);
nor U8551 (N_8551,N_3574,N_236);
xor U8552 (N_8552,N_787,N_4877);
nor U8553 (N_8553,N_3112,N_763);
and U8554 (N_8554,N_3925,N_1709);
nor U8555 (N_8555,N_1113,N_4216);
nor U8556 (N_8556,N_4604,N_3740);
xnor U8557 (N_8557,N_4623,N_950);
or U8558 (N_8558,N_2078,N_1394);
nand U8559 (N_8559,N_895,N_50);
or U8560 (N_8560,N_4483,N_2564);
nor U8561 (N_8561,N_3422,N_3553);
or U8562 (N_8562,N_2666,N_4557);
xor U8563 (N_8563,N_3259,N_3250);
or U8564 (N_8564,N_211,N_3066);
and U8565 (N_8565,N_4415,N_1830);
nand U8566 (N_8566,N_376,N_1428);
nand U8567 (N_8567,N_794,N_3979);
nand U8568 (N_8568,N_2597,N_4328);
nor U8569 (N_8569,N_3803,N_2903);
nand U8570 (N_8570,N_3673,N_2517);
and U8571 (N_8571,N_272,N_4342);
and U8572 (N_8572,N_2490,N_821);
or U8573 (N_8573,N_1167,N_1877);
nand U8574 (N_8574,N_2542,N_4522);
or U8575 (N_8575,N_1510,N_1352);
nand U8576 (N_8576,N_3439,N_3533);
nand U8577 (N_8577,N_1432,N_733);
xor U8578 (N_8578,N_4667,N_4818);
nand U8579 (N_8579,N_1897,N_1673);
nand U8580 (N_8580,N_619,N_1010);
nor U8581 (N_8581,N_3641,N_997);
nand U8582 (N_8582,N_3826,N_1536);
xor U8583 (N_8583,N_2644,N_2889);
xor U8584 (N_8584,N_1533,N_4445);
nor U8585 (N_8585,N_4679,N_4613);
xnor U8586 (N_8586,N_4885,N_4037);
and U8587 (N_8587,N_1198,N_202);
nand U8588 (N_8588,N_4585,N_2550);
nor U8589 (N_8589,N_2001,N_352);
nand U8590 (N_8590,N_2022,N_1965);
nand U8591 (N_8591,N_3260,N_3313);
nand U8592 (N_8592,N_1426,N_2036);
nor U8593 (N_8593,N_2721,N_3045);
or U8594 (N_8594,N_2601,N_2622);
and U8595 (N_8595,N_2674,N_701);
nor U8596 (N_8596,N_2365,N_4303);
nor U8597 (N_8597,N_2358,N_2390);
xnor U8598 (N_8598,N_827,N_2048);
xor U8599 (N_8599,N_4587,N_772);
or U8600 (N_8600,N_4104,N_967);
nor U8601 (N_8601,N_3669,N_4898);
xor U8602 (N_8602,N_3040,N_3583);
or U8603 (N_8603,N_2318,N_2639);
or U8604 (N_8604,N_3628,N_2455);
nor U8605 (N_8605,N_2985,N_2419);
and U8606 (N_8606,N_260,N_2928);
nor U8607 (N_8607,N_833,N_3613);
nor U8608 (N_8608,N_1440,N_1029);
nand U8609 (N_8609,N_2432,N_3462);
or U8610 (N_8610,N_2185,N_780);
or U8611 (N_8611,N_1593,N_1021);
or U8612 (N_8612,N_4735,N_4363);
nand U8613 (N_8613,N_1423,N_499);
nor U8614 (N_8614,N_3391,N_2458);
nor U8615 (N_8615,N_1636,N_1994);
xor U8616 (N_8616,N_377,N_606);
nor U8617 (N_8617,N_1976,N_2646);
nor U8618 (N_8618,N_426,N_2201);
nor U8619 (N_8619,N_1130,N_4404);
nand U8620 (N_8620,N_2101,N_1246);
nor U8621 (N_8621,N_4758,N_1027);
xor U8622 (N_8622,N_3955,N_3122);
nor U8623 (N_8623,N_3608,N_3918);
or U8624 (N_8624,N_3486,N_410);
nand U8625 (N_8625,N_3766,N_1406);
xor U8626 (N_8626,N_3165,N_4533);
nor U8627 (N_8627,N_2679,N_714);
xnor U8628 (N_8628,N_758,N_4066);
or U8629 (N_8629,N_324,N_2113);
nand U8630 (N_8630,N_3635,N_1549);
nand U8631 (N_8631,N_4150,N_1512);
nand U8632 (N_8632,N_3958,N_2294);
or U8633 (N_8633,N_37,N_1622);
or U8634 (N_8634,N_4960,N_3751);
nand U8635 (N_8635,N_400,N_2442);
or U8636 (N_8636,N_4090,N_1031);
nor U8637 (N_8637,N_4247,N_1864);
xor U8638 (N_8638,N_4655,N_3209);
nand U8639 (N_8639,N_2144,N_214);
nor U8640 (N_8640,N_4510,N_1328);
nor U8641 (N_8641,N_3946,N_4441);
xnor U8642 (N_8642,N_4117,N_1151);
nor U8643 (N_8643,N_4711,N_3715);
nand U8644 (N_8644,N_71,N_1553);
xor U8645 (N_8645,N_721,N_2762);
nor U8646 (N_8646,N_2596,N_119);
xor U8647 (N_8647,N_3579,N_65);
xor U8648 (N_8648,N_2269,N_85);
xnor U8649 (N_8649,N_3556,N_168);
and U8650 (N_8650,N_3977,N_3193);
nand U8651 (N_8651,N_2345,N_1679);
nor U8652 (N_8652,N_2493,N_1211);
and U8653 (N_8653,N_4291,N_1550);
nor U8654 (N_8654,N_4866,N_3563);
nand U8655 (N_8655,N_3674,N_2194);
nand U8656 (N_8656,N_3206,N_3224);
nor U8657 (N_8657,N_2651,N_816);
nand U8658 (N_8658,N_829,N_3649);
xnor U8659 (N_8659,N_4601,N_2162);
xnor U8660 (N_8660,N_3523,N_1348);
nor U8661 (N_8661,N_1539,N_1954);
xnor U8662 (N_8662,N_4684,N_4979);
xnor U8663 (N_8663,N_4453,N_3122);
nand U8664 (N_8664,N_3079,N_4472);
xnor U8665 (N_8665,N_2278,N_3565);
nand U8666 (N_8666,N_403,N_1126);
and U8667 (N_8667,N_4610,N_846);
and U8668 (N_8668,N_2480,N_422);
nand U8669 (N_8669,N_1067,N_551);
xor U8670 (N_8670,N_4186,N_3613);
nand U8671 (N_8671,N_4591,N_998);
nand U8672 (N_8672,N_4504,N_1646);
and U8673 (N_8673,N_2770,N_4263);
xnor U8674 (N_8674,N_4815,N_1923);
xnor U8675 (N_8675,N_4781,N_688);
and U8676 (N_8676,N_964,N_1241);
xnor U8677 (N_8677,N_1686,N_2927);
and U8678 (N_8678,N_3710,N_3180);
or U8679 (N_8679,N_3610,N_2352);
and U8680 (N_8680,N_3206,N_4301);
nand U8681 (N_8681,N_4308,N_2975);
nand U8682 (N_8682,N_713,N_888);
nor U8683 (N_8683,N_3549,N_2616);
and U8684 (N_8684,N_972,N_3791);
nor U8685 (N_8685,N_463,N_2025);
and U8686 (N_8686,N_39,N_763);
or U8687 (N_8687,N_3766,N_589);
nor U8688 (N_8688,N_1805,N_2792);
xor U8689 (N_8689,N_2728,N_4157);
nand U8690 (N_8690,N_2920,N_350);
or U8691 (N_8691,N_2600,N_2865);
nand U8692 (N_8692,N_4085,N_4363);
nor U8693 (N_8693,N_4835,N_2814);
xor U8694 (N_8694,N_4318,N_4041);
nor U8695 (N_8695,N_371,N_576);
nand U8696 (N_8696,N_10,N_407);
nor U8697 (N_8697,N_4438,N_3172);
nand U8698 (N_8698,N_2327,N_3806);
nand U8699 (N_8699,N_4910,N_1115);
nor U8700 (N_8700,N_1600,N_3559);
or U8701 (N_8701,N_4524,N_2390);
nand U8702 (N_8702,N_2481,N_2916);
nand U8703 (N_8703,N_317,N_1208);
and U8704 (N_8704,N_2618,N_3342);
nor U8705 (N_8705,N_4626,N_2118);
nor U8706 (N_8706,N_1890,N_3041);
or U8707 (N_8707,N_486,N_4477);
nor U8708 (N_8708,N_853,N_724);
and U8709 (N_8709,N_4707,N_1182);
xor U8710 (N_8710,N_2275,N_4765);
and U8711 (N_8711,N_2041,N_1523);
and U8712 (N_8712,N_1460,N_167);
and U8713 (N_8713,N_3257,N_1358);
and U8714 (N_8714,N_4839,N_3643);
nor U8715 (N_8715,N_3568,N_2822);
nand U8716 (N_8716,N_1648,N_357);
or U8717 (N_8717,N_4753,N_2448);
xor U8718 (N_8718,N_3903,N_2022);
or U8719 (N_8719,N_769,N_81);
and U8720 (N_8720,N_3766,N_3201);
or U8721 (N_8721,N_987,N_1592);
or U8722 (N_8722,N_3191,N_4692);
nand U8723 (N_8723,N_729,N_2819);
or U8724 (N_8724,N_959,N_2449);
and U8725 (N_8725,N_2156,N_3499);
nor U8726 (N_8726,N_1939,N_4381);
nand U8727 (N_8727,N_2483,N_4130);
and U8728 (N_8728,N_3445,N_2799);
xor U8729 (N_8729,N_2376,N_4785);
and U8730 (N_8730,N_2850,N_2);
nor U8731 (N_8731,N_3841,N_4900);
or U8732 (N_8732,N_3000,N_3985);
or U8733 (N_8733,N_3314,N_2154);
nor U8734 (N_8734,N_3466,N_4452);
xor U8735 (N_8735,N_1009,N_224);
or U8736 (N_8736,N_2576,N_1070);
or U8737 (N_8737,N_3218,N_2797);
nand U8738 (N_8738,N_4139,N_3014);
nand U8739 (N_8739,N_4779,N_782);
xnor U8740 (N_8740,N_233,N_3590);
nor U8741 (N_8741,N_299,N_4231);
or U8742 (N_8742,N_4500,N_4781);
xnor U8743 (N_8743,N_1589,N_4410);
nand U8744 (N_8744,N_3382,N_3618);
nor U8745 (N_8745,N_3245,N_3479);
nor U8746 (N_8746,N_2219,N_23);
or U8747 (N_8747,N_1377,N_1016);
nor U8748 (N_8748,N_3151,N_25);
xnor U8749 (N_8749,N_1763,N_3651);
and U8750 (N_8750,N_3323,N_2869);
and U8751 (N_8751,N_1275,N_2386);
xnor U8752 (N_8752,N_1964,N_4850);
and U8753 (N_8753,N_3104,N_3590);
xor U8754 (N_8754,N_48,N_4747);
nand U8755 (N_8755,N_2408,N_1196);
nor U8756 (N_8756,N_2935,N_2410);
nand U8757 (N_8757,N_2413,N_4781);
and U8758 (N_8758,N_1343,N_4040);
or U8759 (N_8759,N_1748,N_2870);
xnor U8760 (N_8760,N_2808,N_3513);
xnor U8761 (N_8761,N_1147,N_2876);
nor U8762 (N_8762,N_3062,N_3945);
or U8763 (N_8763,N_4101,N_3815);
xor U8764 (N_8764,N_4749,N_4938);
and U8765 (N_8765,N_3927,N_2634);
or U8766 (N_8766,N_4556,N_2865);
and U8767 (N_8767,N_3952,N_1378);
nand U8768 (N_8768,N_3105,N_2495);
xor U8769 (N_8769,N_3353,N_3693);
nor U8770 (N_8770,N_2618,N_4527);
xor U8771 (N_8771,N_2670,N_4317);
or U8772 (N_8772,N_2555,N_1785);
nor U8773 (N_8773,N_2912,N_2606);
or U8774 (N_8774,N_2783,N_3685);
xor U8775 (N_8775,N_4694,N_1659);
nand U8776 (N_8776,N_3032,N_2837);
xnor U8777 (N_8777,N_4152,N_1110);
nor U8778 (N_8778,N_1867,N_1745);
or U8779 (N_8779,N_1961,N_3331);
xor U8780 (N_8780,N_4939,N_4853);
and U8781 (N_8781,N_638,N_1198);
and U8782 (N_8782,N_2713,N_750);
or U8783 (N_8783,N_311,N_29);
and U8784 (N_8784,N_3383,N_175);
and U8785 (N_8785,N_72,N_850);
or U8786 (N_8786,N_4658,N_431);
or U8787 (N_8787,N_3421,N_3790);
xor U8788 (N_8788,N_3684,N_3620);
or U8789 (N_8789,N_4170,N_2273);
xnor U8790 (N_8790,N_4538,N_184);
xor U8791 (N_8791,N_2657,N_1574);
or U8792 (N_8792,N_4915,N_3566);
and U8793 (N_8793,N_1746,N_398);
nor U8794 (N_8794,N_4309,N_2433);
and U8795 (N_8795,N_2119,N_763);
nand U8796 (N_8796,N_186,N_1183);
nor U8797 (N_8797,N_4358,N_1781);
and U8798 (N_8798,N_3139,N_1548);
nand U8799 (N_8799,N_2933,N_900);
xnor U8800 (N_8800,N_224,N_4356);
xor U8801 (N_8801,N_955,N_3530);
nand U8802 (N_8802,N_3184,N_2574);
or U8803 (N_8803,N_3042,N_3146);
xor U8804 (N_8804,N_288,N_4692);
and U8805 (N_8805,N_3366,N_4637);
nand U8806 (N_8806,N_3977,N_1113);
and U8807 (N_8807,N_4176,N_4182);
or U8808 (N_8808,N_1968,N_1612);
nand U8809 (N_8809,N_4261,N_2395);
and U8810 (N_8810,N_3529,N_2097);
nand U8811 (N_8811,N_3904,N_2045);
or U8812 (N_8812,N_1209,N_1645);
xnor U8813 (N_8813,N_2374,N_2406);
xnor U8814 (N_8814,N_72,N_1120);
or U8815 (N_8815,N_3071,N_3707);
xor U8816 (N_8816,N_1383,N_126);
xnor U8817 (N_8817,N_1315,N_3652);
or U8818 (N_8818,N_4036,N_4847);
and U8819 (N_8819,N_3378,N_3031);
nand U8820 (N_8820,N_338,N_4795);
nor U8821 (N_8821,N_3580,N_2239);
xnor U8822 (N_8822,N_1586,N_463);
xnor U8823 (N_8823,N_324,N_3791);
or U8824 (N_8824,N_578,N_2700);
nand U8825 (N_8825,N_4411,N_3521);
or U8826 (N_8826,N_3429,N_1658);
nand U8827 (N_8827,N_3707,N_1709);
xnor U8828 (N_8828,N_1879,N_950);
nor U8829 (N_8829,N_313,N_3089);
and U8830 (N_8830,N_2060,N_3624);
nand U8831 (N_8831,N_1212,N_2187);
and U8832 (N_8832,N_1252,N_1493);
xnor U8833 (N_8833,N_716,N_3633);
xor U8834 (N_8834,N_822,N_848);
or U8835 (N_8835,N_111,N_761);
nand U8836 (N_8836,N_1931,N_274);
or U8837 (N_8837,N_3370,N_3829);
or U8838 (N_8838,N_4398,N_270);
xor U8839 (N_8839,N_3692,N_4886);
and U8840 (N_8840,N_3461,N_4688);
nand U8841 (N_8841,N_4170,N_2385);
xor U8842 (N_8842,N_2069,N_1136);
nand U8843 (N_8843,N_1674,N_583);
or U8844 (N_8844,N_892,N_45);
and U8845 (N_8845,N_4134,N_1503);
nand U8846 (N_8846,N_4596,N_1735);
or U8847 (N_8847,N_277,N_628);
or U8848 (N_8848,N_1474,N_2967);
nand U8849 (N_8849,N_3497,N_4545);
or U8850 (N_8850,N_280,N_3780);
nand U8851 (N_8851,N_3433,N_1338);
or U8852 (N_8852,N_2415,N_1445);
xor U8853 (N_8853,N_3242,N_2001);
nand U8854 (N_8854,N_449,N_4449);
or U8855 (N_8855,N_488,N_2573);
or U8856 (N_8856,N_854,N_2442);
or U8857 (N_8857,N_3387,N_2837);
and U8858 (N_8858,N_2541,N_3638);
or U8859 (N_8859,N_3801,N_2109);
and U8860 (N_8860,N_1482,N_4852);
nand U8861 (N_8861,N_3673,N_100);
or U8862 (N_8862,N_2393,N_4928);
nor U8863 (N_8863,N_982,N_3899);
nor U8864 (N_8864,N_3386,N_3833);
xor U8865 (N_8865,N_2671,N_2724);
or U8866 (N_8866,N_391,N_207);
xor U8867 (N_8867,N_484,N_3228);
nor U8868 (N_8868,N_914,N_2691);
or U8869 (N_8869,N_3767,N_242);
nand U8870 (N_8870,N_1581,N_55);
and U8871 (N_8871,N_4487,N_4809);
xnor U8872 (N_8872,N_1438,N_4279);
xnor U8873 (N_8873,N_519,N_1131);
and U8874 (N_8874,N_3941,N_393);
or U8875 (N_8875,N_1688,N_3581);
nand U8876 (N_8876,N_4459,N_2630);
nand U8877 (N_8877,N_4323,N_3487);
and U8878 (N_8878,N_1692,N_14);
or U8879 (N_8879,N_3586,N_4740);
or U8880 (N_8880,N_1676,N_2504);
or U8881 (N_8881,N_4314,N_2278);
nor U8882 (N_8882,N_2173,N_519);
nor U8883 (N_8883,N_1609,N_2769);
nand U8884 (N_8884,N_3364,N_3730);
nor U8885 (N_8885,N_1092,N_1256);
xor U8886 (N_8886,N_980,N_410);
and U8887 (N_8887,N_758,N_3877);
nor U8888 (N_8888,N_4745,N_2449);
nand U8889 (N_8889,N_4572,N_32);
or U8890 (N_8890,N_3761,N_1333);
and U8891 (N_8891,N_4253,N_2975);
or U8892 (N_8892,N_4923,N_1070);
xor U8893 (N_8893,N_498,N_3236);
or U8894 (N_8894,N_2553,N_1887);
nand U8895 (N_8895,N_4442,N_2869);
nor U8896 (N_8896,N_4964,N_545);
nand U8897 (N_8897,N_554,N_1138);
and U8898 (N_8898,N_10,N_4714);
or U8899 (N_8899,N_3744,N_2574);
nand U8900 (N_8900,N_4285,N_3417);
nor U8901 (N_8901,N_2412,N_853);
nand U8902 (N_8902,N_4046,N_210);
nand U8903 (N_8903,N_1460,N_1935);
and U8904 (N_8904,N_4338,N_1230);
and U8905 (N_8905,N_4346,N_1829);
xor U8906 (N_8906,N_394,N_675);
nor U8907 (N_8907,N_515,N_0);
nand U8908 (N_8908,N_1192,N_127);
nand U8909 (N_8909,N_3467,N_546);
xnor U8910 (N_8910,N_3514,N_3658);
nor U8911 (N_8911,N_1189,N_3593);
xnor U8912 (N_8912,N_4133,N_278);
nor U8913 (N_8913,N_3524,N_1897);
or U8914 (N_8914,N_4364,N_2550);
nand U8915 (N_8915,N_3666,N_1403);
nand U8916 (N_8916,N_1525,N_1691);
and U8917 (N_8917,N_2460,N_4403);
nor U8918 (N_8918,N_1164,N_3926);
or U8919 (N_8919,N_1966,N_1308);
or U8920 (N_8920,N_2709,N_2500);
and U8921 (N_8921,N_3263,N_651);
and U8922 (N_8922,N_47,N_4526);
nand U8923 (N_8923,N_4259,N_2096);
nor U8924 (N_8924,N_1776,N_3233);
nor U8925 (N_8925,N_1724,N_787);
or U8926 (N_8926,N_1978,N_75);
xor U8927 (N_8927,N_721,N_2425);
or U8928 (N_8928,N_3026,N_1488);
xnor U8929 (N_8929,N_1626,N_1337);
nor U8930 (N_8930,N_3560,N_4625);
nor U8931 (N_8931,N_2448,N_187);
nand U8932 (N_8932,N_1888,N_796);
or U8933 (N_8933,N_1163,N_3980);
and U8934 (N_8934,N_563,N_3828);
and U8935 (N_8935,N_523,N_61);
or U8936 (N_8936,N_2976,N_1533);
nor U8937 (N_8937,N_2774,N_1083);
and U8938 (N_8938,N_4052,N_598);
or U8939 (N_8939,N_794,N_3327);
nor U8940 (N_8940,N_1675,N_740);
or U8941 (N_8941,N_3886,N_573);
xor U8942 (N_8942,N_4409,N_4162);
and U8943 (N_8943,N_4009,N_1342);
or U8944 (N_8944,N_4635,N_2241);
xor U8945 (N_8945,N_1272,N_3108);
xor U8946 (N_8946,N_3552,N_1946);
nor U8947 (N_8947,N_681,N_2147);
xor U8948 (N_8948,N_4594,N_2053);
nor U8949 (N_8949,N_3578,N_889);
nand U8950 (N_8950,N_587,N_2803);
nor U8951 (N_8951,N_3135,N_2829);
nor U8952 (N_8952,N_2938,N_2857);
xor U8953 (N_8953,N_315,N_4893);
nor U8954 (N_8954,N_1780,N_4671);
xor U8955 (N_8955,N_4613,N_4930);
or U8956 (N_8956,N_3787,N_2646);
nor U8957 (N_8957,N_1295,N_563);
or U8958 (N_8958,N_4271,N_87);
or U8959 (N_8959,N_442,N_4626);
nor U8960 (N_8960,N_3898,N_2944);
or U8961 (N_8961,N_1906,N_4228);
and U8962 (N_8962,N_2442,N_2074);
xnor U8963 (N_8963,N_3453,N_3621);
and U8964 (N_8964,N_4517,N_2348);
and U8965 (N_8965,N_3564,N_4845);
nor U8966 (N_8966,N_3634,N_1126);
nand U8967 (N_8967,N_3327,N_3963);
nand U8968 (N_8968,N_3784,N_746);
xnor U8969 (N_8969,N_2974,N_3470);
nor U8970 (N_8970,N_784,N_2250);
and U8971 (N_8971,N_1398,N_1515);
and U8972 (N_8972,N_1251,N_3963);
and U8973 (N_8973,N_1105,N_4232);
nor U8974 (N_8974,N_4302,N_2209);
and U8975 (N_8975,N_4072,N_3916);
nand U8976 (N_8976,N_4167,N_2201);
nor U8977 (N_8977,N_2896,N_4914);
and U8978 (N_8978,N_4573,N_386);
nand U8979 (N_8979,N_1979,N_1882);
and U8980 (N_8980,N_1189,N_3680);
and U8981 (N_8981,N_2701,N_1453);
nor U8982 (N_8982,N_4371,N_2134);
nand U8983 (N_8983,N_4478,N_737);
or U8984 (N_8984,N_3943,N_1900);
or U8985 (N_8985,N_3060,N_3956);
or U8986 (N_8986,N_1426,N_3829);
nand U8987 (N_8987,N_563,N_3956);
nand U8988 (N_8988,N_838,N_773);
nand U8989 (N_8989,N_2393,N_3027);
and U8990 (N_8990,N_3200,N_3144);
nor U8991 (N_8991,N_2599,N_362);
nand U8992 (N_8992,N_368,N_4591);
xnor U8993 (N_8993,N_983,N_2029);
xor U8994 (N_8994,N_1057,N_794);
and U8995 (N_8995,N_3808,N_1717);
and U8996 (N_8996,N_317,N_3292);
nor U8997 (N_8997,N_3058,N_2612);
or U8998 (N_8998,N_4404,N_3483);
or U8999 (N_8999,N_1374,N_2134);
nand U9000 (N_9000,N_2661,N_576);
xor U9001 (N_9001,N_4703,N_4437);
or U9002 (N_9002,N_4290,N_445);
xor U9003 (N_9003,N_162,N_1952);
xnor U9004 (N_9004,N_4989,N_2625);
and U9005 (N_9005,N_1821,N_4950);
nand U9006 (N_9006,N_3705,N_3875);
xor U9007 (N_9007,N_4060,N_3146);
xnor U9008 (N_9008,N_1279,N_1990);
or U9009 (N_9009,N_3622,N_1133);
and U9010 (N_9010,N_1817,N_1914);
nor U9011 (N_9011,N_443,N_3899);
or U9012 (N_9012,N_4045,N_1548);
xor U9013 (N_9013,N_1856,N_2554);
xor U9014 (N_9014,N_3119,N_363);
xnor U9015 (N_9015,N_3473,N_1344);
nor U9016 (N_9016,N_371,N_2993);
nand U9017 (N_9017,N_3455,N_317);
xor U9018 (N_9018,N_2215,N_675);
xor U9019 (N_9019,N_4486,N_1670);
xor U9020 (N_9020,N_438,N_849);
nor U9021 (N_9021,N_2587,N_1096);
nand U9022 (N_9022,N_2958,N_2070);
or U9023 (N_9023,N_3218,N_4696);
nand U9024 (N_9024,N_4052,N_317);
nand U9025 (N_9025,N_3011,N_4820);
nand U9026 (N_9026,N_1723,N_2549);
nand U9027 (N_9027,N_4130,N_4254);
or U9028 (N_9028,N_50,N_3460);
and U9029 (N_9029,N_1961,N_2251);
nand U9030 (N_9030,N_63,N_3796);
nor U9031 (N_9031,N_997,N_367);
and U9032 (N_9032,N_3365,N_3847);
and U9033 (N_9033,N_1126,N_1836);
nand U9034 (N_9034,N_676,N_206);
xor U9035 (N_9035,N_2392,N_3515);
and U9036 (N_9036,N_2757,N_4289);
nand U9037 (N_9037,N_306,N_2222);
xnor U9038 (N_9038,N_1194,N_1041);
xnor U9039 (N_9039,N_4732,N_1121);
xor U9040 (N_9040,N_3476,N_3708);
nand U9041 (N_9041,N_292,N_3649);
nand U9042 (N_9042,N_4483,N_2680);
and U9043 (N_9043,N_2327,N_1682);
xor U9044 (N_9044,N_4739,N_860);
nand U9045 (N_9045,N_3453,N_2912);
nand U9046 (N_9046,N_807,N_2137);
and U9047 (N_9047,N_2938,N_4853);
nand U9048 (N_9048,N_1881,N_522);
and U9049 (N_9049,N_3792,N_246);
or U9050 (N_9050,N_4442,N_3564);
and U9051 (N_9051,N_3962,N_4395);
or U9052 (N_9052,N_3366,N_3488);
or U9053 (N_9053,N_1886,N_871);
nor U9054 (N_9054,N_2267,N_3258);
xnor U9055 (N_9055,N_2218,N_1306);
and U9056 (N_9056,N_1304,N_133);
and U9057 (N_9057,N_4705,N_4295);
nand U9058 (N_9058,N_1100,N_851);
nor U9059 (N_9059,N_3856,N_4818);
or U9060 (N_9060,N_4075,N_2982);
or U9061 (N_9061,N_2779,N_3898);
and U9062 (N_9062,N_4733,N_3350);
and U9063 (N_9063,N_3092,N_3886);
nand U9064 (N_9064,N_1577,N_2719);
nand U9065 (N_9065,N_449,N_3993);
nand U9066 (N_9066,N_3608,N_3781);
xnor U9067 (N_9067,N_2734,N_4742);
xnor U9068 (N_9068,N_1604,N_865);
and U9069 (N_9069,N_921,N_4589);
nand U9070 (N_9070,N_2345,N_317);
nand U9071 (N_9071,N_4318,N_1065);
nor U9072 (N_9072,N_1936,N_2060);
or U9073 (N_9073,N_3740,N_2393);
and U9074 (N_9074,N_3736,N_1083);
nand U9075 (N_9075,N_3165,N_3831);
and U9076 (N_9076,N_1991,N_3905);
nor U9077 (N_9077,N_4243,N_773);
and U9078 (N_9078,N_236,N_2526);
xor U9079 (N_9079,N_2468,N_1072);
or U9080 (N_9080,N_2975,N_1267);
or U9081 (N_9081,N_4669,N_4333);
xor U9082 (N_9082,N_4538,N_1569);
xor U9083 (N_9083,N_3014,N_2058);
nand U9084 (N_9084,N_2482,N_3517);
or U9085 (N_9085,N_2367,N_1160);
nand U9086 (N_9086,N_2390,N_690);
or U9087 (N_9087,N_1978,N_3328);
and U9088 (N_9088,N_1434,N_1946);
nand U9089 (N_9089,N_1023,N_262);
nand U9090 (N_9090,N_2794,N_4722);
nand U9091 (N_9091,N_3080,N_1928);
nand U9092 (N_9092,N_3766,N_3455);
nor U9093 (N_9093,N_4271,N_2228);
or U9094 (N_9094,N_2087,N_4955);
and U9095 (N_9095,N_2757,N_4578);
nand U9096 (N_9096,N_4401,N_2988);
or U9097 (N_9097,N_2053,N_1375);
nand U9098 (N_9098,N_4714,N_4133);
nor U9099 (N_9099,N_3479,N_1263);
and U9100 (N_9100,N_2159,N_342);
or U9101 (N_9101,N_3529,N_2458);
nor U9102 (N_9102,N_855,N_1983);
and U9103 (N_9103,N_2009,N_1744);
nand U9104 (N_9104,N_3236,N_3508);
nor U9105 (N_9105,N_246,N_4908);
nor U9106 (N_9106,N_2848,N_721);
and U9107 (N_9107,N_3353,N_1429);
xor U9108 (N_9108,N_21,N_4514);
nor U9109 (N_9109,N_1471,N_1863);
or U9110 (N_9110,N_141,N_1210);
and U9111 (N_9111,N_3628,N_571);
nor U9112 (N_9112,N_439,N_2876);
or U9113 (N_9113,N_684,N_4710);
nor U9114 (N_9114,N_2833,N_3257);
nor U9115 (N_9115,N_4398,N_205);
nor U9116 (N_9116,N_82,N_3420);
nand U9117 (N_9117,N_3868,N_1284);
or U9118 (N_9118,N_4706,N_4416);
xnor U9119 (N_9119,N_1125,N_2656);
or U9120 (N_9120,N_483,N_2272);
nand U9121 (N_9121,N_4022,N_3564);
xnor U9122 (N_9122,N_2380,N_1168);
or U9123 (N_9123,N_2084,N_1732);
nor U9124 (N_9124,N_1373,N_1071);
nand U9125 (N_9125,N_3635,N_1684);
and U9126 (N_9126,N_3031,N_4661);
nand U9127 (N_9127,N_3115,N_3034);
or U9128 (N_9128,N_3914,N_2601);
or U9129 (N_9129,N_2804,N_3565);
nor U9130 (N_9130,N_1351,N_1993);
nand U9131 (N_9131,N_4245,N_1700);
and U9132 (N_9132,N_2181,N_1426);
nand U9133 (N_9133,N_360,N_3896);
and U9134 (N_9134,N_2670,N_1834);
or U9135 (N_9135,N_3914,N_2599);
and U9136 (N_9136,N_2540,N_3735);
xnor U9137 (N_9137,N_891,N_1003);
nor U9138 (N_9138,N_1107,N_622);
nor U9139 (N_9139,N_3064,N_230);
and U9140 (N_9140,N_3987,N_1302);
xnor U9141 (N_9141,N_2871,N_711);
and U9142 (N_9142,N_3426,N_1746);
nand U9143 (N_9143,N_1327,N_2467);
xor U9144 (N_9144,N_3740,N_3799);
and U9145 (N_9145,N_4088,N_646);
xnor U9146 (N_9146,N_4886,N_446);
nand U9147 (N_9147,N_1544,N_2644);
and U9148 (N_9148,N_3819,N_2707);
xnor U9149 (N_9149,N_2987,N_3869);
and U9150 (N_9150,N_4127,N_2507);
nor U9151 (N_9151,N_3187,N_123);
and U9152 (N_9152,N_2096,N_752);
nand U9153 (N_9153,N_4807,N_200);
nand U9154 (N_9154,N_4384,N_662);
nor U9155 (N_9155,N_4293,N_1925);
nor U9156 (N_9156,N_1435,N_2475);
nand U9157 (N_9157,N_3152,N_3354);
nand U9158 (N_9158,N_3157,N_3411);
nand U9159 (N_9159,N_1823,N_4855);
or U9160 (N_9160,N_2033,N_1963);
xor U9161 (N_9161,N_995,N_2913);
nor U9162 (N_9162,N_3609,N_3357);
nand U9163 (N_9163,N_212,N_1755);
xnor U9164 (N_9164,N_1507,N_821);
or U9165 (N_9165,N_288,N_105);
and U9166 (N_9166,N_3274,N_2493);
xnor U9167 (N_9167,N_3635,N_2498);
and U9168 (N_9168,N_3470,N_4572);
nand U9169 (N_9169,N_2206,N_1769);
and U9170 (N_9170,N_1063,N_2413);
nor U9171 (N_9171,N_1823,N_415);
nor U9172 (N_9172,N_3679,N_3851);
and U9173 (N_9173,N_4859,N_94);
and U9174 (N_9174,N_2318,N_4119);
and U9175 (N_9175,N_2697,N_2404);
nor U9176 (N_9176,N_2875,N_284);
xnor U9177 (N_9177,N_4527,N_3993);
nor U9178 (N_9178,N_880,N_4052);
or U9179 (N_9179,N_3781,N_4880);
nor U9180 (N_9180,N_1237,N_2);
or U9181 (N_9181,N_4583,N_4207);
nand U9182 (N_9182,N_1192,N_1340);
or U9183 (N_9183,N_948,N_1665);
nor U9184 (N_9184,N_4723,N_2281);
nor U9185 (N_9185,N_2884,N_2799);
nand U9186 (N_9186,N_3616,N_4270);
nand U9187 (N_9187,N_1589,N_819);
and U9188 (N_9188,N_1344,N_4152);
xor U9189 (N_9189,N_4268,N_2235);
or U9190 (N_9190,N_1371,N_3034);
xor U9191 (N_9191,N_1939,N_3480);
nand U9192 (N_9192,N_4035,N_1081);
or U9193 (N_9193,N_3938,N_4516);
and U9194 (N_9194,N_1007,N_3430);
and U9195 (N_9195,N_1489,N_1749);
nor U9196 (N_9196,N_1547,N_2936);
xor U9197 (N_9197,N_4139,N_1006);
or U9198 (N_9198,N_242,N_1138);
or U9199 (N_9199,N_766,N_3188);
xor U9200 (N_9200,N_2699,N_2949);
xor U9201 (N_9201,N_138,N_913);
nand U9202 (N_9202,N_836,N_1916);
and U9203 (N_9203,N_4267,N_718);
nand U9204 (N_9204,N_3423,N_2701);
or U9205 (N_9205,N_2585,N_3006);
xnor U9206 (N_9206,N_3962,N_1101);
xnor U9207 (N_9207,N_1780,N_3795);
xnor U9208 (N_9208,N_2259,N_1874);
xor U9209 (N_9209,N_4872,N_3943);
nor U9210 (N_9210,N_1814,N_548);
and U9211 (N_9211,N_1973,N_4080);
nand U9212 (N_9212,N_3228,N_3928);
xnor U9213 (N_9213,N_1480,N_2680);
nor U9214 (N_9214,N_439,N_1364);
or U9215 (N_9215,N_4575,N_21);
and U9216 (N_9216,N_4318,N_837);
and U9217 (N_9217,N_2748,N_973);
nand U9218 (N_9218,N_4364,N_3913);
nand U9219 (N_9219,N_1584,N_3831);
nor U9220 (N_9220,N_2055,N_4684);
and U9221 (N_9221,N_1018,N_3321);
and U9222 (N_9222,N_1421,N_3776);
nand U9223 (N_9223,N_3332,N_3607);
nand U9224 (N_9224,N_2032,N_1241);
and U9225 (N_9225,N_3664,N_2569);
nand U9226 (N_9226,N_1513,N_1477);
or U9227 (N_9227,N_814,N_2314);
xor U9228 (N_9228,N_576,N_2003);
nand U9229 (N_9229,N_831,N_4111);
nor U9230 (N_9230,N_4738,N_981);
or U9231 (N_9231,N_3816,N_2208);
and U9232 (N_9232,N_1446,N_1972);
nor U9233 (N_9233,N_3247,N_1219);
nor U9234 (N_9234,N_316,N_3488);
and U9235 (N_9235,N_1887,N_618);
nand U9236 (N_9236,N_4866,N_482);
nand U9237 (N_9237,N_2943,N_4089);
nor U9238 (N_9238,N_210,N_726);
nor U9239 (N_9239,N_371,N_3750);
xor U9240 (N_9240,N_2456,N_2134);
xor U9241 (N_9241,N_4684,N_3860);
and U9242 (N_9242,N_1355,N_1290);
or U9243 (N_9243,N_4187,N_3031);
nor U9244 (N_9244,N_4620,N_4208);
xor U9245 (N_9245,N_1914,N_814);
nand U9246 (N_9246,N_1955,N_2196);
xnor U9247 (N_9247,N_485,N_149);
or U9248 (N_9248,N_4074,N_2410);
or U9249 (N_9249,N_179,N_4968);
nand U9250 (N_9250,N_3973,N_1821);
xor U9251 (N_9251,N_1481,N_3062);
and U9252 (N_9252,N_2724,N_1732);
and U9253 (N_9253,N_4742,N_860);
nor U9254 (N_9254,N_2418,N_919);
nand U9255 (N_9255,N_4798,N_2808);
nor U9256 (N_9256,N_4532,N_951);
nand U9257 (N_9257,N_2288,N_1808);
xnor U9258 (N_9258,N_4472,N_2085);
and U9259 (N_9259,N_3669,N_2696);
nand U9260 (N_9260,N_2724,N_4066);
nor U9261 (N_9261,N_1185,N_4020);
nor U9262 (N_9262,N_3924,N_1753);
xor U9263 (N_9263,N_1612,N_1325);
nor U9264 (N_9264,N_4220,N_1082);
and U9265 (N_9265,N_156,N_2332);
nor U9266 (N_9266,N_2856,N_796);
nor U9267 (N_9267,N_591,N_3173);
or U9268 (N_9268,N_3351,N_3612);
nor U9269 (N_9269,N_198,N_3828);
xor U9270 (N_9270,N_1844,N_464);
or U9271 (N_9271,N_556,N_2910);
nand U9272 (N_9272,N_1889,N_3783);
nand U9273 (N_9273,N_135,N_269);
xor U9274 (N_9274,N_2444,N_3760);
nor U9275 (N_9275,N_1493,N_1590);
xnor U9276 (N_9276,N_4666,N_4603);
and U9277 (N_9277,N_4604,N_3996);
nand U9278 (N_9278,N_4032,N_4926);
or U9279 (N_9279,N_485,N_1589);
xnor U9280 (N_9280,N_1929,N_4988);
and U9281 (N_9281,N_1071,N_2078);
nor U9282 (N_9282,N_1888,N_150);
nand U9283 (N_9283,N_3070,N_4272);
nand U9284 (N_9284,N_408,N_2188);
nand U9285 (N_9285,N_772,N_3158);
or U9286 (N_9286,N_4626,N_4316);
xor U9287 (N_9287,N_467,N_2514);
nor U9288 (N_9288,N_4934,N_209);
and U9289 (N_9289,N_1131,N_611);
nand U9290 (N_9290,N_1232,N_4814);
nand U9291 (N_9291,N_1310,N_1226);
nor U9292 (N_9292,N_4230,N_4348);
nor U9293 (N_9293,N_3203,N_84);
xnor U9294 (N_9294,N_1739,N_27);
or U9295 (N_9295,N_150,N_3263);
nand U9296 (N_9296,N_3006,N_771);
nand U9297 (N_9297,N_738,N_549);
and U9298 (N_9298,N_3976,N_3436);
nand U9299 (N_9299,N_1148,N_4466);
or U9300 (N_9300,N_2588,N_3326);
nand U9301 (N_9301,N_4845,N_4736);
nand U9302 (N_9302,N_4441,N_2385);
nor U9303 (N_9303,N_4675,N_1819);
xnor U9304 (N_9304,N_2923,N_4539);
nor U9305 (N_9305,N_2243,N_648);
nor U9306 (N_9306,N_276,N_3618);
or U9307 (N_9307,N_1344,N_2771);
xnor U9308 (N_9308,N_191,N_1121);
xnor U9309 (N_9309,N_4720,N_2253);
nand U9310 (N_9310,N_287,N_3866);
nor U9311 (N_9311,N_4189,N_2282);
nand U9312 (N_9312,N_4673,N_3453);
or U9313 (N_9313,N_4681,N_2575);
or U9314 (N_9314,N_3604,N_4543);
xor U9315 (N_9315,N_589,N_3835);
and U9316 (N_9316,N_592,N_178);
nand U9317 (N_9317,N_4518,N_1816);
or U9318 (N_9318,N_4211,N_3158);
and U9319 (N_9319,N_1242,N_2085);
or U9320 (N_9320,N_144,N_999);
and U9321 (N_9321,N_1012,N_2465);
nor U9322 (N_9322,N_218,N_2644);
or U9323 (N_9323,N_709,N_3362);
nand U9324 (N_9324,N_2578,N_4011);
and U9325 (N_9325,N_225,N_694);
nor U9326 (N_9326,N_3568,N_103);
and U9327 (N_9327,N_3941,N_110);
nand U9328 (N_9328,N_3835,N_406);
or U9329 (N_9329,N_3888,N_3625);
nor U9330 (N_9330,N_1094,N_1623);
nand U9331 (N_9331,N_2513,N_3410);
nor U9332 (N_9332,N_1688,N_1957);
or U9333 (N_9333,N_3718,N_1773);
nor U9334 (N_9334,N_1502,N_1812);
xor U9335 (N_9335,N_1351,N_407);
nor U9336 (N_9336,N_3025,N_4207);
nor U9337 (N_9337,N_4510,N_3852);
nand U9338 (N_9338,N_3477,N_2904);
xnor U9339 (N_9339,N_2843,N_172);
and U9340 (N_9340,N_361,N_2483);
nand U9341 (N_9341,N_3686,N_473);
nor U9342 (N_9342,N_2844,N_1705);
or U9343 (N_9343,N_2753,N_2845);
or U9344 (N_9344,N_451,N_3616);
and U9345 (N_9345,N_1196,N_3227);
nor U9346 (N_9346,N_1819,N_2359);
or U9347 (N_9347,N_352,N_225);
nor U9348 (N_9348,N_4748,N_4057);
xnor U9349 (N_9349,N_1619,N_3663);
nand U9350 (N_9350,N_567,N_359);
nand U9351 (N_9351,N_372,N_3460);
xnor U9352 (N_9352,N_1019,N_3375);
or U9353 (N_9353,N_283,N_4114);
or U9354 (N_9354,N_4354,N_4951);
xnor U9355 (N_9355,N_2718,N_3158);
and U9356 (N_9356,N_73,N_4218);
and U9357 (N_9357,N_1667,N_4888);
nand U9358 (N_9358,N_1559,N_1551);
nor U9359 (N_9359,N_483,N_2256);
or U9360 (N_9360,N_1640,N_1045);
nand U9361 (N_9361,N_999,N_1919);
nand U9362 (N_9362,N_4979,N_753);
nand U9363 (N_9363,N_4987,N_3443);
or U9364 (N_9364,N_2852,N_1455);
nor U9365 (N_9365,N_1701,N_320);
and U9366 (N_9366,N_2513,N_3000);
and U9367 (N_9367,N_4235,N_1013);
nor U9368 (N_9368,N_1257,N_4597);
and U9369 (N_9369,N_3394,N_2926);
or U9370 (N_9370,N_4916,N_2302);
nand U9371 (N_9371,N_594,N_3802);
nor U9372 (N_9372,N_2877,N_1611);
and U9373 (N_9373,N_169,N_3815);
or U9374 (N_9374,N_1432,N_3556);
nor U9375 (N_9375,N_3065,N_1613);
and U9376 (N_9376,N_1789,N_1224);
nor U9377 (N_9377,N_3608,N_1967);
and U9378 (N_9378,N_1419,N_3273);
and U9379 (N_9379,N_2366,N_3982);
xor U9380 (N_9380,N_2014,N_4896);
xnor U9381 (N_9381,N_2975,N_4788);
nor U9382 (N_9382,N_1018,N_1940);
or U9383 (N_9383,N_2796,N_2983);
nor U9384 (N_9384,N_4661,N_4546);
xnor U9385 (N_9385,N_596,N_3247);
xnor U9386 (N_9386,N_12,N_4011);
nand U9387 (N_9387,N_2645,N_1585);
nand U9388 (N_9388,N_3739,N_2762);
nor U9389 (N_9389,N_1866,N_614);
or U9390 (N_9390,N_3780,N_2658);
nand U9391 (N_9391,N_3374,N_3261);
xnor U9392 (N_9392,N_219,N_4420);
and U9393 (N_9393,N_58,N_1233);
or U9394 (N_9394,N_715,N_2073);
or U9395 (N_9395,N_1604,N_440);
xnor U9396 (N_9396,N_381,N_1731);
nor U9397 (N_9397,N_1585,N_1734);
nand U9398 (N_9398,N_204,N_3977);
xor U9399 (N_9399,N_1855,N_3577);
and U9400 (N_9400,N_2438,N_2985);
or U9401 (N_9401,N_1957,N_641);
nand U9402 (N_9402,N_3787,N_2418);
xnor U9403 (N_9403,N_606,N_3063);
or U9404 (N_9404,N_2658,N_506);
nand U9405 (N_9405,N_655,N_4617);
and U9406 (N_9406,N_1670,N_4618);
nand U9407 (N_9407,N_2482,N_3843);
or U9408 (N_9408,N_2026,N_1990);
nor U9409 (N_9409,N_3902,N_248);
xor U9410 (N_9410,N_3965,N_2075);
nand U9411 (N_9411,N_2890,N_3880);
nor U9412 (N_9412,N_4197,N_865);
nor U9413 (N_9413,N_2191,N_2592);
nor U9414 (N_9414,N_2539,N_2560);
or U9415 (N_9415,N_3562,N_3379);
xnor U9416 (N_9416,N_892,N_2858);
nor U9417 (N_9417,N_2558,N_666);
and U9418 (N_9418,N_4395,N_2658);
nand U9419 (N_9419,N_1566,N_3936);
or U9420 (N_9420,N_4369,N_4880);
and U9421 (N_9421,N_3995,N_605);
nor U9422 (N_9422,N_1866,N_3109);
and U9423 (N_9423,N_2257,N_2355);
xnor U9424 (N_9424,N_743,N_2520);
and U9425 (N_9425,N_954,N_3234);
or U9426 (N_9426,N_847,N_1032);
nor U9427 (N_9427,N_206,N_1303);
or U9428 (N_9428,N_2549,N_2308);
or U9429 (N_9429,N_522,N_4304);
nand U9430 (N_9430,N_4023,N_919);
or U9431 (N_9431,N_4310,N_4298);
nor U9432 (N_9432,N_197,N_2377);
nor U9433 (N_9433,N_3887,N_2124);
and U9434 (N_9434,N_4730,N_422);
nand U9435 (N_9435,N_412,N_4098);
nor U9436 (N_9436,N_3690,N_1397);
nand U9437 (N_9437,N_3827,N_2670);
nor U9438 (N_9438,N_3805,N_4709);
xnor U9439 (N_9439,N_3087,N_731);
nor U9440 (N_9440,N_977,N_3652);
xnor U9441 (N_9441,N_4140,N_373);
or U9442 (N_9442,N_438,N_1225);
and U9443 (N_9443,N_1003,N_3496);
xnor U9444 (N_9444,N_1230,N_4210);
nor U9445 (N_9445,N_2195,N_216);
or U9446 (N_9446,N_2609,N_443);
nor U9447 (N_9447,N_3317,N_4169);
nor U9448 (N_9448,N_704,N_3171);
or U9449 (N_9449,N_4227,N_3709);
nor U9450 (N_9450,N_4255,N_3740);
nor U9451 (N_9451,N_1623,N_4679);
and U9452 (N_9452,N_4905,N_237);
xnor U9453 (N_9453,N_2988,N_92);
or U9454 (N_9454,N_2391,N_4303);
nand U9455 (N_9455,N_4590,N_4519);
xnor U9456 (N_9456,N_99,N_2007);
and U9457 (N_9457,N_1898,N_4805);
nand U9458 (N_9458,N_3677,N_1568);
nor U9459 (N_9459,N_2940,N_3994);
and U9460 (N_9460,N_901,N_462);
nor U9461 (N_9461,N_371,N_209);
nand U9462 (N_9462,N_1189,N_2146);
or U9463 (N_9463,N_2508,N_2007);
and U9464 (N_9464,N_392,N_4322);
xnor U9465 (N_9465,N_2477,N_1097);
nor U9466 (N_9466,N_4096,N_4137);
nand U9467 (N_9467,N_4818,N_4033);
and U9468 (N_9468,N_2915,N_1141);
xor U9469 (N_9469,N_2406,N_155);
nor U9470 (N_9470,N_3659,N_3826);
nand U9471 (N_9471,N_1456,N_692);
and U9472 (N_9472,N_835,N_1420);
and U9473 (N_9473,N_381,N_2104);
and U9474 (N_9474,N_2064,N_2393);
nor U9475 (N_9475,N_2634,N_1790);
or U9476 (N_9476,N_1487,N_2636);
and U9477 (N_9477,N_3104,N_1881);
xnor U9478 (N_9478,N_2465,N_3696);
nand U9479 (N_9479,N_4719,N_3962);
or U9480 (N_9480,N_2320,N_2759);
nand U9481 (N_9481,N_4780,N_2178);
nand U9482 (N_9482,N_1077,N_3650);
xor U9483 (N_9483,N_4408,N_2023);
or U9484 (N_9484,N_4209,N_2232);
nand U9485 (N_9485,N_775,N_95);
or U9486 (N_9486,N_3617,N_3185);
or U9487 (N_9487,N_2503,N_4054);
and U9488 (N_9488,N_1223,N_155);
or U9489 (N_9489,N_1020,N_4383);
nand U9490 (N_9490,N_1908,N_916);
xnor U9491 (N_9491,N_1190,N_1131);
xnor U9492 (N_9492,N_993,N_20);
nand U9493 (N_9493,N_3832,N_79);
xnor U9494 (N_9494,N_1649,N_916);
or U9495 (N_9495,N_2774,N_179);
nand U9496 (N_9496,N_4845,N_2523);
nand U9497 (N_9497,N_367,N_3206);
and U9498 (N_9498,N_1032,N_1172);
nor U9499 (N_9499,N_4006,N_1840);
or U9500 (N_9500,N_581,N_3752);
xor U9501 (N_9501,N_392,N_4480);
or U9502 (N_9502,N_2310,N_4652);
nand U9503 (N_9503,N_4403,N_631);
nor U9504 (N_9504,N_920,N_2913);
and U9505 (N_9505,N_2996,N_4514);
and U9506 (N_9506,N_3858,N_3838);
and U9507 (N_9507,N_1863,N_653);
nor U9508 (N_9508,N_392,N_3267);
xnor U9509 (N_9509,N_4951,N_2596);
or U9510 (N_9510,N_4986,N_1170);
nand U9511 (N_9511,N_2372,N_2394);
nor U9512 (N_9512,N_2589,N_688);
and U9513 (N_9513,N_4931,N_527);
and U9514 (N_9514,N_2800,N_3104);
nor U9515 (N_9515,N_2394,N_126);
xnor U9516 (N_9516,N_3096,N_1657);
nor U9517 (N_9517,N_3312,N_3351);
or U9518 (N_9518,N_4157,N_2246);
nor U9519 (N_9519,N_1807,N_1662);
and U9520 (N_9520,N_388,N_4757);
nand U9521 (N_9521,N_3669,N_2530);
nand U9522 (N_9522,N_1304,N_4250);
xnor U9523 (N_9523,N_4972,N_1003);
and U9524 (N_9524,N_4210,N_3613);
nand U9525 (N_9525,N_1153,N_105);
and U9526 (N_9526,N_3264,N_1968);
or U9527 (N_9527,N_1472,N_872);
and U9528 (N_9528,N_3341,N_4829);
or U9529 (N_9529,N_3511,N_1382);
nor U9530 (N_9530,N_2114,N_3220);
and U9531 (N_9531,N_3418,N_4176);
or U9532 (N_9532,N_1340,N_3393);
nand U9533 (N_9533,N_380,N_459);
nand U9534 (N_9534,N_4389,N_1502);
xnor U9535 (N_9535,N_4182,N_1745);
nor U9536 (N_9536,N_697,N_2202);
and U9537 (N_9537,N_3328,N_1219);
nor U9538 (N_9538,N_4584,N_3779);
and U9539 (N_9539,N_868,N_3999);
and U9540 (N_9540,N_121,N_273);
and U9541 (N_9541,N_1034,N_3509);
nand U9542 (N_9542,N_3406,N_921);
nand U9543 (N_9543,N_4588,N_1186);
and U9544 (N_9544,N_2485,N_808);
or U9545 (N_9545,N_1557,N_4712);
nand U9546 (N_9546,N_3918,N_207);
nor U9547 (N_9547,N_4760,N_834);
nand U9548 (N_9548,N_4874,N_2071);
and U9549 (N_9549,N_3388,N_4430);
nor U9550 (N_9550,N_4176,N_2938);
nand U9551 (N_9551,N_3688,N_737);
and U9552 (N_9552,N_4115,N_4592);
nor U9553 (N_9553,N_2064,N_2347);
xnor U9554 (N_9554,N_3833,N_633);
and U9555 (N_9555,N_793,N_2670);
or U9556 (N_9556,N_4726,N_1877);
or U9557 (N_9557,N_3936,N_4160);
xnor U9558 (N_9558,N_3700,N_4239);
nor U9559 (N_9559,N_2060,N_1576);
nand U9560 (N_9560,N_3484,N_3825);
and U9561 (N_9561,N_1904,N_1025);
or U9562 (N_9562,N_2522,N_3840);
xor U9563 (N_9563,N_1134,N_4310);
or U9564 (N_9564,N_3215,N_1972);
nand U9565 (N_9565,N_1585,N_39);
xor U9566 (N_9566,N_347,N_959);
or U9567 (N_9567,N_2928,N_3240);
and U9568 (N_9568,N_843,N_3441);
xnor U9569 (N_9569,N_3424,N_4749);
or U9570 (N_9570,N_2172,N_594);
xnor U9571 (N_9571,N_2982,N_2790);
nand U9572 (N_9572,N_4074,N_4702);
or U9573 (N_9573,N_452,N_138);
xor U9574 (N_9574,N_3332,N_1854);
and U9575 (N_9575,N_1573,N_3874);
or U9576 (N_9576,N_3777,N_36);
nor U9577 (N_9577,N_26,N_4714);
or U9578 (N_9578,N_2145,N_960);
xnor U9579 (N_9579,N_748,N_1169);
nor U9580 (N_9580,N_4768,N_1066);
nor U9581 (N_9581,N_2744,N_2479);
and U9582 (N_9582,N_3074,N_2258);
nor U9583 (N_9583,N_4144,N_2579);
or U9584 (N_9584,N_207,N_1772);
or U9585 (N_9585,N_629,N_2634);
and U9586 (N_9586,N_3264,N_240);
nand U9587 (N_9587,N_1621,N_2809);
nor U9588 (N_9588,N_360,N_4676);
nor U9589 (N_9589,N_132,N_3093);
nand U9590 (N_9590,N_2308,N_3026);
nand U9591 (N_9591,N_3963,N_1065);
nor U9592 (N_9592,N_4494,N_4965);
xor U9593 (N_9593,N_275,N_3055);
nor U9594 (N_9594,N_4993,N_3206);
nand U9595 (N_9595,N_4341,N_538);
and U9596 (N_9596,N_216,N_587);
and U9597 (N_9597,N_2027,N_4210);
nor U9598 (N_9598,N_1524,N_2259);
xnor U9599 (N_9599,N_3004,N_4058);
and U9600 (N_9600,N_1342,N_3451);
and U9601 (N_9601,N_1096,N_940);
xor U9602 (N_9602,N_3855,N_2660);
nand U9603 (N_9603,N_781,N_1004);
or U9604 (N_9604,N_3156,N_137);
and U9605 (N_9605,N_1784,N_3756);
or U9606 (N_9606,N_4808,N_417);
and U9607 (N_9607,N_4879,N_621);
nor U9608 (N_9608,N_1992,N_3666);
and U9609 (N_9609,N_416,N_1554);
nand U9610 (N_9610,N_1570,N_1607);
and U9611 (N_9611,N_278,N_1443);
or U9612 (N_9612,N_4500,N_1114);
xor U9613 (N_9613,N_4506,N_821);
nor U9614 (N_9614,N_1958,N_970);
nor U9615 (N_9615,N_3901,N_4005);
or U9616 (N_9616,N_3766,N_4709);
xor U9617 (N_9617,N_2779,N_2363);
and U9618 (N_9618,N_128,N_3234);
nand U9619 (N_9619,N_990,N_1013);
nand U9620 (N_9620,N_4997,N_2682);
nand U9621 (N_9621,N_3046,N_2501);
nand U9622 (N_9622,N_2663,N_2313);
xnor U9623 (N_9623,N_2754,N_1344);
or U9624 (N_9624,N_941,N_2483);
nand U9625 (N_9625,N_3159,N_3107);
xnor U9626 (N_9626,N_612,N_909);
or U9627 (N_9627,N_1877,N_2513);
xor U9628 (N_9628,N_2306,N_157);
nand U9629 (N_9629,N_3008,N_2064);
or U9630 (N_9630,N_2822,N_4091);
nand U9631 (N_9631,N_1768,N_3223);
nor U9632 (N_9632,N_555,N_3917);
nor U9633 (N_9633,N_1904,N_36);
nand U9634 (N_9634,N_3931,N_3859);
nand U9635 (N_9635,N_4849,N_4500);
or U9636 (N_9636,N_3269,N_943);
nor U9637 (N_9637,N_2817,N_1114);
and U9638 (N_9638,N_468,N_4150);
and U9639 (N_9639,N_3400,N_690);
and U9640 (N_9640,N_258,N_56);
and U9641 (N_9641,N_1039,N_2575);
nand U9642 (N_9642,N_1645,N_3860);
and U9643 (N_9643,N_4236,N_263);
nor U9644 (N_9644,N_1411,N_4598);
xor U9645 (N_9645,N_373,N_2478);
nand U9646 (N_9646,N_721,N_3);
nor U9647 (N_9647,N_2446,N_3827);
nand U9648 (N_9648,N_1530,N_3812);
xnor U9649 (N_9649,N_4268,N_197);
nor U9650 (N_9650,N_3722,N_817);
nor U9651 (N_9651,N_4173,N_674);
nand U9652 (N_9652,N_892,N_4827);
nand U9653 (N_9653,N_1123,N_2685);
and U9654 (N_9654,N_155,N_716);
nor U9655 (N_9655,N_2896,N_1263);
and U9656 (N_9656,N_1129,N_2405);
xnor U9657 (N_9657,N_3291,N_837);
nand U9658 (N_9658,N_51,N_2749);
and U9659 (N_9659,N_2404,N_3669);
xnor U9660 (N_9660,N_3786,N_4664);
xor U9661 (N_9661,N_3120,N_2249);
and U9662 (N_9662,N_3431,N_4489);
nor U9663 (N_9663,N_4470,N_3947);
xor U9664 (N_9664,N_3329,N_3661);
or U9665 (N_9665,N_725,N_3848);
or U9666 (N_9666,N_4832,N_2754);
and U9667 (N_9667,N_791,N_4715);
and U9668 (N_9668,N_419,N_1640);
and U9669 (N_9669,N_1649,N_1753);
or U9670 (N_9670,N_3656,N_637);
nor U9671 (N_9671,N_608,N_3262);
nand U9672 (N_9672,N_1207,N_4129);
or U9673 (N_9673,N_3811,N_1241);
nand U9674 (N_9674,N_2875,N_1792);
nor U9675 (N_9675,N_2873,N_2588);
or U9676 (N_9676,N_577,N_3327);
nor U9677 (N_9677,N_1274,N_2710);
nand U9678 (N_9678,N_89,N_1164);
xnor U9679 (N_9679,N_1361,N_3846);
xor U9680 (N_9680,N_3273,N_529);
and U9681 (N_9681,N_3389,N_2381);
or U9682 (N_9682,N_2000,N_3424);
xor U9683 (N_9683,N_2183,N_673);
or U9684 (N_9684,N_4495,N_3620);
and U9685 (N_9685,N_1125,N_3500);
or U9686 (N_9686,N_1618,N_1988);
nor U9687 (N_9687,N_223,N_4709);
and U9688 (N_9688,N_4331,N_3496);
nor U9689 (N_9689,N_2987,N_4424);
xor U9690 (N_9690,N_3996,N_1384);
or U9691 (N_9691,N_2044,N_1400);
nand U9692 (N_9692,N_3643,N_923);
nor U9693 (N_9693,N_2662,N_4503);
nand U9694 (N_9694,N_1225,N_3352);
nand U9695 (N_9695,N_1191,N_1358);
or U9696 (N_9696,N_2359,N_4942);
or U9697 (N_9697,N_1025,N_4999);
xor U9698 (N_9698,N_2468,N_2780);
or U9699 (N_9699,N_522,N_4420);
or U9700 (N_9700,N_1303,N_342);
and U9701 (N_9701,N_1909,N_4384);
and U9702 (N_9702,N_1965,N_2533);
nand U9703 (N_9703,N_3482,N_2021);
or U9704 (N_9704,N_985,N_1707);
xor U9705 (N_9705,N_2773,N_2503);
nor U9706 (N_9706,N_815,N_492);
xor U9707 (N_9707,N_4864,N_3284);
nand U9708 (N_9708,N_578,N_513);
nor U9709 (N_9709,N_2979,N_1712);
xor U9710 (N_9710,N_3360,N_2984);
xnor U9711 (N_9711,N_572,N_3738);
nor U9712 (N_9712,N_290,N_1317);
nor U9713 (N_9713,N_4432,N_2656);
nand U9714 (N_9714,N_2017,N_4070);
nand U9715 (N_9715,N_3338,N_2527);
or U9716 (N_9716,N_3895,N_1660);
xor U9717 (N_9717,N_4984,N_2439);
and U9718 (N_9718,N_3221,N_4388);
nand U9719 (N_9719,N_2431,N_875);
or U9720 (N_9720,N_1182,N_2152);
and U9721 (N_9721,N_2598,N_1147);
or U9722 (N_9722,N_1610,N_1063);
nor U9723 (N_9723,N_4244,N_1568);
nand U9724 (N_9724,N_2264,N_2667);
or U9725 (N_9725,N_1366,N_344);
or U9726 (N_9726,N_2820,N_2760);
and U9727 (N_9727,N_4568,N_2924);
nand U9728 (N_9728,N_1270,N_3031);
and U9729 (N_9729,N_557,N_2568);
nor U9730 (N_9730,N_3444,N_2979);
nand U9731 (N_9731,N_4820,N_1195);
and U9732 (N_9732,N_4388,N_1381);
and U9733 (N_9733,N_4796,N_508);
nand U9734 (N_9734,N_3402,N_1908);
nor U9735 (N_9735,N_1268,N_2279);
xor U9736 (N_9736,N_1489,N_4409);
nor U9737 (N_9737,N_1193,N_3344);
xor U9738 (N_9738,N_412,N_3841);
nor U9739 (N_9739,N_4987,N_1221);
or U9740 (N_9740,N_2585,N_623);
nand U9741 (N_9741,N_2126,N_3731);
nand U9742 (N_9742,N_2549,N_326);
and U9743 (N_9743,N_2432,N_2214);
or U9744 (N_9744,N_1397,N_2030);
nor U9745 (N_9745,N_2502,N_355);
or U9746 (N_9746,N_83,N_17);
and U9747 (N_9747,N_3309,N_284);
and U9748 (N_9748,N_4563,N_3089);
nand U9749 (N_9749,N_4094,N_2101);
and U9750 (N_9750,N_2805,N_1324);
nand U9751 (N_9751,N_1998,N_3877);
nand U9752 (N_9752,N_3959,N_4483);
and U9753 (N_9753,N_4292,N_3395);
or U9754 (N_9754,N_2457,N_272);
nand U9755 (N_9755,N_3998,N_1943);
xnor U9756 (N_9756,N_1062,N_4370);
and U9757 (N_9757,N_2491,N_1956);
or U9758 (N_9758,N_359,N_2662);
and U9759 (N_9759,N_2802,N_1497);
nand U9760 (N_9760,N_4991,N_4240);
and U9761 (N_9761,N_2804,N_4153);
nor U9762 (N_9762,N_2714,N_668);
nand U9763 (N_9763,N_2230,N_1403);
nor U9764 (N_9764,N_3160,N_3439);
nor U9765 (N_9765,N_1554,N_2853);
xor U9766 (N_9766,N_3897,N_2407);
or U9767 (N_9767,N_4075,N_2705);
xor U9768 (N_9768,N_526,N_393);
xor U9769 (N_9769,N_2977,N_956);
xor U9770 (N_9770,N_2706,N_4272);
nor U9771 (N_9771,N_112,N_2230);
xnor U9772 (N_9772,N_3067,N_4996);
nand U9773 (N_9773,N_2753,N_3341);
xor U9774 (N_9774,N_632,N_1550);
nand U9775 (N_9775,N_2950,N_265);
xor U9776 (N_9776,N_4231,N_1118);
nor U9777 (N_9777,N_3498,N_1306);
nor U9778 (N_9778,N_4000,N_185);
or U9779 (N_9779,N_322,N_184);
nor U9780 (N_9780,N_3589,N_3954);
xnor U9781 (N_9781,N_2426,N_821);
nor U9782 (N_9782,N_4021,N_1745);
nand U9783 (N_9783,N_4194,N_4391);
xor U9784 (N_9784,N_2823,N_4314);
or U9785 (N_9785,N_2451,N_1001);
nand U9786 (N_9786,N_1869,N_4062);
xnor U9787 (N_9787,N_1092,N_3392);
or U9788 (N_9788,N_3245,N_4840);
and U9789 (N_9789,N_2051,N_436);
xor U9790 (N_9790,N_1654,N_3411);
or U9791 (N_9791,N_856,N_2796);
nand U9792 (N_9792,N_1496,N_19);
nor U9793 (N_9793,N_2971,N_1813);
xor U9794 (N_9794,N_3903,N_2368);
or U9795 (N_9795,N_1088,N_141);
xor U9796 (N_9796,N_2717,N_3756);
nor U9797 (N_9797,N_4283,N_3578);
xnor U9798 (N_9798,N_557,N_3931);
xnor U9799 (N_9799,N_2247,N_3744);
nor U9800 (N_9800,N_4265,N_3387);
and U9801 (N_9801,N_4877,N_1949);
nor U9802 (N_9802,N_1678,N_3626);
nor U9803 (N_9803,N_3827,N_4562);
and U9804 (N_9804,N_270,N_3566);
nand U9805 (N_9805,N_2646,N_3810);
nand U9806 (N_9806,N_279,N_1172);
and U9807 (N_9807,N_382,N_1275);
or U9808 (N_9808,N_3898,N_2432);
xor U9809 (N_9809,N_2631,N_2721);
xnor U9810 (N_9810,N_2467,N_4360);
and U9811 (N_9811,N_3450,N_4981);
nor U9812 (N_9812,N_4856,N_4178);
nand U9813 (N_9813,N_44,N_2439);
and U9814 (N_9814,N_4162,N_714);
or U9815 (N_9815,N_4228,N_225);
nor U9816 (N_9816,N_2070,N_817);
nor U9817 (N_9817,N_721,N_1305);
or U9818 (N_9818,N_2071,N_1869);
or U9819 (N_9819,N_1,N_1984);
or U9820 (N_9820,N_4769,N_4408);
xnor U9821 (N_9821,N_4008,N_1793);
nand U9822 (N_9822,N_958,N_111);
xnor U9823 (N_9823,N_1051,N_3044);
and U9824 (N_9824,N_1480,N_2116);
nor U9825 (N_9825,N_618,N_4995);
xor U9826 (N_9826,N_3832,N_367);
or U9827 (N_9827,N_3919,N_519);
and U9828 (N_9828,N_1062,N_2968);
xor U9829 (N_9829,N_4053,N_2460);
xnor U9830 (N_9830,N_196,N_2295);
nor U9831 (N_9831,N_4115,N_4286);
or U9832 (N_9832,N_3533,N_1250);
nor U9833 (N_9833,N_734,N_3725);
or U9834 (N_9834,N_146,N_1175);
xor U9835 (N_9835,N_766,N_1056);
xnor U9836 (N_9836,N_3427,N_2070);
nor U9837 (N_9837,N_528,N_4552);
and U9838 (N_9838,N_698,N_1679);
nand U9839 (N_9839,N_3922,N_1792);
nand U9840 (N_9840,N_1009,N_403);
nand U9841 (N_9841,N_2688,N_4343);
or U9842 (N_9842,N_1297,N_452);
or U9843 (N_9843,N_2184,N_3179);
nand U9844 (N_9844,N_815,N_3110);
xor U9845 (N_9845,N_250,N_3691);
and U9846 (N_9846,N_988,N_1481);
nor U9847 (N_9847,N_3205,N_4721);
or U9848 (N_9848,N_4045,N_3327);
nor U9849 (N_9849,N_4437,N_2263);
nand U9850 (N_9850,N_3036,N_2335);
and U9851 (N_9851,N_4600,N_4227);
nand U9852 (N_9852,N_2534,N_2325);
or U9853 (N_9853,N_1095,N_4639);
nand U9854 (N_9854,N_490,N_4444);
nor U9855 (N_9855,N_2237,N_3286);
and U9856 (N_9856,N_1284,N_835);
or U9857 (N_9857,N_2821,N_3707);
or U9858 (N_9858,N_749,N_3137);
or U9859 (N_9859,N_3984,N_2255);
or U9860 (N_9860,N_1024,N_2340);
and U9861 (N_9861,N_3659,N_1071);
or U9862 (N_9862,N_787,N_2378);
or U9863 (N_9863,N_2151,N_1558);
nor U9864 (N_9864,N_3250,N_2268);
xor U9865 (N_9865,N_4937,N_551);
xor U9866 (N_9866,N_1590,N_192);
nor U9867 (N_9867,N_4397,N_3593);
nand U9868 (N_9868,N_4014,N_709);
or U9869 (N_9869,N_239,N_1608);
xnor U9870 (N_9870,N_3127,N_4419);
nand U9871 (N_9871,N_4019,N_349);
and U9872 (N_9872,N_2905,N_376);
nor U9873 (N_9873,N_1097,N_336);
or U9874 (N_9874,N_4070,N_2435);
or U9875 (N_9875,N_4240,N_3708);
nor U9876 (N_9876,N_4700,N_1271);
or U9877 (N_9877,N_2178,N_1493);
nor U9878 (N_9878,N_4138,N_1959);
nor U9879 (N_9879,N_2081,N_1119);
xor U9880 (N_9880,N_1553,N_213);
and U9881 (N_9881,N_4200,N_803);
nand U9882 (N_9882,N_73,N_4369);
nand U9883 (N_9883,N_3059,N_1138);
nor U9884 (N_9884,N_4434,N_4137);
xnor U9885 (N_9885,N_3301,N_4214);
and U9886 (N_9886,N_4669,N_2637);
or U9887 (N_9887,N_1164,N_1900);
xor U9888 (N_9888,N_4637,N_4422);
xor U9889 (N_9889,N_3040,N_2908);
nor U9890 (N_9890,N_2619,N_1212);
or U9891 (N_9891,N_73,N_3884);
or U9892 (N_9892,N_3957,N_4492);
nand U9893 (N_9893,N_1315,N_595);
or U9894 (N_9894,N_3590,N_4593);
xor U9895 (N_9895,N_87,N_1145);
nand U9896 (N_9896,N_3139,N_4177);
nor U9897 (N_9897,N_4306,N_2660);
nand U9898 (N_9898,N_3569,N_3532);
nand U9899 (N_9899,N_340,N_1082);
and U9900 (N_9900,N_717,N_1706);
xnor U9901 (N_9901,N_4675,N_1624);
xor U9902 (N_9902,N_3466,N_1898);
and U9903 (N_9903,N_4182,N_1970);
nand U9904 (N_9904,N_585,N_1785);
xnor U9905 (N_9905,N_2576,N_4869);
nand U9906 (N_9906,N_2309,N_2843);
and U9907 (N_9907,N_2197,N_2742);
and U9908 (N_9908,N_1524,N_1020);
nor U9909 (N_9909,N_1029,N_4319);
or U9910 (N_9910,N_427,N_4205);
nor U9911 (N_9911,N_1103,N_1829);
and U9912 (N_9912,N_657,N_2268);
nor U9913 (N_9913,N_4486,N_4110);
and U9914 (N_9914,N_1794,N_4274);
or U9915 (N_9915,N_1610,N_3294);
nand U9916 (N_9916,N_3490,N_4435);
or U9917 (N_9917,N_1159,N_2657);
nor U9918 (N_9918,N_1455,N_1960);
xor U9919 (N_9919,N_2988,N_2009);
or U9920 (N_9920,N_268,N_3228);
and U9921 (N_9921,N_4066,N_4513);
xnor U9922 (N_9922,N_2857,N_1785);
and U9923 (N_9923,N_3470,N_2623);
or U9924 (N_9924,N_244,N_1937);
nand U9925 (N_9925,N_3277,N_457);
nand U9926 (N_9926,N_1881,N_4746);
or U9927 (N_9927,N_1199,N_4428);
xor U9928 (N_9928,N_27,N_1878);
or U9929 (N_9929,N_852,N_670);
and U9930 (N_9930,N_3457,N_1477);
or U9931 (N_9931,N_270,N_3610);
or U9932 (N_9932,N_4362,N_429);
nor U9933 (N_9933,N_4498,N_4079);
nand U9934 (N_9934,N_3712,N_4029);
nor U9935 (N_9935,N_4268,N_1821);
or U9936 (N_9936,N_4638,N_3988);
nor U9937 (N_9937,N_3784,N_146);
nor U9938 (N_9938,N_123,N_1941);
nor U9939 (N_9939,N_4108,N_4264);
nor U9940 (N_9940,N_1009,N_64);
nor U9941 (N_9941,N_400,N_1948);
and U9942 (N_9942,N_4753,N_2185);
or U9943 (N_9943,N_2146,N_1560);
or U9944 (N_9944,N_32,N_4239);
and U9945 (N_9945,N_3902,N_1658);
xnor U9946 (N_9946,N_671,N_2392);
or U9947 (N_9947,N_3253,N_1799);
nor U9948 (N_9948,N_2364,N_1505);
or U9949 (N_9949,N_430,N_3208);
and U9950 (N_9950,N_4391,N_1853);
and U9951 (N_9951,N_4086,N_2073);
or U9952 (N_9952,N_341,N_1840);
xor U9953 (N_9953,N_3839,N_729);
and U9954 (N_9954,N_922,N_3743);
and U9955 (N_9955,N_2129,N_4459);
or U9956 (N_9956,N_1080,N_4106);
and U9957 (N_9957,N_590,N_1285);
and U9958 (N_9958,N_1393,N_4534);
and U9959 (N_9959,N_4614,N_1245);
and U9960 (N_9960,N_2876,N_913);
nand U9961 (N_9961,N_2163,N_1118);
nand U9962 (N_9962,N_1904,N_1077);
nor U9963 (N_9963,N_705,N_3234);
nand U9964 (N_9964,N_2193,N_3442);
and U9965 (N_9965,N_3412,N_3579);
nand U9966 (N_9966,N_3252,N_149);
nand U9967 (N_9967,N_3692,N_3376);
or U9968 (N_9968,N_1870,N_3926);
and U9969 (N_9969,N_1648,N_4594);
or U9970 (N_9970,N_2267,N_4845);
and U9971 (N_9971,N_3350,N_3686);
nand U9972 (N_9972,N_1928,N_3583);
or U9973 (N_9973,N_3370,N_2864);
nor U9974 (N_9974,N_4908,N_2291);
nand U9975 (N_9975,N_1960,N_706);
xor U9976 (N_9976,N_3106,N_249);
xnor U9977 (N_9977,N_156,N_1054);
nor U9978 (N_9978,N_842,N_1835);
and U9979 (N_9979,N_4488,N_1524);
or U9980 (N_9980,N_2254,N_4591);
and U9981 (N_9981,N_4536,N_3612);
or U9982 (N_9982,N_3458,N_4709);
nand U9983 (N_9983,N_587,N_188);
xor U9984 (N_9984,N_248,N_2795);
nand U9985 (N_9985,N_4180,N_1176);
xnor U9986 (N_9986,N_2522,N_1475);
or U9987 (N_9987,N_734,N_3062);
or U9988 (N_9988,N_2159,N_415);
or U9989 (N_9989,N_2722,N_2719);
and U9990 (N_9990,N_3107,N_3503);
and U9991 (N_9991,N_3067,N_2156);
nand U9992 (N_9992,N_4557,N_1366);
and U9993 (N_9993,N_2540,N_309);
and U9994 (N_9994,N_349,N_2215);
or U9995 (N_9995,N_2809,N_4876);
and U9996 (N_9996,N_1506,N_2309);
nor U9997 (N_9997,N_4837,N_4419);
xnor U9998 (N_9998,N_3954,N_2349);
nor U9999 (N_9999,N_4370,N_347);
nand U10000 (N_10000,N_9977,N_7333);
nor U10001 (N_10001,N_7149,N_6388);
nor U10002 (N_10002,N_8573,N_5281);
and U10003 (N_10003,N_9696,N_9554);
and U10004 (N_10004,N_9341,N_9706);
and U10005 (N_10005,N_8625,N_9293);
nor U10006 (N_10006,N_5351,N_6052);
and U10007 (N_10007,N_5532,N_9713);
xor U10008 (N_10008,N_9356,N_7674);
xor U10009 (N_10009,N_6498,N_9903);
xnor U10010 (N_10010,N_7820,N_5677);
xor U10011 (N_10011,N_6735,N_8537);
xnor U10012 (N_10012,N_5077,N_5495);
xor U10013 (N_10013,N_6037,N_6552);
xor U10014 (N_10014,N_7195,N_6973);
xnor U10015 (N_10015,N_5953,N_7102);
xnor U10016 (N_10016,N_6674,N_6044);
and U10017 (N_10017,N_9628,N_8549);
and U10018 (N_10018,N_5441,N_9039);
xnor U10019 (N_10019,N_8843,N_6862);
nor U10020 (N_10020,N_5059,N_9883);
nand U10021 (N_10021,N_8788,N_7724);
and U10022 (N_10022,N_6506,N_7637);
xnor U10023 (N_10023,N_8673,N_7980);
nor U10024 (N_10024,N_7666,N_8197);
xor U10025 (N_10025,N_9645,N_7911);
nor U10026 (N_10026,N_6734,N_7434);
xnor U10027 (N_10027,N_7878,N_6134);
xnor U10028 (N_10028,N_8966,N_8050);
nor U10029 (N_10029,N_6744,N_8322);
nand U10030 (N_10030,N_6984,N_7017);
xnor U10031 (N_10031,N_9643,N_5748);
xor U10032 (N_10032,N_7369,N_8959);
and U10033 (N_10033,N_7902,N_5029);
nand U10034 (N_10034,N_9011,N_5116);
nand U10035 (N_10035,N_7209,N_8137);
and U10036 (N_10036,N_5421,N_9391);
and U10037 (N_10037,N_6718,N_8449);
nand U10038 (N_10038,N_9575,N_7470);
xnor U10039 (N_10039,N_6156,N_9567);
nor U10040 (N_10040,N_5669,N_8694);
nor U10041 (N_10041,N_5721,N_8619);
xor U10042 (N_10042,N_8978,N_8266);
nor U10043 (N_10043,N_6036,N_5335);
nand U10044 (N_10044,N_5655,N_6207);
nor U10045 (N_10045,N_8986,N_8205);
xor U10046 (N_10046,N_7711,N_6790);
xor U10047 (N_10047,N_7973,N_9846);
nand U10048 (N_10048,N_6701,N_6869);
nor U10049 (N_10049,N_7979,N_5823);
xnor U10050 (N_10050,N_8662,N_9679);
or U10051 (N_10051,N_8627,N_5924);
or U10052 (N_10052,N_9657,N_5490);
or U10053 (N_10053,N_6126,N_9133);
and U10054 (N_10054,N_7400,N_7321);
or U10055 (N_10055,N_7588,N_8009);
xnor U10056 (N_10056,N_8028,N_9818);
nor U10057 (N_10057,N_8291,N_9754);
or U10058 (N_10058,N_9819,N_6454);
and U10059 (N_10059,N_7393,N_9944);
nor U10060 (N_10060,N_9894,N_6033);
nand U10061 (N_10061,N_9266,N_9904);
and U10062 (N_10062,N_6611,N_5512);
nor U10063 (N_10063,N_5310,N_9017);
nor U10064 (N_10064,N_9562,N_5491);
nor U10065 (N_10065,N_6992,N_5067);
nand U10066 (N_10066,N_5009,N_8841);
xor U10067 (N_10067,N_9003,N_9288);
and U10068 (N_10068,N_7557,N_6909);
nand U10069 (N_10069,N_6408,N_5478);
or U10070 (N_10070,N_9493,N_8073);
xnor U10071 (N_10071,N_9564,N_7316);
and U10072 (N_10072,N_7672,N_7511);
xnor U10073 (N_10073,N_6485,N_9608);
nand U10074 (N_10074,N_9396,N_6315);
xnor U10075 (N_10075,N_9940,N_8482);
nand U10076 (N_10076,N_7319,N_7488);
nand U10077 (N_10077,N_7583,N_5531);
or U10078 (N_10078,N_7160,N_7717);
nand U10079 (N_10079,N_5947,N_9654);
nand U10080 (N_10080,N_5162,N_7448);
nor U10081 (N_10081,N_8140,N_7167);
nor U10082 (N_10082,N_6418,N_8222);
or U10083 (N_10083,N_6121,N_9755);
xor U10084 (N_10084,N_8315,N_8254);
nand U10085 (N_10085,N_9964,N_9782);
or U10086 (N_10086,N_5367,N_7755);
or U10087 (N_10087,N_8761,N_9395);
nor U10088 (N_10088,N_9028,N_5257);
nand U10089 (N_10089,N_6788,N_5633);
xor U10090 (N_10090,N_6957,N_5026);
and U10091 (N_10091,N_9898,N_6583);
xnor U10092 (N_10092,N_8271,N_9868);
or U10093 (N_10093,N_9599,N_7283);
nor U10094 (N_10094,N_8246,N_9587);
or U10095 (N_10095,N_6354,N_5085);
nor U10096 (N_10096,N_9511,N_7453);
nand U10097 (N_10097,N_6251,N_6516);
nand U10098 (N_10098,N_7282,N_9430);
nand U10099 (N_10099,N_7340,N_7406);
nand U10100 (N_10100,N_9647,N_8716);
nand U10101 (N_10101,N_8598,N_8901);
and U10102 (N_10102,N_6980,N_7663);
or U10103 (N_10103,N_6833,N_8683);
nor U10104 (N_10104,N_9066,N_8085);
nor U10105 (N_10105,N_7889,N_8800);
nand U10106 (N_10106,N_5135,N_7940);
nor U10107 (N_10107,N_6279,N_8426);
nor U10108 (N_10108,N_8104,N_5895);
nor U10109 (N_10109,N_6829,N_9121);
xnor U10110 (N_10110,N_6105,N_7301);
xor U10111 (N_10111,N_7744,N_8902);
xnor U10112 (N_10112,N_7915,N_7098);
nor U10113 (N_10113,N_7714,N_9317);
and U10114 (N_10114,N_5913,N_8945);
and U10115 (N_10115,N_6831,N_5352);
xnor U10116 (N_10116,N_7602,N_6358);
nand U10117 (N_10117,N_5774,N_8977);
nor U10118 (N_10118,N_8886,N_9723);
nand U10119 (N_10119,N_6657,N_5368);
and U10120 (N_10120,N_6772,N_8708);
nand U10121 (N_10121,N_7165,N_8014);
nor U10122 (N_10122,N_8102,N_7431);
xnor U10123 (N_10123,N_8988,N_8510);
nand U10124 (N_10124,N_5045,N_6038);
nor U10125 (N_10125,N_7155,N_9744);
nand U10126 (N_10126,N_7025,N_9385);
and U10127 (N_10127,N_6119,N_6386);
nand U10128 (N_10128,N_5056,N_5349);
and U10129 (N_10129,N_9716,N_8590);
or U10130 (N_10130,N_8488,N_8508);
or U10131 (N_10131,N_8388,N_7484);
or U10132 (N_10132,N_7433,N_5568);
xnor U10133 (N_10133,N_6497,N_8161);
nand U10134 (N_10134,N_7849,N_6515);
xnor U10135 (N_10135,N_8259,N_9325);
and U10136 (N_10136,N_6940,N_8791);
nand U10137 (N_10137,N_5951,N_5767);
nor U10138 (N_10138,N_6009,N_6197);
and U10139 (N_10139,N_8998,N_6341);
and U10140 (N_10140,N_9155,N_6474);
or U10141 (N_10141,N_5033,N_9078);
xnor U10142 (N_10142,N_9766,N_6619);
or U10143 (N_10143,N_5459,N_7123);
or U10144 (N_10144,N_9369,N_5603);
nand U10145 (N_10145,N_8642,N_9830);
nand U10146 (N_10146,N_6577,N_6822);
or U10147 (N_10147,N_6417,N_5208);
or U10148 (N_10148,N_9368,N_5207);
nand U10149 (N_10149,N_5647,N_6546);
nand U10150 (N_10150,N_7410,N_9201);
and U10151 (N_10151,N_9565,N_8267);
nor U10152 (N_10152,N_9532,N_6364);
or U10153 (N_10153,N_9153,N_6228);
and U10154 (N_10154,N_8261,N_8826);
or U10155 (N_10155,N_8003,N_5991);
xor U10156 (N_10156,N_9409,N_5835);
or U10157 (N_10157,N_6384,N_9415);
nand U10158 (N_10158,N_6263,N_9033);
or U10159 (N_10159,N_5403,N_7383);
xor U10160 (N_10160,N_6544,N_8145);
or U10161 (N_10161,N_6804,N_7682);
or U10162 (N_10162,N_6131,N_7240);
xnor U10163 (N_10163,N_9949,N_5743);
nor U10164 (N_10164,N_5004,N_9135);
and U10165 (N_10165,N_8965,N_8193);
xnor U10166 (N_10166,N_6265,N_6355);
nand U10167 (N_10167,N_9287,N_8395);
or U10168 (N_10168,N_9476,N_9275);
or U10169 (N_10169,N_6499,N_7416);
or U10170 (N_10170,N_5635,N_8017);
nor U10171 (N_10171,N_9240,N_5016);
xnor U10172 (N_10172,N_6313,N_5866);
xnor U10173 (N_10173,N_9579,N_6893);
nand U10174 (N_10174,N_7062,N_7959);
and U10175 (N_10175,N_9765,N_9259);
nor U10176 (N_10176,N_6343,N_9825);
or U10177 (N_10177,N_7088,N_7845);
and U10178 (N_10178,N_8566,N_5784);
and U10179 (N_10179,N_6588,N_6624);
or U10180 (N_10180,N_7960,N_6304);
xnor U10181 (N_10181,N_9359,N_6334);
and U10182 (N_10182,N_9478,N_7753);
nor U10183 (N_10183,N_6853,N_9453);
and U10184 (N_10184,N_5453,N_6168);
xnor U10185 (N_10185,N_9932,N_6792);
xor U10186 (N_10186,N_9205,N_5267);
and U10187 (N_10187,N_6441,N_5260);
xor U10188 (N_10188,N_7956,N_9618);
or U10189 (N_10189,N_8435,N_8318);
nor U10190 (N_10190,N_8404,N_5676);
or U10191 (N_10191,N_8932,N_5410);
and U10192 (N_10192,N_5668,N_7273);
and U10193 (N_10193,N_5830,N_5671);
xnor U10194 (N_10194,N_5831,N_9538);
nand U10195 (N_10195,N_5732,N_5855);
or U10196 (N_10196,N_7162,N_9590);
or U10197 (N_10197,N_7541,N_6784);
or U10198 (N_10198,N_7379,N_7661);
nor U10199 (N_10199,N_8202,N_9786);
nand U10200 (N_10200,N_9521,N_6953);
nand U10201 (N_10201,N_7859,N_9805);
nand U10202 (N_10202,N_6642,N_6936);
xor U10203 (N_10203,N_5513,N_9530);
and U10204 (N_10204,N_8814,N_6808);
xor U10205 (N_10205,N_7445,N_7730);
or U10206 (N_10206,N_8353,N_9892);
xnor U10207 (N_10207,N_8679,N_6646);
xnor U10208 (N_10208,N_5418,N_5896);
xnor U10209 (N_10209,N_8281,N_8580);
or U10210 (N_10210,N_7260,N_6430);
xor U10211 (N_10211,N_9733,N_8991);
nor U10212 (N_10212,N_6938,N_8136);
and U10213 (N_10213,N_6215,N_6400);
nand U10214 (N_10214,N_7822,N_9620);
nor U10215 (N_10215,N_7352,N_5870);
and U10216 (N_10216,N_5847,N_7177);
or U10217 (N_10217,N_6285,N_9136);
or U10218 (N_10218,N_6634,N_8074);
and U10219 (N_10219,N_7080,N_5003);
nor U10220 (N_10220,N_9228,N_9421);
nand U10221 (N_10221,N_7141,N_8499);
or U10222 (N_10222,N_5193,N_7650);
or U10223 (N_10223,N_8049,N_7110);
and U10224 (N_10224,N_6326,N_5493);
nand U10225 (N_10225,N_8450,N_9172);
and U10226 (N_10226,N_9137,N_6017);
or U10227 (N_10227,N_5219,N_7315);
xnor U10228 (N_10228,N_7462,N_9920);
nor U10229 (N_10229,N_7142,N_5609);
xnor U10230 (N_10230,N_5702,N_7997);
and U10231 (N_10231,N_9206,N_5381);
and U10232 (N_10232,N_7144,N_9907);
xor U10233 (N_10233,N_8408,N_6359);
or U10234 (N_10234,N_8897,N_5355);
or U10235 (N_10235,N_8121,N_9074);
nand U10236 (N_10236,N_5249,N_5889);
nor U10237 (N_10237,N_7656,N_7351);
nor U10238 (N_10238,N_5443,N_9979);
and U10239 (N_10239,N_8111,N_9413);
xor U10240 (N_10240,N_5482,N_8564);
nand U10241 (N_10241,N_8715,N_5894);
nor U10242 (N_10242,N_8782,N_8702);
nand U10243 (N_10243,N_7318,N_7811);
nand U10244 (N_10244,N_6950,N_8024);
nand U10245 (N_10245,N_9473,N_8867);
or U10246 (N_10246,N_6594,N_5999);
or U10247 (N_10247,N_5426,N_9732);
nor U10248 (N_10248,N_5867,N_8703);
xor U10249 (N_10249,N_7314,N_5992);
or U10250 (N_10250,N_9827,N_5806);
or U10251 (N_10251,N_6541,N_6719);
or U10252 (N_10252,N_5018,N_6186);
xor U10253 (N_10253,N_6450,N_7862);
and U10254 (N_10254,N_8002,N_7291);
nor U10255 (N_10255,N_6760,N_8987);
nand U10256 (N_10256,N_5815,N_5522);
xnor U10257 (N_10257,N_7514,N_9635);
nand U10258 (N_10258,N_8106,N_9048);
nand U10259 (N_10259,N_7373,N_5321);
and U10260 (N_10260,N_6231,N_7148);
nand U10261 (N_10261,N_9953,N_8864);
and U10262 (N_10262,N_7872,N_9375);
nor U10263 (N_10263,N_5632,N_7976);
or U10264 (N_10264,N_6060,N_7085);
and U10265 (N_10265,N_6370,N_7636);
or U10266 (N_10266,N_6026,N_5494);
and U10267 (N_10267,N_9310,N_9380);
or U10268 (N_10268,N_6543,N_8176);
nand U10269 (N_10269,N_8997,N_9016);
xnor U10270 (N_10270,N_6380,N_9986);
and U10271 (N_10271,N_6563,N_5254);
and U10272 (N_10272,N_9864,N_5606);
xor U10273 (N_10273,N_8609,N_8755);
nand U10274 (N_10274,N_8075,N_6557);
nand U10275 (N_10275,N_5988,N_5570);
and U10276 (N_10276,N_7800,N_6698);
nand U10277 (N_10277,N_7528,N_9961);
nand U10278 (N_10278,N_9642,N_8393);
xnor U10279 (N_10279,N_9001,N_8554);
nand U10280 (N_10280,N_5837,N_8801);
nor U10281 (N_10281,N_8342,N_6420);
xnor U10282 (N_10282,N_5087,N_9768);
or U10283 (N_10283,N_6658,N_9073);
and U10284 (N_10284,N_6434,N_6129);
xor U10285 (N_10285,N_8718,N_6429);
and U10286 (N_10286,N_8043,N_6495);
and U10287 (N_10287,N_8096,N_9952);
nor U10288 (N_10288,N_5518,N_5472);
xnor U10289 (N_10289,N_9861,N_5339);
nor U10290 (N_10290,N_8006,N_9634);
nor U10291 (N_10291,N_6649,N_7863);
nand U10292 (N_10292,N_7560,N_6564);
or U10293 (N_10293,N_8175,N_7640);
nor U10294 (N_10294,N_9251,N_5042);
and U10295 (N_10295,N_9992,N_5032);
xor U10296 (N_10296,N_7545,N_5585);
and U10297 (N_10297,N_5445,N_9331);
and U10298 (N_10298,N_8407,N_5178);
or U10299 (N_10299,N_6133,N_6989);
xor U10300 (N_10300,N_5083,N_7612);
or U10301 (N_10301,N_7591,N_5943);
nor U10302 (N_10302,N_7215,N_7841);
nor U10303 (N_10303,N_6640,N_9116);
xnor U10304 (N_10304,N_7797,N_9707);
xor U10305 (N_10305,N_9867,N_9609);
nand U10306 (N_10306,N_6751,N_5102);
nand U10307 (N_10307,N_8960,N_8210);
or U10308 (N_10308,N_9728,N_8636);
and U10309 (N_10309,N_9687,N_9708);
or U10310 (N_10310,N_7206,N_8798);
and U10311 (N_10311,N_8836,N_9281);
nor U10312 (N_10312,N_9110,N_9710);
xor U10313 (N_10313,N_8011,N_8904);
nor U10314 (N_10314,N_7227,N_6740);
nand U10315 (N_10315,N_7257,N_6138);
nor U10316 (N_10316,N_5383,N_8078);
xor U10317 (N_10317,N_6725,N_9485);
and U10318 (N_10318,N_9851,N_5353);
xor U10319 (N_10319,N_9556,N_8649);
nor U10320 (N_10320,N_5414,N_7712);
nand U10321 (N_10321,N_6072,N_5678);
and U10322 (N_10322,N_7270,N_9333);
and U10323 (N_10323,N_5558,N_6084);
nand U10324 (N_10324,N_8691,N_8010);
xor U10325 (N_10325,N_5184,N_7665);
and U10326 (N_10326,N_6378,N_5869);
or U10327 (N_10327,N_5496,N_5820);
or U10328 (N_10328,N_6741,N_9462);
nand U10329 (N_10329,N_8628,N_7306);
and U10330 (N_10330,N_8741,N_5460);
and U10331 (N_10331,N_9122,N_8115);
nor U10332 (N_10332,N_9307,N_5757);
or U10333 (N_10333,N_6742,N_5465);
nand U10334 (N_10334,N_9420,N_6502);
and U10335 (N_10335,N_9872,N_6127);
nand U10336 (N_10336,N_9436,N_5680);
and U10337 (N_10337,N_8746,N_8548);
and U10338 (N_10338,N_6510,N_8107);
nor U10339 (N_10339,N_5366,N_5299);
and U10340 (N_10340,N_7829,N_9810);
and U10341 (N_10341,N_5270,N_5529);
nor U10342 (N_10342,N_6030,N_6666);
nor U10343 (N_10343,N_5323,N_9736);
nor U10344 (N_10344,N_8059,N_8976);
nor U10345 (N_10345,N_8958,N_8500);
nor U10346 (N_10346,N_8532,N_8866);
nor U10347 (N_10347,N_6365,N_7212);
xor U10348 (N_10348,N_9603,N_7197);
nand U10349 (N_10349,N_6551,N_8039);
nand U10350 (N_10350,N_7087,N_6726);
nor U10351 (N_10351,N_8432,N_5822);
or U10352 (N_10352,N_6880,N_9551);
nand U10353 (N_10353,N_9966,N_8521);
or U10354 (N_10354,N_8335,N_7895);
nand U10355 (N_10355,N_9871,N_8764);
xor U10356 (N_10356,N_8982,N_5521);
and U10357 (N_10357,N_9541,N_5338);
or U10358 (N_10358,N_9491,N_5780);
xnor U10359 (N_10359,N_7159,N_7440);
or U10360 (N_10360,N_8947,N_5662);
nand U10361 (N_10361,N_6278,N_7733);
or U10362 (N_10362,N_9311,N_8151);
nor U10363 (N_10363,N_7266,N_8112);
and U10364 (N_10364,N_8612,N_8617);
or U10365 (N_10365,N_9247,N_8912);
nor U10366 (N_10366,N_6656,N_6273);
nor U10367 (N_10367,N_5454,N_6071);
nand U10368 (N_10368,N_9548,N_5150);
nor U10369 (N_10369,N_6689,N_9486);
nand U10370 (N_10370,N_7140,N_9046);
xor U10371 (N_10371,N_6514,N_9301);
nor U10372 (N_10372,N_8348,N_7043);
or U10373 (N_10373,N_9831,N_8633);
nor U10374 (N_10374,N_7219,N_9580);
xor U10375 (N_10375,N_5498,N_5995);
and U10376 (N_10376,N_5181,N_7920);
nand U10377 (N_10377,N_9350,N_7499);
xor U10378 (N_10378,N_6043,N_6990);
xor U10379 (N_10379,N_5886,N_7300);
nor U10380 (N_10380,N_9094,N_6196);
xnor U10381 (N_10381,N_5629,N_6211);
nand U10382 (N_10382,N_5579,N_6046);
xor U10383 (N_10383,N_7641,N_8607);
xor U10384 (N_10384,N_7923,N_7883);
nor U10385 (N_10385,N_5956,N_5619);
and U10386 (N_10386,N_5595,N_8084);
xor U10387 (N_10387,N_9455,N_6633);
nor U10388 (N_10388,N_8667,N_5389);
nor U10389 (N_10389,N_5242,N_9272);
or U10390 (N_10390,N_7563,N_5954);
and U10391 (N_10391,N_5564,N_7497);
xnor U10392 (N_10392,N_8457,N_8563);
and U10393 (N_10393,N_7540,N_6103);
or U10394 (N_10394,N_6991,N_8651);
nand U10395 (N_10395,N_5176,N_8870);
or U10396 (N_10396,N_9595,N_6750);
and U10397 (N_10397,N_5824,N_9584);
or U10398 (N_10398,N_5489,N_9132);
xor U10399 (N_10399,N_7093,N_8931);
or U10400 (N_10400,N_7361,N_5255);
or U10401 (N_10401,N_8955,N_6728);
or U10402 (N_10402,N_8778,N_8263);
xnor U10403 (N_10403,N_9925,N_5685);
and U10404 (N_10404,N_9559,N_8774);
nor U10405 (N_10405,N_8400,N_5206);
nor U10406 (N_10406,N_6120,N_8602);
xor U10407 (N_10407,N_7851,N_8226);
or U10408 (N_10408,N_5020,N_8961);
or U10409 (N_10409,N_8313,N_5014);
nor U10410 (N_10410,N_5024,N_5819);
nand U10411 (N_10411,N_9398,N_7426);
xnor U10412 (N_10412,N_5439,N_6224);
nor U10413 (N_10413,N_7624,N_5280);
and U10414 (N_10414,N_5654,N_7597);
and U10415 (N_10415,N_7741,N_5622);
nand U10416 (N_10416,N_7475,N_5795);
xnor U10417 (N_10417,N_5117,N_8295);
nand U10418 (N_10418,N_9169,N_8483);
and U10419 (N_10419,N_7222,N_5705);
xor U10420 (N_10420,N_6255,N_8661);
nor U10421 (N_10421,N_7395,N_6210);
xor U10422 (N_10422,N_7515,N_7450);
xnor U10423 (N_10423,N_5592,N_9522);
nand U10424 (N_10424,N_7824,N_6457);
nand U10425 (N_10425,N_9767,N_8734);
xnor U10426 (N_10426,N_9047,N_9139);
and U10427 (N_10427,N_6377,N_9295);
nor U10428 (N_10428,N_8093,N_9252);
and U10429 (N_10429,N_6931,N_8845);
nand U10430 (N_10430,N_9691,N_8700);
nand U10431 (N_10431,N_8317,N_9249);
and U10432 (N_10432,N_5311,N_7648);
and U10433 (N_10433,N_7983,N_5607);
and U10434 (N_10434,N_7603,N_6058);
or U10435 (N_10435,N_7150,N_7567);
and U10436 (N_10436,N_6855,N_6866);
xor U10437 (N_10437,N_6924,N_6353);
nand U10438 (N_10438,N_9335,N_8726);
nor U10439 (N_10439,N_7628,N_9390);
xor U10440 (N_10440,N_6040,N_9178);
or U10441 (N_10441,N_8098,N_7116);
nand U10442 (N_10442,N_9217,N_8105);
nor U10443 (N_10443,N_7616,N_5904);
or U10444 (N_10444,N_7226,N_5783);
xnor U10445 (N_10445,N_6972,N_8996);
and U10446 (N_10446,N_6444,N_5258);
nand U10447 (N_10447,N_8303,N_6047);
nand U10448 (N_10448,N_7573,N_9809);
or U10449 (N_10449,N_6768,N_9019);
xor U10450 (N_10450,N_9761,N_9013);
nor U10451 (N_10451,N_9214,N_5064);
xnor U10452 (N_10452,N_8561,N_6153);
nor U10453 (N_10453,N_5880,N_8637);
nand U10454 (N_10454,N_9890,N_8477);
nand U10455 (N_10455,N_7089,N_5615);
xnor U10456 (N_10456,N_5086,N_9026);
nor U10457 (N_10457,N_8230,N_7263);
nor U10458 (N_10458,N_6732,N_5958);
nor U10459 (N_10459,N_6714,N_8144);
nand U10460 (N_10460,N_9788,N_7680);
and U10461 (N_10461,N_9185,N_8777);
or U10462 (N_10462,N_6014,N_9915);
xnor U10463 (N_10463,N_7293,N_5183);
nand U10464 (N_10464,N_7008,N_8669);
or U10465 (N_10465,N_6065,N_6535);
xor U10466 (N_10466,N_9489,N_9397);
and U10467 (N_10467,N_9354,N_5745);
nor U10468 (N_10468,N_8126,N_8948);
nor U10469 (N_10469,N_8496,N_7936);
and U10470 (N_10470,N_9020,N_9746);
nand U10471 (N_10471,N_6117,N_6298);
or U10472 (N_10472,N_9082,N_8526);
or U10473 (N_10473,N_8273,N_9985);
xnor U10474 (N_10474,N_5427,N_9842);
xor U10475 (N_10475,N_7981,N_9106);
xor U10476 (N_10476,N_6948,N_8568);
and U10477 (N_10477,N_5985,N_8401);
nand U10478 (N_10478,N_5902,N_9146);
nor U10479 (N_10479,N_7265,N_9219);
nor U10480 (N_10480,N_7925,N_6109);
nand U10481 (N_10481,N_5111,N_7857);
nor U10482 (N_10482,N_7249,N_5799);
xnor U10483 (N_10483,N_6965,N_6975);
nand U10484 (N_10484,N_7117,N_9351);
nand U10485 (N_10485,N_8821,N_9488);
xnor U10486 (N_10486,N_5694,N_8635);
nand U10487 (N_10487,N_7667,N_7558);
nor U10488 (N_10488,N_6262,N_5508);
or U10489 (N_10489,N_8639,N_5306);
and U10490 (N_10490,N_7896,N_9895);
or U10491 (N_10491,N_6686,N_5005);
nand U10492 (N_10492,N_8124,N_9343);
nand U10493 (N_10493,N_7279,N_5081);
or U10494 (N_10494,N_7033,N_5126);
nand U10495 (N_10495,N_5773,N_6045);
nand U10496 (N_10496,N_7813,N_7871);
xor U10497 (N_10497,N_7035,N_6271);
and U10498 (N_10498,N_8489,N_5979);
or U10499 (N_10499,N_6289,N_9794);
xnor U10500 (N_10500,N_5666,N_8540);
or U10501 (N_10501,N_5912,N_7084);
and U10502 (N_10502,N_9757,N_7329);
and U10503 (N_10503,N_9948,N_6569);
and U10504 (N_10504,N_6591,N_5916);
nor U10505 (N_10505,N_6864,N_7646);
nor U10506 (N_10506,N_7012,N_8330);
xor U10507 (N_10507,N_9012,N_7761);
and U10508 (N_10508,N_8983,N_7169);
nand U10509 (N_10509,N_6521,N_6517);
nand U10510 (N_10510,N_9107,N_7028);
and U10511 (N_10511,N_5528,N_9523);
and U10512 (N_10512,N_6356,N_9705);
nor U10513 (N_10513,N_9837,N_8581);
and U10514 (N_10514,N_8707,N_6193);
xor U10515 (N_10515,N_6523,N_5631);
xnor U10516 (N_10516,N_9313,N_7452);
xnor U10517 (N_10517,N_9750,N_8507);
or U10518 (N_10518,N_8560,N_9089);
nor U10519 (N_10519,N_8614,N_5812);
or U10520 (N_10520,N_9246,N_5626);
xor U10521 (N_10521,N_6946,N_5698);
or U10522 (N_10522,N_5645,N_6021);
xor U10523 (N_10523,N_8027,N_9968);
nand U10524 (N_10524,N_7830,N_6886);
or U10525 (N_10525,N_8583,N_5423);
nand U10526 (N_10526,N_8621,N_8909);
xnor U10527 (N_10527,N_7600,N_7783);
nor U10528 (N_10528,N_9899,N_7326);
xnor U10529 (N_10529,N_8490,N_7136);
nor U10530 (N_10530,N_8422,N_9983);
or U10531 (N_10531,N_8156,N_6190);
xor U10532 (N_10532,N_9799,N_7498);
nand U10533 (N_10533,N_9939,N_7099);
xnor U10534 (N_10534,N_9652,N_5090);
nor U10535 (N_10535,N_8768,N_9936);
nand U10536 (N_10536,N_6887,N_8921);
and U10537 (N_10537,N_5834,N_7986);
and U10538 (N_10538,N_9515,N_9216);
or U10539 (N_10539,N_8837,N_9431);
xnor U10540 (N_10540,N_9083,N_8585);
xnor U10541 (N_10541,N_8148,N_8758);
nand U10542 (N_10542,N_9470,N_6696);
or U10543 (N_10543,N_5230,N_5089);
xnor U10544 (N_10544,N_8604,N_9129);
xnor U10545 (N_10545,N_9285,N_7097);
nor U10546 (N_10546,N_5511,N_6573);
and U10547 (N_10547,N_8062,N_7320);
or U10548 (N_10548,N_5017,N_7030);
xnor U10549 (N_10549,N_5112,N_5563);
and U10550 (N_10550,N_5200,N_9057);
xor U10551 (N_10551,N_6295,N_6707);
nand U10552 (N_10552,N_6501,N_6782);
and U10553 (N_10553,N_9265,N_9807);
or U10554 (N_10554,N_9043,N_6132);
or U10555 (N_10555,N_7930,N_9960);
or U10556 (N_10556,N_6362,N_8630);
nand U10557 (N_10557,N_7481,N_9576);
and U10558 (N_10558,N_5218,N_5091);
xor U10559 (N_10559,N_6079,N_5854);
nand U10560 (N_10560,N_7953,N_8249);
xor U10561 (N_10561,N_5105,N_6617);
and U10562 (N_10562,N_9248,N_5238);
and U10563 (N_10563,N_6100,N_9865);
xor U10564 (N_10564,N_7534,N_7942);
or U10565 (N_10565,N_6630,N_6919);
xor U10566 (N_10566,N_9798,N_6099);
or U10567 (N_10567,N_7360,N_6620);
and U10568 (N_10568,N_5620,N_8089);
or U10569 (N_10569,N_5139,N_8239);
and U10570 (N_10570,N_5010,N_5543);
or U10571 (N_10571,N_6200,N_5290);
or U10572 (N_10572,N_7806,N_8443);
nor U10573 (N_10573,N_9933,N_6963);
or U10574 (N_10574,N_9154,N_6220);
and U10575 (N_10575,N_7961,N_6054);
nand U10576 (N_10576,N_9506,N_6246);
nand U10577 (N_10577,N_5970,N_9574);
nand U10578 (N_10578,N_7460,N_5838);
nor U10579 (N_10579,N_9561,N_9404);
and U10580 (N_10580,N_8705,N_8659);
nand U10581 (N_10581,N_7223,N_5334);
nand U10582 (N_10582,N_7304,N_6253);
or U10583 (N_10583,N_5037,N_6242);
and U10584 (N_10584,N_6667,N_8171);
and U10585 (N_10585,N_6459,N_8168);
nand U10586 (N_10586,N_8037,N_6773);
nand U10587 (N_10587,N_7707,N_8858);
xor U10588 (N_10588,N_9338,N_5118);
nor U10589 (N_10589,N_6394,N_5331);
or U10590 (N_10590,N_8131,N_5068);
nor U10591 (N_10591,N_8654,N_5739);
and U10592 (N_10592,N_9682,N_5289);
and U10593 (N_10593,N_8862,N_5533);
and U10594 (N_10594,N_6881,N_5524);
nand U10595 (N_10595,N_5481,N_7173);
xnor U10596 (N_10596,N_8589,N_6934);
or U10597 (N_10597,N_5076,N_8423);
xnor U10598 (N_10598,N_8600,N_8190);
nand U10599 (N_10599,N_7978,N_9414);
or U10600 (N_10600,N_5398,N_5480);
or U10601 (N_10601,N_8257,N_9223);
nand U10602 (N_10602,N_5818,N_6427);
or U10603 (N_10603,N_5177,N_5397);
xor U10604 (N_10604,N_5723,N_7516);
nor U10605 (N_10605,N_7585,N_6456);
and U10606 (N_10606,N_8357,N_5373);
nand U10607 (N_10607,N_7500,N_5315);
nor U10608 (N_10608,N_9834,N_8584);
nor U10609 (N_10609,N_9622,N_6974);
nor U10610 (N_10610,N_7924,N_7193);
nand U10611 (N_10611,N_7539,N_8812);
nor U10612 (N_10612,N_6063,N_5247);
or U10613 (N_10613,N_5237,N_5706);
nand U10614 (N_10614,N_8750,N_7446);
nor U10615 (N_10615,N_8325,N_9922);
nand U10616 (N_10616,N_9261,N_8544);
xor U10617 (N_10617,N_6440,N_5608);
or U10618 (N_10618,N_6366,N_8695);
nand U10619 (N_10619,N_9813,N_5225);
and U10620 (N_10620,N_6241,N_9850);
xor U10621 (N_10621,N_8418,N_6643);
or U10622 (N_10622,N_9832,N_6282);
nor U10623 (N_10623,N_9854,N_7673);
xnor U10624 (N_10624,N_8201,N_5725);
and U10625 (N_10625,N_6811,N_6314);
xor U10626 (N_10626,N_6303,N_7899);
nand U10627 (N_10627,N_8898,N_7425);
nand U10628 (N_10628,N_7066,N_6202);
and U10629 (N_10629,N_5013,N_8398);
and U10630 (N_10630,N_7346,N_9916);
and U10631 (N_10631,N_8293,N_9339);
xor U10632 (N_10632,N_9027,N_5340);
or U10633 (N_10633,N_9802,N_6381);
nand U10634 (N_10634,N_6672,N_7552);
or U10635 (N_10635,N_6256,N_5240);
xor U10636 (N_10636,N_5930,N_9918);
and U10637 (N_10637,N_6488,N_5817);
and U10638 (N_10638,N_5600,N_6536);
or U10639 (N_10639,N_5569,N_6402);
or U10640 (N_10640,N_8433,N_7011);
or U10641 (N_10641,N_9748,N_9475);
nor U10642 (N_10642,N_7258,N_8546);
xnor U10643 (N_10643,N_9034,N_9144);
xnor U10644 (N_10644,N_5914,N_7589);
nand U10645 (N_10645,N_7781,N_5516);
and U10646 (N_10646,N_5634,N_7653);
nand U10647 (N_10647,N_5034,N_8658);
nor U10648 (N_10648,N_8974,N_5848);
nand U10649 (N_10649,N_8877,N_7432);
and U10650 (N_10650,N_5450,N_5798);
and U10651 (N_10651,N_9023,N_7359);
nand U10652 (N_10652,N_7635,N_7613);
xnor U10653 (N_10653,N_8882,N_5874);
and U10654 (N_10654,N_8941,N_6821);
xnor U10655 (N_10655,N_9015,N_6678);
nand U10656 (N_10656,N_8539,N_7568);
nand U10657 (N_10657,N_9243,N_8294);
or U10658 (N_10658,N_8420,N_6392);
or U10659 (N_10659,N_7838,N_8405);
or U10660 (N_10660,N_8459,N_6654);
nand U10661 (N_10661,N_5501,N_8818);
and U10662 (N_10662,N_8493,N_7137);
and U10663 (N_10663,N_5604,N_8735);
nand U10664 (N_10664,N_6906,N_9292);
or U10665 (N_10665,N_6415,N_9008);
and U10666 (N_10666,N_7947,N_9007);
xor U10667 (N_10667,N_5517,N_6452);
or U10668 (N_10668,N_9712,N_7877);
nor U10669 (N_10669,N_8926,N_7700);
and U10670 (N_10670,N_5714,N_7518);
nor U10671 (N_10671,N_5119,N_7536);
and U10672 (N_10672,N_6664,N_9648);
nand U10673 (N_10673,N_9076,N_5591);
xor U10674 (N_10674,N_8306,N_8476);
nor U10675 (N_10675,N_7074,N_5399);
and U10676 (N_10676,N_7120,N_6602);
nand U10677 (N_10677,N_9318,N_7396);
or U10678 (N_10678,N_7928,N_9014);
or U10679 (N_10679,N_5424,N_8200);
or U10680 (N_10680,N_5094,N_6306);
or U10681 (N_10681,N_8032,N_9226);
or U10682 (N_10682,N_7009,N_6307);
nand U10683 (N_10683,N_8615,N_6397);
xor U10684 (N_10684,N_8973,N_5507);
nor U10685 (N_10685,N_8786,N_7145);
and U10686 (N_10686,N_7397,N_5268);
and U10687 (N_10687,N_5394,N_6983);
xnor U10688 (N_10688,N_6425,N_5605);
nor U10689 (N_10689,N_7581,N_7311);
or U10690 (N_10690,N_5222,N_6223);
or U10691 (N_10691,N_6128,N_8822);
xor U10692 (N_10692,N_7517,N_9194);
and U10693 (N_10693,N_8248,N_9588);
nor U10694 (N_10694,N_5807,N_7281);
or U10695 (N_10695,N_5314,N_9969);
xor U10696 (N_10696,N_8354,N_8284);
nand U10697 (N_10697,N_6102,N_6042);
and U10698 (N_10698,N_5565,N_7578);
or U10699 (N_10699,N_9077,N_6093);
or U10700 (N_10700,N_7269,N_7627);
and U10701 (N_10701,N_7449,N_6824);
and U10702 (N_10702,N_7691,N_9602);
nand U10703 (N_10703,N_6130,N_6874);
nor U10704 (N_10704,N_7241,N_7236);
xnor U10705 (N_10705,N_7584,N_9617);
or U10706 (N_10706,N_7428,N_9257);
and U10707 (N_10707,N_7071,N_5859);
nand U10708 (N_10708,N_8238,N_8403);
nor U10709 (N_10709,N_7245,N_6181);
and U10710 (N_10710,N_7023,N_5216);
or U10711 (N_10711,N_6739,N_6051);
nand U10712 (N_10712,N_5862,N_6280);
xor U10713 (N_10713,N_7503,N_6807);
and U10714 (N_10714,N_6865,N_7693);
xor U10715 (N_10715,N_9504,N_5277);
nand U10716 (N_10716,N_9773,N_7494);
nor U10717 (N_10717,N_6540,N_9653);
xor U10718 (N_10718,N_9616,N_7743);
xor U10719 (N_10719,N_5652,N_5214);
or U10720 (N_10720,N_6652,N_9514);
nand U10721 (N_10721,N_5163,N_8298);
or U10722 (N_10722,N_9601,N_9993);
nand U10723 (N_10723,N_8095,N_6013);
and U10724 (N_10724,N_7436,N_5096);
nor U10725 (N_10725,N_7569,N_8344);
or U10726 (N_10726,N_5814,N_9469);
xnor U10727 (N_10727,N_9167,N_8397);
nand U10728 (N_10728,N_7525,N_5011);
or U10729 (N_10729,N_5527,N_5396);
nand U10730 (N_10730,N_9161,N_6873);
or U10731 (N_10731,N_8101,N_8687);
xnor U10732 (N_10732,N_9381,N_9179);
or U10733 (N_10733,N_7399,N_8260);
nand U10734 (N_10734,N_9378,N_7026);
nor U10735 (N_10735,N_6576,N_5582);
and U10736 (N_10736,N_9625,N_5993);
xnor U10737 (N_10737,N_7632,N_7732);
or U10738 (N_10738,N_5552,N_6631);
nor U10739 (N_10739,N_9729,N_8380);
nor U10740 (N_10740,N_7742,N_6482);
nor U10741 (N_10741,N_6311,N_7553);
and U10742 (N_10742,N_5982,N_9545);
or U10743 (N_10743,N_9394,N_8601);
and U10744 (N_10744,N_7772,N_8894);
or U10745 (N_10745,N_7119,N_7919);
xnor U10746 (N_10746,N_7100,N_7621);
and U10747 (N_10747,N_9447,N_8378);
nor U10748 (N_10748,N_5036,N_7343);
nor U10749 (N_10749,N_7655,N_6695);
xor U10750 (N_10750,N_6124,N_8371);
nor U10751 (N_10751,N_8185,N_8276);
and U10752 (N_10752,N_8738,N_7056);
nand U10753 (N_10753,N_5746,N_9693);
nor U10754 (N_10754,N_9720,N_9816);
and U10755 (N_10755,N_5946,N_7404);
nand U10756 (N_10756,N_6235,N_8883);
xor U10757 (N_10757,N_7766,N_6572);
nor U10758 (N_10758,N_5180,N_7782);
xnor U10759 (N_10759,N_5121,N_6943);
nor U10760 (N_10760,N_8183,N_6538);
nand U10761 (N_10761,N_7413,N_6146);
xor U10762 (N_10762,N_8130,N_5878);
and U10763 (N_10763,N_9100,N_7192);
or U10764 (N_10764,N_8964,N_9908);
nand U10765 (N_10765,N_9158,N_6592);
nand U10766 (N_10766,N_6891,N_6858);
or U10767 (N_10767,N_5342,N_9422);
and U10768 (N_10768,N_5079,N_5243);
xor U10769 (N_10769,N_7363,N_7409);
xnor U10770 (N_10770,N_7952,N_8724);
nand U10771 (N_10771,N_8460,N_8848);
and U10772 (N_10772,N_7046,N_8219);
or U10773 (N_10773,N_7414,N_9702);
and U10774 (N_10774,N_5244,N_9600);
or U10775 (N_10775,N_8656,N_5048);
nand U10776 (N_10776,N_6426,N_8929);
or U10777 (N_10777,N_8142,N_5054);
nor U10778 (N_10778,N_5695,N_6222);
and U10779 (N_10779,N_9051,N_6559);
xor U10780 (N_10780,N_9342,N_5341);
or U10781 (N_10781,N_8036,N_7962);
or U10782 (N_10782,N_7190,N_9142);
nand U10783 (N_10783,N_5312,N_5590);
or U10784 (N_10784,N_5857,N_9297);
xor U10785 (N_10785,N_5644,N_9466);
nand U10786 (N_10786,N_7096,N_8216);
xor U10787 (N_10787,N_7587,N_9306);
and U10788 (N_10788,N_9722,N_7681);
and U10789 (N_10789,N_5316,N_9124);
or U10790 (N_10790,N_5209,N_9108);
xor U10791 (N_10791,N_9518,N_5161);
xor U10792 (N_10792,N_8088,N_7729);
and U10793 (N_10793,N_6083,N_8299);
nand U10794 (N_10794,N_6173,N_8307);
nor U10795 (N_10795,N_8531,N_6977);
and U10796 (N_10796,N_6175,N_6323);
nand U10797 (N_10797,N_9875,N_8542);
or U10798 (N_10798,N_9965,N_9357);
xnor U10799 (N_10799,N_7971,N_7055);
and U10800 (N_10800,N_7507,N_6399);
xor U10801 (N_10801,N_5917,N_5891);
xnor U10802 (N_10802,N_8890,N_7284);
and U10803 (N_10803,N_6711,N_5264);
or U10804 (N_10804,N_9147,N_7831);
xnor U10805 (N_10805,N_9593,N_9134);
nor U10806 (N_10806,N_8872,N_8100);
or U10807 (N_10807,N_6140,N_8285);
nor U10808 (N_10808,N_7454,N_5365);
nand U10809 (N_10809,N_5672,N_6023);
nor U10810 (N_10810,N_8158,N_9010);
or U10811 (N_10811,N_5541,N_9069);
and U10812 (N_10812,N_7495,N_8368);
or U10813 (N_10813,N_8569,N_5444);
nand U10814 (N_10814,N_7228,N_8180);
and U10815 (N_10815,N_9709,N_5546);
and U10816 (N_10816,N_9471,N_5813);
and U10817 (N_10817,N_9157,N_7521);
or U10818 (N_10818,N_9340,N_8910);
or U10819 (N_10819,N_5567,N_8984);
or U10820 (N_10820,N_6027,N_6776);
and U10821 (N_10821,N_7463,N_8759);
and U10822 (N_10822,N_9484,N_5259);
or U10823 (N_10823,N_8928,N_6094);
or U10824 (N_10824,N_7734,N_7135);
nand U10825 (N_10825,N_8629,N_9065);
xor U10826 (N_10826,N_6688,N_7234);
xnor U10827 (N_10827,N_5358,N_7286);
nor U10828 (N_10828,N_9283,N_6840);
nor U10829 (N_10829,N_6478,N_5675);
nand U10830 (N_10830,N_9856,N_7353);
or U10831 (N_10831,N_8337,N_7985);
and U10832 (N_10832,N_6997,N_9649);
or U10833 (N_10833,N_9995,N_8513);
nand U10834 (N_10834,N_5274,N_5978);
nor U10835 (N_10835,N_9187,N_7607);
or U10836 (N_10836,N_7842,N_6309);
nand U10837 (N_10837,N_9423,N_6677);
or U10838 (N_10838,N_5069,N_6861);
xnor U10839 (N_10839,N_7917,N_6937);
and U10840 (N_10840,N_5287,N_8213);
or U10841 (N_10841,N_8714,N_9743);
and U10842 (N_10842,N_9118,N_5642);
xnor U10843 (N_10843,N_7562,N_6762);
nand U10844 (N_10844,N_5545,N_8773);
and U10845 (N_10845,N_8099,N_5972);
or U10846 (N_10846,N_7828,N_8680);
nor U10847 (N_10847,N_6275,N_6025);
xor U10848 (N_10848,N_9909,N_9688);
nand U10849 (N_10849,N_7417,N_5653);
nor U10850 (N_10850,N_7214,N_9889);
nor U10851 (N_10851,N_8813,N_7081);
xnor U10852 (N_10852,N_5787,N_5170);
nand U10853 (N_10853,N_8744,N_9527);
xnor U10854 (N_10854,N_7041,N_7061);
nor U10855 (N_10855,N_9321,N_8192);
and U10856 (N_10856,N_5015,N_6590);
or U10857 (N_10857,N_6151,N_8944);
nor U10858 (N_10858,N_8135,N_8456);
and U10859 (N_10859,N_6761,N_7032);
nor U10860 (N_10860,N_8366,N_8824);
xor U10861 (N_10861,N_7021,N_9668);
nand U10862 (N_10862,N_7188,N_5664);
xor U10863 (N_10863,N_7262,N_8040);
nand U10864 (N_10864,N_5228,N_7076);
xor U10865 (N_10865,N_7690,N_9882);
xor U10866 (N_10866,N_6383,N_9598);
xnor U10867 (N_10867,N_5899,N_8301);
nand U10868 (N_10868,N_5486,N_7237);
and U10869 (N_10869,N_5327,N_9542);
or U10870 (N_10870,N_8109,N_5175);
nand U10871 (N_10871,N_6092,N_9156);
nor U10872 (N_10872,N_8365,N_9245);
and U10873 (N_10873,N_8349,N_6316);
nor U10874 (N_10874,N_5893,N_9557);
nand U10875 (N_10875,N_9769,N_7605);
nand U10876 (N_10876,N_5580,N_6823);
nor U10877 (N_10877,N_7309,N_6789);
xor U10878 (N_10878,N_7143,N_7256);
xnor U10879 (N_10879,N_5760,N_9539);
xor U10880 (N_10880,N_6421,N_7934);
and U10881 (N_10881,N_8729,N_9192);
nor U10882 (N_10882,N_8536,N_6797);
nand U10883 (N_10883,N_8339,N_5971);
nor U10884 (N_10884,N_7598,N_6238);
xor U10885 (N_10885,N_5884,N_8925);
nor U10886 (N_10886,N_5292,N_8370);
nor U10887 (N_10887,N_5597,N_7465);
or U10888 (N_10888,N_7336,N_5473);
or U10889 (N_10889,N_6096,N_6185);
nand U10890 (N_10890,N_7054,N_6606);
nand U10891 (N_10891,N_5194,N_8184);
nor U10892 (N_10892,N_8939,N_6661);
and U10893 (N_10893,N_5770,N_6174);
xor U10894 (N_10894,N_6288,N_6160);
nand U10895 (N_10895,N_8772,N_7659);
nor U10896 (N_10896,N_8859,N_7748);
xor U10897 (N_10897,N_7386,N_5802);
or U10898 (N_10898,N_6684,N_6860);
nand U10899 (N_10899,N_6645,N_7713);
and U10900 (N_10900,N_9817,N_5198);
nand U10901 (N_10901,N_5278,N_6328);
and U10902 (N_10902,N_8305,N_7157);
and U10903 (N_10903,N_6428,N_9163);
or U10904 (N_10904,N_9808,N_9897);
or U10905 (N_10905,N_7550,N_8570);
nor U10906 (N_10906,N_8068,N_6056);
and U10907 (N_10907,N_9571,N_5966);
nand U10908 (N_10908,N_8831,N_5925);
or U10909 (N_10909,N_7651,N_5553);
nor U10910 (N_10910,N_7687,N_6746);
nor U10911 (N_10911,N_7182,N_5440);
xnor U10912 (N_10912,N_8058,N_7196);
nand U10913 (N_10913,N_9209,N_8103);
nand U10914 (N_10914,N_9718,N_9572);
or U10915 (N_10915,N_8653,N_5095);
or U10916 (N_10916,N_9316,N_9800);
nor U10917 (N_10917,N_6527,N_7357);
nand U10918 (N_10918,N_8162,N_7790);
nor U10919 (N_10919,N_9513,N_9823);
xor U10920 (N_10920,N_7331,N_7101);
and U10921 (N_10921,N_7795,N_8994);
nand U10922 (N_10922,N_8847,N_8215);
or U10923 (N_10923,N_7106,N_7348);
nor U10924 (N_10924,N_5758,N_8465);
and U10925 (N_10925,N_9719,N_8753);
nor U10926 (N_10926,N_8582,N_7235);
and U10927 (N_10927,N_7114,N_6187);
and U10928 (N_10928,N_8914,N_6737);
and U10929 (N_10929,N_5195,N_7754);
xor U10930 (N_10930,N_6916,N_9271);
nand U10931 (N_10931,N_8447,N_6537);
nor U10932 (N_10932,N_6312,N_5682);
xor U10933 (N_10933,N_8993,N_5151);
nor U10934 (N_10934,N_5266,N_6467);
and U10935 (N_10935,N_9399,N_6812);
nand U10936 (N_10936,N_8878,N_5976);
nor U10937 (N_10937,N_6333,N_7303);
nor U10938 (N_10938,N_5939,N_5159);
nor U10939 (N_10939,N_8529,N_7161);
nand U10940 (N_10940,N_5863,N_5602);
xor U10941 (N_10941,N_6115,N_8979);
xnor U10942 (N_10942,N_6795,N_9703);
nand U10943 (N_10943,N_6783,N_9268);
nand U10944 (N_10944,N_8900,N_5656);
or U10945 (N_10945,N_6844,N_6942);
xor U10946 (N_10946,N_9018,N_8511);
xor U10947 (N_10947,N_5960,N_6139);
xnor U10948 (N_10948,N_8916,N_8278);
and U10949 (N_10949,N_8379,N_5578);
nor U10950 (N_10950,N_5955,N_9432);
and U10951 (N_10951,N_9869,N_5326);
nand U10952 (N_10952,N_5104,N_8070);
and U10953 (N_10953,N_9623,N_9406);
xor U10954 (N_10954,N_8429,N_5663);
or U10955 (N_10955,N_6952,N_7933);
nor U10956 (N_10956,N_7869,N_8072);
nor U10957 (N_10957,N_8906,N_5182);
nand U10958 (N_10958,N_8415,N_5070);
xor U10959 (N_10959,N_8954,N_7296);
or U10960 (N_10960,N_5300,N_8056);
nand U10961 (N_10961,N_8364,N_7519);
nand U10962 (N_10962,N_8747,N_5729);
xor U10963 (N_10963,N_9727,N_8911);
and U10964 (N_10964,N_6925,N_7617);
or U10965 (N_10965,N_6987,N_9190);
or U10966 (N_10966,N_8587,N_7756);
nand U10967 (N_10967,N_5897,N_7954);
and U10968 (N_10968,N_9697,N_5957);
and U10969 (N_10969,N_8711,N_7823);
and U10970 (N_10970,N_9130,N_6321);
nand U10971 (N_10971,N_5092,N_9627);
or U10972 (N_10972,N_6396,N_6061);
nor U10973 (N_10973,N_5557,N_7221);
and U10974 (N_10974,N_7327,N_5406);
or U10975 (N_10975,N_6050,N_6956);
or U10976 (N_10976,N_6363,N_9838);
xnor U10977 (N_10977,N_9152,N_6390);
nand U10978 (N_10978,N_9441,N_6414);
nor U10979 (N_10979,N_9886,N_6188);
and U10980 (N_10980,N_9451,N_5262);
or U10981 (N_10981,N_5905,N_9680);
nor U10982 (N_10982,N_8120,N_6578);
xnor U10983 (N_10983,N_6500,N_6663);
nor U10984 (N_10984,N_6555,N_5735);
and U10985 (N_10985,N_8520,N_6259);
nor U10986 (N_10986,N_5873,N_6612);
and U10987 (N_10987,N_6770,N_7040);
or U10988 (N_10988,N_7932,N_5110);
and U10989 (N_10989,N_5040,N_7965);
nand U10990 (N_10990,N_7057,N_6158);
nand U10991 (N_10991,N_7480,N_6670);
nor U10992 (N_10992,N_9009,N_6089);
nor U10993 (N_10993,N_7194,N_7526);
nor U10994 (N_10994,N_8287,N_5697);
xnor U10995 (N_10995,N_8655,N_6896);
xor U10996 (N_10996,N_9162,N_8309);
nand U10997 (N_10997,N_6722,N_7779);
or U10998 (N_10998,N_7175,N_9277);
and U10999 (N_10999,N_5638,N_6885);
nor U11000 (N_11000,N_7390,N_9210);
xor U11001 (N_11001,N_5587,N_8562);
xor U11002 (N_11002,N_8133,N_6477);
or U11003 (N_11003,N_9494,N_7812);
nand U11004 (N_11004,N_6921,N_5932);
nand U11005 (N_11005,N_8863,N_7854);
or U11006 (N_11006,N_8212,N_9358);
or U11007 (N_11007,N_6830,N_6575);
nand U11008 (N_11008,N_7769,N_8780);
nor U11009 (N_11009,N_5442,N_7199);
xor U11010 (N_11010,N_6320,N_9056);
nor U11011 (N_11011,N_5377,N_5980);
xor U11012 (N_11012,N_6351,N_8341);
or U11013 (N_11013,N_9315,N_7034);
and U11014 (N_11014,N_8664,N_5012);
and U11015 (N_11015,N_5364,N_6439);
nand U11016 (N_11016,N_5539,N_6835);
or U11017 (N_11017,N_6245,N_8021);
and U11018 (N_11018,N_5185,N_6458);
and U11019 (N_11019,N_6524,N_8634);
nor U11020 (N_11020,N_6286,N_5058);
nand U11021 (N_11021,N_8769,N_5593);
xnor U11022 (N_11022,N_9739,N_8970);
or U11023 (N_11023,N_5386,N_8300);
or U11024 (N_11024,N_6729,N_5169);
and U11025 (N_11025,N_8620,N_7213);
nand U11026 (N_11026,N_9324,N_9665);
nor U11027 (N_11027,N_7504,N_8347);
xor U11028 (N_11028,N_9115,N_7966);
xor U11029 (N_11029,N_8328,N_7559);
nand U11030 (N_11030,N_8007,N_5968);
and U11031 (N_11031,N_6753,N_9778);
or U11032 (N_11032,N_8828,N_5052);
nor U11033 (N_11033,N_6125,N_6817);
and U11034 (N_11034,N_6736,N_8374);
nand U11035 (N_11035,N_5120,N_5509);
xnor U11036 (N_11036,N_8644,N_8092);
xor U11037 (N_11037,N_6486,N_9923);
nand U11038 (N_11038,N_8775,N_7610);
nand U11039 (N_11039,N_7660,N_7496);
nand U11040 (N_11040,N_7771,N_9694);
nor U11041 (N_11041,N_5474,N_7994);
nand U11042 (N_11042,N_5236,N_5115);
nor U11043 (N_11043,N_5540,N_5940);
xnor U11044 (N_11044,N_7853,N_5416);
nor U11045 (N_11045,N_7073,N_5900);
and U11046 (N_11046,N_8643,N_8033);
xnor U11047 (N_11047,N_6432,N_6600);
nor U11048 (N_11048,N_6700,N_8611);
and U11049 (N_11049,N_6250,N_5172);
nand U11050 (N_11050,N_7015,N_6928);
nor U11051 (N_11051,N_5384,N_9537);
xnor U11052 (N_11052,N_7415,N_8471);
and U11053 (N_11053,N_6305,N_5229);
nand U11054 (N_11054,N_6548,N_6567);
xnor U11055 (N_11055,N_5888,N_6558);
nand U11056 (N_11056,N_8731,N_9097);
xnor U11057 (N_11057,N_8143,N_6636);
nand U11058 (N_11058,N_6629,N_5554);
and U11059 (N_11059,N_7776,N_9114);
nor U11060 (N_11060,N_6019,N_7419);
nor U11061 (N_11061,N_8308,N_9624);
nand U11062 (N_11062,N_8241,N_6871);
or U11063 (N_11063,N_7307,N_7243);
nor U11064 (N_11064,N_6031,N_9189);
or U11065 (N_11065,N_5153,N_8173);
nor U11066 (N_11066,N_8231,N_7835);
nand U11067 (N_11067,N_5640,N_7412);
nor U11068 (N_11068,N_9059,N_8346);
nand U11069 (N_11069,N_5772,N_9738);
or U11070 (N_11070,N_8188,N_5700);
or U11071 (N_11071,N_8421,N_5476);
nor U11072 (N_11072,N_6929,N_6177);
nand U11073 (N_11073,N_5881,N_7118);
nand U11074 (N_11074,N_7418,N_5898);
xor U11075 (N_11075,N_7887,N_7163);
and U11076 (N_11076,N_7967,N_6150);
or U11077 (N_11077,N_7677,N_9563);
and U11078 (N_11078,N_6491,N_8481);
nand U11079 (N_11079,N_6679,N_6446);
or U11080 (N_11080,N_6443,N_6660);
and U11081 (N_11081,N_7191,N_5929);
and U11082 (N_11082,N_5319,N_9459);
nand U11083 (N_11083,N_6293,N_9286);
or U11084 (N_11084,N_7652,N_9683);
and U11085 (N_11085,N_8666,N_5761);
xnor U11086 (N_11086,N_8438,N_9942);
nor U11087 (N_11087,N_7784,N_7664);
xnor U11088 (N_11088,N_9062,N_8905);
nor U11089 (N_11089,N_5692,N_9467);
or U11090 (N_11090,N_7670,N_9781);
nand U11091 (N_11091,N_5890,N_5514);
or U11092 (N_11092,N_5492,N_5449);
or U11093 (N_11093,N_9930,N_6955);
and U11094 (N_11094,N_7951,N_9320);
nand U11095 (N_11095,N_8384,N_6715);
xor U11096 (N_11096,N_6136,N_8468);
nand U11097 (N_11097,N_7272,N_6329);
or U11098 (N_11098,N_5766,N_5908);
or U11099 (N_11099,N_8995,N_6985);
or U11100 (N_11100,N_9403,N_5754);
and U11101 (N_11101,N_6549,N_6113);
or U11102 (N_11102,N_7310,N_9621);
nand U11103 (N_11103,N_8463,N_9435);
nor U11104 (N_11104,N_7638,N_5030);
nand U11105 (N_11105,N_8915,N_9880);
or U11106 (N_11106,N_6032,N_7538);
nand U11107 (N_11107,N_6994,N_9424);
xnor U11108 (N_11108,N_7325,N_8852);
xnor U11109 (N_11109,N_9885,N_6648);
and U11110 (N_11110,N_9540,N_8166);
or U11111 (N_11111,N_5140,N_6998);
nand U11112 (N_11112,N_7796,N_7362);
xnor U11113 (N_11113,N_9958,N_5425);
and U11114 (N_11114,N_5061,N_6407);
nor U11115 (N_11115,N_7493,N_5594);
nor U11116 (N_11116,N_9938,N_6757);
nand U11117 (N_11117,N_8555,N_5114);
nand U11118 (N_11118,N_7317,N_8097);
or U11119 (N_11119,N_8270,N_6291);
nand U11120 (N_11120,N_5704,N_6856);
xor U11121 (N_11121,N_7794,N_6635);
nor U11122 (N_11122,N_7564,N_5325);
nor U11123 (N_11123,N_9510,N_6261);
xnor U11124 (N_11124,N_9945,N_9760);
or U11125 (N_11125,N_7629,N_7996);
or U11126 (N_11126,N_5318,N_8856);
nor U11127 (N_11127,N_5108,N_6507);
and U11128 (N_11128,N_5448,N_6244);
nand U11129 (N_11129,N_6967,N_5122);
or U11130 (N_11130,N_9253,N_9101);
and U11131 (N_11131,N_8745,N_6628);
nor U11132 (N_11132,N_8419,N_7762);
nor U11133 (N_11133,N_7372,N_7420);
or U11134 (N_11134,N_6743,N_6483);
nor U11135 (N_11135,N_6004,N_6556);
xnor U11136 (N_11136,N_7850,N_9655);
xnor U11137 (N_11137,N_8277,N_8844);
or U11138 (N_11138,N_6020,N_5171);
nand U11139 (N_11139,N_5330,N_6781);
and U11140 (N_11140,N_5948,N_5938);
or U11141 (N_11141,N_5762,N_6239);
nand U11142 (N_11142,N_9759,N_9749);
nand U11143 (N_11143,N_5413,N_8692);
and U11144 (N_11144,N_5372,N_6603);
nor U11145 (N_11145,N_9450,N_7639);
or U11146 (N_11146,N_9973,N_8191);
xnor U11147 (N_11147,N_8937,N_8516);
nor U11148 (N_11148,N_9791,N_5380);
xor U11149 (N_11149,N_8113,N_9113);
nand U11150 (N_11150,N_6713,N_6137);
xnor U11151 (N_11151,N_7131,N_6854);
nor U11152 (N_11152,N_6240,N_8543);
and U11153 (N_11153,N_9195,N_8487);
nor U11154 (N_11154,N_7109,N_7527);
and U11155 (N_11155,N_6201,N_8026);
and U11156 (N_11156,N_8797,N_5868);
and U11157 (N_11157,N_6475,N_5002);
xor U11158 (N_11158,N_7294,N_5329);
nand U11159 (N_11159,N_5050,N_7710);
nand U11160 (N_11160,N_8138,N_7180);
nand U11161 (N_11161,N_6118,N_9388);
and U11162 (N_11162,N_9921,N_7993);
xnor U11163 (N_11163,N_9741,N_9776);
or U11164 (N_11164,N_9032,N_6302);
and U11165 (N_11165,N_5174,N_7977);
and U11166 (N_11166,N_5382,N_6144);
and U11167 (N_11167,N_9232,N_9790);
or U11168 (N_11168,N_9637,N_6838);
xnor U11169 (N_11169,N_7378,N_8530);
and U11170 (N_11170,N_5630,N_5350);
nor U11171 (N_11171,N_5744,N_7299);
nand U11172 (N_11172,N_9411,N_9416);
or U11173 (N_11173,N_8515,N_7341);
or U11174 (N_11174,N_7125,N_5485);
xor U11175 (N_11175,N_7770,N_9444);
or U11176 (N_11176,N_9784,N_8390);
and U11177 (N_11177,N_6632,N_9465);
xnor U11178 (N_11178,N_5660,N_7623);
or U11179 (N_11179,N_5298,N_8233);
nor U11180 (N_11180,N_8336,N_7037);
nor U11181 (N_11181,N_6157,N_7657);
and U11182 (N_11182,N_5269,N_7261);
or U11183 (N_11183,N_7530,N_8603);
and U11184 (N_11184,N_6845,N_5391);
xor U11185 (N_11185,N_7778,N_5548);
or U11186 (N_11186,N_7566,N_5752);
xor U11187 (N_11187,N_9492,N_9982);
nor U11188 (N_11188,N_7437,N_7485);
nor U11189 (N_11189,N_6276,N_9651);
and U11190 (N_11190,N_6361,N_9389);
nor U11191 (N_11191,N_9998,N_9536);
nor U11192 (N_11192,N_7335,N_9663);
nor U11193 (N_11193,N_6775,N_7298);
nand U11194 (N_11194,N_5088,N_7792);
xor U11195 (N_11195,N_6145,N_6810);
or U11196 (N_11196,N_5109,N_9785);
and U11197 (N_11197,N_9166,N_6053);
xnor U11198 (N_11198,N_7429,N_7643);
or U11199 (N_11199,N_6077,N_6803);
nor U11200 (N_11200,N_7695,N_8235);
and U11201 (N_11201,N_8681,N_9615);
nor U11202 (N_11202,N_7764,N_8881);
nor U11203 (N_11203,N_7582,N_7620);
and U11204 (N_11204,N_8820,N_7189);
nand U11205 (N_11205,N_7244,N_7172);
nand U11206 (N_11206,N_8340,N_5261);
and U11207 (N_11207,N_9250,N_9213);
nor U11208 (N_11208,N_5435,N_6008);
nor U11209 (N_11209,N_6237,N_6189);
or U11210 (N_11210,N_8781,N_7267);
nand U11211 (N_11211,N_7683,N_9866);
or U11212 (N_11212,N_7906,N_5500);
nand U11213 (N_11213,N_6607,N_7914);
nand U11214 (N_11214,N_9119,N_7478);
nand U11215 (N_11215,N_5865,N_8766);
xor U11216 (N_11216,N_6947,N_8141);
xnor U11217 (N_11217,N_7604,N_6049);
nor U11218 (N_11218,N_9870,N_8677);
and U11219 (N_11219,N_7059,N_8206);
and U11220 (N_11220,N_9558,N_7264);
nand U11221 (N_11221,N_5202,N_9996);
or U11222 (N_11222,N_6069,N_7248);
or U11223 (N_11223,N_9072,N_7984);
nor U11224 (N_11224,N_9887,N_8717);
nor U11225 (N_11225,N_8290,N_5658);
nor U11226 (N_11226,N_7821,N_8326);
or U11227 (N_11227,N_7113,N_9547);
or U11228 (N_11228,N_6529,N_7474);
and U11229 (N_11229,N_8274,N_8410);
nand U11230 (N_11230,N_8255,N_5438);
or U11231 (N_11231,N_8799,N_6598);
xor U11232 (N_11232,N_5844,N_6203);
xor U11233 (N_11233,N_6815,N_7104);
xnor U11234 (N_11234,N_5387,N_8495);
or U11235 (N_11235,N_9726,N_8740);
nand U11236 (N_11236,N_6720,N_9289);
xnor U11237 (N_11237,N_8949,N_5959);
xnor U11238 (N_11238,N_5803,N_9578);
and U11239 (N_11239,N_7905,N_7407);
nor U11240 (N_11240,N_9606,N_7912);
or U11241 (N_11241,N_6786,N_5583);
xnor U11242 (N_11242,N_8377,N_8559);
nand U11243 (N_11243,N_6406,N_5742);
and U11244 (N_11244,N_8917,N_5790);
or U11245 (N_11245,N_8399,N_7384);
xor U11246 (N_11246,N_6024,N_8675);
nor U11247 (N_11247,N_7804,N_5842);
and U11248 (N_11248,N_5154,N_5130);
and U11249 (N_11249,N_9934,N_8891);
or U11250 (N_11250,N_5961,N_5276);
nand U11251 (N_11251,N_5233,N_9042);
xor U11252 (N_11252,N_8696,N_5405);
xnor U11253 (N_11253,N_7065,N_8522);
nor U11254 (N_11254,N_5156,N_9480);
xnor U11255 (N_11255,N_9820,N_8462);
xnor U11256 (N_11256,N_8579,N_8990);
and U11257 (N_11257,N_9613,N_9783);
and U11258 (N_11258,N_9040,N_7916);
or U11259 (N_11259,N_7798,N_7402);
nand U11260 (N_11260,N_9336,N_8505);
xnor U11261 (N_11261,N_7382,N_7233);
and U11262 (N_11262,N_7229,N_5839);
xor U11263 (N_11263,N_6826,N_5322);
or U11264 (N_11264,N_7701,N_6562);
nand U11265 (N_11265,N_8722,N_5791);
or U11266 (N_11266,N_7592,N_6449);
nand U11267 (N_11267,N_8090,N_9140);
or U11268 (N_11268,N_6481,N_6593);
nor U11269 (N_11269,N_9314,N_8663);
xor U11270 (N_11270,N_9919,N_6325);
nand U11271 (N_11271,N_6894,N_8875);
or U11272 (N_11272,N_5861,N_5304);
nor U11273 (N_11273,N_9955,N_7852);
nor U11274 (N_11274,N_7435,N_5393);
xor U11275 (N_11275,N_6022,N_6073);
and U11276 (N_11276,N_6114,N_8829);
nor U11277 (N_11277,N_8855,N_9127);
or U11278 (N_11278,N_9604,N_5429);
or U11279 (N_11279,N_8728,N_5643);
and U11280 (N_11280,N_8087,N_8174);
nand U11281 (N_11281,N_9900,N_7814);
or U11282 (N_11282,N_7115,N_5099);
or U11283 (N_11283,N_8402,N_6752);
nor U11284 (N_11284,N_6680,N_8956);
nand U11285 (N_11285,N_9184,N_7292);
or U11286 (N_11286,N_9204,N_9061);
nor U11287 (N_11287,N_5417,N_5272);
nor U11288 (N_11288,N_8809,N_9641);
xnor U11289 (N_11289,N_5871,N_6001);
nor U11290 (N_11290,N_8367,N_9299);
nand U11291 (N_11291,N_6368,N_7070);
or U11292 (N_11292,N_6447,N_5066);
or U11293 (N_11293,N_6839,N_6249);
and U11294 (N_11294,N_6209,N_6525);
nor U11295 (N_11295,N_5718,N_7052);
xnor U11296 (N_11296,N_6814,N_5031);
xnor U11297 (N_11297,N_5703,N_5434);
nand U11298 (N_11298,N_9084,N_5618);
nor U11299 (N_11299,N_8550,N_8816);
nor U11300 (N_11300,N_8139,N_6379);
nand U11301 (N_11301,N_5128,N_7083);
nand U11302 (N_11302,N_9839,N_8178);
nor U11303 (N_11303,N_6879,N_5053);
and U11304 (N_11304,N_9569,N_7991);
xor U11305 (N_11305,N_9400,N_8157);
xnor U11306 (N_11306,N_5097,N_6834);
xnor U11307 (N_11307,N_9329,N_7619);
or U11308 (N_11308,N_9638,N_9672);
xnor U11309 (N_11309,N_7858,N_7347);
nor U11310 (N_11310,N_7506,N_7572);
xnor U11311 (N_11311,N_9664,N_7531);
and U11312 (N_11312,N_9597,N_9577);
nor U11313 (N_11313,N_7686,N_6460);
and U11314 (N_11314,N_7356,N_7124);
nor U11315 (N_11315,N_7716,N_8386);
nor U11316 (N_11316,N_9795,N_7376);
or U11317 (N_11317,N_9935,N_7697);
nor U11318 (N_11318,N_8128,N_5055);
nand U11319 (N_11319,N_8289,N_6057);
xor U11320 (N_11320,N_5226,N_5616);
xnor U11321 (N_11321,N_6709,N_5577);
and U11322 (N_11322,N_9636,N_8783);
nand U11323 (N_11323,N_9045,N_5401);
nand U11324 (N_11324,N_9267,N_8169);
nand U11325 (N_11325,N_9626,N_7751);
and U11326 (N_11326,N_9990,N_5168);
and U11327 (N_11327,N_5650,N_6257);
nor U11328 (N_11328,N_7758,N_6579);
or U11329 (N_11329,N_5344,N_6234);
and U11330 (N_11330,N_9290,N_6074);
or U11331 (N_11331,N_6528,N_8119);
and U11332 (N_11332,N_7024,N_6169);
or U11333 (N_11333,N_9236,N_8889);
nand U11334 (N_11334,N_9495,N_6809);
nor U11335 (N_11335,N_5526,N_8022);
or U11336 (N_11336,N_8808,N_9060);
or U11337 (N_11337,N_7208,N_6147);
or U11338 (N_11338,N_7112,N_5044);
nand U11339 (N_11339,N_9803,N_9888);
nor U11340 (N_11340,N_7757,N_6480);
nand U11341 (N_11341,N_9326,N_5887);
nor U11342 (N_11342,N_8616,N_8163);
nor U11343 (N_11343,N_8591,N_9640);
and U11344 (N_11344,N_8968,N_9905);
nor U11345 (N_11345,N_7508,N_8541);
nor U11346 (N_11346,N_5019,N_5717);
and U11347 (N_11347,N_8023,N_9193);
nor U11348 (N_11348,N_5295,N_8094);
xnor U11349 (N_11349,N_5113,N_5840);
nor U11350 (N_11350,N_7505,N_9724);
and U11351 (N_11351,N_5686,N_5920);
nor U11352 (N_11352,N_5098,N_9186);
nor U11353 (N_11353,N_9296,N_6708);
and U11354 (N_11354,N_8252,N_8892);
or U11355 (N_11355,N_8971,N_8556);
xor U11356 (N_11356,N_8689,N_8623);
xnor U11357 (N_11357,N_7535,N_8387);
xnor U11358 (N_11358,N_8187,N_8086);
xnor U11359 (N_11359,N_5728,N_7337);
xor U11360 (N_11360,N_5283,N_8323);
nor U11361 (N_11361,N_9309,N_8713);
nor U11362 (N_11362,N_9848,N_9091);
nor U11363 (N_11363,N_8942,N_6367);
xnor U11364 (N_11364,N_7929,N_8071);
and U11365 (N_11365,N_9835,N_9669);
and U11366 (N_11366,N_6504,N_5504);
and U11367 (N_11367,N_7479,N_5285);
nor U11368 (N_11368,N_8031,N_9278);
xnor U11369 (N_11369,N_7203,N_9490);
xor U11370 (N_11370,N_9363,N_7232);
or U11371 (N_11371,N_5667,N_6143);
or U11372 (N_11372,N_6609,N_6801);
and U11373 (N_11373,N_8838,N_6142);
nor U11374 (N_11374,N_5375,N_9901);
nand U11375 (N_11375,N_7803,N_9183);
xnor U11376 (N_11376,N_5684,N_5586);
xnor U11377 (N_11377,N_9361,N_7785);
nor U11378 (N_11378,N_5688,N_5212);
or U11379 (N_11379,N_7458,N_7884);
or U11380 (N_11380,N_5256,N_8793);
and U11381 (N_11381,N_5451,N_8792);
nand U11382 (N_11382,N_9229,N_6090);
nand U11383 (N_11383,N_8538,N_6571);
and U11384 (N_11384,N_7972,N_7020);
nand U11385 (N_11385,N_8501,N_8125);
nand U11386 (N_11386,N_7274,N_5173);
nand U11387 (N_11387,N_9370,N_9612);
or U11388 (N_11388,N_9212,N_7513);
nor U11389 (N_11389,N_7091,N_7366);
xnor U11390 (N_11390,N_8314,N_9860);
and U11391 (N_11391,N_8077,N_5730);
and U11392 (N_11392,N_6867,N_6978);
nor U11393 (N_11393,N_6319,N_7278);
and U11394 (N_11394,N_5265,N_5963);
xor U11395 (N_11395,N_9731,N_9410);
nor U11396 (N_11396,N_6154,N_7601);
and U11397 (N_11397,N_7866,N_9327);
nor U11398 (N_11398,N_8279,N_8833);
xnor U11399 (N_11399,N_7302,N_7810);
xnor U11400 (N_11400,N_9639,N_6800);
xnor U11401 (N_11401,N_9109,N_8951);
xor U11402 (N_11402,N_7334,N_9058);
or U11403 (N_11403,N_6676,N_6247);
xor U11404 (N_11404,N_6922,N_5793);
and U11405 (N_11405,N_7727,N_5503);
or U11406 (N_11406,N_9125,N_5374);
and U11407 (N_11407,N_6857,N_9774);
nand U11408 (N_11408,N_6825,N_5246);
and U11409 (N_11409,N_8899,N_6101);
nand U11410 (N_11410,N_9978,N_8776);
xnor U11411 (N_11411,N_8588,N_6352);
nand U11412 (N_11412,N_9610,N_9972);
nor U11413 (N_11413,N_9319,N_7231);
and U11414 (N_11414,N_7501,N_7168);
and U11415 (N_11415,N_7004,N_6927);
or U11416 (N_11416,N_6212,N_7726);
nor U11417 (N_11417,N_6108,N_9780);
nor U11418 (N_11418,N_5084,N_8321);
xor U11419 (N_11419,N_8884,N_6706);
and U11420 (N_11420,N_5877,N_6155);
or U11421 (N_11421,N_7625,N_9912);
and U11422 (N_11422,N_9334,N_7013);
xor U11423 (N_11423,N_9721,N_5186);
nor U11424 (N_11424,N_9910,N_5146);
and U11425 (N_11425,N_8369,N_8302);
and U11426 (N_11426,N_5901,N_9811);
and U11427 (N_11427,N_7388,N_7768);
xor U11428 (N_11428,N_8060,N_6595);
xnor U11429 (N_11429,N_5412,N_5039);
and U11430 (N_11430,N_6227,N_5370);
or U11431 (N_11431,N_9959,N_9516);
nor U11432 (N_11432,N_6509,N_6464);
or U11433 (N_11433,N_8880,N_6889);
nand U11434 (N_11434,N_7187,N_9971);
or U11435 (N_11435,N_6369,N_9242);
and U11436 (N_11436,N_8316,N_7174);
or U11437 (N_11437,N_8025,N_9822);
or U11438 (N_11438,N_6340,N_9675);
and U11439 (N_11439,N_5994,N_7002);
or U11440 (N_11440,N_8203,N_5060);
and U11441 (N_11441,N_5407,N_7225);
and U11442 (N_11442,N_5649,N_7216);
and U11443 (N_11443,N_5022,N_6566);
or U11444 (N_11444,N_6589,N_7408);
xnor U11445 (N_11445,N_7839,N_5921);
nand U11446 (N_11446,N_5741,N_7765);
xnor U11447 (N_11447,N_9814,N_7684);
xor U11448 (N_11448,N_5928,N_6198);
or U11449 (N_11449,N_7094,N_9893);
xor U11450 (N_11450,N_6264,N_8132);
and U11451 (N_11451,N_8005,N_6932);
nand U11452 (N_11452,N_6872,N_5165);
xor U11453 (N_11453,N_7220,N_9499);
and U11454 (N_11454,N_7179,N_6455);
nand U11455 (N_11455,N_5253,N_8787);
nand U11456 (N_11456,N_7746,N_6116);
nand U11457 (N_11457,N_6405,N_7963);
nor U11458 (N_11458,N_6284,N_6793);
nand U11459 (N_11459,N_7886,N_6034);
or U11460 (N_11460,N_7392,N_6466);
xnor U11461 (N_11461,N_6550,N_8454);
xor U11462 (N_11462,N_7855,N_9464);
xor U11463 (N_11463,N_6682,N_6398);
nor U11464 (N_11464,N_6923,N_9054);
and U11465 (N_11465,N_9914,N_8343);
nand U11466 (N_11466,N_6843,N_8823);
nand U11467 (N_11467,N_7735,N_9328);
and U11468 (N_11468,N_6758,N_6832);
and U11469 (N_11469,N_8472,N_8320);
or U11470 (N_11470,N_9067,N_5479);
and U11471 (N_11471,N_7129,N_8149);
nand U11472 (N_11472,N_9052,N_8686);
nor U11473 (N_11473,N_6346,N_8757);
or U11474 (N_11474,N_7322,N_8593);
nand U11475 (N_11475,N_5596,N_8268);
xor U11476 (N_11476,N_7846,N_5404);
and U11477 (N_11477,N_7723,N_8802);
xor U11478 (N_11478,N_5965,N_8795);
or U11479 (N_11479,N_9770,N_6469);
or U11480 (N_11480,N_5523,N_8846);
and U11481 (N_11481,N_7308,N_5303);
xor U11482 (N_11482,N_5875,N_7926);
and U11483 (N_11483,N_9105,N_6962);
nor U11484 (N_11484,N_8453,N_8224);
and U11485 (N_11485,N_5670,N_7802);
nand U11486 (N_11486,N_5297,N_9503);
xor U11487 (N_11487,N_9508,N_7608);
or U11488 (N_11488,N_6206,N_6505);
and U11489 (N_11489,N_7799,N_8552);
nor U11490 (N_11490,N_8922,N_5612);
and U11491 (N_11491,N_6176,N_7247);
xnor U11492 (N_11492,N_9756,N_8000);
or U11493 (N_11493,N_8437,N_8727);
nor U11494 (N_11494,N_7833,N_5148);
and U11495 (N_11495,N_6531,N_5273);
xnor U11496 (N_11496,N_9544,N_6621);
and U11497 (N_11497,N_9458,N_5136);
nand U11498 (N_11498,N_7060,N_6828);
nand U11499 (N_11499,N_9237,N_6300);
nor U11500 (N_11500,N_9594,N_5347);
xnor U11501 (N_11501,N_5879,N_5782);
and U11502 (N_11502,N_9412,N_5906);
xnor U11503 (N_11503,N_5469,N_7349);
and U11504 (N_11504,N_5683,N_8506);
xnor U11505 (N_11505,N_6798,N_9360);
and U11506 (N_11506,N_7908,N_8804);
and U11507 (N_11507,N_9279,N_5191);
nor U11508 (N_11508,N_7789,N_9348);
xnor U11509 (N_11509,N_5324,N_9535);
and U11510 (N_11510,N_9445,N_7461);
or U11511 (N_11511,N_6653,N_5308);
nor U11512 (N_11512,N_5998,N_5065);
nand U11513 (N_11513,N_6818,N_5975);
and U11514 (N_11514,N_5455,N_6487);
nand U11515 (N_11515,N_6668,N_5724);
xnor U11516 (N_11516,N_6401,N_9461);
or U11517 (N_11517,N_5251,N_7029);
and U11518 (N_11518,N_6453,N_7078);
and U11519 (N_11519,N_8807,N_5691);
xor U11520 (N_11520,N_5740,N_6230);
xor U11521 (N_11521,N_8041,N_5738);
xnor U11522 (N_11522,N_9112,N_5690);
and U11523 (N_11523,N_8989,N_6841);
nand U11524 (N_11524,N_8887,N_9730);
and U11525 (N_11525,N_5885,N_5008);
or U11526 (N_11526,N_7999,N_5549);
nor U11527 (N_11527,N_6294,N_7128);
and U11528 (N_11528,N_8817,N_5800);
and U11529 (N_11529,N_5205,N_5354);
or U11530 (N_11530,N_9878,N_7571);
xor U11531 (N_11531,N_5221,N_6336);
nand U11532 (N_11532,N_9300,N_9674);
and U11533 (N_11533,N_5833,N_9332);
or U11534 (N_11534,N_9220,N_9479);
nor U11535 (N_11535,N_6954,N_5057);
nand U11536 (N_11536,N_5926,N_9160);
nand U11537 (N_11537,N_5021,N_5751);
nor U11538 (N_11538,N_9884,N_5544);
nand U11539 (N_11539,N_6777,N_5789);
or U11540 (N_11540,N_9762,N_6012);
and U11541 (N_11541,N_9779,N_6199);
nor U11542 (N_11542,N_7486,N_5049);
or U11543 (N_11543,N_9896,N_6584);
nor U11544 (N_11544,N_6623,N_9717);
or U11545 (N_11545,N_7003,N_6694);
nor U11546 (N_11546,N_7176,N_7295);
or U11547 (N_11547,N_5142,N_6605);
or U11548 (N_11548,N_6205,N_6960);
xnor U11549 (N_11549,N_7577,N_6148);
xnor U11550 (N_11550,N_9068,N_7483);
or U11551 (N_11551,N_7544,N_5778);
xor U11552 (N_11552,N_9208,N_9298);
or U11553 (N_11553,N_7645,N_6912);
and U11554 (N_11554,N_7615,N_5124);
or U11555 (N_11555,N_9128,N_8752);
nand U11556 (N_11556,N_6836,N_5952);
or U11557 (N_11557,N_7111,N_6699);
xor U11558 (N_11558,N_6330,N_6195);
or U11559 (N_11559,N_9666,N_7773);
xnor U11560 (N_11560,N_6041,N_6218);
and U11561 (N_11561,N_8406,N_6767);
nor U11562 (N_11562,N_7551,N_7198);
nor U11563 (N_11563,N_7763,N_5456);
nor U11564 (N_11564,N_5190,N_7874);
and U11565 (N_11565,N_9605,N_9151);
and U11566 (N_11566,N_5547,N_9284);
and U11567 (N_11567,N_9956,N_9931);
or U11568 (N_11568,N_5101,N_6915);
or U11569 (N_11569,N_9273,N_8359);
xnor U11570 (N_11570,N_6412,N_5810);
xor U11571 (N_11571,N_5428,N_6015);
nor U11572 (N_11572,N_7894,N_5707);
or U11573 (N_11573,N_5309,N_9812);
nand U11574 (N_11574,N_5846,N_6888);
nand U11575 (N_11575,N_8214,N_8733);
nand U11576 (N_11576,N_7633,N_9260);
and U11577 (N_11577,N_6705,N_8512);
xnor U11578 (N_11578,N_8258,N_6213);
or U11579 (N_11579,N_5197,N_7614);
xor U11580 (N_11580,N_8229,N_5332);
nor U11581 (N_11581,N_7931,N_5797);
nand U11582 (N_11582,N_5934,N_9534);
nand U11583 (N_11583,N_8739,N_6345);
nor U11584 (N_11584,N_8975,N_9714);
xnor U11585 (N_11585,N_9231,N_6697);
nor U11586 (N_11586,N_8389,N_5689);
xor U11587 (N_11587,N_8779,N_8052);
or U11588 (N_11588,N_5786,N_6712);
nor U11589 (N_11589,N_9238,N_5923);
and U11590 (N_11590,N_6344,N_8247);
nor U11591 (N_11591,N_5537,N_7210);
or U11592 (N_11592,N_9312,N_9659);
nand U11593 (N_11593,N_7022,N_9747);
and U11594 (N_11594,N_7913,N_7467);
nor U11595 (N_11595,N_9384,N_6219);
nand U11596 (N_11596,N_7675,N_6622);
or U11597 (N_11597,N_6470,N_8527);
and U11598 (N_11598,N_8204,N_6170);
nor U11599 (N_11599,N_9678,N_9211);
or U11600 (N_11600,N_5832,N_6738);
and U11601 (N_11601,N_8411,N_8803);
xor U11602 (N_11602,N_7276,N_5328);
and U11603 (N_11603,N_7692,N_5990);
nand U11604 (N_11604,N_7158,N_6618);
or U11605 (N_11605,N_5395,N_7512);
or U11606 (N_11606,N_8069,N_7127);
or U11607 (N_11607,N_7937,N_5864);
xnor U11608 (N_11608,N_5041,N_8082);
or U11609 (N_11609,N_8650,N_8035);
or U11610 (N_11610,N_6582,N_9202);
xnor U11611 (N_11611,N_6479,N_5712);
nor U11612 (N_11612,N_8849,N_9123);
xor U11613 (N_11613,N_9408,N_6373);
or U11614 (N_11614,N_9104,N_9962);
and U11615 (N_11615,N_8749,N_6299);
or U11616 (N_11616,N_6349,N_8876);
and U11617 (N_11617,N_7671,N_5716);
xor U11618 (N_11618,N_6419,N_7082);
xor U11619 (N_11619,N_8784,N_9881);
nand U11620 (N_11620,N_7253,N_6914);
or U11621 (N_11621,N_6097,N_7968);
and U11622 (N_11622,N_8351,N_5432);
nor U11623 (N_11623,N_9704,N_8850);
xor U11624 (N_11624,N_5307,N_5411);
and U11625 (N_11625,N_9806,N_9796);
xnor U11626 (N_11626,N_6318,N_8080);
and U11627 (N_11627,N_7058,N_8484);
and U11628 (N_11628,N_8372,N_5430);
nor U11629 (N_11629,N_5166,N_6710);
or U11630 (N_11630,N_7679,N_7464);
xor U11631 (N_11631,N_9215,N_5288);
xnor U11632 (N_11632,N_5771,N_7238);
nand U11633 (N_11633,N_5613,N_9170);
nand U11634 (N_11634,N_5841,N_5360);
nor U11635 (N_11635,N_8504,N_7907);
xor U11636 (N_11636,N_5681,N_6769);
nand U11637 (N_11637,N_5001,N_9858);
or U11638 (N_11638,N_8503,N_6944);
nand U11639 (N_11639,N_9262,N_7491);
and U11640 (N_11640,N_5821,N_7036);
and U11641 (N_11641,N_6754,N_7476);
and U11642 (N_11642,N_5038,N_9815);
nor U11643 (N_11643,N_7736,N_8599);
or U11644 (N_11644,N_6908,N_9758);
nor U11645 (N_11645,N_9826,N_6554);
and U11646 (N_11646,N_6183,N_8409);
nor U11647 (N_11647,N_8575,N_5505);
xor U11648 (N_11648,N_9270,N_9482);
xnor U11649 (N_11649,N_5167,N_8618);
and U11650 (N_11650,N_6850,N_7788);
nor U11651 (N_11651,N_7834,N_6847);
nand U11652 (N_11652,N_7364,N_6779);
or U11653 (N_11653,N_8211,N_6476);
or U11654 (N_11654,N_7970,N_7204);
nand U11655 (N_11655,N_9752,N_9080);
nand U11656 (N_11656,N_7669,N_7576);
xnor U11657 (N_11657,N_9274,N_9963);
nor U11658 (N_11658,N_5392,N_5239);
xnor U11659 (N_11659,N_7898,N_8385);
nor U11660 (N_11660,N_5145,N_6005);
nand U11661 (N_11661,N_6248,N_5575);
nor U11662 (N_11662,N_8311,N_9777);
or U11663 (N_11663,N_5850,N_5935);
and U11664 (N_11664,N_6389,N_6898);
xor U11665 (N_11665,N_9670,N_5792);
or U11666 (N_11666,N_7935,N_6067);
xnor U11667 (N_11667,N_7288,N_9619);
and U11668 (N_11668,N_7827,N_6374);
or U11669 (N_11669,N_9419,N_7146);
or U11670 (N_11670,N_8934,N_8430);
xnor U11671 (N_11671,N_7424,N_7509);
and U11672 (N_11672,N_7870,N_8933);
or U11673 (N_11673,N_5977,N_7077);
xnor U11674 (N_11674,N_7801,N_6883);
nor U11675 (N_11675,N_8638,N_6774);
nand U11676 (N_11676,N_6971,N_7868);
nor U11677 (N_11677,N_6949,N_5074);
xor U11678 (N_11678,N_8440,N_5231);
nand U11679 (N_11679,N_7548,N_8029);
nand U11680 (N_11680,N_6976,N_8189);
or U11681 (N_11681,N_7787,N_8519);
or U11682 (N_11682,N_9364,N_5043);
nor U11683 (N_11683,N_9853,N_5922);
and U11684 (N_11684,N_6082,N_5845);
nor U11685 (N_11685,N_5989,N_7006);
xor U11686 (N_11686,N_7211,N_9111);
or U11687 (N_11687,N_8208,N_9843);
or U11688 (N_11688,N_5464,N_7747);
xnor U11689 (N_11689,N_8608,N_9497);
or U11690 (N_11690,N_7139,N_5962);
nand U11691 (N_11691,N_7909,N_7958);
xor U11692 (N_11692,N_7007,N_5250);
xor U11693 (N_11693,N_9517,N_7892);
nor U11694 (N_11694,N_6970,N_8431);
nor U11695 (N_11695,N_8647,N_9849);
xor U11696 (N_11696,N_7739,N_6565);
and U11697 (N_11697,N_7345,N_7537);
or U11698 (N_11698,N_8830,N_5345);
nor U11699 (N_11699,N_7843,N_7358);
xor U11700 (N_11700,N_6357,N_9081);
nand U11701 (N_11701,N_5858,N_7492);
or U11702 (N_11702,N_6335,N_8227);
and U11703 (N_11703,N_7277,N_9255);
or U11704 (N_11704,N_6553,N_8237);
xor U11705 (N_11705,N_9456,N_8220);
nor U11706 (N_11706,N_5224,N_9244);
nor U11707 (N_11707,N_9701,N_9929);
or U11708 (N_11708,N_8907,N_7411);
and U11709 (N_11709,N_8736,N_8565);
nand U11710 (N_11710,N_8177,N_6416);
nor U11711 (N_11711,N_9425,N_5931);
and U11712 (N_11712,N_5849,N_9512);
nand U11713 (N_11713,N_5188,N_7477);
and U11714 (N_11714,N_7038,N_6229);
xor U11715 (N_11715,N_9366,N_6006);
nor U11716 (N_11716,N_8327,N_7533);
xor U11717 (N_11717,N_6964,N_5601);
or U11718 (N_11718,N_7939,N_7471);
and U11719 (N_11719,N_5103,N_6471);
xnor U11720 (N_11720,N_5836,N_7154);
nand U11721 (N_11721,N_7818,N_5534);
nor U11722 (N_11722,N_5945,N_8498);
xnor U11723 (N_11723,N_5134,N_6110);
nor U11724 (N_11724,N_5187,N_7090);
xnor U11725 (N_11725,N_8646,N_9673);
or U11726 (N_11726,N_7580,N_8491);
nor U11727 (N_11727,N_9196,N_9235);
nand U11728 (N_11728,N_6422,N_6438);
and U11729 (N_11729,N_5282,N_7546);
nand U11730 (N_11730,N_7555,N_5158);
xor U11731 (N_11731,N_7200,N_8671);
or U11732 (N_11732,N_7152,N_9355);
nor U11733 (N_11733,N_5759,N_6986);
xnor U11734 (N_11734,N_7658,N_6717);
nand U11735 (N_11735,N_8819,N_7826);
nor U11736 (N_11736,N_9258,N_9460);
or U11737 (N_11737,N_7459,N_6164);
nand U11738 (N_11738,N_9063,N_7524);
nor U11739 (N_11739,N_6827,N_8825);
nand U11740 (N_11740,N_9029,N_9549);
nand U11741 (N_11741,N_6534,N_8217);
and U11742 (N_11742,N_5599,N_5336);
nand U11743 (N_11743,N_5997,N_5431);
nor U11744 (N_11744,N_7593,N_6281);
nor U11745 (N_11745,N_5624,N_5860);
or U11746 (N_11746,N_7864,N_5665);
or U11747 (N_11747,N_9075,N_9941);
or U11748 (N_11748,N_5611,N_8063);
nand U11749 (N_11749,N_6749,N_8701);
nor U11750 (N_11750,N_9581,N_7344);
nand U11751 (N_11751,N_6172,N_9633);
or U11752 (N_11752,N_6066,N_8475);
or U11753 (N_11753,N_9439,N_8004);
nor U11754 (N_11754,N_8940,N_7532);
and U11755 (N_11755,N_9443,N_9138);
or U11756 (N_11756,N_8055,N_5204);
and U11757 (N_11757,N_5573,N_5674);
xnor U11758 (N_11758,N_9711,N_7469);
nor U11759 (N_11759,N_7398,N_9689);
or U11760 (N_11760,N_9434,N_5986);
xor U11761 (N_11761,N_5192,N_6232);
xor U11762 (N_11762,N_8767,N_8805);
nand U11763 (N_11763,N_7706,N_9891);
or U11764 (N_11764,N_8123,N_7523);
or U11765 (N_11765,N_6413,N_8927);
xnor U11766 (N_11766,N_9349,N_6518);
and U11767 (N_11767,N_5484,N_9725);
nor U11768 (N_11768,N_7044,N_9472);
nor U11769 (N_11769,N_6849,N_8839);
nand U11770 (N_11770,N_8245,N_9191);
xnor U11771 (N_11771,N_9041,N_5571);
nand U11772 (N_11772,N_8770,N_9103);
nor U11773 (N_11773,N_9607,N_8903);
nand U11774 (N_11774,N_7502,N_8962);
and U11775 (N_11775,N_6107,N_7955);
nand U11776 (N_11776,N_8657,N_5073);
xor U11777 (N_11777,N_8811,N_9662);
nand U11778 (N_11778,N_8624,N_6465);
nor U11779 (N_11779,N_5369,N_5763);
nor U11780 (N_11780,N_5402,N_7644);
xnor U11781 (N_11781,N_6959,N_9550);
nor U11782 (N_11782,N_5709,N_6904);
xor U11783 (N_11783,N_7861,N_5673);
nor U11784 (N_11784,N_6461,N_8485);
and U11785 (N_11785,N_6616,N_8114);
and U11786 (N_11786,N_9531,N_5756);
and U11787 (N_11787,N_6785,N_6310);
xnor U11788 (N_11788,N_8551,N_5659);
and U11789 (N_11789,N_6431,N_7901);
nand U11790 (N_11790,N_9050,N_7918);
or U11791 (N_11791,N_6819,N_7715);
xor U11792 (N_11792,N_5346,N_8436);
xnor U11793 (N_11793,N_9468,N_8688);
and U11794 (N_11794,N_9239,N_7860);
nor U11795 (N_11795,N_6863,N_8869);
nor U11796 (N_11796,N_6075,N_5477);
xnor U11797 (N_11797,N_5483,N_9735);
and U11798 (N_11798,N_9592,N_7678);
xnor U11799 (N_11799,N_5696,N_7974);
and U11800 (N_11800,N_9402,N_9989);
nor U11801 (N_11801,N_8796,N_6703);
and U11802 (N_11802,N_9044,N_8417);
nand U11803 (N_11803,N_7594,N_8678);
and U11804 (N_11804,N_9002,N_5446);
and U11805 (N_11805,N_5359,N_9165);
or U11806 (N_11806,N_6681,N_7289);
or U11807 (N_11807,N_5715,N_5851);
nand U11808 (N_11808,N_6765,N_5775);
or U11809 (N_11809,N_9505,N_8534);
xor U11810 (N_11810,N_8873,N_9474);
or U11811 (N_11811,N_7305,N_8794);
nand U11812 (N_11812,N_7328,N_6724);
nand U11813 (N_11813,N_7903,N_6644);
nand U11814 (N_11814,N_6161,N_7556);
and U11815 (N_11815,N_5623,N_9367);
nor U11816 (N_11816,N_6216,N_8054);
xnor U11817 (N_11817,N_8375,N_6999);
or U11818 (N_11818,N_5984,N_8553);
and U11819 (N_11819,N_5141,N_7565);
nand U11820 (N_11820,N_7688,N_5915);
and U11821 (N_11821,N_7522,N_7586);
xnor U11822 (N_11822,N_8042,N_7720);
xnor U11823 (N_11823,N_6730,N_5826);
or U11824 (N_11824,N_8832,N_5152);
or U11825 (N_11825,N_7401,N_8159);
or U11826 (N_11826,N_7444,N_8053);
xnor U11827 (N_11827,N_8012,N_8992);
xor U11828 (N_11828,N_5825,N_7662);
and U11829 (N_11829,N_7069,N_5719);
nand U11830 (N_11830,N_8117,N_5062);
and U11831 (N_11831,N_8199,N_8470);
or U11832 (N_11832,N_6920,N_8721);
xor U11833 (N_11833,N_8018,N_6221);
nand U11834 (N_11834,N_7095,N_9821);
and U11835 (N_11835,N_9859,N_9543);
and U11836 (N_11836,N_5468,N_6016);
or U11837 (N_11837,N_9004,N_8908);
nand U11838 (N_11838,N_5542,N_5129);
and U11839 (N_11839,N_7975,N_9984);
nor U11840 (N_11840,N_5025,N_7708);
nand U11841 (N_11841,N_9970,N_5525);
nand U11842 (N_11842,N_8275,N_8065);
and U11843 (N_11843,N_6996,N_9427);
or U11844 (N_11844,N_8356,N_5217);
xnor U11845 (N_11845,N_5138,N_6410);
and U11846 (N_11846,N_5189,N_5082);
and U11847 (N_11847,N_8046,N_8186);
xnor U11848 (N_11848,N_7885,N_9401);
nand U11849 (N_11849,N_9676,N_7817);
nor U11850 (N_11850,N_6763,N_5263);
xor U11851 (N_11851,N_5726,N_5506);
nor U11852 (N_11852,N_7350,N_6691);
xnor U11853 (N_11853,N_7865,N_5796);
xnor U11854 (N_11854,N_9362,N_8509);
nor U11855 (N_11855,N_5809,N_9035);
nand U11856 (N_11856,N_9997,N_6327);
nand U11857 (N_11857,N_6533,N_8645);
or U11858 (N_11858,N_9999,N_7647);
or U11859 (N_11859,N_9699,N_9546);
xor U11860 (N_11860,N_8723,N_9079);
and U11861 (N_11861,N_6297,N_7938);
nand U11862 (N_11862,N_5271,N_5941);
xor U11863 (N_11863,N_9264,N_5918);
or U11864 (N_11864,N_7982,N_7079);
xnor U11865 (N_11865,N_8720,N_9382);
xnor U11866 (N_11866,N_6561,N_6806);
and U11867 (N_11867,N_7268,N_9070);
nor U11868 (N_11868,N_5275,N_5996);
or U11869 (N_11869,N_6163,N_9233);
and U11870 (N_11870,N_6859,N_6468);
or U11871 (N_11871,N_9585,N_5046);
xnor U11872 (N_11872,N_5555,N_9734);
nor U11873 (N_11873,N_9222,N_9280);
xor U11874 (N_11874,N_7290,N_8413);
or U11875 (N_11875,N_7873,N_6522);
or U11876 (N_11876,N_7990,N_8558);
or U11877 (N_11877,N_6064,N_7132);
xnor U11878 (N_11878,N_6659,N_7063);
xor U11879 (N_11879,N_8223,N_8751);
nor U11880 (N_11880,N_8712,N_5927);
or U11881 (N_11881,N_7447,N_6764);
nor U11882 (N_11882,N_7092,N_5147);
nor U11883 (N_11883,N_5133,N_8478);
xor U11884 (N_11884,N_6910,N_6122);
xnor U11885 (N_11885,N_6687,N_9022);
and U11886 (N_11886,N_8524,N_6000);
xnor U11887 (N_11887,N_5530,N_7836);
or U11888 (N_11888,N_5106,N_6794);
or U11889 (N_11889,N_7561,N_9177);
nand U11890 (N_11890,N_8331,N_5936);
or U11891 (N_11891,N_9698,N_7385);
xnor U11892 (N_11892,N_7722,N_9308);
nor U11893 (N_11893,N_8439,N_8228);
nor U11894 (N_11894,N_9182,N_6217);
nor U11895 (N_11895,N_6135,N_6848);
xor U11896 (N_11896,N_8355,N_8076);
nor U11897 (N_11897,N_6805,N_5794);
xnor U11898 (N_11898,N_9225,N_5627);
nor U11899 (N_11899,N_9496,N_5713);
xnor U11900 (N_11900,N_5419,N_8236);
xor U11901 (N_11901,N_5883,N_9330);
or U11902 (N_11902,N_9877,N_6141);
nand U11903 (N_11903,N_8842,N_6799);
nand U11904 (N_11904,N_6007,N_8358);
or U11905 (N_11905,N_6350,N_6907);
nand U11906 (N_11906,N_7759,N_8597);
xnor U11907 (N_11907,N_7989,N_9552);
and U11908 (N_11908,N_7825,N_6003);
nand U11909 (N_11909,N_6081,N_6080);
xor U11910 (N_11910,N_8209,N_7844);
nor U11911 (N_11911,N_9994,N_9117);
or U11912 (N_11912,N_9143,N_6913);
nand U11913 (N_11913,N_8480,N_8952);
or U11914 (N_11914,N_5461,N_7487);
nor U11915 (N_11915,N_6423,N_7049);
or U11916 (N_11916,N_6702,N_8396);
nor U11917 (N_11917,N_8893,N_7847);
and U11918 (N_11918,N_7405,N_6283);
nor U11919 (N_11919,N_5628,N_9845);
xor U11920 (N_11920,N_6182,N_6433);
nor U11921 (N_11921,N_6969,N_6178);
nor U11922 (N_11922,N_8827,N_7456);
xnor U11923 (N_11923,N_8533,N_6208);
nand U11924 (N_11924,N_6296,N_7867);
nand U11925 (N_11925,N_5737,N_9093);
nand U11926 (N_11926,N_8469,N_5343);
nor U11927 (N_11927,N_8269,N_5808);
and U11928 (N_11928,N_8416,N_8256);
nand U11929 (N_11929,N_9596,N_8242);
nor U11930 (N_11930,N_9276,N_9071);
xor U11931 (N_11931,N_5581,N_6393);
and U11932 (N_11932,N_8207,N_8392);
or U11933 (N_11933,N_6385,N_9631);
nor U11934 (N_11934,N_9085,N_9801);
nand U11935 (N_11935,N_6639,N_6068);
or U11936 (N_11936,N_8250,N_7689);
nand U11937 (N_11937,N_9611,N_9520);
xnor U11938 (N_11938,N_9098,N_8473);
and U11939 (N_11939,N_8632,N_9188);
nand U11940 (N_11940,N_8913,N_5199);
and U11941 (N_11941,N_9031,N_6348);
or U11942 (N_11942,N_7438,N_6716);
xor U11943 (N_11943,N_7694,N_6254);
xnor U11944 (N_11944,N_9025,N_8134);
xnor U11945 (N_11945,N_8690,N_6610);
nor U11946 (N_11946,N_8455,N_6489);
and U11947 (N_11947,N_9365,N_8719);
and U11948 (N_11948,N_9483,N_6878);
and U11949 (N_11949,N_5933,N_9218);
xor U11950 (N_11950,N_6484,N_5363);
nor U11951 (N_11951,N_5241,N_6608);
nor U11952 (N_11952,N_8172,N_9437);
and U11953 (N_11953,N_5909,N_8286);
or U11954 (N_11954,N_5248,N_8652);
nor U11955 (N_11955,N_8091,N_8572);
or U11956 (N_11956,N_6287,N_5333);
xnor U11957 (N_11957,N_7051,N_8874);
nor U11958 (N_11958,N_6587,N_5245);
or U11959 (N_11959,N_5072,N_6424);
or U11960 (N_11960,N_5471,N_5967);
nor U11961 (N_11961,N_6796,N_8665);
and U11962 (N_11962,N_9677,N_9173);
or U11963 (N_11963,N_8251,N_8606);
and U11964 (N_11964,N_8394,N_8479);
and U11965 (N_11965,N_8523,N_7703);
xnor U11966 (N_11966,N_8324,N_7529);
or U11967 (N_11967,N_9917,N_5942);
and U11968 (N_11968,N_9533,N_6820);
and U11969 (N_11969,N_9951,N_7676);
xor U11970 (N_11970,N_9055,N_9038);
and U11971 (N_11971,N_9386,N_7455);
nand U11972 (N_11972,N_7122,N_9126);
nand U11973 (N_11973,N_6693,N_9221);
and U11974 (N_11974,N_5488,N_6627);
nor U11975 (N_11975,N_7718,N_6982);
and U11976 (N_11976,N_7468,N_5409);
and U11977 (N_11977,N_8381,N_7001);
or U11978 (N_11978,N_6816,N_9176);
and U11979 (N_11979,N_7780,N_7685);
and U11980 (N_11980,N_5437,N_5510);
or U11981 (N_11981,N_9241,N_6274);
nor U11982 (N_11982,N_9751,N_9742);
and U11983 (N_11983,N_6911,N_7371);
nand U11984 (N_11984,N_8771,N_9344);
nor U11985 (N_11985,N_6192,N_7890);
or U11986 (N_11986,N_7807,N_7490);
and U11987 (N_11987,N_7218,N_8763);
nand U11988 (N_11988,N_7719,N_9352);
xnor U11989 (N_11989,N_6451,N_6704);
nand U11990 (N_11990,N_9911,N_9376);
xnor U11991 (N_11991,N_9405,N_5433);
or U11992 (N_11992,N_8631,N_7342);
and U11993 (N_11993,N_9498,N_6371);
xor U11994 (N_11994,N_8265,N_6372);
and U11995 (N_11995,N_5420,N_6903);
nor U11996 (N_11996,N_9345,N_8243);
nand U11997 (N_11997,N_8081,N_7856);
nor U11998 (N_11998,N_9477,N_7554);
nand U11999 (N_11999,N_6613,N_9024);
or U12000 (N_12000,N_6901,N_7837);
xor U12001 (N_12001,N_5006,N_8851);
and U12002 (N_12002,N_6545,N_9428);
or U12003 (N_12003,N_6939,N_6882);
or U12004 (N_12004,N_6039,N_5637);
and U12005 (N_12005,N_5574,N_8924);
nor U12006 (N_12006,N_6442,N_8427);
xor U12007 (N_12007,N_7330,N_5317);
xnor U12008 (N_12008,N_5215,N_5155);
nor U12009 (N_12009,N_8710,N_9037);
and U12010 (N_12010,N_5313,N_7313);
nand U12011 (N_12011,N_9452,N_7000);
or U12012 (N_12012,N_6171,N_8155);
nand U12013 (N_12013,N_7876,N_8919);
or U12014 (N_12014,N_8699,N_6260);
or U12015 (N_12015,N_8360,N_8860);
xnor U12016 (N_12016,N_8288,N_9053);
nand U12017 (N_12017,N_8221,N_7987);
nor U12018 (N_12018,N_7848,N_7482);
and U12019 (N_12019,N_8108,N_7542);
xor U12020 (N_12020,N_6290,N_7457);
and U12021 (N_12021,N_8789,N_5882);
xor U12022 (N_12022,N_5520,N_5550);
nor U12023 (N_12023,N_6884,N_8626);
nor U12024 (N_12024,N_7423,N_8517);
or U12025 (N_12025,N_7472,N_6968);
nor U12026 (N_12026,N_6337,N_5750);
nor U12027 (N_12027,N_7067,N_9857);
xnor U12028 (N_12028,N_9323,N_9159);
and U12029 (N_12029,N_7018,N_5301);
nand U12030 (N_12030,N_5708,N_7626);
nand U12031 (N_12031,N_5636,N_5639);
xor U12032 (N_12032,N_8196,N_7259);
xnor U12033 (N_12033,N_6437,N_9906);
xor U12034 (N_12034,N_7184,N_9772);
xnor U12035 (N_12035,N_5589,N_6586);
or U12036 (N_12036,N_7252,N_6028);
or U12037 (N_12037,N_6236,N_6123);
and U12038 (N_12038,N_6149,N_5853);
or U12039 (N_12039,N_6979,N_5769);
nand U12040 (N_12040,N_5785,N_5007);
and U12041 (N_12041,N_7287,N_6059);
and U12042 (N_12042,N_9021,N_5149);
xor U12043 (N_12043,N_6011,N_5969);
nor U12044 (N_12044,N_5390,N_5497);
and U12045 (N_12045,N_7147,N_5949);
and U12046 (N_12046,N_6995,N_8502);
xnor U12047 (N_12047,N_7242,N_8474);
and U12048 (N_12048,N_9449,N_8574);
or U12049 (N_12049,N_6641,N_6585);
or U12050 (N_12050,N_9263,N_5679);
and U12051 (N_12051,N_6532,N_8008);
and U12052 (N_12052,N_7819,N_8391);
xor U12053 (N_12053,N_7473,N_6958);
and U12054 (N_12054,N_5284,N_5776);
xor U12055 (N_12055,N_7170,N_8790);
or U12056 (N_12056,N_9371,N_6159);
or U12057 (N_12057,N_8425,N_6745);
xor U12058 (N_12058,N_8030,N_7570);
xor U12059 (N_12059,N_9347,N_6671);
and U12060 (N_12060,N_8613,N_7945);
and U12061 (N_12061,N_7275,N_9974);
nand U12062 (N_12062,N_8861,N_8748);
nor U12063 (N_12063,N_9501,N_8676);
xor U12064 (N_12064,N_6899,N_6601);
nor U12065 (N_12065,N_6731,N_8016);
and U12066 (N_12066,N_6062,N_5903);
or U12067 (N_12067,N_8972,N_7183);
and U12068 (N_12068,N_8064,N_7737);
nand U12069 (N_12069,N_8038,N_7642);
xor U12070 (N_12070,N_8452,N_7186);
nor U12071 (N_12071,N_9086,N_7832);
xor U12072 (N_12072,N_6542,N_5035);
or U12073 (N_12073,N_5075,N_9197);
and U12074 (N_12074,N_5829,N_7365);
nor U12075 (N_12075,N_8150,N_7654);
nor U12076 (N_12076,N_8885,N_9433);
and U12077 (N_12077,N_8981,N_6966);
xor U12078 (N_12078,N_5731,N_5361);
and U12079 (N_12079,N_7816,N_8198);
xnor U12080 (N_12080,N_9256,N_6258);
nand U12081 (N_12081,N_7900,N_9954);
nand U12082 (N_12082,N_7992,N_9650);
or U12083 (N_12083,N_7904,N_5252);
nor U12084 (N_12084,N_5203,N_9566);
and U12085 (N_12085,N_9715,N_5466);
nand U12086 (N_12086,N_9500,N_6166);
and U12087 (N_12087,N_8110,N_6112);
nand U12088 (N_12088,N_5572,N_8182);
nand U12089 (N_12089,N_9175,N_6723);
nor U12090 (N_12090,N_5376,N_5872);
xnor U12091 (N_12091,N_8362,N_5415);
xor U12092 (N_12092,N_6902,N_5816);
and U12093 (N_12093,N_6076,N_9975);
nor U12094 (N_12094,N_5610,N_5080);
and U12095 (N_12095,N_6503,N_6748);
xnor U12096 (N_12096,N_6382,N_9418);
nor U12097 (N_12097,N_7381,N_5279);
and U12098 (N_12098,N_8127,N_6180);
nor U12099 (N_12099,N_7775,N_5028);
and U12100 (N_12100,N_7618,N_9753);
xnor U12101 (N_12101,N_7368,N_5422);
or U12102 (N_12102,N_7745,N_8412);
and U12103 (N_12103,N_9681,N_9438);
xnor U12104 (N_12104,N_7153,N_6813);
xor U12105 (N_12105,N_5701,N_7750);
or U12106 (N_12106,N_9656,N_6655);
or U12107 (N_12107,N_7297,N_7815);
or U12108 (N_12108,N_8868,N_7312);
or U12109 (N_12109,N_6277,N_6981);
xor U12110 (N_12110,N_9797,N_8262);
xor U12111 (N_12111,N_7048,N_5462);
nor U12112 (N_12112,N_9879,N_9303);
nor U12113 (N_12113,N_5063,N_7178);
nand U12114 (N_12114,N_7649,N_7740);
nand U12115 (N_12115,N_8363,N_5201);
nand U12116 (N_12116,N_6332,N_7207);
nor U12117 (N_12117,N_5107,N_5137);
or U12118 (N_12118,N_8674,N_6683);
and U12119 (N_12119,N_6637,N_8083);
xnor U12120 (N_12120,N_5131,N_6941);
xnor U12121 (N_12121,N_5648,N_8297);
or U12122 (N_12122,N_9740,N_9006);
nor U12123 (N_12123,N_7201,N_9924);
nand U12124 (N_12124,N_9862,N_8920);
nor U12125 (N_12125,N_5071,N_5765);
or U12126 (N_12126,N_6152,N_8668);
and U12127 (N_12127,N_7606,N_5385);
nand U12128 (N_12128,N_7164,N_5223);
nand U12129 (N_12129,N_6322,N_8181);
and U12130 (N_12130,N_7374,N_5291);
nand U12131 (N_12131,N_9525,N_8840);
xnor U12132 (N_12132,N_6665,N_9294);
or U12133 (N_12133,N_8001,N_6615);
xnor U12134 (N_12134,N_5436,N_8567);
nand U12135 (N_12135,N_9095,N_9448);
nor U12136 (N_12136,N_5811,N_8622);
nor U12137 (N_12137,N_8953,N_5047);
or U12138 (N_12138,N_5747,N_8451);
nor U12139 (N_12139,N_5753,N_6733);
nor U12140 (N_12140,N_9291,N_6614);
nor U12141 (N_12141,N_8672,N_7574);
nor U12142 (N_12142,N_9519,N_5559);
or U12143 (N_12143,N_8170,N_9828);
xor U12144 (N_12144,N_7103,N_7271);
nor U12145 (N_12145,N_8545,N_6292);
nor U12146 (N_12146,N_7403,N_7891);
xor U12147 (N_12147,N_5892,N_8232);
nor U12148 (N_12148,N_9644,N_6626);
xor U12149 (N_12149,N_9064,N_6391);
nand U12150 (N_12150,N_8946,N_8051);
or U12151 (N_12151,N_9502,N_9553);
or U12152 (N_12152,N_7549,N_8304);
or U12153 (N_12153,N_6597,N_9928);
nand U12154 (N_12154,N_6747,N_5100);
xor U12155 (N_12155,N_6930,N_7391);
and U12156 (N_12156,N_6404,N_8153);
nand U12157 (N_12157,N_9976,N_5502);
nand U12158 (N_12158,N_8785,N_7441);
nand U12159 (N_12159,N_5768,N_6570);
or U12160 (N_12160,N_9429,N_5710);
nand U12161 (N_12161,N_6342,N_5661);
nor U12162 (N_12162,N_9833,N_8923);
nor U12163 (N_12163,N_6078,N_7599);
nor U12164 (N_12164,N_8333,N_8641);
nor U12165 (N_12165,N_6387,N_5160);
and U12166 (N_12166,N_9181,N_8424);
xnor U12167 (N_12167,N_8444,N_9254);
or U12168 (N_12168,N_9199,N_5987);
xor U12169 (N_12169,N_5519,N_9763);
nand U12170 (N_12170,N_7699,N_6935);
or U12171 (N_12171,N_6851,N_9737);
or U12172 (N_12172,N_6520,N_5294);
and U12173 (N_12173,N_5764,N_8957);
and U12174 (N_12174,N_5458,N_6269);
or U12175 (N_12175,N_8492,N_7875);
nand U12176 (N_12176,N_8466,N_7422);
or U12177 (N_12177,N_8118,N_7949);
xor U12178 (N_12178,N_5843,N_6568);
xnor U12179 (N_12179,N_8547,N_9927);
nor U12180 (N_12180,N_9481,N_5974);
xor U12181 (N_12181,N_8594,N_7045);
nor U12182 (N_12182,N_5356,N_6539);
xnor U12183 (N_12183,N_9230,N_6547);
nand U12184 (N_12184,N_6842,N_9946);
nand U12185 (N_12185,N_9088,N_5362);
xnor U12186 (N_12186,N_7668,N_7728);
or U12187 (N_12187,N_7879,N_9529);
nor U12188 (N_12188,N_6905,N_9840);
nor U12189 (N_12189,N_9793,N_8057);
nor U12190 (N_12190,N_8578,N_9393);
and U12191 (N_12191,N_9926,N_9855);
or U12192 (N_12192,N_5711,N_6086);
or U12193 (N_12193,N_7108,N_9686);
nor U12194 (N_12194,N_6376,N_7016);
xor U12195 (N_12195,N_7367,N_5805);
nand U12196 (N_12196,N_8272,N_5910);
and U12197 (N_12197,N_9947,N_5470);
xor U12198 (N_12198,N_6463,N_8310);
xnor U12199 (N_12199,N_8760,N_5320);
or U12200 (N_12200,N_5463,N_5051);
xnor U12201 (N_12201,N_9457,N_9102);
xor U12202 (N_12202,N_6473,N_9841);
xor U12203 (N_12203,N_6035,N_7696);
nor U12204 (N_12204,N_6162,N_9322);
xnor U12205 (N_12205,N_5211,N_6651);
nand U12206 (N_12206,N_7786,N_7246);
nand U12207 (N_12207,N_8730,N_5348);
and U12208 (N_12208,N_8160,N_6339);
and U12209 (N_12209,N_6897,N_6106);
nor U12210 (N_12210,N_5027,N_9302);
nor U12211 (N_12211,N_5722,N_6347);
nor U12212 (N_12212,N_9305,N_6435);
xor U12213 (N_12213,N_7224,N_6756);
xor U12214 (N_12214,N_5907,N_9614);
and U12215 (N_12215,N_8596,N_7019);
xor U12216 (N_12216,N_7389,N_8765);
nor U12217 (N_12217,N_7752,N_6308);
nor U12218 (N_12218,N_8743,N_5475);
xnor U12219 (N_12219,N_5828,N_6604);
nor U12220 (N_12220,N_5733,N_6204);
and U12221 (N_12221,N_6951,N_5911);
nand U12222 (N_12222,N_6395,N_8704);
xor U12223 (N_12223,N_7944,N_9005);
nor U12224 (N_12224,N_8312,N_9099);
and U12225 (N_12225,N_9980,N_9684);
nor U12226 (N_12226,N_7840,N_9804);
xnor U12227 (N_12227,N_9586,N_6226);
nor U12228 (N_12228,N_8494,N_7014);
and U12229 (N_12229,N_9852,N_7590);
and U12230 (N_12230,N_9372,N_6018);
nor U12231 (N_12231,N_7370,N_6104);
or U12232 (N_12232,N_9337,N_8815);
nor U12233 (N_12233,N_9555,N_5561);
or U12234 (N_12234,N_9131,N_6876);
nand U12235 (N_12235,N_7107,N_6727);
xnor U12236 (N_12236,N_8015,N_8810);
or U12237 (N_12237,N_6317,N_8806);
nor U12238 (N_12238,N_9426,N_6771);
or U12239 (N_12239,N_7893,N_5157);
or U12240 (N_12240,N_8514,N_9824);
nor U12241 (N_12241,N_7181,N_5779);
nand U12242 (N_12242,N_6266,N_5123);
or U12243 (N_12243,N_8373,N_8756);
nand U12244 (N_12244,N_8888,N_7105);
nand U12245 (N_12245,N_8225,N_8709);
nor U12246 (N_12246,N_5164,N_7595);
or U12247 (N_12247,N_8648,N_5736);
xnor U12248 (N_12248,N_7995,N_6755);
xnor U12249 (N_12249,N_6581,N_9874);
or U12250 (N_12250,N_6179,N_8684);
or U12251 (N_12251,N_9180,N_9771);
xor U12252 (N_12252,N_9764,N_6560);
or U12253 (N_12253,N_6519,N_5196);
and U12254 (N_12254,N_6685,N_6759);
nand U12255 (N_12255,N_7609,N_7156);
nor U12256 (N_12256,N_8732,N_5408);
nor U12257 (N_12257,N_8535,N_8334);
and U12258 (N_12258,N_5305,N_7072);
nor U12259 (N_12259,N_8895,N_6988);
or U12260 (N_12260,N_9282,N_9417);
and U12261 (N_12261,N_9967,N_8352);
nor U12262 (N_12262,N_6403,N_8338);
or U12263 (N_12263,N_7702,N_7998);
nand U12264 (N_12264,N_7239,N_7948);
xor U12265 (N_12265,N_9148,N_7010);
and U12266 (N_12266,N_6087,N_7285);
and U12267 (N_12267,N_8164,N_5876);
nand U12268 (N_12268,N_5127,N_6268);
and U12269 (N_12269,N_9507,N_7964);
nor U12270 (N_12270,N_6766,N_5657);
or U12271 (N_12271,N_6511,N_6721);
nand U12272 (N_12272,N_6837,N_5641);
xor U12273 (N_12273,N_6690,N_6184);
nand U12274 (N_12274,N_8044,N_6029);
and U12275 (N_12275,N_8896,N_9789);
or U12276 (N_12276,N_8383,N_9353);
xor U12277 (N_12277,N_5220,N_9407);
nand U12278 (N_12278,N_8282,N_7251);
xnor U12279 (N_12279,N_9745,N_5576);
nor U12280 (N_12280,N_6647,N_8319);
nand U12281 (N_12281,N_9164,N_8834);
xor U12282 (N_12282,N_8935,N_6530);
nor U12283 (N_12283,N_9847,N_9667);
xor U12284 (N_12284,N_9829,N_8152);
and U12285 (N_12285,N_8871,N_6048);
xnor U12286 (N_12286,N_7988,N_8967);
nor U12287 (N_12287,N_7809,N_8950);
nor U12288 (N_12288,N_8067,N_9200);
xor U12289 (N_12289,N_9150,N_9203);
and U12290 (N_12290,N_5625,N_6010);
nor U12291 (N_12291,N_6267,N_8116);
xnor U12292 (N_12292,N_6692,N_9145);
nand U12293 (N_12293,N_9487,N_9629);
nand U12294 (N_12294,N_9943,N_5584);
or U12295 (N_12295,N_7705,N_8640);
nor U12296 (N_12296,N_5378,N_9030);
xor U12297 (N_12297,N_5651,N_8854);
xnor U12298 (N_12298,N_5536,N_6625);
nor U12299 (N_12299,N_5781,N_5538);
xor U12300 (N_12300,N_8693,N_8835);
xnor U12301 (N_12301,N_8079,N_5621);
and U12302 (N_12302,N_5566,N_6574);
xnor U12303 (N_12303,N_7075,N_8943);
nor U12304 (N_12304,N_5617,N_8980);
nor U12305 (N_12305,N_7050,N_8013);
nand U12306 (N_12306,N_7805,N_6870);
nand U12307 (N_12307,N_7731,N_5788);
nand U12308 (N_12308,N_6191,N_9440);
nor U12309 (N_12309,N_9096,N_8280);
or U12310 (N_12310,N_5827,N_6338);
nor U12311 (N_12311,N_8518,N_5371);
nor U12312 (N_12312,N_6890,N_9526);
and U12313 (N_12313,N_8557,N_8467);
xnor U12314 (N_12314,N_9374,N_5535);
nand U12315 (N_12315,N_8382,N_8461);
or U12316 (N_12316,N_9844,N_8047);
and U12317 (N_12317,N_6331,N_6490);
nand U12318 (N_12318,N_7443,N_8670);
xor U12319 (N_12319,N_8571,N_6194);
nor U12320 (N_12320,N_7950,N_5213);
or U12321 (N_12321,N_5125,N_5400);
and U12322 (N_12322,N_7897,N_9387);
xor U12323 (N_12323,N_7631,N_7547);
nor U12324 (N_12324,N_5023,N_9383);
nor U12325 (N_12325,N_7031,N_8610);
or U12326 (N_12326,N_6436,N_6165);
or U12327 (N_12327,N_8195,N_7394);
or U12328 (N_12328,N_6918,N_5919);
and U12329 (N_12329,N_8361,N_9589);
and U12330 (N_12330,N_7255,N_8605);
and U12331 (N_12331,N_5551,N_9049);
or U12332 (N_12332,N_6512,N_9902);
and U12333 (N_12333,N_9090,N_5801);
xor U12334 (N_12334,N_8930,N_5457);
or U12335 (N_12335,N_5000,N_7427);
and U12336 (N_12336,N_5337,N_5950);
nand U12337 (N_12337,N_9000,N_7808);
and U12338 (N_12338,N_7339,N_9661);
and U12339 (N_12339,N_8165,N_9671);
nand U12340 (N_12340,N_7047,N_8376);
nor U12341 (N_12341,N_6411,N_6852);
or U12342 (N_12342,N_6513,N_8762);
nand U12343 (N_12343,N_8685,N_9304);
nor U12344 (N_12344,N_9346,N_6791);
and U12345 (N_12345,N_6252,N_7439);
or U12346 (N_12346,N_9863,N_7738);
nand U12347 (N_12347,N_5856,N_6780);
or U12348 (N_12348,N_8458,N_8497);
nor U12349 (N_12349,N_7185,N_8576);
xor U12350 (N_12350,N_8194,N_5727);
and U12351 (N_12351,N_6095,N_6900);
xnor U12352 (N_12352,N_5804,N_7704);
and U12353 (N_12353,N_9392,N_6961);
xnor U12354 (N_12354,N_8577,N_8244);
and U12355 (N_12355,N_8725,N_7575);
nor U12356 (N_12356,N_7377,N_8865);
and U12357 (N_12357,N_7250,N_5232);
xor U12358 (N_12358,N_5973,N_8122);
nand U12359 (N_12359,N_7622,N_6055);
nand U12360 (N_12360,N_7709,N_8234);
nor U12361 (N_12361,N_7489,N_7171);
xor U12362 (N_12362,N_7380,N_5210);
nand U12363 (N_12363,N_5964,N_7721);
nand U12364 (N_12364,N_8061,N_9036);
xnor U12365 (N_12365,N_7774,N_8434);
and U12366 (N_12366,N_6272,N_7596);
nand U12367 (N_12367,N_9092,N_6675);
xor U12368 (N_12368,N_6917,N_6492);
or U12369 (N_12369,N_8446,N_6445);
and U12370 (N_12370,N_7634,N_6945);
nand U12371 (N_12371,N_7133,N_8969);
xnor U12372 (N_12372,N_9570,N_6868);
or U12373 (N_12373,N_6662,N_6448);
and U12374 (N_12374,N_8034,N_5234);
xnor U12375 (N_12375,N_7882,N_9120);
xor U12376 (N_12376,N_8985,N_9509);
or U12377 (N_12377,N_8218,N_6895);
nand U12378 (N_12378,N_5755,N_9442);
and U12379 (N_12379,N_6508,N_5093);
xor U12380 (N_12380,N_8697,N_5598);
xnor U12381 (N_12381,N_7005,N_7777);
nor U12382 (N_12382,N_8528,N_8445);
xor U12383 (N_12383,N_8592,N_5379);
xnor U12384 (N_12384,N_6088,N_5235);
nand U12385 (N_12385,N_5296,N_8879);
and U12386 (N_12386,N_8167,N_8147);
nor U12387 (N_12387,N_5286,N_5981);
nand U12388 (N_12388,N_7725,N_9981);
xnor U12389 (N_12389,N_8292,N_9913);
xor U12390 (N_12390,N_8963,N_9988);
nor U12391 (N_12391,N_9646,N_7466);
nor U12392 (N_12392,N_9630,N_6462);
and U12393 (N_12393,N_7793,N_8999);
and U12394 (N_12394,N_5388,N_7068);
nand U12395 (N_12395,N_8129,N_7910);
or U12396 (N_12396,N_5734,N_9937);
xor U12397 (N_12397,N_7430,N_6892);
or U12398 (N_12398,N_7941,N_8019);
nand U12399 (N_12399,N_9792,N_5556);
and U12400 (N_12400,N_9454,N_5562);
xor U12401 (N_12401,N_9379,N_8350);
xor U12402 (N_12402,N_5983,N_5944);
or U12403 (N_12403,N_8442,N_5749);
xnor U12404 (N_12404,N_8240,N_9690);
xnor U12405 (N_12405,N_8464,N_7888);
or U12406 (N_12406,N_9591,N_9700);
nand U12407 (N_12407,N_7611,N_7946);
xnor U12408 (N_12408,N_5302,N_9373);
or U12409 (N_12409,N_7202,N_7698);
and U12410 (N_12410,N_9446,N_8742);
and U12411 (N_12411,N_6324,N_6802);
and U12412 (N_12412,N_6650,N_5687);
nor U12413 (N_12413,N_5720,N_7324);
or U12414 (N_12414,N_6085,N_6875);
nor U12415 (N_12415,N_8586,N_6167);
nor U12416 (N_12416,N_6669,N_6877);
nor U12417 (N_12417,N_5452,N_8179);
nand U12418 (N_12418,N_8253,N_9787);
and U12419 (N_12419,N_7027,N_9560);
and U12420 (N_12420,N_8857,N_8918);
or U12421 (N_12421,N_9950,N_7280);
or U12422 (N_12422,N_5937,N_7767);
and U12423 (N_12423,N_7791,N_7130);
or U12424 (N_12424,N_9658,N_6494);
nand U12425 (N_12425,N_9836,N_9087);
nand U12426 (N_12426,N_6993,N_7442);
nor U12427 (N_12427,N_9234,N_5852);
xor U12428 (N_12428,N_7121,N_9141);
or U12429 (N_12429,N_5560,N_9207);
xnor U12430 (N_12430,N_6111,N_8296);
and U12431 (N_12431,N_7217,N_9582);
nand U12432 (N_12432,N_7451,N_9685);
or U12433 (N_12433,N_5487,N_7205);
nand U12434 (N_12434,N_9149,N_5588);
nor U12435 (N_12435,N_6270,N_6496);
nand U12436 (N_12436,N_7355,N_5693);
or U12437 (N_12437,N_6225,N_9987);
or U12438 (N_12438,N_7138,N_8066);
xnor U12439 (N_12439,N_8525,N_7086);
nand U12440 (N_12440,N_8441,N_8936);
xor U12441 (N_12441,N_9269,N_5614);
nand U12442 (N_12442,N_5515,N_8595);
xnor U12443 (N_12443,N_5227,N_7039);
xor U12444 (N_12444,N_7881,N_8853);
xor U12445 (N_12445,N_9695,N_6002);
xnor U12446 (N_12446,N_9573,N_6233);
nor U12447 (N_12447,N_5467,N_7922);
nand U12448 (N_12448,N_7520,N_9528);
and U12449 (N_12449,N_5447,N_8660);
and U12450 (N_12450,N_6472,N_7323);
and U12451 (N_12451,N_8146,N_7579);
nor U12452 (N_12452,N_6301,N_7749);
or U12453 (N_12453,N_9692,N_9224);
nor U12454 (N_12454,N_7375,N_5179);
or U12455 (N_12455,N_9873,N_8428);
nor U12456 (N_12456,N_5293,N_5143);
and U12457 (N_12457,N_9377,N_9463);
nor U12458 (N_12458,N_7921,N_7254);
or U12459 (N_12459,N_9583,N_7042);
and U12460 (N_12460,N_6360,N_6599);
xor U12461 (N_12461,N_6243,N_7927);
and U12462 (N_12462,N_5699,N_6375);
and U12463 (N_12463,N_9171,N_9957);
nand U12464 (N_12464,N_6596,N_9632);
nor U12465 (N_12465,N_6933,N_7332);
nor U12466 (N_12466,N_7969,N_8264);
xnor U12467 (N_12467,N_7354,N_6926);
nand U12468 (N_12468,N_9568,N_8448);
xnor U12469 (N_12469,N_9198,N_8048);
or U12470 (N_12470,N_8332,N_9174);
xnor U12471 (N_12471,N_7338,N_7064);
nor U12472 (N_12472,N_9991,N_7126);
and U12473 (N_12473,N_6091,N_6070);
nor U12474 (N_12474,N_5357,N_9227);
nand U12475 (N_12475,N_5078,N_8698);
xor U12476 (N_12476,N_7543,N_8938);
nand U12477 (N_12477,N_6846,N_5646);
nor U12478 (N_12478,N_6526,N_8283);
nor U12479 (N_12479,N_5499,N_7151);
nor U12480 (N_12480,N_7053,N_7630);
xor U12481 (N_12481,N_8345,N_6638);
nand U12482 (N_12482,N_9876,N_9524);
and U12483 (N_12483,N_8414,N_9775);
or U12484 (N_12484,N_6673,N_6493);
nand U12485 (N_12485,N_8045,N_6214);
or U12486 (N_12486,N_9168,N_7510);
xnor U12487 (N_12487,N_6409,N_8329);
xnor U12488 (N_12488,N_8737,N_8754);
xnor U12489 (N_12489,N_6787,N_7880);
xnor U12490 (N_12490,N_8682,N_7421);
or U12491 (N_12491,N_7943,N_9660);
nand U12492 (N_12492,N_8020,N_8706);
nor U12493 (N_12493,N_8154,N_7166);
or U12494 (N_12494,N_8486,N_7134);
and U12495 (N_12495,N_7957,N_5144);
xnor U12496 (N_12496,N_5132,N_6778);
or U12497 (N_12497,N_7760,N_7387);
nor U12498 (N_12498,N_5777,N_6580);
nor U12499 (N_12499,N_7230,N_6098);
and U12500 (N_12500,N_7945,N_6268);
nand U12501 (N_12501,N_6946,N_6723);
nand U12502 (N_12502,N_9668,N_8988);
or U12503 (N_12503,N_5126,N_5003);
xnor U12504 (N_12504,N_6412,N_9280);
xnor U12505 (N_12505,N_9028,N_5017);
and U12506 (N_12506,N_6975,N_8958);
nor U12507 (N_12507,N_9870,N_5277);
or U12508 (N_12508,N_8192,N_9082);
or U12509 (N_12509,N_6655,N_5166);
nand U12510 (N_12510,N_5647,N_6182);
nor U12511 (N_12511,N_5322,N_9662);
nor U12512 (N_12512,N_6995,N_6561);
nand U12513 (N_12513,N_7262,N_6279);
nand U12514 (N_12514,N_7495,N_5162);
or U12515 (N_12515,N_5646,N_6309);
nor U12516 (N_12516,N_7027,N_6212);
and U12517 (N_12517,N_9326,N_9933);
xnor U12518 (N_12518,N_6607,N_6520);
nand U12519 (N_12519,N_9835,N_7836);
and U12520 (N_12520,N_7845,N_9968);
and U12521 (N_12521,N_8276,N_6068);
xnor U12522 (N_12522,N_5138,N_9706);
or U12523 (N_12523,N_9354,N_9776);
or U12524 (N_12524,N_5240,N_6445);
or U12525 (N_12525,N_9461,N_8414);
xnor U12526 (N_12526,N_7061,N_8014);
nand U12527 (N_12527,N_5561,N_7219);
nand U12528 (N_12528,N_7131,N_9111);
xor U12529 (N_12529,N_8612,N_8771);
nand U12530 (N_12530,N_5634,N_7773);
xor U12531 (N_12531,N_6935,N_8439);
nor U12532 (N_12532,N_8858,N_8746);
or U12533 (N_12533,N_7592,N_7981);
nor U12534 (N_12534,N_7861,N_5058);
nand U12535 (N_12535,N_7307,N_7761);
xor U12536 (N_12536,N_6501,N_7649);
nor U12537 (N_12537,N_7289,N_6544);
or U12538 (N_12538,N_5421,N_9553);
and U12539 (N_12539,N_8099,N_7847);
and U12540 (N_12540,N_9427,N_9127);
xnor U12541 (N_12541,N_5110,N_6921);
and U12542 (N_12542,N_6643,N_9381);
nor U12543 (N_12543,N_6639,N_9727);
or U12544 (N_12544,N_7665,N_8961);
nand U12545 (N_12545,N_5335,N_6718);
xor U12546 (N_12546,N_9380,N_6316);
and U12547 (N_12547,N_5088,N_6314);
and U12548 (N_12548,N_8766,N_6932);
nand U12549 (N_12549,N_8763,N_8128);
and U12550 (N_12550,N_7140,N_5874);
or U12551 (N_12551,N_7149,N_6828);
and U12552 (N_12552,N_8239,N_5464);
and U12553 (N_12553,N_8981,N_5908);
or U12554 (N_12554,N_5240,N_5861);
nand U12555 (N_12555,N_8382,N_7615);
xor U12556 (N_12556,N_9975,N_5529);
nand U12557 (N_12557,N_6542,N_5579);
xor U12558 (N_12558,N_6090,N_7890);
nand U12559 (N_12559,N_5068,N_6646);
nand U12560 (N_12560,N_6151,N_5039);
nand U12561 (N_12561,N_9266,N_7540);
and U12562 (N_12562,N_6552,N_7322);
or U12563 (N_12563,N_9169,N_8009);
and U12564 (N_12564,N_5672,N_6535);
xnor U12565 (N_12565,N_9432,N_8574);
or U12566 (N_12566,N_5707,N_6869);
nand U12567 (N_12567,N_5439,N_7650);
or U12568 (N_12568,N_9571,N_6760);
or U12569 (N_12569,N_9539,N_9284);
or U12570 (N_12570,N_9101,N_9519);
nor U12571 (N_12571,N_7886,N_7160);
nand U12572 (N_12572,N_7916,N_5649);
nand U12573 (N_12573,N_6277,N_6336);
and U12574 (N_12574,N_7626,N_6913);
and U12575 (N_12575,N_8073,N_9688);
xnor U12576 (N_12576,N_9659,N_9460);
or U12577 (N_12577,N_5684,N_6662);
nand U12578 (N_12578,N_6034,N_7982);
or U12579 (N_12579,N_5441,N_5391);
or U12580 (N_12580,N_8902,N_9990);
or U12581 (N_12581,N_5125,N_6022);
nor U12582 (N_12582,N_6599,N_7770);
and U12583 (N_12583,N_9080,N_8887);
nand U12584 (N_12584,N_8177,N_5619);
or U12585 (N_12585,N_5536,N_5350);
and U12586 (N_12586,N_9918,N_5592);
or U12587 (N_12587,N_8551,N_8089);
and U12588 (N_12588,N_6270,N_6099);
nand U12589 (N_12589,N_5841,N_6652);
nand U12590 (N_12590,N_7567,N_8480);
and U12591 (N_12591,N_5104,N_7741);
xor U12592 (N_12592,N_6637,N_9749);
nand U12593 (N_12593,N_7353,N_9999);
xor U12594 (N_12594,N_8408,N_9424);
nand U12595 (N_12595,N_6793,N_7459);
nand U12596 (N_12596,N_7681,N_6507);
and U12597 (N_12597,N_9517,N_9644);
and U12598 (N_12598,N_5189,N_8139);
xnor U12599 (N_12599,N_6306,N_7733);
and U12600 (N_12600,N_7386,N_6966);
nand U12601 (N_12601,N_7638,N_5128);
nand U12602 (N_12602,N_9386,N_5357);
or U12603 (N_12603,N_8058,N_9907);
xor U12604 (N_12604,N_8715,N_6025);
and U12605 (N_12605,N_8906,N_6928);
nor U12606 (N_12606,N_5645,N_8907);
nand U12607 (N_12607,N_9203,N_6024);
xor U12608 (N_12608,N_8748,N_7122);
nor U12609 (N_12609,N_5091,N_9703);
and U12610 (N_12610,N_8448,N_7155);
and U12611 (N_12611,N_5358,N_5523);
nand U12612 (N_12612,N_6050,N_9610);
xnor U12613 (N_12613,N_9662,N_8968);
nand U12614 (N_12614,N_8688,N_5204);
or U12615 (N_12615,N_8871,N_6634);
nor U12616 (N_12616,N_5600,N_6882);
xor U12617 (N_12617,N_7956,N_9463);
nor U12618 (N_12618,N_6331,N_7699);
nor U12619 (N_12619,N_8629,N_5434);
or U12620 (N_12620,N_7155,N_7766);
or U12621 (N_12621,N_6889,N_5199);
nor U12622 (N_12622,N_9054,N_6979);
or U12623 (N_12623,N_5399,N_9114);
or U12624 (N_12624,N_9746,N_7032);
or U12625 (N_12625,N_8200,N_9907);
xnor U12626 (N_12626,N_6566,N_6671);
and U12627 (N_12627,N_5945,N_5025);
xnor U12628 (N_12628,N_6298,N_8057);
nor U12629 (N_12629,N_5214,N_6538);
nor U12630 (N_12630,N_7929,N_6769);
nor U12631 (N_12631,N_8821,N_8566);
and U12632 (N_12632,N_9080,N_7623);
or U12633 (N_12633,N_7388,N_7046);
and U12634 (N_12634,N_9698,N_7120);
xnor U12635 (N_12635,N_7642,N_5810);
or U12636 (N_12636,N_7630,N_8547);
xnor U12637 (N_12637,N_7285,N_5087);
and U12638 (N_12638,N_9702,N_6715);
nor U12639 (N_12639,N_8254,N_6184);
nor U12640 (N_12640,N_7787,N_7363);
nor U12641 (N_12641,N_8824,N_7021);
nor U12642 (N_12642,N_8612,N_5568);
xor U12643 (N_12643,N_8429,N_9714);
and U12644 (N_12644,N_9447,N_9658);
nor U12645 (N_12645,N_9652,N_9828);
xor U12646 (N_12646,N_6416,N_8449);
nand U12647 (N_12647,N_9239,N_6994);
and U12648 (N_12648,N_9193,N_6565);
or U12649 (N_12649,N_7765,N_8584);
nor U12650 (N_12650,N_9267,N_9008);
nand U12651 (N_12651,N_6298,N_5390);
nand U12652 (N_12652,N_6866,N_7220);
xor U12653 (N_12653,N_5220,N_6315);
or U12654 (N_12654,N_5742,N_6599);
or U12655 (N_12655,N_5283,N_7055);
nand U12656 (N_12656,N_5493,N_5760);
or U12657 (N_12657,N_8361,N_7189);
nand U12658 (N_12658,N_5383,N_9726);
xor U12659 (N_12659,N_8379,N_9041);
nor U12660 (N_12660,N_7770,N_9892);
or U12661 (N_12661,N_9230,N_5787);
and U12662 (N_12662,N_9492,N_6044);
xor U12663 (N_12663,N_5191,N_8201);
xnor U12664 (N_12664,N_5974,N_9966);
nand U12665 (N_12665,N_9434,N_8202);
or U12666 (N_12666,N_7552,N_5713);
or U12667 (N_12667,N_5998,N_9447);
nor U12668 (N_12668,N_5687,N_8669);
nor U12669 (N_12669,N_6785,N_9198);
and U12670 (N_12670,N_9624,N_6093);
nand U12671 (N_12671,N_5386,N_9576);
nand U12672 (N_12672,N_5850,N_7268);
nor U12673 (N_12673,N_7923,N_8904);
xnor U12674 (N_12674,N_7663,N_7054);
nand U12675 (N_12675,N_5162,N_6236);
nor U12676 (N_12676,N_9824,N_5569);
xnor U12677 (N_12677,N_5732,N_6208);
nand U12678 (N_12678,N_7624,N_7672);
nand U12679 (N_12679,N_5484,N_5001);
nor U12680 (N_12680,N_5225,N_9274);
xor U12681 (N_12681,N_9818,N_7864);
nand U12682 (N_12682,N_5050,N_8127);
or U12683 (N_12683,N_9580,N_8943);
nor U12684 (N_12684,N_6155,N_9644);
nor U12685 (N_12685,N_9167,N_8433);
or U12686 (N_12686,N_6328,N_9994);
nor U12687 (N_12687,N_9855,N_6027);
nor U12688 (N_12688,N_7009,N_6319);
nand U12689 (N_12689,N_5505,N_6304);
nor U12690 (N_12690,N_6162,N_6888);
nand U12691 (N_12691,N_9760,N_7483);
xor U12692 (N_12692,N_9703,N_9821);
nand U12693 (N_12693,N_7164,N_9694);
nor U12694 (N_12694,N_7756,N_7235);
and U12695 (N_12695,N_9974,N_5155);
xnor U12696 (N_12696,N_9335,N_8893);
and U12697 (N_12697,N_5336,N_8463);
nand U12698 (N_12698,N_5216,N_9672);
nor U12699 (N_12699,N_5292,N_7571);
nor U12700 (N_12700,N_8153,N_9191);
or U12701 (N_12701,N_9274,N_9447);
nand U12702 (N_12702,N_8731,N_6229);
xor U12703 (N_12703,N_5692,N_8518);
nor U12704 (N_12704,N_5708,N_6140);
xor U12705 (N_12705,N_7854,N_9609);
nor U12706 (N_12706,N_9521,N_9243);
nor U12707 (N_12707,N_8048,N_6512);
or U12708 (N_12708,N_7595,N_9359);
xor U12709 (N_12709,N_5229,N_8626);
xor U12710 (N_12710,N_6341,N_5881);
and U12711 (N_12711,N_5664,N_5861);
nand U12712 (N_12712,N_9696,N_7370);
nand U12713 (N_12713,N_7006,N_9545);
nand U12714 (N_12714,N_5408,N_9873);
xnor U12715 (N_12715,N_9942,N_6958);
nor U12716 (N_12716,N_5945,N_7830);
or U12717 (N_12717,N_8437,N_8322);
nand U12718 (N_12718,N_9555,N_7184);
nand U12719 (N_12719,N_9665,N_8277);
nor U12720 (N_12720,N_5348,N_8151);
nand U12721 (N_12721,N_5300,N_8751);
and U12722 (N_12722,N_9624,N_9794);
or U12723 (N_12723,N_8978,N_8294);
or U12724 (N_12724,N_5298,N_9804);
and U12725 (N_12725,N_6137,N_9975);
xnor U12726 (N_12726,N_7030,N_7139);
xnor U12727 (N_12727,N_5656,N_8445);
xor U12728 (N_12728,N_7783,N_7875);
nor U12729 (N_12729,N_5410,N_9773);
xnor U12730 (N_12730,N_5247,N_7659);
and U12731 (N_12731,N_9182,N_9474);
or U12732 (N_12732,N_5829,N_8722);
xnor U12733 (N_12733,N_8155,N_9485);
nor U12734 (N_12734,N_7142,N_9537);
nor U12735 (N_12735,N_9228,N_9274);
nand U12736 (N_12736,N_6277,N_9529);
nand U12737 (N_12737,N_6595,N_6836);
or U12738 (N_12738,N_5457,N_8192);
and U12739 (N_12739,N_5451,N_7112);
nand U12740 (N_12740,N_6130,N_9293);
or U12741 (N_12741,N_9773,N_5197);
and U12742 (N_12742,N_9020,N_8518);
nor U12743 (N_12743,N_5928,N_7899);
nand U12744 (N_12744,N_5640,N_9890);
and U12745 (N_12745,N_9607,N_5430);
nand U12746 (N_12746,N_5463,N_9326);
xor U12747 (N_12747,N_8872,N_8885);
and U12748 (N_12748,N_9969,N_8959);
xnor U12749 (N_12749,N_8171,N_5445);
and U12750 (N_12750,N_5882,N_6065);
and U12751 (N_12751,N_6365,N_6743);
xnor U12752 (N_12752,N_5895,N_7800);
nor U12753 (N_12753,N_6361,N_6283);
nor U12754 (N_12754,N_9663,N_7089);
or U12755 (N_12755,N_5884,N_8324);
xnor U12756 (N_12756,N_9677,N_5186);
xor U12757 (N_12757,N_9925,N_9129);
or U12758 (N_12758,N_9922,N_9231);
xor U12759 (N_12759,N_8005,N_6434);
or U12760 (N_12760,N_6260,N_8430);
nand U12761 (N_12761,N_7908,N_9037);
xnor U12762 (N_12762,N_8754,N_5993);
and U12763 (N_12763,N_6697,N_9348);
or U12764 (N_12764,N_9267,N_8524);
nor U12765 (N_12765,N_8265,N_7449);
and U12766 (N_12766,N_7392,N_6237);
and U12767 (N_12767,N_7090,N_8555);
nand U12768 (N_12768,N_6504,N_9134);
and U12769 (N_12769,N_5863,N_8339);
or U12770 (N_12770,N_7650,N_7117);
xnor U12771 (N_12771,N_7907,N_5811);
and U12772 (N_12772,N_9457,N_5533);
xnor U12773 (N_12773,N_9502,N_5680);
and U12774 (N_12774,N_5434,N_7029);
or U12775 (N_12775,N_8111,N_6484);
or U12776 (N_12776,N_8442,N_5009);
and U12777 (N_12777,N_6359,N_6724);
nor U12778 (N_12778,N_8435,N_8719);
nor U12779 (N_12779,N_5374,N_6740);
xnor U12780 (N_12780,N_5752,N_5702);
or U12781 (N_12781,N_5725,N_5846);
nor U12782 (N_12782,N_7486,N_8862);
or U12783 (N_12783,N_8819,N_8030);
and U12784 (N_12784,N_8377,N_9014);
nor U12785 (N_12785,N_7051,N_6210);
nand U12786 (N_12786,N_7035,N_7653);
or U12787 (N_12787,N_7734,N_9271);
and U12788 (N_12788,N_9069,N_6790);
and U12789 (N_12789,N_6451,N_5192);
nor U12790 (N_12790,N_6075,N_7689);
nor U12791 (N_12791,N_9911,N_7152);
or U12792 (N_12792,N_8053,N_9518);
nor U12793 (N_12793,N_9206,N_6149);
xnor U12794 (N_12794,N_8683,N_9402);
xnor U12795 (N_12795,N_6981,N_9712);
or U12796 (N_12796,N_9305,N_8344);
xor U12797 (N_12797,N_5425,N_7893);
nand U12798 (N_12798,N_5105,N_8307);
nor U12799 (N_12799,N_7152,N_5032);
and U12800 (N_12800,N_6639,N_8402);
or U12801 (N_12801,N_9840,N_6663);
nand U12802 (N_12802,N_5005,N_6027);
nand U12803 (N_12803,N_9842,N_7545);
and U12804 (N_12804,N_8670,N_5772);
and U12805 (N_12805,N_7356,N_6677);
and U12806 (N_12806,N_7984,N_5700);
xor U12807 (N_12807,N_7759,N_9785);
or U12808 (N_12808,N_5776,N_5227);
nor U12809 (N_12809,N_9037,N_8015);
or U12810 (N_12810,N_7787,N_7623);
nor U12811 (N_12811,N_7700,N_6208);
nand U12812 (N_12812,N_8816,N_6727);
xnor U12813 (N_12813,N_6680,N_5641);
or U12814 (N_12814,N_5084,N_6670);
and U12815 (N_12815,N_9309,N_6175);
nor U12816 (N_12816,N_5068,N_8026);
and U12817 (N_12817,N_7384,N_6558);
and U12818 (N_12818,N_7511,N_5314);
xor U12819 (N_12819,N_6123,N_5330);
nand U12820 (N_12820,N_6353,N_7247);
nand U12821 (N_12821,N_6803,N_7789);
and U12822 (N_12822,N_9496,N_8578);
or U12823 (N_12823,N_5314,N_6131);
nor U12824 (N_12824,N_7258,N_6664);
nor U12825 (N_12825,N_8282,N_7002);
nand U12826 (N_12826,N_7106,N_6860);
and U12827 (N_12827,N_7230,N_7667);
xnor U12828 (N_12828,N_9220,N_9183);
nand U12829 (N_12829,N_5834,N_5871);
and U12830 (N_12830,N_5044,N_5876);
xnor U12831 (N_12831,N_9450,N_7175);
nand U12832 (N_12832,N_6905,N_6162);
nor U12833 (N_12833,N_6815,N_5707);
nor U12834 (N_12834,N_8006,N_7340);
xnor U12835 (N_12835,N_9887,N_6552);
nor U12836 (N_12836,N_5350,N_8298);
xor U12837 (N_12837,N_8109,N_9730);
and U12838 (N_12838,N_5168,N_8605);
nand U12839 (N_12839,N_8352,N_9550);
xor U12840 (N_12840,N_5816,N_6664);
xor U12841 (N_12841,N_5206,N_7212);
xor U12842 (N_12842,N_7920,N_6003);
or U12843 (N_12843,N_5082,N_5458);
and U12844 (N_12844,N_6940,N_7930);
or U12845 (N_12845,N_8849,N_7175);
nor U12846 (N_12846,N_9424,N_6577);
nor U12847 (N_12847,N_8481,N_7892);
xnor U12848 (N_12848,N_6618,N_8803);
nor U12849 (N_12849,N_8077,N_8607);
nor U12850 (N_12850,N_5228,N_5965);
xnor U12851 (N_12851,N_8056,N_8335);
nor U12852 (N_12852,N_7394,N_8823);
xor U12853 (N_12853,N_6015,N_6182);
nand U12854 (N_12854,N_9231,N_9049);
and U12855 (N_12855,N_8023,N_9801);
and U12856 (N_12856,N_8717,N_8926);
nand U12857 (N_12857,N_5326,N_9360);
or U12858 (N_12858,N_8125,N_6274);
nand U12859 (N_12859,N_7952,N_9471);
and U12860 (N_12860,N_5853,N_5662);
nand U12861 (N_12861,N_7232,N_8075);
xnor U12862 (N_12862,N_9723,N_7741);
or U12863 (N_12863,N_5132,N_6008);
or U12864 (N_12864,N_5354,N_8705);
nand U12865 (N_12865,N_6035,N_8889);
or U12866 (N_12866,N_7021,N_7426);
nand U12867 (N_12867,N_5791,N_8142);
nor U12868 (N_12868,N_5110,N_6340);
and U12869 (N_12869,N_9111,N_6718);
nor U12870 (N_12870,N_7151,N_9887);
xor U12871 (N_12871,N_6301,N_9615);
nor U12872 (N_12872,N_8968,N_7584);
or U12873 (N_12873,N_8387,N_5784);
xnor U12874 (N_12874,N_6970,N_9749);
and U12875 (N_12875,N_8764,N_8196);
nand U12876 (N_12876,N_8211,N_9551);
or U12877 (N_12877,N_5914,N_6225);
nor U12878 (N_12878,N_5939,N_5106);
and U12879 (N_12879,N_5239,N_9007);
nand U12880 (N_12880,N_5279,N_5177);
nor U12881 (N_12881,N_6612,N_6566);
and U12882 (N_12882,N_7502,N_9225);
nand U12883 (N_12883,N_8738,N_6756);
and U12884 (N_12884,N_5684,N_9740);
and U12885 (N_12885,N_7717,N_5902);
nor U12886 (N_12886,N_9909,N_6125);
nor U12887 (N_12887,N_9974,N_6327);
and U12888 (N_12888,N_5508,N_6369);
and U12889 (N_12889,N_6786,N_8129);
xor U12890 (N_12890,N_9627,N_8439);
nand U12891 (N_12891,N_6002,N_5635);
xor U12892 (N_12892,N_6647,N_8797);
nor U12893 (N_12893,N_9696,N_6360);
xnor U12894 (N_12894,N_9191,N_6130);
and U12895 (N_12895,N_6193,N_5729);
xnor U12896 (N_12896,N_8474,N_7343);
or U12897 (N_12897,N_6458,N_8968);
and U12898 (N_12898,N_7405,N_6888);
nand U12899 (N_12899,N_8971,N_9610);
nand U12900 (N_12900,N_8708,N_6635);
xnor U12901 (N_12901,N_6634,N_7098);
and U12902 (N_12902,N_8765,N_5451);
nand U12903 (N_12903,N_8521,N_6324);
nand U12904 (N_12904,N_5492,N_7265);
nor U12905 (N_12905,N_9094,N_7897);
or U12906 (N_12906,N_7244,N_6331);
and U12907 (N_12907,N_9774,N_5429);
and U12908 (N_12908,N_6007,N_7997);
or U12909 (N_12909,N_6810,N_5971);
nor U12910 (N_12910,N_9610,N_6309);
and U12911 (N_12911,N_7840,N_8672);
and U12912 (N_12912,N_9736,N_6410);
and U12913 (N_12913,N_7946,N_9194);
or U12914 (N_12914,N_7835,N_5001);
and U12915 (N_12915,N_6593,N_6942);
nand U12916 (N_12916,N_5795,N_9014);
nor U12917 (N_12917,N_5002,N_9337);
nor U12918 (N_12918,N_5942,N_7301);
xor U12919 (N_12919,N_6316,N_6102);
nor U12920 (N_12920,N_5947,N_5453);
nor U12921 (N_12921,N_7028,N_9946);
and U12922 (N_12922,N_9752,N_7950);
and U12923 (N_12923,N_6338,N_8306);
or U12924 (N_12924,N_7799,N_8417);
nand U12925 (N_12925,N_6708,N_6642);
nor U12926 (N_12926,N_6649,N_6466);
nand U12927 (N_12927,N_6731,N_7814);
and U12928 (N_12928,N_9195,N_6741);
nand U12929 (N_12929,N_6969,N_7204);
and U12930 (N_12930,N_7216,N_8731);
nand U12931 (N_12931,N_7781,N_8557);
nor U12932 (N_12932,N_5983,N_9936);
and U12933 (N_12933,N_9882,N_5586);
or U12934 (N_12934,N_6033,N_6734);
xnor U12935 (N_12935,N_7174,N_7123);
nand U12936 (N_12936,N_7118,N_8961);
nor U12937 (N_12937,N_6889,N_9479);
nor U12938 (N_12938,N_5466,N_7359);
or U12939 (N_12939,N_9948,N_8127);
or U12940 (N_12940,N_8602,N_9358);
and U12941 (N_12941,N_7416,N_7646);
nor U12942 (N_12942,N_6103,N_7131);
nand U12943 (N_12943,N_7846,N_6333);
nand U12944 (N_12944,N_7987,N_9976);
nand U12945 (N_12945,N_8889,N_8114);
nand U12946 (N_12946,N_8545,N_8491);
and U12947 (N_12947,N_5117,N_8132);
nand U12948 (N_12948,N_6723,N_6862);
or U12949 (N_12949,N_5967,N_7321);
nand U12950 (N_12950,N_9570,N_6550);
or U12951 (N_12951,N_5418,N_5604);
nor U12952 (N_12952,N_6056,N_8611);
xnor U12953 (N_12953,N_7648,N_8174);
or U12954 (N_12954,N_8664,N_8155);
or U12955 (N_12955,N_6930,N_6315);
xnor U12956 (N_12956,N_8941,N_6650);
xnor U12957 (N_12957,N_7430,N_8525);
and U12958 (N_12958,N_7548,N_6666);
or U12959 (N_12959,N_7505,N_5505);
nand U12960 (N_12960,N_5692,N_9529);
nor U12961 (N_12961,N_9965,N_6812);
or U12962 (N_12962,N_7534,N_9292);
and U12963 (N_12963,N_8264,N_5129);
and U12964 (N_12964,N_6002,N_6950);
xor U12965 (N_12965,N_6296,N_9551);
and U12966 (N_12966,N_5306,N_9815);
nor U12967 (N_12967,N_7773,N_8110);
and U12968 (N_12968,N_8011,N_7257);
nor U12969 (N_12969,N_6551,N_7701);
nand U12970 (N_12970,N_5607,N_8554);
or U12971 (N_12971,N_5776,N_6751);
nor U12972 (N_12972,N_9572,N_7144);
nand U12973 (N_12973,N_8647,N_7309);
and U12974 (N_12974,N_7616,N_7003);
xor U12975 (N_12975,N_6428,N_5209);
xor U12976 (N_12976,N_7296,N_9961);
nor U12977 (N_12977,N_6708,N_7765);
nand U12978 (N_12978,N_9595,N_5326);
and U12979 (N_12979,N_8648,N_9073);
nand U12980 (N_12980,N_8824,N_7266);
and U12981 (N_12981,N_9765,N_5587);
nand U12982 (N_12982,N_7339,N_8781);
or U12983 (N_12983,N_6144,N_6047);
nor U12984 (N_12984,N_6079,N_5930);
xnor U12985 (N_12985,N_5696,N_9144);
nand U12986 (N_12986,N_9023,N_7663);
or U12987 (N_12987,N_9546,N_8261);
xor U12988 (N_12988,N_6595,N_9372);
nor U12989 (N_12989,N_7444,N_6498);
and U12990 (N_12990,N_7385,N_9097);
or U12991 (N_12991,N_8427,N_8480);
nand U12992 (N_12992,N_6884,N_7879);
xor U12993 (N_12993,N_5245,N_9976);
or U12994 (N_12994,N_5067,N_8684);
xor U12995 (N_12995,N_9168,N_6261);
or U12996 (N_12996,N_9009,N_7462);
or U12997 (N_12997,N_9916,N_9992);
xnor U12998 (N_12998,N_8419,N_7242);
nor U12999 (N_12999,N_6023,N_7187);
or U13000 (N_13000,N_9047,N_8799);
xor U13001 (N_13001,N_5021,N_9274);
xor U13002 (N_13002,N_9391,N_6932);
xnor U13003 (N_13003,N_5930,N_9453);
nor U13004 (N_13004,N_6818,N_6699);
or U13005 (N_13005,N_9531,N_6176);
and U13006 (N_13006,N_9425,N_5275);
xor U13007 (N_13007,N_9042,N_8133);
nand U13008 (N_13008,N_9790,N_5505);
and U13009 (N_13009,N_7042,N_7096);
xnor U13010 (N_13010,N_9555,N_6332);
and U13011 (N_13011,N_6787,N_8290);
and U13012 (N_13012,N_5253,N_7900);
xnor U13013 (N_13013,N_9105,N_9563);
xnor U13014 (N_13014,N_8341,N_9493);
and U13015 (N_13015,N_7135,N_5161);
or U13016 (N_13016,N_5195,N_9677);
nor U13017 (N_13017,N_6705,N_8379);
nand U13018 (N_13018,N_9430,N_6675);
nand U13019 (N_13019,N_6949,N_8161);
nor U13020 (N_13020,N_9607,N_6248);
nor U13021 (N_13021,N_6548,N_7310);
xnor U13022 (N_13022,N_8198,N_6464);
and U13023 (N_13023,N_7534,N_7792);
or U13024 (N_13024,N_6019,N_8182);
xnor U13025 (N_13025,N_6043,N_8466);
nor U13026 (N_13026,N_5970,N_5417);
or U13027 (N_13027,N_7101,N_5591);
nor U13028 (N_13028,N_5148,N_5578);
or U13029 (N_13029,N_5236,N_8763);
nand U13030 (N_13030,N_9938,N_6574);
nor U13031 (N_13031,N_8502,N_8775);
xnor U13032 (N_13032,N_7559,N_6124);
or U13033 (N_13033,N_5315,N_8627);
and U13034 (N_13034,N_9197,N_7205);
xnor U13035 (N_13035,N_5896,N_7390);
or U13036 (N_13036,N_5473,N_7178);
or U13037 (N_13037,N_8854,N_5532);
and U13038 (N_13038,N_5368,N_8696);
or U13039 (N_13039,N_8027,N_6819);
xnor U13040 (N_13040,N_5086,N_5316);
nand U13041 (N_13041,N_6343,N_6148);
or U13042 (N_13042,N_7751,N_8699);
nor U13043 (N_13043,N_8263,N_5690);
nor U13044 (N_13044,N_5787,N_9113);
nor U13045 (N_13045,N_8071,N_9712);
and U13046 (N_13046,N_5588,N_8133);
nor U13047 (N_13047,N_6482,N_6274);
nor U13048 (N_13048,N_7030,N_5103);
or U13049 (N_13049,N_5347,N_6911);
nor U13050 (N_13050,N_5786,N_9191);
nor U13051 (N_13051,N_5996,N_8607);
or U13052 (N_13052,N_9958,N_8325);
xnor U13053 (N_13053,N_7334,N_9622);
and U13054 (N_13054,N_9185,N_6322);
nor U13055 (N_13055,N_9455,N_8723);
nand U13056 (N_13056,N_5410,N_5379);
and U13057 (N_13057,N_7658,N_5364);
nand U13058 (N_13058,N_6874,N_5689);
xnor U13059 (N_13059,N_5342,N_9239);
and U13060 (N_13060,N_7394,N_8073);
nor U13061 (N_13061,N_8381,N_6983);
or U13062 (N_13062,N_8809,N_5027);
and U13063 (N_13063,N_6351,N_5749);
and U13064 (N_13064,N_5114,N_6340);
nand U13065 (N_13065,N_5676,N_9306);
or U13066 (N_13066,N_7522,N_9554);
xnor U13067 (N_13067,N_9043,N_9623);
nor U13068 (N_13068,N_5094,N_8503);
and U13069 (N_13069,N_7192,N_8547);
nor U13070 (N_13070,N_9524,N_5427);
xor U13071 (N_13071,N_9969,N_7004);
xnor U13072 (N_13072,N_7752,N_6754);
and U13073 (N_13073,N_6837,N_6555);
xnor U13074 (N_13074,N_9263,N_8952);
xnor U13075 (N_13075,N_9085,N_9477);
or U13076 (N_13076,N_6469,N_7629);
or U13077 (N_13077,N_8970,N_9300);
and U13078 (N_13078,N_6963,N_5851);
nor U13079 (N_13079,N_9264,N_7423);
and U13080 (N_13080,N_8114,N_8475);
xnor U13081 (N_13081,N_8167,N_7818);
or U13082 (N_13082,N_9117,N_5746);
xnor U13083 (N_13083,N_5077,N_5138);
xor U13084 (N_13084,N_5130,N_8174);
or U13085 (N_13085,N_8716,N_5841);
nor U13086 (N_13086,N_9239,N_9886);
nand U13087 (N_13087,N_6320,N_8903);
nand U13088 (N_13088,N_7407,N_5656);
nor U13089 (N_13089,N_8806,N_5878);
nand U13090 (N_13090,N_7682,N_6699);
nand U13091 (N_13091,N_7706,N_5490);
or U13092 (N_13092,N_8324,N_7898);
nand U13093 (N_13093,N_9848,N_5204);
or U13094 (N_13094,N_9620,N_8152);
nand U13095 (N_13095,N_5288,N_5649);
or U13096 (N_13096,N_7997,N_9501);
nor U13097 (N_13097,N_6458,N_6322);
nor U13098 (N_13098,N_6472,N_8407);
nand U13099 (N_13099,N_5125,N_7556);
xnor U13100 (N_13100,N_9505,N_8145);
nand U13101 (N_13101,N_7594,N_9910);
nand U13102 (N_13102,N_6899,N_7637);
nor U13103 (N_13103,N_9053,N_6470);
xnor U13104 (N_13104,N_5835,N_8663);
xor U13105 (N_13105,N_6934,N_6614);
or U13106 (N_13106,N_6617,N_5851);
nand U13107 (N_13107,N_5867,N_8416);
xor U13108 (N_13108,N_8493,N_6984);
and U13109 (N_13109,N_7511,N_8431);
xnor U13110 (N_13110,N_8513,N_7909);
xor U13111 (N_13111,N_6164,N_8247);
and U13112 (N_13112,N_7791,N_7214);
or U13113 (N_13113,N_9185,N_5866);
or U13114 (N_13114,N_9154,N_9227);
or U13115 (N_13115,N_6021,N_7818);
and U13116 (N_13116,N_6081,N_8611);
xor U13117 (N_13117,N_6655,N_5037);
nor U13118 (N_13118,N_5651,N_8212);
nand U13119 (N_13119,N_8984,N_6409);
and U13120 (N_13120,N_8155,N_9008);
nor U13121 (N_13121,N_7185,N_9216);
nor U13122 (N_13122,N_6934,N_8992);
nor U13123 (N_13123,N_8064,N_6520);
nand U13124 (N_13124,N_7631,N_9901);
nand U13125 (N_13125,N_8298,N_8257);
and U13126 (N_13126,N_6883,N_8834);
xor U13127 (N_13127,N_7177,N_9328);
nand U13128 (N_13128,N_5483,N_9305);
xnor U13129 (N_13129,N_6280,N_9377);
or U13130 (N_13130,N_7773,N_9998);
nand U13131 (N_13131,N_9779,N_9846);
or U13132 (N_13132,N_6908,N_5102);
or U13133 (N_13133,N_6646,N_8299);
nand U13134 (N_13134,N_9993,N_6967);
xor U13135 (N_13135,N_7023,N_8024);
nor U13136 (N_13136,N_6391,N_6893);
and U13137 (N_13137,N_9847,N_5744);
nand U13138 (N_13138,N_9399,N_5877);
xor U13139 (N_13139,N_5781,N_9084);
nand U13140 (N_13140,N_8011,N_5274);
or U13141 (N_13141,N_7273,N_8710);
nor U13142 (N_13142,N_5230,N_7220);
and U13143 (N_13143,N_7778,N_9754);
nand U13144 (N_13144,N_9746,N_6898);
nor U13145 (N_13145,N_5596,N_5821);
and U13146 (N_13146,N_5887,N_8193);
xor U13147 (N_13147,N_8075,N_8149);
and U13148 (N_13148,N_9356,N_7161);
nand U13149 (N_13149,N_8534,N_7201);
nand U13150 (N_13150,N_7765,N_5469);
or U13151 (N_13151,N_5779,N_7360);
xnor U13152 (N_13152,N_8550,N_7467);
or U13153 (N_13153,N_6408,N_8762);
nand U13154 (N_13154,N_8080,N_8727);
nor U13155 (N_13155,N_9789,N_7472);
and U13156 (N_13156,N_8965,N_8718);
nor U13157 (N_13157,N_7762,N_9326);
xor U13158 (N_13158,N_7489,N_8363);
xor U13159 (N_13159,N_9092,N_9624);
nor U13160 (N_13160,N_5650,N_7191);
nand U13161 (N_13161,N_9265,N_5970);
or U13162 (N_13162,N_9634,N_9924);
nand U13163 (N_13163,N_6369,N_9123);
nand U13164 (N_13164,N_5919,N_7134);
nor U13165 (N_13165,N_6630,N_7331);
and U13166 (N_13166,N_9438,N_6912);
nor U13167 (N_13167,N_6870,N_6937);
or U13168 (N_13168,N_6994,N_7581);
nand U13169 (N_13169,N_9379,N_9524);
xor U13170 (N_13170,N_8318,N_8455);
nor U13171 (N_13171,N_5879,N_7858);
nor U13172 (N_13172,N_5598,N_8193);
and U13173 (N_13173,N_7829,N_6246);
nor U13174 (N_13174,N_5968,N_9214);
nor U13175 (N_13175,N_6127,N_6240);
or U13176 (N_13176,N_9083,N_8072);
nor U13177 (N_13177,N_6752,N_7197);
nand U13178 (N_13178,N_9363,N_7894);
nand U13179 (N_13179,N_8384,N_8070);
xor U13180 (N_13180,N_6239,N_9757);
xnor U13181 (N_13181,N_8816,N_6361);
nor U13182 (N_13182,N_7071,N_8623);
and U13183 (N_13183,N_8507,N_5650);
nand U13184 (N_13184,N_5480,N_5671);
or U13185 (N_13185,N_5267,N_9041);
nor U13186 (N_13186,N_7431,N_6517);
xnor U13187 (N_13187,N_7024,N_5824);
xnor U13188 (N_13188,N_9137,N_8548);
and U13189 (N_13189,N_6359,N_5092);
xor U13190 (N_13190,N_6805,N_6170);
or U13191 (N_13191,N_6382,N_9005);
or U13192 (N_13192,N_8097,N_9562);
nor U13193 (N_13193,N_5268,N_9245);
or U13194 (N_13194,N_9988,N_8645);
nor U13195 (N_13195,N_8849,N_9380);
nor U13196 (N_13196,N_9283,N_8664);
nor U13197 (N_13197,N_7992,N_9869);
xor U13198 (N_13198,N_7095,N_8065);
and U13199 (N_13199,N_9557,N_9411);
and U13200 (N_13200,N_7227,N_9250);
and U13201 (N_13201,N_5318,N_7327);
and U13202 (N_13202,N_8400,N_8438);
and U13203 (N_13203,N_6274,N_6053);
xor U13204 (N_13204,N_8813,N_9483);
nor U13205 (N_13205,N_7177,N_5434);
nand U13206 (N_13206,N_8381,N_6591);
and U13207 (N_13207,N_7486,N_6830);
and U13208 (N_13208,N_7270,N_8318);
nor U13209 (N_13209,N_6627,N_5310);
nor U13210 (N_13210,N_5512,N_9292);
xnor U13211 (N_13211,N_8080,N_8292);
nor U13212 (N_13212,N_6884,N_5613);
nand U13213 (N_13213,N_6528,N_9925);
nand U13214 (N_13214,N_6460,N_5507);
or U13215 (N_13215,N_6393,N_7668);
xnor U13216 (N_13216,N_8414,N_9388);
and U13217 (N_13217,N_7292,N_6480);
or U13218 (N_13218,N_7290,N_7999);
and U13219 (N_13219,N_9146,N_9565);
or U13220 (N_13220,N_7765,N_5099);
and U13221 (N_13221,N_6742,N_7183);
and U13222 (N_13222,N_5586,N_8985);
and U13223 (N_13223,N_8705,N_8551);
xor U13224 (N_13224,N_9403,N_7120);
xor U13225 (N_13225,N_5914,N_6256);
xor U13226 (N_13226,N_6231,N_8664);
or U13227 (N_13227,N_5416,N_5534);
or U13228 (N_13228,N_5566,N_6529);
xnor U13229 (N_13229,N_8654,N_5981);
and U13230 (N_13230,N_7809,N_8242);
nor U13231 (N_13231,N_5806,N_7605);
or U13232 (N_13232,N_8185,N_8776);
and U13233 (N_13233,N_7258,N_7931);
nor U13234 (N_13234,N_9008,N_9846);
nor U13235 (N_13235,N_6141,N_5505);
xnor U13236 (N_13236,N_9603,N_5493);
nand U13237 (N_13237,N_7380,N_7082);
and U13238 (N_13238,N_9485,N_6519);
xnor U13239 (N_13239,N_8532,N_8326);
nor U13240 (N_13240,N_5900,N_9376);
nand U13241 (N_13241,N_9321,N_7522);
and U13242 (N_13242,N_9850,N_6047);
or U13243 (N_13243,N_7544,N_6199);
xor U13244 (N_13244,N_8241,N_5982);
xor U13245 (N_13245,N_8958,N_8054);
or U13246 (N_13246,N_9117,N_7960);
or U13247 (N_13247,N_6264,N_5314);
xor U13248 (N_13248,N_6782,N_9938);
and U13249 (N_13249,N_8844,N_6614);
nor U13250 (N_13250,N_6503,N_7277);
xor U13251 (N_13251,N_5237,N_5807);
nor U13252 (N_13252,N_9683,N_5270);
and U13253 (N_13253,N_9826,N_8371);
nor U13254 (N_13254,N_7172,N_8297);
or U13255 (N_13255,N_9466,N_6086);
or U13256 (N_13256,N_7404,N_8213);
xor U13257 (N_13257,N_6434,N_7939);
xnor U13258 (N_13258,N_9001,N_7318);
and U13259 (N_13259,N_6647,N_8611);
or U13260 (N_13260,N_6538,N_6848);
or U13261 (N_13261,N_7480,N_6930);
and U13262 (N_13262,N_5566,N_8118);
nor U13263 (N_13263,N_8258,N_8519);
or U13264 (N_13264,N_5900,N_6833);
nor U13265 (N_13265,N_5513,N_5499);
nor U13266 (N_13266,N_8517,N_7795);
or U13267 (N_13267,N_5538,N_5221);
and U13268 (N_13268,N_7866,N_5103);
and U13269 (N_13269,N_6824,N_8328);
nand U13270 (N_13270,N_9042,N_6400);
nand U13271 (N_13271,N_9779,N_8249);
or U13272 (N_13272,N_6819,N_8017);
and U13273 (N_13273,N_5190,N_7429);
or U13274 (N_13274,N_5090,N_9022);
or U13275 (N_13275,N_8436,N_5743);
and U13276 (N_13276,N_8248,N_9253);
nand U13277 (N_13277,N_5410,N_6386);
and U13278 (N_13278,N_9795,N_8650);
xor U13279 (N_13279,N_8704,N_5171);
and U13280 (N_13280,N_7867,N_6771);
nand U13281 (N_13281,N_7806,N_7936);
and U13282 (N_13282,N_9299,N_9762);
nand U13283 (N_13283,N_6424,N_7445);
nand U13284 (N_13284,N_8148,N_5361);
and U13285 (N_13285,N_9138,N_8091);
nand U13286 (N_13286,N_7065,N_7634);
or U13287 (N_13287,N_7001,N_8124);
nor U13288 (N_13288,N_5039,N_5678);
nor U13289 (N_13289,N_8785,N_6212);
and U13290 (N_13290,N_5982,N_7102);
or U13291 (N_13291,N_5466,N_9285);
nand U13292 (N_13292,N_6060,N_6750);
nor U13293 (N_13293,N_7119,N_6349);
xor U13294 (N_13294,N_8900,N_5041);
nor U13295 (N_13295,N_6212,N_5723);
and U13296 (N_13296,N_8206,N_9754);
or U13297 (N_13297,N_7007,N_7145);
nor U13298 (N_13298,N_9615,N_6118);
nor U13299 (N_13299,N_9659,N_7882);
xor U13300 (N_13300,N_9242,N_5925);
and U13301 (N_13301,N_5829,N_9562);
xor U13302 (N_13302,N_5372,N_9375);
nand U13303 (N_13303,N_6629,N_7677);
xor U13304 (N_13304,N_6898,N_6112);
and U13305 (N_13305,N_9609,N_6798);
nor U13306 (N_13306,N_7354,N_5548);
nand U13307 (N_13307,N_6242,N_5499);
nand U13308 (N_13308,N_7060,N_6338);
nor U13309 (N_13309,N_8561,N_8321);
nand U13310 (N_13310,N_6325,N_5283);
or U13311 (N_13311,N_9867,N_6450);
and U13312 (N_13312,N_7682,N_5141);
nand U13313 (N_13313,N_6282,N_9108);
xor U13314 (N_13314,N_6732,N_8808);
or U13315 (N_13315,N_8713,N_7929);
and U13316 (N_13316,N_9726,N_5519);
or U13317 (N_13317,N_5089,N_7627);
nor U13318 (N_13318,N_9526,N_6478);
or U13319 (N_13319,N_6155,N_9177);
nor U13320 (N_13320,N_5753,N_6134);
and U13321 (N_13321,N_7275,N_5779);
nor U13322 (N_13322,N_9629,N_9198);
or U13323 (N_13323,N_9773,N_5504);
or U13324 (N_13324,N_8778,N_9293);
or U13325 (N_13325,N_9445,N_6390);
and U13326 (N_13326,N_9272,N_6997);
xnor U13327 (N_13327,N_9615,N_7485);
or U13328 (N_13328,N_6876,N_8696);
xnor U13329 (N_13329,N_6377,N_7985);
or U13330 (N_13330,N_7470,N_6975);
or U13331 (N_13331,N_6452,N_7370);
or U13332 (N_13332,N_7966,N_5425);
nand U13333 (N_13333,N_8827,N_7821);
nand U13334 (N_13334,N_7916,N_9424);
nand U13335 (N_13335,N_9199,N_8023);
nor U13336 (N_13336,N_8940,N_5904);
xnor U13337 (N_13337,N_6241,N_8051);
nor U13338 (N_13338,N_9285,N_5258);
or U13339 (N_13339,N_6201,N_8120);
xnor U13340 (N_13340,N_9690,N_8340);
nand U13341 (N_13341,N_9404,N_7331);
and U13342 (N_13342,N_5700,N_6298);
or U13343 (N_13343,N_8815,N_7476);
or U13344 (N_13344,N_7552,N_6315);
xnor U13345 (N_13345,N_5729,N_8120);
xnor U13346 (N_13346,N_5032,N_9062);
nand U13347 (N_13347,N_6907,N_7588);
or U13348 (N_13348,N_9106,N_7487);
nor U13349 (N_13349,N_5037,N_9743);
nor U13350 (N_13350,N_5727,N_5725);
or U13351 (N_13351,N_9971,N_7809);
and U13352 (N_13352,N_5169,N_7823);
and U13353 (N_13353,N_8035,N_6546);
nand U13354 (N_13354,N_7062,N_9437);
xnor U13355 (N_13355,N_6349,N_8800);
or U13356 (N_13356,N_8260,N_6336);
nor U13357 (N_13357,N_8717,N_8965);
xor U13358 (N_13358,N_6568,N_9686);
xnor U13359 (N_13359,N_5477,N_6537);
nand U13360 (N_13360,N_7323,N_6398);
nor U13361 (N_13361,N_8469,N_7544);
xor U13362 (N_13362,N_8891,N_5280);
nor U13363 (N_13363,N_8354,N_9231);
and U13364 (N_13364,N_8495,N_9468);
nand U13365 (N_13365,N_5569,N_8008);
xor U13366 (N_13366,N_9032,N_9332);
and U13367 (N_13367,N_6352,N_6783);
nor U13368 (N_13368,N_5398,N_7580);
nor U13369 (N_13369,N_9016,N_5108);
and U13370 (N_13370,N_9169,N_5164);
or U13371 (N_13371,N_8807,N_5483);
and U13372 (N_13372,N_6310,N_6904);
xor U13373 (N_13373,N_9335,N_8862);
nand U13374 (N_13374,N_9026,N_7862);
or U13375 (N_13375,N_6970,N_5915);
xor U13376 (N_13376,N_8149,N_6479);
or U13377 (N_13377,N_5183,N_8179);
and U13378 (N_13378,N_7836,N_7178);
xnor U13379 (N_13379,N_8477,N_8684);
and U13380 (N_13380,N_7539,N_5906);
and U13381 (N_13381,N_9162,N_9137);
xor U13382 (N_13382,N_8513,N_5359);
or U13383 (N_13383,N_6515,N_9270);
xor U13384 (N_13384,N_8242,N_9612);
nor U13385 (N_13385,N_8631,N_7291);
and U13386 (N_13386,N_7580,N_5756);
or U13387 (N_13387,N_7740,N_7204);
nor U13388 (N_13388,N_9600,N_8759);
and U13389 (N_13389,N_5863,N_6348);
nand U13390 (N_13390,N_5000,N_6080);
nor U13391 (N_13391,N_7799,N_5256);
nor U13392 (N_13392,N_9822,N_6229);
and U13393 (N_13393,N_5596,N_8503);
or U13394 (N_13394,N_7883,N_7073);
or U13395 (N_13395,N_5881,N_9686);
xnor U13396 (N_13396,N_8176,N_8648);
nor U13397 (N_13397,N_7793,N_8541);
xor U13398 (N_13398,N_7405,N_9206);
or U13399 (N_13399,N_8221,N_8216);
or U13400 (N_13400,N_9393,N_5835);
nand U13401 (N_13401,N_9146,N_5340);
nand U13402 (N_13402,N_8221,N_5908);
nor U13403 (N_13403,N_7992,N_8220);
or U13404 (N_13404,N_5837,N_5159);
or U13405 (N_13405,N_9253,N_9137);
and U13406 (N_13406,N_8113,N_5858);
nor U13407 (N_13407,N_9456,N_9803);
or U13408 (N_13408,N_8019,N_7793);
and U13409 (N_13409,N_9554,N_8919);
or U13410 (N_13410,N_5920,N_5307);
nand U13411 (N_13411,N_6026,N_9785);
and U13412 (N_13412,N_8659,N_9485);
and U13413 (N_13413,N_9157,N_7779);
xnor U13414 (N_13414,N_7356,N_7079);
nand U13415 (N_13415,N_8924,N_8686);
xor U13416 (N_13416,N_8321,N_6731);
xor U13417 (N_13417,N_6068,N_5365);
or U13418 (N_13418,N_5193,N_9175);
nand U13419 (N_13419,N_7114,N_5061);
and U13420 (N_13420,N_6256,N_9802);
or U13421 (N_13421,N_7171,N_5043);
nor U13422 (N_13422,N_7276,N_6208);
nor U13423 (N_13423,N_6547,N_7136);
or U13424 (N_13424,N_8915,N_5713);
nand U13425 (N_13425,N_8803,N_6880);
nor U13426 (N_13426,N_7321,N_9295);
and U13427 (N_13427,N_9023,N_7827);
or U13428 (N_13428,N_9922,N_5271);
nand U13429 (N_13429,N_5701,N_5632);
or U13430 (N_13430,N_7141,N_8408);
nor U13431 (N_13431,N_7231,N_7508);
nor U13432 (N_13432,N_7175,N_7193);
xnor U13433 (N_13433,N_6631,N_7994);
nor U13434 (N_13434,N_7431,N_9541);
xor U13435 (N_13435,N_8951,N_6414);
xor U13436 (N_13436,N_7220,N_7912);
nor U13437 (N_13437,N_6184,N_6653);
nand U13438 (N_13438,N_6559,N_9870);
nor U13439 (N_13439,N_6544,N_9345);
nor U13440 (N_13440,N_9736,N_8780);
or U13441 (N_13441,N_5207,N_9031);
xnor U13442 (N_13442,N_5765,N_6829);
nor U13443 (N_13443,N_7570,N_9264);
xnor U13444 (N_13444,N_6682,N_7461);
nor U13445 (N_13445,N_6183,N_9620);
xor U13446 (N_13446,N_5942,N_5819);
nand U13447 (N_13447,N_7375,N_7533);
xor U13448 (N_13448,N_8642,N_7552);
and U13449 (N_13449,N_8143,N_8623);
nor U13450 (N_13450,N_5010,N_6167);
or U13451 (N_13451,N_5640,N_5385);
nor U13452 (N_13452,N_8943,N_5410);
or U13453 (N_13453,N_9269,N_7138);
xnor U13454 (N_13454,N_8831,N_7099);
or U13455 (N_13455,N_5682,N_9750);
or U13456 (N_13456,N_6873,N_9159);
xor U13457 (N_13457,N_7131,N_9089);
and U13458 (N_13458,N_7663,N_9660);
or U13459 (N_13459,N_6549,N_8467);
xor U13460 (N_13460,N_5722,N_7034);
xnor U13461 (N_13461,N_5527,N_8567);
xor U13462 (N_13462,N_5259,N_5511);
or U13463 (N_13463,N_8784,N_7674);
nor U13464 (N_13464,N_5074,N_8820);
and U13465 (N_13465,N_5389,N_7991);
nand U13466 (N_13466,N_6130,N_6579);
or U13467 (N_13467,N_9765,N_8234);
and U13468 (N_13468,N_6659,N_7178);
nor U13469 (N_13469,N_8461,N_8466);
nand U13470 (N_13470,N_6801,N_7859);
and U13471 (N_13471,N_5078,N_5651);
and U13472 (N_13472,N_9928,N_6110);
nand U13473 (N_13473,N_5564,N_6227);
and U13474 (N_13474,N_5407,N_9034);
nand U13475 (N_13475,N_8927,N_5753);
or U13476 (N_13476,N_5227,N_6179);
nand U13477 (N_13477,N_9722,N_7514);
nor U13478 (N_13478,N_5208,N_7708);
nor U13479 (N_13479,N_7269,N_7363);
nand U13480 (N_13480,N_7398,N_9952);
xnor U13481 (N_13481,N_7971,N_5569);
nor U13482 (N_13482,N_8801,N_8673);
or U13483 (N_13483,N_9062,N_7169);
and U13484 (N_13484,N_5572,N_9467);
xor U13485 (N_13485,N_6110,N_8981);
or U13486 (N_13486,N_5075,N_8449);
nor U13487 (N_13487,N_9960,N_5918);
nor U13488 (N_13488,N_7289,N_5374);
xor U13489 (N_13489,N_8240,N_6637);
xor U13490 (N_13490,N_9003,N_5260);
xor U13491 (N_13491,N_5673,N_6176);
and U13492 (N_13492,N_6523,N_9345);
nand U13493 (N_13493,N_5970,N_9914);
and U13494 (N_13494,N_8393,N_9397);
nor U13495 (N_13495,N_9849,N_6296);
nor U13496 (N_13496,N_8123,N_8717);
and U13497 (N_13497,N_9520,N_6431);
nand U13498 (N_13498,N_7737,N_6949);
or U13499 (N_13499,N_7871,N_7104);
and U13500 (N_13500,N_9254,N_8454);
nor U13501 (N_13501,N_9726,N_9704);
and U13502 (N_13502,N_9754,N_8201);
nor U13503 (N_13503,N_6356,N_8821);
nor U13504 (N_13504,N_6808,N_9994);
xnor U13505 (N_13505,N_6411,N_9290);
and U13506 (N_13506,N_7432,N_9721);
nor U13507 (N_13507,N_6725,N_8889);
nand U13508 (N_13508,N_9189,N_9876);
nor U13509 (N_13509,N_7246,N_8767);
or U13510 (N_13510,N_7867,N_8467);
and U13511 (N_13511,N_9480,N_9119);
nand U13512 (N_13512,N_7952,N_8035);
nor U13513 (N_13513,N_7885,N_6641);
or U13514 (N_13514,N_5989,N_8520);
or U13515 (N_13515,N_5394,N_7259);
and U13516 (N_13516,N_7624,N_8377);
nand U13517 (N_13517,N_7889,N_8009);
and U13518 (N_13518,N_7756,N_7699);
nand U13519 (N_13519,N_9361,N_8036);
nand U13520 (N_13520,N_5408,N_8404);
and U13521 (N_13521,N_5109,N_5708);
or U13522 (N_13522,N_8258,N_5989);
or U13523 (N_13523,N_5486,N_6063);
nand U13524 (N_13524,N_5376,N_9008);
nor U13525 (N_13525,N_5546,N_7004);
nand U13526 (N_13526,N_6653,N_8317);
or U13527 (N_13527,N_5804,N_6519);
xnor U13528 (N_13528,N_5947,N_7698);
or U13529 (N_13529,N_6691,N_8969);
and U13530 (N_13530,N_6916,N_8154);
xor U13531 (N_13531,N_5356,N_9048);
or U13532 (N_13532,N_7029,N_5542);
or U13533 (N_13533,N_8851,N_6860);
xnor U13534 (N_13534,N_6307,N_5981);
nand U13535 (N_13535,N_9257,N_6637);
or U13536 (N_13536,N_6886,N_5077);
nor U13537 (N_13537,N_9700,N_6325);
xor U13538 (N_13538,N_9487,N_8264);
and U13539 (N_13539,N_9679,N_5624);
or U13540 (N_13540,N_8733,N_8875);
nand U13541 (N_13541,N_8665,N_8227);
or U13542 (N_13542,N_5403,N_5472);
or U13543 (N_13543,N_7382,N_5937);
or U13544 (N_13544,N_5569,N_6657);
xnor U13545 (N_13545,N_6479,N_8722);
nor U13546 (N_13546,N_6339,N_9125);
nand U13547 (N_13547,N_8641,N_8151);
and U13548 (N_13548,N_8400,N_9351);
or U13549 (N_13549,N_7290,N_9137);
and U13550 (N_13550,N_6425,N_7900);
nand U13551 (N_13551,N_8347,N_6864);
and U13552 (N_13552,N_5699,N_9356);
and U13553 (N_13553,N_9020,N_6923);
nor U13554 (N_13554,N_6180,N_9667);
xnor U13555 (N_13555,N_6190,N_9169);
nand U13556 (N_13556,N_5384,N_9111);
nor U13557 (N_13557,N_7253,N_9138);
nand U13558 (N_13558,N_6925,N_8337);
nand U13559 (N_13559,N_7194,N_5134);
nor U13560 (N_13560,N_9534,N_5496);
or U13561 (N_13561,N_9043,N_5648);
nand U13562 (N_13562,N_8967,N_5495);
nor U13563 (N_13563,N_9101,N_6868);
xor U13564 (N_13564,N_7495,N_7344);
or U13565 (N_13565,N_9575,N_5141);
nor U13566 (N_13566,N_6192,N_5311);
xor U13567 (N_13567,N_6405,N_5845);
and U13568 (N_13568,N_5438,N_5947);
and U13569 (N_13569,N_9073,N_7382);
nand U13570 (N_13570,N_9717,N_9383);
nand U13571 (N_13571,N_7402,N_6793);
nor U13572 (N_13572,N_5202,N_9048);
xnor U13573 (N_13573,N_7053,N_6877);
and U13574 (N_13574,N_7887,N_9172);
xnor U13575 (N_13575,N_9086,N_7045);
xnor U13576 (N_13576,N_5562,N_5329);
nand U13577 (N_13577,N_7296,N_8707);
nand U13578 (N_13578,N_5869,N_8462);
nor U13579 (N_13579,N_5799,N_7410);
nor U13580 (N_13580,N_6730,N_9433);
nand U13581 (N_13581,N_9208,N_7427);
xnor U13582 (N_13582,N_8461,N_6622);
nor U13583 (N_13583,N_9828,N_5227);
nand U13584 (N_13584,N_6284,N_7064);
or U13585 (N_13585,N_6443,N_7411);
xnor U13586 (N_13586,N_8189,N_6986);
or U13587 (N_13587,N_5690,N_5057);
nor U13588 (N_13588,N_8780,N_7336);
xor U13589 (N_13589,N_5166,N_7330);
or U13590 (N_13590,N_9451,N_9400);
xor U13591 (N_13591,N_7660,N_5215);
xnor U13592 (N_13592,N_8989,N_7712);
and U13593 (N_13593,N_5506,N_6904);
nor U13594 (N_13594,N_5355,N_5382);
nor U13595 (N_13595,N_7266,N_5579);
and U13596 (N_13596,N_5841,N_6280);
nor U13597 (N_13597,N_9336,N_9250);
xor U13598 (N_13598,N_7279,N_9215);
nand U13599 (N_13599,N_5257,N_8663);
nand U13600 (N_13600,N_6020,N_6282);
xnor U13601 (N_13601,N_7590,N_9119);
xnor U13602 (N_13602,N_9418,N_7125);
or U13603 (N_13603,N_8820,N_8928);
and U13604 (N_13604,N_8629,N_9041);
nand U13605 (N_13605,N_7708,N_5967);
or U13606 (N_13606,N_5985,N_5950);
nor U13607 (N_13607,N_7300,N_5303);
and U13608 (N_13608,N_9354,N_9814);
nand U13609 (N_13609,N_8032,N_8710);
nand U13610 (N_13610,N_8498,N_9540);
nand U13611 (N_13611,N_9869,N_6853);
nor U13612 (N_13612,N_9171,N_6536);
and U13613 (N_13613,N_8565,N_8309);
xnor U13614 (N_13614,N_9792,N_6158);
or U13615 (N_13615,N_6309,N_8280);
and U13616 (N_13616,N_9219,N_9152);
and U13617 (N_13617,N_7585,N_6362);
nand U13618 (N_13618,N_7372,N_5564);
nor U13619 (N_13619,N_6581,N_7443);
or U13620 (N_13620,N_9898,N_9922);
or U13621 (N_13621,N_9924,N_7019);
nor U13622 (N_13622,N_6182,N_9743);
xor U13623 (N_13623,N_7058,N_7676);
or U13624 (N_13624,N_6410,N_6944);
nor U13625 (N_13625,N_9214,N_7523);
nor U13626 (N_13626,N_6891,N_9651);
nor U13627 (N_13627,N_9272,N_6220);
or U13628 (N_13628,N_9619,N_9439);
or U13629 (N_13629,N_7817,N_5468);
or U13630 (N_13630,N_9140,N_8659);
nand U13631 (N_13631,N_9594,N_9059);
xnor U13632 (N_13632,N_5739,N_5273);
xor U13633 (N_13633,N_5651,N_9712);
xnor U13634 (N_13634,N_6137,N_6262);
nor U13635 (N_13635,N_7540,N_6717);
xnor U13636 (N_13636,N_8121,N_5047);
and U13637 (N_13637,N_8719,N_5822);
and U13638 (N_13638,N_6558,N_9314);
and U13639 (N_13639,N_8185,N_5321);
and U13640 (N_13640,N_7577,N_8948);
or U13641 (N_13641,N_8457,N_8514);
or U13642 (N_13642,N_8867,N_6322);
xor U13643 (N_13643,N_9304,N_7841);
and U13644 (N_13644,N_5809,N_8913);
nand U13645 (N_13645,N_9378,N_8193);
nand U13646 (N_13646,N_8051,N_8020);
xnor U13647 (N_13647,N_9036,N_7217);
or U13648 (N_13648,N_7423,N_9189);
and U13649 (N_13649,N_5186,N_9597);
nand U13650 (N_13650,N_6514,N_5915);
or U13651 (N_13651,N_6297,N_9057);
xnor U13652 (N_13652,N_6484,N_5627);
or U13653 (N_13653,N_7122,N_9216);
nor U13654 (N_13654,N_7894,N_9008);
xor U13655 (N_13655,N_5123,N_5297);
xor U13656 (N_13656,N_5849,N_7609);
xnor U13657 (N_13657,N_8462,N_8916);
nor U13658 (N_13658,N_8113,N_5458);
nand U13659 (N_13659,N_8597,N_5491);
xor U13660 (N_13660,N_9299,N_9188);
nor U13661 (N_13661,N_8659,N_5966);
xnor U13662 (N_13662,N_6781,N_6848);
or U13663 (N_13663,N_5520,N_7862);
xor U13664 (N_13664,N_8760,N_9932);
nor U13665 (N_13665,N_7647,N_9136);
and U13666 (N_13666,N_8373,N_6242);
xor U13667 (N_13667,N_5835,N_6341);
xor U13668 (N_13668,N_7054,N_7159);
or U13669 (N_13669,N_8568,N_9933);
and U13670 (N_13670,N_7305,N_9468);
nor U13671 (N_13671,N_8455,N_5938);
nor U13672 (N_13672,N_9906,N_9323);
and U13673 (N_13673,N_7911,N_5906);
xor U13674 (N_13674,N_8328,N_6442);
or U13675 (N_13675,N_8599,N_5074);
nor U13676 (N_13676,N_6737,N_6906);
nand U13677 (N_13677,N_6829,N_7715);
and U13678 (N_13678,N_7795,N_6569);
nor U13679 (N_13679,N_8901,N_8563);
xnor U13680 (N_13680,N_8633,N_6233);
and U13681 (N_13681,N_7897,N_8788);
nor U13682 (N_13682,N_8635,N_6145);
nor U13683 (N_13683,N_5144,N_7236);
nand U13684 (N_13684,N_8693,N_8921);
nand U13685 (N_13685,N_6518,N_5859);
and U13686 (N_13686,N_5896,N_9291);
and U13687 (N_13687,N_5765,N_5177);
xor U13688 (N_13688,N_5676,N_6273);
or U13689 (N_13689,N_9777,N_7073);
nor U13690 (N_13690,N_8200,N_9018);
nor U13691 (N_13691,N_9106,N_5119);
nor U13692 (N_13692,N_8582,N_5717);
nand U13693 (N_13693,N_7636,N_7223);
or U13694 (N_13694,N_9697,N_7400);
or U13695 (N_13695,N_8568,N_5619);
or U13696 (N_13696,N_9659,N_6326);
xor U13697 (N_13697,N_6515,N_6972);
nor U13698 (N_13698,N_7220,N_7934);
nand U13699 (N_13699,N_7068,N_8957);
or U13700 (N_13700,N_8403,N_7147);
nand U13701 (N_13701,N_6051,N_9640);
nand U13702 (N_13702,N_5363,N_9643);
nor U13703 (N_13703,N_8998,N_8084);
and U13704 (N_13704,N_7721,N_5270);
nand U13705 (N_13705,N_6454,N_9878);
xor U13706 (N_13706,N_6007,N_9562);
xnor U13707 (N_13707,N_8239,N_8965);
nor U13708 (N_13708,N_6336,N_6196);
nand U13709 (N_13709,N_7802,N_6256);
or U13710 (N_13710,N_7135,N_5498);
xnor U13711 (N_13711,N_8882,N_5255);
nand U13712 (N_13712,N_8772,N_9373);
or U13713 (N_13713,N_9919,N_8725);
xnor U13714 (N_13714,N_6143,N_5834);
nor U13715 (N_13715,N_7880,N_9160);
or U13716 (N_13716,N_5900,N_7023);
or U13717 (N_13717,N_7960,N_9367);
nor U13718 (N_13718,N_6134,N_8911);
nor U13719 (N_13719,N_8314,N_5294);
xor U13720 (N_13720,N_8548,N_9779);
and U13721 (N_13721,N_7535,N_8034);
nor U13722 (N_13722,N_9370,N_5592);
nor U13723 (N_13723,N_8933,N_9107);
and U13724 (N_13724,N_6223,N_5227);
nand U13725 (N_13725,N_8723,N_9252);
nand U13726 (N_13726,N_8373,N_6203);
xnor U13727 (N_13727,N_9181,N_8912);
and U13728 (N_13728,N_9297,N_8018);
and U13729 (N_13729,N_9707,N_8115);
nand U13730 (N_13730,N_7326,N_9417);
nand U13731 (N_13731,N_5954,N_8750);
or U13732 (N_13732,N_5316,N_5198);
nand U13733 (N_13733,N_5642,N_8688);
or U13734 (N_13734,N_6372,N_9448);
nand U13735 (N_13735,N_9873,N_9344);
and U13736 (N_13736,N_8853,N_5496);
nand U13737 (N_13737,N_6656,N_5826);
nand U13738 (N_13738,N_5139,N_7830);
nor U13739 (N_13739,N_9017,N_6105);
and U13740 (N_13740,N_9285,N_7758);
or U13741 (N_13741,N_8499,N_8420);
and U13742 (N_13742,N_8111,N_7211);
nand U13743 (N_13743,N_7901,N_6144);
nor U13744 (N_13744,N_7546,N_6951);
and U13745 (N_13745,N_5393,N_6299);
nor U13746 (N_13746,N_9575,N_9427);
or U13747 (N_13747,N_7295,N_5811);
nand U13748 (N_13748,N_9674,N_9486);
nand U13749 (N_13749,N_7694,N_5972);
nand U13750 (N_13750,N_6121,N_6369);
or U13751 (N_13751,N_8254,N_7617);
nand U13752 (N_13752,N_8817,N_5699);
nand U13753 (N_13753,N_7163,N_6510);
xor U13754 (N_13754,N_6625,N_6677);
xor U13755 (N_13755,N_9293,N_9950);
and U13756 (N_13756,N_5726,N_9736);
or U13757 (N_13757,N_7500,N_7690);
or U13758 (N_13758,N_9656,N_9674);
nor U13759 (N_13759,N_9107,N_8987);
nand U13760 (N_13760,N_9437,N_6754);
xor U13761 (N_13761,N_5918,N_5982);
nor U13762 (N_13762,N_6727,N_9529);
nand U13763 (N_13763,N_5839,N_7909);
nand U13764 (N_13764,N_7318,N_6344);
nand U13765 (N_13765,N_9336,N_8955);
and U13766 (N_13766,N_6230,N_9737);
or U13767 (N_13767,N_5440,N_5708);
and U13768 (N_13768,N_5570,N_5382);
or U13769 (N_13769,N_6084,N_6541);
nand U13770 (N_13770,N_5057,N_5829);
nor U13771 (N_13771,N_7876,N_6599);
xor U13772 (N_13772,N_6382,N_9859);
nand U13773 (N_13773,N_6058,N_8232);
nand U13774 (N_13774,N_7133,N_7834);
or U13775 (N_13775,N_8171,N_5430);
nor U13776 (N_13776,N_9883,N_9244);
nand U13777 (N_13777,N_7551,N_7039);
and U13778 (N_13778,N_9548,N_9925);
nand U13779 (N_13779,N_8665,N_5360);
nand U13780 (N_13780,N_9098,N_6892);
nor U13781 (N_13781,N_5138,N_8889);
nand U13782 (N_13782,N_6807,N_8513);
or U13783 (N_13783,N_5198,N_6263);
nand U13784 (N_13784,N_8878,N_6248);
xnor U13785 (N_13785,N_5293,N_9814);
and U13786 (N_13786,N_8172,N_6093);
xor U13787 (N_13787,N_6043,N_5084);
and U13788 (N_13788,N_6273,N_5819);
nor U13789 (N_13789,N_9592,N_6720);
nand U13790 (N_13790,N_7809,N_7923);
nand U13791 (N_13791,N_7535,N_5912);
or U13792 (N_13792,N_8358,N_6321);
nand U13793 (N_13793,N_9038,N_6126);
nor U13794 (N_13794,N_9454,N_6160);
nand U13795 (N_13795,N_8919,N_9175);
xnor U13796 (N_13796,N_6852,N_7887);
and U13797 (N_13797,N_9702,N_6614);
and U13798 (N_13798,N_7513,N_7994);
and U13799 (N_13799,N_5747,N_6828);
and U13800 (N_13800,N_6658,N_8762);
nor U13801 (N_13801,N_5519,N_8333);
nand U13802 (N_13802,N_5463,N_5086);
nor U13803 (N_13803,N_7303,N_8007);
or U13804 (N_13804,N_7513,N_5991);
xnor U13805 (N_13805,N_6108,N_6589);
and U13806 (N_13806,N_5892,N_6541);
nand U13807 (N_13807,N_6483,N_9535);
nor U13808 (N_13808,N_9982,N_5937);
or U13809 (N_13809,N_7320,N_7485);
nand U13810 (N_13810,N_8655,N_6734);
and U13811 (N_13811,N_9937,N_6993);
and U13812 (N_13812,N_5139,N_8781);
xor U13813 (N_13813,N_6057,N_7819);
or U13814 (N_13814,N_5994,N_7226);
and U13815 (N_13815,N_8567,N_8856);
or U13816 (N_13816,N_9332,N_5979);
nor U13817 (N_13817,N_7279,N_8187);
nand U13818 (N_13818,N_5935,N_5207);
nand U13819 (N_13819,N_7063,N_9171);
xor U13820 (N_13820,N_7762,N_6323);
or U13821 (N_13821,N_6417,N_5192);
nor U13822 (N_13822,N_8735,N_7419);
and U13823 (N_13823,N_9510,N_6372);
and U13824 (N_13824,N_9254,N_8493);
or U13825 (N_13825,N_8341,N_8807);
and U13826 (N_13826,N_9881,N_7398);
nand U13827 (N_13827,N_5066,N_5367);
and U13828 (N_13828,N_5043,N_5748);
nand U13829 (N_13829,N_9648,N_9443);
or U13830 (N_13830,N_8371,N_8539);
and U13831 (N_13831,N_9918,N_7832);
and U13832 (N_13832,N_5440,N_8018);
or U13833 (N_13833,N_9046,N_6090);
and U13834 (N_13834,N_5117,N_9372);
nor U13835 (N_13835,N_7778,N_5201);
xor U13836 (N_13836,N_6490,N_7051);
or U13837 (N_13837,N_6896,N_7567);
nand U13838 (N_13838,N_9367,N_7609);
nor U13839 (N_13839,N_5279,N_9826);
xor U13840 (N_13840,N_6944,N_7046);
nor U13841 (N_13841,N_9769,N_7467);
and U13842 (N_13842,N_8904,N_5361);
nand U13843 (N_13843,N_5220,N_8135);
or U13844 (N_13844,N_6688,N_6351);
xor U13845 (N_13845,N_7983,N_7677);
and U13846 (N_13846,N_5781,N_8923);
or U13847 (N_13847,N_7175,N_6371);
nand U13848 (N_13848,N_6111,N_9126);
and U13849 (N_13849,N_5825,N_6199);
xnor U13850 (N_13850,N_7307,N_8921);
or U13851 (N_13851,N_5443,N_5788);
nand U13852 (N_13852,N_9039,N_5882);
nand U13853 (N_13853,N_8441,N_8052);
or U13854 (N_13854,N_6584,N_7530);
nor U13855 (N_13855,N_7196,N_9023);
nor U13856 (N_13856,N_9358,N_9105);
nand U13857 (N_13857,N_9340,N_8576);
nand U13858 (N_13858,N_7376,N_8446);
nor U13859 (N_13859,N_8566,N_5502);
xnor U13860 (N_13860,N_7572,N_8960);
nor U13861 (N_13861,N_8490,N_7261);
nand U13862 (N_13862,N_7576,N_7790);
nor U13863 (N_13863,N_7617,N_9422);
nand U13864 (N_13864,N_8914,N_5241);
nand U13865 (N_13865,N_6342,N_9140);
nand U13866 (N_13866,N_5859,N_5834);
xor U13867 (N_13867,N_5979,N_5899);
xor U13868 (N_13868,N_7286,N_8478);
or U13869 (N_13869,N_7050,N_6099);
xnor U13870 (N_13870,N_8195,N_5594);
nor U13871 (N_13871,N_8785,N_5250);
and U13872 (N_13872,N_5024,N_6250);
and U13873 (N_13873,N_8174,N_7534);
and U13874 (N_13874,N_7396,N_5995);
nor U13875 (N_13875,N_8436,N_8276);
xor U13876 (N_13876,N_7083,N_8005);
xor U13877 (N_13877,N_8396,N_8405);
or U13878 (N_13878,N_9459,N_7356);
or U13879 (N_13879,N_8225,N_5805);
and U13880 (N_13880,N_9184,N_8526);
nor U13881 (N_13881,N_5576,N_6480);
and U13882 (N_13882,N_9056,N_6204);
and U13883 (N_13883,N_6393,N_5584);
nor U13884 (N_13884,N_7133,N_5567);
nor U13885 (N_13885,N_8059,N_9662);
xor U13886 (N_13886,N_5945,N_7345);
or U13887 (N_13887,N_6031,N_7486);
xnor U13888 (N_13888,N_9996,N_6942);
xnor U13889 (N_13889,N_7129,N_9281);
and U13890 (N_13890,N_6217,N_9581);
nand U13891 (N_13891,N_5400,N_9914);
nand U13892 (N_13892,N_6499,N_8156);
nor U13893 (N_13893,N_6436,N_7903);
and U13894 (N_13894,N_9047,N_5340);
nand U13895 (N_13895,N_7285,N_7498);
xor U13896 (N_13896,N_9560,N_9654);
and U13897 (N_13897,N_5283,N_8080);
nor U13898 (N_13898,N_9641,N_9623);
and U13899 (N_13899,N_5826,N_9984);
xnor U13900 (N_13900,N_5713,N_9743);
nand U13901 (N_13901,N_5590,N_6098);
or U13902 (N_13902,N_5942,N_6778);
nand U13903 (N_13903,N_5733,N_6604);
nand U13904 (N_13904,N_8915,N_6810);
nand U13905 (N_13905,N_9467,N_8681);
or U13906 (N_13906,N_9951,N_8109);
nand U13907 (N_13907,N_8559,N_9498);
xor U13908 (N_13908,N_7693,N_6916);
xnor U13909 (N_13909,N_9296,N_7104);
and U13910 (N_13910,N_5481,N_6972);
nor U13911 (N_13911,N_7702,N_6984);
xnor U13912 (N_13912,N_7470,N_6676);
and U13913 (N_13913,N_9084,N_6738);
or U13914 (N_13914,N_9606,N_7922);
nand U13915 (N_13915,N_8946,N_8722);
xnor U13916 (N_13916,N_9937,N_9345);
xnor U13917 (N_13917,N_5434,N_7712);
nand U13918 (N_13918,N_6954,N_8020);
nor U13919 (N_13919,N_7753,N_6932);
and U13920 (N_13920,N_8943,N_7819);
and U13921 (N_13921,N_9750,N_5849);
xor U13922 (N_13922,N_6182,N_7452);
xnor U13923 (N_13923,N_6548,N_6896);
and U13924 (N_13924,N_8140,N_8781);
and U13925 (N_13925,N_9104,N_6347);
and U13926 (N_13926,N_8948,N_6862);
nor U13927 (N_13927,N_6423,N_8020);
or U13928 (N_13928,N_9563,N_5394);
nand U13929 (N_13929,N_5789,N_7851);
xor U13930 (N_13930,N_8589,N_7948);
xor U13931 (N_13931,N_6270,N_9666);
xor U13932 (N_13932,N_5523,N_6633);
xnor U13933 (N_13933,N_9344,N_8683);
and U13934 (N_13934,N_8856,N_7825);
nor U13935 (N_13935,N_7037,N_6230);
and U13936 (N_13936,N_7177,N_7134);
and U13937 (N_13937,N_7795,N_9605);
nand U13938 (N_13938,N_9912,N_7065);
and U13939 (N_13939,N_6427,N_6138);
or U13940 (N_13940,N_8226,N_9487);
and U13941 (N_13941,N_9418,N_5072);
or U13942 (N_13942,N_7404,N_6979);
and U13943 (N_13943,N_9187,N_9116);
or U13944 (N_13944,N_5520,N_7383);
xnor U13945 (N_13945,N_6608,N_6003);
and U13946 (N_13946,N_5191,N_5350);
and U13947 (N_13947,N_5080,N_7353);
or U13948 (N_13948,N_7788,N_9766);
and U13949 (N_13949,N_9850,N_5056);
or U13950 (N_13950,N_6605,N_9855);
or U13951 (N_13951,N_6061,N_7210);
or U13952 (N_13952,N_8012,N_9568);
or U13953 (N_13953,N_8087,N_5769);
xor U13954 (N_13954,N_5011,N_5178);
nor U13955 (N_13955,N_8855,N_7594);
nand U13956 (N_13956,N_7884,N_8584);
and U13957 (N_13957,N_9815,N_8638);
nand U13958 (N_13958,N_5705,N_8421);
and U13959 (N_13959,N_5338,N_9010);
and U13960 (N_13960,N_7169,N_5999);
and U13961 (N_13961,N_6074,N_7160);
and U13962 (N_13962,N_7641,N_5722);
and U13963 (N_13963,N_9752,N_8080);
nand U13964 (N_13964,N_8397,N_6469);
nor U13965 (N_13965,N_5052,N_6704);
and U13966 (N_13966,N_8702,N_8604);
xnor U13967 (N_13967,N_6039,N_9804);
and U13968 (N_13968,N_6252,N_7404);
nor U13969 (N_13969,N_7906,N_6726);
and U13970 (N_13970,N_8743,N_9744);
nand U13971 (N_13971,N_5656,N_6616);
or U13972 (N_13972,N_6106,N_5797);
nor U13973 (N_13973,N_7209,N_5338);
nand U13974 (N_13974,N_6489,N_5237);
nor U13975 (N_13975,N_7044,N_8599);
or U13976 (N_13976,N_5089,N_6122);
xor U13977 (N_13977,N_9025,N_6323);
or U13978 (N_13978,N_9182,N_6401);
and U13979 (N_13979,N_5272,N_8507);
nand U13980 (N_13980,N_6480,N_8275);
nand U13981 (N_13981,N_5297,N_8195);
and U13982 (N_13982,N_7009,N_6671);
or U13983 (N_13983,N_9618,N_9187);
nor U13984 (N_13984,N_5205,N_6571);
xor U13985 (N_13985,N_6828,N_8105);
nand U13986 (N_13986,N_7699,N_8706);
and U13987 (N_13987,N_5845,N_6650);
nor U13988 (N_13988,N_9414,N_9266);
nor U13989 (N_13989,N_5780,N_7343);
xnor U13990 (N_13990,N_6997,N_5488);
or U13991 (N_13991,N_5276,N_6464);
xnor U13992 (N_13992,N_8833,N_8724);
nand U13993 (N_13993,N_6154,N_6394);
nand U13994 (N_13994,N_8341,N_7621);
nand U13995 (N_13995,N_7711,N_9073);
nor U13996 (N_13996,N_7054,N_6303);
and U13997 (N_13997,N_7528,N_6441);
or U13998 (N_13998,N_9339,N_7651);
and U13999 (N_13999,N_6788,N_5794);
or U14000 (N_14000,N_5235,N_8033);
nor U14001 (N_14001,N_7518,N_8751);
xnor U14002 (N_14002,N_8502,N_5547);
and U14003 (N_14003,N_8147,N_7562);
nor U14004 (N_14004,N_6025,N_6045);
xnor U14005 (N_14005,N_5686,N_7944);
xnor U14006 (N_14006,N_5385,N_9240);
nor U14007 (N_14007,N_7500,N_5618);
and U14008 (N_14008,N_7372,N_7198);
or U14009 (N_14009,N_8228,N_6883);
nand U14010 (N_14010,N_8507,N_6715);
nand U14011 (N_14011,N_5300,N_5256);
or U14012 (N_14012,N_9319,N_5338);
nand U14013 (N_14013,N_8077,N_5461);
nor U14014 (N_14014,N_6172,N_5541);
nand U14015 (N_14015,N_5311,N_9009);
and U14016 (N_14016,N_6833,N_9217);
or U14017 (N_14017,N_5246,N_5731);
xor U14018 (N_14018,N_8333,N_9380);
nand U14019 (N_14019,N_6242,N_5325);
nor U14020 (N_14020,N_5675,N_5336);
or U14021 (N_14021,N_6539,N_8378);
or U14022 (N_14022,N_6110,N_5073);
or U14023 (N_14023,N_7806,N_5596);
nor U14024 (N_14024,N_6319,N_6584);
and U14025 (N_14025,N_6882,N_5154);
or U14026 (N_14026,N_5486,N_5489);
or U14027 (N_14027,N_5554,N_6290);
nand U14028 (N_14028,N_7934,N_7908);
nor U14029 (N_14029,N_7673,N_9746);
nand U14030 (N_14030,N_5841,N_5527);
nor U14031 (N_14031,N_6219,N_8629);
or U14032 (N_14032,N_7651,N_5509);
nor U14033 (N_14033,N_9448,N_9869);
or U14034 (N_14034,N_5494,N_5852);
nor U14035 (N_14035,N_5693,N_8105);
xnor U14036 (N_14036,N_8469,N_5423);
or U14037 (N_14037,N_9040,N_6204);
and U14038 (N_14038,N_8963,N_9834);
xor U14039 (N_14039,N_5465,N_8168);
and U14040 (N_14040,N_8427,N_5513);
or U14041 (N_14041,N_7379,N_8388);
and U14042 (N_14042,N_7890,N_9555);
or U14043 (N_14043,N_7422,N_8135);
xor U14044 (N_14044,N_5985,N_5906);
nor U14045 (N_14045,N_7661,N_7109);
or U14046 (N_14046,N_9194,N_9609);
nor U14047 (N_14047,N_9657,N_9991);
and U14048 (N_14048,N_9492,N_9916);
nand U14049 (N_14049,N_9882,N_8150);
xnor U14050 (N_14050,N_7960,N_5046);
and U14051 (N_14051,N_6009,N_8556);
and U14052 (N_14052,N_5199,N_8657);
nand U14053 (N_14053,N_6601,N_6153);
or U14054 (N_14054,N_5828,N_5781);
xnor U14055 (N_14055,N_7477,N_5611);
nand U14056 (N_14056,N_6417,N_7327);
nand U14057 (N_14057,N_6761,N_8029);
xor U14058 (N_14058,N_9795,N_7062);
nand U14059 (N_14059,N_7629,N_8629);
nor U14060 (N_14060,N_6154,N_5366);
nand U14061 (N_14061,N_5331,N_8787);
nor U14062 (N_14062,N_6001,N_7843);
or U14063 (N_14063,N_7440,N_5961);
or U14064 (N_14064,N_9406,N_8093);
xnor U14065 (N_14065,N_5676,N_7273);
nand U14066 (N_14066,N_6058,N_6178);
or U14067 (N_14067,N_8026,N_6168);
xor U14068 (N_14068,N_9394,N_5706);
or U14069 (N_14069,N_6310,N_6594);
or U14070 (N_14070,N_6933,N_7594);
and U14071 (N_14071,N_9922,N_7471);
nand U14072 (N_14072,N_8990,N_6258);
xor U14073 (N_14073,N_8081,N_7505);
xor U14074 (N_14074,N_7601,N_9363);
xor U14075 (N_14075,N_5901,N_8479);
and U14076 (N_14076,N_7478,N_6000);
nand U14077 (N_14077,N_9277,N_6384);
nand U14078 (N_14078,N_9909,N_5319);
xor U14079 (N_14079,N_8752,N_5849);
and U14080 (N_14080,N_7211,N_5824);
nor U14081 (N_14081,N_6243,N_7606);
xnor U14082 (N_14082,N_7938,N_9876);
xnor U14083 (N_14083,N_6113,N_6376);
nor U14084 (N_14084,N_8447,N_5340);
xor U14085 (N_14085,N_9743,N_9233);
nand U14086 (N_14086,N_8659,N_6166);
xnor U14087 (N_14087,N_9253,N_6089);
or U14088 (N_14088,N_5716,N_6304);
or U14089 (N_14089,N_7707,N_6358);
nor U14090 (N_14090,N_8288,N_5540);
xnor U14091 (N_14091,N_8809,N_7864);
and U14092 (N_14092,N_5074,N_9707);
nor U14093 (N_14093,N_7405,N_6351);
and U14094 (N_14094,N_8055,N_8562);
nor U14095 (N_14095,N_9970,N_6326);
xnor U14096 (N_14096,N_8007,N_5566);
xor U14097 (N_14097,N_7904,N_7866);
and U14098 (N_14098,N_9488,N_5976);
or U14099 (N_14099,N_9443,N_7613);
nor U14100 (N_14100,N_5942,N_9497);
nor U14101 (N_14101,N_9262,N_7452);
or U14102 (N_14102,N_9257,N_9395);
xor U14103 (N_14103,N_5066,N_7939);
nor U14104 (N_14104,N_5293,N_7572);
and U14105 (N_14105,N_7417,N_5542);
and U14106 (N_14106,N_7904,N_9293);
nand U14107 (N_14107,N_8264,N_8695);
xnor U14108 (N_14108,N_5103,N_6094);
and U14109 (N_14109,N_7806,N_7793);
or U14110 (N_14110,N_5742,N_5553);
nor U14111 (N_14111,N_8745,N_8466);
nand U14112 (N_14112,N_6918,N_5669);
nand U14113 (N_14113,N_6254,N_7312);
nand U14114 (N_14114,N_8532,N_9682);
or U14115 (N_14115,N_9815,N_7771);
or U14116 (N_14116,N_6227,N_6142);
and U14117 (N_14117,N_5153,N_6369);
nand U14118 (N_14118,N_6330,N_8068);
xor U14119 (N_14119,N_9432,N_9316);
and U14120 (N_14120,N_6821,N_5690);
nor U14121 (N_14121,N_9473,N_9919);
nor U14122 (N_14122,N_5221,N_7284);
and U14123 (N_14123,N_7374,N_8628);
and U14124 (N_14124,N_7971,N_6411);
and U14125 (N_14125,N_9254,N_9131);
xnor U14126 (N_14126,N_5199,N_9385);
nand U14127 (N_14127,N_6040,N_7574);
xor U14128 (N_14128,N_7719,N_9152);
nor U14129 (N_14129,N_7545,N_9361);
and U14130 (N_14130,N_8275,N_7433);
and U14131 (N_14131,N_7732,N_8151);
nand U14132 (N_14132,N_7967,N_9424);
nor U14133 (N_14133,N_8363,N_6854);
and U14134 (N_14134,N_6786,N_9235);
and U14135 (N_14135,N_8009,N_5170);
or U14136 (N_14136,N_9697,N_9001);
and U14137 (N_14137,N_9858,N_6979);
nand U14138 (N_14138,N_5711,N_5917);
nand U14139 (N_14139,N_5811,N_7460);
or U14140 (N_14140,N_8401,N_6287);
or U14141 (N_14141,N_8834,N_7135);
or U14142 (N_14142,N_7558,N_5923);
and U14143 (N_14143,N_9319,N_8528);
or U14144 (N_14144,N_6125,N_5009);
nor U14145 (N_14145,N_5712,N_5740);
or U14146 (N_14146,N_8415,N_9770);
or U14147 (N_14147,N_9801,N_8866);
xnor U14148 (N_14148,N_7222,N_7067);
nand U14149 (N_14149,N_9032,N_7784);
or U14150 (N_14150,N_7689,N_7046);
nor U14151 (N_14151,N_8021,N_8858);
xnor U14152 (N_14152,N_9260,N_8479);
and U14153 (N_14153,N_7455,N_8452);
and U14154 (N_14154,N_9101,N_9985);
or U14155 (N_14155,N_7579,N_9356);
and U14156 (N_14156,N_7150,N_7311);
or U14157 (N_14157,N_9160,N_7050);
and U14158 (N_14158,N_6322,N_5804);
and U14159 (N_14159,N_5433,N_8182);
or U14160 (N_14160,N_5290,N_7718);
xor U14161 (N_14161,N_9148,N_9384);
nand U14162 (N_14162,N_5447,N_9328);
and U14163 (N_14163,N_7048,N_7137);
nand U14164 (N_14164,N_9997,N_5097);
nand U14165 (N_14165,N_8781,N_6746);
nor U14166 (N_14166,N_7164,N_5180);
xnor U14167 (N_14167,N_8379,N_5276);
xnor U14168 (N_14168,N_6226,N_7131);
nor U14169 (N_14169,N_7729,N_9012);
or U14170 (N_14170,N_8487,N_8113);
nor U14171 (N_14171,N_8215,N_9466);
or U14172 (N_14172,N_9632,N_7523);
and U14173 (N_14173,N_6285,N_9495);
xnor U14174 (N_14174,N_5119,N_5985);
nand U14175 (N_14175,N_6831,N_8922);
and U14176 (N_14176,N_5128,N_7339);
nor U14177 (N_14177,N_8648,N_9453);
or U14178 (N_14178,N_8999,N_7608);
nand U14179 (N_14179,N_6264,N_6185);
and U14180 (N_14180,N_7151,N_9044);
nand U14181 (N_14181,N_8873,N_6663);
and U14182 (N_14182,N_5865,N_8759);
nor U14183 (N_14183,N_5413,N_8854);
xnor U14184 (N_14184,N_9920,N_6316);
or U14185 (N_14185,N_5054,N_7584);
xor U14186 (N_14186,N_9568,N_9588);
or U14187 (N_14187,N_9384,N_5010);
or U14188 (N_14188,N_7742,N_5199);
nor U14189 (N_14189,N_6416,N_5396);
or U14190 (N_14190,N_5642,N_8557);
nand U14191 (N_14191,N_6679,N_9646);
and U14192 (N_14192,N_9572,N_8764);
nor U14193 (N_14193,N_8952,N_5021);
or U14194 (N_14194,N_6613,N_9510);
xnor U14195 (N_14195,N_8664,N_9714);
nand U14196 (N_14196,N_8921,N_6956);
nor U14197 (N_14197,N_9999,N_8981);
nor U14198 (N_14198,N_8401,N_8105);
nand U14199 (N_14199,N_7226,N_5770);
nand U14200 (N_14200,N_8118,N_9889);
nand U14201 (N_14201,N_7901,N_8134);
xor U14202 (N_14202,N_6883,N_9933);
and U14203 (N_14203,N_6470,N_6068);
or U14204 (N_14204,N_7232,N_7977);
xnor U14205 (N_14205,N_9750,N_5753);
and U14206 (N_14206,N_8518,N_8975);
nand U14207 (N_14207,N_9227,N_8641);
nand U14208 (N_14208,N_8520,N_7838);
nand U14209 (N_14209,N_7797,N_7514);
or U14210 (N_14210,N_9644,N_6767);
and U14211 (N_14211,N_7026,N_5035);
or U14212 (N_14212,N_9343,N_6138);
nor U14213 (N_14213,N_6740,N_8355);
nor U14214 (N_14214,N_8683,N_8856);
and U14215 (N_14215,N_7375,N_6210);
xnor U14216 (N_14216,N_5478,N_8505);
nor U14217 (N_14217,N_6151,N_6656);
and U14218 (N_14218,N_7011,N_8010);
and U14219 (N_14219,N_7728,N_9263);
nor U14220 (N_14220,N_8592,N_9667);
nand U14221 (N_14221,N_5108,N_9101);
nor U14222 (N_14222,N_5425,N_7414);
nor U14223 (N_14223,N_5617,N_9894);
nor U14224 (N_14224,N_5960,N_9664);
xor U14225 (N_14225,N_6943,N_7022);
nand U14226 (N_14226,N_8353,N_6619);
and U14227 (N_14227,N_5314,N_5456);
nand U14228 (N_14228,N_6544,N_7641);
or U14229 (N_14229,N_6728,N_6777);
nor U14230 (N_14230,N_9915,N_5286);
nor U14231 (N_14231,N_8461,N_9054);
nor U14232 (N_14232,N_6651,N_8976);
xor U14233 (N_14233,N_8806,N_5344);
and U14234 (N_14234,N_9293,N_5991);
or U14235 (N_14235,N_8380,N_5512);
nand U14236 (N_14236,N_5629,N_7100);
nand U14237 (N_14237,N_5048,N_5750);
and U14238 (N_14238,N_9401,N_9148);
nor U14239 (N_14239,N_5524,N_5568);
or U14240 (N_14240,N_5841,N_7425);
xnor U14241 (N_14241,N_5493,N_8375);
nand U14242 (N_14242,N_5921,N_6623);
xnor U14243 (N_14243,N_5786,N_8148);
nor U14244 (N_14244,N_5216,N_7897);
or U14245 (N_14245,N_6880,N_9599);
nor U14246 (N_14246,N_6077,N_7228);
and U14247 (N_14247,N_8537,N_6526);
nand U14248 (N_14248,N_6318,N_7350);
xnor U14249 (N_14249,N_7292,N_5306);
nand U14250 (N_14250,N_9263,N_5380);
nor U14251 (N_14251,N_9207,N_7753);
nor U14252 (N_14252,N_5923,N_8042);
xor U14253 (N_14253,N_5838,N_9569);
or U14254 (N_14254,N_5424,N_5157);
and U14255 (N_14255,N_5110,N_5173);
or U14256 (N_14256,N_6175,N_5724);
and U14257 (N_14257,N_5251,N_6736);
nor U14258 (N_14258,N_6630,N_7044);
nand U14259 (N_14259,N_6238,N_6314);
nand U14260 (N_14260,N_8551,N_5192);
and U14261 (N_14261,N_5167,N_7150);
nand U14262 (N_14262,N_7466,N_5623);
nor U14263 (N_14263,N_6273,N_6382);
nor U14264 (N_14264,N_8019,N_5837);
xnor U14265 (N_14265,N_9966,N_7761);
nor U14266 (N_14266,N_9538,N_7615);
or U14267 (N_14267,N_5810,N_9801);
nand U14268 (N_14268,N_5635,N_7522);
and U14269 (N_14269,N_5732,N_6445);
nor U14270 (N_14270,N_8880,N_7729);
or U14271 (N_14271,N_9834,N_9499);
or U14272 (N_14272,N_9572,N_7115);
nand U14273 (N_14273,N_9840,N_8403);
or U14274 (N_14274,N_7157,N_6317);
nor U14275 (N_14275,N_7468,N_8362);
nor U14276 (N_14276,N_5756,N_7921);
nand U14277 (N_14277,N_6376,N_5233);
and U14278 (N_14278,N_6258,N_9960);
and U14279 (N_14279,N_9750,N_7006);
nand U14280 (N_14280,N_9600,N_8897);
nand U14281 (N_14281,N_9285,N_7716);
nand U14282 (N_14282,N_8396,N_8565);
xor U14283 (N_14283,N_5426,N_6857);
xor U14284 (N_14284,N_9867,N_6191);
nand U14285 (N_14285,N_6084,N_9212);
xor U14286 (N_14286,N_9290,N_7219);
xor U14287 (N_14287,N_5256,N_6862);
nand U14288 (N_14288,N_6232,N_8951);
and U14289 (N_14289,N_8388,N_7865);
or U14290 (N_14290,N_6769,N_6526);
nand U14291 (N_14291,N_5394,N_6637);
nor U14292 (N_14292,N_5895,N_7829);
xor U14293 (N_14293,N_7267,N_6274);
or U14294 (N_14294,N_7606,N_8557);
and U14295 (N_14295,N_7454,N_7903);
or U14296 (N_14296,N_7340,N_8875);
or U14297 (N_14297,N_5249,N_8237);
xor U14298 (N_14298,N_7356,N_8416);
and U14299 (N_14299,N_9602,N_6457);
nand U14300 (N_14300,N_6611,N_8247);
nand U14301 (N_14301,N_5675,N_6113);
xor U14302 (N_14302,N_8118,N_5074);
and U14303 (N_14303,N_8464,N_5478);
xnor U14304 (N_14304,N_6602,N_6192);
and U14305 (N_14305,N_9256,N_7180);
or U14306 (N_14306,N_5394,N_8064);
or U14307 (N_14307,N_5896,N_7268);
or U14308 (N_14308,N_5513,N_5319);
xor U14309 (N_14309,N_5977,N_7257);
nor U14310 (N_14310,N_7516,N_8610);
nand U14311 (N_14311,N_7707,N_6059);
nor U14312 (N_14312,N_7868,N_5749);
nand U14313 (N_14313,N_9228,N_8056);
xor U14314 (N_14314,N_9672,N_7976);
nand U14315 (N_14315,N_5982,N_5505);
and U14316 (N_14316,N_9782,N_6972);
nor U14317 (N_14317,N_8478,N_9112);
and U14318 (N_14318,N_9801,N_6305);
or U14319 (N_14319,N_8123,N_8188);
xor U14320 (N_14320,N_5150,N_7491);
nand U14321 (N_14321,N_9894,N_8554);
xnor U14322 (N_14322,N_8820,N_6631);
nor U14323 (N_14323,N_9763,N_5780);
nor U14324 (N_14324,N_8390,N_8013);
nand U14325 (N_14325,N_6435,N_7503);
nand U14326 (N_14326,N_9533,N_6164);
xor U14327 (N_14327,N_5505,N_7815);
and U14328 (N_14328,N_9868,N_6081);
xor U14329 (N_14329,N_8131,N_8410);
nand U14330 (N_14330,N_7195,N_9968);
or U14331 (N_14331,N_5267,N_5206);
or U14332 (N_14332,N_5948,N_8115);
xnor U14333 (N_14333,N_5541,N_5834);
nand U14334 (N_14334,N_9516,N_9044);
nand U14335 (N_14335,N_6283,N_5134);
or U14336 (N_14336,N_7436,N_9722);
and U14337 (N_14337,N_9042,N_8498);
nand U14338 (N_14338,N_8839,N_9341);
nand U14339 (N_14339,N_7819,N_8962);
and U14340 (N_14340,N_9911,N_8322);
and U14341 (N_14341,N_6207,N_6964);
nand U14342 (N_14342,N_5983,N_5693);
nor U14343 (N_14343,N_5296,N_6989);
nand U14344 (N_14344,N_6442,N_6627);
or U14345 (N_14345,N_5297,N_9623);
nand U14346 (N_14346,N_5845,N_6524);
nand U14347 (N_14347,N_5963,N_8268);
nor U14348 (N_14348,N_8509,N_9557);
nand U14349 (N_14349,N_5515,N_9782);
nand U14350 (N_14350,N_9248,N_9703);
and U14351 (N_14351,N_8734,N_5907);
nand U14352 (N_14352,N_7263,N_5416);
xnor U14353 (N_14353,N_9111,N_8572);
or U14354 (N_14354,N_9242,N_5940);
xnor U14355 (N_14355,N_6307,N_6021);
and U14356 (N_14356,N_5435,N_9761);
nand U14357 (N_14357,N_5256,N_5347);
or U14358 (N_14358,N_9560,N_5419);
xor U14359 (N_14359,N_5791,N_6492);
and U14360 (N_14360,N_8549,N_9172);
xnor U14361 (N_14361,N_6697,N_6719);
nor U14362 (N_14362,N_6120,N_8530);
xor U14363 (N_14363,N_8347,N_5685);
or U14364 (N_14364,N_5667,N_8460);
and U14365 (N_14365,N_5966,N_5853);
nand U14366 (N_14366,N_5940,N_9279);
or U14367 (N_14367,N_5774,N_8563);
and U14368 (N_14368,N_5271,N_7421);
nor U14369 (N_14369,N_9942,N_9661);
nand U14370 (N_14370,N_7762,N_9568);
nand U14371 (N_14371,N_6322,N_8644);
and U14372 (N_14372,N_8413,N_8883);
and U14373 (N_14373,N_6512,N_9431);
xor U14374 (N_14374,N_8986,N_5824);
nand U14375 (N_14375,N_9833,N_9749);
and U14376 (N_14376,N_5848,N_8268);
or U14377 (N_14377,N_6133,N_5411);
or U14378 (N_14378,N_8217,N_9147);
nor U14379 (N_14379,N_6168,N_7306);
or U14380 (N_14380,N_7518,N_6583);
nor U14381 (N_14381,N_9656,N_8396);
nor U14382 (N_14382,N_9301,N_8379);
and U14383 (N_14383,N_8896,N_8272);
nand U14384 (N_14384,N_7465,N_5434);
xor U14385 (N_14385,N_6771,N_9549);
nor U14386 (N_14386,N_8680,N_5750);
nand U14387 (N_14387,N_8235,N_9111);
and U14388 (N_14388,N_7792,N_9777);
xor U14389 (N_14389,N_5753,N_5179);
or U14390 (N_14390,N_5564,N_9169);
and U14391 (N_14391,N_9619,N_6165);
xor U14392 (N_14392,N_8226,N_5263);
nand U14393 (N_14393,N_9406,N_8781);
xor U14394 (N_14394,N_5480,N_8814);
nor U14395 (N_14395,N_7677,N_9448);
xnor U14396 (N_14396,N_5046,N_8422);
or U14397 (N_14397,N_6822,N_7625);
and U14398 (N_14398,N_9063,N_7131);
xnor U14399 (N_14399,N_8837,N_6950);
nor U14400 (N_14400,N_6200,N_9634);
nor U14401 (N_14401,N_8277,N_9993);
or U14402 (N_14402,N_7905,N_7975);
and U14403 (N_14403,N_6460,N_8884);
nand U14404 (N_14404,N_9734,N_8957);
xnor U14405 (N_14405,N_6790,N_6547);
nand U14406 (N_14406,N_8582,N_9367);
xor U14407 (N_14407,N_7834,N_9773);
nand U14408 (N_14408,N_8925,N_7154);
and U14409 (N_14409,N_7534,N_8959);
and U14410 (N_14410,N_9613,N_8282);
nand U14411 (N_14411,N_6035,N_5909);
xnor U14412 (N_14412,N_9625,N_6325);
nand U14413 (N_14413,N_7330,N_8595);
nand U14414 (N_14414,N_9617,N_7909);
xor U14415 (N_14415,N_8553,N_8787);
nand U14416 (N_14416,N_8556,N_5203);
nor U14417 (N_14417,N_8617,N_5250);
or U14418 (N_14418,N_6349,N_9235);
nor U14419 (N_14419,N_8119,N_5186);
nand U14420 (N_14420,N_6138,N_5402);
nand U14421 (N_14421,N_5335,N_8685);
nor U14422 (N_14422,N_7897,N_5648);
nand U14423 (N_14423,N_5962,N_9962);
nor U14424 (N_14424,N_9671,N_7739);
or U14425 (N_14425,N_6272,N_6093);
xnor U14426 (N_14426,N_8690,N_7850);
xnor U14427 (N_14427,N_8189,N_7736);
nor U14428 (N_14428,N_5759,N_8598);
xor U14429 (N_14429,N_9955,N_8590);
xor U14430 (N_14430,N_9552,N_8135);
nand U14431 (N_14431,N_9657,N_5727);
and U14432 (N_14432,N_7992,N_6297);
nor U14433 (N_14433,N_8804,N_9681);
or U14434 (N_14434,N_8617,N_9149);
xnor U14435 (N_14435,N_7272,N_5397);
nand U14436 (N_14436,N_5160,N_5855);
or U14437 (N_14437,N_6366,N_8356);
or U14438 (N_14438,N_7305,N_5975);
xnor U14439 (N_14439,N_9097,N_7828);
xor U14440 (N_14440,N_8168,N_8323);
nor U14441 (N_14441,N_6791,N_5972);
nand U14442 (N_14442,N_8672,N_8172);
xnor U14443 (N_14443,N_6353,N_8378);
nor U14444 (N_14444,N_6861,N_9762);
or U14445 (N_14445,N_7312,N_5582);
xor U14446 (N_14446,N_9364,N_8895);
nand U14447 (N_14447,N_9860,N_8117);
nor U14448 (N_14448,N_6293,N_5649);
and U14449 (N_14449,N_9210,N_8465);
nor U14450 (N_14450,N_7170,N_9216);
xor U14451 (N_14451,N_8665,N_8274);
xnor U14452 (N_14452,N_8508,N_5694);
and U14453 (N_14453,N_9250,N_8741);
and U14454 (N_14454,N_6541,N_6872);
nor U14455 (N_14455,N_9053,N_6766);
nand U14456 (N_14456,N_8821,N_5683);
or U14457 (N_14457,N_7064,N_5497);
nand U14458 (N_14458,N_8733,N_9669);
xnor U14459 (N_14459,N_5691,N_6931);
or U14460 (N_14460,N_5158,N_8128);
or U14461 (N_14461,N_9789,N_9834);
nor U14462 (N_14462,N_8714,N_9984);
and U14463 (N_14463,N_8331,N_7814);
nor U14464 (N_14464,N_7237,N_6766);
xnor U14465 (N_14465,N_8133,N_5842);
xnor U14466 (N_14466,N_8075,N_9737);
xor U14467 (N_14467,N_9832,N_8728);
and U14468 (N_14468,N_5898,N_8731);
or U14469 (N_14469,N_6543,N_5338);
or U14470 (N_14470,N_8141,N_7120);
or U14471 (N_14471,N_7860,N_8125);
xor U14472 (N_14472,N_6886,N_6162);
nor U14473 (N_14473,N_7787,N_8231);
or U14474 (N_14474,N_9850,N_5053);
nand U14475 (N_14475,N_8303,N_5296);
nor U14476 (N_14476,N_9255,N_6526);
nor U14477 (N_14477,N_9844,N_5629);
nor U14478 (N_14478,N_9829,N_5611);
xnor U14479 (N_14479,N_9470,N_7978);
xnor U14480 (N_14480,N_6669,N_9509);
or U14481 (N_14481,N_8463,N_7222);
nor U14482 (N_14482,N_5543,N_5710);
or U14483 (N_14483,N_6583,N_5399);
and U14484 (N_14484,N_9258,N_8046);
and U14485 (N_14485,N_5331,N_8934);
or U14486 (N_14486,N_5652,N_8988);
and U14487 (N_14487,N_9765,N_8867);
or U14488 (N_14488,N_9846,N_6919);
or U14489 (N_14489,N_6364,N_6755);
xor U14490 (N_14490,N_8160,N_9250);
or U14491 (N_14491,N_6656,N_9719);
and U14492 (N_14492,N_5615,N_5708);
nor U14493 (N_14493,N_5118,N_8586);
or U14494 (N_14494,N_9611,N_7113);
and U14495 (N_14495,N_5557,N_8442);
nand U14496 (N_14496,N_5075,N_8167);
nand U14497 (N_14497,N_8169,N_9319);
and U14498 (N_14498,N_9058,N_5896);
nor U14499 (N_14499,N_5462,N_7566);
and U14500 (N_14500,N_7933,N_9061);
or U14501 (N_14501,N_8377,N_5813);
nor U14502 (N_14502,N_8536,N_6499);
nand U14503 (N_14503,N_8521,N_7174);
nand U14504 (N_14504,N_9876,N_6840);
and U14505 (N_14505,N_9001,N_9123);
or U14506 (N_14506,N_7055,N_7881);
xor U14507 (N_14507,N_5069,N_5039);
nor U14508 (N_14508,N_6082,N_8202);
xnor U14509 (N_14509,N_9175,N_7567);
nand U14510 (N_14510,N_7116,N_5963);
nor U14511 (N_14511,N_7652,N_6214);
xor U14512 (N_14512,N_7856,N_6468);
nand U14513 (N_14513,N_9635,N_9523);
nor U14514 (N_14514,N_7137,N_7070);
or U14515 (N_14515,N_9214,N_8128);
nor U14516 (N_14516,N_5644,N_6633);
xnor U14517 (N_14517,N_6757,N_5247);
nor U14518 (N_14518,N_6651,N_7931);
or U14519 (N_14519,N_5663,N_8515);
xnor U14520 (N_14520,N_8703,N_6372);
nand U14521 (N_14521,N_6377,N_8433);
nor U14522 (N_14522,N_9501,N_8587);
or U14523 (N_14523,N_5073,N_9103);
or U14524 (N_14524,N_7344,N_6713);
and U14525 (N_14525,N_8423,N_9859);
nor U14526 (N_14526,N_8005,N_7421);
nand U14527 (N_14527,N_5232,N_6024);
or U14528 (N_14528,N_8041,N_8800);
and U14529 (N_14529,N_8521,N_8857);
and U14530 (N_14530,N_7542,N_9991);
and U14531 (N_14531,N_8342,N_7357);
xor U14532 (N_14532,N_9936,N_9040);
or U14533 (N_14533,N_6601,N_9969);
nor U14534 (N_14534,N_6274,N_9299);
and U14535 (N_14535,N_9711,N_7440);
and U14536 (N_14536,N_5706,N_7139);
nand U14537 (N_14537,N_5964,N_6180);
xor U14538 (N_14538,N_9389,N_6478);
xor U14539 (N_14539,N_8278,N_8334);
or U14540 (N_14540,N_8651,N_8152);
nand U14541 (N_14541,N_5467,N_9416);
nand U14542 (N_14542,N_7234,N_7228);
xor U14543 (N_14543,N_9745,N_5169);
nand U14544 (N_14544,N_6884,N_6951);
nor U14545 (N_14545,N_8076,N_8557);
or U14546 (N_14546,N_6128,N_6455);
and U14547 (N_14547,N_7100,N_5084);
nand U14548 (N_14548,N_6057,N_9282);
or U14549 (N_14549,N_9281,N_7370);
nand U14550 (N_14550,N_8306,N_5305);
and U14551 (N_14551,N_7212,N_6634);
and U14552 (N_14552,N_8451,N_9582);
and U14553 (N_14553,N_9759,N_7980);
nand U14554 (N_14554,N_8013,N_5274);
nand U14555 (N_14555,N_8244,N_9663);
nor U14556 (N_14556,N_8255,N_6006);
nand U14557 (N_14557,N_8039,N_5927);
and U14558 (N_14558,N_7549,N_8192);
nand U14559 (N_14559,N_9175,N_9308);
xnor U14560 (N_14560,N_6581,N_6979);
nor U14561 (N_14561,N_6312,N_7058);
and U14562 (N_14562,N_9453,N_6201);
or U14563 (N_14563,N_9192,N_9500);
or U14564 (N_14564,N_8131,N_7477);
nor U14565 (N_14565,N_7861,N_9863);
nand U14566 (N_14566,N_7757,N_7773);
and U14567 (N_14567,N_5582,N_6429);
nor U14568 (N_14568,N_9799,N_6537);
and U14569 (N_14569,N_5349,N_8462);
and U14570 (N_14570,N_6392,N_9125);
or U14571 (N_14571,N_8720,N_6619);
or U14572 (N_14572,N_6313,N_9143);
xor U14573 (N_14573,N_7829,N_7410);
nor U14574 (N_14574,N_5203,N_9920);
xnor U14575 (N_14575,N_5617,N_6293);
nand U14576 (N_14576,N_7032,N_9867);
nor U14577 (N_14577,N_5104,N_6812);
or U14578 (N_14578,N_9051,N_6779);
xnor U14579 (N_14579,N_9979,N_5276);
xor U14580 (N_14580,N_7684,N_8291);
and U14581 (N_14581,N_9624,N_7373);
nor U14582 (N_14582,N_7315,N_8060);
and U14583 (N_14583,N_7807,N_5071);
and U14584 (N_14584,N_6466,N_8382);
and U14585 (N_14585,N_9454,N_9667);
nor U14586 (N_14586,N_8557,N_6473);
and U14587 (N_14587,N_8082,N_8021);
xor U14588 (N_14588,N_9794,N_6668);
or U14589 (N_14589,N_6145,N_6113);
nor U14590 (N_14590,N_9477,N_6096);
or U14591 (N_14591,N_8845,N_7936);
or U14592 (N_14592,N_5513,N_6003);
xor U14593 (N_14593,N_6627,N_5255);
nand U14594 (N_14594,N_9457,N_9869);
xnor U14595 (N_14595,N_6113,N_6330);
nor U14596 (N_14596,N_5469,N_6395);
xnor U14597 (N_14597,N_6636,N_9718);
or U14598 (N_14598,N_5860,N_5589);
or U14599 (N_14599,N_9314,N_9115);
and U14600 (N_14600,N_9695,N_6098);
nand U14601 (N_14601,N_9618,N_8103);
or U14602 (N_14602,N_7475,N_6383);
nand U14603 (N_14603,N_9243,N_9540);
nor U14604 (N_14604,N_5259,N_8724);
or U14605 (N_14605,N_9559,N_8396);
xnor U14606 (N_14606,N_7725,N_6304);
or U14607 (N_14607,N_8410,N_6886);
or U14608 (N_14608,N_9828,N_5153);
nor U14609 (N_14609,N_5533,N_6370);
nor U14610 (N_14610,N_9186,N_8888);
nor U14611 (N_14611,N_9755,N_7279);
xnor U14612 (N_14612,N_6852,N_9247);
xnor U14613 (N_14613,N_9511,N_6912);
xor U14614 (N_14614,N_8899,N_6452);
nand U14615 (N_14615,N_9358,N_6471);
nand U14616 (N_14616,N_9099,N_6074);
xnor U14617 (N_14617,N_7196,N_8950);
xnor U14618 (N_14618,N_9638,N_5480);
nor U14619 (N_14619,N_9252,N_5840);
or U14620 (N_14620,N_6360,N_5394);
nor U14621 (N_14621,N_6482,N_9106);
xnor U14622 (N_14622,N_6343,N_9148);
and U14623 (N_14623,N_9380,N_7872);
or U14624 (N_14624,N_8875,N_6137);
or U14625 (N_14625,N_8117,N_7888);
nor U14626 (N_14626,N_6989,N_7583);
and U14627 (N_14627,N_6792,N_9634);
xor U14628 (N_14628,N_7285,N_6298);
nand U14629 (N_14629,N_5214,N_6935);
nand U14630 (N_14630,N_8881,N_9076);
or U14631 (N_14631,N_7537,N_6165);
or U14632 (N_14632,N_6845,N_7692);
xnor U14633 (N_14633,N_9920,N_6592);
and U14634 (N_14634,N_8383,N_8369);
nor U14635 (N_14635,N_9411,N_6110);
or U14636 (N_14636,N_6284,N_9443);
xor U14637 (N_14637,N_7737,N_5408);
xnor U14638 (N_14638,N_8366,N_8647);
xor U14639 (N_14639,N_5057,N_5423);
xor U14640 (N_14640,N_8317,N_7561);
xnor U14641 (N_14641,N_7503,N_7447);
nor U14642 (N_14642,N_7915,N_6810);
or U14643 (N_14643,N_5531,N_9941);
xor U14644 (N_14644,N_5529,N_6822);
nor U14645 (N_14645,N_9711,N_6961);
or U14646 (N_14646,N_6003,N_5441);
nand U14647 (N_14647,N_9593,N_6856);
nor U14648 (N_14648,N_6231,N_7378);
and U14649 (N_14649,N_7412,N_7009);
nor U14650 (N_14650,N_6293,N_6691);
or U14651 (N_14651,N_5917,N_7226);
nand U14652 (N_14652,N_8703,N_6192);
nor U14653 (N_14653,N_6465,N_8840);
or U14654 (N_14654,N_6708,N_6002);
xnor U14655 (N_14655,N_6931,N_6815);
or U14656 (N_14656,N_6172,N_8931);
or U14657 (N_14657,N_9462,N_9991);
nor U14658 (N_14658,N_9177,N_9442);
or U14659 (N_14659,N_9302,N_7448);
and U14660 (N_14660,N_5839,N_6698);
xnor U14661 (N_14661,N_9313,N_7433);
xor U14662 (N_14662,N_6035,N_6074);
and U14663 (N_14663,N_9266,N_9623);
nand U14664 (N_14664,N_8832,N_5260);
and U14665 (N_14665,N_8305,N_8112);
xor U14666 (N_14666,N_8101,N_7113);
xor U14667 (N_14667,N_7006,N_8108);
and U14668 (N_14668,N_8802,N_9744);
nor U14669 (N_14669,N_7822,N_7930);
xnor U14670 (N_14670,N_5563,N_7256);
xnor U14671 (N_14671,N_6135,N_6557);
or U14672 (N_14672,N_7607,N_6849);
or U14673 (N_14673,N_9864,N_9926);
or U14674 (N_14674,N_5504,N_9243);
nand U14675 (N_14675,N_8238,N_9516);
or U14676 (N_14676,N_9599,N_5525);
nand U14677 (N_14677,N_6988,N_6632);
xor U14678 (N_14678,N_6687,N_6250);
and U14679 (N_14679,N_9935,N_7666);
xnor U14680 (N_14680,N_7472,N_7771);
nor U14681 (N_14681,N_5487,N_8354);
nor U14682 (N_14682,N_6557,N_7990);
or U14683 (N_14683,N_5148,N_6103);
nor U14684 (N_14684,N_5380,N_9916);
xor U14685 (N_14685,N_8158,N_6282);
xor U14686 (N_14686,N_9673,N_5204);
nor U14687 (N_14687,N_8494,N_6236);
and U14688 (N_14688,N_8801,N_8958);
and U14689 (N_14689,N_5484,N_5553);
xor U14690 (N_14690,N_6311,N_8779);
nand U14691 (N_14691,N_8312,N_9103);
or U14692 (N_14692,N_5485,N_6631);
nor U14693 (N_14693,N_9540,N_8666);
nor U14694 (N_14694,N_7184,N_5603);
xor U14695 (N_14695,N_7629,N_7212);
nand U14696 (N_14696,N_8996,N_8749);
nand U14697 (N_14697,N_7380,N_7208);
or U14698 (N_14698,N_8664,N_5711);
nor U14699 (N_14699,N_5601,N_9033);
and U14700 (N_14700,N_9908,N_9731);
and U14701 (N_14701,N_5971,N_7530);
nand U14702 (N_14702,N_9990,N_5654);
nand U14703 (N_14703,N_7275,N_9142);
or U14704 (N_14704,N_8381,N_9086);
and U14705 (N_14705,N_8726,N_9695);
nor U14706 (N_14706,N_9345,N_5370);
or U14707 (N_14707,N_5850,N_9162);
or U14708 (N_14708,N_6725,N_8917);
nor U14709 (N_14709,N_7030,N_8001);
and U14710 (N_14710,N_8949,N_5090);
nor U14711 (N_14711,N_5299,N_5136);
nor U14712 (N_14712,N_5647,N_7332);
or U14713 (N_14713,N_9007,N_6910);
xnor U14714 (N_14714,N_9900,N_9867);
nand U14715 (N_14715,N_9427,N_6495);
nor U14716 (N_14716,N_6713,N_9504);
xnor U14717 (N_14717,N_5340,N_5393);
nand U14718 (N_14718,N_5576,N_7227);
nand U14719 (N_14719,N_6600,N_6804);
or U14720 (N_14720,N_6708,N_7576);
xnor U14721 (N_14721,N_9047,N_5231);
nand U14722 (N_14722,N_6985,N_5981);
and U14723 (N_14723,N_5040,N_6432);
xnor U14724 (N_14724,N_8551,N_9729);
and U14725 (N_14725,N_8295,N_7878);
or U14726 (N_14726,N_5151,N_9372);
nor U14727 (N_14727,N_7244,N_9295);
or U14728 (N_14728,N_6385,N_5162);
or U14729 (N_14729,N_8920,N_5965);
or U14730 (N_14730,N_8431,N_5020);
or U14731 (N_14731,N_7313,N_6473);
nor U14732 (N_14732,N_7360,N_6077);
nand U14733 (N_14733,N_8600,N_9578);
or U14734 (N_14734,N_8149,N_5262);
nand U14735 (N_14735,N_5286,N_7348);
nor U14736 (N_14736,N_5595,N_6437);
nand U14737 (N_14737,N_8010,N_9927);
nand U14738 (N_14738,N_7505,N_7912);
nand U14739 (N_14739,N_9006,N_5829);
nor U14740 (N_14740,N_9725,N_8937);
or U14741 (N_14741,N_5492,N_6674);
nand U14742 (N_14742,N_9751,N_7270);
xor U14743 (N_14743,N_5258,N_7980);
xnor U14744 (N_14744,N_9568,N_5381);
nor U14745 (N_14745,N_6014,N_9866);
nand U14746 (N_14746,N_7502,N_9121);
nand U14747 (N_14747,N_7970,N_6747);
and U14748 (N_14748,N_8670,N_5302);
or U14749 (N_14749,N_6283,N_5430);
nand U14750 (N_14750,N_6259,N_5508);
and U14751 (N_14751,N_6452,N_8369);
xor U14752 (N_14752,N_8700,N_9224);
xnor U14753 (N_14753,N_5958,N_5943);
and U14754 (N_14754,N_8229,N_8132);
or U14755 (N_14755,N_6658,N_9416);
xor U14756 (N_14756,N_6756,N_5131);
and U14757 (N_14757,N_9535,N_8453);
and U14758 (N_14758,N_8412,N_6469);
xor U14759 (N_14759,N_7246,N_8400);
nor U14760 (N_14760,N_8574,N_5400);
and U14761 (N_14761,N_8983,N_7642);
xnor U14762 (N_14762,N_8426,N_6749);
nand U14763 (N_14763,N_5559,N_8877);
and U14764 (N_14764,N_9044,N_6776);
nand U14765 (N_14765,N_6784,N_9907);
and U14766 (N_14766,N_6265,N_7969);
nor U14767 (N_14767,N_9151,N_9932);
nor U14768 (N_14768,N_7392,N_9205);
xor U14769 (N_14769,N_7644,N_8814);
nand U14770 (N_14770,N_7778,N_6975);
xor U14771 (N_14771,N_7908,N_5497);
nand U14772 (N_14772,N_5133,N_8877);
nor U14773 (N_14773,N_9796,N_5293);
or U14774 (N_14774,N_7494,N_6317);
or U14775 (N_14775,N_8610,N_7080);
xnor U14776 (N_14776,N_6853,N_5266);
or U14777 (N_14777,N_5336,N_7085);
nand U14778 (N_14778,N_6419,N_8726);
nor U14779 (N_14779,N_5466,N_9940);
nor U14780 (N_14780,N_5643,N_7905);
nand U14781 (N_14781,N_8492,N_5496);
nor U14782 (N_14782,N_8048,N_8389);
xor U14783 (N_14783,N_7921,N_6271);
nand U14784 (N_14784,N_7046,N_9004);
or U14785 (N_14785,N_6252,N_9364);
nand U14786 (N_14786,N_6536,N_8795);
nand U14787 (N_14787,N_5774,N_8993);
or U14788 (N_14788,N_5711,N_7958);
nor U14789 (N_14789,N_5256,N_8069);
nand U14790 (N_14790,N_9789,N_8662);
or U14791 (N_14791,N_9322,N_9625);
nand U14792 (N_14792,N_9743,N_8875);
xor U14793 (N_14793,N_5779,N_5507);
xor U14794 (N_14794,N_5620,N_5454);
xor U14795 (N_14795,N_5699,N_6974);
nand U14796 (N_14796,N_7537,N_9413);
or U14797 (N_14797,N_6085,N_9148);
nand U14798 (N_14798,N_6623,N_5064);
or U14799 (N_14799,N_5830,N_5597);
or U14800 (N_14800,N_8590,N_5362);
xnor U14801 (N_14801,N_7417,N_9963);
and U14802 (N_14802,N_7866,N_9222);
or U14803 (N_14803,N_6381,N_7381);
or U14804 (N_14804,N_9886,N_8138);
nand U14805 (N_14805,N_7375,N_9661);
xor U14806 (N_14806,N_8677,N_8498);
nor U14807 (N_14807,N_6576,N_5483);
xnor U14808 (N_14808,N_9116,N_9823);
nand U14809 (N_14809,N_6604,N_9891);
xnor U14810 (N_14810,N_6366,N_6942);
nor U14811 (N_14811,N_9066,N_6300);
nor U14812 (N_14812,N_7194,N_8603);
xnor U14813 (N_14813,N_6544,N_6608);
nor U14814 (N_14814,N_8385,N_9781);
or U14815 (N_14815,N_8705,N_9566);
and U14816 (N_14816,N_9153,N_6293);
nand U14817 (N_14817,N_5170,N_5629);
nor U14818 (N_14818,N_8672,N_9105);
nor U14819 (N_14819,N_6602,N_6517);
nor U14820 (N_14820,N_8891,N_6514);
and U14821 (N_14821,N_7163,N_8842);
xor U14822 (N_14822,N_7715,N_8423);
and U14823 (N_14823,N_6512,N_5450);
and U14824 (N_14824,N_5303,N_8466);
or U14825 (N_14825,N_9302,N_8504);
nor U14826 (N_14826,N_9981,N_9780);
xor U14827 (N_14827,N_5274,N_6235);
and U14828 (N_14828,N_6148,N_8616);
or U14829 (N_14829,N_7784,N_5210);
nand U14830 (N_14830,N_8963,N_5448);
or U14831 (N_14831,N_8219,N_5289);
xor U14832 (N_14832,N_9770,N_7714);
or U14833 (N_14833,N_9075,N_7945);
xnor U14834 (N_14834,N_5178,N_9344);
xnor U14835 (N_14835,N_6585,N_5988);
or U14836 (N_14836,N_7173,N_6970);
nand U14837 (N_14837,N_9978,N_7439);
nand U14838 (N_14838,N_6039,N_8577);
or U14839 (N_14839,N_5461,N_5776);
or U14840 (N_14840,N_6360,N_8672);
or U14841 (N_14841,N_5276,N_9780);
xnor U14842 (N_14842,N_5843,N_6555);
nand U14843 (N_14843,N_7592,N_7053);
nand U14844 (N_14844,N_6113,N_6533);
and U14845 (N_14845,N_9103,N_6931);
nor U14846 (N_14846,N_9510,N_6160);
nor U14847 (N_14847,N_6495,N_6901);
or U14848 (N_14848,N_7678,N_8101);
nand U14849 (N_14849,N_9652,N_7440);
and U14850 (N_14850,N_9127,N_6400);
nor U14851 (N_14851,N_7785,N_5953);
nand U14852 (N_14852,N_6678,N_8915);
or U14853 (N_14853,N_6512,N_6850);
nand U14854 (N_14854,N_7516,N_8517);
or U14855 (N_14855,N_8335,N_5700);
or U14856 (N_14856,N_9395,N_9383);
xnor U14857 (N_14857,N_5506,N_8962);
nand U14858 (N_14858,N_5706,N_5413);
nand U14859 (N_14859,N_6593,N_8456);
or U14860 (N_14860,N_5626,N_7966);
and U14861 (N_14861,N_8217,N_6396);
nand U14862 (N_14862,N_5949,N_6865);
or U14863 (N_14863,N_6561,N_8607);
nor U14864 (N_14864,N_8670,N_5009);
nor U14865 (N_14865,N_6073,N_9918);
or U14866 (N_14866,N_6892,N_6229);
or U14867 (N_14867,N_5279,N_7040);
or U14868 (N_14868,N_6337,N_5543);
nor U14869 (N_14869,N_6113,N_9681);
xnor U14870 (N_14870,N_5674,N_8402);
nand U14871 (N_14871,N_6158,N_9321);
and U14872 (N_14872,N_7018,N_6806);
nand U14873 (N_14873,N_5734,N_7175);
nor U14874 (N_14874,N_8377,N_8690);
or U14875 (N_14875,N_5002,N_5219);
xnor U14876 (N_14876,N_9157,N_7061);
xnor U14877 (N_14877,N_5965,N_8342);
and U14878 (N_14878,N_6300,N_7213);
or U14879 (N_14879,N_9715,N_9130);
and U14880 (N_14880,N_7151,N_6719);
nand U14881 (N_14881,N_5002,N_8036);
or U14882 (N_14882,N_7055,N_7826);
nand U14883 (N_14883,N_9657,N_9446);
nand U14884 (N_14884,N_5430,N_8247);
and U14885 (N_14885,N_7712,N_8680);
xnor U14886 (N_14886,N_5786,N_6933);
nand U14887 (N_14887,N_5564,N_5024);
and U14888 (N_14888,N_7227,N_5124);
xor U14889 (N_14889,N_8972,N_5799);
and U14890 (N_14890,N_6054,N_5302);
nand U14891 (N_14891,N_5426,N_9297);
or U14892 (N_14892,N_5997,N_9666);
nand U14893 (N_14893,N_8650,N_5381);
and U14894 (N_14894,N_6578,N_9711);
nand U14895 (N_14895,N_7168,N_5284);
nand U14896 (N_14896,N_5478,N_5335);
nor U14897 (N_14897,N_6978,N_5651);
xor U14898 (N_14898,N_8490,N_5974);
or U14899 (N_14899,N_5083,N_8950);
nor U14900 (N_14900,N_9525,N_8072);
nand U14901 (N_14901,N_9401,N_5254);
and U14902 (N_14902,N_9725,N_5600);
and U14903 (N_14903,N_6376,N_9234);
nor U14904 (N_14904,N_7144,N_5607);
nor U14905 (N_14905,N_6319,N_6248);
and U14906 (N_14906,N_8393,N_6957);
nor U14907 (N_14907,N_5519,N_8775);
and U14908 (N_14908,N_6050,N_5191);
nand U14909 (N_14909,N_9024,N_5581);
nand U14910 (N_14910,N_7358,N_9792);
and U14911 (N_14911,N_7140,N_7373);
nor U14912 (N_14912,N_9522,N_8207);
nor U14913 (N_14913,N_9105,N_8547);
nor U14914 (N_14914,N_9061,N_6574);
nand U14915 (N_14915,N_6862,N_5094);
and U14916 (N_14916,N_8395,N_7644);
nor U14917 (N_14917,N_5198,N_9649);
nand U14918 (N_14918,N_5160,N_5434);
nor U14919 (N_14919,N_6636,N_6200);
and U14920 (N_14920,N_9394,N_8143);
or U14921 (N_14921,N_5940,N_5590);
nand U14922 (N_14922,N_6013,N_9071);
or U14923 (N_14923,N_8074,N_9001);
xor U14924 (N_14924,N_6738,N_7105);
nand U14925 (N_14925,N_6289,N_9903);
and U14926 (N_14926,N_7370,N_9791);
nor U14927 (N_14927,N_8962,N_5592);
or U14928 (N_14928,N_7796,N_6938);
or U14929 (N_14929,N_6908,N_7836);
nand U14930 (N_14930,N_8664,N_5261);
xnor U14931 (N_14931,N_7792,N_5402);
xnor U14932 (N_14932,N_9686,N_9561);
nor U14933 (N_14933,N_7432,N_6685);
xor U14934 (N_14934,N_7867,N_6501);
nor U14935 (N_14935,N_8871,N_5478);
nor U14936 (N_14936,N_6365,N_8489);
or U14937 (N_14937,N_5315,N_7617);
xor U14938 (N_14938,N_8306,N_5004);
and U14939 (N_14939,N_7970,N_7021);
or U14940 (N_14940,N_6577,N_5334);
nand U14941 (N_14941,N_5276,N_5696);
and U14942 (N_14942,N_7860,N_6150);
or U14943 (N_14943,N_6217,N_6179);
nand U14944 (N_14944,N_6066,N_7096);
xnor U14945 (N_14945,N_5509,N_5850);
or U14946 (N_14946,N_9351,N_7512);
nor U14947 (N_14947,N_8386,N_8740);
and U14948 (N_14948,N_9512,N_6001);
and U14949 (N_14949,N_8839,N_8213);
and U14950 (N_14950,N_8529,N_6979);
nor U14951 (N_14951,N_7284,N_6188);
nand U14952 (N_14952,N_7900,N_5800);
nor U14953 (N_14953,N_9951,N_6781);
nand U14954 (N_14954,N_8017,N_8477);
or U14955 (N_14955,N_5397,N_8032);
nor U14956 (N_14956,N_9622,N_8569);
nor U14957 (N_14957,N_6253,N_8420);
or U14958 (N_14958,N_9095,N_8511);
xor U14959 (N_14959,N_8656,N_7712);
nand U14960 (N_14960,N_6779,N_5487);
xor U14961 (N_14961,N_7193,N_6616);
xor U14962 (N_14962,N_6586,N_7120);
nor U14963 (N_14963,N_7271,N_9002);
and U14964 (N_14964,N_6785,N_7450);
xnor U14965 (N_14965,N_6184,N_9778);
and U14966 (N_14966,N_5554,N_8521);
nor U14967 (N_14967,N_7369,N_8719);
or U14968 (N_14968,N_6930,N_5750);
xor U14969 (N_14969,N_6306,N_5128);
or U14970 (N_14970,N_9772,N_8958);
nor U14971 (N_14971,N_5956,N_8551);
nor U14972 (N_14972,N_6901,N_7603);
and U14973 (N_14973,N_6847,N_9743);
or U14974 (N_14974,N_6409,N_7641);
nand U14975 (N_14975,N_9276,N_8029);
or U14976 (N_14976,N_9648,N_5449);
nand U14977 (N_14977,N_6032,N_9687);
nand U14978 (N_14978,N_5044,N_5315);
nand U14979 (N_14979,N_8705,N_5084);
or U14980 (N_14980,N_6254,N_5993);
or U14981 (N_14981,N_7696,N_7752);
and U14982 (N_14982,N_7227,N_5154);
and U14983 (N_14983,N_7316,N_9807);
nor U14984 (N_14984,N_9209,N_8249);
nor U14985 (N_14985,N_5436,N_5460);
nand U14986 (N_14986,N_8659,N_5278);
nor U14987 (N_14987,N_8249,N_8429);
or U14988 (N_14988,N_9822,N_7580);
nor U14989 (N_14989,N_7731,N_9528);
nor U14990 (N_14990,N_6539,N_6717);
or U14991 (N_14991,N_6631,N_8590);
nand U14992 (N_14992,N_5239,N_5310);
nand U14993 (N_14993,N_8314,N_7010);
or U14994 (N_14994,N_9488,N_6430);
xnor U14995 (N_14995,N_8900,N_8420);
and U14996 (N_14996,N_8132,N_5038);
xnor U14997 (N_14997,N_7034,N_9646);
nand U14998 (N_14998,N_5669,N_5349);
and U14999 (N_14999,N_6973,N_9486);
nand U15000 (N_15000,N_12709,N_13680);
and U15001 (N_15001,N_11483,N_14187);
nor U15002 (N_15002,N_10080,N_13936);
nor U15003 (N_15003,N_14411,N_14285);
xor U15004 (N_15004,N_13642,N_10854);
or U15005 (N_15005,N_12317,N_10083);
xor U15006 (N_15006,N_14425,N_10898);
xnor U15007 (N_15007,N_12755,N_12809);
or U15008 (N_15008,N_10991,N_12393);
xor U15009 (N_15009,N_10914,N_11889);
xor U15010 (N_15010,N_12209,N_10238);
and U15011 (N_15011,N_12097,N_10593);
or U15012 (N_15012,N_12252,N_10119);
nor U15013 (N_15013,N_14955,N_13119);
or U15014 (N_15014,N_12021,N_14517);
xor U15015 (N_15015,N_11529,N_13044);
and U15016 (N_15016,N_13113,N_14221);
or U15017 (N_15017,N_10353,N_10101);
or U15018 (N_15018,N_14191,N_13894);
nand U15019 (N_15019,N_13814,N_11391);
nor U15020 (N_15020,N_11928,N_12150);
nor U15021 (N_15021,N_10496,N_11805);
nor U15022 (N_15022,N_14541,N_14011);
nand U15023 (N_15023,N_12592,N_14487);
xor U15024 (N_15024,N_11411,N_13861);
nand U15025 (N_15025,N_14749,N_14850);
nand U15026 (N_15026,N_13563,N_11108);
nand U15027 (N_15027,N_11793,N_12259);
or U15028 (N_15028,N_12061,N_13610);
or U15029 (N_15029,N_12300,N_13973);
xnor U15030 (N_15030,N_12348,N_11751);
nand U15031 (N_15031,N_12245,N_13182);
or U15032 (N_15032,N_11451,N_13896);
nor U15033 (N_15033,N_12807,N_11518);
xor U15034 (N_15034,N_12375,N_12437);
nand U15035 (N_15035,N_13067,N_13766);
nor U15036 (N_15036,N_11818,N_10055);
xor U15037 (N_15037,N_10942,N_13104);
xnor U15038 (N_15038,N_11342,N_12666);
nand U15039 (N_15039,N_10528,N_11557);
nand U15040 (N_15040,N_14396,N_10604);
or U15041 (N_15041,N_13638,N_14438);
xnor U15042 (N_15042,N_10035,N_10014);
nor U15043 (N_15043,N_13391,N_12497);
and U15044 (N_15044,N_14325,N_11145);
nor U15045 (N_15045,N_12521,N_11612);
xor U15046 (N_15046,N_11533,N_13477);
nor U15047 (N_15047,N_11707,N_14959);
nor U15048 (N_15048,N_11063,N_12232);
nand U15049 (N_15049,N_12257,N_11511);
nand U15050 (N_15050,N_13041,N_14660);
xnor U15051 (N_15051,N_13575,N_12525);
and U15052 (N_15052,N_10142,N_10387);
or U15053 (N_15053,N_11115,N_10943);
or U15054 (N_15054,N_14873,N_12985);
and U15055 (N_15055,N_11492,N_14563);
xnor U15056 (N_15056,N_13707,N_10997);
and U15057 (N_15057,N_11417,N_14963);
and U15058 (N_15058,N_13652,N_10424);
nor U15059 (N_15059,N_11566,N_12597);
or U15060 (N_15060,N_11610,N_11201);
nand U15061 (N_15061,N_12674,N_13442);
nand U15062 (N_15062,N_14891,N_12760);
or U15063 (N_15063,N_14585,N_10252);
and U15064 (N_15064,N_10558,N_10766);
nand U15065 (N_15065,N_10639,N_14040);
nand U15066 (N_15066,N_11348,N_14962);
xor U15067 (N_15067,N_14856,N_10621);
nand U15068 (N_15068,N_14257,N_11459);
and U15069 (N_15069,N_12585,N_11957);
xor U15070 (N_15070,N_14395,N_12901);
xor U15071 (N_15071,N_14874,N_14414);
nor U15072 (N_15072,N_12098,N_11546);
and U15073 (N_15073,N_10115,N_13753);
xor U15074 (N_15074,N_10598,N_13636);
and U15075 (N_15075,N_13414,N_13979);
and U15076 (N_15076,N_13154,N_14900);
and U15077 (N_15077,N_13915,N_10715);
nand U15078 (N_15078,N_10732,N_10539);
xnor U15079 (N_15079,N_13673,N_14499);
nor U15080 (N_15080,N_11318,N_14201);
nand U15081 (N_15081,N_12382,N_11992);
or U15082 (N_15082,N_12189,N_10156);
and U15083 (N_15083,N_14952,N_10931);
xnor U15084 (N_15084,N_13721,N_11346);
and U15085 (N_15085,N_11013,N_11171);
nor U15086 (N_15086,N_14837,N_11895);
nor U15087 (N_15087,N_10106,N_11905);
nand U15088 (N_15088,N_12886,N_10426);
or U15089 (N_15089,N_13746,N_10999);
nand U15090 (N_15090,N_14810,N_11690);
nand U15091 (N_15091,N_11917,N_12899);
or U15092 (N_15092,N_13165,N_12840);
nand U15093 (N_15093,N_11066,N_14078);
xnor U15094 (N_15094,N_10792,N_10546);
and U15095 (N_15095,N_11271,N_10367);
and U15096 (N_15096,N_14394,N_10913);
or U15097 (N_15097,N_14491,N_12333);
or U15098 (N_15098,N_12904,N_13460);
or U15099 (N_15099,N_10578,N_12212);
nand U15100 (N_15100,N_10004,N_11971);
xnor U15101 (N_15101,N_14882,N_12764);
nand U15102 (N_15102,N_12472,N_14233);
and U15103 (N_15103,N_14675,N_10308);
or U15104 (N_15104,N_14186,N_12279);
nand U15105 (N_15105,N_10318,N_11980);
nand U15106 (N_15106,N_10232,N_13978);
or U15107 (N_15107,N_11939,N_10215);
nand U15108 (N_15108,N_13306,N_11831);
xor U15109 (N_15109,N_11230,N_14919);
nand U15110 (N_15110,N_14113,N_10489);
and U15111 (N_15111,N_14562,N_11626);
nor U15112 (N_15112,N_10276,N_14474);
nand U15113 (N_15113,N_12483,N_13678);
nand U15114 (N_15114,N_11532,N_10372);
nor U15115 (N_15115,N_12862,N_13988);
nor U15116 (N_15116,N_13102,N_12128);
or U15117 (N_15117,N_11363,N_11096);
xnor U15118 (N_15118,N_11400,N_13161);
nand U15119 (N_15119,N_11296,N_14983);
and U15120 (N_15120,N_14840,N_10843);
or U15121 (N_15121,N_11328,N_11397);
or U15122 (N_15122,N_14447,N_11899);
or U15123 (N_15123,N_10319,N_12532);
and U15124 (N_15124,N_14575,N_11195);
or U15125 (N_15125,N_13732,N_12767);
nor U15126 (N_15126,N_10587,N_12707);
nand U15127 (N_15127,N_11186,N_13186);
and U15128 (N_15128,N_14182,N_13074);
nor U15129 (N_15129,N_13889,N_11068);
nand U15130 (N_15130,N_14321,N_11906);
nor U15131 (N_15131,N_10124,N_11437);
xnor U15132 (N_15132,N_11945,N_14344);
or U15133 (N_15133,N_14202,N_12491);
xor U15134 (N_15134,N_10342,N_13334);
nor U15135 (N_15135,N_14366,N_14542);
and U15136 (N_15136,N_10916,N_14076);
xnor U15137 (N_15137,N_13938,N_11742);
nor U15138 (N_15138,N_12339,N_12648);
xor U15139 (N_15139,N_10311,N_14164);
or U15140 (N_15140,N_11754,N_12217);
nor U15141 (N_15141,N_11938,N_13534);
or U15142 (N_15142,N_12170,N_12253);
nand U15143 (N_15143,N_13819,N_14323);
xnor U15144 (N_15144,N_14105,N_10956);
or U15145 (N_15145,N_10248,N_10551);
or U15146 (N_15146,N_13543,N_13954);
xnor U15147 (N_15147,N_11460,N_11026);
nand U15148 (N_15148,N_10389,N_11470);
or U15149 (N_15149,N_11501,N_11399);
nand U15150 (N_15150,N_11785,N_12636);
nor U15151 (N_15151,N_10378,N_11517);
or U15152 (N_15152,N_14420,N_14427);
xnor U15153 (N_15153,N_13462,N_13629);
and U15154 (N_15154,N_12896,N_10657);
nand U15155 (N_15155,N_10325,N_12396);
nor U15156 (N_15156,N_13576,N_13810);
nor U15157 (N_15157,N_10563,N_14482);
xnor U15158 (N_15158,N_12271,N_14039);
and U15159 (N_15159,N_11314,N_10729);
or U15160 (N_15160,N_13676,N_14915);
nand U15161 (N_15161,N_10859,N_12032);
or U15162 (N_15162,N_14974,N_14489);
nand U15163 (N_15163,N_13091,N_14507);
and U15164 (N_15164,N_11668,N_13635);
nand U15165 (N_15165,N_11847,N_13445);
xnor U15166 (N_15166,N_14304,N_11119);
and U15167 (N_15167,N_13371,N_13960);
and U15168 (N_15168,N_10240,N_13363);
xor U15169 (N_15169,N_12815,N_12584);
nor U15170 (N_15170,N_14203,N_12751);
nand U15171 (N_15171,N_13572,N_11011);
nand U15172 (N_15172,N_14716,N_11367);
xor U15173 (N_15173,N_13486,N_13424);
xor U15174 (N_15174,N_10706,N_14155);
and U15175 (N_15175,N_14197,N_14393);
nand U15176 (N_15176,N_12605,N_12941);
nor U15177 (N_15177,N_13398,N_10397);
or U15178 (N_15178,N_10036,N_14049);
or U15179 (N_15179,N_12559,N_11739);
or U15180 (N_15180,N_12802,N_14226);
and U15181 (N_15181,N_10521,N_13305);
xor U15182 (N_15182,N_10716,N_10767);
xnor U15183 (N_15183,N_13167,N_13244);
or U15184 (N_15184,N_12040,N_10815);
xnor U15185 (N_15185,N_12052,N_11476);
xnor U15186 (N_15186,N_10335,N_14118);
nor U15187 (N_15187,N_14373,N_14050);
xnor U15188 (N_15188,N_12177,N_14583);
and U15189 (N_15189,N_10865,N_14827);
nor U15190 (N_15190,N_11364,N_10011);
or U15191 (N_15191,N_10282,N_12413);
and U15192 (N_15192,N_13911,N_13366);
xor U15193 (N_15193,N_13408,N_14194);
nand U15194 (N_15194,N_13929,N_11819);
or U15195 (N_15195,N_13361,N_12397);
or U15196 (N_15196,N_13857,N_10057);
xor U15197 (N_15197,N_11773,N_11269);
xor U15198 (N_15198,N_12745,N_11242);
and U15199 (N_15199,N_10993,N_12550);
nand U15200 (N_15200,N_14645,N_13280);
or U15201 (N_15201,N_12658,N_14608);
nor U15202 (N_15202,N_13079,N_14467);
nor U15203 (N_15203,N_12590,N_11873);
and U15204 (N_15204,N_12384,N_13177);
xnor U15205 (N_15205,N_11383,N_14656);
or U15206 (N_15206,N_13441,N_12882);
and U15207 (N_15207,N_14894,N_10233);
or U15208 (N_15208,N_11140,N_12220);
and U15209 (N_15209,N_13518,N_11556);
xor U15210 (N_15210,N_13139,N_11260);
and U15211 (N_15211,N_11658,N_14719);
nor U15212 (N_15212,N_10484,N_13666);
xor U15213 (N_15213,N_14041,N_10464);
nand U15214 (N_15214,N_12965,N_13654);
xnor U15215 (N_15215,N_10110,N_10269);
and U15216 (N_15216,N_14433,N_14907);
or U15217 (N_15217,N_13722,N_13415);
and U15218 (N_15218,N_12304,N_10681);
xor U15219 (N_15219,N_13701,N_13842);
xor U15220 (N_15220,N_10895,N_11516);
nor U15221 (N_15221,N_10994,N_11620);
nor U15222 (N_15222,N_11777,N_12612);
nor U15223 (N_15223,N_10901,N_14858);
nand U15224 (N_15224,N_14851,N_13342);
and U15225 (N_15225,N_13005,N_10794);
xor U15226 (N_15226,N_14984,N_13568);
nand U15227 (N_15227,N_11832,N_13376);
xnor U15228 (N_15228,N_12889,N_14215);
and U15229 (N_15229,N_11904,N_14609);
xnor U15230 (N_15230,N_13796,N_14966);
xor U15231 (N_15231,N_11169,N_10358);
and U15232 (N_15232,N_12318,N_14244);
nand U15233 (N_15233,N_13852,N_14413);
or U15234 (N_15234,N_14745,N_14695);
nand U15235 (N_15235,N_14193,N_11107);
xor U15236 (N_15236,N_10870,N_14811);
or U15237 (N_15237,N_13550,N_11490);
and U15238 (N_15238,N_14328,N_13142);
xnor U15239 (N_15239,N_10301,N_13172);
xor U15240 (N_15240,N_11049,N_12763);
nand U15241 (N_15241,N_13492,N_13858);
or U15242 (N_15242,N_13937,N_11868);
nand U15243 (N_15243,N_11596,N_11875);
nor U15244 (N_15244,N_11276,N_14409);
nand U15245 (N_15245,N_11023,N_13608);
nand U15246 (N_15246,N_12439,N_14713);
nand U15247 (N_15247,N_14574,N_13625);
and U15248 (N_15248,N_11554,N_12218);
or U15249 (N_15249,N_11019,N_11046);
nand U15250 (N_15250,N_13360,N_14453);
nor U15251 (N_15251,N_13515,N_13659);
nor U15252 (N_15252,N_11942,N_11192);
nor U15253 (N_15253,N_13147,N_11376);
or U15254 (N_15254,N_13045,N_13193);
and U15255 (N_15255,N_10965,N_14623);
nand U15256 (N_15256,N_14890,N_12961);
xnor U15257 (N_15257,N_12544,N_10869);
or U15258 (N_15258,N_11993,N_11016);
nand U15259 (N_15259,N_14122,N_11129);
and U15260 (N_15260,N_10940,N_10316);
or U15261 (N_15261,N_12208,N_11666);
nand U15262 (N_15262,N_11159,N_14119);
or U15263 (N_15263,N_10400,N_12919);
nand U15264 (N_15264,N_13315,N_14587);
xnor U15265 (N_15265,N_11587,N_13781);
and U15266 (N_15266,N_10212,N_12219);
xnor U15267 (N_15267,N_13418,N_13088);
xor U15268 (N_15268,N_14147,N_13548);
nand U15269 (N_15269,N_12131,N_12710);
nand U15270 (N_15270,N_11193,N_11547);
nand U15271 (N_15271,N_13591,N_14471);
and U15272 (N_15272,N_14722,N_12504);
nand U15273 (N_15273,N_13019,N_12376);
xnor U15274 (N_15274,N_12204,N_12969);
nor U15275 (N_15275,N_14917,N_12461);
and U15276 (N_15276,N_11443,N_11814);
xnor U15277 (N_15277,N_13913,N_14756);
nand U15278 (N_15278,N_12383,N_11220);
and U15279 (N_15279,N_13413,N_14978);
and U15280 (N_15280,N_11584,N_14841);
nor U15281 (N_15281,N_14450,N_11007);
nor U15282 (N_15282,N_12144,N_14376);
or U15283 (N_15283,N_12067,N_10637);
or U15284 (N_15284,N_14343,N_13435);
and U15285 (N_15285,N_14712,N_11680);
nor U15286 (N_15286,N_12990,N_12546);
nand U15287 (N_15287,N_14140,N_10608);
nor U15288 (N_15288,N_10281,N_11360);
or U15289 (N_15289,N_10343,N_12020);
or U15290 (N_15290,N_14691,N_13597);
and U15291 (N_15291,N_12782,N_13864);
nor U15292 (N_15292,N_11252,N_10878);
nor U15293 (N_15293,N_10157,N_11325);
or U15294 (N_15294,N_14292,N_10911);
nor U15295 (N_15295,N_13833,N_13836);
nor U15296 (N_15296,N_14424,N_14560);
nand U15297 (N_15297,N_11249,N_11368);
nor U15298 (N_15298,N_12870,N_12018);
nand U15299 (N_15299,N_13250,N_12885);
xnor U15300 (N_15300,N_13918,N_12008);
and U15301 (N_15301,N_10191,N_13464);
or U15302 (N_15302,N_14115,N_13326);
xor U15303 (N_15303,N_14198,N_10884);
xor U15304 (N_15304,N_13290,N_13195);
nand U15305 (N_15305,N_12999,N_10957);
nor U15306 (N_15306,N_11564,N_13544);
or U15307 (N_15307,N_12288,N_11381);
nand U15308 (N_15308,N_12856,N_11614);
and U15309 (N_15309,N_13373,N_12494);
and U15310 (N_15310,N_12028,N_12010);
xnor U15311 (N_15311,N_10763,N_11839);
nor U15312 (N_15312,N_12250,N_12200);
or U15313 (N_15313,N_12599,N_11312);
xor U15314 (N_15314,N_10505,N_12153);
and U15315 (N_15315,N_14108,N_11306);
nand U15316 (N_15316,N_11983,N_10032);
and U15317 (N_15317,N_14689,N_10396);
and U15318 (N_15318,N_12869,N_12754);
nor U15319 (N_15319,N_13344,N_12110);
xor U15320 (N_15320,N_10034,N_13633);
nand U15321 (N_15321,N_12068,N_12959);
nor U15322 (N_15322,N_11461,N_11864);
and U15323 (N_15323,N_12613,N_10431);
nand U15324 (N_15324,N_10229,N_13689);
nand U15325 (N_15325,N_12244,N_14670);
nor U15326 (N_15326,N_11613,N_10892);
nor U15327 (N_15327,N_11630,N_11560);
or U15328 (N_15328,N_14071,N_12326);
or U15329 (N_15329,N_10117,N_11469);
nor U15330 (N_15330,N_14999,N_13377);
xnor U15331 (N_15331,N_11734,N_10885);
or U15332 (N_15332,N_10172,N_12074);
or U15333 (N_15333,N_11317,N_13825);
nand U15334 (N_15334,N_11618,N_11057);
and U15335 (N_15335,N_13856,N_14853);
nor U15336 (N_15336,N_14473,N_13510);
xnor U15337 (N_15337,N_10019,N_10167);
and U15338 (N_15338,N_10073,N_14755);
xnor U15339 (N_15339,N_14596,N_12643);
nand U15340 (N_15340,N_12179,N_11663);
or U15341 (N_15341,N_11062,N_13974);
nor U15342 (N_15342,N_11624,N_10921);
nand U15343 (N_15343,N_13577,N_14975);
xor U15344 (N_15344,N_11361,N_12617);
xor U15345 (N_15345,N_10201,N_11878);
nand U15346 (N_15346,N_14251,N_14145);
nand U15347 (N_15347,N_13688,N_14143);
nor U15348 (N_15348,N_11806,N_14322);
nand U15349 (N_15349,N_12495,N_13010);
nand U15350 (N_15350,N_11721,N_12205);
or U15351 (N_15351,N_14238,N_10460);
xnor U15352 (N_15352,N_14653,N_10473);
nor U15353 (N_15353,N_13089,N_12265);
nor U15354 (N_15354,N_11728,N_14248);
nand U15355 (N_15355,N_10404,N_12829);
and U15356 (N_15356,N_12766,N_14058);
nand U15357 (N_15357,N_12139,N_11148);
nand U15358 (N_15358,N_11711,N_11081);
nor U15359 (N_15359,N_14782,N_14472);
xnor U15360 (N_15360,N_10278,N_13981);
nand U15361 (N_15361,N_12850,N_12680);
and U15362 (N_15362,N_11432,N_12411);
nand U15363 (N_15363,N_14311,N_13444);
or U15364 (N_15364,N_14214,N_11857);
nor U15365 (N_15365,N_10907,N_14514);
or U15366 (N_15366,N_13349,N_13209);
and U15367 (N_15367,N_13097,N_14175);
or U15368 (N_15368,N_14730,N_10809);
nor U15369 (N_15369,N_13788,N_10193);
xor U15370 (N_15370,N_11452,N_10271);
and U15371 (N_15371,N_12556,N_14402);
and U15372 (N_15372,N_13994,N_10540);
and U15373 (N_15373,N_10824,N_11619);
nand U15374 (N_15374,N_11415,N_14530);
nand U15375 (N_15375,N_11485,N_12852);
and U15376 (N_15376,N_10206,N_13986);
nor U15377 (N_15377,N_13776,N_10091);
nand U15378 (N_15378,N_11930,N_10437);
nand U15379 (N_15379,N_14668,N_10021);
and U15380 (N_15380,N_11332,N_11822);
nand U15381 (N_15381,N_14786,N_13525);
xor U15382 (N_15382,N_13712,N_11695);
nor U15383 (N_15383,N_11457,N_10723);
or U15384 (N_15384,N_12423,N_10568);
nor U15385 (N_15385,N_10453,N_14696);
nand U15386 (N_15386,N_12444,N_10696);
or U15387 (N_15387,N_11055,N_14877);
and U15388 (N_15388,N_12857,N_10970);
or U15389 (N_15389,N_10985,N_14488);
or U15390 (N_15390,N_10700,N_10938);
and U15391 (N_15391,N_10328,N_13860);
xnor U15392 (N_15392,N_13479,N_12635);
xor U15393 (N_15393,N_11682,N_12462);
and U15394 (N_15394,N_10982,N_13109);
nand U15395 (N_15395,N_10192,N_12490);
or U15396 (N_15396,N_14911,N_11984);
xnor U15397 (N_15397,N_10651,N_13924);
and U15398 (N_15398,N_13192,N_10564);
nand U15399 (N_15399,N_12112,N_12484);
nand U15400 (N_15400,N_13768,N_12343);
or U15401 (N_15401,N_12569,N_10631);
or U15402 (N_15402,N_11125,N_11319);
nor U15403 (N_15403,N_10031,N_11309);
nand U15404 (N_15404,N_12792,N_14511);
xor U15405 (N_15405,N_14815,N_11716);
and U15406 (N_15406,N_12331,N_11416);
or U15407 (N_15407,N_12656,N_10310);
nor U15408 (N_15408,N_10586,N_14616);
xnor U15409 (N_15409,N_12352,N_13411);
nor U15410 (N_15410,N_11410,N_13669);
and U15411 (N_15411,N_14602,N_10623);
nand U15412 (N_15412,N_12302,N_14531);
nand U15413 (N_15413,N_11392,N_13660);
nor U15414 (N_15414,N_12264,N_11288);
and U15415 (N_15415,N_10990,N_13145);
nand U15416 (N_15416,N_13399,N_14033);
xor U15417 (N_15417,N_11586,N_11458);
and U15418 (N_15418,N_12781,N_13352);
nor U15419 (N_15419,N_14318,N_12420);
nand U15420 (N_15420,N_12665,N_10573);
xor U15421 (N_15421,N_12795,N_14951);
and U15422 (N_15422,N_12513,N_11580);
nand U15423 (N_15423,N_13813,N_12626);
nand U15424 (N_15424,N_13007,N_11241);
and U15425 (N_15425,N_14205,N_14947);
xnor U15426 (N_15426,N_14230,N_13811);
and U15427 (N_15427,N_10027,N_13599);
or U15428 (N_15428,N_13595,N_11528);
or U15429 (N_15429,N_12696,N_11499);
nor U15430 (N_15430,N_11922,N_11217);
and U15431 (N_15431,N_10002,N_13557);
and U15432 (N_15432,N_13033,N_14766);
or U15433 (N_15433,N_14522,N_14348);
nor U15434 (N_15434,N_13950,N_10214);
xnor U15435 (N_15435,N_12142,N_11093);
and U15436 (N_15436,N_11446,N_14994);
or U15437 (N_15437,N_13370,N_10811);
nor U15438 (N_15438,N_14943,N_10407);
xnor U15439 (N_15439,N_14445,N_13272);
or U15440 (N_15440,N_14658,N_10509);
nor U15441 (N_15441,N_12037,N_13545);
or U15442 (N_15442,N_12402,N_13153);
nor U15443 (N_15443,N_14229,N_10354);
xor U15444 (N_15444,N_10769,N_10111);
nor U15445 (N_15445,N_11261,N_12057);
nand U15446 (N_15446,N_12310,N_10144);
and U15447 (N_15447,N_14030,N_13395);
xnor U15448 (N_15448,N_14377,N_13631);
xnor U15449 (N_15449,N_10848,N_10090);
or U15450 (N_15450,N_14448,N_11280);
and U15451 (N_15451,N_13928,N_13345);
nand U15452 (N_15452,N_12733,N_11522);
and U15453 (N_15453,N_10636,N_13696);
xnor U15454 (N_15454,N_11048,N_10054);
xnor U15455 (N_15455,N_14480,N_14498);
nand U15456 (N_15456,N_13314,N_11588);
xor U15457 (N_15457,N_11717,N_11943);
and U15458 (N_15458,N_11335,N_11882);
nand U15459 (N_15459,N_12534,N_12711);
or U15460 (N_15460,N_13336,N_14000);
or U15461 (N_15461,N_11884,N_14410);
nand U15462 (N_15462,N_10145,N_10261);
and U15463 (N_15463,N_10690,N_14778);
or U15464 (N_15464,N_12202,N_14080);
nor U15465 (N_15465,N_14572,N_10567);
xor U15466 (N_15466,N_13751,N_13920);
xnor U15467 (N_15467,N_14612,N_12638);
and U15468 (N_15468,N_10390,N_13419);
or U15469 (N_15469,N_10391,N_11106);
and U15470 (N_15470,N_11000,N_12313);
or U15471 (N_15471,N_11462,N_13100);
nand U15472 (N_15472,N_13767,N_10522);
xor U15473 (N_15473,N_13425,N_14967);
nand U15474 (N_15474,N_13728,N_12778);
nor U15475 (N_15475,N_12868,N_14478);
xnor U15476 (N_15476,N_12269,N_13485);
or U15477 (N_15477,N_11975,N_12194);
nor U15478 (N_15478,N_13521,N_14624);
or U15479 (N_15479,N_11480,N_14534);
xnor U15480 (N_15480,N_10043,N_11341);
and U15481 (N_15481,N_13480,N_14854);
nor U15482 (N_15482,N_10996,N_13573);
xnor U15483 (N_15483,N_14960,N_11635);
nand U15484 (N_15484,N_13733,N_10543);
and U15485 (N_15485,N_13129,N_10712);
or U15486 (N_15486,N_11272,N_10738);
xnor U15487 (N_15487,N_12718,N_10289);
and U15488 (N_15488,N_14546,N_14405);
and U15489 (N_15489,N_12842,N_11725);
and U15490 (N_15490,N_10719,N_12602);
or U15491 (N_15491,N_12299,N_10702);
or U15492 (N_15492,N_13199,N_10000);
xor U15493 (N_15493,N_11175,N_12233);
or U15494 (N_15494,N_12828,N_12975);
and U15495 (N_15495,N_10658,N_12373);
nor U15496 (N_15496,N_12404,N_11097);
xnor U15497 (N_15497,N_13762,N_11911);
nand U15498 (N_15498,N_10634,N_13252);
xor U15499 (N_15499,N_12188,N_11827);
or U15500 (N_15500,N_13763,N_10989);
xnor U15501 (N_15501,N_13212,N_11653);
nor U15502 (N_15502,N_13423,N_11498);
xor U15503 (N_15503,N_11578,N_10136);
or U15504 (N_15504,N_13771,N_10671);
xor U15505 (N_15505,N_12837,N_14104);
or U15506 (N_15506,N_12511,N_10655);
or U15507 (N_15507,N_11503,N_14737);
nor U15508 (N_15508,N_11014,N_11550);
and U15509 (N_15509,N_10065,N_14089);
or U15510 (N_15510,N_13012,N_10129);
nand U15511 (N_15511,N_14986,N_12516);
nand U15512 (N_15512,N_10958,N_11623);
nand U15513 (N_15513,N_11599,N_11041);
and U15514 (N_15514,N_11138,N_14267);
or U15515 (N_15515,N_12447,N_11648);
xor U15516 (N_15516,N_13229,N_12762);
and U15517 (N_15517,N_13821,N_13261);
xnor U15518 (N_15518,N_13009,N_14195);
nand U15519 (N_15519,N_12742,N_12957);
or U15520 (N_15520,N_14176,N_13906);
nand U15521 (N_15521,N_14264,N_11797);
nor U15522 (N_15522,N_14048,N_10613);
nor U15523 (N_15523,N_12818,N_14687);
nand U15524 (N_15524,N_10647,N_11820);
and U15525 (N_15525,N_12640,N_13245);
xnor U15526 (N_15526,N_14893,N_11852);
nand U15527 (N_15527,N_11086,N_11173);
xor U15528 (N_15528,N_10359,N_13222);
and U15529 (N_15529,N_12800,N_10694);
and U15530 (N_15530,N_14772,N_14086);
xnor U15531 (N_15531,N_13606,N_11172);
or U15532 (N_15532,N_10932,N_12621);
and U15533 (N_15533,N_11909,N_14601);
or U15534 (N_15534,N_14110,N_12314);
and U15535 (N_15535,N_10751,N_11888);
nor U15536 (N_15536,N_14746,N_11702);
nand U15537 (N_15537,N_10360,N_10590);
nand U15538 (N_15538,N_12560,N_13122);
or U15539 (N_15539,N_11300,N_12858);
and U15540 (N_15540,N_10306,N_12705);
and U15541 (N_15541,N_11244,N_12216);
nand U15542 (N_15542,N_14533,N_10605);
and U15543 (N_15543,N_14726,N_14421);
xor U15544 (N_15544,N_14934,N_12044);
xnor U15545 (N_15545,N_11150,N_12871);
xnor U15546 (N_15546,N_10695,N_13824);
nand U15547 (N_15547,N_11127,N_10917);
xnor U15548 (N_15548,N_10333,N_14760);
nand U15549 (N_15549,N_11549,N_10779);
xnor U15550 (N_15550,N_10363,N_14068);
and U15551 (N_15551,N_10494,N_12429);
or U15552 (N_15552,N_11641,N_11429);
or U15553 (N_15553,N_12111,N_13134);
nor U15554 (N_15554,N_10374,N_11935);
xor U15555 (N_15555,N_14734,N_14092);
and U15556 (N_15556,N_12251,N_10255);
xnor U15557 (N_15557,N_14005,N_10733);
and U15558 (N_15558,N_10980,N_10329);
nand U15559 (N_15559,N_10234,N_11430);
nand U15560 (N_15560,N_10210,N_12174);
nor U15561 (N_15561,N_14682,N_14382);
or U15562 (N_15562,N_12756,N_10530);
or U15563 (N_15563,N_10152,N_13389);
nand U15564 (N_15564,N_10197,N_10915);
and U15565 (N_15565,N_11199,N_10490);
or U15566 (N_15566,N_12893,N_13589);
and U15567 (N_15567,N_12369,N_12798);
or U15568 (N_15568,N_10195,N_10768);
or U15569 (N_15569,N_13524,N_13698);
and U15570 (N_15570,N_10813,N_12723);
nor U15571 (N_15571,N_13082,N_12035);
or U15572 (N_15572,N_10170,N_12457);
or U15573 (N_15573,N_12670,N_12775);
nand U15574 (N_15574,N_11440,N_12254);
nor U15575 (N_15575,N_13761,N_13432);
xnor U15576 (N_15576,N_11779,N_14385);
and U15577 (N_15577,N_12971,N_14392);
nand U15578 (N_15578,N_13919,N_11575);
nand U15579 (N_15579,N_13709,N_12996);
nor U15580 (N_15580,N_14277,N_10442);
or U15581 (N_15581,N_14234,N_13130);
and U15582 (N_15582,N_13469,N_12844);
or U15583 (N_15583,N_11104,N_11606);
nor U15584 (N_15584,N_13816,N_13394);
xnor U15585 (N_15585,N_11025,N_12133);
nor U15586 (N_15586,N_10114,N_10075);
or U15587 (N_15587,N_13171,N_11365);
and U15588 (N_15588,N_13191,N_12738);
xor U15589 (N_15589,N_11694,N_10393);
nor U15590 (N_15590,N_10737,N_14996);
and U15591 (N_15591,N_13687,N_10939);
nand U15592 (N_15592,N_13230,N_13693);
nand U15593 (N_15593,N_13992,N_14503);
or U15594 (N_15594,N_12262,N_12826);
xor U15595 (N_15595,N_10469,N_11863);
xnor U15596 (N_15596,N_11593,N_13381);
nor U15597 (N_15597,N_10532,N_12529);
and U15598 (N_15598,N_13844,N_13308);
and U15599 (N_15599,N_10285,N_11530);
and U15600 (N_15600,N_12861,N_13076);
and U15601 (N_15601,N_11128,N_14003);
and U15602 (N_15602,N_10413,N_10417);
nor U15603 (N_15603,N_10334,N_13173);
and U15604 (N_15604,N_13253,N_13708);
and U15605 (N_15605,N_11581,N_14153);
and U15606 (N_15606,N_13329,N_12753);
nor U15607 (N_15607,N_10904,N_14626);
xnor U15608 (N_15608,N_13710,N_10514);
and U15609 (N_15609,N_12647,N_11880);
or U15610 (N_15610,N_12692,N_10243);
xnor U15611 (N_15611,N_13517,N_10804);
xor U15612 (N_15612,N_13787,N_12810);
and U15613 (N_15613,N_13714,N_14685);
xnor U15614 (N_15614,N_11114,N_11423);
xnor U15615 (N_15615,N_12972,N_11126);
xnor U15616 (N_15616,N_11629,N_13065);
xor U15617 (N_15617,N_10614,N_11585);
nor U15618 (N_15618,N_12672,N_14426);
and U15619 (N_15619,N_14428,N_12575);
nand U15620 (N_15620,N_12874,N_12943);
and U15621 (N_15621,N_12046,N_14881);
nor U15622 (N_15622,N_10100,N_14942);
and U15623 (N_15623,N_12163,N_12240);
xor U15624 (N_15624,N_12860,N_13406);
nand U15625 (N_15625,N_11589,N_12747);
nor U15626 (N_15626,N_11170,N_10659);
nand U15627 (N_15627,N_12684,N_12566);
and U15628 (N_15628,N_12679,N_14116);
nand U15629 (N_15629,N_14898,N_12758);
nand U15630 (N_15630,N_10246,N_10887);
xnor U15631 (N_15631,N_13051,N_13022);
xor U15632 (N_15632,N_12506,N_13135);
or U15633 (N_15633,N_10787,N_10033);
nor U15634 (N_15634,N_11780,N_12549);
xnor U15635 (N_15635,N_12587,N_11123);
and U15636 (N_15636,N_14139,N_10883);
nor U15637 (N_15637,N_12031,N_14293);
and U15638 (N_15638,N_14946,N_14527);
or U15639 (N_15639,N_13546,N_14024);
and U15640 (N_15640,N_11932,N_10448);
xor U15641 (N_15641,N_14061,N_13302);
or U15642 (N_15642,N_14305,N_10178);
nand U15643 (N_15643,N_11187,N_11953);
and U15644 (N_15644,N_10734,N_13111);
or U15645 (N_15645,N_10436,N_14930);
nor U15646 (N_15646,N_12083,N_10153);
and U15647 (N_15647,N_12425,N_13584);
xnor U15648 (N_15648,N_14725,N_11386);
nand U15649 (N_15649,N_14804,N_11924);
nand U15650 (N_15650,N_13240,N_13726);
and U15651 (N_15651,N_10162,N_13313);
or U15652 (N_15652,N_12921,N_11937);
nor U15653 (N_15653,N_10833,N_10351);
xor U15654 (N_15654,N_12374,N_13723);
nor U15655 (N_15655,N_11036,N_12702);
or U15656 (N_15656,N_13217,N_12016);
nand U15657 (N_15657,N_13211,N_13180);
nand U15658 (N_15658,N_13379,N_12315);
and U15659 (N_15659,N_10365,N_14192);
xnor U15660 (N_15660,N_10796,N_10425);
xnor U15661 (N_15661,N_14905,N_11978);
or U15662 (N_15662,N_14029,N_12719);
nand U15663 (N_15663,N_12249,N_10948);
or U15664 (N_15664,N_13155,N_13574);
and U15665 (N_15665,N_14275,N_14055);
nor U15666 (N_15666,N_13739,N_14761);
nand U15667 (N_15667,N_14700,N_13392);
xnor U15668 (N_15668,N_14126,N_13047);
or U15669 (N_15669,N_10835,N_14240);
and U15670 (N_15670,N_10380,N_11266);
or U15671 (N_15671,N_12421,N_13291);
nor U15672 (N_15672,N_10429,N_10666);
nand U15673 (N_15673,N_10406,N_14916);
nor U15674 (N_15674,N_12392,N_10896);
and U15675 (N_15675,N_11676,N_12161);
or U15676 (N_15676,N_13020,N_11414);
nor U15677 (N_15677,N_14095,N_14286);
nand U15678 (N_15678,N_14013,N_13677);
nor U15679 (N_15679,N_12363,N_10474);
xnor U15680 (N_15680,N_13895,N_10332);
nand U15681 (N_15681,N_11277,N_13143);
nand U15682 (N_15682,N_14678,N_14308);
nand U15683 (N_15683,N_11234,N_10231);
or U15684 (N_15684,N_11344,N_14209);
nand U15685 (N_15685,N_13436,N_10776);
xnor U15686 (N_15686,N_12562,N_14995);
nand U15687 (N_15687,N_12958,N_12059);
nor U15688 (N_15688,N_12581,N_11157);
and U15689 (N_15689,N_11667,N_13138);
nand U15690 (N_15690,N_12750,N_14625);
nor U15691 (N_15691,N_11426,N_12668);
nand U15692 (N_15692,N_13283,N_12694);
nor U15693 (N_15693,N_10998,N_12281);
nand U15694 (N_15694,N_13164,N_13468);
xnor U15695 (N_15695,N_14389,N_12501);
and U15696 (N_15696,N_13341,N_14628);
nand U15697 (N_15697,N_11849,N_10973);
or U15698 (N_15698,N_11855,N_10542);
and U15699 (N_15699,N_12002,N_11539);
and U15700 (N_15700,N_12100,N_11508);
nor U15701 (N_15701,N_11685,N_12607);
nand U15702 (N_15702,N_13892,N_14157);
or U15703 (N_15703,N_10745,N_10962);
and U15704 (N_15704,N_12618,N_12805);
nand U15705 (N_15705,N_12428,N_12833);
nand U15706 (N_15706,N_14066,N_11449);
or U15707 (N_15707,N_13133,N_10402);
nor U15708 (N_15708,N_13001,N_13736);
nor U15709 (N_15709,N_11401,N_12542);
and U15710 (N_15710,N_11946,N_14903);
xnor U15711 (N_15711,N_14582,N_13704);
nor U15712 (N_15712,N_12596,N_13472);
xnor U15713 (N_15713,N_13927,N_12897);
nand U15714 (N_15714,N_12731,N_14159);
nand U15715 (N_15715,N_14836,N_14440);
nand U15716 (N_15716,N_13359,N_13949);
or U15717 (N_15717,N_10561,N_10290);
nor U15718 (N_15718,N_12606,N_10772);
and U15719 (N_15719,N_14298,N_14870);
xor U15720 (N_15720,N_10220,N_11670);
and U15721 (N_15721,N_10286,N_11047);
xnor U15722 (N_15722,N_13925,N_10668);
nand U15723 (N_15723,N_13241,N_13630);
and U15724 (N_15724,N_13806,N_10412);
nor U15725 (N_15725,N_11771,N_13731);
and U15726 (N_15726,N_10188,N_13433);
and U15727 (N_15727,N_10077,N_14958);
nor U15728 (N_15728,N_11017,N_12051);
xnor U15729 (N_15729,N_13096,N_11408);
nand U15730 (N_15730,N_10548,N_13874);
xnor U15731 (N_15731,N_14154,N_12888);
and U15732 (N_15732,N_12699,N_10735);
xnor U15733 (N_15733,N_12434,N_11279);
nor U15734 (N_15734,N_11582,N_11105);
xnor U15735 (N_15735,N_11526,N_14557);
or U15736 (N_15736,N_13879,N_13117);
or U15737 (N_15737,N_13935,N_13031);
or U15738 (N_15738,N_13637,N_10477);
xor U15739 (N_15739,N_12043,N_13105);
nor U15740 (N_15740,N_12214,N_10967);
or U15741 (N_15741,N_11069,N_13656);
nand U15742 (N_15742,N_12164,N_12371);
and U15743 (N_15743,N_10482,N_10919);
and U15744 (N_15744,N_13207,N_12450);
or U15745 (N_15745,N_12716,N_11848);
nand U15746 (N_15746,N_14538,N_10410);
nand U15747 (N_15747,N_13609,N_11072);
or U15748 (N_15748,N_14632,N_13756);
and U15749 (N_15749,N_14792,N_12713);
xor U15750 (N_15750,N_12268,N_12014);
or U15751 (N_15751,N_13318,N_12308);
and U15752 (N_15752,N_12728,N_12878);
and U15753 (N_15753,N_12048,N_13962);
and U15754 (N_15754,N_10687,N_14255);
nand U15755 (N_15755,N_11902,N_14295);
or U15756 (N_15756,N_11650,N_13064);
nand U15757 (N_15757,N_13646,N_12960);
nor U15758 (N_15758,N_13613,N_13279);
nand U15759 (N_15759,N_12688,N_11710);
nor U15760 (N_15760,N_14185,N_12305);
nor U15761 (N_15761,N_12737,N_12746);
and U15762 (N_15762,N_11345,N_10805);
and U15763 (N_15763,N_14988,N_12830);
or U15764 (N_15764,N_11375,N_12955);
and U15765 (N_15765,N_12739,N_14156);
nor U15766 (N_15766,N_10630,N_14398);
nand U15767 (N_15767,N_10762,N_12686);
or U15768 (N_15768,N_13116,N_10284);
nor U15769 (N_15769,N_12964,N_10827);
and U15770 (N_15770,N_14539,N_10314);
or U15771 (N_15771,N_13287,N_14969);
or U15772 (N_15772,N_13124,N_11372);
nand U15773 (N_15773,N_14589,N_13887);
nand U15774 (N_15774,N_12065,N_11183);
xor U15775 (N_15775,N_11552,N_11627);
or U15776 (N_15776,N_10799,N_13456);
xnor U15777 (N_15777,N_10293,N_14866);
nor U15778 (N_15778,N_10899,N_10633);
nand U15779 (N_15779,N_12910,N_11168);
nand U15780 (N_15780,N_12600,N_12221);
nor U15781 (N_15781,N_12956,N_13488);
and U15782 (N_15782,N_14351,N_12645);
nor U15783 (N_15783,N_13234,N_10463);
nand U15784 (N_15784,N_14739,N_10134);
or U15785 (N_15785,N_14509,N_11222);
and U15786 (N_15786,N_13274,N_14485);
nor U15787 (N_15787,N_13190,N_11862);
or U15788 (N_15788,N_10643,N_10455);
nand U15789 (N_15789,N_13541,N_10562);
nor U15790 (N_15790,N_12446,N_13720);
and U15791 (N_15791,N_10691,N_11144);
nand U15792 (N_15792,N_10099,N_11898);
or U15793 (N_15793,N_13567,N_10750);
or U15794 (N_15794,N_11789,N_14619);
nand U15795 (N_15795,N_14657,N_13554);
or U15796 (N_15796,N_14569,N_12017);
and U15797 (N_15797,N_12646,N_13547);
nand U15798 (N_15798,N_12106,N_14661);
nor U15799 (N_15799,N_11355,N_10791);
xor U15800 (N_15800,N_12611,N_11866);
nor U15801 (N_15801,N_12788,N_13218);
nand U15802 (N_15802,N_14412,N_11436);
and U15803 (N_15803,N_11027,N_13691);
or U15804 (N_15804,N_11211,N_10797);
and U15805 (N_15805,N_10265,N_13090);
or U15806 (N_15806,N_10495,N_12637);
or U15807 (N_15807,N_10493,N_14740);
nand U15808 (N_15808,N_12986,N_11512);
or U15809 (N_15809,N_14180,N_14641);
or U15810 (N_15810,N_13899,N_10368);
nor U15811 (N_15811,N_14060,N_11197);
or U15812 (N_15812,N_12385,N_13977);
xor U15813 (N_15813,N_11531,N_10150);
nand U15814 (N_15814,N_12512,N_12193);
nand U15815 (N_15815,N_10761,N_13325);
nand U15816 (N_15816,N_12845,N_11665);
xor U15817 (N_15817,N_14206,N_10470);
nor U15818 (N_15818,N_10467,N_14222);
xnor U15819 (N_15819,N_12741,N_10140);
xor U15820 (N_15820,N_10975,N_12055);
nand U15821 (N_15821,N_10018,N_11224);
xnor U15822 (N_15822,N_11358,N_14475);
or U15823 (N_15823,N_12379,N_14387);
nand U15824 (N_15824,N_11139,N_13422);
nand U15825 (N_15825,N_12791,N_10447);
nor U15826 (N_15826,N_11464,N_10009);
xor U15827 (N_15827,N_12145,N_10571);
nand U15828 (N_15828,N_13036,N_11625);
xor U15829 (N_15829,N_10610,N_10336);
or U15830 (N_15830,N_12045,N_11085);
nor U15831 (N_15831,N_12920,N_13686);
xnor U15832 (N_15832,N_10291,N_12578);
and U15833 (N_15833,N_11894,N_12812);
nor U15834 (N_15834,N_12071,N_14936);
nand U15835 (N_15835,N_13586,N_13428);
or U15836 (N_15836,N_10947,N_11094);
xor U15837 (N_15837,N_13410,N_11723);
or U15838 (N_15838,N_10008,N_14094);
xnor U15839 (N_15839,N_10337,N_13611);
and U15840 (N_15840,N_10686,N_12146);
nor U15841 (N_15841,N_13727,N_14697);
nor U15842 (N_15842,N_13148,N_13916);
xnor U15843 (N_15843,N_10267,N_14249);
nand U15844 (N_15844,N_14123,N_12477);
xor U15845 (N_15845,N_12287,N_14130);
nand U15846 (N_15846,N_10597,N_14524);
and U15847 (N_15847,N_10774,N_12238);
nor U15848 (N_15848,N_11854,N_13431);
nor U15849 (N_15849,N_14950,N_14004);
and U15850 (N_15850,N_13281,N_13848);
nand U15851 (N_15851,N_10222,N_12717);
or U15852 (N_15852,N_11311,N_13482);
nor U15853 (N_15853,N_11910,N_14120);
or U15854 (N_15854,N_13539,N_11239);
or U15855 (N_15855,N_14604,N_10462);
or U15856 (N_15856,N_14816,N_13474);
and U15857 (N_15857,N_11649,N_14436);
xnor U15858 (N_15858,N_12176,N_13466);
xor U15859 (N_15859,N_10208,N_13324);
nand U15860 (N_15860,N_11326,N_12915);
or U15861 (N_15861,N_13098,N_14314);
or U15862 (N_15862,N_10758,N_14785);
or U15863 (N_15863,N_11524,N_10127);
or U15864 (N_15864,N_13156,N_11605);
nand U15865 (N_15865,N_13989,N_10519);
nand U15866 (N_15866,N_11463,N_13043);
nor U15867 (N_15867,N_11302,N_10133);
nand U15868 (N_15868,N_10603,N_10247);
or U15869 (N_15869,N_12768,N_13968);
xnor U15870 (N_15870,N_13255,N_14860);
or U15871 (N_15871,N_13276,N_11726);
and U15872 (N_15872,N_12881,N_11800);
nand U15873 (N_15873,N_12681,N_12855);
nand U15874 (N_15874,N_13094,N_13522);
or U15875 (N_15875,N_14468,N_12316);
or U15876 (N_15876,N_13772,N_13667);
nand U15877 (N_15877,N_14458,N_11914);
or U15878 (N_15878,N_10341,N_14899);
and U15879 (N_15879,N_13463,N_11903);
xor U15880 (N_15880,N_14590,N_14225);
nor U15881 (N_15881,N_13914,N_11010);
xor U15882 (N_15882,N_13309,N_14466);
nand U15883 (N_15883,N_14158,N_12086);
and U15884 (N_15884,N_14603,N_11824);
xnor U15885 (N_15885,N_12949,N_14662);
xnor U15886 (N_15886,N_12030,N_14769);
and U15887 (N_15887,N_12604,N_14497);
or U15888 (N_15888,N_13888,N_12866);
and U15889 (N_15889,N_13719,N_14415);
nand U15890 (N_15890,N_13556,N_10771);
xor U15891 (N_15891,N_13817,N_14977);
and U15892 (N_15892,N_12565,N_10945);
nand U15893 (N_15893,N_12784,N_13828);
and U15894 (N_15894,N_11536,N_14709);
nor U15895 (N_15895,N_11194,N_11379);
nor U15896 (N_15896,N_14549,N_12357);
xnor U15897 (N_15897,N_14163,N_14565);
nand U15898 (N_15898,N_13459,N_10656);
xor U15899 (N_15899,N_14243,N_14883);
and U15900 (N_15900,N_12522,N_10632);
and U15901 (N_15901,N_14397,N_10619);
and U15902 (N_15902,N_13740,N_14272);
or U15903 (N_15903,N_11058,N_10912);
nand U15904 (N_15904,N_11374,N_10617);
or U15905 (N_15905,N_10299,N_11813);
nand U15906 (N_15906,N_13206,N_12586);
xor U15907 (N_15907,N_13627,N_14199);
or U15908 (N_15908,N_12474,N_11960);
nand U15909 (N_15909,N_14706,N_11558);
nand U15910 (N_15910,N_10795,N_13531);
and U15911 (N_15911,N_14954,N_11237);
xor U15912 (N_15912,N_10755,N_12589);
nand U15913 (N_15913,N_13598,N_13150);
and U15914 (N_15914,N_10478,N_14085);
or U15915 (N_15915,N_14738,N_10984);
and U15916 (N_15916,N_13396,N_10882);
xnor U15917 (N_15917,N_10064,N_11340);
nor U15918 (N_15918,N_12942,N_10679);
xor U15919 (N_15919,N_11413,N_10928);
xor U15920 (N_15920,N_12700,N_12729);
or U15921 (N_15921,N_12355,N_14399);
and U15922 (N_15922,N_14403,N_10902);
nand U15923 (N_15923,N_10118,N_14332);
or U15924 (N_15924,N_12258,N_11907);
nor U15925 (N_15925,N_13618,N_11651);
nor U15926 (N_15926,N_14501,N_11405);
xnor U15927 (N_15927,N_11100,N_13930);
and U15928 (N_15928,N_10891,N_12278);
and U15929 (N_15929,N_10120,N_11098);
or U15930 (N_15930,N_14213,N_10535);
or U15931 (N_15931,N_11616,N_10327);
and U15932 (N_15932,N_13219,N_10812);
or U15933 (N_15933,N_13227,N_10823);
and U15934 (N_15934,N_10151,N_11142);
nor U15935 (N_15935,N_14372,N_11323);
xor U15936 (N_15936,N_13015,N_10506);
nor U15937 (N_15937,N_13267,N_13670);
nand U15938 (N_15938,N_12107,N_13061);
or U15939 (N_15939,N_10629,N_11352);
nor U15940 (N_15940,N_10486,N_13416);
nand U15941 (N_15941,N_12938,N_14570);
nor U15942 (N_15942,N_11404,N_10262);
or U15943 (N_15943,N_13348,N_11520);
xor U15944 (N_15944,N_13042,N_13002);
xor U15945 (N_15945,N_13063,N_14852);
or U15946 (N_15946,N_14721,N_14861);
nor U15947 (N_15947,N_14620,N_14017);
and U15948 (N_15948,N_12603,N_12465);
nand U15949 (N_15949,N_11577,N_10508);
nand U15950 (N_15950,N_14797,N_13075);
nand U15951 (N_15951,N_12211,N_14371);
nand U15952 (N_15952,N_14417,N_14897);
and U15953 (N_15953,N_12928,N_14989);
or U15954 (N_15954,N_14002,N_14506);
and U15955 (N_15955,N_13316,N_11555);
nand U15956 (N_15956,N_13144,N_12445);
xor U15957 (N_15957,N_11741,N_13943);
nand U15958 (N_15958,N_11445,N_13901);
nor U15959 (N_15959,N_11163,N_12452);
xor U15960 (N_15960,N_14912,N_10109);
nand U15961 (N_15961,N_12261,N_10566);
xor U15962 (N_15962,N_12984,N_11258);
xor U15963 (N_15963,N_10868,N_10362);
nor U15964 (N_15964,N_10307,N_12991);
and U15965 (N_15965,N_14390,N_14525);
nor U15966 (N_15966,N_13328,N_10625);
nor U15967 (N_15967,N_10624,N_10048);
xnor U15968 (N_15968,N_14207,N_10373);
nor U15969 (N_15969,N_13303,N_10839);
and U15970 (N_15970,N_11321,N_11770);
xor U15971 (N_15971,N_11331,N_10644);
or U15972 (N_15972,N_14006,N_11743);
nor U15973 (N_15973,N_10132,N_10040);
or U15974 (N_15974,N_10092,N_14865);
nor U15975 (N_15975,N_11767,N_12077);
or U15976 (N_15976,N_13832,N_13265);
xnor U15977 (N_15977,N_13439,N_11604);
and U15978 (N_15978,N_11740,N_10801);
nand U15979 (N_15979,N_10175,N_13118);
nand U15980 (N_15980,N_14261,N_12081);
and U15981 (N_15981,N_11535,N_11356);
xor U15982 (N_15982,N_10646,N_12312);
nor U15983 (N_15983,N_12895,N_13580);
or U15984 (N_15984,N_13420,N_11080);
nor U15985 (N_15985,N_14069,N_13587);
nor U15986 (N_15986,N_10392,N_14054);
xor U15987 (N_15987,N_10071,N_12864);
nor U15988 (N_15988,N_12029,N_11167);
nand U15989 (N_15989,N_11545,N_14694);
xnor U15990 (N_15990,N_11656,N_10983);
nor U15991 (N_15991,N_11840,N_13163);
xor U15992 (N_15992,N_10275,N_10516);
and U15993 (N_15993,N_11687,N_13301);
nand U15994 (N_15994,N_14088,N_13831);
nand U15995 (N_15995,N_14454,N_11647);
or U15996 (N_15996,N_11913,N_14965);
or U15997 (N_15997,N_12783,N_12873);
nand U15998 (N_15998,N_14329,N_11719);
nand U15999 (N_15999,N_13185,N_11264);
nor U16000 (N_16000,N_10399,N_12790);
and U16001 (N_16001,N_14464,N_14568);
xor U16002 (N_16002,N_11307,N_11844);
nor U16003 (N_16003,N_13758,N_10274);
and U16004 (N_16004,N_12940,N_11421);
nand U16005 (N_16005,N_13931,N_11071);
xor U16006 (N_16006,N_11486,N_12405);
xor U16007 (N_16007,N_12554,N_13058);
and U16008 (N_16008,N_11064,N_13049);
xor U16009 (N_16009,N_12580,N_12831);
and U16010 (N_16010,N_11031,N_11964);
nor U16011 (N_16011,N_11583,N_14364);
nand U16012 (N_16012,N_12242,N_14592);
nor U16013 (N_16013,N_10849,N_14843);
nor U16014 (N_16014,N_11986,N_14599);
or U16015 (N_16015,N_12282,N_13476);
nand U16016 (N_16016,N_10782,N_12832);
nor U16017 (N_16017,N_11890,N_11493);
xor U16018 (N_16018,N_12027,N_12486);
and U16019 (N_16019,N_12009,N_10163);
or U16020 (N_16020,N_13795,N_11290);
nand U16021 (N_16021,N_13016,N_12510);
xnor U16022 (N_16022,N_13834,N_10909);
or U16023 (N_16023,N_12094,N_12579);
nor U16024 (N_16024,N_13237,N_13278);
nand U16025 (N_16025,N_14669,N_14477);
and U16026 (N_16026,N_14607,N_12406);
or U16027 (N_16027,N_10841,N_13277);
xnor U16028 (N_16028,N_11679,N_14762);
nor U16029 (N_16029,N_10104,N_10349);
and U16030 (N_16030,N_11196,N_12162);
nor U16031 (N_16031,N_12064,N_14217);
nor U16032 (N_16032,N_10675,N_11645);
nand U16033 (N_16033,N_13717,N_10081);
nor U16034 (N_16034,N_12892,N_11887);
nand U16035 (N_16035,N_12994,N_13473);
nor U16036 (N_16036,N_12793,N_11592);
nand U16037 (N_16037,N_14673,N_11997);
or U16038 (N_16038,N_10221,N_11009);
xnor U16039 (N_16039,N_11689,N_12243);
nand U16040 (N_16040,N_11534,N_11136);
nor U16041 (N_16041,N_13026,N_11891);
or U16042 (N_16042,N_14750,N_11236);
or U16043 (N_16043,N_12900,N_12395);
nor U16044 (N_16044,N_14875,N_12966);
nor U16045 (N_16045,N_14422,N_11843);
nor U16046 (N_16046,N_14361,N_14902);
nand U16047 (N_16047,N_11152,N_11750);
and U16048 (N_16048,N_12533,N_12496);
and U16049 (N_16049,N_10294,N_14241);
or U16050 (N_16050,N_13059,N_14971);
or U16051 (N_16051,N_13604,N_14925);
xor U16052 (N_16052,N_13380,N_11424);
or U16053 (N_16053,N_12473,N_10599);
or U16054 (N_16054,N_13818,N_14901);
xor U16055 (N_16055,N_13417,N_10023);
xor U16056 (N_16056,N_14165,N_10434);
or U16057 (N_16057,N_12433,N_14724);
nor U16058 (N_16058,N_14309,N_10244);
and U16059 (N_16059,N_14845,N_12488);
and U16060 (N_16060,N_13322,N_14991);
xor U16061 (N_16061,N_12400,N_14714);
nor U16062 (N_16062,N_14743,N_11920);
xnor U16063 (N_16063,N_12255,N_14341);
and U16064 (N_16064,N_13297,N_14007);
xor U16065 (N_16065,N_11731,N_10978);
xnor U16066 (N_16066,N_12283,N_14839);
nor U16067 (N_16067,N_13829,N_13312);
or U16068 (N_16068,N_14269,N_13797);
xnor U16069 (N_16069,N_12024,N_13737);
and U16070 (N_16070,N_14849,N_11856);
and U16071 (N_16071,N_12482,N_11951);
nand U16072 (N_16072,N_11177,N_11686);
nor U16073 (N_16073,N_11468,N_13101);
nand U16074 (N_16074,N_11305,N_12982);
nand U16075 (N_16075,N_12989,N_10324);
and U16076 (N_16076,N_11652,N_13759);
nand U16077 (N_16077,N_14611,N_13976);
xnor U16078 (N_16078,N_13014,N_12049);
and U16079 (N_16079,N_10834,N_12247);
and U16080 (N_16080,N_14654,N_10596);
nor U16081 (N_16081,N_14354,N_10479);
nor U16082 (N_16082,N_13025,N_12273);
and U16083 (N_16083,N_11837,N_14144);
nand U16084 (N_16084,N_13003,N_10838);
xnor U16085 (N_16085,N_13233,N_14150);
and U16086 (N_16086,N_12372,N_13401);
or U16087 (N_16087,N_13700,N_10030);
and U16088 (N_16088,N_14168,N_12104);
xnor U16089 (N_16089,N_14228,N_10003);
xor U16090 (N_16090,N_13258,N_14057);
and U16091 (N_16091,N_12712,N_14429);
or U16092 (N_16092,N_13137,N_12448);
nand U16093 (N_16093,N_11122,N_14016);
nand U16094 (N_16094,N_10102,N_10765);
or U16095 (N_16095,N_11791,N_12248);
nor U16096 (N_16096,N_11403,N_10296);
nor U16097 (N_16097,N_14733,N_11185);
or U16098 (N_16098,N_10673,N_14288);
nor U16099 (N_16099,N_12736,N_10422);
nor U16100 (N_16100,N_10272,N_13443);
and U16101 (N_16101,N_10465,N_12182);
nand U16102 (N_16102,N_12114,N_11603);
and U16103 (N_16103,N_12571,N_12777);
and U16104 (N_16104,N_11801,N_10653);
xnor U16105 (N_16105,N_12341,N_11617);
xnor U16106 (N_16106,N_10481,N_14339);
xor U16107 (N_16107,N_14418,N_14564);
and U16108 (N_16108,N_11223,N_14271);
xnor U16109 (N_16109,N_12963,N_12993);
or U16110 (N_16110,N_12848,N_12786);
xnor U16111 (N_16111,N_12319,N_11484);
xnor U16112 (N_16112,N_13451,N_14106);
nor U16113 (N_16113,N_11782,N_10047);
nor U16114 (N_16114,N_14586,N_12417);
or U16115 (N_16115,N_11853,N_10577);
xnor U16116 (N_16116,N_12466,N_12801);
xnor U16117 (N_16117,N_14924,N_14134);
or U16118 (N_16118,N_10297,N_13655);
nand U16119 (N_16119,N_10020,N_10303);
nor U16120 (N_16120,N_10697,N_12011);
nand U16121 (N_16121,N_11958,N_13987);
and U16122 (N_16122,N_11515,N_14188);
nor U16123 (N_16123,N_12872,N_12295);
or U16124 (N_16124,N_10840,N_13013);
nand U16125 (N_16125,N_14821,N_10058);
and U16126 (N_16126,N_11941,N_10322);
and U16127 (N_16127,N_13718,N_13777);
xnor U16128 (N_16128,N_10317,N_13146);
and U16129 (N_16129,N_11703,N_11044);
nand U16130 (N_16130,N_14566,N_11622);
or U16131 (N_16131,N_14617,N_12698);
and U16132 (N_16132,N_10026,N_12056);
nand U16133 (N_16133,N_13387,N_13760);
or U16134 (N_16134,N_10042,N_14913);
nor U16135 (N_16135,N_10717,N_12335);
and U16136 (N_16136,N_11313,N_10930);
nor U16137 (N_16137,N_14333,N_12701);
xor U16138 (N_16138,N_11297,N_10476);
xor U16139 (N_16139,N_14282,N_11514);
nor U16140 (N_16140,N_10198,N_10537);
nand U16141 (N_16141,N_13214,N_14559);
and U16142 (N_16142,N_10534,N_11398);
and U16143 (N_16143,N_10107,N_13647);
and U16144 (N_16144,N_12080,N_11833);
or U16145 (N_16145,N_14336,N_12697);
and U16146 (N_16146,N_10747,N_12576);
nor U16147 (N_16147,N_12123,N_10421);
and U16148 (N_16148,N_10524,N_10583);
or U16149 (N_16149,N_10602,N_13822);
nor U16150 (N_16150,N_14310,N_13340);
or U16151 (N_16151,N_11389,N_13452);
or U16152 (N_16152,N_10722,N_14404);
and U16153 (N_16153,N_12527,N_11816);
or U16154 (N_16154,N_12946,N_11137);
and U16155 (N_16155,N_13125,N_12902);
or U16156 (N_16156,N_14606,N_13337);
and U16157 (N_16157,N_10357,N_14035);
and U16158 (N_16158,N_12998,N_12722);
xnor U16159 (N_16159,N_10383,N_14067);
or U16160 (N_16160,N_13333,N_12360);
xnor U16161 (N_16161,N_11963,N_10029);
or U16162 (N_16162,N_10411,N_14796);
xnor U16163 (N_16163,N_13048,N_13499);
or U16164 (N_16164,N_10502,N_13826);
or U16165 (N_16165,N_13735,N_12015);
or U16166 (N_16166,N_14181,N_10485);
nand U16167 (N_16167,N_13000,N_11251);
nor U16168 (N_16168,N_14099,N_10304);
and U16169 (N_16169,N_10183,N_13536);
and U16170 (N_16170,N_14794,N_12660);
nor U16171 (N_16171,N_12345,N_11565);
and U16172 (N_16172,N_11472,N_14888);
xor U16173 (N_16173,N_13196,N_10439);
nand U16174 (N_16174,N_14504,N_13294);
nor U16175 (N_16175,N_14111,N_12634);
or U16176 (N_16176,N_13275,N_11339);
xnor U16177 (N_16177,N_14190,N_13178);
or U16178 (N_16178,N_10955,N_11402);
xnor U16179 (N_16179,N_13385,N_11354);
nand U16180 (N_16180,N_11900,N_14982);
xor U16181 (N_16181,N_12192,N_14407);
xnor U16182 (N_16182,N_10305,N_14508);
nor U16183 (N_16183,N_11758,N_12683);
nor U16184 (N_16184,N_10775,N_10196);
nor U16185 (N_16185,N_10628,N_12796);
and U16186 (N_16186,N_13353,N_12236);
and U16187 (N_16187,N_14388,N_14513);
xor U16188 (N_16188,N_14763,N_13980);
nor U16189 (N_16189,N_14892,N_14072);
nand U16190 (N_16190,N_11543,N_11133);
xnor U16191 (N_16191,N_11040,N_13957);
nand U16192 (N_16192,N_11250,N_14781);
and U16193 (N_16193,N_13357,N_14972);
or U16194 (N_16194,N_11757,N_11892);
xor U16195 (N_16195,N_14842,N_10388);
or U16196 (N_16196,N_10836,N_10589);
or U16197 (N_16197,N_12476,N_12368);
or U16198 (N_16198,N_10039,N_14505);
nor U16199 (N_16199,N_12364,N_11735);
and U16200 (N_16200,N_11968,N_11600);
or U16201 (N_16201,N_14374,N_12438);
nor U16202 (N_16202,N_13285,N_10186);
xnor U16203 (N_16203,N_14200,N_10028);
nor U16204 (N_16204,N_11985,N_11732);
nand U16205 (N_16205,N_14872,N_13921);
xor U16206 (N_16206,N_14567,N_14481);
and U16207 (N_16207,N_13775,N_12443);
nand U16208 (N_16208,N_14833,N_13115);
and U16209 (N_16209,N_12744,N_13535);
nand U16210 (N_16210,N_12642,N_10986);
nand U16211 (N_16211,N_11454,N_13744);
or U16212 (N_16212,N_13141,N_13823);
xnor U16213 (N_16213,N_14280,N_14751);
and U16214 (N_16214,N_11184,N_13780);
nor U16215 (N_16215,N_13745,N_13493);
and U16216 (N_16216,N_12669,N_10867);
nor U16217 (N_16217,N_10123,N_13128);
xnor U16218 (N_16218,N_12130,N_12469);
nor U16219 (N_16219,N_11267,N_14728);
or U16220 (N_16220,N_12190,N_10184);
or U16221 (N_16221,N_14717,N_12186);
and U16222 (N_16222,N_11221,N_14895);
nand U16223 (N_16223,N_13256,N_10260);
xor U16224 (N_16224,N_10046,N_12854);
or U16225 (N_16225,N_11559,N_13223);
xor U16226 (N_16226,N_14461,N_11684);
nor U16227 (N_16227,N_12779,N_13513);
xor U16228 (N_16228,N_11067,N_10069);
xnor U16229 (N_16229,N_13961,N_13849);
xor U16230 (N_16230,N_12073,N_13438);
and U16231 (N_16231,N_14065,N_10006);
nand U16232 (N_16232,N_10538,N_11294);
and U16233 (N_16233,N_11794,N_10445);
nor U16234 (N_16234,N_10025,N_14536);
xnor U16235 (N_16235,N_13282,N_12226);
and U16236 (N_16236,N_10352,N_12992);
nand U16237 (N_16237,N_12347,N_12004);
or U16238 (N_16238,N_13959,N_13236);
xor U16239 (N_16239,N_12906,N_10078);
and U16240 (N_16240,N_11799,N_14077);
nand U16241 (N_16241,N_14081,N_14731);
nand U16242 (N_16242,N_10742,N_12806);
or U16243 (N_16243,N_14819,N_13402);
nor U16244 (N_16244,N_11644,N_11509);
or U16245 (N_16245,N_10263,N_13632);
nand U16246 (N_16246,N_11353,N_10130);
xor U16247 (N_16247,N_10591,N_14302);
or U16248 (N_16248,N_10141,N_14652);
and U16249 (N_16249,N_12539,N_11746);
or U16250 (N_16250,N_11639,N_11506);
xor U16251 (N_16251,N_14693,N_13407);
or U16252 (N_16252,N_11931,N_13103);
and U16253 (N_16253,N_14708,N_13815);
and U16254 (N_16254,N_10818,N_10529);
xnor U16255 (N_16255,N_14795,N_13908);
xor U16256 (N_16256,N_14993,N_10581);
nand U16257 (N_16257,N_11143,N_12196);
nand U16258 (N_16258,N_11925,N_13198);
nand U16259 (N_16259,N_12849,N_14476);
nand U16260 (N_16260,N_11790,N_11809);
xnor U16261 (N_16261,N_10155,N_11956);
and U16262 (N_16262,N_11696,N_11776);
or U16263 (N_16263,N_14223,N_14279);
nand U16264 (N_16264,N_13210,N_11632);
nor U16265 (N_16265,N_12013,N_12508);
xor U16266 (N_16266,N_10545,N_13321);
nand U16267 (N_16267,N_13354,N_10976);
xor U16268 (N_16268,N_14125,N_13868);
nand U16269 (N_16269,N_10068,N_10202);
nor U16270 (N_16270,N_12804,N_11798);
or U16271 (N_16271,N_14790,N_11631);
or U16272 (N_16272,N_13862,N_10225);
xor U16273 (N_16273,N_14496,N_10128);
and U16274 (N_16274,N_11477,N_14141);
or U16275 (N_16275,N_14754,N_13500);
nand U16276 (N_16276,N_14803,N_14941);
and U16277 (N_16277,N_11573,N_12460);
nor U16278 (N_16278,N_10205,N_13457);
nor U16279 (N_16279,N_11453,N_13809);
xor U16280 (N_16280,N_10223,N_12687);
nand U16281 (N_16281,N_14441,N_12334);
nand U16282 (N_16282,N_12026,N_12184);
and U16283 (N_16283,N_11973,N_12407);
or U16284 (N_16284,N_13066,N_12937);
and U16285 (N_16285,N_13215,N_14528);
or U16286 (N_16286,N_11934,N_10264);
and U16287 (N_16287,N_11253,N_10498);
xor U16288 (N_16288,N_13725,N_11835);
and U16289 (N_16289,N_12165,N_10600);
nand U16290 (N_16290,N_10226,N_12875);
and U16291 (N_16291,N_10458,N_13592);
xor U16292 (N_16292,N_11212,N_13769);
or U16293 (N_16293,N_14664,N_13481);
nand U16294 (N_16294,N_13271,N_14008);
xor U16295 (N_16295,N_11829,N_14800);
or U16296 (N_16296,N_13679,N_12732);
nand U16297 (N_16297,N_12078,N_11214);
nand U16298 (N_16298,N_11155,N_11936);
or U16299 (N_16299,N_14742,N_14046);
or U16300 (N_16300,N_12320,N_12524);
nand U16301 (N_16301,N_14297,N_12160);
nor U16302 (N_16302,N_11753,N_12289);
and U16303 (N_16303,N_14629,N_12601);
xor U16304 (N_16304,N_11876,N_14367);
and U16305 (N_16305,N_10218,N_14128);
or U16306 (N_16306,N_13034,N_11952);
xor U16307 (N_16307,N_12136,N_10569);
xnor U16308 (N_16308,N_11919,N_13454);
nand U16309 (N_16309,N_13697,N_11308);
nor U16310 (N_16310,N_11003,N_13741);
xnor U16311 (N_16311,N_11507,N_12492);
or U16312 (N_16312,N_14976,N_10580);
xnor U16313 (N_16313,N_11646,N_14117);
nand U16314 (N_16314,N_13225,N_10253);
nand U16315 (N_16315,N_12453,N_13453);
nor U16316 (N_16316,N_11705,N_12301);
nand U16317 (N_16317,N_11994,N_12734);
nand U16318 (N_16318,N_13800,N_13738);
or U16319 (N_16319,N_14835,N_10168);
xnor U16320 (N_16320,N_14059,N_13224);
or U16321 (N_16321,N_10070,N_10199);
and U16322 (N_16322,N_13910,N_14446);
xnor U16323 (N_16323,N_11838,N_10770);
or U16324 (N_16324,N_11489,N_10929);
and U16325 (N_16325,N_11488,N_14515);
xnor U16326 (N_16326,N_11116,N_14812);
nor U16327 (N_16327,N_14702,N_12505);
or U16328 (N_16328,N_12945,N_10227);
or U16329 (N_16329,N_14219,N_12908);
or U16330 (N_16330,N_10888,N_11674);
nand U16331 (N_16331,N_11988,N_14232);
nand U16332 (N_16332,N_12324,N_11881);
xnor U16333 (N_16333,N_13523,N_14239);
xnor U16334 (N_16334,N_12410,N_11435);
xnor U16335 (N_16335,N_13711,N_14757);
nor U16336 (N_16336,N_11481,N_10871);
nand U16337 (N_16337,N_11427,N_14184);
and U16338 (N_16338,N_10067,N_12644);
nor U16339 (N_16339,N_12129,N_14622);
nor U16340 (N_16340,N_12773,N_14774);
nor U16341 (N_16341,N_10338,N_12297);
xor U16342 (N_16342,N_11688,N_10085);
xor U16343 (N_16343,N_13087,N_14075);
nand U16344 (N_16344,N_13993,N_12087);
nor U16345 (N_16345,N_10951,N_10798);
or U16346 (N_16346,N_11349,N_14889);
and U16347 (N_16347,N_14805,N_10076);
nor U16348 (N_16348,N_13802,N_12515);
xor U16349 (N_16349,N_14814,N_14663);
nand U16350 (N_16350,N_10483,N_14171);
xor U16351 (N_16351,N_11478,N_11747);
nand U16352 (N_16352,N_13773,N_11132);
nand U16353 (N_16353,N_13841,N_13159);
or U16354 (N_16354,N_12125,N_14551);
nor U16355 (N_16355,N_13877,N_10512);
and U16356 (N_16356,N_10680,N_10250);
xor U16357 (N_16357,N_14324,N_13505);
nor U16358 (N_16358,N_12388,N_13114);
nand U16359 (N_16359,N_14613,N_11265);
nand U16360 (N_16360,N_10454,N_14510);
and U16361 (N_16361,N_13805,N_13093);
and U16362 (N_16362,N_14832,N_13160);
xnor U16363 (N_16363,N_11409,N_14146);
xor U16364 (N_16364,N_14416,N_11538);
or U16365 (N_16365,N_11642,N_13083);
xor U16366 (N_16366,N_13170,N_14265);
or U16367 (N_16367,N_12102,N_13404);
nand U16368 (N_16368,N_11706,N_13078);
nor U16369 (N_16369,N_12903,N_10640);
or U16370 (N_16370,N_14486,N_14183);
or U16371 (N_16371,N_12155,N_14093);
and U16372 (N_16372,N_13549,N_13909);
nand U16373 (N_16373,N_14926,N_12463);
nor U16374 (N_16374,N_10098,N_12655);
nor U16375 (N_16375,N_10725,N_11038);
nor U16376 (N_16376,N_12076,N_12914);
nand U16377 (N_16377,N_13685,N_13351);
or U16378 (N_16378,N_10430,N_10224);
xnor U16379 (N_16379,N_10953,N_14419);
and U16380 (N_16380,N_11595,N_12811);
xor U16381 (N_16381,N_10280,N_14294);
xor U16382 (N_16382,N_10704,N_10432);
xor U16383 (N_16383,N_13690,N_13286);
and U16384 (N_16384,N_11675,N_13675);
and U16385 (N_16385,N_13785,N_11204);
xnor U16386 (N_16386,N_14787,N_14362);
nor U16387 (N_16387,N_14923,N_14457);
nand U16388 (N_16388,N_12610,N_11786);
nand U16389 (N_16389,N_14813,N_12277);
or U16390 (N_16390,N_14345,N_10936);
xor U16391 (N_16391,N_12630,N_12230);
xnor U16392 (N_16392,N_13046,N_10350);
or U16393 (N_16393,N_12272,N_12122);
xor U16394 (N_16394,N_14615,N_11102);
xnor U16395 (N_16395,N_12109,N_14701);
nor U16396 (N_16396,N_11061,N_10001);
nand U16397 (N_16397,N_10743,N_12430);
or U16398 (N_16398,N_11301,N_11043);
or U16399 (N_16399,N_12359,N_11315);
xor U16400 (N_16400,N_13990,N_12624);
or U16401 (N_16401,N_10517,N_12140);
nand U16402 (N_16402,N_14680,N_12715);
nor U16403 (N_16403,N_11428,N_12330);
xor U16404 (N_16404,N_10292,N_10187);
nor U16405 (N_16405,N_12475,N_14863);
or U16406 (N_16406,N_12366,N_14493);
and U16407 (N_16407,N_10471,N_12436);
nor U16408 (N_16408,N_12390,N_11256);
or U16409 (N_16409,N_12115,N_12286);
or U16410 (N_16410,N_12062,N_13273);
xnor U16411 (N_16411,N_14138,N_13634);
or U16412 (N_16412,N_13368,N_13538);
and U16413 (N_16413,N_12158,N_10103);
xor U16414 (N_16414,N_10356,N_10677);
and U16415 (N_16415,N_11896,N_13798);
xor U16416 (N_16416,N_10044,N_13881);
nor U16417 (N_16417,N_11465,N_12327);
xor U16418 (N_16418,N_10061,N_12322);
nor U16419 (N_16419,N_14502,N_14047);
nand U16420 (N_16420,N_10169,N_13483);
xnor U16421 (N_16421,N_13221,N_13440);
or U16422 (N_16422,N_13956,N_10415);
nor U16423 (N_16423,N_10933,N_12678);
nor U16424 (N_16424,N_14363,N_13942);
and U16425 (N_16425,N_14469,N_10072);
nor U16426 (N_16426,N_11324,N_11494);
nor U16427 (N_16427,N_14079,N_14135);
nand U16428 (N_16428,N_12789,N_11979);
or U16429 (N_16429,N_14434,N_13615);
xnor U16430 (N_16430,N_12431,N_12973);
nor U16431 (N_16431,N_12178,N_10475);
and U16432 (N_16432,N_10844,N_11764);
xnor U16433 (N_16433,N_14764,N_12489);
nand U16434 (N_16434,N_13859,N_12116);
nor U16435 (N_16435,N_12367,N_10283);
nor U16436 (N_16436,N_10154,N_11787);
nor U16437 (N_16437,N_13448,N_11227);
nand U16438 (N_16438,N_12652,N_11859);
and U16439 (N_16439,N_13235,N_13029);
or U16440 (N_16440,N_11343,N_10816);
xor U16441 (N_16441,N_14009,N_14063);
xnor U16442 (N_16442,N_10825,N_13106);
and U16443 (N_16443,N_12478,N_12907);
xor U16444 (N_16444,N_13487,N_13330);
or U16445 (N_16445,N_13866,N_11537);
and U16446 (N_16446,N_12487,N_14631);
xnor U16447 (N_16447,N_10386,N_13607);
and U16448 (N_16448,N_10847,N_12408);
xor U16449 (N_16449,N_13335,N_12075);
nor U16450 (N_16450,N_10576,N_12284);
nor U16451 (N_16451,N_10627,N_10685);
nand U16452 (N_16452,N_11860,N_10300);
and U16453 (N_16453,N_10480,N_13504);
nor U16454 (N_16454,N_13355,N_10701);
nor U16455 (N_16455,N_14964,N_10560);
nand U16456 (N_16456,N_13070,N_14576);
nand U16457 (N_16457,N_11295,N_14430);
or U16458 (N_16458,N_12530,N_13900);
nor U16459 (N_16459,N_13820,N_10960);
nor U16460 (N_16460,N_11778,N_12119);
nor U16461 (N_16461,N_10857,N_11289);
nand U16462 (N_16462,N_11886,N_14627);
or U16463 (N_16463,N_10862,N_11004);
xor U16464 (N_16464,N_11748,N_12859);
nor U16465 (N_16465,N_10855,N_11927);
xor U16466 (N_16466,N_10910,N_14299);
xor U16467 (N_16467,N_14152,N_13085);
nand U16468 (N_16468,N_10518,N_13683);
nor U16469 (N_16469,N_10213,N_12213);
and U16470 (N_16470,N_12365,N_11134);
and U16471 (N_16471,N_13213,N_11054);
or U16472 (N_16472,N_11156,N_14012);
xor U16473 (N_16473,N_14340,N_14876);
and U16474 (N_16474,N_13953,N_13447);
or U16475 (N_16475,N_11200,N_10698);
and U16476 (N_16476,N_12730,N_11713);
xnor U16477 (N_16477,N_14166,N_13694);
nand U16478 (N_16478,N_11788,N_13903);
and U16479 (N_16479,N_12468,N_13729);
and U16480 (N_16480,N_14021,N_10499);
and U16481 (N_16481,N_10236,N_10401);
nand U16482 (N_16482,N_13490,N_14644);
nand U16483 (N_16483,N_13713,N_10963);
nor U16484 (N_16484,N_13175,N_12632);
or U16485 (N_16485,N_13705,N_11160);
or U16486 (N_16486,N_11158,N_10135);
xor U16487 (N_16487,N_11969,N_11028);
or U16488 (N_16488,N_14767,N_11141);
nand U16489 (N_16489,N_13491,N_12997);
and U16490 (N_16490,N_12567,N_12416);
nand U16491 (N_16491,N_13749,N_12442);
or U16492 (N_16492,N_14296,N_13540);
or U16493 (N_16493,N_12306,N_11654);
nor U16494 (N_16494,N_14571,N_14189);
or U16495 (N_16495,N_11135,N_11523);
nand U16496 (N_16496,N_13260,N_12704);
or U16497 (N_16497,N_10331,N_10084);
nand U16498 (N_16498,N_10611,N_13870);
nand U16499 (N_16499,N_10382,N_10394);
or U16500 (N_16500,N_13897,N_10851);
and U16501 (N_16501,N_13730,N_11083);
nand U16502 (N_16502,N_11149,N_13702);
and U16503 (N_16503,N_14732,N_10981);
and U16504 (N_16504,N_10556,N_11636);
and U16505 (N_16505,N_13060,N_12148);
xor U16506 (N_16506,N_10971,N_11059);
and U16507 (N_16507,N_14973,N_13622);
xnor U16508 (N_16508,N_13867,N_10819);
xnor U16509 (N_16509,N_12835,N_10257);
xnor U16510 (N_16510,N_14210,N_13934);
nand U16511 (N_16511,N_14526,N_14018);
nand U16512 (N_16512,N_13516,N_10320);
nand U16513 (N_16513,N_12931,N_13801);
or U16514 (N_16514,N_11733,N_14051);
nand U16515 (N_16515,N_11283,N_14479);
xor U16516 (N_16516,N_11467,N_10491);
nor U16517 (N_16517,N_10649,N_11024);
and U16518 (N_16518,N_13204,N_13397);
nor U16519 (N_16519,N_10935,N_14579);
nor U16520 (N_16520,N_10595,N_11240);
nand U16521 (N_16521,N_14073,N_11113);
nor U16522 (N_16522,N_10926,N_11926);
nand U16523 (N_16523,N_11008,N_10313);
or U16524 (N_16524,N_10757,N_11109);
or U16525 (N_16525,N_11095,N_14287);
xnor U16526 (N_16526,N_14581,N_14683);
xor U16527 (N_16527,N_14765,N_10800);
and U16528 (N_16528,N_13027,N_14038);
nand U16529 (N_16529,N_10312,N_12353);
nor U16530 (N_16530,N_14970,N_13367);
nor U16531 (N_16531,N_12651,N_13764);
nor U16532 (N_16532,N_12180,N_11456);
nor U16533 (N_16533,N_10511,N_14490);
or U16534 (N_16534,N_12096,N_14247);
nand U16535 (N_16535,N_10074,N_12309);
or U16536 (N_16536,N_10820,N_11117);
or U16537 (N_16537,N_14100,N_14204);
nor U16538 (N_16538,N_10923,N_14052);
xor U16539 (N_16539,N_10897,N_11278);
and U16540 (N_16540,N_14857,N_10408);
nor U16541 (N_16541,N_14640,N_12936);
or U16542 (N_16542,N_12276,N_14600);
xnor U16543 (N_16543,N_10143,N_10949);
xor U16544 (N_16544,N_14259,N_11090);
and U16545 (N_16545,N_12441,N_11247);
nand U16546 (N_16546,N_12950,N_12771);
xor U16547 (N_16547,N_13623,N_13843);
nor U16548 (N_16548,N_14770,N_14741);
and U16549 (N_16549,N_14256,N_14129);
nor U16550 (N_16550,N_13475,N_10693);
nor U16551 (N_16551,N_11916,N_11022);
xor U16552 (N_16552,N_12502,N_14331);
or U16553 (N_16553,N_14151,N_10022);
and U16554 (N_16554,N_10384,N_11291);
nand U16555 (N_16555,N_10544,N_12909);
nand U16556 (N_16556,N_13640,N_12458);
and U16557 (N_16557,N_10918,N_13590);
xor U16558 (N_16558,N_10880,N_10288);
xor U16559 (N_16559,N_12157,N_14829);
xor U16560 (N_16560,N_11812,N_13496);
nor U16561 (N_16561,N_12398,N_14594);
nor U16562 (N_16562,N_12593,N_13149);
nor U16563 (N_16563,N_12540,N_11078);
or U16564 (N_16564,N_12967,N_10650);
xor U16565 (N_16565,N_14867,N_14019);
or U16566 (N_16566,N_13151,N_10251);
xor U16567 (N_16567,N_11299,N_13890);
or U16568 (N_16568,N_13671,N_12235);
xor U16569 (N_16569,N_10149,N_13596);
and U16570 (N_16570,N_11395,N_11225);
nor U16571 (N_16571,N_12113,N_14789);
nor U16572 (N_16572,N_14802,N_10013);
xnor U16573 (N_16573,N_13926,N_12422);
nor U16574 (N_16574,N_11406,N_10995);
nor U16575 (N_16575,N_11691,N_12167);
xnor U16576 (N_16576,N_12595,N_11921);
or U16577 (N_16577,N_13559,N_13247);
nor U16578 (N_16578,N_11015,N_12925);
or U16579 (N_16579,N_10419,N_14809);
nor U16580 (N_16580,N_14886,N_10969);
and U16581 (N_16581,N_13885,N_13715);
and U16582 (N_16582,N_13458,N_14637);
or U16583 (N_16583,N_11474,N_11245);
nand U16584 (N_16584,N_11215,N_11438);
nor U16585 (N_16585,N_12329,N_10674);
or U16586 (N_16586,N_11834,N_14707);
and U16587 (N_16587,N_14258,N_14735);
nand U16588 (N_16588,N_14273,N_12307);
xnor U16589 (N_16589,N_11697,N_12614);
xor U16590 (N_16590,N_11304,N_13651);
or U16591 (N_16591,N_14718,N_14651);
xnor U16592 (N_16592,N_11867,N_12470);
and U16593 (N_16593,N_12727,N_14824);
nor U16594 (N_16594,N_14705,N_14459);
or U16595 (N_16595,N_11448,N_14597);
and U16596 (N_16596,N_13593,N_14650);
xnor U16597 (N_16597,N_14532,N_11967);
nand U16598 (N_16598,N_11274,N_10753);
xor U16599 (N_16599,N_11475,N_11394);
xnor U16600 (N_16600,N_10592,N_11977);
nand U16601 (N_16601,N_10108,N_12038);
and U16602 (N_16602,N_11219,N_10817);
xor U16603 (N_16603,N_12847,N_14346);
xor U16604 (N_16604,N_12583,N_12134);
nand U16605 (N_16605,N_14494,N_13239);
xnor U16606 (N_16606,N_12340,N_12743);
and U16607 (N_16607,N_11455,N_10622);
nand U16608 (N_16608,N_11482,N_11213);
xnor U16609 (N_16609,N_13975,N_10531);
and U16610 (N_16610,N_14179,N_10266);
xor U16611 (N_16611,N_10456,N_14045);
nor U16612 (N_16612,N_12817,N_10395);
nor U16613 (N_16613,N_14218,N_12185);
and U16614 (N_16614,N_13965,N_12432);
and U16615 (N_16615,N_12748,N_13205);
xor U16616 (N_16616,N_12001,N_14262);
xor U16617 (N_16617,N_12924,N_14655);
and U16618 (N_16618,N_11052,N_14573);
or U16619 (N_16619,N_14939,N_14847);
xnor U16620 (N_16620,N_14020,N_12616);
or U16621 (N_16621,N_13905,N_12336);
nand U16622 (N_16622,N_13875,N_13107);
and U16623 (N_16623,N_14736,N_12765);
nor U16624 (N_16624,N_11370,N_10323);
nand U16625 (N_16625,N_10954,N_13569);
and U16626 (N_16626,N_12821,N_11699);
xor U16627 (N_16627,N_13383,N_12759);
xor U16628 (N_16628,N_13251,N_10585);
nor U16629 (N_16629,N_11310,N_11729);
nand U16630 (N_16630,N_11810,N_13023);
or U16631 (N_16631,N_14444,N_10507);
or U16632 (N_16632,N_10663,N_10207);
or U16633 (N_16633,N_10428,N_12147);
nor U16634 (N_16634,N_10752,N_10258);
or U16635 (N_16635,N_13619,N_10052);
or U16636 (N_16636,N_13484,N_13174);
nand U16637 (N_16637,N_13778,N_14775);
or U16638 (N_16638,N_12962,N_14010);
nand U16639 (N_16639,N_10339,N_11029);
and U16640 (N_16640,N_14859,N_12415);
nor U16641 (N_16641,N_14001,N_10547);
xor U16642 (N_16642,N_12493,N_11387);
or U16643 (N_16643,N_14922,N_12485);
nand U16644 (N_16644,N_13188,N_12695);
xnor U16645 (N_16645,N_11422,N_10159);
xnor U16646 (N_16646,N_12677,N_13682);
nor U16647 (N_16647,N_12568,N_13081);
xnor U16648 (N_16648,N_11738,N_10094);
nor U16649 (N_16649,N_13757,N_12380);
nor U16650 (N_16650,N_13232,N_13966);
or U16651 (N_16651,N_14681,N_12053);
or U16652 (N_16652,N_13863,N_14540);
nand U16653 (N_16653,N_10850,N_12851);
nor U16654 (N_16654,N_13692,N_14961);
and U16655 (N_16655,N_12757,N_13947);
xnor U16656 (N_16656,N_11795,N_14384);
nand U16657 (N_16657,N_11808,N_12827);
nor U16658 (N_16658,N_12121,N_10739);
xnor U16659 (N_16659,N_11933,N_10721);
xor U16660 (N_16660,N_10050,N_13792);
xnor U16661 (N_16661,N_13450,N_10554);
and U16662 (N_16662,N_14442,N_12370);
nor U16663 (N_16663,N_11661,N_14028);
xnor U16664 (N_16664,N_13319,N_12922);
or U16665 (N_16665,N_14319,N_11803);
nor U16666 (N_16666,N_12050,N_12523);
and U16667 (N_16667,N_11845,N_11303);
or U16668 (N_16668,N_10185,N_11769);
nand U16669 (N_16669,N_10340,N_13624);
and U16670 (N_16670,N_12234,N_12820);
or U16671 (N_16671,N_12321,N_10711);
or U16672 (N_16672,N_13498,N_10541);
nand U16673 (N_16673,N_10714,N_14818);
nor U16674 (N_16674,N_14799,N_11961);
nand U16675 (N_16675,N_10452,N_10217);
nor U16676 (N_16676,N_13018,N_11692);
nand U16677 (N_16677,N_13350,N_14170);
nor U16678 (N_16678,N_13054,N_12846);
or U16679 (N_16679,N_12519,N_12979);
xor U16680 (N_16680,N_12838,N_12041);
or U16681 (N_16681,N_10056,N_11815);
xnor U16682 (N_16682,N_13555,N_10379);
nor U16683 (N_16683,N_12912,N_13812);
or U16684 (N_16684,N_13553,N_13603);
nand U16685 (N_16685,N_11420,N_11851);
or U16686 (N_16686,N_10699,N_10703);
nor U16687 (N_16687,N_11371,N_12210);
nand U16688 (N_16688,N_11572,N_14887);
nand U16689 (N_16689,N_10638,N_14990);
or U16690 (N_16690,N_12229,N_14690);
or U16691 (N_16691,N_12918,N_13527);
nor U16692 (N_16692,N_10832,N_10946);
and U16693 (N_16693,N_10872,N_14776);
xor U16694 (N_16694,N_10173,N_14704);
nand U16695 (N_16695,N_14452,N_11745);
nor U16696 (N_16696,N_11990,N_14359);
nand U16697 (N_16697,N_14064,N_12499);
nor U16698 (N_16698,N_12543,N_14227);
and U16699 (N_16699,N_13126,N_11497);
and U16700 (N_16700,N_11923,N_12662);
and U16701 (N_16701,N_12377,N_10588);
or U16702 (N_16702,N_12890,N_12797);
and U16703 (N_16703,N_12239,N_11736);
and U16704 (N_16704,N_12292,N_14748);
nor U16705 (N_16705,N_11359,N_11590);
xor U16706 (N_16706,N_14391,N_13552);
nand U16707 (N_16707,N_14879,N_11781);
nand U16708 (N_16708,N_10579,N_12127);
nand U16709 (N_16709,N_10689,N_13053);
and U16710 (N_16710,N_10443,N_11846);
and U16711 (N_16711,N_13600,N_12270);
nor U16712 (N_16712,N_14236,N_13388);
nand U16713 (N_16713,N_11673,N_14711);
xor U16714 (N_16714,N_11775,N_12507);
or U16715 (N_16715,N_10950,N_11737);
nor U16716 (N_16716,N_10147,N_12126);
nor U16717 (N_16717,N_13343,N_12199);
nand U16718 (N_16718,N_13662,N_11431);
nand U16719 (N_16719,N_13971,N_13356);
or U16720 (N_16720,N_11473,N_11574);
nor U16721 (N_16721,N_10860,N_13996);
and U16722 (N_16722,N_10900,N_12952);
and U16723 (N_16723,N_14483,N_14132);
and U16724 (N_16724,N_11287,N_13917);
nor U16725 (N_16725,N_11817,N_14980);
and U16726 (N_16726,N_13092,N_13375);
nor U16727 (N_16727,N_10097,N_11154);
nand U16728 (N_16728,N_11334,N_10330);
and U16729 (N_16729,N_12619,N_12808);
or U16730 (N_16730,N_14577,N_13226);
xor U16731 (N_16731,N_11885,N_10418);
xor U16732 (N_16732,N_12042,N_12843);
nor U16733 (N_16733,N_12033,N_13621);
nor U16734 (N_16734,N_10786,N_11042);
nor U16735 (N_16735,N_12913,N_14822);
nand U16736 (N_16736,N_12451,N_12231);
and U16737 (N_16737,N_13426,N_10814);
nor U16738 (N_16738,N_14327,N_12577);
or U16739 (N_16739,N_10472,N_14074);
nand U16740 (N_16740,N_11708,N_11870);
or U16741 (N_16741,N_11634,N_14598);
and U16742 (N_16742,N_14906,N_12787);
and U16743 (N_16743,N_14044,N_10309);
xor U16744 (N_16744,N_11998,N_12822);
or U16745 (N_16745,N_12641,N_10146);
and U16746 (N_16746,N_13648,N_12120);
xor U16747 (N_16747,N_14437,N_14908);
xnor U16748 (N_16748,N_11525,N_10016);
nor U16749 (N_16749,N_11179,N_12036);
nand U16750 (N_16750,N_12403,N_12019);
or U16751 (N_16751,N_14160,N_10641);
and U16752 (N_16752,N_14878,N_13846);
nand U16753 (N_16753,N_14710,N_10242);
or U16754 (N_16754,N_13248,N_14278);
or U16755 (N_16755,N_13434,N_12479);
or U16756 (N_16756,N_11615,N_14588);
nand U16757 (N_16757,N_14997,N_10992);
xnor U16758 (N_16758,N_12573,N_11203);
or U16759 (N_16759,N_13296,N_12291);
or U16760 (N_16760,N_10893,N_10808);
and U16761 (N_16761,N_13084,N_11897);
and U16762 (N_16762,N_13933,N_13883);
nor U16763 (N_16763,N_12898,N_14307);
nand U16764 (N_16764,N_13152,N_13674);
or U16765 (N_16765,N_12761,N_14715);
and U16766 (N_16766,N_14944,N_14470);
nand U16767 (N_16767,N_10211,N_13786);
xnor U16768 (N_16768,N_14987,N_12323);
and U16769 (N_16769,N_11330,N_12419);
or U16770 (N_16770,N_12108,N_12141);
xor U16771 (N_16771,N_14196,N_13203);
nand U16772 (N_16772,N_13661,N_12649);
or U16773 (N_16773,N_10051,N_14646);
nand U16774 (N_16774,N_11563,N_11561);
nor U16775 (N_16775,N_11087,N_12929);
and U16776 (N_16776,N_12285,N_10059);
or U16777 (N_16777,N_13077,N_11570);
and U16778 (N_16778,N_11908,N_11210);
or U16779 (N_16779,N_11146,N_12412);
xor U16780 (N_16780,N_10688,N_10165);
nand U16781 (N_16781,N_10449,N_10952);
or U16782 (N_16782,N_10866,N_12197);
nand U16783 (N_16783,N_12039,N_13967);
nand U16784 (N_16784,N_11384,N_11821);
xnor U16785 (N_16785,N_14303,N_14558);
nand U16786 (N_16786,N_11976,N_11198);
xor U16787 (N_16787,N_13123,N_13202);
and U16788 (N_16788,N_12693,N_10459);
or U16789 (N_16789,N_14136,N_12084);
xor U16790 (N_16790,N_12724,N_10684);
and U16791 (N_16791,N_14449,N_10616);
xnor U16792 (N_16792,N_12399,N_11541);
nand U16793 (N_16793,N_14618,N_10287);
xor U16794 (N_16794,N_12570,N_14688);
or U16795 (N_16795,N_13838,N_11496);
nor U16796 (N_16796,N_10450,N_13558);
xor U16797 (N_16797,N_11715,N_10241);
xor U16798 (N_16798,N_13358,N_11444);
or U16799 (N_16799,N_10626,N_11293);
xnor U16800 (N_16800,N_10122,N_14406);
nand U16801 (N_16801,N_13386,N_12191);
and U16802 (N_16802,N_14783,N_13311);
nand U16803 (N_16803,N_10903,N_11164);
nand U16804 (N_16804,N_14561,N_13099);
and U16805 (N_16805,N_14699,N_12007);
or U16806 (N_16806,N_14727,N_13127);
or U16807 (N_16807,N_12455,N_13964);
xnor U16808 (N_16808,N_12070,N_10398);
nand U16809 (N_16809,N_11825,N_12378);
or U16810 (N_16810,N_12561,N_14025);
xor U16811 (N_16811,N_10326,N_13528);
nor U16812 (N_16812,N_10667,N_10793);
nor U16813 (N_16813,N_11712,N_13489);
xor U16814 (N_16814,N_11257,N_12987);
nor U16815 (N_16815,N_10536,N_13782);
and U16816 (N_16816,N_12467,N_13982);
or U16817 (N_16817,N_13657,N_10730);
xor U16818 (N_16818,N_12022,N_12006);
and U16819 (N_16819,N_13939,N_14686);
xor U16820 (N_16820,N_11768,N_12916);
nor U16821 (N_16821,N_13269,N_13639);
or U16822 (N_16822,N_13904,N_12557);
and U16823 (N_16823,N_10759,N_12337);
and U16824 (N_16824,N_13072,N_14634);
or U16825 (N_16825,N_13907,N_10553);
nand U16826 (N_16826,N_11915,N_10789);
nand U16827 (N_16827,N_11292,N_10137);
nor U16828 (N_16828,N_11337,N_14788);
xnor U16829 (N_16829,N_10049,N_11407);
nor U16830 (N_16830,N_13984,N_13307);
nor U16831 (N_16831,N_13231,N_12883);
nand U16832 (N_16832,N_14910,N_14649);
or U16833 (N_16833,N_12103,N_10194);
nand U16834 (N_16834,N_12401,N_14768);
nand U16835 (N_16835,N_14747,N_12358);
nor U16836 (N_16836,N_11883,N_11640);
nor U16837 (N_16837,N_13393,N_12720);
nand U16838 (N_16838,N_12706,N_11759);
xor U16839 (N_16839,N_12418,N_12280);
and U16840 (N_16840,N_14235,N_14516);
and U16841 (N_16841,N_11441,N_11796);
xnor U16842 (N_16842,N_14368,N_14036);
xor U16843 (N_16843,N_11275,N_14109);
and U16844 (N_16844,N_11762,N_14920);
or U16845 (N_16845,N_14605,N_14124);
nor U16846 (N_16846,N_10922,N_14102);
and U16847 (N_16847,N_14083,N_13594);
and U16848 (N_16848,N_13197,N_12926);
nor U16849 (N_16849,N_14777,N_10405);
nand U16850 (N_16850,N_13384,N_12137);
or U16851 (N_16851,N_12294,N_13184);
nor U16852 (N_16852,N_12005,N_10549);
nand U16853 (N_16853,N_10672,N_14798);
nand U16854 (N_16854,N_14884,N_12689);
and U16855 (N_16855,N_12223,N_13257);
nand U16856 (N_16856,N_11045,N_12622);
xor U16857 (N_16857,N_14806,N_12066);
or U16858 (N_16858,N_14666,N_10461);
or U16859 (N_16859,N_12293,N_12000);
and U16860 (N_16860,N_14648,N_14313);
or U16861 (N_16861,N_11598,N_12260);
nand U16862 (N_16862,N_13617,N_12675);
and U16863 (N_16863,N_12346,N_14547);
or U16864 (N_16864,N_14268,N_13922);
and U16865 (N_16865,N_14684,N_12726);
and U16866 (N_16866,N_11001,N_12168);
and U16867 (N_16867,N_14643,N_14317);
nand U16868 (N_16868,N_10810,N_14090);
nand U16869 (N_16869,N_10181,N_13958);
xor U16870 (N_16870,N_11232,N_14379);
or U16871 (N_16871,N_14027,N_14342);
xor U16872 (N_16872,N_10890,N_10235);
nand U16873 (N_16873,N_11755,N_10347);
nand U16874 (N_16874,N_11396,N_14252);
and U16875 (N_16875,N_12391,N_14928);
and U16876 (N_16876,N_13409,N_13243);
nand U16877 (N_16877,N_11772,N_14266);
xnor U16878 (N_16878,N_14312,N_11542);
or U16879 (N_16879,N_12774,N_14580);
or U16880 (N_16880,N_10615,N_10964);
xor U16881 (N_16881,N_12661,N_14070);
or U16882 (N_16882,N_10116,N_11763);
and U16883 (N_16883,N_14855,N_14520);
nand U16884 (N_16884,N_11021,N_14484);
nor U16885 (N_16885,N_14759,N_11693);
and U16886 (N_16886,N_14432,N_13028);
nor U16887 (N_16887,N_10705,N_11579);
nor U16888 (N_16888,N_11949,N_13839);
nor U16889 (N_16889,N_14315,N_10662);
nor U16890 (N_16890,N_10138,N_13437);
xnor U16891 (N_16891,N_11151,N_13069);
nor U16892 (N_16892,N_13583,N_13194);
and U16893 (N_16893,N_11804,N_10754);
xor U16894 (N_16894,N_12175,N_12794);
and U16895 (N_16895,N_12088,N_13703);
nor U16896 (N_16896,N_12132,N_13120);
and U16897 (N_16897,N_14169,N_14284);
and U16898 (N_16898,N_12296,N_10864);
or U16899 (N_16899,N_13465,N_11850);
and U16900 (N_16900,N_11548,N_12685);
nor U16901 (N_16901,N_10451,N_11347);
xor U16902 (N_16902,N_10837,N_11190);
nor U16903 (N_16903,N_10877,N_11576);
and U16904 (N_16904,N_10664,N_11669);
xnor U16905 (N_16905,N_11698,N_12657);
and U16906 (N_16906,N_13497,N_12714);
xor U16907 (N_16907,N_12025,N_11982);
or U16908 (N_16908,N_13653,N_13136);
and U16909 (N_16909,N_13970,N_11385);
and U16910 (N_16910,N_11591,N_13784);
nand U16911 (N_16911,N_10361,N_13752);
xor U16912 (N_16912,N_10277,N_12003);
nor U16913 (N_16913,N_11471,N_12536);
nor U16914 (N_16914,N_11974,N_14465);
xnor U16915 (N_16915,N_13991,N_12414);
or U16916 (N_16916,N_11861,N_14245);
and U16917 (N_16917,N_11180,N_10806);
nand U16918 (N_16918,N_13032,N_11955);
nand U16919 (N_16919,N_12311,N_12500);
nor U16920 (N_16920,N_12537,N_14107);
or U16921 (N_16921,N_13902,N_10842);
xor U16922 (N_16922,N_11270,N_10601);
xor U16923 (N_16923,N_10966,N_11479);
xor U16924 (N_16924,N_12183,N_11659);
xnor U16925 (N_16925,N_10510,N_11188);
nor U16926 (N_16926,N_13886,N_13035);
nand U16927 (N_16927,N_11035,N_14871);
nand U16928 (N_16928,N_12813,N_14723);
xor U16929 (N_16929,N_11147,N_12143);
or U16930 (N_16930,N_12927,N_12799);
nand U16931 (N_16931,N_11286,N_13249);
or U16932 (N_16932,N_10279,N_10527);
and U16933 (N_16933,N_12682,N_14435);
or U16934 (N_16934,N_12356,N_14885);
and U16935 (N_16935,N_13403,N_14355);
nor U16936 (N_16936,N_14082,N_10420);
or U16937 (N_16937,N_12911,N_14784);
nor U16938 (N_16938,N_13791,N_12135);
nand U16939 (N_16939,N_13835,N_13382);
or U16940 (N_16940,N_12877,N_12691);
xnor U16941 (N_16941,N_11962,N_12528);
xor U16942 (N_16942,N_14720,N_13095);
xor U16943 (N_16943,N_10315,N_10160);
nor U16944 (N_16944,N_13876,N_13514);
xnor U16945 (N_16945,N_12939,N_12023);
and U16946 (N_16946,N_13390,N_13570);
xor U16947 (N_16947,N_12983,N_11996);
xor U16948 (N_16948,N_13663,N_12152);
nand U16949 (N_16949,N_12923,N_10612);
or U16950 (N_16950,N_13664,N_14773);
nor U16951 (N_16951,N_11959,N_10268);
or U16952 (N_16952,N_13220,N_14554);
xor U16953 (N_16953,N_13140,N_11513);
and U16954 (N_16954,N_11076,N_14161);
nor U16955 (N_16955,N_14981,N_10446);
nand U16956 (N_16956,N_14868,N_10790);
nor U16957 (N_16957,N_13338,N_12166);
or U16958 (N_16958,N_12387,N_10066);
or U16959 (N_16959,N_13803,N_12381);
nor U16960 (N_16960,N_14306,N_14729);
xnor U16961 (N_16961,N_11246,N_10807);
nor U16962 (N_16962,N_11567,N_10440);
or U16963 (N_16963,N_10259,N_11940);
nor U16964 (N_16964,N_10852,N_11425);
xor U16965 (N_16965,N_12935,N_14638);
nor U16966 (N_16966,N_14353,N_10683);
nor U16967 (N_16967,N_10740,N_12865);
xnor U16968 (N_16968,N_12776,N_12389);
or U16969 (N_16969,N_14208,N_13494);
and U16970 (N_16970,N_10927,N_10784);
nor U16971 (N_16971,N_10785,N_11672);
or U16972 (N_16972,N_10894,N_13157);
xor U16973 (N_16973,N_13582,N_12552);
or U16974 (N_16974,N_11701,N_11879);
xor U16975 (N_16975,N_11033,N_13644);
or U16976 (N_16976,N_11784,N_12514);
xor U16977 (N_16977,N_10348,N_10635);
or U16978 (N_16978,N_11369,N_14263);
nand U16979 (N_16979,N_14337,N_13259);
nor U16980 (N_16980,N_11638,N_12349);
nand U16981 (N_16981,N_14014,N_10190);
xnor U16982 (N_16982,N_11718,N_10974);
or U16983 (N_16983,N_14523,N_10741);
nand U16984 (N_16984,N_14929,N_12725);
nor U16985 (N_16985,N_10500,N_13037);
xor U16986 (N_16986,N_13169,N_14246);
nand U16987 (N_16987,N_11228,N_13050);
or U16988 (N_16988,N_10017,N_14545);
or U16989 (N_16989,N_11442,N_11182);
nor U16990 (N_16990,N_11207,N_10618);
and U16991 (N_16991,N_10979,N_14330);
or U16992 (N_16992,N_11495,N_11828);
and U16993 (N_16993,N_14753,N_11948);
or U16994 (N_16994,N_14026,N_12225);
nor U16995 (N_16995,N_12995,N_10376);
and U16996 (N_16996,N_14949,N_11765);
and U16997 (N_16997,N_10941,N_11206);
or U16998 (N_16998,N_11322,N_11419);
nand U16999 (N_16999,N_10642,N_13011);
and U17000 (N_17000,N_12266,N_10254);
xnor U17001 (N_17001,N_11079,N_10237);
or U17002 (N_17002,N_14358,N_10087);
and U17003 (N_17003,N_12703,N_14862);
nor U17004 (N_17004,N_13270,N_11226);
xor U17005 (N_17005,N_13176,N_10427);
xnor U17006 (N_17006,N_14097,N_13021);
nor U17007 (N_17007,N_13537,N_10381);
nor U17008 (N_17008,N_13421,N_11131);
xnor U17009 (N_17009,N_14744,N_10053);
nor U17010 (N_17010,N_13400,N_14237);
nand U17011 (N_17011,N_13471,N_13299);
and U17012 (N_17012,N_12981,N_11811);
xor U17013 (N_17013,N_10744,N_11807);
and U17014 (N_17014,N_11744,N_14543);
or U17015 (N_17015,N_14462,N_10781);
and U17016 (N_17016,N_13837,N_12454);
nand U17017 (N_17017,N_14142,N_14820);
nand U17018 (N_17018,N_11628,N_13665);
nand U17019 (N_17019,N_13254,N_11544);
xor U17020 (N_17020,N_14349,N_14103);
nand U17021 (N_17021,N_10944,N_12834);
nand U17022 (N_17022,N_14127,N_10139);
or U17023 (N_17023,N_10924,N_10038);
nor U17024 (N_17024,N_12520,N_10416);
nand U17025 (N_17025,N_13288,N_10126);
and U17026 (N_17026,N_10829,N_11912);
and U17027 (N_17027,N_11378,N_10444);
nor U17028 (N_17028,N_10853,N_13052);
and U17029 (N_17029,N_12206,N_10780);
and U17030 (N_17030,N_10773,N_10010);
nand U17031 (N_17031,N_13228,N_11235);
or U17032 (N_17032,N_13850,N_14780);
nor U17033 (N_17033,N_12531,N_13643);
xnor U17034 (N_17034,N_13374,N_11388);
and U17035 (N_17035,N_13320,N_11991);
nor U17036 (N_17036,N_11671,N_13339);
nand U17037 (N_17037,N_11189,N_12639);
and U17038 (N_17038,N_11070,N_13378);
xnor U17039 (N_17039,N_13995,N_14665);
or U17040 (N_17040,N_11989,N_14752);
nor U17041 (N_17041,N_13501,N_13430);
and U17042 (N_17042,N_13502,N_14918);
and U17043 (N_17043,N_14831,N_10063);
xnor U17044 (N_17044,N_10515,N_13871);
nor U17045 (N_17045,N_12089,N_13585);
and U17046 (N_17046,N_10565,N_10731);
and U17047 (N_17047,N_10230,N_10216);
nand U17048 (N_17048,N_14023,N_11089);
or U17049 (N_17049,N_10423,N_10620);
or U17050 (N_17050,N_11944,N_10086);
and U17051 (N_17051,N_10661,N_10606);
nor U17052 (N_17052,N_10371,N_12588);
and U17053 (N_17053,N_11995,N_10728);
xnor U17054 (N_17054,N_10468,N_12951);
or U17055 (N_17055,N_11020,N_10645);
xnor U17056 (N_17056,N_14352,N_10582);
nor U17057 (N_17057,N_14274,N_11263);
and U17058 (N_17058,N_14455,N_14381);
nand U17059 (N_17059,N_13509,N_11929);
xor U17060 (N_17060,N_13923,N_14276);
xnor U17061 (N_17061,N_11002,N_11161);
and U17062 (N_17062,N_10219,N_10760);
nand U17063 (N_17063,N_12054,N_13263);
nor U17064 (N_17064,N_14300,N_10273);
and U17065 (N_17065,N_13131,N_10520);
and U17066 (N_17066,N_12409,N_11502);
nand U17067 (N_17067,N_11947,N_13292);
or U17068 (N_17068,N_11683,N_10270);
nand U17069 (N_17069,N_13520,N_14495);
nor U17070 (N_17070,N_11774,N_12498);
xor U17071 (N_17071,N_13166,N_14834);
xnor U17072 (N_17072,N_10764,N_12172);
xor U17073 (N_17073,N_11965,N_14676);
nor U17074 (N_17074,N_12628,N_10082);
and U17075 (N_17075,N_14281,N_12853);
xnor U17076 (N_17076,N_14844,N_13601);
and U17077 (N_17077,N_10905,N_10802);
xnor U17078 (N_17078,N_12631,N_11766);
nor U17079 (N_17079,N_13779,N_11166);
and U17080 (N_17080,N_12948,N_11118);
nand U17081 (N_17081,N_13412,N_13071);
xnor U17082 (N_17082,N_13461,N_10575);
and U17083 (N_17083,N_11527,N_14220);
nor U17084 (N_17084,N_13179,N_14178);
nand U17085 (N_17085,N_14846,N_12171);
and U17086 (N_17086,N_10555,N_12526);
xor U17087 (N_17087,N_11053,N_14621);
nor U17088 (N_17088,N_12350,N_13467);
nor U17089 (N_17089,N_12954,N_14133);
xor U17090 (N_17090,N_13566,N_12654);
and U17091 (N_17091,N_10594,N_11393);
nand U17092 (N_17092,N_12503,N_14091);
and U17093 (N_17093,N_11229,N_10501);
and U17094 (N_17094,N_11749,N_13940);
or U17095 (N_17095,N_10096,N_10345);
xnor U17096 (N_17096,N_13446,N_12328);
or U17097 (N_17097,N_12151,N_11130);
and U17098 (N_17098,N_13242,N_12047);
nor U17099 (N_17099,N_11602,N_12082);
and U17100 (N_17100,N_14253,N_12456);
xnor U17101 (N_17101,N_12627,N_13565);
or U17102 (N_17102,N_12085,N_14914);
and U17103 (N_17103,N_12623,N_10492);
and U17104 (N_17104,N_12749,N_14121);
nand U17105 (N_17105,N_10777,N_13855);
and U17106 (N_17106,N_10435,N_10988);
nand U17107 (N_17107,N_12608,N_14326);
and U17108 (N_17108,N_13331,N_10708);
or U17109 (N_17109,N_11205,N_14224);
nor U17110 (N_17110,N_14932,N_14909);
xor U17111 (N_17111,N_11111,N_14177);
nor U17112 (N_17112,N_11005,N_12803);
xor U17113 (N_17113,N_10968,N_12263);
nor U17114 (N_17114,N_10961,N_13108);
or U17115 (N_17115,N_12582,N_13470);
nand U17116 (N_17116,N_14630,N_13216);
xnor U17117 (N_17117,N_12224,N_10041);
xnor U17118 (N_17118,N_10256,N_10908);
nand U17119 (N_17119,N_11637,N_11056);
or U17120 (N_17120,N_14556,N_11051);
xnor U17121 (N_17121,N_12944,N_14347);
nor U17122 (N_17122,N_12201,N_12976);
or U17123 (N_17123,N_11607,N_13588);
or U17124 (N_17124,N_13840,N_11176);
or U17125 (N_17125,N_13672,N_11178);
or U17126 (N_17126,N_11050,N_10972);
nand U17127 (N_17127,N_12891,N_11551);
and U17128 (N_17128,N_11826,N_11433);
nor U17129 (N_17129,N_11568,N_14791);
nand U17130 (N_17130,N_14830,N_13983);
xnor U17131 (N_17131,N_12101,N_12517);
xnor U17132 (N_17132,N_14548,N_12735);
nor U17133 (N_17133,N_10131,N_13793);
nor U17134 (N_17134,N_10720,N_12274);
nor U17135 (N_17135,N_13372,N_10015);
nor U17136 (N_17136,N_14935,N_12426);
or U17137 (N_17137,N_10822,N_13332);
nand U17138 (N_17138,N_14043,N_11709);
nand U17139 (N_17139,N_11092,N_12222);
or U17140 (N_17140,N_11865,N_13181);
xnor U17141 (N_17141,N_11569,N_13427);
or U17142 (N_17142,N_12932,N_12541);
nor U17143 (N_17143,N_11439,N_12947);
nand U17144 (N_17144,N_12095,N_12058);
nand U17145 (N_17145,N_10648,N_11110);
nand U17146 (N_17146,N_11714,N_13132);
nor U17147 (N_17147,N_11350,N_13062);
nor U17148 (N_17148,N_11273,N_13794);
or U17149 (N_17149,N_13649,N_12676);
or U17150 (N_17150,N_11101,N_11621);
nand U17151 (N_17151,N_11609,N_12207);
nand U17152 (N_17152,N_14460,N_12471);
or U17153 (N_17153,N_11316,N_13529);
and U17154 (N_17154,N_11664,N_12917);
nor U17155 (N_17155,N_11643,N_14463);
xor U17156 (N_17156,N_10607,N_13268);
or U17157 (N_17157,N_12060,N_11039);
nand U17158 (N_17158,N_11285,N_11540);
nand U17159 (N_17159,N_10959,N_11871);
and U17160 (N_17160,N_11366,N_10652);
nand U17161 (N_17161,N_11103,N_10889);
or U17162 (N_17162,N_13187,N_13262);
nand U17163 (N_17163,N_12079,N_13804);
or U17164 (N_17164,N_14647,N_12977);
nand U17165 (N_17165,N_14096,N_12551);
nor U17166 (N_17166,N_10660,N_12481);
and U17167 (N_17167,N_12887,N_14378);
and U17168 (N_17168,N_13830,N_14537);
nand U17169 (N_17169,N_10987,N_12354);
nor U17170 (N_17170,N_13086,N_14301);
and U17171 (N_17171,N_14335,N_11657);
nand U17172 (N_17172,N_11893,N_10879);
nand U17173 (N_17173,N_14380,N_13056);
and U17174 (N_17174,N_11662,N_11724);
or U17175 (N_17175,N_11505,N_13295);
and U17176 (N_17176,N_14254,N_13530);
or U17177 (N_17177,N_10552,N_11282);
xnor U17178 (N_17178,N_13873,N_11700);
and U17179 (N_17179,N_12721,N_13369);
nor U17180 (N_17180,N_11181,N_13997);
nor U17181 (N_17181,N_11362,N_11681);
nor U17182 (N_17182,N_12620,N_13004);
nand U17183 (N_17183,N_13364,N_13681);
nand U17184 (N_17184,N_14216,N_13264);
xor U17185 (N_17185,N_12740,N_11677);
and U17186 (N_17186,N_11073,N_13742);
and U17187 (N_17187,N_11519,N_10179);
and U17188 (N_17188,N_12825,N_10180);
or U17189 (N_17189,N_13512,N_11248);
or U17190 (N_17190,N_14369,N_10863);
or U17191 (N_17191,N_14985,N_12823);
nor U17192 (N_17192,N_13110,N_13743);
xnor U17193 (N_17193,N_11727,N_10249);
nand U17194 (N_17194,N_11336,N_13201);
xnor U17195 (N_17195,N_13847,N_11660);
nor U17196 (N_17196,N_12841,N_11874);
or U17197 (N_17197,N_12615,N_10873);
xnor U17198 (N_17198,N_14817,N_12535);
or U17199 (N_17199,N_14439,N_12667);
and U17200 (N_17200,N_13616,N_13807);
nor U17201 (N_17201,N_10756,N_11088);
and U17202 (N_17202,N_14927,N_13765);
or U17203 (N_17203,N_14550,N_12338);
and U17204 (N_17204,N_12138,N_13158);
nand U17205 (N_17205,N_14131,N_12342);
nor U17206 (N_17206,N_14375,N_12980);
nor U17207 (N_17207,N_11633,N_14408);
and U17208 (N_17208,N_13429,N_11329);
xnor U17209 (N_17209,N_12884,N_13614);
and U17210 (N_17210,N_11298,N_13641);
xnor U17211 (N_17211,N_11390,N_10523);
and U17212 (N_17212,N_10174,N_12105);
xnor U17213 (N_17213,N_14172,N_10012);
xor U17214 (N_17214,N_14826,N_14779);
nor U17215 (N_17215,N_14838,N_12594);
nor U17216 (N_17216,N_11562,N_11611);
and U17217 (N_17217,N_12708,N_10525);
nand U17218 (N_17218,N_11901,N_11380);
nor U17219 (N_17219,N_12880,N_14383);
or U17220 (N_17220,N_13057,N_10189);
xor U17221 (N_17221,N_12625,N_14848);
nand U17222 (N_17222,N_12256,N_14316);
or U17223 (N_17223,N_12361,N_13882);
and U17224 (N_17224,N_10366,N_11802);
and U17225 (N_17225,N_10821,N_13238);
and U17226 (N_17226,N_14211,N_14992);
nor U17227 (N_17227,N_12930,N_14031);
nor U17228 (N_17228,N_11950,N_10024);
xor U17229 (N_17229,N_10441,N_13808);
nand U17230 (N_17230,N_11466,N_11601);
nor U17231 (N_17231,N_14948,N_11281);
nand U17232 (N_17232,N_14979,N_13039);
xnor U17233 (N_17233,N_12653,N_14521);
nand U17234 (N_17234,N_10364,N_14401);
or U17235 (N_17235,N_14535,N_12752);
and U17236 (N_17236,N_13605,N_12237);
xor U17237 (N_17237,N_10095,N_10858);
nand U17238 (N_17238,N_10161,N_14320);
nor U17239 (N_17239,N_12780,N_11121);
xor U17240 (N_17240,N_13851,N_13951);
and U17241 (N_17241,N_11836,N_10497);
xnor U17242 (N_17242,N_13162,N_14679);
nand U17243 (N_17243,N_11338,N_12673);
nand U17244 (N_17244,N_12091,N_10112);
or U17245 (N_17245,N_13266,N_11597);
nor U17246 (N_17246,N_11722,N_13932);
nand U17247 (N_17247,N_14578,N_14360);
or U17248 (N_17248,N_12934,N_11720);
and U17249 (N_17249,N_14357,N_12545);
nor U17250 (N_17250,N_12227,N_12424);
nand U17251 (N_17251,N_11491,N_10466);
nor U17252 (N_17252,N_11553,N_11382);
or U17253 (N_17253,N_12876,N_10906);
nor U17254 (N_17254,N_12298,N_11202);
and U17255 (N_17255,N_13564,N_14456);
or U17256 (N_17256,N_10513,N_11075);
xnor U17257 (N_17257,N_13941,N_12563);
nand U17258 (N_17258,N_12093,N_13168);
nand U17259 (N_17259,N_12012,N_14823);
nor U17260 (N_17260,N_13626,N_14101);
nand U17261 (N_17261,N_10171,N_13346);
or U17262 (N_17262,N_12867,N_10925);
and U17263 (N_17263,N_13790,N_14921);
or U17264 (N_17264,N_11704,N_10574);
or U17265 (N_17265,N_14828,N_11412);
or U17266 (N_17266,N_10089,N_11165);
xor U17267 (N_17267,N_12241,N_14451);
and U17268 (N_17268,N_13774,N_10093);
xor U17269 (N_17269,N_14529,N_10749);
nand U17270 (N_17270,N_10403,N_12659);
or U17271 (N_17271,N_10344,N_14137);
or U17272 (N_17272,N_13969,N_11208);
xnor U17273 (N_17273,N_13068,N_14677);
nand U17274 (N_17274,N_14087,N_11877);
xor U17275 (N_17275,N_13298,N_10856);
nor U17276 (N_17276,N_14610,N_12069);
nand U17277 (N_17277,N_12894,N_11842);
nor U17278 (N_17278,N_13495,N_10409);
nand U17279 (N_17279,N_10239,N_14674);
nor U17280 (N_17280,N_12555,N_13121);
and U17281 (N_17281,N_11012,N_11091);
nand U17282 (N_17282,N_11084,N_12118);
or U17283 (N_17283,N_13511,N_14386);
xor U17284 (N_17284,N_14022,N_13030);
nand U17285 (N_17285,N_11268,N_12154);
xnor U17286 (N_17286,N_12564,N_12769);
xor U17287 (N_17287,N_10875,N_11124);
nand U17288 (N_17288,N_13284,N_12509);
nand U17289 (N_17289,N_13952,N_11112);
and U17290 (N_17290,N_14290,N_13362);
and U17291 (N_17291,N_10088,N_11254);
nor U17292 (N_17292,N_10778,N_12362);
and U17293 (N_17293,N_11037,N_14173);
or U17294 (N_17294,N_10920,N_10125);
nor U17295 (N_17295,N_10121,N_10438);
nand U17296 (N_17296,N_14112,N_13055);
nand U17297 (N_17297,N_13854,N_10105);
and U17298 (N_17298,N_12547,N_14270);
nand U17299 (N_17299,N_12863,N_11783);
nand U17300 (N_17300,N_13898,N_10846);
and U17301 (N_17301,N_10718,N_10346);
or U17302 (N_17302,N_12664,N_14162);
and U17303 (N_17303,N_12149,N_11153);
and U17304 (N_17304,N_11357,N_13628);
nand U17305 (N_17305,N_10557,N_11760);
or U17306 (N_17306,N_11218,N_13747);
nand U17307 (N_17307,N_13955,N_14595);
xor U17308 (N_17308,N_10874,N_13112);
nand U17309 (N_17309,N_10682,N_11259);
and U17310 (N_17310,N_10713,N_10079);
and U17311 (N_17311,N_14032,N_14667);
xor U17312 (N_17312,N_14639,N_14338);
xor U17313 (N_17313,N_10503,N_12978);
xnor U17314 (N_17314,N_11655,N_13317);
xor U17315 (N_17315,N_14614,N_12203);
and U17316 (N_17316,N_14808,N_13827);
nor U17317 (N_17317,N_14642,N_10876);
or U17318 (N_17318,N_12785,N_13507);
nand U17319 (N_17319,N_10861,N_14242);
or U17320 (N_17320,N_14512,N_11018);
or U17321 (N_17321,N_12609,N_13946);
xnor U17322 (N_17322,N_11447,N_12548);
xor U17323 (N_17323,N_12181,N_12090);
xor U17324 (N_17324,N_14940,N_12819);
and U17325 (N_17325,N_11521,N_11373);
and U17326 (N_17326,N_10550,N_10709);
nand U17327 (N_17327,N_12879,N_11032);
nor U17328 (N_17328,N_12816,N_14431);
and U17329 (N_17329,N_10164,N_10457);
nor U17330 (N_17330,N_13945,N_13449);
or U17331 (N_17331,N_14555,N_12629);
and U17332 (N_17332,N_10200,N_10934);
or U17333 (N_17333,N_10182,N_14659);
xor U17334 (N_17334,N_11841,N_10176);
and U17335 (N_17335,N_13869,N_10177);
nor U17336 (N_17336,N_14671,N_11191);
xor U17337 (N_17337,N_14869,N_11255);
nand U17338 (N_17338,N_11987,N_14758);
nor U17339 (N_17339,N_12633,N_10533);
or U17340 (N_17340,N_10609,N_13532);
and U17341 (N_17341,N_12092,N_10321);
xor U17342 (N_17342,N_10748,N_14053);
xnor U17343 (N_17343,N_10158,N_13783);
or U17344 (N_17344,N_13853,N_10433);
or U17345 (N_17345,N_11327,N_14212);
xor U17346 (N_17346,N_10669,N_10831);
or U17347 (N_17347,N_10559,N_12464);
nor U17348 (N_17348,N_13073,N_12591);
and U17349 (N_17349,N_10707,N_11571);
xor U17350 (N_17350,N_14492,N_12351);
nor U17351 (N_17351,N_10302,N_12650);
or U17352 (N_17352,N_10726,N_11174);
nand U17353 (N_17353,N_14864,N_13562);
or U17354 (N_17354,N_13006,N_12228);
nor U17355 (N_17355,N_10377,N_13542);
or U17356 (N_17356,N_13695,N_12427);
xnor U17357 (N_17357,N_13750,N_13008);
nor U17358 (N_17358,N_12124,N_14591);
or U17359 (N_17359,N_10570,N_13533);
nor U17360 (N_17360,N_14703,N_13755);
or U17361 (N_17361,N_12449,N_10572);
xnor U17362 (N_17362,N_10204,N_14518);
or U17363 (N_17363,N_11872,N_10385);
or U17364 (N_17364,N_13405,N_12671);
nor U17365 (N_17365,N_11510,N_14231);
nor U17366 (N_17366,N_10881,N_14931);
or U17367 (N_17367,N_13944,N_14933);
or U17368 (N_17368,N_13293,N_10113);
or U17369 (N_17369,N_10060,N_10678);
and U17370 (N_17370,N_10803,N_11074);
xor U17371 (N_17371,N_12953,N_11162);
nor U17372 (N_17372,N_14672,N_12156);
nor U17373 (N_17373,N_11231,N_13770);
and U17374 (N_17374,N_12275,N_11966);
nand U17375 (N_17375,N_12303,N_12459);
and U17376 (N_17376,N_14370,N_14945);
and U17377 (N_17377,N_14552,N_13310);
nand U17378 (N_17378,N_14056,N_12215);
nand U17379 (N_17379,N_12440,N_10370);
and U17380 (N_17380,N_13040,N_14260);
nand U17381 (N_17381,N_13189,N_11869);
nand U17382 (N_17382,N_14289,N_11233);
or U17383 (N_17383,N_12574,N_10062);
nand U17384 (N_17384,N_10584,N_11434);
xnor U17385 (N_17385,N_13561,N_13645);
or U17386 (N_17386,N_12518,N_11216);
xnor U17387 (N_17387,N_10037,N_10203);
or U17388 (N_17388,N_11418,N_14793);
and U17389 (N_17389,N_10676,N_12246);
nand U17390 (N_17390,N_10783,N_12970);
xor U17391 (N_17391,N_12772,N_13327);
and U17392 (N_17392,N_13551,N_11060);
xnor U17393 (N_17393,N_14084,N_13799);
xnor U17394 (N_17394,N_13865,N_12173);
and U17395 (N_17395,N_14174,N_12435);
and U17396 (N_17396,N_12553,N_12836);
and U17397 (N_17397,N_11830,N_11752);
xnor U17398 (N_17398,N_12267,N_14291);
nand U17399 (N_17399,N_11487,N_13872);
and U17400 (N_17400,N_13581,N_10007);
nand U17401 (N_17401,N_11792,N_11981);
nor U17402 (N_17402,N_10665,N_10005);
or U17403 (N_17403,N_11678,N_10727);
or U17404 (N_17404,N_13508,N_13891);
nor U17405 (N_17405,N_13080,N_14938);
xnor U17406 (N_17406,N_13880,N_13985);
and U17407 (N_17407,N_14042,N_13503);
xor U17408 (N_17408,N_10937,N_12905);
nand U17409 (N_17409,N_10209,N_13998);
nor U17410 (N_17410,N_13972,N_11450);
nor U17411 (N_17411,N_11608,N_12187);
xnor U17412 (N_17412,N_12538,N_10487);
or U17413 (N_17413,N_14825,N_11082);
xnor U17414 (N_17414,N_13289,N_13845);
or U17415 (N_17415,N_12169,N_14167);
nor U17416 (N_17416,N_13024,N_14037);
nor U17417 (N_17417,N_14544,N_14998);
or U17418 (N_17418,N_12332,N_10166);
nor U17419 (N_17419,N_12072,N_11065);
or U17420 (N_17420,N_12974,N_12968);
xor U17421 (N_17421,N_14937,N_13754);
or U17422 (N_17422,N_13455,N_12480);
and U17423 (N_17423,N_11504,N_13578);
nor U17424 (N_17424,N_13571,N_14334);
and U17425 (N_17425,N_12344,N_13999);
xor U17426 (N_17426,N_11730,N_12690);
nor U17427 (N_17427,N_10826,N_11970);
nor U17428 (N_17428,N_12117,N_10830);
nor U17429 (N_17429,N_14423,N_10692);
or U17430 (N_17430,N_10045,N_11030);
xor U17431 (N_17431,N_13684,N_13246);
xnor U17432 (N_17432,N_14356,N_14114);
xnor U17433 (N_17433,N_12325,N_13300);
nor U17434 (N_17434,N_14593,N_13724);
nor U17435 (N_17435,N_14771,N_12572);
nor U17436 (N_17436,N_14443,N_14956);
and U17437 (N_17437,N_13208,N_12839);
xnor U17438 (N_17438,N_10504,N_11333);
or U17439 (N_17439,N_14957,N_14365);
xnor U17440 (N_17440,N_12159,N_13519);
and U17441 (N_17441,N_14636,N_11238);
or U17442 (N_17442,N_11858,N_12063);
and U17443 (N_17443,N_12099,N_10746);
nor U17444 (N_17444,N_12598,N_10654);
nand U17445 (N_17445,N_10355,N_11500);
or U17446 (N_17446,N_12195,N_11351);
xnor U17447 (N_17447,N_13716,N_14801);
and U17448 (N_17448,N_11262,N_13365);
nand U17449 (N_17449,N_14698,N_12663);
or U17450 (N_17450,N_13323,N_11243);
and U17451 (N_17451,N_13620,N_11320);
or U17452 (N_17452,N_11034,N_13706);
or U17453 (N_17453,N_12198,N_13560);
xor U17454 (N_17454,N_13347,N_13884);
nand U17455 (N_17455,N_10414,N_14880);
and U17456 (N_17456,N_13612,N_14400);
nor U17457 (N_17457,N_11209,N_11594);
or U17458 (N_17458,N_13748,N_14635);
xor U17459 (N_17459,N_14584,N_12558);
nor U17460 (N_17460,N_13200,N_14015);
nor U17461 (N_17461,N_13963,N_10845);
nor U17462 (N_17462,N_12394,N_10724);
xor U17463 (N_17463,N_13658,N_11954);
and U17464 (N_17464,N_13478,N_10369);
and U17465 (N_17465,N_13893,N_14350);
and U17466 (N_17466,N_12386,N_14034);
or U17467 (N_17467,N_13699,N_13948);
nor U17468 (N_17468,N_14149,N_10228);
nor U17469 (N_17469,N_13650,N_10710);
xnor U17470 (N_17470,N_13526,N_14553);
or U17471 (N_17471,N_10670,N_10977);
and U17472 (N_17472,N_11918,N_10298);
or U17473 (N_17473,N_11077,N_14062);
or U17474 (N_17474,N_13668,N_13183);
xor U17475 (N_17475,N_11284,N_11120);
and U17476 (N_17476,N_11756,N_12290);
and U17477 (N_17477,N_11999,N_10886);
xor U17478 (N_17478,N_14098,N_11006);
nor U17479 (N_17479,N_14250,N_11099);
or U17480 (N_17480,N_13506,N_10788);
nand U17481 (N_17481,N_14633,N_14807);
and U17482 (N_17482,N_10526,N_10375);
or U17483 (N_17483,N_12034,N_11823);
nor U17484 (N_17484,N_10295,N_12988);
xnor U17485 (N_17485,N_14896,N_11972);
xnor U17486 (N_17486,N_14968,N_13579);
nor U17487 (N_17487,N_13602,N_14904);
and U17488 (N_17488,N_14283,N_12824);
and U17489 (N_17489,N_11761,N_12814);
nor U17490 (N_17490,N_13789,N_13038);
nor U17491 (N_17491,N_10736,N_14692);
or U17492 (N_17492,N_14500,N_10245);
or U17493 (N_17493,N_10148,N_10828);
nand U17494 (N_17494,N_12933,N_14148);
and U17495 (N_17495,N_13017,N_12770);
nand U17496 (N_17496,N_14953,N_13878);
and U17497 (N_17497,N_13912,N_10488);
nand U17498 (N_17498,N_13304,N_11377);
nand U17499 (N_17499,N_13734,N_14519);
xnor U17500 (N_17500,N_13833,N_12515);
nor U17501 (N_17501,N_14219,N_10319);
nor U17502 (N_17502,N_13428,N_11157);
nor U17503 (N_17503,N_11376,N_14049);
xnor U17504 (N_17504,N_11495,N_11282);
and U17505 (N_17505,N_11623,N_12397);
or U17506 (N_17506,N_14889,N_10297);
nor U17507 (N_17507,N_10726,N_12403);
xnor U17508 (N_17508,N_10050,N_13949);
or U17509 (N_17509,N_11181,N_14593);
or U17510 (N_17510,N_14866,N_12040);
nand U17511 (N_17511,N_13857,N_14633);
xnor U17512 (N_17512,N_11583,N_14426);
xor U17513 (N_17513,N_11969,N_11219);
xnor U17514 (N_17514,N_11087,N_12542);
xor U17515 (N_17515,N_11295,N_11731);
and U17516 (N_17516,N_10676,N_12694);
and U17517 (N_17517,N_10891,N_14634);
xor U17518 (N_17518,N_10054,N_10529);
xor U17519 (N_17519,N_14438,N_13444);
and U17520 (N_17520,N_12065,N_11885);
nand U17521 (N_17521,N_13507,N_10951);
nor U17522 (N_17522,N_13021,N_10016);
and U17523 (N_17523,N_13197,N_11000);
and U17524 (N_17524,N_11949,N_14974);
or U17525 (N_17525,N_12735,N_11800);
and U17526 (N_17526,N_11598,N_11862);
xor U17527 (N_17527,N_12437,N_10605);
xnor U17528 (N_17528,N_10833,N_11555);
xor U17529 (N_17529,N_14172,N_12479);
and U17530 (N_17530,N_14476,N_11445);
nand U17531 (N_17531,N_13935,N_11186);
and U17532 (N_17532,N_13918,N_13421);
or U17533 (N_17533,N_12288,N_12972);
and U17534 (N_17534,N_10842,N_12395);
or U17535 (N_17535,N_10154,N_12606);
and U17536 (N_17536,N_10366,N_11871);
and U17537 (N_17537,N_11341,N_11850);
nor U17538 (N_17538,N_10495,N_11613);
nor U17539 (N_17539,N_11889,N_14623);
and U17540 (N_17540,N_14923,N_14204);
nand U17541 (N_17541,N_10932,N_10265);
nor U17542 (N_17542,N_12652,N_13865);
xor U17543 (N_17543,N_11849,N_11566);
nand U17544 (N_17544,N_11921,N_11496);
and U17545 (N_17545,N_10211,N_10220);
nor U17546 (N_17546,N_10588,N_11542);
and U17547 (N_17547,N_14509,N_12190);
and U17548 (N_17548,N_11729,N_11461);
nor U17549 (N_17549,N_10531,N_11184);
nor U17550 (N_17550,N_13634,N_12464);
nor U17551 (N_17551,N_10982,N_10720);
nor U17552 (N_17552,N_13647,N_14912);
xor U17553 (N_17553,N_11194,N_14780);
nor U17554 (N_17554,N_12848,N_14836);
or U17555 (N_17555,N_13078,N_11353);
nor U17556 (N_17556,N_14057,N_10178);
nand U17557 (N_17557,N_13206,N_11356);
and U17558 (N_17558,N_12164,N_11591);
nand U17559 (N_17559,N_11036,N_14776);
and U17560 (N_17560,N_12682,N_14216);
and U17561 (N_17561,N_12287,N_13495);
xor U17562 (N_17562,N_13147,N_10783);
xnor U17563 (N_17563,N_13964,N_11752);
xor U17564 (N_17564,N_13182,N_11562);
nor U17565 (N_17565,N_11847,N_12228);
nand U17566 (N_17566,N_13751,N_10968);
or U17567 (N_17567,N_10659,N_14826);
or U17568 (N_17568,N_13900,N_11390);
or U17569 (N_17569,N_10263,N_11390);
nor U17570 (N_17570,N_10391,N_11935);
and U17571 (N_17571,N_14406,N_12431);
xor U17572 (N_17572,N_12608,N_13156);
and U17573 (N_17573,N_11451,N_11259);
or U17574 (N_17574,N_11761,N_12173);
nor U17575 (N_17575,N_10128,N_14949);
nand U17576 (N_17576,N_10770,N_13421);
nor U17577 (N_17577,N_12730,N_13154);
nand U17578 (N_17578,N_11743,N_14065);
nand U17579 (N_17579,N_13592,N_14791);
nor U17580 (N_17580,N_13904,N_14107);
nor U17581 (N_17581,N_11249,N_11478);
xnor U17582 (N_17582,N_14651,N_14966);
nor U17583 (N_17583,N_10193,N_12619);
xor U17584 (N_17584,N_10096,N_14143);
or U17585 (N_17585,N_10371,N_11911);
and U17586 (N_17586,N_11909,N_12802);
and U17587 (N_17587,N_13412,N_10650);
nor U17588 (N_17588,N_12765,N_14878);
nand U17589 (N_17589,N_14671,N_14255);
or U17590 (N_17590,N_14554,N_14249);
or U17591 (N_17591,N_12520,N_12557);
or U17592 (N_17592,N_13588,N_14825);
xnor U17593 (N_17593,N_12324,N_12125);
nor U17594 (N_17594,N_10184,N_14672);
nor U17595 (N_17595,N_10108,N_13421);
xor U17596 (N_17596,N_14153,N_12303);
or U17597 (N_17597,N_11007,N_14798);
and U17598 (N_17598,N_10333,N_14140);
or U17599 (N_17599,N_12544,N_10078);
nand U17600 (N_17600,N_12117,N_11454);
nor U17601 (N_17601,N_14137,N_11089);
nand U17602 (N_17602,N_10832,N_14101);
and U17603 (N_17603,N_14729,N_14952);
xnor U17604 (N_17604,N_12720,N_10340);
and U17605 (N_17605,N_12500,N_11934);
xor U17606 (N_17606,N_10251,N_11286);
nor U17607 (N_17607,N_11745,N_11639);
nand U17608 (N_17608,N_11636,N_14838);
nor U17609 (N_17609,N_14005,N_13898);
nor U17610 (N_17610,N_10896,N_11538);
xnor U17611 (N_17611,N_10676,N_14569);
and U17612 (N_17612,N_10038,N_14703);
nand U17613 (N_17613,N_10483,N_14258);
xor U17614 (N_17614,N_14728,N_13201);
nand U17615 (N_17615,N_12118,N_10938);
xor U17616 (N_17616,N_13131,N_12799);
or U17617 (N_17617,N_14305,N_12555);
and U17618 (N_17618,N_11124,N_10509);
xor U17619 (N_17619,N_10472,N_11134);
or U17620 (N_17620,N_11356,N_12716);
or U17621 (N_17621,N_10193,N_11485);
and U17622 (N_17622,N_10809,N_13046);
xor U17623 (N_17623,N_13729,N_12302);
nand U17624 (N_17624,N_10343,N_12544);
or U17625 (N_17625,N_12317,N_10701);
or U17626 (N_17626,N_12501,N_11316);
or U17627 (N_17627,N_13425,N_12867);
xor U17628 (N_17628,N_14381,N_14228);
and U17629 (N_17629,N_12017,N_10377);
nand U17630 (N_17630,N_12679,N_14781);
or U17631 (N_17631,N_13613,N_11832);
or U17632 (N_17632,N_13442,N_11858);
or U17633 (N_17633,N_14317,N_14118);
nand U17634 (N_17634,N_11719,N_10583);
nor U17635 (N_17635,N_14337,N_13115);
xor U17636 (N_17636,N_14765,N_10436);
xor U17637 (N_17637,N_11730,N_11359);
nor U17638 (N_17638,N_13966,N_13098);
and U17639 (N_17639,N_10401,N_10213);
and U17640 (N_17640,N_10132,N_10520);
and U17641 (N_17641,N_14075,N_12019);
and U17642 (N_17642,N_13916,N_13503);
nor U17643 (N_17643,N_13809,N_13837);
nand U17644 (N_17644,N_14828,N_12189);
xor U17645 (N_17645,N_14759,N_11475);
nor U17646 (N_17646,N_13588,N_11123);
nand U17647 (N_17647,N_10041,N_10564);
and U17648 (N_17648,N_14022,N_10294);
nand U17649 (N_17649,N_11086,N_10737);
or U17650 (N_17650,N_14616,N_10164);
or U17651 (N_17651,N_10695,N_12384);
nand U17652 (N_17652,N_10289,N_14659);
or U17653 (N_17653,N_14955,N_10601);
xor U17654 (N_17654,N_12871,N_14215);
or U17655 (N_17655,N_14965,N_10429);
or U17656 (N_17656,N_13633,N_13347);
and U17657 (N_17657,N_13811,N_13906);
nor U17658 (N_17658,N_13334,N_12826);
xnor U17659 (N_17659,N_13492,N_13181);
nor U17660 (N_17660,N_11360,N_13129);
nor U17661 (N_17661,N_12799,N_10697);
xnor U17662 (N_17662,N_10564,N_10339);
nor U17663 (N_17663,N_12324,N_11448);
or U17664 (N_17664,N_11073,N_10722);
xor U17665 (N_17665,N_10436,N_11856);
or U17666 (N_17666,N_12117,N_10356);
or U17667 (N_17667,N_14733,N_12469);
or U17668 (N_17668,N_10363,N_14386);
or U17669 (N_17669,N_13573,N_10140);
or U17670 (N_17670,N_12112,N_11278);
and U17671 (N_17671,N_10894,N_11348);
nor U17672 (N_17672,N_10637,N_10056);
xnor U17673 (N_17673,N_10871,N_11030);
xnor U17674 (N_17674,N_13646,N_13076);
xnor U17675 (N_17675,N_14623,N_13399);
xor U17676 (N_17676,N_10294,N_11314);
nor U17677 (N_17677,N_12289,N_14836);
nor U17678 (N_17678,N_11314,N_14216);
and U17679 (N_17679,N_10961,N_10504);
or U17680 (N_17680,N_11032,N_12769);
xor U17681 (N_17681,N_13211,N_11075);
and U17682 (N_17682,N_11639,N_13840);
nor U17683 (N_17683,N_11571,N_14551);
and U17684 (N_17684,N_11710,N_10985);
xor U17685 (N_17685,N_14138,N_13379);
nand U17686 (N_17686,N_10040,N_11179);
and U17687 (N_17687,N_14141,N_11725);
nor U17688 (N_17688,N_12766,N_14064);
and U17689 (N_17689,N_11208,N_10868);
or U17690 (N_17690,N_12916,N_10549);
or U17691 (N_17691,N_13434,N_13000);
nand U17692 (N_17692,N_10298,N_13952);
or U17693 (N_17693,N_12581,N_14682);
nor U17694 (N_17694,N_13728,N_12450);
nand U17695 (N_17695,N_13776,N_10850);
xnor U17696 (N_17696,N_12668,N_10488);
nand U17697 (N_17697,N_14084,N_10107);
nor U17698 (N_17698,N_11748,N_11461);
and U17699 (N_17699,N_13950,N_14730);
nor U17700 (N_17700,N_13277,N_13670);
or U17701 (N_17701,N_14315,N_11122);
xor U17702 (N_17702,N_14580,N_11265);
xnor U17703 (N_17703,N_12299,N_14559);
nand U17704 (N_17704,N_14112,N_11119);
nand U17705 (N_17705,N_12330,N_10304);
nor U17706 (N_17706,N_13457,N_12822);
nor U17707 (N_17707,N_14035,N_12183);
xor U17708 (N_17708,N_12676,N_14454);
xor U17709 (N_17709,N_13711,N_12488);
nor U17710 (N_17710,N_12920,N_10215);
nand U17711 (N_17711,N_13099,N_14134);
xor U17712 (N_17712,N_12114,N_11956);
nand U17713 (N_17713,N_11563,N_11181);
or U17714 (N_17714,N_13760,N_10129);
xnor U17715 (N_17715,N_11733,N_10685);
nand U17716 (N_17716,N_11818,N_13571);
and U17717 (N_17717,N_14855,N_14549);
nand U17718 (N_17718,N_10351,N_11454);
xor U17719 (N_17719,N_11832,N_12380);
nor U17720 (N_17720,N_13503,N_11116);
nand U17721 (N_17721,N_14892,N_14029);
nand U17722 (N_17722,N_14126,N_10615);
nand U17723 (N_17723,N_10481,N_12303);
nor U17724 (N_17724,N_14310,N_14530);
and U17725 (N_17725,N_12380,N_12586);
xor U17726 (N_17726,N_14448,N_11022);
nand U17727 (N_17727,N_11079,N_12788);
and U17728 (N_17728,N_14193,N_10313);
or U17729 (N_17729,N_11479,N_11624);
xnor U17730 (N_17730,N_13954,N_10186);
nor U17731 (N_17731,N_14404,N_14576);
nand U17732 (N_17732,N_10922,N_10405);
nand U17733 (N_17733,N_13092,N_11679);
nor U17734 (N_17734,N_10331,N_12508);
nand U17735 (N_17735,N_13212,N_12375);
and U17736 (N_17736,N_11153,N_11274);
and U17737 (N_17737,N_11990,N_10671);
and U17738 (N_17738,N_14635,N_12586);
and U17739 (N_17739,N_14627,N_14635);
nand U17740 (N_17740,N_10612,N_13055);
and U17741 (N_17741,N_11558,N_11276);
and U17742 (N_17742,N_12835,N_10333);
or U17743 (N_17743,N_11536,N_13100);
nor U17744 (N_17744,N_10388,N_13403);
and U17745 (N_17745,N_13938,N_14928);
or U17746 (N_17746,N_10079,N_12385);
and U17747 (N_17747,N_11352,N_14188);
xor U17748 (N_17748,N_11508,N_13547);
nand U17749 (N_17749,N_13089,N_11803);
nand U17750 (N_17750,N_13453,N_11867);
xor U17751 (N_17751,N_12005,N_14524);
nand U17752 (N_17752,N_14518,N_12861);
or U17753 (N_17753,N_13345,N_10751);
and U17754 (N_17754,N_14387,N_11621);
nand U17755 (N_17755,N_13323,N_11480);
nor U17756 (N_17756,N_14803,N_14389);
or U17757 (N_17757,N_10288,N_12500);
xor U17758 (N_17758,N_10814,N_14558);
xor U17759 (N_17759,N_12152,N_13833);
and U17760 (N_17760,N_10488,N_11778);
and U17761 (N_17761,N_12322,N_14950);
and U17762 (N_17762,N_13901,N_13988);
nand U17763 (N_17763,N_12054,N_12521);
xnor U17764 (N_17764,N_13730,N_13888);
nor U17765 (N_17765,N_11949,N_11274);
and U17766 (N_17766,N_11469,N_12723);
nand U17767 (N_17767,N_14388,N_13401);
xnor U17768 (N_17768,N_10855,N_11635);
xnor U17769 (N_17769,N_11354,N_11562);
xor U17770 (N_17770,N_11687,N_12470);
nand U17771 (N_17771,N_10446,N_13795);
or U17772 (N_17772,N_13280,N_10867);
and U17773 (N_17773,N_11971,N_11322);
and U17774 (N_17774,N_10824,N_12771);
xnor U17775 (N_17775,N_12923,N_11667);
xor U17776 (N_17776,N_10848,N_10284);
nand U17777 (N_17777,N_10498,N_13844);
and U17778 (N_17778,N_10441,N_12284);
nor U17779 (N_17779,N_11610,N_14645);
xnor U17780 (N_17780,N_13049,N_11893);
xor U17781 (N_17781,N_14237,N_13883);
or U17782 (N_17782,N_12187,N_12125);
nor U17783 (N_17783,N_13456,N_10040);
and U17784 (N_17784,N_12413,N_14079);
xnor U17785 (N_17785,N_11234,N_11875);
nand U17786 (N_17786,N_10156,N_12187);
and U17787 (N_17787,N_10887,N_12918);
or U17788 (N_17788,N_12079,N_10526);
and U17789 (N_17789,N_12369,N_14747);
xor U17790 (N_17790,N_12324,N_10514);
or U17791 (N_17791,N_14090,N_12380);
and U17792 (N_17792,N_14045,N_14941);
and U17793 (N_17793,N_10353,N_11880);
nor U17794 (N_17794,N_14357,N_10632);
or U17795 (N_17795,N_14820,N_12486);
xnor U17796 (N_17796,N_14108,N_10409);
and U17797 (N_17797,N_12344,N_10842);
xnor U17798 (N_17798,N_13659,N_10119);
and U17799 (N_17799,N_11256,N_13951);
nand U17800 (N_17800,N_10590,N_13150);
xor U17801 (N_17801,N_13712,N_11815);
or U17802 (N_17802,N_10268,N_12106);
or U17803 (N_17803,N_13881,N_12029);
xnor U17804 (N_17804,N_10865,N_13967);
and U17805 (N_17805,N_13259,N_11455);
and U17806 (N_17806,N_11081,N_10704);
and U17807 (N_17807,N_12356,N_13846);
nand U17808 (N_17808,N_12645,N_13708);
xor U17809 (N_17809,N_11058,N_14581);
and U17810 (N_17810,N_11578,N_12468);
and U17811 (N_17811,N_12296,N_14418);
or U17812 (N_17812,N_13802,N_11058);
xnor U17813 (N_17813,N_13561,N_14713);
nor U17814 (N_17814,N_13937,N_11402);
nor U17815 (N_17815,N_10487,N_11754);
or U17816 (N_17816,N_12501,N_11523);
and U17817 (N_17817,N_10876,N_10277);
or U17818 (N_17818,N_14765,N_11249);
or U17819 (N_17819,N_14464,N_10843);
and U17820 (N_17820,N_10074,N_14808);
or U17821 (N_17821,N_11241,N_14194);
xor U17822 (N_17822,N_14136,N_11688);
or U17823 (N_17823,N_10929,N_13395);
nor U17824 (N_17824,N_13641,N_10536);
nand U17825 (N_17825,N_14738,N_14672);
or U17826 (N_17826,N_14502,N_10240);
xor U17827 (N_17827,N_11889,N_13541);
nor U17828 (N_17828,N_11557,N_12905);
xnor U17829 (N_17829,N_11695,N_11395);
or U17830 (N_17830,N_14994,N_14828);
and U17831 (N_17831,N_13436,N_12085);
nor U17832 (N_17832,N_10056,N_10806);
or U17833 (N_17833,N_14256,N_14614);
or U17834 (N_17834,N_12107,N_13696);
or U17835 (N_17835,N_14912,N_14543);
and U17836 (N_17836,N_14109,N_10983);
xor U17837 (N_17837,N_13670,N_14712);
and U17838 (N_17838,N_11363,N_13831);
or U17839 (N_17839,N_10780,N_12783);
and U17840 (N_17840,N_13896,N_10174);
and U17841 (N_17841,N_11924,N_14110);
xor U17842 (N_17842,N_13148,N_14088);
xor U17843 (N_17843,N_13711,N_12841);
nand U17844 (N_17844,N_14129,N_14942);
nand U17845 (N_17845,N_12934,N_11294);
and U17846 (N_17846,N_14164,N_11561);
or U17847 (N_17847,N_12760,N_11118);
xnor U17848 (N_17848,N_12181,N_12060);
xnor U17849 (N_17849,N_14977,N_14628);
nor U17850 (N_17850,N_12905,N_12924);
nor U17851 (N_17851,N_14569,N_11915);
or U17852 (N_17852,N_11429,N_10878);
xnor U17853 (N_17853,N_12467,N_12990);
or U17854 (N_17854,N_12228,N_10884);
nand U17855 (N_17855,N_10208,N_14846);
xor U17856 (N_17856,N_13944,N_13817);
or U17857 (N_17857,N_12884,N_14148);
and U17858 (N_17858,N_10291,N_10880);
or U17859 (N_17859,N_12928,N_12707);
nor U17860 (N_17860,N_10192,N_14054);
or U17861 (N_17861,N_12486,N_13167);
and U17862 (N_17862,N_10196,N_12496);
nand U17863 (N_17863,N_10155,N_14054);
or U17864 (N_17864,N_13199,N_14387);
nand U17865 (N_17865,N_11485,N_13081);
and U17866 (N_17866,N_10533,N_12233);
and U17867 (N_17867,N_10550,N_11632);
nand U17868 (N_17868,N_13058,N_10180);
xnor U17869 (N_17869,N_12568,N_11768);
xor U17870 (N_17870,N_14971,N_13443);
and U17871 (N_17871,N_10141,N_14089);
and U17872 (N_17872,N_11191,N_14230);
xor U17873 (N_17873,N_11482,N_11069);
or U17874 (N_17874,N_12951,N_10592);
nand U17875 (N_17875,N_11249,N_10610);
nor U17876 (N_17876,N_10233,N_13999);
xor U17877 (N_17877,N_11857,N_14796);
nand U17878 (N_17878,N_12815,N_10862);
and U17879 (N_17879,N_12436,N_13624);
or U17880 (N_17880,N_13576,N_13950);
nor U17881 (N_17881,N_10123,N_11821);
or U17882 (N_17882,N_11336,N_12453);
nor U17883 (N_17883,N_13943,N_13848);
nor U17884 (N_17884,N_14255,N_11467);
and U17885 (N_17885,N_10304,N_10211);
xnor U17886 (N_17886,N_11372,N_13183);
and U17887 (N_17887,N_11350,N_14520);
nor U17888 (N_17888,N_10483,N_11048);
or U17889 (N_17889,N_14717,N_14776);
and U17890 (N_17890,N_11571,N_14911);
and U17891 (N_17891,N_13567,N_11092);
xor U17892 (N_17892,N_10142,N_11277);
nand U17893 (N_17893,N_10567,N_11728);
nor U17894 (N_17894,N_10566,N_10548);
nand U17895 (N_17895,N_13289,N_13037);
and U17896 (N_17896,N_13974,N_12081);
and U17897 (N_17897,N_14252,N_11192);
nand U17898 (N_17898,N_13076,N_11348);
nand U17899 (N_17899,N_12702,N_13858);
xnor U17900 (N_17900,N_12742,N_14346);
or U17901 (N_17901,N_14031,N_12695);
or U17902 (N_17902,N_11990,N_13402);
and U17903 (N_17903,N_11365,N_11790);
nor U17904 (N_17904,N_11065,N_11882);
xnor U17905 (N_17905,N_12100,N_14703);
nor U17906 (N_17906,N_14660,N_12498);
nor U17907 (N_17907,N_12370,N_11735);
nor U17908 (N_17908,N_14234,N_11726);
nor U17909 (N_17909,N_12564,N_11976);
nand U17910 (N_17910,N_14144,N_14973);
and U17911 (N_17911,N_12504,N_13964);
and U17912 (N_17912,N_12296,N_11882);
xor U17913 (N_17913,N_12432,N_10496);
and U17914 (N_17914,N_10011,N_14703);
or U17915 (N_17915,N_11736,N_11624);
xor U17916 (N_17916,N_13277,N_13598);
nand U17917 (N_17917,N_12963,N_11738);
nor U17918 (N_17918,N_14586,N_11536);
and U17919 (N_17919,N_14602,N_13087);
or U17920 (N_17920,N_10363,N_13052);
nor U17921 (N_17921,N_11334,N_10263);
xor U17922 (N_17922,N_13270,N_12210);
and U17923 (N_17923,N_12895,N_14088);
nor U17924 (N_17924,N_12686,N_12430);
xor U17925 (N_17925,N_12816,N_13522);
nand U17926 (N_17926,N_11437,N_11818);
and U17927 (N_17927,N_11348,N_14536);
nor U17928 (N_17928,N_14934,N_12622);
or U17929 (N_17929,N_14092,N_11473);
xnor U17930 (N_17930,N_13643,N_12107);
xor U17931 (N_17931,N_11256,N_14702);
and U17932 (N_17932,N_10740,N_12826);
and U17933 (N_17933,N_10029,N_12834);
nand U17934 (N_17934,N_13746,N_12660);
and U17935 (N_17935,N_13338,N_14460);
nor U17936 (N_17936,N_12238,N_13012);
xor U17937 (N_17937,N_11937,N_13102);
nand U17938 (N_17938,N_11275,N_10841);
nand U17939 (N_17939,N_12052,N_10112);
nor U17940 (N_17940,N_13889,N_13119);
xnor U17941 (N_17941,N_10171,N_11717);
or U17942 (N_17942,N_12391,N_12555);
or U17943 (N_17943,N_14707,N_12569);
xor U17944 (N_17944,N_12512,N_10562);
xor U17945 (N_17945,N_12570,N_12063);
or U17946 (N_17946,N_11051,N_12638);
xor U17947 (N_17947,N_11543,N_14227);
xnor U17948 (N_17948,N_11059,N_12759);
xnor U17949 (N_17949,N_14762,N_10261);
or U17950 (N_17950,N_14745,N_10026);
xor U17951 (N_17951,N_13409,N_12873);
and U17952 (N_17952,N_11134,N_12056);
or U17953 (N_17953,N_14638,N_10331);
or U17954 (N_17954,N_11015,N_14446);
xnor U17955 (N_17955,N_12980,N_14167);
or U17956 (N_17956,N_11862,N_14763);
nor U17957 (N_17957,N_14334,N_12578);
nand U17958 (N_17958,N_11033,N_13747);
nor U17959 (N_17959,N_11084,N_12836);
and U17960 (N_17960,N_12127,N_13446);
and U17961 (N_17961,N_10081,N_10438);
xor U17962 (N_17962,N_10874,N_14838);
nand U17963 (N_17963,N_12108,N_10469);
xor U17964 (N_17964,N_14965,N_14484);
or U17965 (N_17965,N_11658,N_11737);
xnor U17966 (N_17966,N_10899,N_11344);
or U17967 (N_17967,N_12883,N_11562);
nor U17968 (N_17968,N_14630,N_10444);
nand U17969 (N_17969,N_10389,N_11751);
and U17970 (N_17970,N_14258,N_14329);
and U17971 (N_17971,N_10641,N_11337);
nand U17972 (N_17972,N_12072,N_13975);
xor U17973 (N_17973,N_14702,N_13210);
or U17974 (N_17974,N_14368,N_11621);
xor U17975 (N_17975,N_12657,N_14422);
and U17976 (N_17976,N_11659,N_10995);
nand U17977 (N_17977,N_12562,N_10299);
and U17978 (N_17978,N_11299,N_12758);
or U17979 (N_17979,N_13732,N_13481);
or U17980 (N_17980,N_14594,N_14279);
xor U17981 (N_17981,N_13777,N_14491);
nand U17982 (N_17982,N_14569,N_13144);
nand U17983 (N_17983,N_13733,N_14136);
nand U17984 (N_17984,N_11384,N_10965);
nand U17985 (N_17985,N_12965,N_14610);
and U17986 (N_17986,N_10982,N_11895);
or U17987 (N_17987,N_14360,N_10588);
and U17988 (N_17988,N_12709,N_13069);
nand U17989 (N_17989,N_12493,N_10926);
nand U17990 (N_17990,N_10363,N_13902);
xnor U17991 (N_17991,N_13945,N_13704);
or U17992 (N_17992,N_14081,N_14584);
or U17993 (N_17993,N_11481,N_10698);
and U17994 (N_17994,N_14484,N_10334);
or U17995 (N_17995,N_13232,N_14662);
nor U17996 (N_17996,N_13621,N_11462);
nand U17997 (N_17997,N_14403,N_12707);
or U17998 (N_17998,N_11164,N_14320);
and U17999 (N_17999,N_14028,N_10194);
or U18000 (N_18000,N_13783,N_13916);
xor U18001 (N_18001,N_12236,N_14443);
xor U18002 (N_18002,N_14529,N_14011);
or U18003 (N_18003,N_12932,N_12791);
or U18004 (N_18004,N_11793,N_12276);
nor U18005 (N_18005,N_13416,N_14721);
and U18006 (N_18006,N_10711,N_11065);
nor U18007 (N_18007,N_10212,N_13511);
nor U18008 (N_18008,N_13732,N_14354);
or U18009 (N_18009,N_10878,N_14027);
and U18010 (N_18010,N_12700,N_11137);
or U18011 (N_18011,N_10616,N_12202);
nor U18012 (N_18012,N_10512,N_11231);
or U18013 (N_18013,N_14894,N_12796);
or U18014 (N_18014,N_10742,N_13102);
nand U18015 (N_18015,N_13484,N_10265);
nand U18016 (N_18016,N_12991,N_14983);
nand U18017 (N_18017,N_13808,N_14177);
nor U18018 (N_18018,N_14871,N_13620);
nor U18019 (N_18019,N_10095,N_14894);
and U18020 (N_18020,N_13189,N_14695);
nor U18021 (N_18021,N_12257,N_14064);
or U18022 (N_18022,N_12574,N_11845);
xor U18023 (N_18023,N_13062,N_10817);
or U18024 (N_18024,N_13203,N_10840);
and U18025 (N_18025,N_14343,N_12412);
xor U18026 (N_18026,N_13178,N_13416);
xnor U18027 (N_18027,N_14141,N_10196);
nor U18028 (N_18028,N_13926,N_13370);
and U18029 (N_18029,N_14615,N_10184);
or U18030 (N_18030,N_14538,N_12203);
or U18031 (N_18031,N_12176,N_14439);
nor U18032 (N_18032,N_11072,N_12658);
nor U18033 (N_18033,N_14535,N_13265);
nand U18034 (N_18034,N_13735,N_11234);
xor U18035 (N_18035,N_11918,N_13104);
xnor U18036 (N_18036,N_12461,N_12426);
or U18037 (N_18037,N_12429,N_11885);
nand U18038 (N_18038,N_11352,N_12726);
nand U18039 (N_18039,N_14219,N_12327);
xor U18040 (N_18040,N_12302,N_11660);
and U18041 (N_18041,N_13084,N_11393);
nor U18042 (N_18042,N_13779,N_14406);
or U18043 (N_18043,N_12162,N_14042);
and U18044 (N_18044,N_10677,N_11881);
xnor U18045 (N_18045,N_14902,N_11948);
or U18046 (N_18046,N_13178,N_12659);
or U18047 (N_18047,N_11126,N_10099);
nor U18048 (N_18048,N_14945,N_10057);
and U18049 (N_18049,N_11740,N_14859);
xor U18050 (N_18050,N_12643,N_12055);
nand U18051 (N_18051,N_11014,N_12868);
nor U18052 (N_18052,N_12559,N_10563);
nor U18053 (N_18053,N_11068,N_13831);
and U18054 (N_18054,N_11587,N_10211);
and U18055 (N_18055,N_13434,N_14860);
or U18056 (N_18056,N_11915,N_12519);
and U18057 (N_18057,N_14194,N_10707);
nor U18058 (N_18058,N_12636,N_11738);
nand U18059 (N_18059,N_13881,N_14984);
or U18060 (N_18060,N_11606,N_12870);
or U18061 (N_18061,N_14392,N_14276);
and U18062 (N_18062,N_10094,N_10325);
xnor U18063 (N_18063,N_11241,N_11055);
xnor U18064 (N_18064,N_14440,N_10291);
nor U18065 (N_18065,N_14096,N_12034);
or U18066 (N_18066,N_11901,N_14346);
or U18067 (N_18067,N_13549,N_12076);
nand U18068 (N_18068,N_12326,N_13393);
nor U18069 (N_18069,N_12987,N_13852);
xnor U18070 (N_18070,N_10542,N_13792);
xor U18071 (N_18071,N_14407,N_14197);
xnor U18072 (N_18072,N_12864,N_12213);
xor U18073 (N_18073,N_13666,N_14116);
xnor U18074 (N_18074,N_12490,N_13456);
and U18075 (N_18075,N_11725,N_10605);
or U18076 (N_18076,N_13456,N_14076);
and U18077 (N_18077,N_11525,N_10970);
or U18078 (N_18078,N_13573,N_13989);
nand U18079 (N_18079,N_12708,N_11004);
or U18080 (N_18080,N_14435,N_10192);
nor U18081 (N_18081,N_11658,N_12702);
and U18082 (N_18082,N_11597,N_14694);
nand U18083 (N_18083,N_13728,N_10749);
nor U18084 (N_18084,N_10597,N_10432);
and U18085 (N_18085,N_10850,N_11680);
nor U18086 (N_18086,N_11465,N_11756);
or U18087 (N_18087,N_11040,N_14727);
or U18088 (N_18088,N_11869,N_12276);
xnor U18089 (N_18089,N_14567,N_14243);
nor U18090 (N_18090,N_10669,N_10236);
nor U18091 (N_18091,N_10995,N_12003);
nor U18092 (N_18092,N_13426,N_12842);
or U18093 (N_18093,N_12359,N_12690);
or U18094 (N_18094,N_10751,N_13611);
nor U18095 (N_18095,N_11186,N_12531);
nand U18096 (N_18096,N_10730,N_12459);
xnor U18097 (N_18097,N_12267,N_13101);
nand U18098 (N_18098,N_11821,N_10086);
xor U18099 (N_18099,N_13717,N_11419);
or U18100 (N_18100,N_10115,N_11977);
nor U18101 (N_18101,N_14682,N_13504);
or U18102 (N_18102,N_12385,N_14800);
or U18103 (N_18103,N_13163,N_12134);
nand U18104 (N_18104,N_13836,N_14711);
xnor U18105 (N_18105,N_13595,N_14009);
xnor U18106 (N_18106,N_13229,N_12227);
xnor U18107 (N_18107,N_13441,N_11158);
nand U18108 (N_18108,N_14368,N_11494);
or U18109 (N_18109,N_11760,N_14567);
or U18110 (N_18110,N_13018,N_12900);
and U18111 (N_18111,N_12836,N_12234);
nor U18112 (N_18112,N_10656,N_13447);
or U18113 (N_18113,N_11779,N_10921);
nor U18114 (N_18114,N_11570,N_12978);
nand U18115 (N_18115,N_11411,N_12335);
xor U18116 (N_18116,N_12048,N_14051);
nor U18117 (N_18117,N_11580,N_13171);
and U18118 (N_18118,N_11133,N_13258);
or U18119 (N_18119,N_12365,N_10455);
nand U18120 (N_18120,N_13524,N_11047);
and U18121 (N_18121,N_13228,N_10010);
or U18122 (N_18122,N_10475,N_13871);
nor U18123 (N_18123,N_13725,N_10220);
or U18124 (N_18124,N_10377,N_12388);
xnor U18125 (N_18125,N_10426,N_10819);
and U18126 (N_18126,N_11877,N_10548);
nand U18127 (N_18127,N_12143,N_11241);
xor U18128 (N_18128,N_10602,N_10311);
or U18129 (N_18129,N_11086,N_10025);
nor U18130 (N_18130,N_12792,N_12012);
and U18131 (N_18131,N_12780,N_11111);
nand U18132 (N_18132,N_11752,N_12528);
nand U18133 (N_18133,N_14684,N_12713);
and U18134 (N_18134,N_11510,N_11377);
nor U18135 (N_18135,N_12026,N_14421);
xnor U18136 (N_18136,N_13236,N_13245);
and U18137 (N_18137,N_12034,N_11400);
xor U18138 (N_18138,N_10291,N_11675);
nor U18139 (N_18139,N_11169,N_14226);
nor U18140 (N_18140,N_14203,N_10475);
nor U18141 (N_18141,N_14808,N_12255);
xnor U18142 (N_18142,N_14106,N_12237);
or U18143 (N_18143,N_10423,N_14149);
nor U18144 (N_18144,N_13414,N_11487);
xnor U18145 (N_18145,N_10719,N_11017);
nor U18146 (N_18146,N_14113,N_13996);
nor U18147 (N_18147,N_10047,N_12183);
or U18148 (N_18148,N_10783,N_12053);
nor U18149 (N_18149,N_11179,N_10426);
nor U18150 (N_18150,N_12023,N_14345);
or U18151 (N_18151,N_14864,N_12370);
nand U18152 (N_18152,N_13685,N_14623);
nor U18153 (N_18153,N_12809,N_10471);
xor U18154 (N_18154,N_14434,N_14825);
or U18155 (N_18155,N_14721,N_11006);
and U18156 (N_18156,N_11933,N_14284);
or U18157 (N_18157,N_14959,N_12344);
xnor U18158 (N_18158,N_13022,N_12718);
or U18159 (N_18159,N_10439,N_13853);
nor U18160 (N_18160,N_14862,N_13153);
and U18161 (N_18161,N_10413,N_11798);
xor U18162 (N_18162,N_13852,N_10704);
or U18163 (N_18163,N_11954,N_11347);
or U18164 (N_18164,N_13512,N_13414);
xnor U18165 (N_18165,N_14003,N_10045);
and U18166 (N_18166,N_11751,N_10195);
nand U18167 (N_18167,N_11066,N_14337);
nand U18168 (N_18168,N_10191,N_12322);
nor U18169 (N_18169,N_10984,N_12382);
or U18170 (N_18170,N_10995,N_10841);
xnor U18171 (N_18171,N_10508,N_12206);
and U18172 (N_18172,N_11981,N_13671);
and U18173 (N_18173,N_11519,N_14786);
and U18174 (N_18174,N_12876,N_11169);
and U18175 (N_18175,N_13692,N_13089);
or U18176 (N_18176,N_12614,N_13221);
or U18177 (N_18177,N_10470,N_13787);
and U18178 (N_18178,N_14165,N_13688);
or U18179 (N_18179,N_11534,N_11317);
nor U18180 (N_18180,N_14036,N_14094);
and U18181 (N_18181,N_10592,N_14869);
or U18182 (N_18182,N_10820,N_12341);
nand U18183 (N_18183,N_11755,N_13509);
or U18184 (N_18184,N_13868,N_11941);
and U18185 (N_18185,N_14632,N_13242);
or U18186 (N_18186,N_12914,N_10501);
xor U18187 (N_18187,N_14459,N_14393);
xnor U18188 (N_18188,N_14238,N_14695);
and U18189 (N_18189,N_11543,N_14944);
or U18190 (N_18190,N_14635,N_10717);
or U18191 (N_18191,N_12635,N_13160);
and U18192 (N_18192,N_14013,N_12175);
or U18193 (N_18193,N_12001,N_10278);
nand U18194 (N_18194,N_13663,N_10779);
or U18195 (N_18195,N_13591,N_13014);
nor U18196 (N_18196,N_12237,N_14738);
nor U18197 (N_18197,N_12505,N_13918);
xnor U18198 (N_18198,N_13902,N_13704);
nor U18199 (N_18199,N_14513,N_14481);
nand U18200 (N_18200,N_11002,N_11099);
and U18201 (N_18201,N_14092,N_11614);
nand U18202 (N_18202,N_11879,N_14932);
nor U18203 (N_18203,N_14589,N_12234);
or U18204 (N_18204,N_14785,N_13118);
or U18205 (N_18205,N_12300,N_11073);
nand U18206 (N_18206,N_12597,N_13514);
nand U18207 (N_18207,N_11160,N_14685);
nand U18208 (N_18208,N_11904,N_14767);
xor U18209 (N_18209,N_11269,N_11626);
and U18210 (N_18210,N_11191,N_13333);
and U18211 (N_18211,N_10012,N_14588);
or U18212 (N_18212,N_14020,N_12606);
nand U18213 (N_18213,N_10842,N_12071);
and U18214 (N_18214,N_11005,N_14549);
or U18215 (N_18215,N_11335,N_13285);
and U18216 (N_18216,N_14757,N_14436);
xor U18217 (N_18217,N_14247,N_11064);
xor U18218 (N_18218,N_13201,N_14278);
nand U18219 (N_18219,N_13948,N_11903);
nand U18220 (N_18220,N_14463,N_11484);
or U18221 (N_18221,N_11916,N_14457);
xor U18222 (N_18222,N_12535,N_11485);
or U18223 (N_18223,N_12462,N_10612);
and U18224 (N_18224,N_11948,N_14613);
nor U18225 (N_18225,N_13944,N_13955);
xor U18226 (N_18226,N_12746,N_12174);
nand U18227 (N_18227,N_12484,N_13943);
nand U18228 (N_18228,N_10469,N_14788);
nor U18229 (N_18229,N_13743,N_11757);
and U18230 (N_18230,N_10827,N_14995);
and U18231 (N_18231,N_13539,N_13238);
nand U18232 (N_18232,N_14597,N_11432);
nor U18233 (N_18233,N_14115,N_11570);
and U18234 (N_18234,N_13102,N_12424);
xnor U18235 (N_18235,N_12854,N_11697);
nor U18236 (N_18236,N_12029,N_13874);
nand U18237 (N_18237,N_13324,N_11625);
nor U18238 (N_18238,N_10665,N_14430);
nor U18239 (N_18239,N_14086,N_13407);
and U18240 (N_18240,N_13996,N_11357);
xor U18241 (N_18241,N_14881,N_13043);
or U18242 (N_18242,N_14033,N_14305);
nor U18243 (N_18243,N_10610,N_14473);
nor U18244 (N_18244,N_14744,N_13733);
nor U18245 (N_18245,N_11423,N_10460);
xor U18246 (N_18246,N_11671,N_13129);
and U18247 (N_18247,N_11843,N_12737);
or U18248 (N_18248,N_13896,N_12036);
nor U18249 (N_18249,N_13479,N_13588);
or U18250 (N_18250,N_10411,N_10960);
nand U18251 (N_18251,N_11588,N_12572);
or U18252 (N_18252,N_11921,N_11431);
or U18253 (N_18253,N_13876,N_12685);
and U18254 (N_18254,N_11522,N_13329);
or U18255 (N_18255,N_10753,N_12725);
nand U18256 (N_18256,N_12173,N_12325);
and U18257 (N_18257,N_14936,N_11203);
or U18258 (N_18258,N_14786,N_13827);
nor U18259 (N_18259,N_10781,N_13445);
nor U18260 (N_18260,N_10368,N_14091);
xor U18261 (N_18261,N_10269,N_14261);
or U18262 (N_18262,N_11062,N_14242);
nand U18263 (N_18263,N_12016,N_14594);
and U18264 (N_18264,N_11078,N_13326);
nor U18265 (N_18265,N_13087,N_11816);
nor U18266 (N_18266,N_14786,N_11375);
nand U18267 (N_18267,N_13248,N_11166);
and U18268 (N_18268,N_13398,N_11621);
nand U18269 (N_18269,N_10320,N_10838);
nand U18270 (N_18270,N_13345,N_10002);
nand U18271 (N_18271,N_13736,N_11115);
or U18272 (N_18272,N_10848,N_11278);
nor U18273 (N_18273,N_14374,N_12424);
xnor U18274 (N_18274,N_14877,N_10813);
xor U18275 (N_18275,N_13295,N_14238);
nor U18276 (N_18276,N_12415,N_10910);
xnor U18277 (N_18277,N_12784,N_14542);
nand U18278 (N_18278,N_14344,N_14759);
and U18279 (N_18279,N_13702,N_14282);
or U18280 (N_18280,N_11286,N_10501);
xor U18281 (N_18281,N_11220,N_14284);
and U18282 (N_18282,N_13873,N_12233);
nand U18283 (N_18283,N_14901,N_10704);
nand U18284 (N_18284,N_11899,N_13169);
nor U18285 (N_18285,N_13145,N_12742);
and U18286 (N_18286,N_12598,N_14199);
xnor U18287 (N_18287,N_10918,N_11151);
or U18288 (N_18288,N_14181,N_11835);
nand U18289 (N_18289,N_10425,N_11817);
and U18290 (N_18290,N_13597,N_11552);
and U18291 (N_18291,N_13695,N_13354);
xnor U18292 (N_18292,N_11231,N_11727);
and U18293 (N_18293,N_12077,N_14560);
nand U18294 (N_18294,N_13292,N_14215);
nand U18295 (N_18295,N_11314,N_10932);
xnor U18296 (N_18296,N_12497,N_10723);
nor U18297 (N_18297,N_11767,N_11484);
nor U18298 (N_18298,N_13182,N_13280);
and U18299 (N_18299,N_10204,N_14268);
nor U18300 (N_18300,N_13074,N_10305);
nor U18301 (N_18301,N_11577,N_12189);
nor U18302 (N_18302,N_10456,N_13170);
or U18303 (N_18303,N_12697,N_11750);
nor U18304 (N_18304,N_12796,N_14956);
and U18305 (N_18305,N_13156,N_10237);
nor U18306 (N_18306,N_12373,N_12726);
and U18307 (N_18307,N_14005,N_10504);
nor U18308 (N_18308,N_11069,N_11279);
xor U18309 (N_18309,N_12641,N_12040);
and U18310 (N_18310,N_11882,N_13630);
and U18311 (N_18311,N_13152,N_11443);
or U18312 (N_18312,N_12774,N_10607);
nor U18313 (N_18313,N_11539,N_11845);
or U18314 (N_18314,N_11806,N_14374);
and U18315 (N_18315,N_13910,N_10181);
nand U18316 (N_18316,N_12856,N_13735);
xnor U18317 (N_18317,N_13809,N_12373);
xnor U18318 (N_18318,N_11885,N_11530);
and U18319 (N_18319,N_13680,N_10995);
nor U18320 (N_18320,N_14517,N_14520);
nor U18321 (N_18321,N_14186,N_12275);
or U18322 (N_18322,N_12362,N_13806);
or U18323 (N_18323,N_12471,N_14335);
or U18324 (N_18324,N_14214,N_14705);
nor U18325 (N_18325,N_12498,N_11315);
nand U18326 (N_18326,N_13966,N_12667);
and U18327 (N_18327,N_10559,N_10169);
and U18328 (N_18328,N_13032,N_12257);
or U18329 (N_18329,N_14293,N_13410);
and U18330 (N_18330,N_11531,N_14080);
and U18331 (N_18331,N_10108,N_14938);
xor U18332 (N_18332,N_14337,N_10379);
or U18333 (N_18333,N_13818,N_11643);
and U18334 (N_18334,N_10145,N_10950);
nor U18335 (N_18335,N_11734,N_10824);
nand U18336 (N_18336,N_13927,N_14207);
or U18337 (N_18337,N_10201,N_13568);
xnor U18338 (N_18338,N_12164,N_14529);
nand U18339 (N_18339,N_10645,N_11225);
nand U18340 (N_18340,N_11950,N_14497);
nor U18341 (N_18341,N_10451,N_10268);
and U18342 (N_18342,N_13373,N_10572);
nor U18343 (N_18343,N_10688,N_13438);
nor U18344 (N_18344,N_14397,N_12147);
or U18345 (N_18345,N_10842,N_10831);
or U18346 (N_18346,N_11101,N_10342);
and U18347 (N_18347,N_12872,N_11017);
nand U18348 (N_18348,N_13715,N_12976);
nand U18349 (N_18349,N_10722,N_10354);
or U18350 (N_18350,N_12609,N_10870);
nor U18351 (N_18351,N_13075,N_10272);
or U18352 (N_18352,N_12961,N_12946);
nor U18353 (N_18353,N_13007,N_11704);
xnor U18354 (N_18354,N_13449,N_13436);
nand U18355 (N_18355,N_10353,N_14956);
nand U18356 (N_18356,N_10412,N_14640);
xnor U18357 (N_18357,N_13879,N_10328);
xnor U18358 (N_18358,N_14486,N_11058);
or U18359 (N_18359,N_13743,N_13445);
nor U18360 (N_18360,N_14045,N_12941);
nor U18361 (N_18361,N_13927,N_13872);
nor U18362 (N_18362,N_13417,N_11889);
or U18363 (N_18363,N_10968,N_10453);
and U18364 (N_18364,N_13757,N_14378);
nand U18365 (N_18365,N_14351,N_10158);
and U18366 (N_18366,N_10298,N_13333);
nand U18367 (N_18367,N_13714,N_13081);
nand U18368 (N_18368,N_11219,N_12975);
nand U18369 (N_18369,N_14485,N_14629);
and U18370 (N_18370,N_12257,N_11527);
nand U18371 (N_18371,N_12617,N_10641);
and U18372 (N_18372,N_12149,N_11926);
or U18373 (N_18373,N_11865,N_12619);
or U18374 (N_18374,N_14279,N_11527);
nor U18375 (N_18375,N_11488,N_13549);
nand U18376 (N_18376,N_14352,N_13931);
nor U18377 (N_18377,N_12208,N_14083);
and U18378 (N_18378,N_13785,N_14558);
nand U18379 (N_18379,N_11277,N_10708);
nand U18380 (N_18380,N_11768,N_13173);
or U18381 (N_18381,N_13230,N_11926);
nor U18382 (N_18382,N_10198,N_11180);
nand U18383 (N_18383,N_13771,N_12378);
nand U18384 (N_18384,N_12542,N_13518);
or U18385 (N_18385,N_12802,N_11547);
nand U18386 (N_18386,N_10398,N_11126);
or U18387 (N_18387,N_10246,N_11569);
nand U18388 (N_18388,N_13731,N_12157);
or U18389 (N_18389,N_14371,N_10236);
nand U18390 (N_18390,N_10043,N_14825);
and U18391 (N_18391,N_13199,N_12686);
or U18392 (N_18392,N_14242,N_13481);
or U18393 (N_18393,N_13486,N_14988);
nand U18394 (N_18394,N_12280,N_10505);
xor U18395 (N_18395,N_14928,N_13336);
xor U18396 (N_18396,N_14843,N_14769);
or U18397 (N_18397,N_12849,N_14580);
and U18398 (N_18398,N_13012,N_13180);
and U18399 (N_18399,N_10829,N_12946);
xnor U18400 (N_18400,N_14703,N_14574);
xnor U18401 (N_18401,N_11857,N_10149);
and U18402 (N_18402,N_11031,N_14733);
and U18403 (N_18403,N_10440,N_12055);
and U18404 (N_18404,N_11433,N_12330);
and U18405 (N_18405,N_11829,N_11657);
or U18406 (N_18406,N_14715,N_13719);
or U18407 (N_18407,N_12360,N_12773);
or U18408 (N_18408,N_12806,N_12401);
nor U18409 (N_18409,N_11460,N_12659);
or U18410 (N_18410,N_10523,N_12089);
or U18411 (N_18411,N_14008,N_13303);
or U18412 (N_18412,N_11739,N_13238);
nand U18413 (N_18413,N_14587,N_10831);
xor U18414 (N_18414,N_13403,N_12892);
or U18415 (N_18415,N_10650,N_11353);
and U18416 (N_18416,N_13021,N_12109);
and U18417 (N_18417,N_13656,N_14144);
nor U18418 (N_18418,N_14259,N_14143);
or U18419 (N_18419,N_10306,N_11334);
and U18420 (N_18420,N_13555,N_12231);
or U18421 (N_18421,N_12219,N_10020);
nand U18422 (N_18422,N_13237,N_12913);
nor U18423 (N_18423,N_13006,N_14588);
nand U18424 (N_18424,N_13415,N_13584);
nand U18425 (N_18425,N_14976,N_10244);
nand U18426 (N_18426,N_13642,N_10556);
nand U18427 (N_18427,N_13863,N_14785);
nor U18428 (N_18428,N_11321,N_12748);
nand U18429 (N_18429,N_13660,N_11126);
nand U18430 (N_18430,N_11066,N_13862);
nor U18431 (N_18431,N_11735,N_10468);
nand U18432 (N_18432,N_12904,N_10271);
nand U18433 (N_18433,N_14312,N_12341);
xor U18434 (N_18434,N_14724,N_14444);
nor U18435 (N_18435,N_10199,N_13727);
or U18436 (N_18436,N_14282,N_12912);
nand U18437 (N_18437,N_13597,N_13473);
nand U18438 (N_18438,N_12293,N_10084);
or U18439 (N_18439,N_11051,N_14633);
xnor U18440 (N_18440,N_14194,N_12900);
xnor U18441 (N_18441,N_11345,N_14455);
and U18442 (N_18442,N_13436,N_11323);
or U18443 (N_18443,N_10601,N_11421);
and U18444 (N_18444,N_12149,N_10303);
and U18445 (N_18445,N_10173,N_10783);
xor U18446 (N_18446,N_12530,N_11447);
or U18447 (N_18447,N_12635,N_14150);
nor U18448 (N_18448,N_12604,N_12614);
nand U18449 (N_18449,N_13255,N_14579);
xor U18450 (N_18450,N_13850,N_11709);
and U18451 (N_18451,N_14688,N_14951);
and U18452 (N_18452,N_12188,N_11951);
or U18453 (N_18453,N_12317,N_10077);
nor U18454 (N_18454,N_11046,N_11821);
nor U18455 (N_18455,N_13250,N_11128);
xor U18456 (N_18456,N_13491,N_12784);
nand U18457 (N_18457,N_11332,N_13912);
or U18458 (N_18458,N_12177,N_14105);
and U18459 (N_18459,N_14137,N_11112);
nand U18460 (N_18460,N_14034,N_13556);
and U18461 (N_18461,N_11923,N_10733);
and U18462 (N_18462,N_14636,N_11302);
or U18463 (N_18463,N_10857,N_11774);
nor U18464 (N_18464,N_11145,N_13658);
xor U18465 (N_18465,N_13900,N_10117);
xor U18466 (N_18466,N_10340,N_10173);
or U18467 (N_18467,N_13592,N_11704);
xnor U18468 (N_18468,N_13636,N_12424);
nor U18469 (N_18469,N_13933,N_13161);
nor U18470 (N_18470,N_11047,N_14766);
nand U18471 (N_18471,N_14156,N_14657);
nand U18472 (N_18472,N_10197,N_13667);
and U18473 (N_18473,N_12302,N_10378);
nand U18474 (N_18474,N_11699,N_13340);
and U18475 (N_18475,N_12133,N_10887);
and U18476 (N_18476,N_13710,N_11641);
nand U18477 (N_18477,N_10368,N_11594);
xnor U18478 (N_18478,N_11203,N_13179);
and U18479 (N_18479,N_12191,N_11111);
nor U18480 (N_18480,N_10249,N_10418);
nor U18481 (N_18481,N_11325,N_10658);
nor U18482 (N_18482,N_12427,N_11547);
nand U18483 (N_18483,N_13479,N_14628);
nor U18484 (N_18484,N_13613,N_13920);
nor U18485 (N_18485,N_11072,N_13076);
nand U18486 (N_18486,N_13924,N_12232);
nor U18487 (N_18487,N_13473,N_11785);
xor U18488 (N_18488,N_13369,N_12265);
nand U18489 (N_18489,N_14445,N_12665);
and U18490 (N_18490,N_11682,N_12509);
and U18491 (N_18491,N_10490,N_11216);
nor U18492 (N_18492,N_12306,N_11700);
xnor U18493 (N_18493,N_12988,N_14298);
nand U18494 (N_18494,N_10887,N_12393);
nor U18495 (N_18495,N_12205,N_10346);
xnor U18496 (N_18496,N_14827,N_12215);
nor U18497 (N_18497,N_12091,N_10505);
nand U18498 (N_18498,N_11452,N_13392);
or U18499 (N_18499,N_10474,N_13949);
nor U18500 (N_18500,N_14024,N_12492);
or U18501 (N_18501,N_11924,N_13785);
nor U18502 (N_18502,N_12814,N_14364);
or U18503 (N_18503,N_12290,N_11612);
nand U18504 (N_18504,N_14516,N_14601);
and U18505 (N_18505,N_11584,N_14806);
nor U18506 (N_18506,N_14625,N_13524);
nor U18507 (N_18507,N_13122,N_12761);
nand U18508 (N_18508,N_11949,N_12818);
nor U18509 (N_18509,N_12809,N_14048);
and U18510 (N_18510,N_11862,N_12895);
or U18511 (N_18511,N_11949,N_11390);
nor U18512 (N_18512,N_12297,N_10332);
or U18513 (N_18513,N_12923,N_10959);
and U18514 (N_18514,N_10513,N_13391);
xnor U18515 (N_18515,N_12996,N_14428);
and U18516 (N_18516,N_13377,N_11152);
nand U18517 (N_18517,N_14723,N_10490);
nor U18518 (N_18518,N_12460,N_14172);
nand U18519 (N_18519,N_10179,N_12519);
nand U18520 (N_18520,N_10386,N_10804);
and U18521 (N_18521,N_10314,N_10675);
and U18522 (N_18522,N_13990,N_10953);
and U18523 (N_18523,N_14003,N_11558);
nor U18524 (N_18524,N_10391,N_14678);
or U18525 (N_18525,N_12061,N_11330);
xnor U18526 (N_18526,N_14169,N_13897);
nor U18527 (N_18527,N_10906,N_14677);
and U18528 (N_18528,N_14999,N_14426);
and U18529 (N_18529,N_14915,N_13655);
or U18530 (N_18530,N_12791,N_10495);
nor U18531 (N_18531,N_12260,N_12121);
nor U18532 (N_18532,N_10482,N_12046);
xnor U18533 (N_18533,N_14129,N_11740);
nand U18534 (N_18534,N_14647,N_11837);
and U18535 (N_18535,N_14533,N_12236);
nor U18536 (N_18536,N_11511,N_12710);
nor U18537 (N_18537,N_12632,N_12253);
and U18538 (N_18538,N_10468,N_13310);
or U18539 (N_18539,N_12730,N_13996);
or U18540 (N_18540,N_13047,N_10357);
nor U18541 (N_18541,N_13574,N_11405);
nor U18542 (N_18542,N_12304,N_14520);
nor U18543 (N_18543,N_14450,N_13038);
xnor U18544 (N_18544,N_13528,N_13886);
xnor U18545 (N_18545,N_11279,N_12796);
and U18546 (N_18546,N_11653,N_11199);
nor U18547 (N_18547,N_14494,N_14186);
xor U18548 (N_18548,N_11075,N_11965);
and U18549 (N_18549,N_11854,N_14022);
and U18550 (N_18550,N_13050,N_14174);
nand U18551 (N_18551,N_12701,N_10184);
nor U18552 (N_18552,N_11345,N_14373);
nand U18553 (N_18553,N_14367,N_14882);
nand U18554 (N_18554,N_12035,N_12275);
nor U18555 (N_18555,N_13905,N_14498);
nor U18556 (N_18556,N_13788,N_11121);
nor U18557 (N_18557,N_14588,N_10583);
xor U18558 (N_18558,N_14337,N_14649);
nor U18559 (N_18559,N_11336,N_13736);
and U18560 (N_18560,N_12538,N_10100);
nand U18561 (N_18561,N_14186,N_12666);
and U18562 (N_18562,N_11183,N_14466);
nand U18563 (N_18563,N_13557,N_12308);
and U18564 (N_18564,N_12561,N_10828);
and U18565 (N_18565,N_14024,N_14451);
xnor U18566 (N_18566,N_12697,N_10680);
and U18567 (N_18567,N_14919,N_12930);
or U18568 (N_18568,N_13649,N_10377);
and U18569 (N_18569,N_10625,N_12260);
or U18570 (N_18570,N_12908,N_11374);
nand U18571 (N_18571,N_14913,N_12193);
nand U18572 (N_18572,N_11006,N_14531);
nor U18573 (N_18573,N_11291,N_11964);
nand U18574 (N_18574,N_10370,N_14362);
and U18575 (N_18575,N_13537,N_14493);
and U18576 (N_18576,N_14685,N_10033);
and U18577 (N_18577,N_12123,N_13099);
nor U18578 (N_18578,N_14783,N_13834);
xnor U18579 (N_18579,N_12269,N_10213);
nor U18580 (N_18580,N_10753,N_10273);
nand U18581 (N_18581,N_11945,N_11724);
nand U18582 (N_18582,N_11720,N_13740);
or U18583 (N_18583,N_13799,N_10793);
xor U18584 (N_18584,N_13765,N_10964);
nor U18585 (N_18585,N_12986,N_14202);
nand U18586 (N_18586,N_11907,N_13452);
xnor U18587 (N_18587,N_11954,N_11524);
and U18588 (N_18588,N_14032,N_13084);
nand U18589 (N_18589,N_12065,N_10194);
or U18590 (N_18590,N_11944,N_13259);
nor U18591 (N_18591,N_11815,N_13782);
or U18592 (N_18592,N_14477,N_12952);
xor U18593 (N_18593,N_12877,N_13444);
xnor U18594 (N_18594,N_10427,N_12945);
nand U18595 (N_18595,N_10999,N_10492);
xnor U18596 (N_18596,N_10804,N_14937);
xor U18597 (N_18597,N_11070,N_13566);
and U18598 (N_18598,N_11565,N_10358);
xor U18599 (N_18599,N_13080,N_13783);
and U18600 (N_18600,N_12183,N_12445);
or U18601 (N_18601,N_13096,N_11364);
or U18602 (N_18602,N_12260,N_10119);
and U18603 (N_18603,N_12929,N_11154);
and U18604 (N_18604,N_14060,N_14966);
nor U18605 (N_18605,N_10141,N_14984);
and U18606 (N_18606,N_14214,N_14669);
and U18607 (N_18607,N_14031,N_14883);
xnor U18608 (N_18608,N_12001,N_13245);
or U18609 (N_18609,N_13946,N_11487);
xnor U18610 (N_18610,N_13701,N_12520);
nand U18611 (N_18611,N_12845,N_13715);
or U18612 (N_18612,N_10421,N_10772);
or U18613 (N_18613,N_10727,N_11175);
or U18614 (N_18614,N_11463,N_11966);
nor U18615 (N_18615,N_13749,N_10195);
or U18616 (N_18616,N_14785,N_14042);
and U18617 (N_18617,N_12194,N_13113);
nand U18618 (N_18618,N_11420,N_14806);
nor U18619 (N_18619,N_11192,N_12236);
or U18620 (N_18620,N_10392,N_14656);
xnor U18621 (N_18621,N_12062,N_14820);
and U18622 (N_18622,N_14819,N_10861);
nand U18623 (N_18623,N_14470,N_13331);
nor U18624 (N_18624,N_11906,N_12757);
nand U18625 (N_18625,N_10288,N_13497);
xnor U18626 (N_18626,N_14875,N_12639);
nand U18627 (N_18627,N_13457,N_14043);
or U18628 (N_18628,N_11345,N_10733);
or U18629 (N_18629,N_11885,N_10417);
nor U18630 (N_18630,N_10727,N_12682);
nor U18631 (N_18631,N_14151,N_12675);
nor U18632 (N_18632,N_10700,N_12760);
and U18633 (N_18633,N_14337,N_10173);
and U18634 (N_18634,N_12394,N_13732);
and U18635 (N_18635,N_11438,N_10473);
or U18636 (N_18636,N_12837,N_13699);
nor U18637 (N_18637,N_10978,N_14952);
and U18638 (N_18638,N_10103,N_10645);
or U18639 (N_18639,N_10178,N_13415);
nor U18640 (N_18640,N_11310,N_14568);
nor U18641 (N_18641,N_11059,N_10875);
nor U18642 (N_18642,N_11568,N_11991);
nand U18643 (N_18643,N_10234,N_14438);
nor U18644 (N_18644,N_14839,N_12808);
or U18645 (N_18645,N_13578,N_12880);
xor U18646 (N_18646,N_13484,N_13908);
and U18647 (N_18647,N_13810,N_12275);
xor U18648 (N_18648,N_12004,N_13302);
xor U18649 (N_18649,N_14348,N_14128);
nand U18650 (N_18650,N_14810,N_10383);
xor U18651 (N_18651,N_12861,N_10334);
nand U18652 (N_18652,N_13630,N_11870);
nand U18653 (N_18653,N_10575,N_11967);
nor U18654 (N_18654,N_11055,N_11413);
or U18655 (N_18655,N_14339,N_10767);
xnor U18656 (N_18656,N_11086,N_11225);
and U18657 (N_18657,N_12352,N_13485);
or U18658 (N_18658,N_11763,N_14678);
xor U18659 (N_18659,N_13779,N_12513);
and U18660 (N_18660,N_12607,N_14588);
xor U18661 (N_18661,N_14253,N_14584);
and U18662 (N_18662,N_13920,N_11004);
xnor U18663 (N_18663,N_12913,N_11191);
or U18664 (N_18664,N_14326,N_11215);
nor U18665 (N_18665,N_14006,N_12041);
nand U18666 (N_18666,N_10829,N_11766);
or U18667 (N_18667,N_14663,N_12859);
and U18668 (N_18668,N_10619,N_10827);
or U18669 (N_18669,N_11063,N_12222);
nor U18670 (N_18670,N_12094,N_13484);
nand U18671 (N_18671,N_12371,N_10754);
or U18672 (N_18672,N_11016,N_13184);
nand U18673 (N_18673,N_14082,N_10423);
nor U18674 (N_18674,N_10709,N_13031);
and U18675 (N_18675,N_12342,N_11995);
and U18676 (N_18676,N_13308,N_11352);
nand U18677 (N_18677,N_14605,N_13579);
or U18678 (N_18678,N_13395,N_13458);
nand U18679 (N_18679,N_11437,N_10261);
and U18680 (N_18680,N_13033,N_10123);
nand U18681 (N_18681,N_12085,N_14215);
and U18682 (N_18682,N_10281,N_14734);
xor U18683 (N_18683,N_12106,N_13200);
or U18684 (N_18684,N_14752,N_14939);
and U18685 (N_18685,N_14830,N_11052);
or U18686 (N_18686,N_10007,N_12669);
and U18687 (N_18687,N_13404,N_14478);
or U18688 (N_18688,N_10250,N_13325);
nand U18689 (N_18689,N_13971,N_10385);
nand U18690 (N_18690,N_11678,N_12874);
and U18691 (N_18691,N_12437,N_13275);
xor U18692 (N_18692,N_12852,N_11621);
nor U18693 (N_18693,N_11105,N_13282);
xor U18694 (N_18694,N_14876,N_12754);
or U18695 (N_18695,N_13724,N_14332);
xnor U18696 (N_18696,N_12305,N_14032);
or U18697 (N_18697,N_12821,N_11803);
xor U18698 (N_18698,N_10163,N_11125);
nor U18699 (N_18699,N_11520,N_14140);
nand U18700 (N_18700,N_11750,N_13413);
xnor U18701 (N_18701,N_12540,N_13505);
xor U18702 (N_18702,N_11114,N_12728);
or U18703 (N_18703,N_13419,N_11716);
and U18704 (N_18704,N_12582,N_10360);
nor U18705 (N_18705,N_10931,N_10089);
xor U18706 (N_18706,N_13637,N_10497);
xor U18707 (N_18707,N_12716,N_11999);
xor U18708 (N_18708,N_13927,N_14708);
nand U18709 (N_18709,N_11558,N_11721);
and U18710 (N_18710,N_13114,N_11063);
xor U18711 (N_18711,N_10386,N_13372);
nor U18712 (N_18712,N_10020,N_11493);
xor U18713 (N_18713,N_13890,N_10098);
nand U18714 (N_18714,N_13836,N_13333);
xor U18715 (N_18715,N_13397,N_14422);
and U18716 (N_18716,N_11418,N_12369);
nor U18717 (N_18717,N_10171,N_12057);
and U18718 (N_18718,N_12128,N_14998);
nand U18719 (N_18719,N_11249,N_13247);
nand U18720 (N_18720,N_13116,N_11448);
or U18721 (N_18721,N_11935,N_11475);
nor U18722 (N_18722,N_10738,N_12121);
or U18723 (N_18723,N_12303,N_10138);
or U18724 (N_18724,N_14766,N_12515);
nand U18725 (N_18725,N_10368,N_10858);
xnor U18726 (N_18726,N_11012,N_12640);
nand U18727 (N_18727,N_11930,N_12994);
and U18728 (N_18728,N_14031,N_13421);
nand U18729 (N_18729,N_11755,N_10523);
and U18730 (N_18730,N_12309,N_13081);
nor U18731 (N_18731,N_13405,N_13670);
nor U18732 (N_18732,N_11948,N_10435);
xnor U18733 (N_18733,N_14506,N_12387);
and U18734 (N_18734,N_10040,N_11105);
nor U18735 (N_18735,N_14477,N_10127);
or U18736 (N_18736,N_10187,N_12809);
nand U18737 (N_18737,N_11621,N_11052);
and U18738 (N_18738,N_13551,N_14129);
or U18739 (N_18739,N_10781,N_10630);
nand U18740 (N_18740,N_10632,N_14251);
nor U18741 (N_18741,N_10686,N_14638);
xor U18742 (N_18742,N_10537,N_14310);
nor U18743 (N_18743,N_10062,N_14934);
or U18744 (N_18744,N_11994,N_13899);
xnor U18745 (N_18745,N_10516,N_10015);
nor U18746 (N_18746,N_12117,N_11893);
and U18747 (N_18747,N_12571,N_11963);
or U18748 (N_18748,N_12193,N_13014);
xnor U18749 (N_18749,N_13175,N_13246);
and U18750 (N_18750,N_11406,N_13087);
and U18751 (N_18751,N_11849,N_12415);
nand U18752 (N_18752,N_10184,N_13699);
nor U18753 (N_18753,N_11608,N_11207);
nor U18754 (N_18754,N_10082,N_14554);
nor U18755 (N_18755,N_13924,N_13861);
or U18756 (N_18756,N_10419,N_13482);
nor U18757 (N_18757,N_13688,N_13589);
nor U18758 (N_18758,N_13764,N_10678);
and U18759 (N_18759,N_13373,N_10614);
nor U18760 (N_18760,N_14574,N_10149);
xnor U18761 (N_18761,N_14767,N_13902);
and U18762 (N_18762,N_13179,N_11429);
xor U18763 (N_18763,N_11865,N_12626);
nand U18764 (N_18764,N_12362,N_11889);
xnor U18765 (N_18765,N_13680,N_11254);
nand U18766 (N_18766,N_13052,N_13938);
or U18767 (N_18767,N_11211,N_12378);
nor U18768 (N_18768,N_11873,N_11154);
nor U18769 (N_18769,N_14417,N_12824);
xnor U18770 (N_18770,N_10780,N_10177);
nor U18771 (N_18771,N_11076,N_10919);
and U18772 (N_18772,N_13115,N_11973);
xor U18773 (N_18773,N_12634,N_11747);
xor U18774 (N_18774,N_10161,N_12647);
nor U18775 (N_18775,N_12273,N_11470);
xor U18776 (N_18776,N_11777,N_14224);
and U18777 (N_18777,N_14770,N_14976);
and U18778 (N_18778,N_12669,N_12332);
nor U18779 (N_18779,N_12514,N_14767);
xor U18780 (N_18780,N_10021,N_13280);
nor U18781 (N_18781,N_13893,N_13694);
or U18782 (N_18782,N_12069,N_13180);
or U18783 (N_18783,N_13866,N_12691);
and U18784 (N_18784,N_13958,N_10098);
and U18785 (N_18785,N_13454,N_14767);
nand U18786 (N_18786,N_11096,N_10229);
and U18787 (N_18787,N_11580,N_10748);
or U18788 (N_18788,N_11008,N_13747);
or U18789 (N_18789,N_11948,N_14470);
and U18790 (N_18790,N_12894,N_13964);
nor U18791 (N_18791,N_11751,N_11067);
nor U18792 (N_18792,N_14475,N_10861);
nor U18793 (N_18793,N_12958,N_10769);
xnor U18794 (N_18794,N_14092,N_13813);
and U18795 (N_18795,N_10278,N_13329);
nand U18796 (N_18796,N_10810,N_14990);
or U18797 (N_18797,N_12655,N_14346);
nor U18798 (N_18798,N_14906,N_11436);
nand U18799 (N_18799,N_13407,N_14453);
and U18800 (N_18800,N_10923,N_11825);
and U18801 (N_18801,N_12437,N_11154);
xor U18802 (N_18802,N_12015,N_11265);
and U18803 (N_18803,N_10395,N_10030);
xnor U18804 (N_18804,N_10580,N_10690);
and U18805 (N_18805,N_11916,N_14737);
or U18806 (N_18806,N_12902,N_12451);
xor U18807 (N_18807,N_10606,N_12575);
nor U18808 (N_18808,N_12847,N_13072);
and U18809 (N_18809,N_12200,N_13140);
and U18810 (N_18810,N_11612,N_11456);
xor U18811 (N_18811,N_12844,N_10776);
nand U18812 (N_18812,N_12241,N_14639);
nor U18813 (N_18813,N_11782,N_11423);
and U18814 (N_18814,N_13103,N_13922);
and U18815 (N_18815,N_13569,N_13782);
or U18816 (N_18816,N_13461,N_11230);
and U18817 (N_18817,N_14961,N_11936);
xnor U18818 (N_18818,N_10669,N_11373);
xor U18819 (N_18819,N_12817,N_11897);
or U18820 (N_18820,N_11348,N_13242);
xor U18821 (N_18821,N_10616,N_10085);
nand U18822 (N_18822,N_12815,N_11643);
xnor U18823 (N_18823,N_14526,N_11336);
nand U18824 (N_18824,N_14265,N_12759);
or U18825 (N_18825,N_12232,N_11882);
or U18826 (N_18826,N_10159,N_12788);
and U18827 (N_18827,N_10190,N_12852);
nor U18828 (N_18828,N_11041,N_14783);
nor U18829 (N_18829,N_14098,N_10357);
xnor U18830 (N_18830,N_14110,N_13216);
xor U18831 (N_18831,N_12147,N_14109);
or U18832 (N_18832,N_10195,N_11486);
nand U18833 (N_18833,N_13812,N_12999);
or U18834 (N_18834,N_14550,N_14336);
nand U18835 (N_18835,N_11177,N_12868);
nor U18836 (N_18836,N_14239,N_12458);
nand U18837 (N_18837,N_14174,N_13096);
and U18838 (N_18838,N_12519,N_11165);
nor U18839 (N_18839,N_12107,N_12964);
or U18840 (N_18840,N_11790,N_13944);
or U18841 (N_18841,N_11194,N_12528);
nor U18842 (N_18842,N_11889,N_13009);
nand U18843 (N_18843,N_12576,N_11801);
and U18844 (N_18844,N_12874,N_12774);
and U18845 (N_18845,N_14301,N_11337);
or U18846 (N_18846,N_13387,N_12130);
xnor U18847 (N_18847,N_13284,N_11965);
nand U18848 (N_18848,N_11351,N_10010);
or U18849 (N_18849,N_11453,N_11069);
xnor U18850 (N_18850,N_13699,N_12131);
or U18851 (N_18851,N_13065,N_13272);
nand U18852 (N_18852,N_14130,N_10398);
nor U18853 (N_18853,N_12120,N_12376);
nand U18854 (N_18854,N_13024,N_14715);
and U18855 (N_18855,N_12890,N_14940);
xnor U18856 (N_18856,N_10158,N_13830);
nor U18857 (N_18857,N_13246,N_14247);
and U18858 (N_18858,N_13815,N_14559);
nand U18859 (N_18859,N_11515,N_13526);
xor U18860 (N_18860,N_13663,N_10895);
and U18861 (N_18861,N_11950,N_10858);
and U18862 (N_18862,N_12513,N_14034);
nand U18863 (N_18863,N_12612,N_11201);
nor U18864 (N_18864,N_12413,N_11605);
xor U18865 (N_18865,N_10111,N_12967);
nor U18866 (N_18866,N_12658,N_10268);
or U18867 (N_18867,N_12851,N_12131);
and U18868 (N_18868,N_11689,N_13724);
or U18869 (N_18869,N_12476,N_12776);
nand U18870 (N_18870,N_14676,N_13041);
xor U18871 (N_18871,N_12518,N_12340);
and U18872 (N_18872,N_12279,N_14315);
and U18873 (N_18873,N_12989,N_11539);
xnor U18874 (N_18874,N_13079,N_13287);
xnor U18875 (N_18875,N_10961,N_14875);
and U18876 (N_18876,N_14804,N_13015);
xnor U18877 (N_18877,N_11822,N_13845);
xnor U18878 (N_18878,N_11340,N_11712);
nand U18879 (N_18879,N_11712,N_11378);
nor U18880 (N_18880,N_12671,N_13852);
or U18881 (N_18881,N_12558,N_13345);
or U18882 (N_18882,N_11700,N_12307);
nand U18883 (N_18883,N_14891,N_11839);
xor U18884 (N_18884,N_12444,N_11956);
xnor U18885 (N_18885,N_10141,N_14703);
nand U18886 (N_18886,N_14978,N_12385);
xnor U18887 (N_18887,N_12882,N_14398);
or U18888 (N_18888,N_12164,N_10583);
xor U18889 (N_18889,N_11669,N_11880);
xor U18890 (N_18890,N_12927,N_13785);
nor U18891 (N_18891,N_10026,N_11790);
xnor U18892 (N_18892,N_14090,N_14313);
or U18893 (N_18893,N_14386,N_13934);
nand U18894 (N_18894,N_10551,N_11243);
nand U18895 (N_18895,N_14008,N_10184);
or U18896 (N_18896,N_14632,N_13618);
xor U18897 (N_18897,N_13116,N_14880);
nor U18898 (N_18898,N_10281,N_10958);
nand U18899 (N_18899,N_11302,N_10936);
nand U18900 (N_18900,N_13415,N_12428);
nor U18901 (N_18901,N_10580,N_10578);
nand U18902 (N_18902,N_10477,N_10878);
nand U18903 (N_18903,N_13167,N_13477);
nor U18904 (N_18904,N_12345,N_10249);
xnor U18905 (N_18905,N_10244,N_12076);
nand U18906 (N_18906,N_10214,N_14136);
or U18907 (N_18907,N_12365,N_12532);
and U18908 (N_18908,N_10719,N_10092);
nor U18909 (N_18909,N_12759,N_10168);
nor U18910 (N_18910,N_12201,N_12491);
or U18911 (N_18911,N_12836,N_12938);
xor U18912 (N_18912,N_13836,N_14441);
or U18913 (N_18913,N_13182,N_13760);
nand U18914 (N_18914,N_14281,N_13950);
or U18915 (N_18915,N_11583,N_12318);
and U18916 (N_18916,N_10704,N_10604);
nor U18917 (N_18917,N_13773,N_13231);
nand U18918 (N_18918,N_14360,N_13917);
nor U18919 (N_18919,N_11963,N_12098);
nand U18920 (N_18920,N_10211,N_10392);
nand U18921 (N_18921,N_10394,N_13544);
or U18922 (N_18922,N_13357,N_11146);
and U18923 (N_18923,N_13791,N_11854);
nand U18924 (N_18924,N_11762,N_14450);
or U18925 (N_18925,N_14454,N_10140);
xnor U18926 (N_18926,N_11884,N_13661);
xor U18927 (N_18927,N_13162,N_13719);
or U18928 (N_18928,N_14632,N_12103);
nor U18929 (N_18929,N_10494,N_12551);
or U18930 (N_18930,N_14612,N_12252);
or U18931 (N_18931,N_11814,N_10938);
nand U18932 (N_18932,N_12265,N_13400);
xnor U18933 (N_18933,N_13047,N_12683);
or U18934 (N_18934,N_13406,N_11686);
nand U18935 (N_18935,N_13613,N_11743);
xnor U18936 (N_18936,N_12295,N_11539);
or U18937 (N_18937,N_12820,N_11464);
nor U18938 (N_18938,N_12807,N_12429);
nor U18939 (N_18939,N_11284,N_11390);
nand U18940 (N_18940,N_10561,N_10164);
and U18941 (N_18941,N_11130,N_11629);
nand U18942 (N_18942,N_10427,N_12265);
or U18943 (N_18943,N_11697,N_11530);
and U18944 (N_18944,N_14496,N_13597);
nor U18945 (N_18945,N_11219,N_12996);
nand U18946 (N_18946,N_10230,N_11913);
xor U18947 (N_18947,N_12799,N_10715);
xnor U18948 (N_18948,N_13045,N_10459);
nand U18949 (N_18949,N_11107,N_13252);
nand U18950 (N_18950,N_14381,N_10109);
xnor U18951 (N_18951,N_11567,N_12873);
nor U18952 (N_18952,N_13028,N_13199);
or U18953 (N_18953,N_10097,N_12912);
nor U18954 (N_18954,N_12976,N_14044);
nand U18955 (N_18955,N_10788,N_13119);
nand U18956 (N_18956,N_14428,N_14091);
xnor U18957 (N_18957,N_12382,N_11388);
xor U18958 (N_18958,N_11029,N_12061);
xnor U18959 (N_18959,N_14839,N_10547);
nand U18960 (N_18960,N_11300,N_10639);
xor U18961 (N_18961,N_11472,N_14530);
nor U18962 (N_18962,N_11227,N_14193);
nand U18963 (N_18963,N_11916,N_11864);
and U18964 (N_18964,N_13550,N_14131);
nor U18965 (N_18965,N_10770,N_14695);
nor U18966 (N_18966,N_12765,N_14494);
and U18967 (N_18967,N_14526,N_11972);
and U18968 (N_18968,N_14509,N_10800);
xor U18969 (N_18969,N_10995,N_14288);
nor U18970 (N_18970,N_13175,N_10901);
xor U18971 (N_18971,N_14235,N_14221);
and U18972 (N_18972,N_14037,N_14277);
xnor U18973 (N_18973,N_12655,N_14292);
nand U18974 (N_18974,N_14656,N_11890);
and U18975 (N_18975,N_10596,N_11621);
nand U18976 (N_18976,N_12317,N_12732);
and U18977 (N_18977,N_11776,N_14250);
nand U18978 (N_18978,N_10801,N_10441);
or U18979 (N_18979,N_13675,N_10686);
xnor U18980 (N_18980,N_11178,N_13434);
nand U18981 (N_18981,N_14360,N_12210);
and U18982 (N_18982,N_10979,N_11048);
and U18983 (N_18983,N_10425,N_14471);
nor U18984 (N_18984,N_12151,N_13433);
xor U18985 (N_18985,N_11462,N_10563);
nand U18986 (N_18986,N_10472,N_11248);
and U18987 (N_18987,N_12608,N_10512);
or U18988 (N_18988,N_14748,N_14144);
xor U18989 (N_18989,N_13010,N_13841);
or U18990 (N_18990,N_10255,N_13608);
nand U18991 (N_18991,N_12503,N_13627);
nor U18992 (N_18992,N_11981,N_14591);
and U18993 (N_18993,N_10516,N_14762);
nor U18994 (N_18994,N_14886,N_14307);
nor U18995 (N_18995,N_10047,N_13047);
and U18996 (N_18996,N_11815,N_14162);
and U18997 (N_18997,N_12892,N_11987);
nand U18998 (N_18998,N_12076,N_11715);
xor U18999 (N_18999,N_10946,N_10234);
or U19000 (N_19000,N_14669,N_13286);
and U19001 (N_19001,N_14310,N_12515);
nor U19002 (N_19002,N_10156,N_13400);
or U19003 (N_19003,N_10705,N_12758);
nand U19004 (N_19004,N_12231,N_14552);
or U19005 (N_19005,N_13922,N_11736);
or U19006 (N_19006,N_12837,N_11225);
or U19007 (N_19007,N_12587,N_13003);
xnor U19008 (N_19008,N_12289,N_13256);
and U19009 (N_19009,N_13702,N_11268);
nand U19010 (N_19010,N_12268,N_14869);
xnor U19011 (N_19011,N_14814,N_13178);
nor U19012 (N_19012,N_10524,N_14346);
nor U19013 (N_19013,N_13200,N_10425);
nand U19014 (N_19014,N_14662,N_13921);
nor U19015 (N_19015,N_10658,N_14136);
nor U19016 (N_19016,N_10488,N_12993);
and U19017 (N_19017,N_10782,N_11231);
nand U19018 (N_19018,N_13754,N_11446);
nor U19019 (N_19019,N_10333,N_10701);
or U19020 (N_19020,N_14413,N_12292);
and U19021 (N_19021,N_11066,N_10479);
xor U19022 (N_19022,N_11236,N_13064);
or U19023 (N_19023,N_12681,N_12542);
nor U19024 (N_19024,N_14297,N_13226);
nand U19025 (N_19025,N_13805,N_14748);
and U19026 (N_19026,N_10016,N_13917);
nand U19027 (N_19027,N_12910,N_11488);
nand U19028 (N_19028,N_14192,N_12891);
and U19029 (N_19029,N_11382,N_11330);
nor U19030 (N_19030,N_10193,N_10434);
nor U19031 (N_19031,N_11758,N_12912);
nor U19032 (N_19032,N_10811,N_14718);
nor U19033 (N_19033,N_11389,N_14908);
nand U19034 (N_19034,N_14516,N_10051);
nand U19035 (N_19035,N_13735,N_10090);
and U19036 (N_19036,N_11213,N_13498);
and U19037 (N_19037,N_13826,N_12690);
nor U19038 (N_19038,N_14371,N_12542);
nand U19039 (N_19039,N_14669,N_11450);
or U19040 (N_19040,N_12543,N_13718);
xor U19041 (N_19041,N_13781,N_11901);
or U19042 (N_19042,N_11760,N_14309);
nand U19043 (N_19043,N_12359,N_12486);
xnor U19044 (N_19044,N_13422,N_13899);
and U19045 (N_19045,N_10168,N_10667);
and U19046 (N_19046,N_11517,N_10841);
xor U19047 (N_19047,N_10778,N_11590);
or U19048 (N_19048,N_14716,N_13103);
or U19049 (N_19049,N_10265,N_11664);
nor U19050 (N_19050,N_14285,N_12917);
xor U19051 (N_19051,N_12191,N_14380);
or U19052 (N_19052,N_13830,N_13299);
and U19053 (N_19053,N_13725,N_14882);
nor U19054 (N_19054,N_13904,N_10166);
nor U19055 (N_19055,N_13474,N_13454);
and U19056 (N_19056,N_14477,N_11609);
or U19057 (N_19057,N_14809,N_14262);
nand U19058 (N_19058,N_13139,N_11408);
or U19059 (N_19059,N_11456,N_13698);
nor U19060 (N_19060,N_12242,N_10547);
nand U19061 (N_19061,N_14218,N_12964);
xnor U19062 (N_19062,N_11572,N_14448);
and U19063 (N_19063,N_10184,N_10745);
or U19064 (N_19064,N_10200,N_13409);
nand U19065 (N_19065,N_10317,N_11507);
nor U19066 (N_19066,N_10124,N_11780);
nand U19067 (N_19067,N_11724,N_13234);
nand U19068 (N_19068,N_12574,N_10278);
xor U19069 (N_19069,N_13173,N_10371);
nor U19070 (N_19070,N_14485,N_14266);
and U19071 (N_19071,N_14814,N_13078);
nor U19072 (N_19072,N_12418,N_14986);
and U19073 (N_19073,N_13606,N_14579);
and U19074 (N_19074,N_14553,N_10338);
or U19075 (N_19075,N_14232,N_10775);
or U19076 (N_19076,N_10054,N_12599);
and U19077 (N_19077,N_14012,N_13462);
xor U19078 (N_19078,N_13026,N_10155);
nor U19079 (N_19079,N_13694,N_12825);
nand U19080 (N_19080,N_11925,N_14277);
nor U19081 (N_19081,N_10017,N_11593);
nor U19082 (N_19082,N_10585,N_12832);
and U19083 (N_19083,N_13570,N_14597);
nor U19084 (N_19084,N_13093,N_13591);
or U19085 (N_19085,N_13163,N_11422);
or U19086 (N_19086,N_10561,N_14361);
or U19087 (N_19087,N_13931,N_11298);
nor U19088 (N_19088,N_10764,N_12691);
nor U19089 (N_19089,N_11624,N_13084);
or U19090 (N_19090,N_11298,N_11888);
and U19091 (N_19091,N_10157,N_14275);
or U19092 (N_19092,N_13409,N_11108);
nand U19093 (N_19093,N_12873,N_14013);
xor U19094 (N_19094,N_10126,N_11225);
nand U19095 (N_19095,N_11485,N_10231);
xor U19096 (N_19096,N_10826,N_10641);
or U19097 (N_19097,N_10668,N_10733);
or U19098 (N_19098,N_12548,N_14304);
xnor U19099 (N_19099,N_13209,N_14125);
nor U19100 (N_19100,N_11682,N_13738);
xnor U19101 (N_19101,N_10211,N_11428);
or U19102 (N_19102,N_12625,N_11726);
and U19103 (N_19103,N_14334,N_13035);
xnor U19104 (N_19104,N_14263,N_11324);
xnor U19105 (N_19105,N_12330,N_12447);
and U19106 (N_19106,N_13597,N_10657);
and U19107 (N_19107,N_11257,N_13605);
xnor U19108 (N_19108,N_11422,N_13843);
and U19109 (N_19109,N_13618,N_13389);
or U19110 (N_19110,N_14641,N_10272);
or U19111 (N_19111,N_13039,N_13652);
nor U19112 (N_19112,N_13854,N_13525);
xnor U19113 (N_19113,N_11985,N_12910);
xor U19114 (N_19114,N_10274,N_10541);
nor U19115 (N_19115,N_13639,N_14775);
nor U19116 (N_19116,N_14639,N_14049);
and U19117 (N_19117,N_13796,N_10491);
or U19118 (N_19118,N_12916,N_14688);
nand U19119 (N_19119,N_13401,N_12106);
and U19120 (N_19120,N_10257,N_10785);
nor U19121 (N_19121,N_13563,N_12375);
xnor U19122 (N_19122,N_13860,N_13388);
nor U19123 (N_19123,N_12466,N_13601);
nand U19124 (N_19124,N_14976,N_10137);
nand U19125 (N_19125,N_11755,N_11006);
or U19126 (N_19126,N_11639,N_11624);
and U19127 (N_19127,N_12920,N_12688);
nor U19128 (N_19128,N_12305,N_11210);
or U19129 (N_19129,N_13095,N_13909);
nand U19130 (N_19130,N_14478,N_13572);
or U19131 (N_19131,N_13149,N_14748);
xor U19132 (N_19132,N_10085,N_10456);
or U19133 (N_19133,N_12389,N_13597);
nand U19134 (N_19134,N_14884,N_13019);
nand U19135 (N_19135,N_13415,N_10233);
xor U19136 (N_19136,N_14691,N_12363);
and U19137 (N_19137,N_12571,N_13647);
or U19138 (N_19138,N_11893,N_12791);
or U19139 (N_19139,N_13907,N_13262);
xor U19140 (N_19140,N_11049,N_14341);
or U19141 (N_19141,N_11057,N_14902);
xnor U19142 (N_19142,N_14355,N_11083);
nand U19143 (N_19143,N_13489,N_13813);
xor U19144 (N_19144,N_12645,N_10547);
nor U19145 (N_19145,N_10921,N_10889);
xnor U19146 (N_19146,N_12585,N_13514);
and U19147 (N_19147,N_11172,N_10209);
nand U19148 (N_19148,N_10944,N_11490);
or U19149 (N_19149,N_12060,N_10980);
xor U19150 (N_19150,N_13304,N_10440);
nand U19151 (N_19151,N_13800,N_10303);
xor U19152 (N_19152,N_13043,N_10628);
or U19153 (N_19153,N_13668,N_11837);
or U19154 (N_19154,N_13272,N_10877);
and U19155 (N_19155,N_11848,N_12383);
or U19156 (N_19156,N_12991,N_14031);
xor U19157 (N_19157,N_14588,N_12547);
xor U19158 (N_19158,N_10816,N_13176);
or U19159 (N_19159,N_14745,N_10680);
nand U19160 (N_19160,N_13250,N_12302);
nand U19161 (N_19161,N_11127,N_11089);
nand U19162 (N_19162,N_13640,N_11653);
xnor U19163 (N_19163,N_13043,N_13738);
or U19164 (N_19164,N_14076,N_14414);
nand U19165 (N_19165,N_12867,N_12718);
nand U19166 (N_19166,N_11258,N_13004);
and U19167 (N_19167,N_11831,N_10120);
nand U19168 (N_19168,N_13340,N_14398);
or U19169 (N_19169,N_10704,N_12668);
or U19170 (N_19170,N_10857,N_14494);
nor U19171 (N_19171,N_13296,N_13501);
and U19172 (N_19172,N_11572,N_14011);
nand U19173 (N_19173,N_14106,N_14910);
nand U19174 (N_19174,N_10121,N_10424);
and U19175 (N_19175,N_12139,N_12059);
xnor U19176 (N_19176,N_12118,N_11061);
nand U19177 (N_19177,N_12302,N_14191);
nand U19178 (N_19178,N_14645,N_10991);
and U19179 (N_19179,N_12104,N_13214);
and U19180 (N_19180,N_13602,N_14264);
and U19181 (N_19181,N_12473,N_13391);
nor U19182 (N_19182,N_14749,N_10658);
nand U19183 (N_19183,N_10508,N_13072);
xor U19184 (N_19184,N_14280,N_10247);
nor U19185 (N_19185,N_13908,N_14391);
nor U19186 (N_19186,N_14322,N_11725);
and U19187 (N_19187,N_10649,N_13097);
nor U19188 (N_19188,N_13689,N_14649);
or U19189 (N_19189,N_13470,N_13169);
nor U19190 (N_19190,N_13982,N_10248);
xor U19191 (N_19191,N_13787,N_12668);
xor U19192 (N_19192,N_11908,N_11891);
and U19193 (N_19193,N_13461,N_11560);
and U19194 (N_19194,N_14727,N_11670);
nor U19195 (N_19195,N_13313,N_10222);
or U19196 (N_19196,N_11721,N_11569);
nor U19197 (N_19197,N_14522,N_13679);
nor U19198 (N_19198,N_14319,N_11834);
nor U19199 (N_19199,N_13059,N_14985);
and U19200 (N_19200,N_12780,N_12899);
nand U19201 (N_19201,N_11062,N_10396);
or U19202 (N_19202,N_14564,N_11281);
or U19203 (N_19203,N_14623,N_10943);
or U19204 (N_19204,N_10567,N_14127);
or U19205 (N_19205,N_11893,N_11071);
nand U19206 (N_19206,N_14764,N_13684);
nand U19207 (N_19207,N_12676,N_12205);
xor U19208 (N_19208,N_14599,N_11137);
nor U19209 (N_19209,N_14058,N_10103);
and U19210 (N_19210,N_12179,N_13519);
and U19211 (N_19211,N_10976,N_11840);
xnor U19212 (N_19212,N_11052,N_12616);
xnor U19213 (N_19213,N_10301,N_13649);
nand U19214 (N_19214,N_10189,N_10163);
or U19215 (N_19215,N_12614,N_13086);
nor U19216 (N_19216,N_14919,N_14287);
or U19217 (N_19217,N_12362,N_13138);
or U19218 (N_19218,N_13317,N_14480);
nor U19219 (N_19219,N_10316,N_11177);
and U19220 (N_19220,N_12733,N_13240);
nand U19221 (N_19221,N_14410,N_14078);
xnor U19222 (N_19222,N_13573,N_11349);
nor U19223 (N_19223,N_12818,N_14194);
xor U19224 (N_19224,N_10058,N_14381);
xor U19225 (N_19225,N_12386,N_14624);
or U19226 (N_19226,N_12534,N_10952);
nor U19227 (N_19227,N_13886,N_11816);
or U19228 (N_19228,N_13290,N_10085);
nor U19229 (N_19229,N_12819,N_12366);
nor U19230 (N_19230,N_14395,N_11166);
nand U19231 (N_19231,N_10037,N_10153);
nor U19232 (N_19232,N_10401,N_12836);
or U19233 (N_19233,N_12949,N_14404);
nor U19234 (N_19234,N_13161,N_10382);
nor U19235 (N_19235,N_10557,N_10325);
nor U19236 (N_19236,N_12645,N_13393);
and U19237 (N_19237,N_10633,N_13111);
or U19238 (N_19238,N_11264,N_11323);
or U19239 (N_19239,N_11394,N_11773);
nand U19240 (N_19240,N_13995,N_12007);
nor U19241 (N_19241,N_14101,N_13113);
or U19242 (N_19242,N_11561,N_14154);
xnor U19243 (N_19243,N_10107,N_14030);
nor U19244 (N_19244,N_12732,N_10105);
nor U19245 (N_19245,N_10884,N_11932);
xnor U19246 (N_19246,N_14098,N_11972);
nand U19247 (N_19247,N_10102,N_11350);
nand U19248 (N_19248,N_13057,N_11175);
xnor U19249 (N_19249,N_13176,N_13846);
xor U19250 (N_19250,N_12493,N_11928);
and U19251 (N_19251,N_10390,N_13953);
nor U19252 (N_19252,N_14536,N_10411);
nor U19253 (N_19253,N_10723,N_14497);
nand U19254 (N_19254,N_11917,N_11551);
nand U19255 (N_19255,N_14445,N_10806);
nor U19256 (N_19256,N_14801,N_14718);
or U19257 (N_19257,N_14447,N_12793);
xnor U19258 (N_19258,N_10762,N_14839);
nand U19259 (N_19259,N_14278,N_12328);
or U19260 (N_19260,N_11538,N_14947);
nand U19261 (N_19261,N_14837,N_13966);
nor U19262 (N_19262,N_10033,N_11917);
nand U19263 (N_19263,N_14810,N_12677);
nor U19264 (N_19264,N_12940,N_13733);
and U19265 (N_19265,N_13770,N_12033);
and U19266 (N_19266,N_13849,N_13563);
or U19267 (N_19267,N_13841,N_11337);
or U19268 (N_19268,N_14261,N_12426);
nand U19269 (N_19269,N_11918,N_10187);
nor U19270 (N_19270,N_12357,N_14610);
xnor U19271 (N_19271,N_14019,N_13057);
nor U19272 (N_19272,N_13987,N_14663);
nand U19273 (N_19273,N_13855,N_14452);
nor U19274 (N_19274,N_12567,N_14470);
xnor U19275 (N_19275,N_10858,N_12061);
nand U19276 (N_19276,N_10378,N_12395);
or U19277 (N_19277,N_10252,N_12461);
or U19278 (N_19278,N_10319,N_11848);
and U19279 (N_19279,N_11318,N_11959);
nor U19280 (N_19280,N_11699,N_14974);
nor U19281 (N_19281,N_11562,N_13802);
nand U19282 (N_19282,N_11961,N_14624);
nand U19283 (N_19283,N_10338,N_12412);
or U19284 (N_19284,N_13589,N_13057);
and U19285 (N_19285,N_10909,N_11646);
and U19286 (N_19286,N_10829,N_10872);
and U19287 (N_19287,N_11176,N_13087);
and U19288 (N_19288,N_10023,N_13655);
nand U19289 (N_19289,N_12055,N_14178);
nand U19290 (N_19290,N_12741,N_14861);
and U19291 (N_19291,N_12082,N_13281);
or U19292 (N_19292,N_14384,N_12281);
xor U19293 (N_19293,N_11363,N_14122);
nor U19294 (N_19294,N_12106,N_13603);
or U19295 (N_19295,N_13272,N_11849);
nand U19296 (N_19296,N_10337,N_10889);
nand U19297 (N_19297,N_12766,N_10091);
and U19298 (N_19298,N_10940,N_14488);
xnor U19299 (N_19299,N_14035,N_12902);
nor U19300 (N_19300,N_11095,N_14978);
and U19301 (N_19301,N_10302,N_10814);
nor U19302 (N_19302,N_10098,N_13931);
nor U19303 (N_19303,N_14558,N_12404);
nand U19304 (N_19304,N_11841,N_11790);
xor U19305 (N_19305,N_14218,N_13612);
or U19306 (N_19306,N_12946,N_14969);
nor U19307 (N_19307,N_14775,N_12866);
nor U19308 (N_19308,N_12054,N_14779);
nand U19309 (N_19309,N_10320,N_14245);
nor U19310 (N_19310,N_13561,N_13241);
or U19311 (N_19311,N_11741,N_12581);
xor U19312 (N_19312,N_14594,N_10453);
or U19313 (N_19313,N_10491,N_10645);
nor U19314 (N_19314,N_11411,N_14401);
nor U19315 (N_19315,N_10003,N_11679);
nand U19316 (N_19316,N_11134,N_14463);
nand U19317 (N_19317,N_11643,N_10369);
or U19318 (N_19318,N_14165,N_11855);
and U19319 (N_19319,N_12856,N_13076);
nor U19320 (N_19320,N_14790,N_14677);
nor U19321 (N_19321,N_11345,N_14025);
nand U19322 (N_19322,N_10857,N_10255);
and U19323 (N_19323,N_12641,N_13144);
and U19324 (N_19324,N_11671,N_11033);
nor U19325 (N_19325,N_11373,N_14021);
or U19326 (N_19326,N_10023,N_12324);
xnor U19327 (N_19327,N_12244,N_11474);
nor U19328 (N_19328,N_13872,N_12266);
and U19329 (N_19329,N_12150,N_12323);
or U19330 (N_19330,N_13048,N_13334);
and U19331 (N_19331,N_13869,N_13136);
nor U19332 (N_19332,N_11012,N_13901);
nor U19333 (N_19333,N_10305,N_11809);
and U19334 (N_19334,N_13509,N_10000);
or U19335 (N_19335,N_13890,N_14161);
or U19336 (N_19336,N_12423,N_14532);
nor U19337 (N_19337,N_10306,N_12685);
nand U19338 (N_19338,N_14076,N_10169);
xnor U19339 (N_19339,N_14525,N_13799);
xnor U19340 (N_19340,N_10776,N_14470);
or U19341 (N_19341,N_14075,N_11159);
nand U19342 (N_19342,N_13850,N_10311);
and U19343 (N_19343,N_11763,N_11009);
nor U19344 (N_19344,N_13517,N_12123);
xnor U19345 (N_19345,N_14013,N_11194);
or U19346 (N_19346,N_13316,N_13565);
or U19347 (N_19347,N_14243,N_13765);
and U19348 (N_19348,N_14815,N_13433);
or U19349 (N_19349,N_13036,N_10818);
and U19350 (N_19350,N_14141,N_13191);
nor U19351 (N_19351,N_10369,N_13128);
xnor U19352 (N_19352,N_14614,N_13733);
nand U19353 (N_19353,N_13650,N_14667);
xor U19354 (N_19354,N_11813,N_14010);
nand U19355 (N_19355,N_11191,N_12460);
nand U19356 (N_19356,N_12485,N_12709);
and U19357 (N_19357,N_10368,N_11780);
or U19358 (N_19358,N_14758,N_11173);
and U19359 (N_19359,N_10622,N_10413);
nand U19360 (N_19360,N_13746,N_10419);
or U19361 (N_19361,N_14120,N_13812);
nand U19362 (N_19362,N_13895,N_12940);
or U19363 (N_19363,N_10318,N_12070);
nand U19364 (N_19364,N_13081,N_11744);
nor U19365 (N_19365,N_14684,N_10928);
xor U19366 (N_19366,N_12041,N_13313);
and U19367 (N_19367,N_13852,N_11841);
nor U19368 (N_19368,N_13675,N_13256);
nor U19369 (N_19369,N_13263,N_14530);
or U19370 (N_19370,N_10866,N_13957);
xor U19371 (N_19371,N_10739,N_12865);
or U19372 (N_19372,N_10429,N_13707);
xnor U19373 (N_19373,N_11886,N_12690);
nand U19374 (N_19374,N_14432,N_11186);
and U19375 (N_19375,N_10387,N_12209);
nand U19376 (N_19376,N_10526,N_13174);
and U19377 (N_19377,N_13714,N_11082);
nor U19378 (N_19378,N_14213,N_14643);
xnor U19379 (N_19379,N_14934,N_10613);
nand U19380 (N_19380,N_14150,N_13659);
and U19381 (N_19381,N_10726,N_11833);
nand U19382 (N_19382,N_10691,N_11397);
xor U19383 (N_19383,N_10504,N_10716);
nand U19384 (N_19384,N_13946,N_11064);
xor U19385 (N_19385,N_13092,N_12910);
nand U19386 (N_19386,N_12065,N_14975);
xnor U19387 (N_19387,N_12593,N_12858);
nand U19388 (N_19388,N_11881,N_14865);
and U19389 (N_19389,N_14035,N_10294);
or U19390 (N_19390,N_13664,N_14210);
nand U19391 (N_19391,N_12409,N_13952);
xor U19392 (N_19392,N_13887,N_11153);
nor U19393 (N_19393,N_11497,N_13690);
xor U19394 (N_19394,N_11565,N_12270);
or U19395 (N_19395,N_10865,N_12588);
xnor U19396 (N_19396,N_14000,N_10119);
and U19397 (N_19397,N_11460,N_14207);
xnor U19398 (N_19398,N_10195,N_10720);
xnor U19399 (N_19399,N_11112,N_10879);
or U19400 (N_19400,N_12254,N_13357);
nor U19401 (N_19401,N_14156,N_14592);
nor U19402 (N_19402,N_10809,N_13335);
and U19403 (N_19403,N_13091,N_14065);
nor U19404 (N_19404,N_11716,N_14231);
nand U19405 (N_19405,N_11531,N_11017);
xor U19406 (N_19406,N_13175,N_10593);
xnor U19407 (N_19407,N_11351,N_14397);
or U19408 (N_19408,N_11336,N_13453);
xnor U19409 (N_19409,N_11585,N_13051);
or U19410 (N_19410,N_10102,N_11570);
nor U19411 (N_19411,N_14382,N_13208);
and U19412 (N_19412,N_11634,N_12577);
xnor U19413 (N_19413,N_10700,N_11498);
or U19414 (N_19414,N_11027,N_13904);
or U19415 (N_19415,N_11767,N_13237);
nand U19416 (N_19416,N_10367,N_12515);
nor U19417 (N_19417,N_12735,N_12927);
nor U19418 (N_19418,N_12530,N_13859);
or U19419 (N_19419,N_11853,N_10328);
and U19420 (N_19420,N_10471,N_10723);
or U19421 (N_19421,N_10053,N_12048);
and U19422 (N_19422,N_12553,N_13877);
nand U19423 (N_19423,N_11192,N_13183);
or U19424 (N_19424,N_14409,N_13007);
xnor U19425 (N_19425,N_10713,N_11439);
nor U19426 (N_19426,N_13393,N_12157);
or U19427 (N_19427,N_10034,N_12260);
or U19428 (N_19428,N_14103,N_11556);
and U19429 (N_19429,N_10796,N_12959);
nand U19430 (N_19430,N_10094,N_14699);
xnor U19431 (N_19431,N_14905,N_14052);
nor U19432 (N_19432,N_10127,N_10571);
and U19433 (N_19433,N_14535,N_13024);
xor U19434 (N_19434,N_12110,N_11428);
or U19435 (N_19435,N_11037,N_10870);
nand U19436 (N_19436,N_12187,N_10186);
nor U19437 (N_19437,N_10564,N_12392);
and U19438 (N_19438,N_10494,N_13140);
and U19439 (N_19439,N_12182,N_14439);
and U19440 (N_19440,N_13660,N_14817);
nand U19441 (N_19441,N_14165,N_14029);
and U19442 (N_19442,N_10928,N_12015);
nand U19443 (N_19443,N_10877,N_10417);
xnor U19444 (N_19444,N_12268,N_11741);
and U19445 (N_19445,N_10912,N_14328);
and U19446 (N_19446,N_11871,N_12564);
nor U19447 (N_19447,N_11078,N_12742);
and U19448 (N_19448,N_10133,N_11329);
nand U19449 (N_19449,N_10690,N_12797);
or U19450 (N_19450,N_12955,N_10383);
nor U19451 (N_19451,N_14478,N_10056);
nand U19452 (N_19452,N_12839,N_11082);
or U19453 (N_19453,N_12371,N_11451);
xor U19454 (N_19454,N_10247,N_14658);
and U19455 (N_19455,N_10997,N_11922);
and U19456 (N_19456,N_12762,N_14601);
and U19457 (N_19457,N_10841,N_12648);
and U19458 (N_19458,N_12531,N_10672);
xnor U19459 (N_19459,N_13304,N_14803);
and U19460 (N_19460,N_11855,N_13503);
nor U19461 (N_19461,N_11401,N_13565);
nand U19462 (N_19462,N_10324,N_12794);
nor U19463 (N_19463,N_10919,N_13545);
nand U19464 (N_19464,N_14009,N_11362);
or U19465 (N_19465,N_12449,N_10909);
and U19466 (N_19466,N_14200,N_14760);
and U19467 (N_19467,N_11758,N_14665);
or U19468 (N_19468,N_14555,N_13259);
or U19469 (N_19469,N_12052,N_14094);
nor U19470 (N_19470,N_13606,N_12169);
nor U19471 (N_19471,N_14082,N_11348);
xnor U19472 (N_19472,N_14142,N_14211);
or U19473 (N_19473,N_14902,N_11459);
or U19474 (N_19474,N_13320,N_13030);
or U19475 (N_19475,N_11245,N_13815);
nor U19476 (N_19476,N_11759,N_12327);
and U19477 (N_19477,N_13948,N_10508);
or U19478 (N_19478,N_12591,N_11050);
nor U19479 (N_19479,N_12653,N_10410);
and U19480 (N_19480,N_12918,N_12406);
nor U19481 (N_19481,N_10417,N_13478);
and U19482 (N_19482,N_14298,N_13918);
xnor U19483 (N_19483,N_13477,N_11557);
and U19484 (N_19484,N_13701,N_12285);
xor U19485 (N_19485,N_12299,N_10986);
nor U19486 (N_19486,N_12033,N_12558);
nor U19487 (N_19487,N_11653,N_12584);
or U19488 (N_19488,N_13668,N_12873);
or U19489 (N_19489,N_10665,N_11289);
xnor U19490 (N_19490,N_11566,N_12481);
nor U19491 (N_19491,N_10918,N_14860);
nor U19492 (N_19492,N_11586,N_11324);
xnor U19493 (N_19493,N_13370,N_14761);
nor U19494 (N_19494,N_14911,N_12560);
xnor U19495 (N_19495,N_11430,N_10849);
nand U19496 (N_19496,N_10049,N_12219);
or U19497 (N_19497,N_12101,N_13397);
nor U19498 (N_19498,N_14837,N_14828);
nor U19499 (N_19499,N_14642,N_10919);
nand U19500 (N_19500,N_13812,N_13127);
xnor U19501 (N_19501,N_12457,N_11470);
or U19502 (N_19502,N_14509,N_12573);
xnor U19503 (N_19503,N_13612,N_13417);
and U19504 (N_19504,N_10945,N_10122);
nand U19505 (N_19505,N_11716,N_13608);
nor U19506 (N_19506,N_13380,N_12012);
and U19507 (N_19507,N_14171,N_12724);
nor U19508 (N_19508,N_13950,N_10572);
or U19509 (N_19509,N_13895,N_14015);
or U19510 (N_19510,N_13969,N_10123);
or U19511 (N_19511,N_14341,N_11027);
nor U19512 (N_19512,N_11570,N_10544);
and U19513 (N_19513,N_10869,N_10506);
nor U19514 (N_19514,N_10242,N_12587);
and U19515 (N_19515,N_13208,N_10211);
and U19516 (N_19516,N_12408,N_13085);
nor U19517 (N_19517,N_10931,N_11061);
and U19518 (N_19518,N_13610,N_14306);
or U19519 (N_19519,N_12956,N_11682);
or U19520 (N_19520,N_11950,N_10908);
nand U19521 (N_19521,N_12600,N_14300);
nand U19522 (N_19522,N_13498,N_13156);
or U19523 (N_19523,N_13007,N_14444);
nor U19524 (N_19524,N_12686,N_13064);
or U19525 (N_19525,N_13578,N_14605);
or U19526 (N_19526,N_12647,N_12606);
nor U19527 (N_19527,N_13945,N_12278);
nor U19528 (N_19528,N_13617,N_13273);
nor U19529 (N_19529,N_12182,N_12610);
or U19530 (N_19530,N_14442,N_11332);
nand U19531 (N_19531,N_10252,N_14619);
or U19532 (N_19532,N_14311,N_10841);
xnor U19533 (N_19533,N_10360,N_12261);
or U19534 (N_19534,N_12658,N_13648);
nand U19535 (N_19535,N_12509,N_13451);
xor U19536 (N_19536,N_13817,N_12942);
xnor U19537 (N_19537,N_13603,N_10955);
and U19538 (N_19538,N_11298,N_12401);
nand U19539 (N_19539,N_10927,N_14527);
nor U19540 (N_19540,N_13547,N_13640);
nor U19541 (N_19541,N_11779,N_14383);
nor U19542 (N_19542,N_11889,N_13291);
xor U19543 (N_19543,N_12520,N_13118);
or U19544 (N_19544,N_12025,N_12883);
xnor U19545 (N_19545,N_13738,N_14129);
nor U19546 (N_19546,N_14096,N_12040);
and U19547 (N_19547,N_10727,N_10227);
nand U19548 (N_19548,N_12275,N_12670);
nand U19549 (N_19549,N_14455,N_11539);
nand U19550 (N_19550,N_14592,N_13946);
and U19551 (N_19551,N_14939,N_10864);
nor U19552 (N_19552,N_10579,N_14858);
nand U19553 (N_19553,N_10527,N_10375);
and U19554 (N_19554,N_11561,N_14853);
nand U19555 (N_19555,N_14658,N_11180);
nor U19556 (N_19556,N_12887,N_12906);
xnor U19557 (N_19557,N_14662,N_11570);
nand U19558 (N_19558,N_14536,N_10716);
nor U19559 (N_19559,N_10277,N_12964);
nand U19560 (N_19560,N_14811,N_14739);
nand U19561 (N_19561,N_14066,N_10856);
or U19562 (N_19562,N_14512,N_12009);
xnor U19563 (N_19563,N_14988,N_12802);
xnor U19564 (N_19564,N_10158,N_14081);
xnor U19565 (N_19565,N_13357,N_12494);
and U19566 (N_19566,N_13267,N_10262);
and U19567 (N_19567,N_10254,N_10932);
nand U19568 (N_19568,N_11520,N_10613);
and U19569 (N_19569,N_12942,N_11917);
nand U19570 (N_19570,N_11710,N_14539);
nand U19571 (N_19571,N_10619,N_14499);
and U19572 (N_19572,N_13442,N_13579);
nand U19573 (N_19573,N_13165,N_14001);
nor U19574 (N_19574,N_10378,N_13639);
or U19575 (N_19575,N_14266,N_11157);
nor U19576 (N_19576,N_14851,N_14055);
nand U19577 (N_19577,N_11423,N_13762);
or U19578 (N_19578,N_11619,N_10227);
or U19579 (N_19579,N_12935,N_10715);
or U19580 (N_19580,N_10924,N_11148);
nor U19581 (N_19581,N_10280,N_12962);
xor U19582 (N_19582,N_12103,N_11801);
nor U19583 (N_19583,N_13031,N_12267);
and U19584 (N_19584,N_12858,N_10590);
xor U19585 (N_19585,N_10920,N_10784);
or U19586 (N_19586,N_14851,N_11272);
nor U19587 (N_19587,N_12342,N_13549);
xnor U19588 (N_19588,N_10364,N_14653);
nor U19589 (N_19589,N_13713,N_14930);
nand U19590 (N_19590,N_13663,N_10995);
xor U19591 (N_19591,N_13093,N_11894);
nand U19592 (N_19592,N_12768,N_14418);
or U19593 (N_19593,N_10866,N_12771);
xnor U19594 (N_19594,N_14548,N_11811);
nor U19595 (N_19595,N_14462,N_10028);
xor U19596 (N_19596,N_14165,N_14592);
nor U19597 (N_19597,N_10567,N_13527);
and U19598 (N_19598,N_13123,N_11141);
and U19599 (N_19599,N_12315,N_12704);
nor U19600 (N_19600,N_10712,N_12498);
xor U19601 (N_19601,N_10551,N_12782);
nand U19602 (N_19602,N_12993,N_13139);
and U19603 (N_19603,N_13288,N_11045);
nor U19604 (N_19604,N_14342,N_14818);
nand U19605 (N_19605,N_12767,N_13724);
nor U19606 (N_19606,N_11870,N_13588);
nor U19607 (N_19607,N_10088,N_13959);
nand U19608 (N_19608,N_11306,N_10823);
nor U19609 (N_19609,N_10640,N_11334);
or U19610 (N_19610,N_14646,N_14703);
and U19611 (N_19611,N_11623,N_14091);
nor U19612 (N_19612,N_11497,N_14509);
and U19613 (N_19613,N_10987,N_12223);
or U19614 (N_19614,N_10997,N_12203);
nor U19615 (N_19615,N_10605,N_14382);
and U19616 (N_19616,N_12746,N_10533);
nand U19617 (N_19617,N_14772,N_11767);
or U19618 (N_19618,N_12872,N_10591);
nand U19619 (N_19619,N_13965,N_10043);
nor U19620 (N_19620,N_13881,N_14189);
or U19621 (N_19621,N_10869,N_13604);
or U19622 (N_19622,N_12166,N_12835);
nand U19623 (N_19623,N_13641,N_14605);
or U19624 (N_19624,N_14748,N_14883);
xnor U19625 (N_19625,N_10369,N_11365);
nor U19626 (N_19626,N_14742,N_11056);
and U19627 (N_19627,N_14399,N_12888);
nand U19628 (N_19628,N_11446,N_11174);
nand U19629 (N_19629,N_14148,N_12550);
xor U19630 (N_19630,N_10462,N_10465);
and U19631 (N_19631,N_11696,N_14835);
nor U19632 (N_19632,N_10158,N_11277);
nand U19633 (N_19633,N_14688,N_14544);
nand U19634 (N_19634,N_14130,N_11539);
nor U19635 (N_19635,N_12138,N_11877);
nor U19636 (N_19636,N_14887,N_13506);
xor U19637 (N_19637,N_11476,N_13220);
xor U19638 (N_19638,N_10885,N_12900);
nand U19639 (N_19639,N_13120,N_12206);
or U19640 (N_19640,N_11360,N_13323);
or U19641 (N_19641,N_11063,N_10730);
nand U19642 (N_19642,N_13084,N_14787);
nand U19643 (N_19643,N_10844,N_12512);
xor U19644 (N_19644,N_12848,N_13694);
or U19645 (N_19645,N_14920,N_10816);
nand U19646 (N_19646,N_10533,N_14551);
nand U19647 (N_19647,N_10832,N_10392);
nand U19648 (N_19648,N_12539,N_11209);
nand U19649 (N_19649,N_10345,N_10374);
nand U19650 (N_19650,N_13860,N_12419);
nor U19651 (N_19651,N_10054,N_11014);
and U19652 (N_19652,N_11395,N_10394);
xnor U19653 (N_19653,N_14280,N_10914);
nand U19654 (N_19654,N_12240,N_11552);
xnor U19655 (N_19655,N_10171,N_11619);
nor U19656 (N_19656,N_11582,N_12260);
nand U19657 (N_19657,N_13109,N_14183);
xor U19658 (N_19658,N_10848,N_11279);
or U19659 (N_19659,N_13051,N_14417);
nand U19660 (N_19660,N_12560,N_14325);
nand U19661 (N_19661,N_12472,N_14598);
nor U19662 (N_19662,N_13406,N_10842);
nand U19663 (N_19663,N_11521,N_13402);
or U19664 (N_19664,N_12436,N_12632);
nand U19665 (N_19665,N_11400,N_14849);
nor U19666 (N_19666,N_10298,N_12107);
and U19667 (N_19667,N_11022,N_13761);
nand U19668 (N_19668,N_14073,N_12572);
xnor U19669 (N_19669,N_11386,N_12426);
nor U19670 (N_19670,N_13564,N_10497);
nand U19671 (N_19671,N_12881,N_11390);
nor U19672 (N_19672,N_11342,N_14557);
nor U19673 (N_19673,N_12970,N_12846);
nand U19674 (N_19674,N_14274,N_14033);
nand U19675 (N_19675,N_10714,N_13664);
xnor U19676 (N_19676,N_13668,N_11224);
or U19677 (N_19677,N_14886,N_14333);
nand U19678 (N_19678,N_12469,N_12107);
nand U19679 (N_19679,N_14054,N_11881);
xnor U19680 (N_19680,N_13686,N_10170);
xor U19681 (N_19681,N_12689,N_10694);
nand U19682 (N_19682,N_11579,N_13062);
and U19683 (N_19683,N_10070,N_11123);
xor U19684 (N_19684,N_11639,N_13229);
or U19685 (N_19685,N_12249,N_13443);
xnor U19686 (N_19686,N_14779,N_13066);
nand U19687 (N_19687,N_13175,N_12218);
nor U19688 (N_19688,N_14221,N_10806);
or U19689 (N_19689,N_10526,N_10601);
and U19690 (N_19690,N_10247,N_12746);
nand U19691 (N_19691,N_13156,N_10340);
and U19692 (N_19692,N_10106,N_14806);
xor U19693 (N_19693,N_11747,N_13032);
or U19694 (N_19694,N_13836,N_12472);
and U19695 (N_19695,N_12938,N_13294);
or U19696 (N_19696,N_10107,N_12544);
nor U19697 (N_19697,N_10494,N_12755);
nand U19698 (N_19698,N_14066,N_11140);
xor U19699 (N_19699,N_14433,N_12290);
xor U19700 (N_19700,N_11814,N_14098);
nor U19701 (N_19701,N_14336,N_11715);
and U19702 (N_19702,N_12592,N_13035);
nor U19703 (N_19703,N_13156,N_12980);
and U19704 (N_19704,N_10449,N_11377);
nor U19705 (N_19705,N_12279,N_14905);
xor U19706 (N_19706,N_14547,N_11970);
xnor U19707 (N_19707,N_13851,N_10620);
xnor U19708 (N_19708,N_13959,N_14477);
nand U19709 (N_19709,N_14239,N_11604);
or U19710 (N_19710,N_12479,N_12631);
nand U19711 (N_19711,N_14249,N_14529);
xor U19712 (N_19712,N_14761,N_10635);
or U19713 (N_19713,N_13454,N_14766);
xnor U19714 (N_19714,N_12162,N_12014);
xnor U19715 (N_19715,N_11252,N_13033);
nor U19716 (N_19716,N_11397,N_14922);
or U19717 (N_19717,N_14302,N_11908);
nand U19718 (N_19718,N_13630,N_13244);
xor U19719 (N_19719,N_12586,N_10176);
nand U19720 (N_19720,N_13685,N_10654);
nor U19721 (N_19721,N_14901,N_11158);
nor U19722 (N_19722,N_13293,N_11999);
nand U19723 (N_19723,N_14933,N_13814);
or U19724 (N_19724,N_11326,N_13926);
xnor U19725 (N_19725,N_13551,N_11380);
nor U19726 (N_19726,N_12054,N_14474);
nor U19727 (N_19727,N_10059,N_12747);
nand U19728 (N_19728,N_12744,N_11856);
and U19729 (N_19729,N_12389,N_11600);
and U19730 (N_19730,N_10536,N_10118);
and U19731 (N_19731,N_11704,N_13849);
nor U19732 (N_19732,N_12292,N_12231);
xor U19733 (N_19733,N_14746,N_13261);
and U19734 (N_19734,N_13391,N_12658);
nor U19735 (N_19735,N_14530,N_13060);
nor U19736 (N_19736,N_11470,N_11523);
xnor U19737 (N_19737,N_13421,N_13148);
nand U19738 (N_19738,N_14911,N_14616);
xnor U19739 (N_19739,N_10380,N_10907);
or U19740 (N_19740,N_14024,N_12279);
nand U19741 (N_19741,N_10344,N_10449);
nand U19742 (N_19742,N_10097,N_14321);
xnor U19743 (N_19743,N_12803,N_11114);
xnor U19744 (N_19744,N_11848,N_12785);
xnor U19745 (N_19745,N_14115,N_10970);
or U19746 (N_19746,N_12868,N_10744);
and U19747 (N_19747,N_10513,N_10762);
nor U19748 (N_19748,N_12765,N_11370);
nor U19749 (N_19749,N_11157,N_12625);
and U19750 (N_19750,N_11019,N_11674);
nand U19751 (N_19751,N_11093,N_10016);
nand U19752 (N_19752,N_11546,N_10545);
nor U19753 (N_19753,N_12126,N_12799);
and U19754 (N_19754,N_10713,N_13686);
nand U19755 (N_19755,N_14206,N_10129);
nand U19756 (N_19756,N_13935,N_13619);
or U19757 (N_19757,N_12762,N_12144);
nor U19758 (N_19758,N_12203,N_10447);
nor U19759 (N_19759,N_14856,N_13612);
nor U19760 (N_19760,N_13796,N_10341);
nand U19761 (N_19761,N_10832,N_12421);
or U19762 (N_19762,N_13604,N_13589);
xnor U19763 (N_19763,N_11925,N_13981);
and U19764 (N_19764,N_14855,N_10035);
nand U19765 (N_19765,N_13985,N_12836);
and U19766 (N_19766,N_13387,N_14477);
and U19767 (N_19767,N_12878,N_10606);
or U19768 (N_19768,N_10479,N_11840);
nand U19769 (N_19769,N_14129,N_10196);
and U19770 (N_19770,N_12828,N_12623);
and U19771 (N_19771,N_10505,N_10339);
nor U19772 (N_19772,N_12005,N_11627);
or U19773 (N_19773,N_13382,N_13718);
nor U19774 (N_19774,N_14913,N_10589);
xor U19775 (N_19775,N_13185,N_12850);
or U19776 (N_19776,N_11355,N_13719);
nand U19777 (N_19777,N_12483,N_12086);
or U19778 (N_19778,N_10318,N_12751);
nand U19779 (N_19779,N_11449,N_13247);
nor U19780 (N_19780,N_14370,N_12044);
nand U19781 (N_19781,N_11983,N_12408);
xor U19782 (N_19782,N_10957,N_13330);
nand U19783 (N_19783,N_12169,N_11446);
and U19784 (N_19784,N_12278,N_11354);
and U19785 (N_19785,N_11962,N_12697);
xnor U19786 (N_19786,N_11653,N_11189);
or U19787 (N_19787,N_13721,N_11755);
nand U19788 (N_19788,N_10950,N_10306);
nor U19789 (N_19789,N_12893,N_12116);
xor U19790 (N_19790,N_12299,N_10734);
and U19791 (N_19791,N_11986,N_14648);
and U19792 (N_19792,N_11983,N_11013);
nand U19793 (N_19793,N_11331,N_10886);
and U19794 (N_19794,N_10371,N_13629);
and U19795 (N_19795,N_14641,N_10160);
or U19796 (N_19796,N_14887,N_14693);
nor U19797 (N_19797,N_10676,N_14660);
nand U19798 (N_19798,N_11879,N_12795);
nor U19799 (N_19799,N_13781,N_12509);
xnor U19800 (N_19800,N_12307,N_10659);
nor U19801 (N_19801,N_12373,N_10845);
or U19802 (N_19802,N_13424,N_13989);
xnor U19803 (N_19803,N_13044,N_11203);
nand U19804 (N_19804,N_14131,N_14519);
nor U19805 (N_19805,N_10084,N_10712);
and U19806 (N_19806,N_10343,N_11436);
nand U19807 (N_19807,N_10044,N_12677);
nor U19808 (N_19808,N_12199,N_12803);
nand U19809 (N_19809,N_14757,N_12322);
xnor U19810 (N_19810,N_11506,N_14073);
xnor U19811 (N_19811,N_14612,N_13359);
nand U19812 (N_19812,N_11587,N_13516);
nand U19813 (N_19813,N_11147,N_10688);
or U19814 (N_19814,N_14335,N_11791);
and U19815 (N_19815,N_10504,N_13639);
nor U19816 (N_19816,N_12722,N_14000);
nand U19817 (N_19817,N_10275,N_10697);
or U19818 (N_19818,N_11502,N_10384);
nand U19819 (N_19819,N_12446,N_12874);
nor U19820 (N_19820,N_13263,N_13674);
and U19821 (N_19821,N_10433,N_14391);
and U19822 (N_19822,N_11417,N_10058);
and U19823 (N_19823,N_10380,N_10725);
and U19824 (N_19824,N_12364,N_12842);
xnor U19825 (N_19825,N_10325,N_13614);
xor U19826 (N_19826,N_12463,N_14529);
and U19827 (N_19827,N_10216,N_10056);
or U19828 (N_19828,N_12362,N_12122);
and U19829 (N_19829,N_10991,N_11536);
or U19830 (N_19830,N_10237,N_11175);
nor U19831 (N_19831,N_12378,N_13438);
and U19832 (N_19832,N_14219,N_11774);
nor U19833 (N_19833,N_10404,N_12636);
nor U19834 (N_19834,N_10582,N_10108);
and U19835 (N_19835,N_12737,N_11916);
nor U19836 (N_19836,N_14774,N_10048);
or U19837 (N_19837,N_13055,N_14553);
xor U19838 (N_19838,N_10102,N_10191);
and U19839 (N_19839,N_10381,N_13139);
and U19840 (N_19840,N_12726,N_11069);
and U19841 (N_19841,N_12729,N_11218);
nor U19842 (N_19842,N_11540,N_12021);
or U19843 (N_19843,N_10532,N_10982);
nand U19844 (N_19844,N_12115,N_13674);
or U19845 (N_19845,N_12251,N_10479);
and U19846 (N_19846,N_12299,N_11135);
or U19847 (N_19847,N_14283,N_10186);
nand U19848 (N_19848,N_14964,N_11230);
xor U19849 (N_19849,N_13980,N_10685);
and U19850 (N_19850,N_10339,N_10433);
or U19851 (N_19851,N_13500,N_10070);
nor U19852 (N_19852,N_13101,N_14270);
or U19853 (N_19853,N_10070,N_12636);
xnor U19854 (N_19854,N_11878,N_11976);
or U19855 (N_19855,N_11575,N_14187);
and U19856 (N_19856,N_13460,N_14859);
nor U19857 (N_19857,N_12935,N_10004);
xnor U19858 (N_19858,N_10862,N_12663);
nor U19859 (N_19859,N_12628,N_13296);
xnor U19860 (N_19860,N_10283,N_14315);
and U19861 (N_19861,N_11151,N_11760);
nand U19862 (N_19862,N_12188,N_12799);
xor U19863 (N_19863,N_11108,N_11989);
nor U19864 (N_19864,N_11112,N_13064);
xnor U19865 (N_19865,N_10433,N_14184);
and U19866 (N_19866,N_10028,N_14426);
xor U19867 (N_19867,N_10333,N_13196);
and U19868 (N_19868,N_11392,N_11893);
nand U19869 (N_19869,N_14896,N_10027);
and U19870 (N_19870,N_14029,N_12004);
nand U19871 (N_19871,N_14740,N_10744);
and U19872 (N_19872,N_10879,N_10712);
or U19873 (N_19873,N_12919,N_13838);
nand U19874 (N_19874,N_11592,N_11222);
or U19875 (N_19875,N_14930,N_10060);
or U19876 (N_19876,N_12598,N_11028);
nand U19877 (N_19877,N_12461,N_11634);
and U19878 (N_19878,N_10550,N_14003);
nor U19879 (N_19879,N_14032,N_11324);
nand U19880 (N_19880,N_13538,N_12848);
and U19881 (N_19881,N_14111,N_10080);
nand U19882 (N_19882,N_12965,N_13474);
or U19883 (N_19883,N_11258,N_13663);
nor U19884 (N_19884,N_12040,N_12716);
nor U19885 (N_19885,N_11847,N_11124);
xnor U19886 (N_19886,N_14087,N_10756);
or U19887 (N_19887,N_12792,N_14944);
nand U19888 (N_19888,N_11401,N_10259);
xor U19889 (N_19889,N_10894,N_10652);
xnor U19890 (N_19890,N_14793,N_14133);
and U19891 (N_19891,N_12684,N_10757);
xnor U19892 (N_19892,N_11660,N_11188);
and U19893 (N_19893,N_14574,N_11307);
and U19894 (N_19894,N_13136,N_12299);
xor U19895 (N_19895,N_10759,N_13646);
nand U19896 (N_19896,N_11676,N_14961);
and U19897 (N_19897,N_12466,N_14527);
nand U19898 (N_19898,N_11195,N_13808);
nor U19899 (N_19899,N_14480,N_10701);
or U19900 (N_19900,N_13523,N_13434);
and U19901 (N_19901,N_10818,N_14641);
nand U19902 (N_19902,N_14020,N_12973);
nand U19903 (N_19903,N_12974,N_14125);
xnor U19904 (N_19904,N_13356,N_13195);
and U19905 (N_19905,N_12770,N_11749);
nor U19906 (N_19906,N_14184,N_14549);
nand U19907 (N_19907,N_11352,N_13110);
or U19908 (N_19908,N_12729,N_11765);
xor U19909 (N_19909,N_11571,N_11750);
or U19910 (N_19910,N_10547,N_13238);
xor U19911 (N_19911,N_13257,N_11565);
nor U19912 (N_19912,N_14763,N_14285);
xnor U19913 (N_19913,N_13514,N_14185);
or U19914 (N_19914,N_13546,N_11045);
nor U19915 (N_19915,N_14303,N_11496);
nand U19916 (N_19916,N_12809,N_14557);
nor U19917 (N_19917,N_11137,N_12527);
or U19918 (N_19918,N_12664,N_14248);
nor U19919 (N_19919,N_12030,N_10414);
and U19920 (N_19920,N_11446,N_13435);
and U19921 (N_19921,N_14603,N_12881);
nand U19922 (N_19922,N_11540,N_14118);
xor U19923 (N_19923,N_12035,N_12941);
nor U19924 (N_19924,N_14208,N_13784);
or U19925 (N_19925,N_11418,N_10992);
nand U19926 (N_19926,N_12694,N_12629);
and U19927 (N_19927,N_10611,N_12996);
and U19928 (N_19928,N_11997,N_11172);
or U19929 (N_19929,N_14942,N_12558);
nor U19930 (N_19930,N_14122,N_10096);
nor U19931 (N_19931,N_14410,N_13222);
or U19932 (N_19932,N_11526,N_11488);
nand U19933 (N_19933,N_14329,N_14388);
or U19934 (N_19934,N_13202,N_10110);
nor U19935 (N_19935,N_13452,N_10109);
xnor U19936 (N_19936,N_11239,N_10394);
nor U19937 (N_19937,N_10669,N_14137);
nand U19938 (N_19938,N_12666,N_13934);
nor U19939 (N_19939,N_12679,N_11934);
and U19940 (N_19940,N_13106,N_10091);
nor U19941 (N_19941,N_14689,N_10630);
nor U19942 (N_19942,N_12685,N_13589);
nand U19943 (N_19943,N_10451,N_13650);
nand U19944 (N_19944,N_10526,N_12092);
nor U19945 (N_19945,N_12909,N_11381);
and U19946 (N_19946,N_14530,N_12944);
and U19947 (N_19947,N_13283,N_13513);
nor U19948 (N_19948,N_12536,N_10801);
nand U19949 (N_19949,N_13366,N_13309);
nor U19950 (N_19950,N_10639,N_10202);
xor U19951 (N_19951,N_11533,N_14486);
and U19952 (N_19952,N_14957,N_11347);
nor U19953 (N_19953,N_13988,N_12939);
nor U19954 (N_19954,N_10219,N_14271);
nor U19955 (N_19955,N_12985,N_10000);
nor U19956 (N_19956,N_14147,N_12883);
nor U19957 (N_19957,N_12875,N_11926);
nor U19958 (N_19958,N_14250,N_14420);
nand U19959 (N_19959,N_11231,N_13853);
and U19960 (N_19960,N_10324,N_13722);
nand U19961 (N_19961,N_14263,N_11530);
or U19962 (N_19962,N_10220,N_13834);
and U19963 (N_19963,N_13710,N_14252);
or U19964 (N_19964,N_13853,N_12498);
xor U19965 (N_19965,N_13651,N_14787);
xor U19966 (N_19966,N_11659,N_14602);
nor U19967 (N_19967,N_13639,N_14584);
or U19968 (N_19968,N_10314,N_10895);
xnor U19969 (N_19969,N_14443,N_11124);
nand U19970 (N_19970,N_10064,N_14298);
nor U19971 (N_19971,N_12381,N_13047);
or U19972 (N_19972,N_11989,N_12526);
nor U19973 (N_19973,N_14409,N_13172);
nand U19974 (N_19974,N_12659,N_14707);
xnor U19975 (N_19975,N_10714,N_13146);
and U19976 (N_19976,N_11335,N_13378);
or U19977 (N_19977,N_14216,N_14941);
xor U19978 (N_19978,N_10029,N_12885);
nor U19979 (N_19979,N_14406,N_13070);
or U19980 (N_19980,N_13317,N_13983);
xor U19981 (N_19981,N_14575,N_10252);
and U19982 (N_19982,N_10360,N_13002);
xnor U19983 (N_19983,N_14394,N_14904);
or U19984 (N_19984,N_13674,N_13667);
xnor U19985 (N_19985,N_11752,N_13444);
or U19986 (N_19986,N_11506,N_10890);
nand U19987 (N_19987,N_14408,N_14963);
and U19988 (N_19988,N_14103,N_11594);
or U19989 (N_19989,N_12776,N_11829);
and U19990 (N_19990,N_11507,N_12530);
xor U19991 (N_19991,N_13041,N_14153);
nand U19992 (N_19992,N_14807,N_13670);
or U19993 (N_19993,N_14062,N_12854);
xor U19994 (N_19994,N_12543,N_13221);
and U19995 (N_19995,N_10439,N_10924);
nand U19996 (N_19996,N_11583,N_11401);
xnor U19997 (N_19997,N_14706,N_10414);
or U19998 (N_19998,N_14487,N_10559);
or U19999 (N_19999,N_10402,N_12922);
and U20000 (N_20000,N_19865,N_18964);
or U20001 (N_20001,N_19230,N_19703);
and U20002 (N_20002,N_16409,N_18788);
or U20003 (N_20003,N_19925,N_16395);
and U20004 (N_20004,N_17158,N_18388);
or U20005 (N_20005,N_19275,N_16877);
nor U20006 (N_20006,N_18160,N_16189);
nand U20007 (N_20007,N_16083,N_15546);
or U20008 (N_20008,N_16448,N_17202);
or U20009 (N_20009,N_15264,N_16958);
or U20010 (N_20010,N_15058,N_17809);
xor U20011 (N_20011,N_17175,N_15166);
and U20012 (N_20012,N_17242,N_17481);
or U20013 (N_20013,N_15277,N_18099);
or U20014 (N_20014,N_17174,N_15377);
xnor U20015 (N_20015,N_16068,N_16124);
or U20016 (N_20016,N_19611,N_17664);
or U20017 (N_20017,N_19086,N_19376);
and U20018 (N_20018,N_17182,N_19503);
and U20019 (N_20019,N_17070,N_19721);
nand U20020 (N_20020,N_19734,N_18248);
xnor U20021 (N_20021,N_18566,N_16560);
xor U20022 (N_20022,N_15821,N_18480);
nor U20023 (N_20023,N_16884,N_19638);
xnor U20024 (N_20024,N_16981,N_18330);
nand U20025 (N_20025,N_15543,N_19619);
nor U20026 (N_20026,N_18932,N_16322);
xor U20027 (N_20027,N_19766,N_16949);
nand U20028 (N_20028,N_19365,N_15693);
and U20029 (N_20029,N_17600,N_17616);
xor U20030 (N_20030,N_18325,N_18571);
or U20031 (N_20031,N_17763,N_19218);
xor U20032 (N_20032,N_15274,N_16330);
and U20033 (N_20033,N_15729,N_16233);
nor U20034 (N_20034,N_17048,N_17354);
or U20035 (N_20035,N_17312,N_16631);
nand U20036 (N_20036,N_15341,N_15353);
nand U20037 (N_20037,N_18395,N_19440);
or U20038 (N_20038,N_15698,N_16250);
and U20039 (N_20039,N_15326,N_18637);
or U20040 (N_20040,N_16253,N_18112);
or U20041 (N_20041,N_18491,N_16519);
xor U20042 (N_20042,N_15452,N_17759);
xor U20043 (N_20043,N_15763,N_18088);
xnor U20044 (N_20044,N_18920,N_17138);
xor U20045 (N_20045,N_15263,N_17478);
and U20046 (N_20046,N_15589,N_16353);
nor U20047 (N_20047,N_18155,N_16853);
or U20048 (N_20048,N_19396,N_18505);
and U20049 (N_20049,N_17404,N_15169);
xor U20050 (N_20050,N_15883,N_15554);
or U20051 (N_20051,N_19383,N_17698);
nand U20052 (N_20052,N_19778,N_15290);
or U20053 (N_20053,N_17011,N_18953);
xnor U20054 (N_20054,N_17090,N_17653);
xnor U20055 (N_20055,N_15598,N_19319);
and U20056 (N_20056,N_18403,N_18811);
xnor U20057 (N_20057,N_16643,N_18245);
and U20058 (N_20058,N_17876,N_18537);
or U20059 (N_20059,N_16416,N_19296);
or U20060 (N_20060,N_16137,N_17502);
nor U20061 (N_20061,N_17310,N_18456);
and U20062 (N_20062,N_18674,N_15932);
xor U20063 (N_20063,N_18848,N_18093);
xor U20064 (N_20064,N_17890,N_17435);
xnor U20065 (N_20065,N_16116,N_18853);
nor U20066 (N_20066,N_16864,N_16451);
nor U20067 (N_20067,N_17888,N_18520);
or U20068 (N_20068,N_18079,N_16428);
xor U20069 (N_20069,N_18760,N_18063);
nand U20070 (N_20070,N_16086,N_15715);
xnor U20071 (N_20071,N_19404,N_17430);
and U20072 (N_20072,N_15671,N_15023);
or U20073 (N_20073,N_16869,N_18377);
nor U20074 (N_20074,N_15603,N_16708);
or U20075 (N_20075,N_17540,N_16754);
and U20076 (N_20076,N_19502,N_18771);
xnor U20077 (N_20077,N_16815,N_15762);
nor U20078 (N_20078,N_19018,N_18924);
or U20079 (N_20079,N_18777,N_16932);
and U20080 (N_20080,N_15300,N_19189);
xnor U20081 (N_20081,N_17582,N_17299);
xor U20082 (N_20082,N_17285,N_17046);
nor U20083 (N_20083,N_15292,N_16044);
xor U20084 (N_20084,N_18247,N_15031);
xnor U20085 (N_20085,N_17902,N_16022);
and U20086 (N_20086,N_16952,N_16273);
xor U20087 (N_20087,N_16348,N_15876);
nand U20088 (N_20088,N_18043,N_18738);
nor U20089 (N_20089,N_19781,N_16766);
xnor U20090 (N_20090,N_15923,N_15520);
or U20091 (N_20091,N_17190,N_15634);
xor U20092 (N_20092,N_15740,N_16750);
nor U20093 (N_20093,N_15756,N_16435);
xnor U20094 (N_20094,N_19536,N_19884);
or U20095 (N_20095,N_18747,N_17020);
or U20096 (N_20096,N_17837,N_17055);
and U20097 (N_20097,N_15230,N_18751);
or U20098 (N_20098,N_15366,N_15015);
nor U20099 (N_20099,N_19273,N_17840);
nor U20100 (N_20100,N_17019,N_19799);
nand U20101 (N_20101,N_18225,N_19194);
or U20102 (N_20102,N_18148,N_15094);
xnor U20103 (N_20103,N_19163,N_16729);
nand U20104 (N_20104,N_16597,N_18399);
or U20105 (N_20105,N_16039,N_19268);
nand U20106 (N_20106,N_19643,N_15103);
nor U20107 (N_20107,N_15832,N_15065);
or U20108 (N_20108,N_15802,N_17007);
nor U20109 (N_20109,N_18487,N_19452);
xnor U20110 (N_20110,N_16531,N_16025);
xnor U20111 (N_20111,N_19171,N_16668);
and U20112 (N_20112,N_17379,N_18194);
or U20113 (N_20113,N_18312,N_17091);
nor U20114 (N_20114,N_15751,N_19022);
nand U20115 (N_20115,N_19629,N_19288);
nand U20116 (N_20116,N_19001,N_19354);
nor U20117 (N_20117,N_15610,N_19696);
nor U20118 (N_20118,N_19886,N_18867);
xnor U20119 (N_20119,N_19133,N_19762);
nand U20120 (N_20120,N_19264,N_18511);
xor U20121 (N_20121,N_19728,N_16179);
or U20122 (N_20122,N_15632,N_19314);
and U20123 (N_20123,N_16702,N_19172);
xor U20124 (N_20124,N_15018,N_18797);
nand U20125 (N_20125,N_18359,N_17668);
nor U20126 (N_20126,N_18367,N_17586);
xor U20127 (N_20127,N_17437,N_19716);
and U20128 (N_20128,N_17014,N_17128);
nor U20129 (N_20129,N_16413,N_17716);
and U20130 (N_20130,N_18052,N_17735);
nand U20131 (N_20131,N_18922,N_19689);
xor U20132 (N_20132,N_18936,N_18598);
nand U20133 (N_20133,N_19692,N_17306);
xor U20134 (N_20134,N_17415,N_15393);
nor U20135 (N_20135,N_18426,N_16183);
xor U20136 (N_20136,N_18128,N_19775);
or U20137 (N_20137,N_16899,N_19564);
or U20138 (N_20138,N_18364,N_19910);
and U20139 (N_20139,N_18529,N_17359);
or U20140 (N_20140,N_15078,N_18648);
nor U20141 (N_20141,N_17395,N_16064);
or U20142 (N_20142,N_15423,N_19802);
and U20143 (N_20143,N_16477,N_18933);
or U20144 (N_20144,N_19379,N_18031);
and U20145 (N_20145,N_18821,N_17205);
or U20146 (N_20146,N_16184,N_17804);
or U20147 (N_20147,N_18672,N_15303);
or U20148 (N_20148,N_18217,N_16020);
xor U20149 (N_20149,N_17580,N_16517);
nand U20150 (N_20150,N_18834,N_19213);
nand U20151 (N_20151,N_18739,N_18996);
nor U20152 (N_20152,N_16092,N_15146);
nor U20153 (N_20153,N_15800,N_16218);
nor U20154 (N_20154,N_19289,N_15443);
nor U20155 (N_20155,N_19677,N_18113);
or U20156 (N_20156,N_18501,N_18595);
nand U20157 (N_20157,N_17471,N_15448);
or U20158 (N_20158,N_16276,N_19008);
or U20159 (N_20159,N_15468,N_19615);
and U20160 (N_20160,N_17695,N_18370);
xnor U20161 (N_20161,N_18409,N_15316);
or U20162 (N_20162,N_17723,N_17749);
xnor U20163 (N_20163,N_18096,N_17513);
and U20164 (N_20164,N_15935,N_16028);
nand U20165 (N_20165,N_15337,N_17343);
nor U20166 (N_20166,N_16031,N_19670);
or U20167 (N_20167,N_19113,N_17271);
xor U20168 (N_20168,N_17758,N_15760);
and U20169 (N_20169,N_19399,N_16714);
nand U20170 (N_20170,N_18697,N_18471);
and U20171 (N_20171,N_16040,N_16512);
nor U20172 (N_20172,N_15831,N_18220);
and U20173 (N_20173,N_16673,N_16625);
or U20174 (N_20174,N_15330,N_18846);
xor U20175 (N_20175,N_15828,N_19057);
nand U20176 (N_20176,N_16538,N_18743);
or U20177 (N_20177,N_17040,N_19249);
nand U20178 (N_20178,N_17741,N_17703);
nor U20179 (N_20179,N_18274,N_17536);
or U20180 (N_20180,N_18348,N_18277);
and U20181 (N_20181,N_16169,N_15373);
or U20182 (N_20182,N_15385,N_15497);
nand U20183 (N_20183,N_16872,N_19836);
or U20184 (N_20184,N_17670,N_18551);
and U20185 (N_20185,N_17448,N_17053);
nand U20186 (N_20186,N_15363,N_17887);
xnor U20187 (N_20187,N_19998,N_15574);
nand U20188 (N_20188,N_16893,N_18067);
or U20189 (N_20189,N_17498,N_19408);
or U20190 (N_20190,N_19582,N_19477);
or U20191 (N_20191,N_19167,N_15289);
xor U20192 (N_20192,N_16989,N_18304);
and U20193 (N_20193,N_18926,N_15812);
nand U20194 (N_20194,N_18038,N_15674);
nand U20195 (N_20195,N_16835,N_18818);
or U20196 (N_20196,N_15985,N_16879);
nand U20197 (N_20197,N_17697,N_15327);
nor U20198 (N_20198,N_17144,N_18550);
nand U20199 (N_20199,N_16946,N_18822);
and U20200 (N_20200,N_19980,N_17596);
xnor U20201 (N_20201,N_16104,N_19370);
nand U20202 (N_20202,N_16687,N_16108);
xnor U20203 (N_20203,N_17232,N_18151);
xor U20204 (N_20204,N_15437,N_17491);
or U20205 (N_20205,N_19139,N_16171);
and U20206 (N_20206,N_15072,N_17026);
xnor U20207 (N_20207,N_19904,N_17511);
xnor U20208 (N_20208,N_17520,N_19655);
nor U20209 (N_20209,N_16763,N_17439);
nor U20210 (N_20210,N_19606,N_17146);
and U20211 (N_20211,N_19870,N_19843);
nand U20212 (N_20212,N_17259,N_19149);
or U20213 (N_20213,N_15323,N_16050);
nand U20214 (N_20214,N_16805,N_17489);
or U20215 (N_20215,N_19384,N_16466);
or U20216 (N_20216,N_15466,N_15051);
xnor U20217 (N_20217,N_18283,N_15946);
xnor U20218 (N_20218,N_15990,N_19495);
and U20219 (N_20219,N_19512,N_19410);
xor U20220 (N_20220,N_17677,N_16450);
nand U20221 (N_20221,N_17017,N_16377);
or U20222 (N_20222,N_15734,N_16870);
xor U20223 (N_20223,N_15608,N_16890);
nor U20224 (N_20224,N_17462,N_18955);
or U20225 (N_20225,N_18673,N_15162);
and U20226 (N_20226,N_15336,N_16595);
or U20227 (N_20227,N_18954,N_19530);
and U20228 (N_20228,N_19271,N_15255);
or U20229 (N_20229,N_16186,N_16299);
or U20230 (N_20230,N_18706,N_17279);
nand U20231 (N_20231,N_17975,N_16764);
nand U20232 (N_20232,N_18150,N_15392);
xor U20233 (N_20233,N_15583,N_17323);
xor U20234 (N_20234,N_16749,N_15676);
and U20235 (N_20235,N_17391,N_16412);
nor U20236 (N_20236,N_17376,N_15662);
and U20237 (N_20237,N_19517,N_17911);
or U20238 (N_20238,N_17100,N_17367);
and U20239 (N_20239,N_17204,N_18035);
xor U20240 (N_20240,N_17332,N_19484);
nor U20241 (N_20241,N_19053,N_18786);
xor U20242 (N_20242,N_15982,N_18346);
and U20243 (N_20243,N_18272,N_15248);
nand U20244 (N_20244,N_18689,N_17225);
xnor U20245 (N_20245,N_19509,N_16120);
and U20246 (N_20246,N_18732,N_17342);
nand U20247 (N_20247,N_18990,N_17823);
or U20248 (N_20248,N_15979,N_17244);
nand U20249 (N_20249,N_16420,N_18089);
nor U20250 (N_20250,N_15971,N_18513);
and U20251 (N_20251,N_18881,N_17521);
xor U20252 (N_20252,N_18361,N_15957);
nand U20253 (N_20253,N_17874,N_17029);
nor U20254 (N_20254,N_16289,N_19921);
nand U20255 (N_20255,N_17083,N_19780);
or U20256 (N_20256,N_16453,N_16368);
xnor U20257 (N_20257,N_17743,N_17865);
and U20258 (N_20258,N_19824,N_16204);
xnor U20259 (N_20259,N_15987,N_16166);
or U20260 (N_20260,N_16343,N_16030);
or U20261 (N_20261,N_15396,N_18948);
xnor U20262 (N_20262,N_16640,N_19659);
xnor U20263 (N_20263,N_19878,N_16839);
or U20264 (N_20264,N_19191,N_19343);
or U20265 (N_20265,N_15747,N_16681);
xnor U20266 (N_20266,N_17004,N_16284);
nand U20267 (N_20267,N_16755,N_19990);
or U20268 (N_20268,N_16215,N_17124);
and U20269 (N_20269,N_19604,N_17964);
and U20270 (N_20270,N_19393,N_17387);
nand U20271 (N_20271,N_15048,N_19345);
xnor U20272 (N_20272,N_17431,N_15688);
xor U20273 (N_20273,N_17099,N_15805);
xnor U20274 (N_20274,N_17917,N_17103);
nand U20275 (N_20275,N_18707,N_16619);
nand U20276 (N_20276,N_16536,N_16962);
xor U20277 (N_20277,N_17424,N_15759);
xnor U20278 (N_20278,N_17413,N_15252);
nand U20279 (N_20279,N_16012,N_17635);
nand U20280 (N_20280,N_17684,N_19797);
and U20281 (N_20281,N_17351,N_15722);
nor U20282 (N_20282,N_16878,N_17024);
nor U20283 (N_20283,N_19342,N_17127);
nand U20284 (N_20284,N_16280,N_19568);
nand U20285 (N_20285,N_18898,N_16144);
and U20286 (N_20286,N_16267,N_15680);
nor U20287 (N_20287,N_19885,N_15943);
or U20288 (N_20288,N_19202,N_16277);
xnor U20289 (N_20289,N_16142,N_16868);
nor U20290 (N_20290,N_17618,N_16198);
nand U20291 (N_20291,N_19767,N_16844);
xnor U20292 (N_20292,N_17729,N_16709);
and U20293 (N_20293,N_15198,N_19551);
nand U20294 (N_20294,N_16898,N_16222);
or U20295 (N_20295,N_16281,N_19784);
nand U20296 (N_20296,N_16846,N_19806);
or U20297 (N_20297,N_15884,N_18423);
xor U20298 (N_20298,N_18561,N_15530);
and U20299 (N_20299,N_19589,N_15477);
nor U20300 (N_20300,N_19763,N_18579);
nand U20301 (N_20301,N_15531,N_18839);
xnor U20302 (N_20302,N_18265,N_15942);
nor U20303 (N_20303,N_18616,N_19764);
or U20304 (N_20304,N_16762,N_17167);
xor U20305 (N_20305,N_16534,N_19438);
nor U20306 (N_20306,N_15324,N_16954);
nand U20307 (N_20307,N_18017,N_17012);
and U20308 (N_20308,N_15056,N_18087);
xor U20309 (N_20309,N_15552,N_19088);
xnor U20310 (N_20310,N_16133,N_16817);
and U20311 (N_20311,N_17968,N_17614);
and U20312 (N_20312,N_17518,N_18758);
nor U20313 (N_20313,N_15352,N_16596);
and U20314 (N_20314,N_16489,N_17549);
xnor U20315 (N_20315,N_18020,N_16360);
or U20316 (N_20316,N_18912,N_17571);
or U20317 (N_20317,N_17620,N_19673);
or U20318 (N_20318,N_19465,N_16779);
and U20319 (N_20319,N_15120,N_15081);
or U20320 (N_20320,N_18719,N_16747);
nor U20321 (N_20321,N_19363,N_18903);
xor U20322 (N_20322,N_19842,N_19476);
or U20323 (N_20323,N_18240,N_19160);
or U20324 (N_20324,N_18583,N_15781);
xnor U20325 (N_20325,N_19923,N_16618);
and U20326 (N_20326,N_19786,N_15716);
and U20327 (N_20327,N_17896,N_15718);
nor U20328 (N_20328,N_16892,N_16583);
nand U20329 (N_20329,N_16592,N_16337);
nand U20330 (N_20330,N_16228,N_19602);
or U20331 (N_20331,N_18547,N_19050);
xnor U20332 (N_20332,N_15210,N_17276);
nand U20333 (N_20333,N_17609,N_19588);
or U20334 (N_20334,N_17702,N_16014);
and U20335 (N_20335,N_18290,N_17639);
or U20336 (N_20336,N_19029,N_17534);
or U20337 (N_20337,N_17330,N_18145);
nor U20338 (N_20338,N_18273,N_17066);
nand U20339 (N_20339,N_17084,N_18022);
and U20340 (N_20340,N_16473,N_17957);
nand U20341 (N_20341,N_19546,N_18663);
nor U20342 (N_20342,N_18215,N_19795);
or U20343 (N_20343,N_15492,N_16243);
or U20344 (N_20344,N_15964,N_16589);
and U20345 (N_20345,N_17708,N_18257);
and U20346 (N_20346,N_15167,N_15232);
or U20347 (N_20347,N_16479,N_16076);
nand U20348 (N_20348,N_16069,N_18327);
and U20349 (N_20349,N_18252,N_18255);
nor U20350 (N_20350,N_16901,N_18901);
nand U20351 (N_20351,N_15461,N_18407);
nand U20352 (N_20352,N_19028,N_16793);
nor U20353 (N_20353,N_18917,N_15629);
and U20354 (N_20354,N_15890,N_17254);
or U20355 (N_20355,N_17188,N_18018);
nand U20356 (N_20356,N_17522,N_18195);
nor U20357 (N_20357,N_16045,N_16568);
or U20358 (N_20358,N_15064,N_15627);
nand U20359 (N_20359,N_15914,N_18941);
nor U20360 (N_20360,N_16692,N_15795);
nand U20361 (N_20361,N_19403,N_17104);
nor U20362 (N_20362,N_19196,N_15374);
or U20363 (N_20363,N_17470,N_17465);
nand U20364 (N_20364,N_16153,N_18517);
nor U20365 (N_20365,N_18587,N_16100);
nor U20366 (N_20366,N_16398,N_17531);
nor U20367 (N_20367,N_19958,N_19467);
nor U20368 (N_20368,N_19963,N_17234);
or U20369 (N_20369,N_18496,N_19510);
nand U20370 (N_20370,N_17422,N_19894);
nand U20371 (N_20371,N_16672,N_18165);
xor U20372 (N_20372,N_15311,N_18639);
and U20373 (N_20373,N_16552,N_16737);
nand U20374 (N_20374,N_16252,N_18559);
and U20375 (N_20375,N_19811,N_17933);
nor U20376 (N_20376,N_18082,N_17371);
nand U20377 (N_20377,N_15547,N_16049);
or U20378 (N_20378,N_18385,N_18457);
nor U20379 (N_20379,N_15476,N_16671);
or U20380 (N_20380,N_19906,N_15107);
nor U20381 (N_20381,N_18085,N_16140);
nand U20382 (N_20382,N_18642,N_15049);
nand U20383 (N_20383,N_15359,N_18769);
xor U20384 (N_20384,N_18657,N_18001);
xnor U20385 (N_20385,N_17514,N_17222);
or U20386 (N_20386,N_17171,N_15029);
nand U20387 (N_20387,N_17613,N_16738);
or U20388 (N_20388,N_15223,N_17409);
nor U20389 (N_20389,N_15165,N_18794);
or U20390 (N_20390,N_19428,N_15891);
and U20391 (N_20391,N_17984,N_18524);
or U20392 (N_20392,N_18804,N_19649);
or U20393 (N_20393,N_18815,N_17889);
nand U20394 (N_20394,N_18560,N_19859);
nor U20395 (N_20395,N_15463,N_19197);
or U20396 (N_20396,N_15727,N_16224);
xor U20397 (N_20397,N_16249,N_16862);
nor U20398 (N_20398,N_19826,N_15604);
or U20399 (N_20399,N_15398,N_18928);
or U20400 (N_20400,N_16888,N_19298);
xnor U20401 (N_20401,N_19175,N_15572);
or U20402 (N_20402,N_17878,N_17784);
nand U20403 (N_20403,N_19491,N_15758);
and U20404 (N_20404,N_19310,N_16543);
xnor U20405 (N_20405,N_18966,N_16383);
or U20406 (N_20406,N_17986,N_15007);
or U20407 (N_20407,N_17834,N_19475);
xnor U20408 (N_20408,N_18649,N_17480);
xor U20409 (N_20409,N_19093,N_19875);
or U20410 (N_20410,N_18959,N_19624);
and U20411 (N_20411,N_17594,N_17794);
xor U20412 (N_20412,N_15471,N_18937);
xnor U20413 (N_20413,N_15160,N_15282);
or U20414 (N_20414,N_17787,N_17721);
nand U20415 (N_20415,N_18836,N_15057);
and U20416 (N_20416,N_16130,N_16203);
nand U20417 (N_20417,N_15912,N_19812);
or U20418 (N_20418,N_15666,N_18305);
xnor U20419 (N_20419,N_18424,N_15069);
xor U20420 (N_20420,N_17606,N_16430);
nor U20421 (N_20421,N_16753,N_17251);
nand U20422 (N_20422,N_19572,N_18459);
nor U20423 (N_20423,N_15453,N_17864);
xnor U20424 (N_20424,N_17654,N_19256);
and U20425 (N_20425,N_15937,N_19660);
or U20426 (N_20426,N_15550,N_16988);
nor U20427 (N_20427,N_16361,N_17230);
or U20428 (N_20428,N_16079,N_18746);
and U20429 (N_20429,N_17111,N_18962);
or U20430 (N_20430,N_17647,N_18957);
or U20431 (N_20431,N_15692,N_15147);
xor U20432 (N_20432,N_18952,N_18332);
nor U20433 (N_20433,N_16355,N_19426);
nor U20434 (N_20434,N_15809,N_18329);
xnor U20435 (N_20435,N_17059,N_19173);
nand U20436 (N_20436,N_16999,N_18092);
xnor U20437 (N_20437,N_19941,N_17243);
nor U20438 (N_20438,N_19874,N_17325);
and U20439 (N_20439,N_16669,N_18814);
nor U20440 (N_20440,N_19773,N_16822);
xnor U20441 (N_20441,N_16721,N_16964);
nor U20442 (N_20442,N_19107,N_15947);
or U20443 (N_20443,N_17803,N_15062);
nor U20444 (N_20444,N_17765,N_18380);
and U20445 (N_20445,N_17235,N_17773);
nor U20446 (N_20446,N_19744,N_18864);
and U20447 (N_20447,N_15008,N_16567);
nor U20448 (N_20448,N_18466,N_18791);
nand U20449 (N_20449,N_19136,N_16930);
or U20450 (N_20450,N_15999,N_19844);
nand U20451 (N_20451,N_19158,N_17621);
nand U20452 (N_20452,N_15206,N_16471);
xnor U20453 (N_20453,N_17901,N_18632);
or U20454 (N_20454,N_16371,N_15174);
xor U20455 (N_20455,N_18726,N_19614);
nand U20456 (N_20456,N_19713,N_19879);
or U20457 (N_20457,N_19285,N_16953);
xnor U20458 (N_20458,N_19062,N_18103);
and U20459 (N_20459,N_16863,N_16160);
and U20460 (N_20460,N_16118,N_16929);
and U20461 (N_20461,N_18429,N_16802);
or U20462 (N_20462,N_19608,N_18282);
nand U20463 (N_20463,N_19776,N_15214);
xor U20464 (N_20464,N_19449,N_17996);
xnor U20465 (N_20465,N_18866,N_19258);
or U20466 (N_20466,N_18365,N_16035);
xor U20467 (N_20467,N_17566,N_15141);
and U20468 (N_20468,N_18737,N_19593);
xor U20469 (N_20469,N_17212,N_15288);
xor U20470 (N_20470,N_17372,N_16637);
nand U20471 (N_20471,N_16774,N_17515);
or U20472 (N_20472,N_15075,N_15012);
nand U20473 (N_20473,N_15409,N_16278);
xnor U20474 (N_20474,N_17678,N_19240);
or U20475 (N_20475,N_19684,N_17288);
xnor U20476 (N_20476,N_18203,N_15976);
or U20477 (N_20477,N_16182,N_17622);
and U20478 (N_20478,N_16696,N_17718);
and U20479 (N_20479,N_16515,N_17042);
nand U20480 (N_20480,N_15867,N_18609);
and U20481 (N_20481,N_17807,N_15266);
xnor U20482 (N_20482,N_15743,N_17361);
nand U20483 (N_20483,N_17704,N_15389);
or U20484 (N_20484,N_16176,N_18944);
xor U20485 (N_20485,N_18554,N_19900);
or U20486 (N_20486,N_17134,N_18764);
and U20487 (N_20487,N_19892,N_16043);
nand U20488 (N_20488,N_18897,N_17088);
and U20489 (N_20489,N_18373,N_16024);
nor U20490 (N_20490,N_19094,N_18582);
nand U20491 (N_20491,N_18993,N_17630);
or U20492 (N_20492,N_18268,N_17875);
or U20493 (N_20493,N_19199,N_15293);
nor U20494 (N_20494,N_15505,N_15527);
or U20495 (N_20495,N_18224,N_17688);
xnor U20496 (N_20496,N_15670,N_17727);
nor U20497 (N_20497,N_16758,N_19566);
and U20498 (N_20498,N_17368,N_17877);
or U20499 (N_20499,N_19430,N_18242);
or U20500 (N_20500,N_15306,N_18512);
nand U20501 (N_20501,N_17971,N_19722);
nand U20502 (N_20502,N_18398,N_15027);
nand U20503 (N_20503,N_19731,N_15365);
and U20504 (N_20504,N_16865,N_16942);
xnor U20505 (N_20505,N_15844,N_18885);
or U20506 (N_20506,N_15164,N_17049);
or U20507 (N_20507,N_18384,N_15155);
xor U20508 (N_20508,N_19397,N_19928);
nand U20509 (N_20509,N_17063,N_17044);
nor U20510 (N_20510,N_16480,N_19235);
nor U20511 (N_20511,N_17880,N_19697);
nand U20512 (N_20512,N_15667,N_15536);
or U20513 (N_20513,N_19981,N_16813);
xor U20514 (N_20514,N_19882,N_15772);
nor U20515 (N_20515,N_15845,N_17927);
nor U20516 (N_20516,N_16173,N_17812);
nand U20517 (N_20517,N_17665,N_15860);
or U20518 (N_20518,N_16296,N_19312);
xnor U20519 (N_20519,N_17912,N_17976);
nor U20520 (N_20520,N_18845,N_15577);
and U20521 (N_20521,N_18484,N_15564);
xor U20522 (N_20522,N_15349,N_15479);
nor U20523 (N_20523,N_19936,N_19849);
and U20524 (N_20524,N_17140,N_19031);
nand U20525 (N_20525,N_16496,N_15892);
xor U20526 (N_20526,N_16264,N_16190);
nor U20527 (N_20527,N_18942,N_17092);
nor U20528 (N_20528,N_17564,N_19006);
nor U20529 (N_20529,N_15467,N_17497);
xor U20530 (N_20530,N_18350,N_16410);
nand U20531 (N_20531,N_16492,N_16101);
xor U20532 (N_20532,N_17038,N_15247);
xor U20533 (N_20533,N_19803,N_16828);
or U20534 (N_20534,N_18392,N_16503);
nand U20535 (N_20535,N_15991,N_18289);
nand U20536 (N_20536,N_15254,N_16994);
or U20537 (N_20537,N_17130,N_17426);
and U20538 (N_20538,N_19535,N_15244);
xnor U20539 (N_20539,N_19048,N_18795);
xor U20540 (N_20540,N_18080,N_15291);
xnor U20541 (N_20541,N_19101,N_17320);
and U20542 (N_20542,N_19544,N_16251);
nand U20543 (N_20543,N_18324,N_15158);
nand U20544 (N_20544,N_19297,N_15132);
nand U20545 (N_20545,N_19307,N_15131);
xor U20546 (N_20546,N_16513,N_15825);
or U20547 (N_20547,N_19690,N_18024);
nor U20548 (N_20548,N_17484,N_18125);
and U20549 (N_20549,N_17855,N_19902);
and U20550 (N_20550,N_18023,N_16620);
and U20551 (N_20551,N_18231,N_18754);
and U20552 (N_20552,N_17151,N_19417);
and U20553 (N_20553,N_18431,N_16905);
or U20554 (N_20554,N_19742,N_15469);
nand U20555 (N_20555,N_16563,N_18950);
xor U20556 (N_20556,N_19035,N_15636);
xnor U20557 (N_20557,N_19400,N_17400);
xnor U20558 (N_20558,N_15019,N_17460);
nand U20559 (N_20559,N_18120,N_19445);
xnor U20560 (N_20560,N_17916,N_16293);
nor U20561 (N_20561,N_18345,N_15362);
xnor U20562 (N_20562,N_15977,N_18907);
and U20563 (N_20563,N_15807,N_17687);
nand U20564 (N_20564,N_19060,N_19047);
nand U20565 (N_20565,N_19529,N_19077);
or U20566 (N_20566,N_17005,N_19487);
xor U20567 (N_20567,N_15231,N_16551);
nor U20568 (N_20568,N_19729,N_18600);
nor U20569 (N_20569,N_19574,N_17858);
or U20570 (N_20570,N_19371,N_15719);
or U20571 (N_20571,N_16418,N_18721);
xor U20572 (N_20572,N_18351,N_17782);
xnor U20573 (N_20573,N_19225,N_16849);
nor U20574 (N_20574,N_18157,N_16759);
or U20575 (N_20575,N_15871,N_16365);
xnor U20576 (N_20576,N_17344,N_17095);
xor U20577 (N_20577,N_15405,N_18382);
nand U20578 (N_20578,N_16180,N_18455);
nor U20579 (N_20579,N_18275,N_17421);
nand U20580 (N_20580,N_16824,N_15310);
xor U20581 (N_20581,N_15243,N_19951);
and U20582 (N_20582,N_18177,N_19243);
and U20583 (N_20583,N_17378,N_16686);
nand U20584 (N_20584,N_15669,N_19041);
xor U20585 (N_20585,N_17560,N_18021);
xor U20586 (N_20586,N_19702,N_17457);
or U20587 (N_20587,N_17179,N_18141);
nand U20588 (N_20588,N_17977,N_15499);
and U20589 (N_20589,N_17475,N_19671);
xor U20590 (N_20590,N_19032,N_15642);
nor U20591 (N_20591,N_17573,N_18360);
nand U20592 (N_20592,N_16232,N_15768);
or U20593 (N_20593,N_17646,N_17990);
or U20594 (N_20594,N_18847,N_16831);
xnor U20595 (N_20595,N_18536,N_19575);
nand U20596 (N_20596,N_15881,N_15707);
nor U20597 (N_20597,N_17793,N_15744);
and U20598 (N_20598,N_19519,N_16990);
or U20599 (N_20599,N_17073,N_17045);
xnor U20600 (N_20600,N_18467,N_18874);
xor U20601 (N_20601,N_17852,N_16550);
nand U20602 (N_20602,N_18636,N_16210);
and U20603 (N_20603,N_16174,N_18546);
xor U20604 (N_20604,N_15983,N_18976);
nor U20605 (N_20605,N_18216,N_18658);
xor U20606 (N_20606,N_18333,N_17148);
and U20607 (N_20607,N_16579,N_16629);
nand U20608 (N_20608,N_18212,N_19771);
and U20609 (N_20609,N_18435,N_19768);
or U20610 (N_20610,N_18988,N_19034);
nand U20611 (N_20611,N_19110,N_15414);
nor U20612 (N_20612,N_16085,N_15897);
nor U20613 (N_20613,N_16810,N_15149);
nand U20614 (N_20614,N_16366,N_19953);
nand U20615 (N_20615,N_15542,N_16334);
nor U20616 (N_20616,N_15140,N_15411);
and U20617 (N_20617,N_17919,N_15833);
and U20618 (N_20618,N_19155,N_18383);
nand U20619 (N_20619,N_18149,N_15364);
nand U20620 (N_20620,N_18544,N_18712);
or U20621 (N_20621,N_15655,N_19454);
and U20622 (N_20622,N_15503,N_15921);
or U20623 (N_20623,N_17006,N_15089);
nand U20624 (N_20624,N_16297,N_16227);
and U20625 (N_20625,N_15489,N_17181);
nand U20626 (N_20626,N_15509,N_16483);
or U20627 (N_20627,N_15261,N_17969);
nor U20628 (N_20628,N_19108,N_16982);
or U20629 (N_20629,N_15071,N_19866);
xor U20630 (N_20630,N_15339,N_18410);
and U20631 (N_20631,N_16925,N_18521);
nor U20632 (N_20632,N_15368,N_19971);
xnor U20633 (N_20633,N_16260,N_19747);
or U20634 (N_20634,N_18340,N_17231);
or U20635 (N_20635,N_15319,N_19015);
or U20636 (N_20636,N_18347,N_16414);
xor U20637 (N_20637,N_16987,N_18577);
xnor U20638 (N_20638,N_16794,N_19633);
nor U20639 (N_20639,N_18756,N_19681);
nor U20640 (N_20640,N_18631,N_18136);
nor U20641 (N_20641,N_19738,N_19667);
or U20642 (N_20642,N_19385,N_16840);
xnor U20643 (N_20643,N_19694,N_17168);
and U20644 (N_20644,N_15568,N_16847);
or U20645 (N_20645,N_19709,N_18971);
and U20646 (N_20646,N_15705,N_19112);
or U20647 (N_20647,N_16419,N_17450);
nand U20648 (N_20648,N_15478,N_18807);
and U20649 (N_20649,N_15725,N_17681);
nor U20650 (N_20650,N_15115,N_19748);
nand U20651 (N_20651,N_16722,N_18730);
nor U20652 (N_20652,N_19903,N_19045);
xor U20653 (N_20653,N_19051,N_18066);
or U20654 (N_20654,N_18931,N_17335);
xor U20655 (N_20655,N_17319,N_17227);
nand U20656 (N_20656,N_19024,N_16301);
or U20657 (N_20657,N_18323,N_19291);
xor U20658 (N_20658,N_18253,N_16984);
or U20659 (N_20659,N_19931,N_15429);
xnor U20660 (N_20660,N_18184,N_17533);
and U20661 (N_20661,N_18530,N_16128);
and U20662 (N_20662,N_15464,N_19381);
and U20663 (N_20663,N_17322,N_19209);
and U20664 (N_20664,N_15639,N_19933);
and U20665 (N_20665,N_15189,N_19959);
or U20666 (N_20666,N_16388,N_18138);
nand U20667 (N_20667,N_18711,N_18121);
and U20668 (N_20668,N_15403,N_18902);
xor U20669 (N_20669,N_17016,N_16547);
nand U20670 (N_20670,N_16736,N_19373);
nor U20671 (N_20671,N_15548,N_16587);
and U20672 (N_20672,N_16175,N_19964);
nor U20673 (N_20673,N_15567,N_17429);
nor U20674 (N_20674,N_16812,N_18132);
nor U20675 (N_20675,N_17009,N_19909);
and U20676 (N_20676,N_18201,N_18027);
xnor U20677 (N_20677,N_15804,N_17187);
xor U20678 (N_20678,N_18202,N_15724);
nor U20679 (N_20679,N_19915,N_15450);
nor U20680 (N_20680,N_18129,N_17753);
xnor U20681 (N_20681,N_19206,N_17085);
nand U20682 (N_20682,N_16188,N_18303);
and U20683 (N_20683,N_18056,N_19068);
nand U20684 (N_20684,N_18989,N_16308);
xnor U20685 (N_20685,N_16098,N_17412);
xor U20686 (N_20686,N_19207,N_19676);
nor U20687 (N_20687,N_15672,N_15177);
nand U20688 (N_20688,N_16187,N_15868);
and U20689 (N_20689,N_17458,N_17924);
nor U20690 (N_20690,N_16380,N_15838);
and U20691 (N_20691,N_15824,N_19000);
nand U20692 (N_20692,N_17318,N_16823);
or U20693 (N_20693,N_16306,N_19505);
nand U20694 (N_20694,N_15088,N_19276);
xor U20695 (N_20695,N_15585,N_18523);
xor U20696 (N_20696,N_19995,N_19863);
nor U20697 (N_20697,N_15428,N_15501);
xor U20698 (N_20698,N_18655,N_19355);
xor U20699 (N_20699,N_16927,N_17443);
nor U20700 (N_20700,N_17693,N_16279);
or U20701 (N_20701,N_19358,N_15712);
nor U20702 (N_20702,N_19717,N_16422);
nor U20703 (N_20703,N_18285,N_16112);
xor U20704 (N_20704,N_16647,N_17768);
xor U20705 (N_20705,N_17137,N_16756);
nor U20706 (N_20706,N_17894,N_15026);
nor U20707 (N_20707,N_18570,N_19080);
nor U20708 (N_20708,N_16417,N_18854);
nor U20709 (N_20709,N_16682,N_19165);
nand U20710 (N_20710,N_17064,N_19064);
xnor U20711 (N_20711,N_15687,N_18379);
nand U20712 (N_20712,N_18033,N_15010);
and U20713 (N_20713,N_18016,N_16320);
and U20714 (N_20714,N_17283,N_19216);
xnor U20715 (N_20715,N_15789,N_16499);
and U20716 (N_20716,N_15434,N_19456);
nand U20717 (N_20717,N_19985,N_16246);
or U20718 (N_20718,N_16986,N_16465);
nor U20719 (N_20719,N_19751,N_15938);
or U20720 (N_20720,N_18307,N_17419);
nor U20721 (N_20721,N_15590,N_18588);
nand U20722 (N_20722,N_19313,N_15766);
xor U20723 (N_20723,N_19949,N_18679);
xor U20724 (N_20724,N_15276,N_18541);
nor U20725 (N_20725,N_17455,N_19912);
and U20726 (N_20726,N_19516,N_16339);
or U20727 (N_20727,N_17551,N_15931);
or U20728 (N_20728,N_16730,N_16569);
and U20729 (N_20729,N_15637,N_15765);
or U20730 (N_20730,N_19800,N_15318);
nor U20731 (N_20731,N_17791,N_18048);
xor U20732 (N_20732,N_19883,N_17802);
nand U20733 (N_20733,N_19628,N_18281);
or U20734 (N_20734,N_19665,N_15581);
and U20735 (N_20735,N_18805,N_19121);
xnor U20736 (N_20736,N_16167,N_16918);
xor U20737 (N_20737,N_16875,N_16216);
nor U20738 (N_20738,N_19309,N_16271);
nand U20739 (N_20739,N_16578,N_17463);
nor U20740 (N_20740,N_18614,N_17201);
nand U20741 (N_20741,N_18450,N_17304);
or U20742 (N_20742,N_16716,N_15313);
and U20743 (N_20743,N_15854,N_18538);
xor U20744 (N_20744,N_19796,N_16735);
or U20745 (N_20745,N_19241,N_17795);
or U20746 (N_20746,N_17701,N_18186);
and U20747 (N_20747,N_18870,N_15630);
and U20748 (N_20748,N_16765,N_18452);
and U20749 (N_20749,N_17944,N_15969);
or U20750 (N_20750,N_15055,N_18698);
or U20751 (N_20751,N_19020,N_18770);
or U20752 (N_20752,N_18790,N_19102);
nand U20753 (N_20753,N_16785,N_18784);
nor U20754 (N_20754,N_17028,N_17456);
xnor U20755 (N_20755,N_15895,N_19816);
xnor U20756 (N_20756,N_17001,N_19790);
nor U20757 (N_20757,N_17745,N_17923);
and U20758 (N_20758,N_15645,N_15347);
nand U20759 (N_20759,N_15170,N_17872);
nor U20760 (N_20760,N_15822,N_18652);
xnor U20761 (N_20761,N_15579,N_17256);
xnor U20762 (N_20762,N_17301,N_16516);
xor U20763 (N_20763,N_19553,N_17196);
and U20764 (N_20764,N_17278,N_18482);
and U20765 (N_20765,N_19550,N_17886);
nor U20766 (N_20766,N_18704,N_18401);
nor U20767 (N_20767,N_18199,N_18209);
nor U20768 (N_20768,N_17710,N_19919);
and U20769 (N_20769,N_16786,N_18972);
nor U20770 (N_20770,N_18724,N_17122);
nand U20771 (N_20771,N_16819,N_19346);
nand U20772 (N_20772,N_19613,N_16294);
xor U20773 (N_20773,N_15329,N_18635);
and U20774 (N_20774,N_19339,N_18694);
or U20775 (N_20775,N_16649,N_16979);
nor U20776 (N_20776,N_17185,N_18925);
or U20777 (N_20777,N_19735,N_16633);
nand U20778 (N_20778,N_16969,N_18140);
nor U20779 (N_20779,N_18562,N_18534);
nor U20780 (N_20780,N_18943,N_16664);
or U20781 (N_20781,N_15958,N_16950);
nor U20782 (N_20782,N_17810,N_19232);
and U20783 (N_20783,N_17814,N_18667);
and U20784 (N_20784,N_15661,N_19737);
or U20785 (N_20785,N_18008,N_15843);
nand U20786 (N_20786,N_15379,N_18827);
xnor U20787 (N_20787,N_16700,N_17373);
nand U20788 (N_20788,N_17528,N_15037);
xnor U20789 (N_20789,N_18154,N_16341);
and U20790 (N_20790,N_16303,N_16641);
xor U20791 (N_20791,N_18683,N_18439);
nor U20792 (N_20792,N_18660,N_18389);
or U20793 (N_20793,N_15638,N_18668);
nand U20794 (N_20794,N_17764,N_19164);
nand U20795 (N_20795,N_16523,N_16352);
xnor U20796 (N_20796,N_16185,N_18418);
nand U20797 (N_20797,N_18474,N_19617);
nor U20798 (N_20798,N_15001,N_19607);
and U20799 (N_20799,N_15721,N_18623);
or U20800 (N_20800,N_19814,N_17266);
nand U20801 (N_20801,N_18497,N_18842);
xnor U20802 (N_20802,N_15475,N_19049);
nor U20803 (N_20803,N_18427,N_17268);
nor U20804 (N_20804,N_17221,N_18865);
nor U20805 (N_20805,N_19187,N_19533);
and U20806 (N_20806,N_15893,N_15928);
or U20807 (N_20807,N_18180,N_18861);
xnor U20808 (N_20808,N_16914,N_18032);
xnor U20809 (N_20809,N_16207,N_16948);
and U20810 (N_20810,N_15128,N_16542);
and U20811 (N_20811,N_17317,N_18887);
xnor U20812 (N_20812,N_18072,N_18097);
nor U20813 (N_20813,N_17113,N_19727);
nor U20814 (N_20814,N_19987,N_18011);
nor U20815 (N_20815,N_15416,N_16789);
nor U20816 (N_20816,N_16093,N_19600);
or U20817 (N_20817,N_16559,N_19471);
or U20818 (N_20818,N_19097,N_19054);
xor U20819 (N_20819,N_15419,N_19782);
xnor U20820 (N_20820,N_16195,N_18299);
or U20821 (N_20821,N_15617,N_17525);
xor U20822 (N_20822,N_16887,N_19065);
and U20823 (N_20823,N_19950,N_16268);
and U20824 (N_20824,N_18083,N_15650);
xor U20825 (N_20825,N_18844,N_17047);
nand U20826 (N_20826,N_15267,N_19743);
or U20827 (N_20827,N_16406,N_17145);
and U20828 (N_20828,N_16162,N_19140);
or U20829 (N_20829,N_15124,N_19161);
nor U20830 (N_20830,N_17147,N_17107);
xnor U20831 (N_20831,N_17568,N_18593);
or U20832 (N_20832,N_19730,N_19578);
xor U20833 (N_20833,N_19236,N_19897);
nand U20834 (N_20834,N_19375,N_15228);
and U20835 (N_20835,N_18802,N_15053);
or U20836 (N_20836,N_18986,N_18510);
and U20837 (N_20837,N_19195,N_17574);
nand U20838 (N_20838,N_17022,N_17989);
and U20839 (N_20839,N_18034,N_16060);
nand U20840 (N_20840,N_16070,N_18028);
nor U20841 (N_20841,N_15656,N_19351);
xnor U20842 (N_20842,N_17381,N_17652);
and U20843 (N_20843,N_19052,N_16013);
xor U20844 (N_20844,N_19401,N_18946);
xnor U20845 (N_20845,N_17483,N_17605);
or U20846 (N_20846,N_19168,N_19605);
xor U20847 (N_20847,N_16056,N_18581);
nand U20848 (N_20848,N_18101,N_18046);
xor U20849 (N_20849,N_19994,N_18979);
nand U20850 (N_20850,N_18223,N_18708);
nor U20851 (N_20851,N_15205,N_16775);
nand U20852 (N_20852,N_15767,N_15493);
nor U20853 (N_20853,N_15872,N_15866);
xor U20854 (N_20854,N_17248,N_18569);
nor U20855 (N_20855,N_18575,N_16710);
nand U20856 (N_20856,N_16421,N_15328);
xor U20857 (N_20857,N_19466,N_17255);
xnor U20858 (N_20858,N_16606,N_19637);
xnor U20859 (N_20859,N_19215,N_15559);
nand U20860 (N_20860,N_17565,N_18750);
and U20861 (N_20861,N_16245,N_16208);
or U20862 (N_20862,N_17993,N_17966);
and U20863 (N_20863,N_19328,N_18376);
xnor U20864 (N_20864,N_17500,N_15101);
and U20865 (N_20865,N_15644,N_18042);
and U20866 (N_20866,N_19525,N_19040);
nand U20867 (N_20867,N_16469,N_17643);
nand U20868 (N_20868,N_19156,N_15899);
nor U20869 (N_20869,N_15494,N_15067);
xnor U20870 (N_20870,N_15780,N_15848);
or U20871 (N_20871,N_19657,N_15445);
xor U20872 (N_20872,N_15668,N_18896);
and U20873 (N_20873,N_16292,N_16707);
and U20874 (N_20874,N_19152,N_19965);
or U20875 (N_20875,N_17003,N_18331);
or U20876 (N_20876,N_16129,N_18628);
and U20877 (N_20877,N_16842,N_16727);
and U20878 (N_20878,N_18135,N_19873);
or U20879 (N_20879,N_15151,N_16158);
or U20880 (N_20880,N_17673,N_15221);
xor U20881 (N_20881,N_15387,N_19669);
nor U20882 (N_20882,N_18156,N_17291);
nand U20883 (N_20883,N_19740,N_15686);
nand U20884 (N_20884,N_19753,N_18167);
xor U20885 (N_20885,N_18328,N_18515);
and U20886 (N_20886,N_18051,N_17080);
nor U20887 (N_20887,N_15272,N_17870);
nand U20888 (N_20888,N_19090,N_17177);
and U20889 (N_20889,N_15989,N_15126);
nor U20890 (N_20890,N_15506,N_18076);
xor U20891 (N_20891,N_19966,N_15195);
or U20892 (N_20892,N_17416,N_15704);
xnor U20893 (N_20893,N_18929,N_15591);
xor U20894 (N_20894,N_15761,N_16533);
and U20895 (N_20895,N_15507,N_16392);
or U20896 (N_20896,N_19185,N_16234);
nor U20897 (N_20897,N_19126,N_19061);
nor U20898 (N_20898,N_19398,N_17656);
nand U20899 (N_20899,N_17868,N_17767);
nor U20900 (N_20900,N_15521,N_15102);
or U20901 (N_20901,N_17495,N_16199);
xnor U20902 (N_20902,N_18514,N_17780);
or U20903 (N_20903,N_16405,N_16141);
nand U20904 (N_20904,N_17298,N_16123);
nor U20905 (N_20905,N_15532,N_19943);
xnor U20906 (N_20906,N_16393,N_18182);
and U20907 (N_20907,N_17240,N_17619);
nor U20908 (N_20908,N_18213,N_19992);
nand U20909 (N_20909,N_16478,N_17761);
nor U20910 (N_20910,N_17736,N_17757);
nor U20911 (N_20911,N_17504,N_19182);
and U20912 (N_20912,N_18464,N_19070);
xnor U20913 (N_20913,N_16581,N_19815);
nand U20914 (N_20914,N_16363,N_19058);
or U20915 (N_20915,N_18873,N_17863);
or U20916 (N_20916,N_17707,N_19148);
nand U20917 (N_20917,N_16440,N_19674);
xor U20918 (N_20918,N_19967,N_18984);
nor U20919 (N_20919,N_19829,N_17593);
nand U20920 (N_20920,N_19099,N_18237);
and U20921 (N_20921,N_18869,N_16720);
or U20922 (N_20922,N_17258,N_18301);
and U20923 (N_20923,N_18065,N_16781);
nor U20924 (N_20924,N_15857,N_15541);
or U20925 (N_20925,N_17474,N_17294);
xor U20926 (N_20926,N_17210,N_16541);
nand U20927 (N_20927,N_19792,N_16010);
xnor U20928 (N_20928,N_19798,N_15746);
and U20929 (N_20929,N_17341,N_16571);
nor U20930 (N_20930,N_18686,N_17072);
nor U20931 (N_20931,N_15184,N_15888);
or U20932 (N_20932,N_17472,N_16980);
nand U20933 (N_20933,N_17199,N_18838);
and U20934 (N_20934,N_15114,N_17034);
nand U20935 (N_20935,N_19229,N_17089);
nand U20936 (N_20936,N_19434,N_19573);
and U20937 (N_20937,N_19267,N_19183);
nand U20938 (N_20938,N_16963,N_19890);
or U20939 (N_20939,N_16827,N_16411);
and U20940 (N_20940,N_17948,N_17496);
or U20941 (N_20941,N_19079,N_17592);
xnor U20942 (N_20942,N_18783,N_18664);
and U20943 (N_20943,N_15413,N_19359);
and U20944 (N_20944,N_19277,N_15817);
nor U20945 (N_20945,N_15915,N_16327);
xnor U20946 (N_20946,N_17928,N_19260);
xnor U20947 (N_20947,N_19076,N_19071);
or U20948 (N_20948,N_17746,N_15551);
and U20949 (N_20949,N_19407,N_15204);
nor U20950 (N_20950,N_16603,N_19957);
and U20951 (N_20951,N_15441,N_16937);
nand U20952 (N_20952,N_15218,N_19823);
or U20953 (N_20953,N_18094,N_15565);
and U20954 (N_20954,N_15901,N_15190);
and U20955 (N_20955,N_17337,N_15209);
or U20956 (N_20956,N_18852,N_18723);
or U20957 (N_20957,N_18539,N_17224);
nand U20958 (N_20958,N_15827,N_18127);
nor U20959 (N_20959,N_17657,N_18995);
and U20960 (N_20960,N_18644,N_15305);
nor U20961 (N_20961,N_19711,N_17954);
nand U20962 (N_20962,N_16432,N_17074);
xor U20963 (N_20963,N_16018,N_16367);
xnor U20964 (N_20964,N_19693,N_17557);
or U20965 (N_20965,N_18883,N_17396);
xnor U20966 (N_20966,N_19201,N_16066);
nor U20967 (N_20967,N_19115,N_19046);
nor U20968 (N_20968,N_18286,N_18041);
and U20969 (N_20969,N_18214,N_15998);
or U20970 (N_20970,N_16238,N_16090);
nor U20971 (N_20971,N_17690,N_19646);
nor U20972 (N_20972,N_15731,N_17191);
or U20973 (N_20973,N_16359,N_18287);
nor U20974 (N_20974,N_16401,N_17032);
xnor U20975 (N_20975,N_16266,N_17336);
nor U20976 (N_20976,N_19493,N_19618);
nor U20977 (N_20977,N_15145,N_19389);
xnor U20978 (N_20978,N_15834,N_16726);
or U20979 (N_20979,N_19712,N_15343);
and U20980 (N_20980,N_19636,N_15348);
and U20981 (N_20981,N_16938,N_15249);
nor U20982 (N_20982,N_15540,N_19119);
and U20983 (N_20983,N_15333,N_18447);
nand U20984 (N_20984,N_16706,N_18412);
xor U20985 (N_20985,N_15250,N_18126);
nand U20986 (N_20986,N_16705,N_17842);
nand U20987 (N_20987,N_19733,N_15451);
and U20988 (N_20988,N_19233,N_16788);
or U20989 (N_20989,N_15122,N_17428);
and U20990 (N_20990,N_19431,N_18576);
nor U20991 (N_20991,N_19482,N_19968);
nand U20992 (N_20992,N_16497,N_19914);
and U20993 (N_20993,N_17420,N_17153);
and U20994 (N_20994,N_18573,N_19378);
nand U20995 (N_20995,N_15325,N_17799);
xor U20996 (N_20996,N_18119,N_18479);
and U20997 (N_20997,N_18173,N_19706);
or U20998 (N_20998,N_18516,N_16509);
or U20999 (N_20999,N_18279,N_16915);
or U21000 (N_21000,N_15404,N_19680);
and U21001 (N_21001,N_17056,N_16325);
nor U21002 (N_21002,N_15059,N_17731);
xor U21003 (N_21003,N_15997,N_19736);
nor U21004 (N_21004,N_19418,N_15601);
xor U21005 (N_21005,N_18624,N_15516);
nand U21006 (N_21006,N_19009,N_18705);
xnor U21007 (N_21007,N_17300,N_19299);
xor U21008 (N_21008,N_18991,N_19324);
and U21009 (N_21009,N_18826,N_18454);
nor U21010 (N_21010,N_16632,N_15090);
nand U21011 (N_21011,N_15003,N_16580);
xor U21012 (N_21012,N_15307,N_18205);
nand U21013 (N_21013,N_16230,N_18422);
and U21014 (N_21014,N_17662,N_16441);
or U21015 (N_21015,N_16313,N_16147);
nand U21016 (N_21016,N_16902,N_17030);
and U21017 (N_21017,N_18690,N_18780);
nor U21018 (N_21018,N_15320,N_17108);
nor U21019 (N_21019,N_16382,N_18735);
nor U21020 (N_21020,N_16399,N_15402);
and U21021 (N_21021,N_17824,N_19612);
and U21022 (N_21022,N_18297,N_19262);
nor U21023 (N_21023,N_16959,N_18860);
nor U21024 (N_21024,N_15953,N_17732);
xor U21025 (N_21025,N_18564,N_16248);
or U21026 (N_21026,N_15433,N_16826);
nor U21027 (N_21027,N_19871,N_16391);
nand U21028 (N_21028,N_15211,N_19069);
or U21029 (N_21029,N_19745,N_16777);
xnor U21030 (N_21030,N_18956,N_18146);
nor U21031 (N_21031,N_15125,N_15677);
nand U21032 (N_21032,N_17831,N_17938);
or U21033 (N_21033,N_19565,N_15797);
nand U21034 (N_21034,N_16518,N_19012);
xnor U21035 (N_21035,N_19424,N_19538);
xnor U21036 (N_21036,N_15042,N_15424);
xor U21037 (N_21037,N_17241,N_16659);
xnor U21038 (N_21038,N_15280,N_17081);
nor U21039 (N_21039,N_19754,N_17778);
or U21040 (N_21040,N_16454,N_16825);
nor U21041 (N_21041,N_15224,N_16787);
or U21042 (N_21042,N_15726,N_17157);
nor U21043 (N_21043,N_16798,N_16321);
nand U21044 (N_21044,N_19783,N_19146);
and U21045 (N_21045,N_16057,N_19360);
nand U21046 (N_21046,N_18900,N_17037);
nor U21047 (N_21047,N_16078,N_17854);
nor U21048 (N_21048,N_16146,N_18077);
nor U21049 (N_21049,N_15959,N_19461);
or U21050 (N_21050,N_15382,N_18913);
nor U21051 (N_21051,N_19837,N_19290);
nand U21052 (N_21052,N_19714,N_15454);
and U21053 (N_21053,N_18356,N_19221);
nor U21054 (N_21054,N_15217,N_15654);
or U21055 (N_21055,N_18292,N_16290);
xnor U21056 (N_21056,N_16939,N_19392);
nand U21057 (N_21057,N_16042,N_15755);
nand U21058 (N_21058,N_18879,N_18084);
xor U21059 (N_21059,N_15076,N_19898);
nand U21060 (N_21060,N_19227,N_16694);
or U21061 (N_21061,N_15044,N_17714);
or U21062 (N_21062,N_19228,N_15874);
or U21063 (N_21063,N_18493,N_19939);
xnor U21064 (N_21064,N_15033,N_17633);
nor U21065 (N_21065,N_19004,N_18819);
nor U21066 (N_21066,N_16850,N_17329);
and U21067 (N_21067,N_19922,N_17226);
or U21068 (N_21068,N_17811,N_16549);
and U21069 (N_21069,N_19340,N_17105);
nand U21070 (N_21070,N_19656,N_16265);
xor U21071 (N_21071,N_17334,N_15080);
or U21072 (N_21072,N_19416,N_17451);
or U21073 (N_21073,N_17583,N_19969);
xor U21074 (N_21074,N_15576,N_16645);
and U21075 (N_21075,N_17357,N_19622);
xnor U21076 (N_21076,N_18638,N_18967);
or U21077 (N_21077,N_17305,N_19142);
or U21078 (N_21078,N_16691,N_17467);
xor U21079 (N_21079,N_18293,N_15215);
nor U21080 (N_21080,N_15182,N_18181);
nor U21081 (N_21081,N_17349,N_19494);
and U21082 (N_21082,N_17493,N_19255);
xnor U21083 (N_21083,N_17383,N_18613);
or U21084 (N_21084,N_15519,N_18599);
nor U21085 (N_21085,N_17682,N_15593);
nand U21086 (N_21086,N_15257,N_19526);
xor U21087 (N_21087,N_17951,N_15995);
nand U21088 (N_21088,N_16718,N_19306);
nor U21089 (N_21089,N_16970,N_17820);
and U21090 (N_21090,N_19770,N_16704);
nor U21091 (N_21091,N_15152,N_15039);
or U21092 (N_21092,N_19926,N_16688);
nor U21093 (N_21093,N_17667,N_19122);
xnor U21094 (N_21094,N_18729,N_17943);
and U21095 (N_21095,N_16138,N_19929);
or U21096 (N_21096,N_16032,N_19834);
and U21097 (N_21097,N_19700,N_18665);
or U21098 (N_21098,N_17796,N_16095);
and U21099 (N_21099,N_18375,N_19924);
nand U21100 (N_21100,N_15907,N_18271);
nand U21101 (N_21101,N_16433,N_17442);
xor U21102 (N_21102,N_17607,N_18381);
or U21103 (N_21103,N_19833,N_19537);
or U21104 (N_21104,N_16426,N_15186);
xor U21105 (N_21105,N_16007,N_17973);
nor U21106 (N_21106,N_17097,N_18700);
and U21107 (N_21107,N_18574,N_19860);
or U21108 (N_21108,N_17015,N_15605);
xnor U21109 (N_21109,N_18317,N_16110);
nor U21110 (N_21110,N_19986,N_19096);
nor U21111 (N_21111,N_17280,N_17331);
or U21112 (N_21112,N_19804,N_18851);
or U21113 (N_21113,N_15104,N_18404);
nand U21114 (N_21114,N_17436,N_19237);
nand U21115 (N_21115,N_15878,N_17010);
nand U21116 (N_21116,N_16936,N_16712);
nor U21117 (N_21117,N_17906,N_19425);
or U21118 (N_21118,N_18444,N_16125);
nand U21119 (N_21119,N_18400,N_17669);
nor U21120 (N_21120,N_15367,N_17546);
xor U21121 (N_21121,N_16973,N_18781);
xor U21122 (N_21122,N_19303,N_15621);
and U21123 (N_21123,N_17098,N_19380);
or U21124 (N_21124,N_17838,N_15787);
xor U21125 (N_21125,N_18107,N_18608);
xnor U21126 (N_21126,N_18081,N_17591);
nor U21127 (N_21127,N_16594,N_15614);
xnor U21128 (N_21128,N_17469,N_19682);
or U21129 (N_21129,N_16883,N_17587);
nor U21130 (N_21130,N_18163,N_18720);
nand U21131 (N_21131,N_16396,N_19506);
and U21132 (N_21132,N_17720,N_18886);
or U21133 (N_21133,N_16576,N_15030);
or U21134 (N_21134,N_18374,N_19543);
nand U21135 (N_21135,N_15047,N_19409);
nand U21136 (N_21136,N_17236,N_16782);
or U21137 (N_21137,N_19948,N_17355);
nor U21138 (N_21138,N_18899,N_17101);
and U21139 (N_21139,N_18262,N_17338);
or U21140 (N_21140,N_18263,N_16242);
or U21141 (N_21141,N_17661,N_15262);
and U21142 (N_21142,N_15354,N_15684);
nor U21143 (N_21143,N_15561,N_19350);
nand U21144 (N_21144,N_16455,N_17267);
and U21145 (N_21145,N_15776,N_17295);
and U21146 (N_21146,N_19542,N_15006);
nor U21147 (N_21147,N_15517,N_18086);
xnor U21148 (N_21148,N_18905,N_15369);
xnor U21149 (N_21149,N_18968,N_15199);
nand U21150 (N_21150,N_18468,N_19248);
and U21151 (N_21151,N_18158,N_17577);
nor U21152 (N_21152,N_19501,N_17023);
nand U21153 (N_21153,N_16833,N_18390);
xor U21154 (N_21154,N_17043,N_15435);
nand U21155 (N_21155,N_17548,N_18820);
or U21156 (N_21156,N_16285,N_16261);
nor U21157 (N_21157,N_18558,N_19441);
xor U21158 (N_21158,N_19308,N_17393);
xnor U21159 (N_21159,N_17425,N_19756);
xnor U21160 (N_21160,N_15229,N_17447);
or U21161 (N_21161,N_15082,N_16554);
and U21162 (N_21162,N_16394,N_18923);
nor U21163 (N_21163,N_16263,N_19124);
and U21164 (N_21164,N_19868,N_16350);
xor U21165 (N_21165,N_19341,N_19078);
nand U21166 (N_21166,N_19809,N_15588);
and U21167 (N_21167,N_18945,N_19979);
xor U21168 (N_21168,N_16239,N_15779);
xor U21169 (N_21169,N_18229,N_15287);
nor U21170 (N_21170,N_16305,N_18441);
and U21171 (N_21171,N_18185,N_16094);
nor U21172 (N_21172,N_17296,N_16860);
nand U21173 (N_21173,N_15819,N_18193);
or U21174 (N_21174,N_19287,N_17615);
nand U21175 (N_21175,N_19422,N_15077);
and U21176 (N_21176,N_18872,N_18787);
nand U21177 (N_21177,N_16660,N_19016);
nand U21178 (N_21178,N_19545,N_18591);
nand U21179 (N_21179,N_15980,N_18030);
or U21180 (N_21180,N_15421,N_15618);
nor U21181 (N_21181,N_15296,N_17789);
nand U21182 (N_21182,N_16269,N_15764);
nor U21183 (N_21183,N_18518,N_15529);
and U21184 (N_21184,N_16231,N_16924);
and U21185 (N_21185,N_16934,N_15474);
nand U21186 (N_21186,N_18578,N_18070);
or U21187 (N_21187,N_16636,N_18300);
nor U21188 (N_21188,N_17830,N_19527);
nand U21189 (N_21189,N_16971,N_17816);
and U21190 (N_21190,N_19222,N_15380);
nand U21191 (N_21191,N_17189,N_15741);
nor U21192 (N_21192,N_19881,N_19023);
and U21193 (N_21193,N_16558,N_19305);
xor U21194 (N_21194,N_16745,N_15646);
or U21195 (N_21195,N_18799,N_19496);
xnor U21196 (N_21196,N_19474,N_15401);
nor U21197 (N_21197,N_18997,N_18894);
or U21198 (N_21198,N_18829,N_15034);
or U21199 (N_21199,N_15150,N_19917);
nor U21200 (N_21200,N_19204,N_19479);
nand U21201 (N_21201,N_17907,N_16588);
and U21202 (N_21202,N_16181,N_19066);
or U21203 (N_21203,N_15814,N_17775);
nand U21204 (N_21204,N_17308,N_18437);
xnor U21205 (N_21205,N_15933,N_17569);
or U21206 (N_21206,N_18054,N_18159);
or U21207 (N_21207,N_16820,N_15622);
or U21208 (N_21208,N_15188,N_15111);
nor U21209 (N_21209,N_19153,N_17114);
nor U21210 (N_21210,N_19552,N_16213);
and U21211 (N_21211,N_15163,N_19203);
nor U21212 (N_21212,N_18047,N_19180);
nand U21213 (N_21213,N_16859,N_17211);
nand U21214 (N_21214,N_15022,N_15631);
nor U21215 (N_21215,N_15653,N_19338);
xnor U21216 (N_21216,N_17992,N_16221);
xor U21217 (N_21217,N_17109,N_16799);
nor U21218 (N_21218,N_18095,N_16006);
nor U21219 (N_21219,N_15242,N_19323);
and U21220 (N_21220,N_19570,N_16425);
or U21221 (N_21221,N_19451,N_16241);
nor U21222 (N_21222,N_17509,N_15967);
nor U21223 (N_21223,N_16535,N_17261);
and U21224 (N_21224,N_15426,N_15728);
and U21225 (N_21225,N_16540,N_15384);
or U21226 (N_21226,N_17939,N_19030);
nor U21227 (N_21227,N_17905,N_18006);
nand U21228 (N_21228,N_16041,N_19623);
and U21229 (N_21229,N_17558,N_15175);
nand U21230 (N_21230,N_19485,N_15085);
or U21231 (N_21231,N_16757,N_15253);
and U21232 (N_21232,N_18434,N_15268);
or U21233 (N_21233,N_17120,N_15988);
nand U21234 (N_21234,N_17488,N_19143);
or U21235 (N_21235,N_19301,N_15818);
and U21236 (N_21236,N_17170,N_19292);
nor U21237 (N_21237,N_17847,N_18227);
nand U21238 (N_21238,N_18408,N_15701);
xnor U21239 (N_21239,N_19361,N_18837);
xnor U21240 (N_21240,N_15508,N_18676);
xor U21241 (N_21241,N_19200,N_19205);
or U21242 (N_21242,N_18162,N_17754);
nand U21243 (N_21243,N_16062,N_16644);
and U21244 (N_21244,N_15240,N_19579);
nand U21245 (N_21245,N_17149,N_15970);
nand U21246 (N_21246,N_17974,N_19231);
nand U21247 (N_21247,N_19190,N_15087);
xor U21248 (N_21248,N_16135,N_17062);
xor U21249 (N_21249,N_15607,N_18934);
nand U21250 (N_21250,N_19432,N_18440);
nor U21251 (N_21251,N_19584,N_15301);
nand U21252 (N_21252,N_18741,N_15898);
nor U21253 (N_21253,N_15440,N_19198);
and U21254 (N_21254,N_18321,N_15383);
and U21255 (N_21255,N_18508,N_16502);
or U21256 (N_21256,N_19524,N_17479);
and U21257 (N_21257,N_18659,N_15139);
xnor U21258 (N_21258,N_17186,N_15714);
nor U21259 (N_21259,N_15690,N_15484);
or U21260 (N_21260,N_19920,N_16575);
nand U21261 (N_21261,N_18472,N_19857);
nand U21262 (N_21262,N_17284,N_17156);
nand U21263 (N_21263,N_16544,N_18363);
and U21264 (N_21264,N_15361,N_19571);
nand U21265 (N_21265,N_15447,N_17277);
nand U21266 (N_21266,N_19368,N_18254);
and U21267 (N_21267,N_18010,N_16780);
xnor U21268 (N_21268,N_18104,N_19514);
nand U21269 (N_21269,N_15108,N_15786);
or U21270 (N_21270,N_15308,N_15865);
and U21271 (N_21271,N_19013,N_18572);
nand U21272 (N_21272,N_19678,N_16074);
xor U21273 (N_21273,N_16058,N_18563);
and U21274 (N_21274,N_16599,N_17711);
nand U21275 (N_21275,N_16498,N_17542);
nor U21276 (N_21276,N_19014,N_15098);
nor U21277 (N_21277,N_17747,N_18486);
and U21278 (N_21278,N_16956,N_17247);
or U21279 (N_21279,N_17193,N_16600);
or U21280 (N_21280,N_18091,N_17808);
nor U21281 (N_21281,N_16837,N_18335);
or U21282 (N_21282,N_18590,N_18406);
nand U21283 (N_21283,N_17313,N_19521);
and U21284 (N_21284,N_18651,N_19651);
and U21285 (N_21285,N_15395,N_16818);
nand U21286 (N_21286,N_16452,N_16105);
nor U21287 (N_21287,N_18442,N_18102);
nor U21288 (N_21288,N_17102,N_15945);
and U21289 (N_21289,N_19675,N_15201);
and U21290 (N_21290,N_16476,N_17215);
nor U21291 (N_21291,N_17464,N_15882);
nor U21292 (N_21292,N_15091,N_16690);
or U21293 (N_21293,N_16667,N_18528);
nor U21294 (N_21294,N_15432,N_17184);
nor U21295 (N_21295,N_19642,N_17885);
nand U21296 (N_21296,N_17402,N_17829);
xor U21297 (N_21297,N_15302,N_18565);
or U21298 (N_21298,N_19726,N_15420);
or U21299 (N_21299,N_15279,N_16314);
or U21300 (N_21300,N_19757,N_16896);
and U21301 (N_21301,N_15925,N_17817);
and U21302 (N_21302,N_17166,N_16287);
and U21303 (N_21303,N_15697,N_19867);
nor U21304 (N_21304,N_15372,N_19794);
nand U21305 (N_21305,N_16626,N_17648);
nand U21306 (N_21306,N_16627,N_18414);
nor U21307 (N_21307,N_18280,N_19534);
or U21308 (N_21308,N_15703,N_17867);
and U21309 (N_21309,N_18421,N_16487);
or U21310 (N_21310,N_19443,N_16566);
nor U21311 (N_21311,N_15137,N_18250);
or U21312 (N_21312,N_15939,N_18734);
and U21313 (N_21313,N_19037,N_16298);
nand U21314 (N_21314,N_19658,N_17203);
and U21315 (N_21315,N_16201,N_19405);
and U21316 (N_21316,N_17069,N_19429);
and U21317 (N_21317,N_15399,N_19188);
nand U21318 (N_21318,N_15920,N_18825);
or U21319 (N_21319,N_15500,N_17453);
xnor U21320 (N_21320,N_16219,N_17686);
xnor U21321 (N_21321,N_15371,N_17501);
xnor U21322 (N_21322,N_15013,N_19081);
nor U21323 (N_21323,N_16624,N_15465);
and U21324 (N_21324,N_15949,N_17559);
nand U21325 (N_21325,N_17370,N_17908);
nand U21326 (N_21326,N_15841,N_15573);
nor U21327 (N_21327,N_17742,N_17399);
and U21328 (N_21328,N_19984,N_17123);
nor U21329 (N_21329,N_18677,N_19852);
xnor U21330 (N_21330,N_16495,N_19072);
xor U21331 (N_21331,N_17627,N_15934);
or U21332 (N_21332,N_17575,N_16177);
or U21333 (N_21333,N_15283,N_15153);
or U21334 (N_21334,N_18369,N_17292);
nand U21335 (N_21335,N_18235,N_17126);
nor U21336 (N_21336,N_15643,N_18696);
and U21337 (N_21337,N_18413,N_16119);
xnor U21338 (N_21338,N_19846,N_16310);
and U21339 (N_21339,N_17289,N_18291);
or U21340 (N_21340,N_15275,N_18004);
xnor U21341 (N_21341,N_17485,N_19286);
or U21342 (N_21342,N_16164,N_19253);
or U21343 (N_21343,N_19162,N_18981);
nand U21344 (N_21344,N_16944,N_16689);
nor U21345 (N_21345,N_18005,N_16375);
xor U21346 (N_21346,N_19293,N_16680);
nand U21347 (N_21347,N_19905,N_15213);
and U21348 (N_21348,N_16565,N_16212);
or U21349 (N_21349,N_18585,N_19459);
or U21350 (N_21350,N_15406,N_16214);
xnor U21351 (N_21351,N_18397,N_18982);
xnor U21352 (N_21352,N_19469,N_16071);
nor U21353 (N_21353,N_15678,N_19234);
xnor U21354 (N_21354,N_19085,N_18478);
or U21355 (N_21355,N_17660,N_19698);
or U21356 (N_21356,N_17176,N_17835);
nor U21357 (N_21357,N_18187,N_16475);
nor U21358 (N_21358,N_19528,N_18152);
nor U21359 (N_21359,N_19820,N_17209);
and U21360 (N_21360,N_16429,N_16657);
nand U21361 (N_21361,N_17963,N_16159);
xor U21362 (N_21362,N_18909,N_16957);
and U21363 (N_21363,N_17617,N_16928);
xnor U21364 (N_21364,N_18812,N_16059);
or U21365 (N_21365,N_16769,N_16082);
nand U21366 (N_21366,N_19937,N_19490);
nand U21367 (N_21367,N_15386,N_16965);
or U21368 (N_21368,N_15083,N_15273);
or U21369 (N_21369,N_17273,N_19723);
xor U21370 (N_21370,N_19083,N_16132);
and U21371 (N_21371,N_16917,N_15648);
nor U21372 (N_21372,N_15777,N_15235);
and U21373 (N_21373,N_18210,N_16312);
nor U21374 (N_21374,N_18877,N_19019);
nand U21375 (N_21375,N_15470,N_18320);
nand U21376 (N_21376,N_17165,N_18816);
nand U21377 (N_21377,N_19141,N_18792);
or U21378 (N_21378,N_19105,N_19916);
nand U21379 (N_21379,N_18653,N_17579);
and U21380 (N_21380,N_19847,N_17384);
xnor U21381 (N_21381,N_15351,N_18745);
nand U21382 (N_21382,N_19025,N_16741);
and U21383 (N_21383,N_19580,N_19074);
xor U21384 (N_21384,N_19887,N_17910);
or U21385 (N_21385,N_16439,N_19036);
and U21386 (N_21386,N_19787,N_19598);
nand U21387 (N_21387,N_18813,N_18469);
xor U21388 (N_21388,N_18502,N_19176);
or U21389 (N_21389,N_18947,N_15317);
or U21390 (N_21390,N_17988,N_19210);
or U21391 (N_21391,N_15412,N_16724);
xnor U21392 (N_21392,N_15612,N_16616);
nand U21393 (N_21393,N_19927,N_19504);
xor U21394 (N_21394,N_15095,N_18904);
xnor U21395 (N_21395,N_15609,N_16378);
nand U21396 (N_21396,N_15823,N_17363);
or U21397 (N_21397,N_18654,N_16026);
xnor U21398 (N_21398,N_17822,N_18987);
or U21399 (N_21399,N_16003,N_18276);
xnor U21400 (N_21400,N_16564,N_19759);
nor U21401 (N_21401,N_19569,N_19707);
and U21402 (N_21402,N_16670,N_15571);
nand U21403 (N_21403,N_16845,N_18211);
xor U21404 (N_21404,N_16102,N_18425);
and U21405 (N_21405,N_15862,N_15570);
xnor U21406 (N_21406,N_17972,N_16635);
or U21407 (N_21407,N_16663,N_16650);
xor U21408 (N_21408,N_18951,N_15052);
nand U21409 (N_21409,N_19366,N_19977);
nor U21410 (N_21410,N_15702,N_19330);
nor U21411 (N_21411,N_18603,N_16037);
nand U21412 (N_21412,N_18270,N_16562);
nor U21413 (N_21413,N_17685,N_15258);
xor U21414 (N_21414,N_18473,N_15473);
nand U21415 (N_21415,N_19329,N_19098);
or U21416 (N_21416,N_18007,N_18371);
nor U21417 (N_21417,N_17879,N_18106);
nand U21418 (N_21418,N_16282,N_17892);
nand U21419 (N_21419,N_15099,N_17734);
xor U21420 (N_21420,N_19577,N_17658);
nor U21421 (N_21421,N_19118,N_16318);
nand U21422 (N_21422,N_18134,N_16202);
or U21423 (N_21423,N_18117,N_16658);
and U21424 (N_21424,N_17375,N_16630);
and U21425 (N_21425,N_18824,N_19320);
nand U21426 (N_21426,N_17550,N_19647);
or U21427 (N_21427,N_18226,N_17362);
nand U21428 (N_21428,N_15109,N_17532);
and U21429 (N_21429,N_15563,N_19758);
nand U21430 (N_21430,N_15219,N_16061);
nand U21431 (N_21431,N_18939,N_18059);
nand U21432 (N_21432,N_16089,N_17625);
nor U21433 (N_21433,N_15004,N_16797);
nand U21434 (N_21434,N_15513,N_16005);
nor U21435 (N_21435,N_17407,N_17347);
and U21436 (N_21436,N_15647,N_17405);
nor U21437 (N_21437,N_18483,N_15685);
xor U21438 (N_21438,N_16300,N_18037);
nor U21439 (N_21439,N_15569,N_17649);
and U21440 (N_21440,N_15344,N_16760);
nor U21441 (N_21441,N_17645,N_15950);
and U21442 (N_21442,N_16107,N_19104);
nor U21443 (N_21443,N_18840,N_16461);
or U21444 (N_21444,N_18495,N_15599);
nand U21445 (N_21445,N_19192,N_17985);
xnor U21446 (N_21446,N_17857,N_17756);
nand U21447 (N_21447,N_17121,N_16109);
or U21448 (N_21448,N_19444,N_19151);
nand U21449 (N_21449,N_18542,N_16402);
and U21450 (N_21450,N_15863,N_19486);
nand U21451 (N_21451,N_17486,N_16654);
nor U21452 (N_21452,N_15815,N_17651);
or U21453 (N_21453,N_15009,N_16168);
and U21454 (N_21454,N_16795,N_15745);
or U21455 (N_21455,N_16317,N_19845);
nor U21456 (N_21456,N_16574,N_19531);
nand U21457 (N_21457,N_15793,N_17952);
nand U21458 (N_21458,N_18342,N_18519);
nand U21459 (N_21459,N_18918,N_17352);
xor U21460 (N_21460,N_19858,N_17380);
nor U21461 (N_21461,N_17717,N_18540);
nand U21462 (N_21462,N_15187,N_19567);
or U21463 (N_21463,N_18949,N_18752);
nand U21464 (N_21464,N_15850,N_19254);
nor U21465 (N_21465,N_15105,N_17152);
and U21466 (N_21466,N_15853,N_15782);
nor U21467 (N_21467,N_16148,N_15375);
or U21468 (N_21468,N_15233,N_16445);
nor U21469 (N_21469,N_18334,N_18420);
and U21470 (N_21470,N_16773,N_19499);
nand U21471 (N_21471,N_18402,N_19464);
nor U21472 (N_21472,N_15752,N_15093);
nand U21473 (N_21473,N_16335,N_17777);
nand U21474 (N_21474,N_15488,N_16270);
xor U21475 (N_21475,N_17719,N_19554);
nor U21476 (N_21476,N_17290,N_17307);
and U21477 (N_21477,N_17826,N_17949);
xnor U21478 (N_21478,N_16464,N_15839);
and U21479 (N_21479,N_18850,N_19295);
nor U21480 (N_21480,N_16063,N_19832);
or U21481 (N_21481,N_19166,N_18453);
nor U21482 (N_21482,N_16446,N_16354);
and U21483 (N_21483,N_18629,N_18662);
and U21484 (N_21484,N_19488,N_19460);
xnor U21485 (N_21485,N_17328,N_17538);
nand U21486 (N_21486,N_18071,N_17077);
nand U21487 (N_21487,N_16081,N_17866);
nand U21488 (N_21488,N_16791,N_19934);
and U21489 (N_21489,N_16556,N_17087);
nand U21490 (N_21490,N_17516,N_16017);
nand U21491 (N_21491,N_18393,N_18733);
nor U21492 (N_21492,N_16415,N_15525);
nor U21493 (N_21493,N_15294,N_15512);
nand U21494 (N_21494,N_15407,N_17118);
and U21495 (N_21495,N_17790,N_18098);
and U21496 (N_21496,N_16832,N_19279);
nor U21497 (N_21497,N_18785,N_18716);
xor U21498 (N_21498,N_15783,N_18025);
or U21499 (N_21499,N_19765,N_17250);
nor U21500 (N_21500,N_17360,N_19626);
nor U21501 (N_21501,N_17125,N_18882);
nor U21502 (N_21502,N_15334,N_17110);
and U21503 (N_21503,N_17733,N_18620);
or U21504 (N_21504,N_19725,N_18763);
and U21505 (N_21505,N_18115,N_16456);
or U21506 (N_21506,N_16033,N_19561);
and U21507 (N_21507,N_16768,N_19251);
xnor U21508 (N_21508,N_15558,N_19226);
or U21509 (N_21509,N_15877,N_17339);
nor U21510 (N_21510,N_19877,N_15260);
or U21511 (N_21511,N_15159,N_19507);
and U21512 (N_21512,N_17194,N_16397);
and U21513 (N_21513,N_17057,N_17086);
nor U21514 (N_21514,N_17946,N_17505);
nor U21515 (N_21515,N_19817,N_17106);
nand U21516 (N_21516,N_18490,N_17856);
or U21517 (N_21517,N_19455,N_17925);
nand U21518 (N_21518,N_17932,N_18432);
xor U21519 (N_21519,N_19415,N_19468);
nand U21520 (N_21520,N_18661,N_19779);
nor U21521 (N_21521,N_18796,N_19558);
nand U21522 (N_21522,N_15378,N_17705);
nor U21523 (N_21523,N_19369,N_17129);
nand U21524 (N_21524,N_17827,N_19739);
xor U21525 (N_21525,N_19145,N_19131);
xor U21526 (N_21526,N_17663,N_19819);
xor U21527 (N_21527,N_15858,N_17853);
xnor U21528 (N_21528,N_18765,N_18808);
nor U21529 (N_21529,N_15236,N_16871);
and U21530 (N_21530,N_15956,N_19856);
xor U21531 (N_21531,N_15116,N_17257);
and U21532 (N_21532,N_17264,N_16357);
or U21533 (N_21533,N_15994,N_15073);
and U21534 (N_21534,N_19433,N_19005);
xnor U21535 (N_21535,N_16529,N_15855);
nand U21536 (N_21536,N_15390,N_16906);
or U21537 (N_21537,N_15024,N_15984);
nor U21538 (N_21538,N_18889,N_19810);
nor U21539 (N_21539,N_15785,N_17961);
nor U21540 (N_21540,N_18366,N_16038);
and U21541 (N_21541,N_15459,N_15121);
nor U21542 (N_21542,N_15649,N_16628);
nor U21543 (N_21543,N_19630,N_15808);
nand U21544 (N_21544,N_17410,N_18567);
xor U21545 (N_21545,N_17666,N_18416);
nand U21546 (N_21546,N_17392,N_18592);
xnor U21547 (N_21547,N_15522,N_18687);
xor U21548 (N_21548,N_16572,N_15106);
xnor U21549 (N_21549,N_19954,N_18915);
or U21550 (N_21550,N_17263,N_19245);
and U21551 (N_21551,N_19772,N_17348);
and U21552 (N_21552,N_19893,N_18108);
nor U21553 (N_21553,N_17570,N_15910);
nand U21554 (N_21554,N_15903,N_17052);
nand U21555 (N_21555,N_15251,N_16767);
xor U21556 (N_21556,N_19492,N_15050);
and U21557 (N_21557,N_18669,N_17346);
and U21558 (N_21558,N_17859,N_19988);
nor U21559 (N_21559,N_16295,N_19272);
nor U21560 (N_21560,N_19586,N_15118);
nor U21561 (N_21561,N_18015,N_15679);
nand U21562 (N_21562,N_15472,N_19664);
or U21563 (N_21563,N_18940,N_19515);
and U21564 (N_21564,N_18057,N_16331);
xnor U21565 (N_21565,N_18169,N_19453);
and U21566 (N_21566,N_15246,N_15880);
nor U21567 (N_21567,N_19114,N_16876);
and U21568 (N_21568,N_17076,N_15538);
nor U21569 (N_21569,N_18171,N_15930);
or U21570 (N_21570,N_17724,N_18172);
or U21571 (N_21571,N_16311,N_16913);
nand U21572 (N_21572,N_19335,N_19876);
or U21573 (N_21573,N_15284,N_16501);
nand U21574 (N_21574,N_18175,N_18200);
nor U21575 (N_21575,N_19601,N_17365);
and U21576 (N_21576,N_15070,N_15431);
or U21577 (N_21577,N_16165,N_19315);
and U21578 (N_21578,N_15068,N_17444);
and U21579 (N_21579,N_16874,N_18391);
xnor U21580 (N_21580,N_16237,N_19134);
xor U21581 (N_21581,N_17340,N_19634);
nor U21582 (N_21582,N_16016,N_15861);
or U21583 (N_21583,N_15578,N_18710);
xnor U21584 (N_21584,N_19472,N_18168);
xor U21585 (N_21585,N_18709,N_17237);
or U21586 (N_21586,N_18586,N_15792);
nor U21587 (N_21587,N_17139,N_18116);
xnor U21588 (N_21588,N_17272,N_15748);
or U21589 (N_21589,N_19807,N_16903);
and U21590 (N_21590,N_19184,N_16880);
xor U21591 (N_21591,N_15417,N_15534);
and U21592 (N_21592,N_17297,N_19174);
or U21593 (N_21593,N_16408,N_19952);
and U21594 (N_21594,N_17706,N_19822);
or U21595 (N_21595,N_17597,N_17206);
and U21596 (N_21596,N_15142,N_16821);
or U21597 (N_21597,N_17632,N_19840);
nor U21598 (N_21598,N_17269,N_15524);
or U21599 (N_21599,N_17543,N_17603);
nand U21600 (N_21600,N_16553,N_16921);
xor U21601 (N_21601,N_17213,N_19413);
nand U21602 (N_21602,N_15020,N_19724);
nor U21603 (N_21603,N_18130,N_16695);
nor U21604 (N_21604,N_15811,N_17978);
and U21605 (N_21605,N_19789,N_18417);
nor U21606 (N_21606,N_15196,N_16156);
and U21607 (N_21607,N_16462,N_18509);
xor U21608 (N_21608,N_17303,N_19522);
nand U21609 (N_21609,N_16191,N_15769);
or U21610 (N_21610,N_16612,N_16000);
xnor U21611 (N_21611,N_17700,N_18789);
nand U21612 (N_21612,N_15025,N_15788);
nor U21613 (N_21613,N_16852,N_17762);
xnor U21614 (N_21614,N_17282,N_18153);
and U21615 (N_21615,N_16866,N_19746);
nor U21616 (N_21616,N_17508,N_17433);
xnor U21617 (N_21617,N_19095,N_16073);
and U21618 (N_21618,N_17945,N_19193);
and U21619 (N_21619,N_18718,N_17260);
or U21620 (N_21620,N_19450,N_15295);
and U21621 (N_21621,N_18533,N_19300);
xnor U21622 (N_21622,N_15226,N_17008);
nor U21623 (N_21623,N_15397,N_16054);
and U21624 (N_21624,N_17983,N_15775);
nor U21625 (N_21625,N_18604,N_16911);
or U21626 (N_21626,N_18183,N_17035);
nand U21627 (N_21627,N_16951,N_18161);
and U21628 (N_21628,N_19720,N_17180);
xnor U21629 (N_21629,N_19419,N_16172);
or U21630 (N_21630,N_15717,N_18264);
or U21631 (N_21631,N_18314,N_15485);
nor U21632 (N_21632,N_18002,N_17423);
and U21633 (N_21633,N_15739,N_19266);
or U21634 (N_21634,N_16683,N_17713);
xor U21635 (N_21635,N_17843,N_15906);
xnor U21636 (N_21636,N_16858,N_16742);
and U21637 (N_21637,N_18166,N_18313);
xor U21638 (N_21638,N_15657,N_18354);
or U21639 (N_21639,N_18650,N_15723);
xor U21640 (N_21640,N_15418,N_19367);
nand U21641 (N_21641,N_16346,N_15238);
xor U21642 (N_21642,N_16867,N_18506);
nor U21643 (N_21643,N_17750,N_16598);
xor U21644 (N_21644,N_16351,N_16008);
and U21645 (N_21645,N_16192,N_19688);
nor U21646 (N_21646,N_17523,N_16676);
nand U21647 (N_21647,N_15856,N_15816);
xnor U21648 (N_21648,N_18748,N_15086);
and U21649 (N_21649,N_18914,N_18596);
nand U21650 (N_21650,N_16236,N_16484);
nor U21651 (N_21651,N_16151,N_16307);
and U21652 (N_21652,N_16490,N_18641);
xnor U21653 (N_21653,N_19170,N_15974);
or U21654 (N_21654,N_15909,N_15625);
or U21655 (N_21655,N_18557,N_18232);
nor U21656 (N_21656,N_17862,N_18191);
and U21657 (N_21657,N_18302,N_18960);
nand U21658 (N_21658,N_17556,N_16099);
and U21659 (N_21659,N_16374,N_18553);
nand U21660 (N_21660,N_15178,N_15360);
nand U21661 (N_21661,N_15144,N_18617);
and U21662 (N_21662,N_17142,N_15774);
nand U21663 (N_21663,N_18916,N_18688);
nand U21664 (N_21664,N_16209,N_15208);
nor U21665 (N_21665,N_15148,N_17454);
nor U21666 (N_21666,N_18124,N_15859);
and U21667 (N_21667,N_17774,N_15952);
xnor U21668 (N_21668,N_17262,N_17689);
and U21669 (N_21669,N_17219,N_15555);
nand U21670 (N_21670,N_18736,N_18556);
or U21671 (N_21671,N_16524,N_17612);
nor U21672 (N_21672,N_18646,N_16001);
nor U21673 (N_21673,N_16460,N_15270);
nor U21674 (N_21674,N_16947,N_16154);
and U21675 (N_21675,N_17934,N_15490);
nand U21676 (N_21676,N_16537,N_15710);
xor U21677 (N_21677,N_17722,N_16304);
nand U21678 (N_21678,N_19548,N_15963);
nor U21679 (N_21679,N_19390,N_17699);
and U21680 (N_21680,N_16834,N_15315);
or U21681 (N_21681,N_15917,N_16638);
and U21682 (N_21682,N_17979,N_17610);
xor U21683 (N_21683,N_16933,N_17624);
xnor U21684 (N_21684,N_19316,N_15079);
xnor U21685 (N_21685,N_18111,N_17197);
and U21686 (N_21686,N_18123,N_15156);
nor U21687 (N_21687,N_15682,N_15200);
nand U21688 (N_21688,N_16103,N_18612);
nor U21689 (N_21689,N_17818,N_16943);
or U21690 (N_21690,N_18147,N_15596);
nand U21691 (N_21691,N_17848,N_18494);
nand U21692 (N_21692,N_15790,N_18433);
and U21693 (N_21693,N_18525,N_16333);
or U21694 (N_21694,N_19244,N_19217);
xnor U21695 (N_21695,N_17861,N_15191);
nor U21696 (N_21696,N_15400,N_16256);
nand U21697 (N_21697,N_19344,N_18969);
and U21698 (N_21698,N_17913,N_16746);
or U21699 (N_21699,N_19563,N_19850);
xor U21700 (N_21700,N_17216,N_19337);
xor U21701 (N_21701,N_19641,N_17562);
or U21702 (N_21702,N_17155,N_16247);
nand U21703 (N_21703,N_17432,N_16804);
or U21704 (N_21704,N_16508,N_19523);
nor U21705 (N_21705,N_15852,N_17781);
nor U21706 (N_21706,N_19043,N_18768);
or U21707 (N_21707,N_17229,N_16725);
nand U21708 (N_21708,N_16733,N_17060);
or U21709 (N_21709,N_18806,N_19364);
and U21710 (N_21710,N_15635,N_18498);
nand U21711 (N_21711,N_18256,N_19889);
and U21712 (N_21712,N_16894,N_19181);
or U21713 (N_21713,N_18463,N_17445);
or U21714 (N_21714,N_16907,N_19710);
nand U21715 (N_21715,N_17602,N_16528);
or U21716 (N_21716,N_19695,N_15346);
xor U21717 (N_21717,N_19947,N_15207);
and U21718 (N_21718,N_16229,N_18105);
and U21719 (N_21719,N_15061,N_17832);
nor U21720 (N_21720,N_19075,N_19635);
or U21721 (N_21721,N_15202,N_18841);
nor U21722 (N_21722,N_16257,N_17941);
and U21723 (N_21723,N_19632,N_16642);
xor U21724 (N_21724,N_18310,N_16972);
and U21725 (N_21725,N_16557,N_15922);
and U21726 (N_21726,N_17169,N_16740);
nor U21727 (N_21727,N_15457,N_19511);
or U21728 (N_21728,N_15130,N_17846);
nand U21729 (N_21729,N_16851,N_17995);
nand U21730 (N_21730,N_18196,N_15544);
xor U21731 (N_21731,N_17737,N_16900);
xnor U21732 (N_21732,N_17921,N_19239);
nor U21733 (N_21733,N_15620,N_17786);
nand U21734 (N_21734,N_18378,N_17578);
xnor U21735 (N_21735,N_16369,N_16593);
and U21736 (N_21736,N_17636,N_19394);
and U21737 (N_21737,N_17675,N_16912);
or U21738 (N_21738,N_17991,N_19835);
or U21739 (N_21739,N_17650,N_19120);
xor U21740 (N_21740,N_15986,N_17093);
xor U21741 (N_21741,N_16916,N_19594);
or U21742 (N_21742,N_16424,N_18326);
or U21743 (N_21743,N_17563,N_15566);
or U21744 (N_21744,N_18294,N_16703);
xnor U21745 (N_21745,N_16065,N_17519);
nand U21746 (N_21746,N_18625,N_18012);
nor U21747 (N_21747,N_19087,N_18767);
nor U21748 (N_21748,N_16886,N_16053);
and U21749 (N_21749,N_16751,N_16829);
nand U21750 (N_21750,N_15664,N_16274);
or U21751 (N_21751,N_18164,N_18691);
nor U21752 (N_21752,N_16021,N_15681);
xor U21753 (N_21753,N_18060,N_18766);
nand U21754 (N_21754,N_18026,N_18249);
nor U21755 (N_21755,N_17133,N_16548);
nor U21756 (N_21756,N_18040,N_16381);
or U21757 (N_21757,N_19463,N_16345);
or U21758 (N_21758,N_19259,N_16922);
or U21759 (N_21759,N_18715,N_18190);
xnor U21760 (N_21760,N_17183,N_19147);
nor U21761 (N_21761,N_15908,N_18114);
or U21762 (N_21762,N_16468,N_16803);
nor U21763 (N_21763,N_19055,N_18621);
and U21764 (N_21764,N_16131,N_18833);
nor U21765 (N_21765,N_17446,N_18053);
or U21766 (N_21766,N_18415,N_15584);
xnor U21767 (N_21767,N_19760,N_16974);
nand U21768 (N_21768,N_17539,N_17364);
nor U21769 (N_21769,N_15063,N_16935);
nor U21770 (N_21770,N_17200,N_18078);
nand U21771 (N_21771,N_16783,N_16843);
or U21772 (N_21772,N_17997,N_17960);
nor U21773 (N_21773,N_18910,N_16114);
nor U21774 (N_21774,N_16051,N_18857);
nor U21775 (N_21775,N_16790,N_17740);
nor U21776 (N_21776,N_17914,N_19498);
xor U21777 (N_21777,N_16732,N_17541);
and U21778 (N_21778,N_16522,N_19353);
or U21779 (N_21779,N_18062,N_19128);
or U21780 (N_21780,N_19541,N_18744);
nor U21781 (N_21781,N_18958,N_17554);
or U21782 (N_21782,N_17477,N_18800);
nand U21783 (N_21783,N_19627,N_19129);
nand U21784 (N_21784,N_19039,N_16488);
xnor U21785 (N_21785,N_15381,N_19223);
nor U21786 (N_21786,N_17025,N_17692);
and U21787 (N_21787,N_16084,N_17252);
xnor U21788 (N_21788,N_17461,N_15700);
and U21789 (N_21789,N_16926,N_18449);
nor U21790 (N_21790,N_16761,N_16272);
xnor U21791 (N_21791,N_19938,N_19327);
nand U21792 (N_21792,N_19154,N_19989);
nor U21793 (N_21793,N_17725,N_15194);
nand U21794 (N_21794,N_19326,N_15770);
and U21795 (N_21795,N_19027,N_16526);
nor U21796 (N_21796,N_16244,N_17748);
or U21797 (N_21797,N_19978,N_15683);
and U21798 (N_21798,N_18499,N_16861);
nor U21799 (N_21799,N_19848,N_19851);
xor U21800 (N_21800,N_16792,N_18368);
nand U21801 (N_21801,N_15695,N_15875);
or U21802 (N_21802,N_18446,N_18068);
nand U21803 (N_21803,N_17797,N_19513);
xnor U21804 (N_21804,N_16976,N_15455);
nand U21805 (N_21805,N_19616,N_18221);
or U21806 (N_21806,N_19935,N_17641);
and U21807 (N_21807,N_18888,N_15157);
nor U21808 (N_21808,N_18228,N_19269);
nand U21809 (N_21809,N_17390,N_16444);
nor U21810 (N_21810,N_17058,N_15017);
nor U21811 (N_21811,N_16403,N_19261);
and U21812 (N_21812,N_15966,N_19793);
xnor U21813 (N_21813,N_17537,N_19895);
or U21814 (N_21814,N_15582,N_17195);
or U21815 (N_21815,N_17752,N_15619);
nor U21816 (N_21816,N_16485,N_15791);
nand U21817 (N_21817,N_15597,N_16605);
nand U21818 (N_21818,N_19839,N_17813);
and U21819 (N_21819,N_19532,N_18670);
and U21820 (N_21820,N_19362,N_17208);
nand U21821 (N_21821,N_17281,N_18727);
and U21822 (N_21822,N_16155,N_18633);
and U21823 (N_21823,N_16611,N_16614);
nor U21824 (N_21824,N_19830,N_19092);
or U21825 (N_21825,N_17726,N_18618);
xor U21826 (N_21826,N_18462,N_19247);
or U21827 (N_21827,N_16197,N_18911);
xnor U21828 (N_21828,N_16196,N_15732);
nor U21829 (N_21829,N_15626,N_17806);
xnor U21830 (N_21830,N_19686,N_18394);
nand U21831 (N_21831,N_17595,N_19825);
or U21832 (N_21832,N_17173,N_18862);
and U21833 (N_21833,N_15350,N_17659);
and U21834 (N_21834,N_17233,N_15594);
nor U21835 (N_21835,N_18198,N_19983);
nor U21836 (N_21836,N_15771,N_19653);
nand U21837 (N_21837,N_18061,N_16494);
xor U21838 (N_21838,N_15265,N_17869);
nor U21839 (N_21839,N_15000,N_15481);
xnor U21840 (N_21840,N_16662,N_18284);
nand U21841 (N_21841,N_15299,N_19808);
nor U21842 (N_21842,N_15192,N_18749);
or U21843 (N_21843,N_15237,N_16376);
xor U21844 (N_21844,N_15496,N_15689);
xnor U21845 (N_21845,N_18699,N_16481);
nand U21846 (N_21846,N_19813,N_16225);
or U21847 (N_21847,N_16122,N_16463);
or U21848 (N_21848,N_17851,N_18680);
and U21849 (N_21849,N_15549,N_15794);
or U21850 (N_21850,N_16438,N_17389);
or U21851 (N_21851,N_19976,N_18895);
xnor U21852 (N_21852,N_17709,N_15742);
nor U21853 (N_21853,N_19106,N_15502);
nor U21854 (N_21854,N_18445,N_16075);
and U21855 (N_21855,N_19138,N_18532);
and U21856 (N_21856,N_19179,N_18892);
or U21857 (N_21857,N_17051,N_16941);
nor U21858 (N_21858,N_18500,N_17909);
or U21859 (N_21859,N_18919,N_15973);
or U21860 (N_21860,N_19067,N_18634);
nor U21861 (N_21861,N_18935,N_15870);
and U21862 (N_21862,N_16623,N_17572);
nand U21863 (N_21863,N_19955,N_17873);
nand U21864 (N_21864,N_18685,N_18675);
xnor U21865 (N_21865,N_17942,N_15355);
nand U21866 (N_21866,N_16500,N_17821);
nand U21867 (N_21867,N_15706,N_16004);
or U21868 (N_21868,N_15338,N_18692);
xor U21869 (N_21869,N_16113,N_19208);
nand U21870 (N_21870,N_16115,N_18267);
nand U21871 (N_21871,N_17459,N_16582);
or U21872 (N_21872,N_17482,N_15097);
nand U21873 (N_21873,N_15996,N_16023);
or U21874 (N_21874,N_16015,N_19940);
nor U21875 (N_21875,N_16211,N_15046);
nand U21876 (N_21876,N_19011,N_16127);
and U21877 (N_21877,N_16801,N_17000);
nor U21878 (N_21878,N_17680,N_18489);
or U21879 (N_21879,N_18983,N_19073);
nand U21880 (N_21880,N_17959,N_15911);
xor U21881 (N_21881,N_18522,N_17377);
xor U21882 (N_21882,N_18075,N_16992);
nand U21883 (N_21883,N_18137,N_15112);
nand U21884 (N_21884,N_18073,N_17039);
nand U21885 (N_21885,N_15560,N_19891);
and U21886 (N_21886,N_15972,N_16674);
nor U21887 (N_21887,N_18492,N_19302);
xnor U21888 (N_21888,N_18460,N_16442);
or U21889 (N_21889,N_17096,N_17937);
nand U21890 (N_21890,N_16193,N_18436);
and U21891 (N_21891,N_17825,N_18477);
nor U21892 (N_21892,N_19719,N_16080);
and U21893 (N_21893,N_17712,N_19331);
and U21894 (N_21894,N_18880,N_18318);
or U21895 (N_21895,N_18288,N_17314);
xnor U21896 (N_21896,N_15449,N_19970);
nand U21897 (N_21897,N_17884,N_19672);
or U21898 (N_21898,N_18978,N_19038);
nand U21899 (N_21899,N_18197,N_15730);
and U21900 (N_21900,N_17274,N_15358);
and U21901 (N_21901,N_19645,N_15498);
and U21902 (N_21902,N_18258,N_17771);
nand U21903 (N_21903,N_19556,N_17466);
xnor U21904 (N_21904,N_16055,N_16545);
and U21905 (N_21905,N_16811,N_15143);
nand U21906 (N_21906,N_18206,N_17898);
nor U21907 (N_21907,N_17785,N_16684);
nand U21908 (N_21908,N_15978,N_16240);
or U21909 (N_21909,N_18430,N_16966);
nand U21910 (N_21910,N_16739,N_16097);
and U21911 (N_21911,N_17841,N_17441);
or U21912 (N_21912,N_15038,N_19683);
nand U21913 (N_21913,N_16808,N_16291);
or U21914 (N_21914,N_17078,N_15129);
xor U21915 (N_21915,N_16609,N_17953);
nor U21916 (N_21916,N_19930,N_19932);
nand U21917 (N_21917,N_17628,N_19123);
xor U21918 (N_21918,N_16283,N_16255);
or U21919 (N_21919,N_18243,N_18133);
and U21920 (N_21920,N_16555,N_18069);
or U21921 (N_21921,N_17150,N_17366);
nor U21922 (N_21922,N_18742,N_16491);
or U21923 (N_21923,N_15197,N_17054);
nor U21924 (N_21924,N_15168,N_15458);
xor U21925 (N_21925,N_18695,N_17249);
xnor U21926 (N_21926,N_17981,N_18640);
nor U21927 (N_21927,N_19420,N_16106);
or U21928 (N_21928,N_18428,N_19374);
nand U21929 (N_21929,N_19610,N_15225);
and U21930 (N_21930,N_19265,N_15773);
nor U21931 (N_21931,N_15014,N_15439);
nand U21932 (N_21932,N_18000,N_16651);
xor U21933 (N_21933,N_19750,N_19872);
and U21934 (N_21934,N_15595,N_17068);
and U21935 (N_21935,N_15181,N_18219);
and U21936 (N_21936,N_15526,N_16940);
or U21937 (N_21937,N_18597,N_17545);
xnor U21938 (N_21938,N_19282,N_15138);
and U21939 (N_21939,N_17798,N_18476);
nand U21940 (N_21940,N_17499,N_15896);
nor U21941 (N_21941,N_15849,N_17218);
or U21942 (N_21942,N_16349,N_16220);
nor U21943 (N_21943,N_16881,N_18809);
or U21944 (N_21944,N_17131,N_19311);
and U21945 (N_21945,N_19540,N_18315);
or U21946 (N_21946,N_15864,N_17819);
and U21947 (N_21947,N_19278,N_15425);
xnor U21948 (N_21948,N_16437,N_15335);
and U21949 (N_21949,N_17027,N_18823);
xnor U21950 (N_21950,N_19962,N_15040);
xor U21951 (N_21951,N_18610,N_16685);
or U21952 (N_21952,N_15011,N_18531);
xor U21953 (N_21953,N_15733,N_16772);
and U21954 (N_21954,N_18372,N_19997);
nor U21955 (N_21955,N_16776,N_17893);
nor U21956 (N_21956,N_15332,N_15633);
and U21957 (N_21957,N_17162,N_16713);
nand U21958 (N_21958,N_19853,N_19458);
or U21959 (N_21959,N_18358,N_15297);
xnor U21960 (N_21960,N_15962,N_15394);
or U21961 (N_21961,N_16699,N_16539);
or U21962 (N_21962,N_15309,N_19652);
and U21963 (N_21963,N_17940,N_16134);
nor U21964 (N_21964,N_15537,N_17895);
and U21965 (N_21965,N_16796,N_18339);
nand U21966 (N_21966,N_16648,N_15640);
xor U21967 (N_21967,N_15757,N_15836);
nand U21968 (N_21968,N_16046,N_19137);
or U21969 (N_21969,N_17783,N_17503);
or U21970 (N_21970,N_17967,N_16358);
xor U21971 (N_21971,N_19395,N_18144);
nand U21972 (N_21972,N_15616,N_16328);
xnor U21973 (N_21973,N_17918,N_17270);
and U21974 (N_21974,N_17544,N_18678);
xor U21975 (N_21975,N_17994,N_15951);
or U21976 (N_21976,N_19590,N_18858);
nand U21977 (N_21977,N_17067,N_15216);
xor U21978 (N_21978,N_15487,N_18740);
or U21979 (N_21979,N_16591,N_18266);
nand U21980 (N_21980,N_15092,N_16993);
nand U21981 (N_21981,N_17369,N_15778);
or U21982 (N_21982,N_18859,N_17315);
xor U21983 (N_21983,N_19888,N_15227);
xor U21984 (N_21984,N_17922,N_16149);
xor U21985 (N_21985,N_19599,N_16329);
nand U21986 (N_21986,N_17018,N_19520);
xnor U21987 (N_21987,N_18828,N_16584);
and U21988 (N_21988,N_15851,N_15298);
nand U21989 (N_21989,N_15357,N_17311);
and U21990 (N_21990,N_18234,N_18938);
and U21991 (N_21991,N_15918,N_19679);
nor U21992 (N_21992,N_19336,N_17326);
and U21993 (N_21993,N_18656,N_16029);
nand U21994 (N_21994,N_17253,N_19774);
nand U21995 (N_21995,N_18192,N_18755);
xnor U21996 (N_21996,N_15913,N_19150);
and U21997 (N_21997,N_17112,N_19755);
and U21998 (N_21998,N_15002,N_16072);
and U21999 (N_21999,N_17965,N_17589);
and U22000 (N_22000,N_16436,N_15342);
or U22001 (N_22001,N_18725,N_15045);
and U22002 (N_22002,N_16036,N_19386);
and U22003 (N_22003,N_15286,N_19089);
nor U22004 (N_22004,N_17691,N_18090);
and U22005 (N_22005,N_16955,N_15438);
and U22006 (N_22006,N_15345,N_17584);
nor U22007 (N_22007,N_18233,N_19907);
or U22008 (N_22008,N_18605,N_17164);
and U22009 (N_22009,N_18260,N_19880);
nand U22010 (N_22010,N_19010,N_19687);
and U22011 (N_22011,N_16697,N_19304);
xnor U22012 (N_22012,N_15846,N_15486);
or U22013 (N_22013,N_19111,N_16977);
xor U22014 (N_22014,N_19457,N_19356);
and U22015 (N_22015,N_15799,N_16608);
xnor U22016 (N_22016,N_15810,N_17623);
nor U22017 (N_22017,N_16447,N_15183);
nor U22018 (N_22018,N_15356,N_17013);
nand U22019 (N_22019,N_16288,N_17440);
and U22020 (N_22020,N_18298,N_17468);
and U22021 (N_22021,N_16504,N_17388);
xnor U22022 (N_22022,N_16254,N_15944);
or U22023 (N_22023,N_16978,N_18362);
xor U22024 (N_22024,N_18386,N_15660);
and U22025 (N_22025,N_16857,N_18451);
nand U22026 (N_22026,N_19827,N_18830);
or U22027 (N_22027,N_19821,N_18779);
xor U22028 (N_22028,N_17286,N_17776);
nor U22029 (N_22029,N_18868,N_15696);
and U22030 (N_22030,N_18703,N_15830);
nand U22031 (N_22031,N_18875,N_17828);
xor U22032 (N_22032,N_18855,N_19414);
nand U22033 (N_22033,N_17903,N_15889);
or U22034 (N_22034,N_15651,N_19896);
and U22035 (N_22035,N_15885,N_17715);
or U22036 (N_22036,N_18050,N_19224);
xor U22037 (N_22037,N_17640,N_16373);
and U22038 (N_22038,N_19220,N_17552);
nand U22039 (N_22039,N_16546,N_17094);
xor U22040 (N_22040,N_15220,N_18238);
nor U22041 (N_22041,N_16431,N_16088);
nand U22042 (N_22042,N_16778,N_15203);
xor U22043 (N_22043,N_18475,N_19084);
nor U22044 (N_22044,N_19446,N_17394);
or U22045 (N_22045,N_19631,N_18316);
xor U22046 (N_22046,N_19685,N_15180);
and U22047 (N_22047,N_16139,N_18774);
or U22048 (N_22048,N_16885,N_17836);
or U22049 (N_22049,N_16744,N_18208);
xnor U22050 (N_22050,N_17845,N_18798);
or U22051 (N_22051,N_15699,N_18843);
or U22052 (N_22052,N_19388,N_19402);
nand U22053 (N_22053,N_17547,N_16895);
or U22054 (N_22054,N_18832,N_16482);
xor U22055 (N_22055,N_16854,N_18055);
and U22056 (N_22056,N_18396,N_18259);
xnor U22057 (N_22057,N_18856,N_16770);
or U22058 (N_22058,N_18999,N_19644);
or U22059 (N_22059,N_18131,N_19332);
nor U22060 (N_22060,N_17631,N_15460);
xor U22061 (N_22061,N_16715,N_19555);
nand U22062 (N_22062,N_17629,N_17744);
or U22063 (N_22063,N_18974,N_18810);
nor U22064 (N_22064,N_15084,N_15720);
and U22065 (N_22065,N_15902,N_17788);
nor U22066 (N_22066,N_18170,N_18549);
xnor U22067 (N_22067,N_16096,N_15796);
xnor U22068 (N_22068,N_15005,N_15446);
and U22069 (N_22069,N_18775,N_19591);
xnor U22070 (N_22070,N_15553,N_17987);
xnor U22071 (N_22071,N_15060,N_18003);
or U22072 (N_22072,N_18064,N_18470);
nor U22073 (N_22073,N_15410,N_16121);
and U22074 (N_22074,N_19972,N_19576);
nand U22075 (N_22075,N_16470,N_18545);
nand U22076 (N_22076,N_19387,N_19169);
and U22077 (N_22077,N_16806,N_16809);
nor U22078 (N_22078,N_15624,N_18930);
nand U22079 (N_22079,N_19059,N_15611);
xnor U22080 (N_22080,N_17414,N_18757);
or U22081 (N_22081,N_17936,N_19242);
and U22082 (N_22082,N_17178,N_17555);
xnor U22083 (N_22083,N_15179,N_18548);
nor U22084 (N_22084,N_16387,N_17839);
or U22085 (N_22085,N_18977,N_17931);
or U22086 (N_22086,N_17136,N_18443);
nand U22087 (N_22087,N_18337,N_15312);
nor U22088 (N_22088,N_18013,N_16157);
or U22089 (N_22089,N_18611,N_17881);
nand U22090 (N_22090,N_17449,N_17487);
xnor U22091 (N_22091,N_15259,N_18793);
xor U22092 (N_22092,N_15096,N_19650);
nor U22093 (N_22093,N_15562,N_15873);
and U22094 (N_22094,N_15919,N_16983);
nand U22095 (N_22095,N_17739,N_16507);
xor U22096 (N_22096,N_15281,N_18338);
and U22097 (N_22097,N_15837,N_17608);
nor U22098 (N_22098,N_17172,N_17434);
nor U22099 (N_22099,N_16923,N_16771);
xor U22100 (N_22100,N_16047,N_16370);
and U22101 (N_22101,N_16111,N_18761);
xnor U22102 (N_22102,N_16891,N_18296);
or U22103 (N_22103,N_19861,N_16675);
xnor U22104 (N_22104,N_18178,N_17507);
or U22105 (N_22105,N_18876,N_18045);
nor U22106 (N_22106,N_19442,N_15694);
xnor U22107 (N_22107,N_15658,N_18619);
xor U22108 (N_22108,N_17302,N_17980);
and U22109 (N_22109,N_16223,N_16800);
xnor U22110 (N_22110,N_19666,N_16525);
nor U22111 (N_22111,N_17915,N_15135);
nor U22112 (N_22112,N_17198,N_18306);
or U22113 (N_22113,N_15940,N_15391);
and U22114 (N_22114,N_16530,N_16145);
nor U22115 (N_22115,N_17132,N_19913);
xnor U22116 (N_22116,N_17159,N_17021);
xnor U22117 (N_22117,N_16459,N_15222);
xor U22118 (N_22118,N_16347,N_16302);
nand U22119 (N_22119,N_15600,N_17061);
xor U22120 (N_22120,N_16678,N_17386);
nand U22121 (N_22121,N_15926,N_18448);
nor U22122 (N_22122,N_16364,N_15234);
and U22123 (N_22123,N_18176,N_16607);
or U22124 (N_22124,N_15965,N_15784);
nand U22125 (N_22125,N_18921,N_16506);
or U22126 (N_22126,N_17833,N_18244);
or U22127 (N_22127,N_16262,N_19246);
and U22128 (N_22128,N_17655,N_17671);
xnor U22129 (N_22129,N_17576,N_19483);
nand U22130 (N_22130,N_15043,N_15136);
nor U22131 (N_22131,N_16848,N_19130);
nor U22132 (N_22132,N_17529,N_16615);
and U22133 (N_22133,N_15436,N_19317);
nand U22134 (N_22134,N_19581,N_17490);
xnor U22135 (N_22135,N_16991,N_18526);
and U22136 (N_22136,N_19349,N_16472);
or U22137 (N_22137,N_18236,N_16570);
or U22138 (N_22138,N_19470,N_17494);
and U22139 (N_22139,N_18908,N_16711);
and U22140 (N_22140,N_19117,N_18782);
nand U22141 (N_22141,N_18504,N_18341);
nor U22142 (N_22142,N_18973,N_19423);
and U22143 (N_22143,N_15539,N_19761);
or U22144 (N_22144,N_18039,N_17245);
nand U22145 (N_22145,N_18772,N_17275);
nand U22146 (N_22146,N_15750,N_17397);
and U22147 (N_22147,N_18728,N_16205);
nor U22148 (N_22148,N_19718,N_19412);
nor U22149 (N_22149,N_19831,N_19841);
xor U22150 (N_22150,N_18405,N_15587);
and U22151 (N_22151,N_17002,N_17223);
nand U22152 (N_22152,N_16235,N_18110);
and U22153 (N_22153,N_15961,N_18884);
nor U22154 (N_22154,N_15900,N_19333);
or U22155 (N_22155,N_17738,N_19100);
and U22156 (N_22156,N_15036,N_18269);
and U22157 (N_22157,N_19732,N_18682);
or U22158 (N_22158,N_19347,N_15580);
nor U22159 (N_22159,N_16882,N_18975);
xnor U22160 (N_22160,N_17766,N_16474);
nand U22161 (N_22161,N_18702,N_18049);
nor U22162 (N_22162,N_15376,N_18552);
xor U22163 (N_22163,N_15556,N_17353);
and U22164 (N_22164,N_19116,N_16573);
nand U22165 (N_22165,N_18074,N_15916);
or U22166 (N_22166,N_16998,N_16034);
nand U22167 (N_22167,N_19125,N_18308);
or U22168 (N_22168,N_16362,N_17239);
or U22169 (N_22169,N_17438,N_16855);
xor U22170 (N_22170,N_17950,N_17324);
xor U22171 (N_22171,N_15557,N_18207);
and U22172 (N_22172,N_16561,N_19063);
or U22173 (N_22173,N_19435,N_19186);
or U22174 (N_22174,N_15123,N_18589);
or U22175 (N_22175,N_15993,N_19691);
and U22176 (N_22176,N_15924,N_18994);
xnor U22177 (N_22177,N_16997,N_19411);
nand U22178 (N_22178,N_18681,N_19439);
or U22179 (N_22179,N_16841,N_17031);
nand U22180 (N_22180,N_17849,N_19640);
nor U22181 (N_22181,N_17751,N_17427);
nand U22182 (N_22182,N_19127,N_15415);
nor U22183 (N_22183,N_16407,N_16136);
xor U22184 (N_22184,N_15133,N_18684);
and U22185 (N_22185,N_15110,N_17601);
and U22186 (N_22186,N_17246,N_16505);
or U22187 (N_22187,N_19489,N_19918);
xnor U22188 (N_22188,N_18543,N_19518);
nand U22189 (N_22189,N_19583,N_19911);
and U22190 (N_22190,N_19283,N_19270);
xnor U22191 (N_22191,N_18778,N_15444);
nand U22192 (N_22192,N_19238,N_18122);
nor U22193 (N_22193,N_19017,N_16960);
and U22194 (N_22194,N_18204,N_19159);
nand U22195 (N_22195,N_17585,N_18036);
nand U22196 (N_22196,N_17882,N_18594);
and U22197 (N_22197,N_16027,N_17634);
nand U22198 (N_22198,N_15074,N_16217);
nand U22199 (N_22199,N_17891,N_16385);
xor U22200 (N_22200,N_16389,N_15269);
nand U22201 (N_22201,N_15331,N_16653);
nand U22202 (N_22202,N_17041,N_16332);
nand U22203 (N_22203,N_17116,N_18503);
or U22204 (N_22204,N_19263,N_15545);
nand U22205 (N_22205,N_15835,N_16356);
or U22206 (N_22206,N_18179,N_19473);
nor U22207 (N_22207,N_16379,N_19596);
nand U22208 (N_22208,N_17850,N_15826);
nand U22209 (N_22209,N_16404,N_19741);
nand U22210 (N_22210,N_16807,N_17904);
nor U22211 (N_22211,N_16324,N_19294);
nor U22212 (N_22212,N_15675,N_16087);
and U22213 (N_22213,N_15041,N_19280);
nand U22214 (N_22214,N_18143,N_16340);
nand U22215 (N_22215,N_17385,N_18507);
and U22216 (N_22216,N_19352,N_15606);
nor U22217 (N_22217,N_15673,N_17920);
nand U22218 (N_22218,N_17408,N_15948);
and U22219 (N_22219,N_17926,N_15927);
and U22220 (N_22220,N_15709,N_19620);
nor U22221 (N_22221,N_15749,N_19322);
or U22222 (N_22222,N_19785,N_17970);
and U22223 (N_22223,N_19609,N_15016);
nor U22224 (N_22224,N_18246,N_17050);
nand U22225 (N_22225,N_19044,N_15321);
nor U22226 (N_22226,N_17517,N_15523);
nor U22227 (N_22227,N_17526,N_16995);
nor U22228 (N_22228,N_18352,N_15735);
or U22229 (N_22229,N_15430,N_17598);
nor U22230 (N_22230,N_17871,N_18835);
nand U22231 (N_22231,N_15514,N_18773);
nand U22232 (N_22232,N_16985,N_16873);
nor U22233 (N_22233,N_19478,N_16126);
nand U22234 (N_22234,N_18009,N_19559);
nand U22235 (N_22235,N_17135,N_17860);
xor U22236 (N_22236,N_19109,N_19406);
or U22237 (N_22237,N_16258,N_17356);
nand U22238 (N_22238,N_15035,N_18189);
xnor U22239 (N_22239,N_16920,N_19436);
nand U22240 (N_22240,N_18014,N_19791);
nor U22241 (N_22241,N_19103,N_15511);
xor U22242 (N_22242,N_18355,N_16427);
and U22243 (N_22243,N_17075,N_19421);
and U22244 (N_22244,N_18295,N_17760);
nor U22245 (N_22245,N_16002,N_18142);
or U22246 (N_22246,N_19481,N_16344);
nand U22247 (N_22247,N_19250,N_16617);
nor U22248 (N_22248,N_17287,N_17358);
and U22249 (N_22249,N_17581,N_17418);
xnor U22250 (N_22250,N_19007,N_16816);
and U22251 (N_22251,N_16152,N_18309);
and U22252 (N_22252,N_19862,N_15894);
and U22253 (N_22253,N_17999,N_17805);
xor U22254 (N_22254,N_16458,N_16904);
xnor U22255 (N_22255,N_15491,N_19212);
nand U22256 (N_22256,N_18626,N_18645);
xnor U22257 (N_22257,N_15652,N_16814);
xnor U22258 (N_22258,N_17883,N_17192);
nor U22259 (N_22259,N_16521,N_15161);
and U22260 (N_22260,N_18759,N_19621);
nand U22261 (N_22261,N_19975,N_16206);
or U22262 (N_22262,N_17117,N_15737);
xnor U22263 (N_22263,N_19157,N_15185);
nor U22264 (N_22264,N_18527,N_19982);
or U22265 (N_22265,N_18630,N_18762);
or U22266 (N_22266,N_17382,N_19281);
nand U22267 (N_22267,N_15054,N_17982);
and U22268 (N_22268,N_19704,N_17535);
xnor U22269 (N_22269,N_19805,N_18251);
and U22270 (N_22270,N_18357,N_16909);
xnor U22271 (N_22271,N_18893,N_15456);
nand U22272 (N_22272,N_16731,N_17604);
xnor U22273 (N_22273,N_15462,N_15736);
or U22274 (N_22274,N_17588,N_16585);
or U22275 (N_22275,N_18831,N_16945);
nor U22276 (N_22276,N_16652,N_16728);
or U22277 (N_22277,N_15847,N_15066);
xnor U22278 (N_22278,N_15613,N_16610);
xor U22279 (N_22279,N_17611,N_19585);
xor U22280 (N_22280,N_18411,N_15955);
nand U22281 (N_22281,N_18965,N_17079);
nor U22282 (N_22282,N_15408,N_16275);
xor U22283 (N_22283,N_18890,N_16338);
or U22284 (N_22284,N_16748,N_19348);
nand U22285 (N_22285,N_19177,N_15954);
and U22286 (N_22286,N_16259,N_17955);
and U22287 (N_22287,N_15245,N_17374);
and U22288 (N_22288,N_18817,N_16527);
nor U22289 (N_22289,N_15981,N_18643);
nand U22290 (N_22290,N_16752,N_18241);
and U22291 (N_22291,N_15340,N_16639);
nand U22292 (N_22292,N_16467,N_18584);
xor U22293 (N_22293,N_16443,N_16372);
nand U22294 (N_22294,N_16117,N_18717);
and U22295 (N_22295,N_18714,N_18139);
nand U22296 (N_22296,N_16510,N_18481);
xor U22297 (N_22297,N_18555,N_15941);
nor U22298 (N_22298,N_19945,N_17792);
xor U22299 (N_22299,N_19427,N_16996);
and U22300 (N_22300,N_17163,N_17801);
nor U22301 (N_22301,N_15840,N_18731);
and U22302 (N_22302,N_16067,N_15968);
xnor U22303 (N_22303,N_16656,N_15803);
or U22304 (N_22304,N_17772,N_19991);
xor U22305 (N_22305,N_17398,N_15172);
nor U22306 (N_22306,N_15869,N_18666);
nand U22307 (N_22307,N_19769,N_19855);
nor U22308 (N_22308,N_16226,N_16655);
nor U22309 (N_22309,N_19818,N_15241);
and U22310 (N_22310,N_15641,N_17512);
nand U22311 (N_22311,N_15711,N_16784);
or U22312 (N_22312,N_19178,N_17530);
nand U22313 (N_22313,N_17143,N_19597);
or U22314 (N_22314,N_18970,N_16048);
nand U22315 (N_22315,N_19357,N_15615);
or U22316 (N_22316,N_15691,N_19587);
or U22317 (N_22317,N_17683,N_17036);
and U22318 (N_22318,N_15442,N_19257);
nand U22319 (N_22319,N_16931,N_19603);
or U22320 (N_22320,N_15388,N_15239);
xnor U22321 (N_22321,N_18465,N_15753);
and U22322 (N_22322,N_18387,N_18218);
xor U22323 (N_22323,N_17899,N_16384);
or U22324 (N_22324,N_16897,N_19318);
and U22325 (N_22325,N_17694,N_17900);
xnor U22326 (N_22326,N_16390,N_15535);
xor U22327 (N_22327,N_15528,N_15975);
nor U22328 (N_22328,N_19663,N_17844);
and U22329 (N_22329,N_18109,N_17321);
or U22330 (N_22330,N_17082,N_15798);
and U22331 (N_22331,N_18602,N_17524);
or U22332 (N_22332,N_15154,N_15813);
nor U22333 (N_22333,N_18535,N_15504);
or U22334 (N_22334,N_19908,N_15960);
nand U22335 (N_22335,N_19219,N_19701);
and U22336 (N_22336,N_18058,N_15842);
nand U22337 (N_22337,N_17728,N_15021);
nor U22338 (N_22338,N_19993,N_18992);
and U22339 (N_22339,N_15533,N_15278);
nor U22340 (N_22340,N_15518,N_16052);
and U22341 (N_22341,N_19033,N_16342);
or U22342 (N_22342,N_15119,N_19699);
nor U22343 (N_22343,N_19497,N_18019);
or U22344 (N_22344,N_15708,N_19500);
and U22345 (N_22345,N_16968,N_18485);
and U22346 (N_22346,N_17769,N_16830);
nand U22347 (N_22347,N_19274,N_15820);
and U22348 (N_22348,N_17510,N_16194);
xnor U22349 (N_22349,N_15515,N_18998);
or U22350 (N_22350,N_16919,N_19854);
nor U22351 (N_22351,N_19557,N_19284);
or U22352 (N_22352,N_17956,N_16613);
nand U22353 (N_22353,N_15032,N_19547);
nor U22354 (N_22354,N_17958,N_18458);
and U22355 (N_22355,N_15304,N_16326);
nor U22356 (N_22356,N_17929,N_17590);
and U22357 (N_22357,N_16150,N_15176);
and U22358 (N_22358,N_19708,N_15193);
or U22359 (N_22359,N_18891,N_18419);
nor U22360 (N_22360,N_17599,N_15427);
and U22361 (N_22361,N_16908,N_18029);
and U22362 (N_22362,N_19973,N_18606);
nor U22363 (N_22363,N_17345,N_16449);
xnor U22364 (N_22364,N_19002,N_16836);
and U22365 (N_22365,N_19661,N_17154);
and U22366 (N_22366,N_19508,N_19942);
or U22367 (N_22367,N_17672,N_16634);
nand U22368 (N_22368,N_19960,N_16743);
or U22369 (N_22369,N_15482,N_19462);
xnor U22370 (N_22370,N_18801,N_19648);
nand U22371 (N_22371,N_16434,N_17473);
nand U22372 (N_22372,N_17930,N_16856);
nor U22373 (N_22373,N_19801,N_17333);
nand U22374 (N_22374,N_18188,N_16693);
or U22375 (N_22375,N_16200,N_16646);
and U22376 (N_22376,N_16009,N_15028);
nand U22377 (N_22377,N_15171,N_18753);
nand U22378 (N_22378,N_16889,N_15314);
nor U22379 (N_22379,N_15271,N_18580);
nor U22380 (N_22380,N_16400,N_18118);
xnor U22381 (N_22381,N_19974,N_19321);
xor U22382 (N_22382,N_18627,N_16178);
nor U22383 (N_22383,N_19869,N_17567);
or U22384 (N_22384,N_18322,N_15173);
nor U22385 (N_22385,N_15322,N_16601);
and U22386 (N_22386,N_19021,N_19662);
nor U22387 (N_22387,N_18803,N_19946);
and U22388 (N_22388,N_16163,N_17561);
or U22389 (N_22389,N_16336,N_19639);
nor U22390 (N_22390,N_19539,N_18671);
nor U22391 (N_22391,N_16961,N_19480);
xnor U22392 (N_22392,N_16734,N_18230);
and U22393 (N_22393,N_18927,N_17350);
xnor U22394 (N_22394,N_19144,N_18222);
and U22395 (N_22395,N_15713,N_17161);
xnor U22396 (N_22396,N_19549,N_19777);
nor U22397 (N_22397,N_15592,N_19752);
nor U22398 (N_22398,N_18701,N_17492);
nand U22399 (N_22399,N_17214,N_16701);
xor U22400 (N_22400,N_15936,N_15929);
or U22401 (N_22401,N_16665,N_15738);
nor U22402 (N_22402,N_18980,N_19377);
and U22403 (N_22403,N_18174,N_17033);
nor U22404 (N_22404,N_18044,N_19082);
xor U22405 (N_22405,N_17815,N_15370);
nor U22406 (N_22406,N_19864,N_16698);
nand U22407 (N_22407,N_17452,N_18963);
or U22408 (N_22408,N_17642,N_17071);
xnor U22409 (N_22409,N_16457,N_16723);
nand U22410 (N_22410,N_17401,N_18871);
xnor U22411 (N_22411,N_17476,N_17309);
xnor U22412 (N_22412,N_16679,N_19901);
and U22413 (N_22413,N_18343,N_17417);
or U22414 (N_22414,N_19003,N_17800);
and U22415 (N_22415,N_18622,N_15100);
nor U22416 (N_22416,N_19595,N_18261);
or U22417 (N_22417,N_18311,N_15495);
nor U22418 (N_22418,N_15992,N_15113);
nor U22419 (N_22419,N_16677,N_15127);
nand U22420 (N_22420,N_16309,N_18615);
xnor U22421 (N_22421,N_16386,N_15285);
and U22422 (N_22422,N_16514,N_18319);
nor U22423 (N_22423,N_17644,N_15480);
nor U22424 (N_22424,N_17220,N_17265);
nand U22425 (N_22425,N_16661,N_15134);
xor U22426 (N_22426,N_16967,N_16319);
and U22427 (N_22427,N_17696,N_18722);
nor U22428 (N_22428,N_18336,N_17160);
nor U22429 (N_22429,N_19211,N_15663);
nor U22430 (N_22430,N_19715,N_18849);
or U22431 (N_22431,N_17228,N_19391);
xnor U22432 (N_22432,N_16486,N_16622);
and U22433 (N_22433,N_16520,N_16621);
nand U22434 (N_22434,N_19999,N_17674);
xnor U22435 (N_22435,N_17779,N_19334);
and U22436 (N_22436,N_17897,N_18239);
xor U22437 (N_22437,N_16011,N_19214);
and U22438 (N_22438,N_19132,N_16719);
and U22439 (N_22439,N_18601,N_17238);
nor U22440 (N_22440,N_17406,N_19592);
nand U22441 (N_22441,N_17935,N_18878);
nand U22442 (N_22442,N_15665,N_17770);
or U22443 (N_22443,N_16717,N_17679);
or U22444 (N_22444,N_16316,N_16602);
nor U22445 (N_22445,N_16666,N_15904);
nor U22446 (N_22446,N_19042,N_17403);
or U22447 (N_22447,N_19654,N_15212);
or U22448 (N_22448,N_18438,N_15879);
nor U22449 (N_22449,N_19828,N_16019);
nor U22450 (N_22450,N_18607,N_17065);
or U22451 (N_22451,N_17998,N_19382);
or U22452 (N_22452,N_15602,N_17527);
and U22453 (N_22453,N_19838,N_19372);
or U22454 (N_22454,N_19956,N_15422);
or U22455 (N_22455,N_16586,N_15801);
and U22456 (N_22456,N_18100,N_19899);
nor U22457 (N_22457,N_16077,N_17316);
xor U22458 (N_22458,N_17638,N_16532);
xnor U22459 (N_22459,N_19749,N_18278);
and U22460 (N_22460,N_15887,N_17962);
or U22461 (N_22461,N_15905,N_18906);
or U22462 (N_22462,N_15117,N_18961);
nor U22463 (N_22463,N_16423,N_16493);
nand U22464 (N_22464,N_18461,N_15628);
or U22465 (N_22465,N_18647,N_16910);
nand U22466 (N_22466,N_16161,N_17327);
and U22467 (N_22467,N_19625,N_18693);
xnor U22468 (N_22468,N_16590,N_17115);
and U22469 (N_22469,N_15754,N_16170);
nand U22470 (N_22470,N_18349,N_19447);
nand U22471 (N_22471,N_15586,N_19135);
xor U22472 (N_22472,N_16091,N_18713);
nand U22473 (N_22473,N_15806,N_19705);
and U22474 (N_22474,N_15510,N_17141);
nand U22475 (N_22475,N_17207,N_17553);
or U22476 (N_22476,N_19944,N_18353);
or U22477 (N_22477,N_17217,N_15886);
or U22478 (N_22478,N_16577,N_15575);
or U22479 (N_22479,N_17119,N_17411);
or U22480 (N_22480,N_18863,N_16143);
or U22481 (N_22481,N_19560,N_17755);
or U22482 (N_22482,N_18488,N_19056);
and U22483 (N_22483,N_18568,N_16286);
xor U22484 (N_22484,N_15829,N_17947);
and U22485 (N_22485,N_16975,N_18985);
xor U22486 (N_22486,N_17637,N_17730);
nor U22487 (N_22487,N_19091,N_19325);
xnor U22488 (N_22488,N_19788,N_17676);
xor U22489 (N_22489,N_19448,N_19562);
and U22490 (N_22490,N_19668,N_19437);
nor U22491 (N_22491,N_19026,N_15623);
nor U22492 (N_22492,N_17506,N_15659);
xnor U22493 (N_22493,N_17293,N_16604);
xnor U22494 (N_22494,N_17626,N_15483);
nor U22495 (N_22495,N_16511,N_18344);
nand U22496 (N_22496,N_16315,N_19961);
nor U22497 (N_22497,N_19996,N_16838);
or U22498 (N_22498,N_16323,N_15256);
nor U22499 (N_22499,N_18776,N_19252);
or U22500 (N_22500,N_16433,N_17788);
xnor U22501 (N_22501,N_18350,N_18586);
and U22502 (N_22502,N_16756,N_17484);
and U22503 (N_22503,N_16477,N_18419);
xor U22504 (N_22504,N_15531,N_15950);
xor U22505 (N_22505,N_19634,N_18336);
nor U22506 (N_22506,N_15204,N_19778);
nor U22507 (N_22507,N_19166,N_18050);
nand U22508 (N_22508,N_19058,N_18806);
xnor U22509 (N_22509,N_17515,N_16822);
nor U22510 (N_22510,N_17182,N_19615);
or U22511 (N_22511,N_17138,N_17161);
xor U22512 (N_22512,N_18341,N_16874);
xnor U22513 (N_22513,N_19670,N_19835);
and U22514 (N_22514,N_19328,N_15576);
nor U22515 (N_22515,N_15312,N_18709);
xnor U22516 (N_22516,N_19960,N_19808);
and U22517 (N_22517,N_15474,N_15664);
nand U22518 (N_22518,N_18600,N_18603);
xnor U22519 (N_22519,N_15442,N_17481);
or U22520 (N_22520,N_17111,N_15856);
nor U22521 (N_22521,N_19831,N_16530);
nor U22522 (N_22522,N_16987,N_16931);
nand U22523 (N_22523,N_17608,N_18775);
and U22524 (N_22524,N_18710,N_19832);
nor U22525 (N_22525,N_18641,N_15637);
and U22526 (N_22526,N_15117,N_17331);
xor U22527 (N_22527,N_19757,N_19741);
nand U22528 (N_22528,N_15328,N_17948);
xnor U22529 (N_22529,N_18240,N_18425);
nand U22530 (N_22530,N_19091,N_16318);
or U22531 (N_22531,N_17059,N_15342);
nor U22532 (N_22532,N_18531,N_16797);
nand U22533 (N_22533,N_15937,N_17431);
nand U22534 (N_22534,N_17177,N_19023);
and U22535 (N_22535,N_17812,N_15573);
and U22536 (N_22536,N_18088,N_16643);
nand U22537 (N_22537,N_15257,N_15583);
xor U22538 (N_22538,N_17972,N_15443);
xor U22539 (N_22539,N_15126,N_19861);
or U22540 (N_22540,N_19795,N_17514);
nor U22541 (N_22541,N_15442,N_15512);
nand U22542 (N_22542,N_19048,N_15917);
xnor U22543 (N_22543,N_16684,N_15319);
xnor U22544 (N_22544,N_19367,N_17653);
nor U22545 (N_22545,N_15589,N_18697);
nand U22546 (N_22546,N_18691,N_18309);
or U22547 (N_22547,N_18857,N_15033);
xnor U22548 (N_22548,N_19312,N_17319);
nand U22549 (N_22549,N_16661,N_15924);
xnor U22550 (N_22550,N_17324,N_19671);
xnor U22551 (N_22551,N_19451,N_17763);
or U22552 (N_22552,N_16987,N_18810);
and U22553 (N_22553,N_19732,N_15465);
nor U22554 (N_22554,N_17467,N_16774);
nand U22555 (N_22555,N_18165,N_15473);
xor U22556 (N_22556,N_17438,N_17373);
and U22557 (N_22557,N_19277,N_17953);
or U22558 (N_22558,N_16218,N_17573);
and U22559 (N_22559,N_17369,N_16417);
nand U22560 (N_22560,N_15139,N_17762);
nor U22561 (N_22561,N_16574,N_17920);
nor U22562 (N_22562,N_15462,N_18195);
and U22563 (N_22563,N_16337,N_17600);
nor U22564 (N_22564,N_18851,N_15853);
xor U22565 (N_22565,N_16162,N_18509);
xnor U22566 (N_22566,N_17968,N_18059);
xor U22567 (N_22567,N_17379,N_19934);
nor U22568 (N_22568,N_17087,N_15691);
xnor U22569 (N_22569,N_19429,N_17599);
or U22570 (N_22570,N_19530,N_17903);
or U22571 (N_22571,N_19557,N_19541);
and U22572 (N_22572,N_18189,N_16899);
or U22573 (N_22573,N_18320,N_15977);
nor U22574 (N_22574,N_16973,N_19470);
nor U22575 (N_22575,N_16567,N_18412);
nor U22576 (N_22576,N_18041,N_18682);
or U22577 (N_22577,N_16192,N_19779);
or U22578 (N_22578,N_19837,N_19077);
nand U22579 (N_22579,N_16278,N_16840);
or U22580 (N_22580,N_19767,N_15640);
or U22581 (N_22581,N_19858,N_18591);
nor U22582 (N_22582,N_19050,N_18382);
nor U22583 (N_22583,N_19609,N_16378);
and U22584 (N_22584,N_17495,N_18555);
or U22585 (N_22585,N_15007,N_15975);
nand U22586 (N_22586,N_19866,N_16128);
nand U22587 (N_22587,N_17412,N_16953);
nor U22588 (N_22588,N_19840,N_15026);
and U22589 (N_22589,N_16438,N_18594);
or U22590 (N_22590,N_17928,N_19219);
nor U22591 (N_22591,N_17682,N_18181);
xor U22592 (N_22592,N_19529,N_18691);
or U22593 (N_22593,N_18280,N_18431);
and U22594 (N_22594,N_15824,N_17193);
or U22595 (N_22595,N_18116,N_19194);
nand U22596 (N_22596,N_16771,N_17558);
and U22597 (N_22597,N_17884,N_19879);
xor U22598 (N_22598,N_18648,N_15830);
and U22599 (N_22599,N_16067,N_19432);
nand U22600 (N_22600,N_15234,N_18320);
or U22601 (N_22601,N_16375,N_18880);
nand U22602 (N_22602,N_18444,N_15181);
nor U22603 (N_22603,N_16390,N_15802);
or U22604 (N_22604,N_19725,N_18346);
nor U22605 (N_22605,N_16518,N_18222);
xnor U22606 (N_22606,N_19195,N_17097);
or U22607 (N_22607,N_16134,N_19064);
nor U22608 (N_22608,N_15369,N_19216);
xor U22609 (N_22609,N_19055,N_16966);
nor U22610 (N_22610,N_17968,N_18470);
xnor U22611 (N_22611,N_16972,N_18689);
xnor U22612 (N_22612,N_17647,N_17993);
nand U22613 (N_22613,N_17321,N_16139);
or U22614 (N_22614,N_16995,N_15184);
nand U22615 (N_22615,N_18054,N_16563);
and U22616 (N_22616,N_16683,N_15402);
and U22617 (N_22617,N_19106,N_16229);
nand U22618 (N_22618,N_15920,N_19288);
and U22619 (N_22619,N_16490,N_15857);
and U22620 (N_22620,N_17003,N_16832);
nand U22621 (N_22621,N_15648,N_16467);
nor U22622 (N_22622,N_16271,N_15569);
and U22623 (N_22623,N_19351,N_16062);
nand U22624 (N_22624,N_15895,N_16892);
and U22625 (N_22625,N_16451,N_18511);
nor U22626 (N_22626,N_19996,N_17519);
xnor U22627 (N_22627,N_16334,N_18971);
xor U22628 (N_22628,N_15966,N_19442);
xor U22629 (N_22629,N_16660,N_17543);
and U22630 (N_22630,N_19282,N_15879);
or U22631 (N_22631,N_18309,N_17716);
or U22632 (N_22632,N_15723,N_18878);
xor U22633 (N_22633,N_17722,N_18504);
or U22634 (N_22634,N_16880,N_15305);
and U22635 (N_22635,N_19364,N_16510);
or U22636 (N_22636,N_18736,N_19235);
or U22637 (N_22637,N_17221,N_17117);
nor U22638 (N_22638,N_15545,N_16432);
xor U22639 (N_22639,N_15104,N_15184);
nor U22640 (N_22640,N_15600,N_16729);
nor U22641 (N_22641,N_18662,N_18129);
and U22642 (N_22642,N_18150,N_16842);
xnor U22643 (N_22643,N_18855,N_16113);
nor U22644 (N_22644,N_16961,N_19536);
or U22645 (N_22645,N_16141,N_15755);
nand U22646 (N_22646,N_19652,N_18360);
and U22647 (N_22647,N_15315,N_17321);
nand U22648 (N_22648,N_15711,N_17777);
or U22649 (N_22649,N_15521,N_17554);
or U22650 (N_22650,N_15313,N_15533);
xnor U22651 (N_22651,N_17199,N_17625);
or U22652 (N_22652,N_19364,N_17614);
or U22653 (N_22653,N_19901,N_17163);
xor U22654 (N_22654,N_19654,N_17718);
and U22655 (N_22655,N_16198,N_18547);
nor U22656 (N_22656,N_16238,N_19977);
and U22657 (N_22657,N_17622,N_19028);
nor U22658 (N_22658,N_18742,N_15491);
nor U22659 (N_22659,N_16534,N_17606);
xor U22660 (N_22660,N_17163,N_16679);
xnor U22661 (N_22661,N_15386,N_18156);
nor U22662 (N_22662,N_19576,N_17457);
nand U22663 (N_22663,N_19231,N_16725);
nand U22664 (N_22664,N_15238,N_15867);
xor U22665 (N_22665,N_19840,N_16594);
xor U22666 (N_22666,N_17853,N_15957);
xnor U22667 (N_22667,N_16896,N_16734);
nor U22668 (N_22668,N_19848,N_15138);
nor U22669 (N_22669,N_15179,N_17859);
or U22670 (N_22670,N_18264,N_18466);
nand U22671 (N_22671,N_16731,N_15097);
nand U22672 (N_22672,N_18015,N_16364);
or U22673 (N_22673,N_19649,N_19843);
nor U22674 (N_22674,N_15436,N_18782);
nor U22675 (N_22675,N_17094,N_18806);
xnor U22676 (N_22676,N_15545,N_16404);
nand U22677 (N_22677,N_15953,N_19514);
and U22678 (N_22678,N_15700,N_16614);
nand U22679 (N_22679,N_19925,N_16512);
and U22680 (N_22680,N_17225,N_17588);
nor U22681 (N_22681,N_19352,N_19524);
xor U22682 (N_22682,N_19914,N_17319);
or U22683 (N_22683,N_17743,N_18472);
or U22684 (N_22684,N_15319,N_18121);
nand U22685 (N_22685,N_19591,N_19511);
nand U22686 (N_22686,N_17885,N_18528);
or U22687 (N_22687,N_17243,N_18817);
nor U22688 (N_22688,N_16700,N_17818);
nand U22689 (N_22689,N_18323,N_17923);
nor U22690 (N_22690,N_17285,N_17951);
xor U22691 (N_22691,N_15918,N_18496);
xor U22692 (N_22692,N_18491,N_19234);
nor U22693 (N_22693,N_18301,N_15014);
and U22694 (N_22694,N_18415,N_18140);
nand U22695 (N_22695,N_19390,N_15271);
nand U22696 (N_22696,N_18766,N_15506);
xnor U22697 (N_22697,N_18501,N_17801);
xor U22698 (N_22698,N_18129,N_15384);
and U22699 (N_22699,N_15004,N_15428);
nor U22700 (N_22700,N_16849,N_18433);
nor U22701 (N_22701,N_18341,N_17874);
xor U22702 (N_22702,N_16209,N_18737);
nand U22703 (N_22703,N_18209,N_17809);
nor U22704 (N_22704,N_15683,N_19601);
nor U22705 (N_22705,N_16245,N_16655);
and U22706 (N_22706,N_16459,N_17914);
nand U22707 (N_22707,N_18566,N_15298);
nor U22708 (N_22708,N_17795,N_16425);
nor U22709 (N_22709,N_15253,N_19055);
and U22710 (N_22710,N_17818,N_17734);
nand U22711 (N_22711,N_19627,N_17521);
nand U22712 (N_22712,N_18337,N_19790);
xnor U22713 (N_22713,N_19884,N_15641);
nor U22714 (N_22714,N_18592,N_16607);
or U22715 (N_22715,N_19476,N_16327);
nand U22716 (N_22716,N_17199,N_16890);
or U22717 (N_22717,N_19587,N_16808);
xor U22718 (N_22718,N_15791,N_19480);
or U22719 (N_22719,N_19945,N_15656);
or U22720 (N_22720,N_16537,N_16532);
nor U22721 (N_22721,N_18039,N_15958);
nand U22722 (N_22722,N_15031,N_18848);
nor U22723 (N_22723,N_16548,N_17780);
nand U22724 (N_22724,N_16658,N_15688);
or U22725 (N_22725,N_19554,N_15238);
xnor U22726 (N_22726,N_16454,N_15259);
and U22727 (N_22727,N_17701,N_17881);
nand U22728 (N_22728,N_15500,N_15607);
or U22729 (N_22729,N_17644,N_19823);
xor U22730 (N_22730,N_17800,N_17466);
nor U22731 (N_22731,N_18520,N_16914);
xor U22732 (N_22732,N_15667,N_17405);
and U22733 (N_22733,N_17905,N_19012);
or U22734 (N_22734,N_17120,N_15629);
nor U22735 (N_22735,N_19776,N_15562);
and U22736 (N_22736,N_18191,N_17570);
xnor U22737 (N_22737,N_18529,N_17071);
and U22738 (N_22738,N_19436,N_18805);
xnor U22739 (N_22739,N_17874,N_15367);
and U22740 (N_22740,N_19058,N_16261);
and U22741 (N_22741,N_19661,N_15133);
nand U22742 (N_22742,N_18314,N_19430);
xor U22743 (N_22743,N_18656,N_16571);
nand U22744 (N_22744,N_16074,N_17113);
nor U22745 (N_22745,N_19841,N_15724);
nor U22746 (N_22746,N_15743,N_16925);
xnor U22747 (N_22747,N_16437,N_15846);
xnor U22748 (N_22748,N_17285,N_18678);
or U22749 (N_22749,N_17180,N_16113);
xor U22750 (N_22750,N_19645,N_16585);
nand U22751 (N_22751,N_18316,N_19048);
xor U22752 (N_22752,N_15971,N_19823);
or U22753 (N_22753,N_16686,N_18192);
nand U22754 (N_22754,N_15738,N_16030);
and U22755 (N_22755,N_15383,N_16290);
nand U22756 (N_22756,N_15966,N_17112);
and U22757 (N_22757,N_19971,N_19698);
nor U22758 (N_22758,N_18885,N_16129);
or U22759 (N_22759,N_16992,N_15319);
and U22760 (N_22760,N_17209,N_17426);
nand U22761 (N_22761,N_18667,N_19266);
xnor U22762 (N_22762,N_19847,N_17909);
or U22763 (N_22763,N_18081,N_19057);
nor U22764 (N_22764,N_18658,N_15051);
and U22765 (N_22765,N_16256,N_16833);
or U22766 (N_22766,N_19301,N_16621);
nor U22767 (N_22767,N_18728,N_15498);
xnor U22768 (N_22768,N_16783,N_15914);
xor U22769 (N_22769,N_18452,N_15241);
xnor U22770 (N_22770,N_19519,N_16796);
xnor U22771 (N_22771,N_18346,N_17724);
and U22772 (N_22772,N_15766,N_15956);
nor U22773 (N_22773,N_15173,N_16765);
nor U22774 (N_22774,N_17695,N_16670);
or U22775 (N_22775,N_15409,N_15509);
nor U22776 (N_22776,N_18535,N_17714);
and U22777 (N_22777,N_19770,N_17790);
xnor U22778 (N_22778,N_17009,N_18285);
nand U22779 (N_22779,N_15371,N_19418);
nand U22780 (N_22780,N_15278,N_15479);
xor U22781 (N_22781,N_18817,N_19524);
xnor U22782 (N_22782,N_17589,N_17694);
and U22783 (N_22783,N_17837,N_17456);
nand U22784 (N_22784,N_17878,N_16576);
and U22785 (N_22785,N_15943,N_18517);
or U22786 (N_22786,N_19706,N_16696);
nor U22787 (N_22787,N_15449,N_15859);
nand U22788 (N_22788,N_18004,N_18099);
or U22789 (N_22789,N_16778,N_16477);
and U22790 (N_22790,N_15638,N_16445);
nor U22791 (N_22791,N_18191,N_17386);
or U22792 (N_22792,N_17444,N_16316);
nor U22793 (N_22793,N_18941,N_17845);
nor U22794 (N_22794,N_15884,N_16382);
xnor U22795 (N_22795,N_19387,N_15561);
nand U22796 (N_22796,N_15489,N_17289);
nor U22797 (N_22797,N_17994,N_18241);
nand U22798 (N_22798,N_17201,N_19543);
nor U22799 (N_22799,N_17051,N_18232);
xnor U22800 (N_22800,N_17864,N_17566);
or U22801 (N_22801,N_18875,N_16256);
nand U22802 (N_22802,N_19700,N_17876);
or U22803 (N_22803,N_19109,N_18012);
or U22804 (N_22804,N_17070,N_15900);
or U22805 (N_22805,N_15569,N_16637);
and U22806 (N_22806,N_16428,N_16677);
nor U22807 (N_22807,N_18659,N_15733);
nand U22808 (N_22808,N_16040,N_17153);
xor U22809 (N_22809,N_15712,N_18244);
xor U22810 (N_22810,N_19688,N_16578);
xnor U22811 (N_22811,N_16214,N_17013);
or U22812 (N_22812,N_16645,N_16931);
or U22813 (N_22813,N_18483,N_16766);
or U22814 (N_22814,N_16087,N_16439);
and U22815 (N_22815,N_15130,N_15375);
nor U22816 (N_22816,N_18992,N_16318);
nor U22817 (N_22817,N_17556,N_18701);
or U22818 (N_22818,N_18824,N_18862);
or U22819 (N_22819,N_15047,N_19397);
and U22820 (N_22820,N_16866,N_15451);
nor U22821 (N_22821,N_19427,N_15313);
nand U22822 (N_22822,N_15991,N_15381);
nand U22823 (N_22823,N_17679,N_19099);
xnor U22824 (N_22824,N_17166,N_19617);
nand U22825 (N_22825,N_18967,N_19372);
and U22826 (N_22826,N_18014,N_17799);
nor U22827 (N_22827,N_16132,N_16817);
nor U22828 (N_22828,N_19885,N_18596);
nand U22829 (N_22829,N_19390,N_15640);
and U22830 (N_22830,N_18470,N_18158);
nand U22831 (N_22831,N_18435,N_15637);
or U22832 (N_22832,N_19382,N_17181);
xnor U22833 (N_22833,N_19961,N_18672);
xor U22834 (N_22834,N_18618,N_16731);
nor U22835 (N_22835,N_16086,N_16791);
xor U22836 (N_22836,N_19709,N_15568);
xnor U22837 (N_22837,N_18974,N_15505);
nand U22838 (N_22838,N_19725,N_15426);
nand U22839 (N_22839,N_18886,N_17179);
and U22840 (N_22840,N_16401,N_17667);
nand U22841 (N_22841,N_16150,N_18264);
nor U22842 (N_22842,N_18080,N_18876);
xor U22843 (N_22843,N_16126,N_17762);
nor U22844 (N_22844,N_15601,N_16183);
nand U22845 (N_22845,N_17459,N_17617);
nand U22846 (N_22846,N_18364,N_19657);
or U22847 (N_22847,N_16046,N_19897);
xor U22848 (N_22848,N_16883,N_18113);
nor U22849 (N_22849,N_16901,N_16001);
xnor U22850 (N_22850,N_18165,N_19546);
xnor U22851 (N_22851,N_19297,N_15353);
xnor U22852 (N_22852,N_15498,N_15962);
and U22853 (N_22853,N_19111,N_15707);
and U22854 (N_22854,N_16633,N_18972);
nand U22855 (N_22855,N_15239,N_16519);
nand U22856 (N_22856,N_19738,N_16463);
xor U22857 (N_22857,N_15630,N_15813);
and U22858 (N_22858,N_17178,N_15179);
nand U22859 (N_22859,N_17407,N_16252);
or U22860 (N_22860,N_19114,N_18966);
xor U22861 (N_22861,N_16795,N_19844);
or U22862 (N_22862,N_17025,N_19378);
and U22863 (N_22863,N_16829,N_16121);
nand U22864 (N_22864,N_19468,N_18786);
nand U22865 (N_22865,N_17668,N_15186);
nor U22866 (N_22866,N_18842,N_19134);
and U22867 (N_22867,N_15667,N_17158);
xor U22868 (N_22868,N_18472,N_18276);
and U22869 (N_22869,N_19801,N_17608);
and U22870 (N_22870,N_17393,N_18012);
nand U22871 (N_22871,N_19834,N_17757);
or U22872 (N_22872,N_19831,N_15030);
nor U22873 (N_22873,N_16666,N_16635);
or U22874 (N_22874,N_15417,N_16733);
nand U22875 (N_22875,N_16212,N_16441);
and U22876 (N_22876,N_17100,N_16821);
xor U22877 (N_22877,N_15786,N_15555);
or U22878 (N_22878,N_15917,N_19843);
and U22879 (N_22879,N_18567,N_19890);
nand U22880 (N_22880,N_19156,N_17111);
nor U22881 (N_22881,N_18421,N_18953);
or U22882 (N_22882,N_17250,N_19751);
and U22883 (N_22883,N_16966,N_17550);
nand U22884 (N_22884,N_17183,N_17638);
and U22885 (N_22885,N_16091,N_18770);
or U22886 (N_22886,N_15447,N_15472);
nand U22887 (N_22887,N_18410,N_15418);
nor U22888 (N_22888,N_18962,N_18249);
xnor U22889 (N_22889,N_17375,N_17800);
and U22890 (N_22890,N_17137,N_18850);
nor U22891 (N_22891,N_17899,N_17257);
or U22892 (N_22892,N_19826,N_17061);
and U22893 (N_22893,N_19290,N_18776);
nor U22894 (N_22894,N_15076,N_18268);
nor U22895 (N_22895,N_17758,N_17155);
nand U22896 (N_22896,N_16521,N_15782);
xnor U22897 (N_22897,N_15368,N_17773);
and U22898 (N_22898,N_15161,N_18660);
and U22899 (N_22899,N_17337,N_15160);
xor U22900 (N_22900,N_18589,N_15931);
nand U22901 (N_22901,N_18591,N_17684);
or U22902 (N_22902,N_17797,N_16308);
and U22903 (N_22903,N_17181,N_17027);
nand U22904 (N_22904,N_18023,N_18522);
xor U22905 (N_22905,N_17634,N_18011);
xnor U22906 (N_22906,N_17729,N_17979);
or U22907 (N_22907,N_15316,N_17791);
nor U22908 (N_22908,N_15017,N_19400);
and U22909 (N_22909,N_17902,N_17745);
nand U22910 (N_22910,N_17382,N_16266);
nor U22911 (N_22911,N_17416,N_18502);
or U22912 (N_22912,N_19526,N_15321);
or U22913 (N_22913,N_15175,N_17715);
or U22914 (N_22914,N_15119,N_19236);
nor U22915 (N_22915,N_15627,N_19890);
or U22916 (N_22916,N_18521,N_16348);
or U22917 (N_22917,N_17285,N_16162);
xnor U22918 (N_22918,N_19284,N_18673);
nand U22919 (N_22919,N_19183,N_15521);
nand U22920 (N_22920,N_15588,N_15189);
xnor U22921 (N_22921,N_18295,N_19238);
nor U22922 (N_22922,N_18424,N_16934);
or U22923 (N_22923,N_19404,N_19387);
xor U22924 (N_22924,N_17358,N_19400);
and U22925 (N_22925,N_19848,N_19904);
or U22926 (N_22926,N_19855,N_16352);
nand U22927 (N_22927,N_18008,N_19986);
and U22928 (N_22928,N_18932,N_16339);
nor U22929 (N_22929,N_16997,N_19209);
xor U22930 (N_22930,N_15503,N_15458);
or U22931 (N_22931,N_16224,N_19509);
and U22932 (N_22932,N_15789,N_15486);
nand U22933 (N_22933,N_18629,N_17936);
and U22934 (N_22934,N_16979,N_15276);
nand U22935 (N_22935,N_19304,N_15444);
nand U22936 (N_22936,N_15146,N_17518);
or U22937 (N_22937,N_19784,N_15119);
nand U22938 (N_22938,N_15302,N_18753);
nor U22939 (N_22939,N_17458,N_15901);
and U22940 (N_22940,N_16253,N_15120);
and U22941 (N_22941,N_17904,N_17722);
xnor U22942 (N_22942,N_18329,N_19828);
xnor U22943 (N_22943,N_15162,N_19008);
nand U22944 (N_22944,N_17066,N_19205);
nand U22945 (N_22945,N_16758,N_18235);
or U22946 (N_22946,N_19702,N_19181);
or U22947 (N_22947,N_19066,N_18901);
xor U22948 (N_22948,N_15896,N_17278);
and U22949 (N_22949,N_18443,N_18127);
or U22950 (N_22950,N_17477,N_16913);
nor U22951 (N_22951,N_15715,N_16414);
nor U22952 (N_22952,N_16146,N_18112);
and U22953 (N_22953,N_16029,N_15385);
nor U22954 (N_22954,N_19441,N_16628);
and U22955 (N_22955,N_19523,N_17395);
and U22956 (N_22956,N_15630,N_18997);
nand U22957 (N_22957,N_18738,N_17069);
or U22958 (N_22958,N_17173,N_18273);
nand U22959 (N_22959,N_16131,N_18875);
nor U22960 (N_22960,N_19310,N_17909);
or U22961 (N_22961,N_16485,N_19331);
or U22962 (N_22962,N_16988,N_16737);
nor U22963 (N_22963,N_18932,N_19558);
nand U22964 (N_22964,N_19115,N_19337);
nand U22965 (N_22965,N_16530,N_18174);
nand U22966 (N_22966,N_18388,N_16017);
nand U22967 (N_22967,N_17475,N_15886);
or U22968 (N_22968,N_15716,N_16553);
and U22969 (N_22969,N_17549,N_16043);
nand U22970 (N_22970,N_15769,N_15261);
or U22971 (N_22971,N_19128,N_15007);
xnor U22972 (N_22972,N_18801,N_16012);
and U22973 (N_22973,N_16661,N_15183);
xnor U22974 (N_22974,N_17968,N_16596);
nor U22975 (N_22975,N_16029,N_15293);
or U22976 (N_22976,N_19616,N_19550);
or U22977 (N_22977,N_17148,N_16042);
nand U22978 (N_22978,N_16767,N_18649);
nor U22979 (N_22979,N_18386,N_17041);
and U22980 (N_22980,N_15805,N_17676);
or U22981 (N_22981,N_17258,N_19298);
and U22982 (N_22982,N_15431,N_15121);
or U22983 (N_22983,N_15228,N_18547);
nand U22984 (N_22984,N_16549,N_17100);
or U22985 (N_22985,N_16989,N_15183);
nor U22986 (N_22986,N_18720,N_18288);
nor U22987 (N_22987,N_15570,N_15169);
or U22988 (N_22988,N_19580,N_15508);
and U22989 (N_22989,N_19739,N_19882);
and U22990 (N_22990,N_17140,N_17094);
xor U22991 (N_22991,N_17683,N_18507);
and U22992 (N_22992,N_17608,N_17757);
xnor U22993 (N_22993,N_16735,N_15797);
and U22994 (N_22994,N_16121,N_15450);
and U22995 (N_22995,N_19499,N_15226);
xnor U22996 (N_22996,N_18736,N_16601);
xor U22997 (N_22997,N_17872,N_15539);
nand U22998 (N_22998,N_16296,N_16695);
and U22999 (N_22999,N_19739,N_19194);
nand U23000 (N_23000,N_18759,N_19711);
nand U23001 (N_23001,N_15320,N_18988);
and U23002 (N_23002,N_15798,N_18215);
nand U23003 (N_23003,N_17176,N_15760);
xnor U23004 (N_23004,N_17049,N_16505);
nor U23005 (N_23005,N_17092,N_16766);
nor U23006 (N_23006,N_15745,N_19114);
nand U23007 (N_23007,N_19086,N_19119);
xor U23008 (N_23008,N_18885,N_15365);
and U23009 (N_23009,N_17910,N_17531);
and U23010 (N_23010,N_17032,N_18579);
nor U23011 (N_23011,N_19161,N_18082);
or U23012 (N_23012,N_18723,N_18189);
and U23013 (N_23013,N_19899,N_15593);
nor U23014 (N_23014,N_15417,N_15195);
xor U23015 (N_23015,N_17004,N_18296);
xor U23016 (N_23016,N_19785,N_15033);
xnor U23017 (N_23017,N_15173,N_18486);
nor U23018 (N_23018,N_16676,N_19842);
or U23019 (N_23019,N_18560,N_15814);
or U23020 (N_23020,N_18270,N_19450);
xnor U23021 (N_23021,N_16085,N_18365);
and U23022 (N_23022,N_16392,N_17719);
nand U23023 (N_23023,N_19685,N_19442);
or U23024 (N_23024,N_18303,N_16429);
nor U23025 (N_23025,N_18189,N_15327);
xnor U23026 (N_23026,N_16920,N_18134);
or U23027 (N_23027,N_15665,N_18428);
and U23028 (N_23028,N_19417,N_16596);
nand U23029 (N_23029,N_19494,N_19000);
xor U23030 (N_23030,N_16933,N_17743);
and U23031 (N_23031,N_15396,N_17536);
or U23032 (N_23032,N_18107,N_16012);
and U23033 (N_23033,N_16120,N_18372);
and U23034 (N_23034,N_18283,N_16768);
nor U23035 (N_23035,N_19768,N_19892);
nand U23036 (N_23036,N_17407,N_16026);
xor U23037 (N_23037,N_19754,N_19432);
nand U23038 (N_23038,N_18690,N_17544);
nor U23039 (N_23039,N_19227,N_16052);
nand U23040 (N_23040,N_16220,N_16610);
and U23041 (N_23041,N_15302,N_16100);
nand U23042 (N_23042,N_18914,N_19504);
nor U23043 (N_23043,N_16442,N_19686);
and U23044 (N_23044,N_18675,N_16975);
xnor U23045 (N_23045,N_16030,N_16909);
xnor U23046 (N_23046,N_15275,N_19147);
nor U23047 (N_23047,N_17923,N_19153);
nand U23048 (N_23048,N_15106,N_19044);
nor U23049 (N_23049,N_15911,N_16563);
and U23050 (N_23050,N_16096,N_16775);
nand U23051 (N_23051,N_15081,N_17638);
or U23052 (N_23052,N_15010,N_17491);
or U23053 (N_23053,N_15276,N_17867);
nor U23054 (N_23054,N_16619,N_15304);
xor U23055 (N_23055,N_19949,N_19228);
nand U23056 (N_23056,N_17317,N_19523);
nor U23057 (N_23057,N_15729,N_17595);
or U23058 (N_23058,N_15543,N_16768);
xnor U23059 (N_23059,N_15091,N_16239);
and U23060 (N_23060,N_19855,N_16575);
nand U23061 (N_23061,N_18207,N_16474);
or U23062 (N_23062,N_17387,N_18870);
nor U23063 (N_23063,N_18505,N_16993);
nand U23064 (N_23064,N_15374,N_16668);
xor U23065 (N_23065,N_16506,N_18801);
or U23066 (N_23066,N_17934,N_19747);
nand U23067 (N_23067,N_16978,N_18000);
xnor U23068 (N_23068,N_17227,N_17979);
xnor U23069 (N_23069,N_19129,N_19887);
nor U23070 (N_23070,N_17039,N_17133);
or U23071 (N_23071,N_17062,N_18826);
nor U23072 (N_23072,N_15791,N_15096);
nor U23073 (N_23073,N_19684,N_16945);
or U23074 (N_23074,N_17779,N_16070);
or U23075 (N_23075,N_15965,N_17866);
and U23076 (N_23076,N_18686,N_15972);
nor U23077 (N_23077,N_16501,N_16991);
or U23078 (N_23078,N_15605,N_15004);
nor U23079 (N_23079,N_15723,N_19397);
and U23080 (N_23080,N_19344,N_17424);
and U23081 (N_23081,N_18604,N_16364);
and U23082 (N_23082,N_16679,N_19858);
and U23083 (N_23083,N_19141,N_18007);
nand U23084 (N_23084,N_17607,N_15935);
nor U23085 (N_23085,N_17382,N_16905);
xor U23086 (N_23086,N_19995,N_17434);
nand U23087 (N_23087,N_19261,N_19439);
nand U23088 (N_23088,N_18228,N_16973);
xnor U23089 (N_23089,N_19840,N_18210);
and U23090 (N_23090,N_19196,N_16037);
and U23091 (N_23091,N_16797,N_18724);
or U23092 (N_23092,N_18615,N_16896);
nand U23093 (N_23093,N_17931,N_17522);
nand U23094 (N_23094,N_19053,N_18328);
nand U23095 (N_23095,N_15916,N_15412);
or U23096 (N_23096,N_17584,N_19211);
and U23097 (N_23097,N_16161,N_18946);
nand U23098 (N_23098,N_18253,N_19679);
nor U23099 (N_23099,N_17743,N_17423);
xor U23100 (N_23100,N_15015,N_15829);
nand U23101 (N_23101,N_15966,N_17566);
nor U23102 (N_23102,N_16259,N_17817);
nand U23103 (N_23103,N_16929,N_16804);
or U23104 (N_23104,N_17980,N_19537);
nor U23105 (N_23105,N_15876,N_17027);
xnor U23106 (N_23106,N_17135,N_16187);
or U23107 (N_23107,N_18501,N_19161);
and U23108 (N_23108,N_15107,N_15182);
nor U23109 (N_23109,N_15169,N_18239);
xnor U23110 (N_23110,N_15661,N_18419);
xor U23111 (N_23111,N_17918,N_15883);
nand U23112 (N_23112,N_19524,N_17639);
nand U23113 (N_23113,N_19915,N_15885);
nor U23114 (N_23114,N_19536,N_16011);
nor U23115 (N_23115,N_16188,N_19486);
and U23116 (N_23116,N_15993,N_17200);
and U23117 (N_23117,N_15758,N_19327);
or U23118 (N_23118,N_17026,N_18959);
xnor U23119 (N_23119,N_15079,N_18376);
and U23120 (N_23120,N_18745,N_19104);
xnor U23121 (N_23121,N_19415,N_16885);
nor U23122 (N_23122,N_17126,N_15710);
nand U23123 (N_23123,N_19477,N_17520);
nor U23124 (N_23124,N_18527,N_15249);
nor U23125 (N_23125,N_19306,N_19493);
or U23126 (N_23126,N_19508,N_15674);
nor U23127 (N_23127,N_17664,N_15986);
or U23128 (N_23128,N_18364,N_15135);
and U23129 (N_23129,N_15464,N_18598);
nand U23130 (N_23130,N_16785,N_17048);
nor U23131 (N_23131,N_15493,N_18692);
and U23132 (N_23132,N_17285,N_18117);
and U23133 (N_23133,N_16818,N_19065);
and U23134 (N_23134,N_15473,N_19144);
nor U23135 (N_23135,N_19805,N_17245);
and U23136 (N_23136,N_18709,N_18226);
nand U23137 (N_23137,N_16010,N_16931);
nor U23138 (N_23138,N_15496,N_19001);
nor U23139 (N_23139,N_18853,N_17219);
or U23140 (N_23140,N_18285,N_19874);
xnor U23141 (N_23141,N_15836,N_19708);
or U23142 (N_23142,N_15878,N_15103);
xor U23143 (N_23143,N_15867,N_15110);
nand U23144 (N_23144,N_15616,N_15465);
or U23145 (N_23145,N_16976,N_19843);
or U23146 (N_23146,N_16405,N_19828);
xor U23147 (N_23147,N_16761,N_17198);
xnor U23148 (N_23148,N_19935,N_15137);
xor U23149 (N_23149,N_15054,N_18177);
nor U23150 (N_23150,N_15985,N_15301);
or U23151 (N_23151,N_17200,N_17089);
xnor U23152 (N_23152,N_19975,N_18650);
nand U23153 (N_23153,N_15646,N_17144);
xor U23154 (N_23154,N_16195,N_16428);
nand U23155 (N_23155,N_18006,N_17013);
nand U23156 (N_23156,N_17699,N_19242);
and U23157 (N_23157,N_15312,N_15058);
xor U23158 (N_23158,N_15576,N_16470);
nand U23159 (N_23159,N_16938,N_15479);
xor U23160 (N_23160,N_17432,N_18240);
and U23161 (N_23161,N_19260,N_18986);
and U23162 (N_23162,N_16984,N_19459);
or U23163 (N_23163,N_15624,N_19666);
nand U23164 (N_23164,N_16274,N_18114);
and U23165 (N_23165,N_17520,N_16646);
nor U23166 (N_23166,N_19564,N_19518);
nor U23167 (N_23167,N_16466,N_15624);
nand U23168 (N_23168,N_19994,N_16995);
nor U23169 (N_23169,N_18974,N_19396);
and U23170 (N_23170,N_15431,N_19035);
nand U23171 (N_23171,N_18780,N_17635);
or U23172 (N_23172,N_18923,N_17638);
xor U23173 (N_23173,N_17631,N_15522);
nor U23174 (N_23174,N_18192,N_15490);
and U23175 (N_23175,N_19250,N_19341);
or U23176 (N_23176,N_17101,N_17011);
or U23177 (N_23177,N_18483,N_19943);
nand U23178 (N_23178,N_19112,N_19289);
and U23179 (N_23179,N_17553,N_18966);
and U23180 (N_23180,N_15565,N_17897);
nor U23181 (N_23181,N_19339,N_19718);
nor U23182 (N_23182,N_15309,N_19044);
and U23183 (N_23183,N_17903,N_18787);
xnor U23184 (N_23184,N_17110,N_16626);
nand U23185 (N_23185,N_15407,N_18254);
nand U23186 (N_23186,N_17915,N_18487);
nand U23187 (N_23187,N_15283,N_18073);
xnor U23188 (N_23188,N_18860,N_16503);
and U23189 (N_23189,N_15769,N_16207);
xor U23190 (N_23190,N_18592,N_16328);
or U23191 (N_23191,N_19354,N_17881);
and U23192 (N_23192,N_19681,N_17488);
nor U23193 (N_23193,N_17207,N_16231);
nor U23194 (N_23194,N_18130,N_16717);
or U23195 (N_23195,N_19031,N_15655);
nand U23196 (N_23196,N_18216,N_16492);
or U23197 (N_23197,N_17793,N_15181);
nand U23198 (N_23198,N_15065,N_19619);
and U23199 (N_23199,N_16459,N_19990);
nor U23200 (N_23200,N_16727,N_15866);
nor U23201 (N_23201,N_18724,N_19032);
and U23202 (N_23202,N_16253,N_19314);
nand U23203 (N_23203,N_19578,N_19765);
nand U23204 (N_23204,N_17391,N_17623);
nand U23205 (N_23205,N_16528,N_15815);
nor U23206 (N_23206,N_17780,N_17226);
nor U23207 (N_23207,N_17967,N_17626);
nand U23208 (N_23208,N_18535,N_18853);
xnor U23209 (N_23209,N_18214,N_19531);
nor U23210 (N_23210,N_16922,N_16539);
nor U23211 (N_23211,N_17225,N_15174);
and U23212 (N_23212,N_16969,N_16710);
nor U23213 (N_23213,N_15644,N_19870);
nor U23214 (N_23214,N_19822,N_17079);
or U23215 (N_23215,N_16189,N_18104);
nor U23216 (N_23216,N_16058,N_16989);
nand U23217 (N_23217,N_16456,N_19507);
nor U23218 (N_23218,N_16824,N_17068);
and U23219 (N_23219,N_18265,N_19686);
nand U23220 (N_23220,N_18799,N_17614);
xor U23221 (N_23221,N_15500,N_17223);
or U23222 (N_23222,N_15119,N_16415);
and U23223 (N_23223,N_19635,N_17259);
nand U23224 (N_23224,N_17429,N_16798);
xnor U23225 (N_23225,N_19867,N_19582);
nand U23226 (N_23226,N_19608,N_16775);
and U23227 (N_23227,N_15252,N_19527);
and U23228 (N_23228,N_17894,N_16858);
and U23229 (N_23229,N_19838,N_17412);
and U23230 (N_23230,N_17236,N_17192);
nand U23231 (N_23231,N_19364,N_19380);
or U23232 (N_23232,N_18273,N_18114);
nor U23233 (N_23233,N_19336,N_16036);
xnor U23234 (N_23234,N_18588,N_19610);
and U23235 (N_23235,N_16353,N_16680);
or U23236 (N_23236,N_17825,N_19874);
and U23237 (N_23237,N_16622,N_17576);
or U23238 (N_23238,N_18647,N_15832);
xor U23239 (N_23239,N_17783,N_19456);
or U23240 (N_23240,N_16732,N_17702);
nand U23241 (N_23241,N_18469,N_16731);
or U23242 (N_23242,N_15722,N_16314);
nand U23243 (N_23243,N_18306,N_19478);
or U23244 (N_23244,N_18343,N_18584);
and U23245 (N_23245,N_19763,N_16770);
xor U23246 (N_23246,N_16446,N_17091);
xor U23247 (N_23247,N_16236,N_16487);
nor U23248 (N_23248,N_17818,N_15285);
nor U23249 (N_23249,N_15087,N_19128);
or U23250 (N_23250,N_15561,N_15041);
nand U23251 (N_23251,N_17783,N_17344);
and U23252 (N_23252,N_19550,N_15800);
or U23253 (N_23253,N_19712,N_17049);
or U23254 (N_23254,N_19455,N_18440);
xnor U23255 (N_23255,N_17883,N_17897);
and U23256 (N_23256,N_18966,N_18743);
nand U23257 (N_23257,N_17485,N_15482);
nand U23258 (N_23258,N_17844,N_15903);
or U23259 (N_23259,N_17053,N_19997);
and U23260 (N_23260,N_19415,N_18847);
nor U23261 (N_23261,N_18045,N_15713);
nand U23262 (N_23262,N_16443,N_17778);
or U23263 (N_23263,N_15130,N_19744);
nand U23264 (N_23264,N_17842,N_15343);
nor U23265 (N_23265,N_16636,N_16734);
nand U23266 (N_23266,N_17921,N_17479);
and U23267 (N_23267,N_15599,N_15180);
nor U23268 (N_23268,N_18853,N_18116);
xnor U23269 (N_23269,N_16847,N_16349);
and U23270 (N_23270,N_17877,N_18609);
nand U23271 (N_23271,N_17885,N_18989);
nand U23272 (N_23272,N_18707,N_17075);
xor U23273 (N_23273,N_19253,N_19191);
and U23274 (N_23274,N_18149,N_17599);
or U23275 (N_23275,N_17836,N_19343);
and U23276 (N_23276,N_19115,N_18457);
nor U23277 (N_23277,N_16692,N_15928);
xnor U23278 (N_23278,N_15051,N_15326);
or U23279 (N_23279,N_17611,N_18699);
or U23280 (N_23280,N_18869,N_17745);
or U23281 (N_23281,N_15296,N_16538);
nand U23282 (N_23282,N_17508,N_18024);
nor U23283 (N_23283,N_17587,N_15294);
or U23284 (N_23284,N_17149,N_19977);
xnor U23285 (N_23285,N_16089,N_18621);
and U23286 (N_23286,N_15121,N_16129);
and U23287 (N_23287,N_15589,N_18232);
nor U23288 (N_23288,N_16287,N_18376);
xnor U23289 (N_23289,N_18506,N_17275);
or U23290 (N_23290,N_18283,N_16272);
nor U23291 (N_23291,N_16251,N_16744);
and U23292 (N_23292,N_18541,N_19320);
nand U23293 (N_23293,N_15202,N_16117);
xnor U23294 (N_23294,N_18146,N_19573);
xor U23295 (N_23295,N_15212,N_19475);
xor U23296 (N_23296,N_15329,N_16719);
or U23297 (N_23297,N_18230,N_15474);
nor U23298 (N_23298,N_19467,N_18166);
nand U23299 (N_23299,N_17405,N_17961);
nand U23300 (N_23300,N_18909,N_17663);
xnor U23301 (N_23301,N_19981,N_17793);
nor U23302 (N_23302,N_18103,N_15664);
or U23303 (N_23303,N_17840,N_18081);
nor U23304 (N_23304,N_15548,N_16965);
nor U23305 (N_23305,N_18559,N_18522);
or U23306 (N_23306,N_16489,N_16967);
xor U23307 (N_23307,N_16331,N_17292);
nand U23308 (N_23308,N_18605,N_18773);
xor U23309 (N_23309,N_15817,N_16138);
nor U23310 (N_23310,N_15131,N_18172);
or U23311 (N_23311,N_15697,N_19011);
and U23312 (N_23312,N_15932,N_15917);
and U23313 (N_23313,N_19752,N_16900);
xor U23314 (N_23314,N_17844,N_16983);
xnor U23315 (N_23315,N_15711,N_15438);
xor U23316 (N_23316,N_18609,N_19433);
or U23317 (N_23317,N_15507,N_18898);
and U23318 (N_23318,N_16389,N_15611);
nor U23319 (N_23319,N_19075,N_17718);
and U23320 (N_23320,N_18921,N_15707);
and U23321 (N_23321,N_18195,N_17414);
and U23322 (N_23322,N_15686,N_15138);
xor U23323 (N_23323,N_19909,N_18403);
or U23324 (N_23324,N_18307,N_19269);
or U23325 (N_23325,N_18349,N_19830);
or U23326 (N_23326,N_15849,N_18916);
nand U23327 (N_23327,N_18069,N_18131);
nand U23328 (N_23328,N_16507,N_19861);
and U23329 (N_23329,N_18322,N_19498);
nor U23330 (N_23330,N_16944,N_15785);
and U23331 (N_23331,N_15891,N_17957);
nor U23332 (N_23332,N_16382,N_15198);
xor U23333 (N_23333,N_16721,N_17838);
xnor U23334 (N_23334,N_19532,N_16429);
xnor U23335 (N_23335,N_19552,N_19868);
nand U23336 (N_23336,N_15334,N_15550);
xnor U23337 (N_23337,N_15958,N_17207);
or U23338 (N_23338,N_15183,N_19135);
xor U23339 (N_23339,N_18773,N_18158);
nor U23340 (N_23340,N_18371,N_18592);
or U23341 (N_23341,N_18668,N_15328);
or U23342 (N_23342,N_19110,N_16570);
or U23343 (N_23343,N_17771,N_19253);
nand U23344 (N_23344,N_15740,N_15776);
or U23345 (N_23345,N_17981,N_15650);
nor U23346 (N_23346,N_15364,N_17331);
nand U23347 (N_23347,N_19898,N_19185);
xnor U23348 (N_23348,N_18591,N_17679);
xor U23349 (N_23349,N_19063,N_19548);
xor U23350 (N_23350,N_18857,N_17628);
xnor U23351 (N_23351,N_19243,N_18082);
nand U23352 (N_23352,N_19947,N_17341);
nand U23353 (N_23353,N_15005,N_19122);
nand U23354 (N_23354,N_15074,N_19879);
or U23355 (N_23355,N_15146,N_18944);
or U23356 (N_23356,N_16739,N_15772);
nand U23357 (N_23357,N_19585,N_18464);
nor U23358 (N_23358,N_16457,N_15613);
and U23359 (N_23359,N_16708,N_19302);
xor U23360 (N_23360,N_16683,N_19589);
xnor U23361 (N_23361,N_15284,N_16653);
xor U23362 (N_23362,N_18234,N_17604);
nand U23363 (N_23363,N_15887,N_19093);
nand U23364 (N_23364,N_18691,N_19019);
nand U23365 (N_23365,N_16628,N_17680);
nor U23366 (N_23366,N_19380,N_19566);
and U23367 (N_23367,N_18674,N_19781);
nand U23368 (N_23368,N_15821,N_18725);
and U23369 (N_23369,N_15486,N_18244);
nor U23370 (N_23370,N_17707,N_19408);
nand U23371 (N_23371,N_17196,N_16963);
nor U23372 (N_23372,N_15239,N_18848);
nor U23373 (N_23373,N_17403,N_18132);
or U23374 (N_23374,N_15121,N_15663);
nand U23375 (N_23375,N_16424,N_16390);
nor U23376 (N_23376,N_15552,N_18161);
xnor U23377 (N_23377,N_18155,N_19197);
nand U23378 (N_23378,N_16796,N_17574);
nor U23379 (N_23379,N_17907,N_17352);
or U23380 (N_23380,N_19992,N_17993);
nand U23381 (N_23381,N_15616,N_16748);
and U23382 (N_23382,N_19972,N_16639);
nor U23383 (N_23383,N_18987,N_17335);
xnor U23384 (N_23384,N_19246,N_15172);
nor U23385 (N_23385,N_15000,N_17676);
xnor U23386 (N_23386,N_17581,N_19817);
xor U23387 (N_23387,N_19978,N_19755);
xor U23388 (N_23388,N_19036,N_18549);
xnor U23389 (N_23389,N_19019,N_18911);
xor U23390 (N_23390,N_19126,N_16494);
and U23391 (N_23391,N_18459,N_16142);
nor U23392 (N_23392,N_18361,N_19992);
xnor U23393 (N_23393,N_15360,N_15451);
or U23394 (N_23394,N_15069,N_16136);
nand U23395 (N_23395,N_18665,N_18732);
and U23396 (N_23396,N_15338,N_17386);
or U23397 (N_23397,N_18698,N_18126);
and U23398 (N_23398,N_19144,N_17067);
or U23399 (N_23399,N_19652,N_16769);
and U23400 (N_23400,N_16660,N_18162);
or U23401 (N_23401,N_16964,N_16335);
and U23402 (N_23402,N_18741,N_19497);
nand U23403 (N_23403,N_17154,N_15188);
xor U23404 (N_23404,N_15993,N_15559);
or U23405 (N_23405,N_16104,N_16937);
xnor U23406 (N_23406,N_15823,N_15142);
xor U23407 (N_23407,N_19173,N_18706);
nand U23408 (N_23408,N_17565,N_15781);
nor U23409 (N_23409,N_16196,N_15099);
nand U23410 (N_23410,N_16001,N_16384);
nor U23411 (N_23411,N_16107,N_17026);
and U23412 (N_23412,N_17996,N_16890);
or U23413 (N_23413,N_19115,N_18110);
nor U23414 (N_23414,N_19875,N_16835);
xor U23415 (N_23415,N_17955,N_16133);
or U23416 (N_23416,N_16034,N_19231);
xor U23417 (N_23417,N_18452,N_18819);
nand U23418 (N_23418,N_16159,N_18608);
and U23419 (N_23419,N_16976,N_15390);
xnor U23420 (N_23420,N_19883,N_16064);
xnor U23421 (N_23421,N_18373,N_15456);
or U23422 (N_23422,N_15427,N_19655);
xor U23423 (N_23423,N_15925,N_17672);
or U23424 (N_23424,N_19808,N_18830);
xnor U23425 (N_23425,N_19552,N_19852);
nor U23426 (N_23426,N_16751,N_17726);
nand U23427 (N_23427,N_15417,N_18757);
nor U23428 (N_23428,N_17620,N_18499);
or U23429 (N_23429,N_19791,N_18021);
and U23430 (N_23430,N_15149,N_19192);
nor U23431 (N_23431,N_18918,N_15897);
nor U23432 (N_23432,N_16020,N_16677);
and U23433 (N_23433,N_19527,N_19178);
nor U23434 (N_23434,N_15955,N_17932);
xnor U23435 (N_23435,N_19964,N_15944);
xor U23436 (N_23436,N_17363,N_17601);
xnor U23437 (N_23437,N_18092,N_16414);
and U23438 (N_23438,N_18682,N_15142);
and U23439 (N_23439,N_17035,N_19980);
nand U23440 (N_23440,N_18222,N_15993);
or U23441 (N_23441,N_19063,N_19359);
nor U23442 (N_23442,N_17601,N_17595);
nand U23443 (N_23443,N_19703,N_17660);
xor U23444 (N_23444,N_15368,N_17161);
nand U23445 (N_23445,N_17099,N_16629);
nor U23446 (N_23446,N_18803,N_16064);
xor U23447 (N_23447,N_15394,N_17039);
xnor U23448 (N_23448,N_17454,N_16443);
or U23449 (N_23449,N_19239,N_19773);
nor U23450 (N_23450,N_19184,N_16141);
nor U23451 (N_23451,N_18389,N_18941);
nand U23452 (N_23452,N_19458,N_18036);
xor U23453 (N_23453,N_19810,N_15976);
or U23454 (N_23454,N_16232,N_16615);
nor U23455 (N_23455,N_15697,N_15906);
nand U23456 (N_23456,N_16471,N_17682);
nor U23457 (N_23457,N_17534,N_17973);
xor U23458 (N_23458,N_18889,N_18936);
nor U23459 (N_23459,N_16166,N_18766);
xnor U23460 (N_23460,N_15039,N_15887);
xnor U23461 (N_23461,N_19561,N_18480);
xor U23462 (N_23462,N_19877,N_17544);
nor U23463 (N_23463,N_16638,N_17998);
and U23464 (N_23464,N_16028,N_18471);
or U23465 (N_23465,N_17255,N_17757);
nand U23466 (N_23466,N_15534,N_17118);
and U23467 (N_23467,N_17004,N_15939);
or U23468 (N_23468,N_15941,N_16909);
xnor U23469 (N_23469,N_16884,N_17629);
or U23470 (N_23470,N_15442,N_18226);
nand U23471 (N_23471,N_19991,N_18590);
xnor U23472 (N_23472,N_15962,N_17737);
xnor U23473 (N_23473,N_15748,N_19773);
nand U23474 (N_23474,N_16214,N_17688);
xor U23475 (N_23475,N_15503,N_15239);
xnor U23476 (N_23476,N_17117,N_15510);
nand U23477 (N_23477,N_16381,N_18939);
or U23478 (N_23478,N_18034,N_19331);
and U23479 (N_23479,N_19861,N_15181);
nand U23480 (N_23480,N_18843,N_15506);
nor U23481 (N_23481,N_17342,N_18197);
xnor U23482 (N_23482,N_19690,N_17031);
nor U23483 (N_23483,N_18434,N_18786);
and U23484 (N_23484,N_15894,N_18079);
xor U23485 (N_23485,N_16326,N_15967);
nor U23486 (N_23486,N_18736,N_18387);
nor U23487 (N_23487,N_18823,N_16658);
nor U23488 (N_23488,N_17536,N_19111);
or U23489 (N_23489,N_18405,N_15685);
nor U23490 (N_23490,N_16248,N_18911);
nand U23491 (N_23491,N_15667,N_17881);
or U23492 (N_23492,N_18839,N_19610);
or U23493 (N_23493,N_19406,N_16503);
and U23494 (N_23494,N_19262,N_15002);
xnor U23495 (N_23495,N_18451,N_18764);
xor U23496 (N_23496,N_19172,N_18273);
or U23497 (N_23497,N_18291,N_18504);
xor U23498 (N_23498,N_17294,N_19679);
or U23499 (N_23499,N_19493,N_15289);
and U23500 (N_23500,N_15478,N_19522);
xor U23501 (N_23501,N_18886,N_19376);
nand U23502 (N_23502,N_15183,N_19822);
nor U23503 (N_23503,N_15176,N_19314);
or U23504 (N_23504,N_18867,N_15279);
or U23505 (N_23505,N_17026,N_18466);
or U23506 (N_23506,N_18203,N_17297);
xnor U23507 (N_23507,N_19335,N_15225);
and U23508 (N_23508,N_15045,N_19799);
or U23509 (N_23509,N_17360,N_16603);
xor U23510 (N_23510,N_15045,N_18452);
xnor U23511 (N_23511,N_15038,N_18824);
nor U23512 (N_23512,N_15367,N_16192);
nand U23513 (N_23513,N_19891,N_16252);
and U23514 (N_23514,N_15822,N_17098);
nor U23515 (N_23515,N_19016,N_19202);
or U23516 (N_23516,N_18011,N_17277);
and U23517 (N_23517,N_17896,N_19250);
xor U23518 (N_23518,N_15180,N_19017);
xnor U23519 (N_23519,N_17284,N_19380);
and U23520 (N_23520,N_17274,N_19292);
or U23521 (N_23521,N_16562,N_17669);
nor U23522 (N_23522,N_18428,N_16593);
xor U23523 (N_23523,N_15891,N_19801);
and U23524 (N_23524,N_15413,N_16317);
and U23525 (N_23525,N_15245,N_17169);
nand U23526 (N_23526,N_19759,N_16811);
nor U23527 (N_23527,N_18890,N_15133);
or U23528 (N_23528,N_16711,N_17535);
nor U23529 (N_23529,N_15244,N_18817);
or U23530 (N_23530,N_19424,N_18733);
or U23531 (N_23531,N_16617,N_16718);
nand U23532 (N_23532,N_17947,N_18846);
and U23533 (N_23533,N_15320,N_18997);
or U23534 (N_23534,N_17294,N_15707);
nand U23535 (N_23535,N_17167,N_15426);
nor U23536 (N_23536,N_16589,N_15920);
and U23537 (N_23537,N_18691,N_19292);
nor U23538 (N_23538,N_16804,N_15864);
nor U23539 (N_23539,N_18417,N_19066);
nand U23540 (N_23540,N_18789,N_15494);
or U23541 (N_23541,N_15306,N_18768);
xor U23542 (N_23542,N_17948,N_15006);
xor U23543 (N_23543,N_16081,N_18648);
nand U23544 (N_23544,N_18985,N_19448);
nand U23545 (N_23545,N_15458,N_18106);
xor U23546 (N_23546,N_19327,N_17415);
and U23547 (N_23547,N_17619,N_19170);
or U23548 (N_23548,N_17364,N_18770);
nor U23549 (N_23549,N_15234,N_16075);
or U23550 (N_23550,N_16596,N_17799);
or U23551 (N_23551,N_19094,N_15685);
nand U23552 (N_23552,N_18415,N_15203);
nor U23553 (N_23553,N_15657,N_16134);
and U23554 (N_23554,N_19631,N_15070);
nand U23555 (N_23555,N_15483,N_19083);
and U23556 (N_23556,N_16477,N_17027);
xor U23557 (N_23557,N_16722,N_15492);
nor U23558 (N_23558,N_16013,N_19991);
xor U23559 (N_23559,N_16960,N_15988);
xnor U23560 (N_23560,N_15312,N_19091);
xnor U23561 (N_23561,N_17673,N_18823);
nor U23562 (N_23562,N_19486,N_17812);
and U23563 (N_23563,N_18909,N_17293);
or U23564 (N_23564,N_15959,N_18777);
nor U23565 (N_23565,N_17126,N_19738);
or U23566 (N_23566,N_19990,N_19669);
and U23567 (N_23567,N_15313,N_18279);
or U23568 (N_23568,N_17668,N_17429);
nor U23569 (N_23569,N_19868,N_16539);
nand U23570 (N_23570,N_17410,N_19408);
xnor U23571 (N_23571,N_19777,N_19593);
or U23572 (N_23572,N_15677,N_16043);
nand U23573 (N_23573,N_18896,N_18201);
nor U23574 (N_23574,N_18596,N_15577);
nand U23575 (N_23575,N_18536,N_16682);
and U23576 (N_23576,N_17371,N_18612);
or U23577 (N_23577,N_19661,N_15404);
nand U23578 (N_23578,N_15566,N_17357);
or U23579 (N_23579,N_18901,N_17476);
nand U23580 (N_23580,N_15783,N_19578);
or U23581 (N_23581,N_17817,N_18731);
nor U23582 (N_23582,N_15060,N_19471);
nand U23583 (N_23583,N_19392,N_16741);
nand U23584 (N_23584,N_16256,N_18891);
nand U23585 (N_23585,N_19846,N_17951);
and U23586 (N_23586,N_16994,N_16441);
nor U23587 (N_23587,N_19962,N_19222);
and U23588 (N_23588,N_18331,N_16439);
xor U23589 (N_23589,N_15541,N_16802);
and U23590 (N_23590,N_19339,N_16090);
or U23591 (N_23591,N_15999,N_15829);
and U23592 (N_23592,N_16998,N_15129);
xnor U23593 (N_23593,N_16354,N_19815);
and U23594 (N_23594,N_19180,N_15468);
xor U23595 (N_23595,N_17405,N_16288);
nand U23596 (N_23596,N_19781,N_18696);
or U23597 (N_23597,N_17462,N_15254);
and U23598 (N_23598,N_18683,N_18075);
or U23599 (N_23599,N_18581,N_18265);
xor U23600 (N_23600,N_19930,N_17818);
nand U23601 (N_23601,N_16818,N_15953);
nand U23602 (N_23602,N_17886,N_16245);
nor U23603 (N_23603,N_17545,N_19892);
or U23604 (N_23604,N_15784,N_19422);
xor U23605 (N_23605,N_17093,N_19138);
xor U23606 (N_23606,N_19953,N_15185);
or U23607 (N_23607,N_17557,N_18334);
nand U23608 (N_23608,N_17183,N_19697);
or U23609 (N_23609,N_17292,N_19286);
nor U23610 (N_23610,N_15206,N_16210);
or U23611 (N_23611,N_16167,N_17843);
nor U23612 (N_23612,N_17312,N_16010);
nor U23613 (N_23613,N_18792,N_16333);
nand U23614 (N_23614,N_16922,N_16742);
and U23615 (N_23615,N_16216,N_18209);
nor U23616 (N_23616,N_15345,N_15681);
and U23617 (N_23617,N_16241,N_16874);
nand U23618 (N_23618,N_17913,N_19293);
xnor U23619 (N_23619,N_16273,N_18613);
or U23620 (N_23620,N_16327,N_16371);
xnor U23621 (N_23621,N_18758,N_16251);
or U23622 (N_23622,N_17017,N_16073);
or U23623 (N_23623,N_18706,N_17903);
nand U23624 (N_23624,N_18926,N_17263);
and U23625 (N_23625,N_16545,N_15280);
or U23626 (N_23626,N_17736,N_19388);
nand U23627 (N_23627,N_19969,N_17817);
nor U23628 (N_23628,N_16843,N_17555);
and U23629 (N_23629,N_19928,N_19803);
nor U23630 (N_23630,N_19437,N_16514);
nand U23631 (N_23631,N_15465,N_15248);
nand U23632 (N_23632,N_18533,N_18774);
or U23633 (N_23633,N_16070,N_19357);
and U23634 (N_23634,N_19774,N_15101);
or U23635 (N_23635,N_19978,N_18671);
nor U23636 (N_23636,N_16551,N_19057);
xor U23637 (N_23637,N_17330,N_19144);
nor U23638 (N_23638,N_17034,N_19610);
or U23639 (N_23639,N_15072,N_19713);
nand U23640 (N_23640,N_19532,N_18344);
nand U23641 (N_23641,N_19375,N_15346);
nand U23642 (N_23642,N_19724,N_15926);
nand U23643 (N_23643,N_17659,N_19687);
and U23644 (N_23644,N_16428,N_15734);
nand U23645 (N_23645,N_19218,N_17958);
and U23646 (N_23646,N_16881,N_16403);
and U23647 (N_23647,N_17770,N_19229);
xor U23648 (N_23648,N_15791,N_15493);
xnor U23649 (N_23649,N_19424,N_17994);
nor U23650 (N_23650,N_18190,N_15479);
nand U23651 (N_23651,N_19886,N_17434);
or U23652 (N_23652,N_17582,N_18101);
xor U23653 (N_23653,N_15658,N_19579);
nand U23654 (N_23654,N_16261,N_16351);
nor U23655 (N_23655,N_16722,N_15940);
xor U23656 (N_23656,N_15735,N_17778);
xnor U23657 (N_23657,N_18714,N_15674);
nand U23658 (N_23658,N_17046,N_17028);
nand U23659 (N_23659,N_16596,N_16104);
nand U23660 (N_23660,N_19794,N_19070);
nor U23661 (N_23661,N_18221,N_17735);
and U23662 (N_23662,N_15874,N_19926);
xnor U23663 (N_23663,N_17064,N_19420);
nand U23664 (N_23664,N_19762,N_17709);
or U23665 (N_23665,N_17129,N_19390);
or U23666 (N_23666,N_18644,N_17315);
nand U23667 (N_23667,N_15384,N_19115);
nand U23668 (N_23668,N_18957,N_19783);
xnor U23669 (N_23669,N_19490,N_18439);
nand U23670 (N_23670,N_17608,N_16370);
and U23671 (N_23671,N_16297,N_16247);
nand U23672 (N_23672,N_19407,N_18405);
nand U23673 (N_23673,N_19302,N_15611);
nand U23674 (N_23674,N_19843,N_15597);
or U23675 (N_23675,N_16083,N_18122);
and U23676 (N_23676,N_18990,N_15432);
nand U23677 (N_23677,N_15224,N_15913);
and U23678 (N_23678,N_17032,N_17669);
nand U23679 (N_23679,N_16435,N_17138);
and U23680 (N_23680,N_18005,N_19107);
or U23681 (N_23681,N_19132,N_15034);
nand U23682 (N_23682,N_17117,N_15364);
or U23683 (N_23683,N_18406,N_15968);
or U23684 (N_23684,N_18335,N_18894);
nand U23685 (N_23685,N_16786,N_16970);
or U23686 (N_23686,N_16492,N_17368);
and U23687 (N_23687,N_15304,N_16719);
and U23688 (N_23688,N_18494,N_16208);
nor U23689 (N_23689,N_15425,N_16916);
nand U23690 (N_23690,N_15512,N_18342);
nand U23691 (N_23691,N_15341,N_18213);
and U23692 (N_23692,N_16991,N_15671);
and U23693 (N_23693,N_15873,N_17887);
xnor U23694 (N_23694,N_17425,N_19769);
or U23695 (N_23695,N_18534,N_17066);
nor U23696 (N_23696,N_18585,N_19153);
and U23697 (N_23697,N_15598,N_15002);
or U23698 (N_23698,N_15792,N_16129);
and U23699 (N_23699,N_17038,N_16455);
nand U23700 (N_23700,N_18930,N_17357);
nand U23701 (N_23701,N_16815,N_19191);
nand U23702 (N_23702,N_18372,N_16359);
xor U23703 (N_23703,N_15330,N_18172);
xor U23704 (N_23704,N_19337,N_17141);
nor U23705 (N_23705,N_17368,N_16844);
or U23706 (N_23706,N_15117,N_15743);
nor U23707 (N_23707,N_18980,N_17623);
nor U23708 (N_23708,N_15075,N_17261);
nand U23709 (N_23709,N_18363,N_17130);
or U23710 (N_23710,N_19119,N_19685);
xor U23711 (N_23711,N_15045,N_15537);
xor U23712 (N_23712,N_16189,N_16035);
or U23713 (N_23713,N_15049,N_18257);
or U23714 (N_23714,N_19956,N_18110);
nor U23715 (N_23715,N_19018,N_17727);
xnor U23716 (N_23716,N_15037,N_17825);
xor U23717 (N_23717,N_15306,N_19924);
and U23718 (N_23718,N_16345,N_19663);
and U23719 (N_23719,N_17093,N_19117);
and U23720 (N_23720,N_16337,N_16542);
xnor U23721 (N_23721,N_15900,N_16840);
or U23722 (N_23722,N_19036,N_17571);
nor U23723 (N_23723,N_16039,N_19432);
nand U23724 (N_23724,N_15598,N_17086);
nand U23725 (N_23725,N_17885,N_18305);
and U23726 (N_23726,N_15502,N_19815);
nand U23727 (N_23727,N_16886,N_19105);
nand U23728 (N_23728,N_19540,N_18002);
or U23729 (N_23729,N_19081,N_15587);
xnor U23730 (N_23730,N_15737,N_19677);
nand U23731 (N_23731,N_17099,N_18065);
xor U23732 (N_23732,N_19169,N_17650);
xnor U23733 (N_23733,N_19469,N_18069);
nand U23734 (N_23734,N_16488,N_15296);
nor U23735 (N_23735,N_18384,N_17853);
nor U23736 (N_23736,N_16238,N_19768);
nand U23737 (N_23737,N_19339,N_18266);
and U23738 (N_23738,N_19261,N_17996);
or U23739 (N_23739,N_16034,N_18685);
xor U23740 (N_23740,N_17096,N_19349);
xor U23741 (N_23741,N_19111,N_18836);
or U23742 (N_23742,N_18938,N_16370);
or U23743 (N_23743,N_18345,N_17220);
or U23744 (N_23744,N_17105,N_16970);
nor U23745 (N_23745,N_15882,N_17818);
or U23746 (N_23746,N_16779,N_18941);
nor U23747 (N_23747,N_16458,N_15129);
or U23748 (N_23748,N_15483,N_17046);
nand U23749 (N_23749,N_17775,N_17617);
nand U23750 (N_23750,N_16954,N_18139);
and U23751 (N_23751,N_18695,N_15437);
nor U23752 (N_23752,N_18118,N_17383);
nor U23753 (N_23753,N_17467,N_16517);
nand U23754 (N_23754,N_15626,N_19956);
xor U23755 (N_23755,N_17962,N_18102);
xnor U23756 (N_23756,N_17760,N_15342);
nand U23757 (N_23757,N_18785,N_15879);
and U23758 (N_23758,N_17395,N_18926);
or U23759 (N_23759,N_15637,N_15325);
xnor U23760 (N_23760,N_18800,N_15546);
and U23761 (N_23761,N_17067,N_16180);
or U23762 (N_23762,N_15318,N_16083);
xnor U23763 (N_23763,N_19681,N_15223);
nand U23764 (N_23764,N_19363,N_15719);
or U23765 (N_23765,N_17844,N_16805);
nand U23766 (N_23766,N_19523,N_18947);
xor U23767 (N_23767,N_16213,N_16112);
nor U23768 (N_23768,N_18011,N_16650);
or U23769 (N_23769,N_19684,N_16860);
xnor U23770 (N_23770,N_16650,N_16544);
and U23771 (N_23771,N_19524,N_17747);
nor U23772 (N_23772,N_18059,N_16095);
nor U23773 (N_23773,N_18533,N_18307);
nand U23774 (N_23774,N_16629,N_15549);
xor U23775 (N_23775,N_17180,N_17541);
nand U23776 (N_23776,N_15710,N_17124);
nand U23777 (N_23777,N_15111,N_19229);
nor U23778 (N_23778,N_18982,N_16234);
nand U23779 (N_23779,N_18337,N_17175);
xnor U23780 (N_23780,N_19912,N_15666);
nand U23781 (N_23781,N_15516,N_19990);
nor U23782 (N_23782,N_19658,N_15582);
xnor U23783 (N_23783,N_16154,N_15202);
and U23784 (N_23784,N_18624,N_19949);
nand U23785 (N_23785,N_16511,N_16252);
xor U23786 (N_23786,N_17375,N_16706);
nand U23787 (N_23787,N_19280,N_15740);
xnor U23788 (N_23788,N_18744,N_19910);
nor U23789 (N_23789,N_17970,N_16820);
xnor U23790 (N_23790,N_15298,N_18873);
nor U23791 (N_23791,N_16691,N_16034);
nor U23792 (N_23792,N_15101,N_17931);
nor U23793 (N_23793,N_17250,N_18225);
and U23794 (N_23794,N_17596,N_19495);
xnor U23795 (N_23795,N_16587,N_19899);
xnor U23796 (N_23796,N_17332,N_19859);
nor U23797 (N_23797,N_19657,N_17835);
xnor U23798 (N_23798,N_16639,N_19102);
nand U23799 (N_23799,N_18076,N_17201);
nand U23800 (N_23800,N_17830,N_15828);
or U23801 (N_23801,N_18382,N_16185);
nand U23802 (N_23802,N_19877,N_18503);
nand U23803 (N_23803,N_19616,N_16038);
nor U23804 (N_23804,N_17341,N_19776);
xor U23805 (N_23805,N_15794,N_16276);
nor U23806 (N_23806,N_17265,N_18549);
and U23807 (N_23807,N_15911,N_17516);
nand U23808 (N_23808,N_19202,N_16089);
xor U23809 (N_23809,N_18029,N_16122);
or U23810 (N_23810,N_17606,N_15079);
nand U23811 (N_23811,N_16629,N_19202);
or U23812 (N_23812,N_19673,N_16242);
nor U23813 (N_23813,N_15645,N_17997);
nor U23814 (N_23814,N_19678,N_16382);
or U23815 (N_23815,N_18858,N_19973);
nand U23816 (N_23816,N_17016,N_16639);
xor U23817 (N_23817,N_17645,N_16204);
nand U23818 (N_23818,N_18087,N_19005);
nor U23819 (N_23819,N_19377,N_19794);
and U23820 (N_23820,N_15289,N_17667);
xor U23821 (N_23821,N_16598,N_19220);
and U23822 (N_23822,N_16194,N_17721);
nand U23823 (N_23823,N_19039,N_16345);
or U23824 (N_23824,N_17443,N_15829);
nor U23825 (N_23825,N_19144,N_19657);
xnor U23826 (N_23826,N_17390,N_19868);
nand U23827 (N_23827,N_17639,N_19788);
and U23828 (N_23828,N_16894,N_18207);
nand U23829 (N_23829,N_17953,N_16787);
and U23830 (N_23830,N_18075,N_18858);
nand U23831 (N_23831,N_15582,N_16889);
or U23832 (N_23832,N_16049,N_18081);
xnor U23833 (N_23833,N_18349,N_18782);
xor U23834 (N_23834,N_19339,N_19939);
nand U23835 (N_23835,N_15639,N_15265);
and U23836 (N_23836,N_15211,N_18490);
and U23837 (N_23837,N_16477,N_16977);
xnor U23838 (N_23838,N_17481,N_17850);
nand U23839 (N_23839,N_18633,N_16355);
nor U23840 (N_23840,N_17479,N_16984);
or U23841 (N_23841,N_17031,N_18283);
nor U23842 (N_23842,N_19689,N_19234);
nand U23843 (N_23843,N_18744,N_19233);
or U23844 (N_23844,N_16930,N_18560);
and U23845 (N_23845,N_16378,N_16331);
and U23846 (N_23846,N_15961,N_15204);
xor U23847 (N_23847,N_19927,N_16449);
xnor U23848 (N_23848,N_16592,N_15480);
nor U23849 (N_23849,N_15210,N_19491);
xor U23850 (N_23850,N_17448,N_15034);
nor U23851 (N_23851,N_18714,N_15221);
xor U23852 (N_23852,N_18476,N_15572);
and U23853 (N_23853,N_16091,N_15224);
xor U23854 (N_23854,N_15455,N_15512);
or U23855 (N_23855,N_17407,N_17063);
and U23856 (N_23856,N_15075,N_15968);
or U23857 (N_23857,N_17797,N_17235);
nor U23858 (N_23858,N_19622,N_17920);
and U23859 (N_23859,N_15232,N_17905);
or U23860 (N_23860,N_19800,N_17272);
or U23861 (N_23861,N_16795,N_15676);
nand U23862 (N_23862,N_18432,N_17547);
nor U23863 (N_23863,N_17107,N_16999);
nand U23864 (N_23864,N_16179,N_15911);
xnor U23865 (N_23865,N_16763,N_17768);
xor U23866 (N_23866,N_18820,N_15176);
nand U23867 (N_23867,N_15441,N_16518);
and U23868 (N_23868,N_19853,N_17312);
or U23869 (N_23869,N_15068,N_17208);
and U23870 (N_23870,N_17087,N_19321);
nor U23871 (N_23871,N_16415,N_15576);
or U23872 (N_23872,N_16782,N_17996);
xnor U23873 (N_23873,N_16350,N_18661);
nor U23874 (N_23874,N_16089,N_18947);
nor U23875 (N_23875,N_19148,N_15518);
nor U23876 (N_23876,N_17984,N_15432);
or U23877 (N_23877,N_15926,N_16401);
xnor U23878 (N_23878,N_18383,N_15648);
xnor U23879 (N_23879,N_16893,N_19278);
or U23880 (N_23880,N_16717,N_18631);
nor U23881 (N_23881,N_19580,N_19717);
nor U23882 (N_23882,N_17512,N_18599);
and U23883 (N_23883,N_17917,N_17876);
xor U23884 (N_23884,N_16296,N_17161);
xor U23885 (N_23885,N_15924,N_15312);
and U23886 (N_23886,N_17862,N_16252);
and U23887 (N_23887,N_17822,N_15835);
nand U23888 (N_23888,N_18016,N_18720);
and U23889 (N_23889,N_18487,N_17883);
xor U23890 (N_23890,N_17942,N_15792);
or U23891 (N_23891,N_17237,N_17101);
nor U23892 (N_23892,N_18054,N_19607);
nand U23893 (N_23893,N_18610,N_15645);
or U23894 (N_23894,N_19139,N_15223);
xnor U23895 (N_23895,N_17042,N_16335);
and U23896 (N_23896,N_18249,N_16147);
or U23897 (N_23897,N_18056,N_19728);
nand U23898 (N_23898,N_19125,N_19407);
nand U23899 (N_23899,N_18278,N_16836);
nor U23900 (N_23900,N_17366,N_18466);
xor U23901 (N_23901,N_17259,N_16752);
nor U23902 (N_23902,N_18803,N_19998);
xor U23903 (N_23903,N_19626,N_18770);
nor U23904 (N_23904,N_15107,N_16811);
and U23905 (N_23905,N_18187,N_16828);
or U23906 (N_23906,N_19144,N_18540);
xnor U23907 (N_23907,N_15253,N_16683);
nor U23908 (N_23908,N_19531,N_19696);
nand U23909 (N_23909,N_15282,N_19316);
and U23910 (N_23910,N_18795,N_16421);
or U23911 (N_23911,N_17850,N_16296);
nand U23912 (N_23912,N_19303,N_15203);
nand U23913 (N_23913,N_18757,N_18765);
or U23914 (N_23914,N_15802,N_17907);
xor U23915 (N_23915,N_15892,N_17899);
and U23916 (N_23916,N_15800,N_18863);
or U23917 (N_23917,N_16299,N_17479);
xnor U23918 (N_23918,N_16144,N_19846);
nand U23919 (N_23919,N_18786,N_18005);
and U23920 (N_23920,N_18075,N_19138);
nor U23921 (N_23921,N_19112,N_15184);
and U23922 (N_23922,N_15884,N_17536);
nand U23923 (N_23923,N_18170,N_17217);
nor U23924 (N_23924,N_19084,N_16693);
nand U23925 (N_23925,N_15952,N_15402);
xnor U23926 (N_23926,N_19547,N_16521);
xor U23927 (N_23927,N_16457,N_18606);
and U23928 (N_23928,N_18692,N_17397);
and U23929 (N_23929,N_15680,N_18195);
and U23930 (N_23930,N_16393,N_19614);
nor U23931 (N_23931,N_19010,N_18477);
xnor U23932 (N_23932,N_18725,N_17107);
xor U23933 (N_23933,N_19968,N_16839);
or U23934 (N_23934,N_15266,N_19150);
and U23935 (N_23935,N_17480,N_18815);
or U23936 (N_23936,N_16119,N_19277);
nor U23937 (N_23937,N_19857,N_17479);
nor U23938 (N_23938,N_17856,N_19410);
nor U23939 (N_23939,N_18269,N_18512);
nor U23940 (N_23940,N_15346,N_17739);
nor U23941 (N_23941,N_15015,N_16888);
nor U23942 (N_23942,N_19927,N_19354);
xor U23943 (N_23943,N_15824,N_16116);
nor U23944 (N_23944,N_18808,N_19295);
nand U23945 (N_23945,N_18127,N_16435);
and U23946 (N_23946,N_17274,N_16669);
xnor U23947 (N_23947,N_17905,N_15081);
xor U23948 (N_23948,N_19013,N_17332);
xnor U23949 (N_23949,N_18533,N_16916);
nand U23950 (N_23950,N_16801,N_19068);
nand U23951 (N_23951,N_18623,N_15820);
nor U23952 (N_23952,N_18894,N_18836);
or U23953 (N_23953,N_15652,N_15496);
or U23954 (N_23954,N_15696,N_18383);
or U23955 (N_23955,N_19311,N_17921);
nand U23956 (N_23956,N_18580,N_16993);
or U23957 (N_23957,N_18408,N_16764);
xnor U23958 (N_23958,N_19373,N_15409);
or U23959 (N_23959,N_15168,N_19718);
or U23960 (N_23960,N_15590,N_16217);
nand U23961 (N_23961,N_17293,N_15942);
nor U23962 (N_23962,N_16057,N_18407);
and U23963 (N_23963,N_19610,N_18960);
nor U23964 (N_23964,N_15937,N_18572);
nand U23965 (N_23965,N_16913,N_17453);
nor U23966 (N_23966,N_17899,N_17035);
and U23967 (N_23967,N_18583,N_18384);
or U23968 (N_23968,N_15739,N_16405);
or U23969 (N_23969,N_18029,N_19385);
or U23970 (N_23970,N_17782,N_18584);
xor U23971 (N_23971,N_15025,N_18074);
or U23972 (N_23972,N_16899,N_16498);
and U23973 (N_23973,N_16086,N_18738);
nand U23974 (N_23974,N_19670,N_19145);
or U23975 (N_23975,N_19620,N_17285);
nor U23976 (N_23976,N_18748,N_15371);
xor U23977 (N_23977,N_16522,N_17544);
xor U23978 (N_23978,N_18499,N_16034);
xor U23979 (N_23979,N_17923,N_17021);
xnor U23980 (N_23980,N_18749,N_18378);
nor U23981 (N_23981,N_16298,N_16486);
nand U23982 (N_23982,N_17522,N_17258);
xnor U23983 (N_23983,N_18397,N_16220);
nor U23984 (N_23984,N_16592,N_18884);
nor U23985 (N_23985,N_17715,N_17961);
nor U23986 (N_23986,N_19279,N_18771);
nor U23987 (N_23987,N_16921,N_16316);
xor U23988 (N_23988,N_17103,N_19644);
or U23989 (N_23989,N_15039,N_15182);
and U23990 (N_23990,N_18713,N_18553);
nor U23991 (N_23991,N_19506,N_17033);
nor U23992 (N_23992,N_17353,N_18536);
xnor U23993 (N_23993,N_18745,N_15180);
or U23994 (N_23994,N_15386,N_16597);
nor U23995 (N_23995,N_17218,N_16703);
or U23996 (N_23996,N_17948,N_17255);
nor U23997 (N_23997,N_15586,N_17411);
nand U23998 (N_23998,N_19127,N_18043);
or U23999 (N_23999,N_17802,N_15372);
nand U24000 (N_24000,N_16200,N_16493);
and U24001 (N_24001,N_18722,N_18312);
nor U24002 (N_24002,N_17759,N_17983);
nand U24003 (N_24003,N_19382,N_16974);
or U24004 (N_24004,N_16646,N_17595);
xor U24005 (N_24005,N_19182,N_15595);
nand U24006 (N_24006,N_17298,N_17919);
nor U24007 (N_24007,N_16707,N_15576);
nor U24008 (N_24008,N_16336,N_17774);
or U24009 (N_24009,N_16871,N_18874);
xnor U24010 (N_24010,N_16652,N_16626);
xnor U24011 (N_24011,N_19582,N_19329);
and U24012 (N_24012,N_18315,N_17078);
xnor U24013 (N_24013,N_18706,N_18242);
or U24014 (N_24014,N_19554,N_16244);
and U24015 (N_24015,N_17700,N_18445);
xnor U24016 (N_24016,N_17421,N_18543);
xnor U24017 (N_24017,N_15972,N_17031);
nand U24018 (N_24018,N_17446,N_16727);
nor U24019 (N_24019,N_16881,N_19009);
nand U24020 (N_24020,N_16775,N_16578);
nor U24021 (N_24021,N_17480,N_18645);
and U24022 (N_24022,N_15418,N_18563);
or U24023 (N_24023,N_18624,N_15290);
nor U24024 (N_24024,N_16456,N_18565);
xnor U24025 (N_24025,N_17979,N_17395);
nand U24026 (N_24026,N_19694,N_16998);
or U24027 (N_24027,N_17569,N_19070);
xnor U24028 (N_24028,N_18749,N_15997);
xor U24029 (N_24029,N_15565,N_15725);
or U24030 (N_24030,N_16466,N_19811);
and U24031 (N_24031,N_19154,N_18308);
nor U24032 (N_24032,N_18619,N_19476);
nand U24033 (N_24033,N_15144,N_18054);
nand U24034 (N_24034,N_15511,N_15789);
nor U24035 (N_24035,N_18768,N_15460);
or U24036 (N_24036,N_18644,N_17389);
or U24037 (N_24037,N_19058,N_15434);
xnor U24038 (N_24038,N_18908,N_18418);
or U24039 (N_24039,N_15157,N_18921);
nand U24040 (N_24040,N_19437,N_18691);
nand U24041 (N_24041,N_17679,N_18033);
nand U24042 (N_24042,N_17428,N_16722);
xnor U24043 (N_24043,N_19988,N_19285);
xor U24044 (N_24044,N_19391,N_16353);
nand U24045 (N_24045,N_19805,N_15676);
xor U24046 (N_24046,N_18428,N_18653);
and U24047 (N_24047,N_17658,N_18220);
nor U24048 (N_24048,N_17067,N_15533);
or U24049 (N_24049,N_16764,N_16400);
or U24050 (N_24050,N_16639,N_17958);
xnor U24051 (N_24051,N_16397,N_15439);
nor U24052 (N_24052,N_18987,N_15443);
nand U24053 (N_24053,N_19602,N_16970);
or U24054 (N_24054,N_18296,N_18123);
nand U24055 (N_24055,N_16795,N_16213);
or U24056 (N_24056,N_15297,N_16298);
xor U24057 (N_24057,N_17046,N_19819);
nand U24058 (N_24058,N_15312,N_17039);
xnor U24059 (N_24059,N_18506,N_16198);
nand U24060 (N_24060,N_18274,N_15078);
xnor U24061 (N_24061,N_19385,N_17725);
or U24062 (N_24062,N_18013,N_19719);
nand U24063 (N_24063,N_17591,N_15309);
nand U24064 (N_24064,N_15351,N_16328);
and U24065 (N_24065,N_17101,N_18730);
or U24066 (N_24066,N_19287,N_18021);
xnor U24067 (N_24067,N_17758,N_15903);
nand U24068 (N_24068,N_19592,N_19015);
xor U24069 (N_24069,N_15125,N_15523);
nor U24070 (N_24070,N_19061,N_15141);
nor U24071 (N_24071,N_18057,N_16674);
or U24072 (N_24072,N_16731,N_16676);
nor U24073 (N_24073,N_18282,N_17290);
xor U24074 (N_24074,N_16758,N_16731);
nor U24075 (N_24075,N_19376,N_15546);
and U24076 (N_24076,N_15091,N_15858);
and U24077 (N_24077,N_18490,N_18103);
and U24078 (N_24078,N_17500,N_18712);
or U24079 (N_24079,N_17154,N_17550);
and U24080 (N_24080,N_15858,N_16508);
nor U24081 (N_24081,N_19127,N_16132);
nor U24082 (N_24082,N_19245,N_18320);
nand U24083 (N_24083,N_15945,N_15192);
nor U24084 (N_24084,N_19649,N_17578);
and U24085 (N_24085,N_18876,N_19662);
and U24086 (N_24086,N_19901,N_17955);
xnor U24087 (N_24087,N_19137,N_18197);
or U24088 (N_24088,N_16221,N_18651);
or U24089 (N_24089,N_19855,N_15878);
or U24090 (N_24090,N_16954,N_18697);
and U24091 (N_24091,N_18291,N_17048);
and U24092 (N_24092,N_16900,N_17234);
nand U24093 (N_24093,N_16799,N_15751);
nand U24094 (N_24094,N_15851,N_18673);
and U24095 (N_24095,N_17670,N_18573);
xnor U24096 (N_24096,N_19069,N_16808);
xnor U24097 (N_24097,N_18090,N_16601);
or U24098 (N_24098,N_15057,N_19048);
nor U24099 (N_24099,N_15709,N_18391);
or U24100 (N_24100,N_19822,N_15475);
nand U24101 (N_24101,N_18874,N_16031);
or U24102 (N_24102,N_19352,N_17820);
xnor U24103 (N_24103,N_18748,N_15805);
or U24104 (N_24104,N_15941,N_19987);
xnor U24105 (N_24105,N_15764,N_16299);
and U24106 (N_24106,N_17790,N_15418);
and U24107 (N_24107,N_18640,N_18621);
xnor U24108 (N_24108,N_16238,N_15443);
and U24109 (N_24109,N_19013,N_16005);
and U24110 (N_24110,N_15844,N_16497);
xnor U24111 (N_24111,N_15527,N_17185);
nor U24112 (N_24112,N_15862,N_18835);
and U24113 (N_24113,N_15572,N_16395);
and U24114 (N_24114,N_17488,N_17828);
nor U24115 (N_24115,N_16266,N_16452);
nor U24116 (N_24116,N_16502,N_19334);
nand U24117 (N_24117,N_15414,N_17235);
and U24118 (N_24118,N_16857,N_18689);
nor U24119 (N_24119,N_15270,N_19545);
or U24120 (N_24120,N_16008,N_16592);
or U24121 (N_24121,N_16444,N_15696);
and U24122 (N_24122,N_17817,N_16728);
nor U24123 (N_24123,N_15252,N_16547);
and U24124 (N_24124,N_17818,N_17539);
or U24125 (N_24125,N_18972,N_15853);
xor U24126 (N_24126,N_19900,N_16342);
nand U24127 (N_24127,N_16389,N_16086);
nor U24128 (N_24128,N_16992,N_19993);
xnor U24129 (N_24129,N_17672,N_16696);
or U24130 (N_24130,N_19194,N_17237);
or U24131 (N_24131,N_16973,N_16449);
xor U24132 (N_24132,N_17147,N_18945);
nand U24133 (N_24133,N_17050,N_15036);
and U24134 (N_24134,N_18020,N_19986);
and U24135 (N_24135,N_16932,N_19934);
and U24136 (N_24136,N_17110,N_15205);
or U24137 (N_24137,N_18256,N_17916);
xor U24138 (N_24138,N_19777,N_18366);
nand U24139 (N_24139,N_15784,N_18041);
xnor U24140 (N_24140,N_16551,N_18802);
nand U24141 (N_24141,N_17394,N_18577);
nor U24142 (N_24142,N_15147,N_19106);
xnor U24143 (N_24143,N_16920,N_18401);
nand U24144 (N_24144,N_15062,N_16491);
nor U24145 (N_24145,N_16926,N_15015);
nor U24146 (N_24146,N_15443,N_15629);
or U24147 (N_24147,N_15329,N_18084);
and U24148 (N_24148,N_16288,N_15520);
or U24149 (N_24149,N_18848,N_18810);
xnor U24150 (N_24150,N_15415,N_19942);
nand U24151 (N_24151,N_16233,N_17669);
xor U24152 (N_24152,N_15617,N_19957);
or U24153 (N_24153,N_18072,N_15725);
or U24154 (N_24154,N_19668,N_19870);
and U24155 (N_24155,N_18683,N_19963);
nor U24156 (N_24156,N_19420,N_19346);
or U24157 (N_24157,N_15620,N_17556);
xnor U24158 (N_24158,N_16708,N_19091);
xnor U24159 (N_24159,N_16617,N_17159);
or U24160 (N_24160,N_16529,N_16742);
nand U24161 (N_24161,N_18731,N_18619);
and U24162 (N_24162,N_19683,N_19792);
or U24163 (N_24163,N_17672,N_19202);
nand U24164 (N_24164,N_19735,N_17113);
xor U24165 (N_24165,N_16016,N_18593);
xor U24166 (N_24166,N_15212,N_17198);
or U24167 (N_24167,N_16165,N_16109);
and U24168 (N_24168,N_15816,N_18618);
xor U24169 (N_24169,N_16753,N_19713);
xnor U24170 (N_24170,N_15968,N_18215);
and U24171 (N_24171,N_15508,N_17441);
xnor U24172 (N_24172,N_19356,N_16380);
or U24173 (N_24173,N_18882,N_18812);
nand U24174 (N_24174,N_17494,N_16157);
xnor U24175 (N_24175,N_19725,N_17741);
nand U24176 (N_24176,N_18292,N_18854);
xor U24177 (N_24177,N_19269,N_18624);
or U24178 (N_24178,N_16823,N_17527);
or U24179 (N_24179,N_16920,N_19455);
xnor U24180 (N_24180,N_17493,N_16783);
or U24181 (N_24181,N_16605,N_16671);
nor U24182 (N_24182,N_15699,N_19804);
xnor U24183 (N_24183,N_18652,N_18271);
or U24184 (N_24184,N_15932,N_15362);
or U24185 (N_24185,N_18563,N_17415);
or U24186 (N_24186,N_15528,N_18760);
nor U24187 (N_24187,N_16062,N_15707);
and U24188 (N_24188,N_17072,N_17609);
xor U24189 (N_24189,N_17758,N_18472);
xnor U24190 (N_24190,N_16703,N_16372);
nor U24191 (N_24191,N_15569,N_17686);
nand U24192 (N_24192,N_15535,N_17246);
nor U24193 (N_24193,N_17573,N_15240);
or U24194 (N_24194,N_17607,N_19728);
nor U24195 (N_24195,N_16835,N_19365);
xnor U24196 (N_24196,N_17888,N_19251);
and U24197 (N_24197,N_18735,N_15463);
nor U24198 (N_24198,N_18130,N_15240);
nand U24199 (N_24199,N_18585,N_19850);
nor U24200 (N_24200,N_16059,N_15738);
nand U24201 (N_24201,N_15076,N_19765);
or U24202 (N_24202,N_15483,N_17664);
nand U24203 (N_24203,N_15274,N_15496);
nor U24204 (N_24204,N_15076,N_19420);
nor U24205 (N_24205,N_17205,N_15144);
and U24206 (N_24206,N_17837,N_19998);
or U24207 (N_24207,N_18886,N_16691);
nor U24208 (N_24208,N_17478,N_19987);
nor U24209 (N_24209,N_18373,N_18178);
xnor U24210 (N_24210,N_17320,N_15598);
nand U24211 (N_24211,N_18893,N_16044);
xor U24212 (N_24212,N_15408,N_18434);
nor U24213 (N_24213,N_18400,N_17440);
and U24214 (N_24214,N_19844,N_18423);
nor U24215 (N_24215,N_16747,N_18215);
and U24216 (N_24216,N_16541,N_18991);
or U24217 (N_24217,N_16066,N_17247);
and U24218 (N_24218,N_16310,N_18217);
nor U24219 (N_24219,N_18314,N_15881);
nand U24220 (N_24220,N_16871,N_19346);
nand U24221 (N_24221,N_16811,N_19499);
or U24222 (N_24222,N_16451,N_15867);
and U24223 (N_24223,N_18421,N_15077);
nor U24224 (N_24224,N_16577,N_15375);
nand U24225 (N_24225,N_19398,N_16188);
nand U24226 (N_24226,N_17490,N_16078);
nand U24227 (N_24227,N_18272,N_16895);
and U24228 (N_24228,N_15092,N_17834);
and U24229 (N_24229,N_17579,N_15269);
and U24230 (N_24230,N_18220,N_16797);
nand U24231 (N_24231,N_18248,N_16357);
xor U24232 (N_24232,N_16310,N_17167);
nand U24233 (N_24233,N_16897,N_15499);
xor U24234 (N_24234,N_18220,N_19064);
or U24235 (N_24235,N_16126,N_16887);
xor U24236 (N_24236,N_16538,N_19314);
and U24237 (N_24237,N_19768,N_17728);
nor U24238 (N_24238,N_17055,N_18831);
xnor U24239 (N_24239,N_18030,N_17500);
or U24240 (N_24240,N_16917,N_19126);
and U24241 (N_24241,N_17559,N_15546);
and U24242 (N_24242,N_15807,N_18881);
nand U24243 (N_24243,N_18635,N_16943);
and U24244 (N_24244,N_19295,N_17589);
or U24245 (N_24245,N_16970,N_17783);
xor U24246 (N_24246,N_16469,N_18162);
nand U24247 (N_24247,N_18087,N_18674);
and U24248 (N_24248,N_15242,N_17450);
nor U24249 (N_24249,N_17918,N_18987);
and U24250 (N_24250,N_18774,N_15349);
or U24251 (N_24251,N_17213,N_16364);
and U24252 (N_24252,N_19983,N_19318);
and U24253 (N_24253,N_16363,N_17573);
nor U24254 (N_24254,N_16515,N_19028);
and U24255 (N_24255,N_18480,N_16835);
xnor U24256 (N_24256,N_16860,N_15098);
xor U24257 (N_24257,N_18236,N_17050);
xnor U24258 (N_24258,N_18700,N_19175);
nand U24259 (N_24259,N_16614,N_15924);
or U24260 (N_24260,N_16988,N_19345);
or U24261 (N_24261,N_15768,N_18056);
nand U24262 (N_24262,N_16564,N_19354);
or U24263 (N_24263,N_15371,N_15511);
or U24264 (N_24264,N_17797,N_15160);
or U24265 (N_24265,N_17286,N_19602);
nand U24266 (N_24266,N_16990,N_16828);
xnor U24267 (N_24267,N_17062,N_19044);
or U24268 (N_24268,N_17882,N_18432);
and U24269 (N_24269,N_19111,N_17051);
and U24270 (N_24270,N_19598,N_16634);
xnor U24271 (N_24271,N_19365,N_17737);
or U24272 (N_24272,N_16956,N_17793);
or U24273 (N_24273,N_17790,N_16537);
nand U24274 (N_24274,N_18181,N_15554);
and U24275 (N_24275,N_17683,N_18394);
nand U24276 (N_24276,N_16973,N_19768);
nor U24277 (N_24277,N_18991,N_16482);
and U24278 (N_24278,N_19060,N_16287);
and U24279 (N_24279,N_15137,N_18472);
nor U24280 (N_24280,N_18555,N_16920);
or U24281 (N_24281,N_15708,N_19008);
or U24282 (N_24282,N_19415,N_19439);
or U24283 (N_24283,N_18253,N_18904);
and U24284 (N_24284,N_17833,N_16493);
nand U24285 (N_24285,N_17249,N_17533);
nor U24286 (N_24286,N_18752,N_17496);
xnor U24287 (N_24287,N_18009,N_17088);
and U24288 (N_24288,N_15845,N_16753);
nand U24289 (N_24289,N_18302,N_15827);
and U24290 (N_24290,N_18821,N_16120);
nand U24291 (N_24291,N_15859,N_16895);
xor U24292 (N_24292,N_17795,N_19844);
nand U24293 (N_24293,N_19918,N_16853);
nor U24294 (N_24294,N_16791,N_19916);
xor U24295 (N_24295,N_16573,N_17964);
nand U24296 (N_24296,N_17133,N_15077);
nand U24297 (N_24297,N_18899,N_15821);
and U24298 (N_24298,N_15142,N_19682);
and U24299 (N_24299,N_19824,N_15647);
and U24300 (N_24300,N_17651,N_19686);
nor U24301 (N_24301,N_18868,N_15548);
xnor U24302 (N_24302,N_16202,N_17336);
xor U24303 (N_24303,N_15458,N_17590);
and U24304 (N_24304,N_16194,N_15001);
xnor U24305 (N_24305,N_18852,N_15429);
or U24306 (N_24306,N_17515,N_15763);
and U24307 (N_24307,N_17372,N_17021);
or U24308 (N_24308,N_17807,N_15606);
and U24309 (N_24309,N_16030,N_17552);
or U24310 (N_24310,N_19964,N_19665);
and U24311 (N_24311,N_15508,N_16878);
and U24312 (N_24312,N_18374,N_17515);
xor U24313 (N_24313,N_18054,N_19218);
and U24314 (N_24314,N_18247,N_16507);
and U24315 (N_24315,N_16225,N_19563);
nand U24316 (N_24316,N_19041,N_15631);
xor U24317 (N_24317,N_18994,N_18002);
xor U24318 (N_24318,N_19220,N_18851);
and U24319 (N_24319,N_15585,N_15124);
or U24320 (N_24320,N_17702,N_15375);
and U24321 (N_24321,N_19544,N_19319);
nand U24322 (N_24322,N_15277,N_16300);
and U24323 (N_24323,N_19296,N_17748);
xor U24324 (N_24324,N_18986,N_19977);
nand U24325 (N_24325,N_19101,N_18858);
or U24326 (N_24326,N_19782,N_18508);
xor U24327 (N_24327,N_16450,N_18811);
and U24328 (N_24328,N_16064,N_17373);
xnor U24329 (N_24329,N_18537,N_15286);
xor U24330 (N_24330,N_17622,N_17042);
nor U24331 (N_24331,N_18347,N_19653);
or U24332 (N_24332,N_19632,N_17230);
and U24333 (N_24333,N_18110,N_16972);
nand U24334 (N_24334,N_15007,N_16358);
xnor U24335 (N_24335,N_16605,N_15172);
or U24336 (N_24336,N_17357,N_18706);
nor U24337 (N_24337,N_18691,N_16011);
nor U24338 (N_24338,N_15943,N_15227);
nand U24339 (N_24339,N_17529,N_19049);
xor U24340 (N_24340,N_16737,N_15990);
and U24341 (N_24341,N_15036,N_19548);
or U24342 (N_24342,N_16081,N_15951);
or U24343 (N_24343,N_17243,N_16929);
nor U24344 (N_24344,N_19315,N_18699);
and U24345 (N_24345,N_15049,N_18433);
and U24346 (N_24346,N_17860,N_15337);
xor U24347 (N_24347,N_19539,N_18786);
nor U24348 (N_24348,N_17455,N_16366);
nor U24349 (N_24349,N_17283,N_16157);
nand U24350 (N_24350,N_16684,N_15938);
or U24351 (N_24351,N_18558,N_18441);
and U24352 (N_24352,N_19357,N_15793);
xnor U24353 (N_24353,N_19994,N_18837);
xor U24354 (N_24354,N_18516,N_19535);
and U24355 (N_24355,N_16570,N_15021);
nand U24356 (N_24356,N_15581,N_18615);
and U24357 (N_24357,N_19885,N_17026);
nor U24358 (N_24358,N_15919,N_18702);
or U24359 (N_24359,N_17478,N_18340);
or U24360 (N_24360,N_18333,N_16590);
nor U24361 (N_24361,N_17459,N_15034);
xnor U24362 (N_24362,N_17222,N_15912);
nor U24363 (N_24363,N_18481,N_18838);
xor U24364 (N_24364,N_16064,N_18703);
nor U24365 (N_24365,N_19299,N_18464);
nor U24366 (N_24366,N_18287,N_17286);
nand U24367 (N_24367,N_15217,N_15268);
or U24368 (N_24368,N_15257,N_16542);
or U24369 (N_24369,N_18074,N_17987);
nor U24370 (N_24370,N_19602,N_17859);
or U24371 (N_24371,N_16964,N_17397);
or U24372 (N_24372,N_19412,N_19609);
xor U24373 (N_24373,N_17309,N_19511);
nor U24374 (N_24374,N_18440,N_16405);
nand U24375 (N_24375,N_18531,N_17331);
nor U24376 (N_24376,N_17674,N_19311);
nor U24377 (N_24377,N_17805,N_18702);
nor U24378 (N_24378,N_18840,N_16710);
xnor U24379 (N_24379,N_18334,N_18590);
nand U24380 (N_24380,N_18744,N_17499);
nor U24381 (N_24381,N_17132,N_16765);
nor U24382 (N_24382,N_19500,N_17777);
nor U24383 (N_24383,N_15323,N_15894);
or U24384 (N_24384,N_19391,N_18753);
nand U24385 (N_24385,N_17442,N_15327);
or U24386 (N_24386,N_18347,N_18774);
or U24387 (N_24387,N_15534,N_15416);
or U24388 (N_24388,N_16499,N_15193);
nor U24389 (N_24389,N_16288,N_16469);
xnor U24390 (N_24390,N_16721,N_15053);
and U24391 (N_24391,N_19421,N_19225);
and U24392 (N_24392,N_16590,N_16232);
xnor U24393 (N_24393,N_16076,N_16276);
or U24394 (N_24394,N_17209,N_19912);
or U24395 (N_24395,N_17625,N_18601);
and U24396 (N_24396,N_18495,N_17153);
or U24397 (N_24397,N_17570,N_15752);
nor U24398 (N_24398,N_16855,N_18515);
nor U24399 (N_24399,N_18658,N_18647);
nand U24400 (N_24400,N_16410,N_17599);
or U24401 (N_24401,N_15134,N_18416);
and U24402 (N_24402,N_19246,N_18253);
xnor U24403 (N_24403,N_19165,N_18646);
xnor U24404 (N_24404,N_18575,N_19108);
xor U24405 (N_24405,N_19512,N_17394);
xor U24406 (N_24406,N_17617,N_16025);
or U24407 (N_24407,N_19042,N_16605);
xor U24408 (N_24408,N_18412,N_15818);
and U24409 (N_24409,N_18119,N_15390);
nor U24410 (N_24410,N_15318,N_16104);
nand U24411 (N_24411,N_19801,N_16441);
or U24412 (N_24412,N_18821,N_17971);
nand U24413 (N_24413,N_17941,N_17099);
or U24414 (N_24414,N_18501,N_17195);
and U24415 (N_24415,N_16167,N_18949);
and U24416 (N_24416,N_17375,N_16614);
and U24417 (N_24417,N_16655,N_19066);
nand U24418 (N_24418,N_19050,N_17230);
or U24419 (N_24419,N_15064,N_18864);
or U24420 (N_24420,N_19294,N_16270);
nand U24421 (N_24421,N_18619,N_17308);
and U24422 (N_24422,N_15917,N_16357);
or U24423 (N_24423,N_17231,N_18598);
xor U24424 (N_24424,N_15500,N_16605);
nor U24425 (N_24425,N_15658,N_18432);
nand U24426 (N_24426,N_17944,N_19012);
or U24427 (N_24427,N_15899,N_17170);
nor U24428 (N_24428,N_18051,N_16334);
xor U24429 (N_24429,N_19819,N_16928);
nor U24430 (N_24430,N_16747,N_17379);
nor U24431 (N_24431,N_15134,N_15314);
xor U24432 (N_24432,N_17319,N_16169);
and U24433 (N_24433,N_16254,N_18214);
nor U24434 (N_24434,N_15782,N_17242);
or U24435 (N_24435,N_16889,N_15393);
xor U24436 (N_24436,N_19634,N_16327);
or U24437 (N_24437,N_17858,N_15411);
nand U24438 (N_24438,N_16038,N_17583);
nor U24439 (N_24439,N_18300,N_15389);
xor U24440 (N_24440,N_19200,N_19058);
nand U24441 (N_24441,N_18833,N_19070);
nor U24442 (N_24442,N_17765,N_16876);
and U24443 (N_24443,N_18714,N_16426);
nor U24444 (N_24444,N_17584,N_15700);
nand U24445 (N_24445,N_17560,N_18421);
nand U24446 (N_24446,N_18453,N_18146);
and U24447 (N_24447,N_18955,N_19598);
nor U24448 (N_24448,N_19847,N_17007);
nand U24449 (N_24449,N_17293,N_15048);
nor U24450 (N_24450,N_15473,N_15601);
nand U24451 (N_24451,N_17199,N_15047);
nor U24452 (N_24452,N_18129,N_15825);
nor U24453 (N_24453,N_18093,N_17758);
and U24454 (N_24454,N_19646,N_17758);
or U24455 (N_24455,N_19822,N_17691);
and U24456 (N_24456,N_19474,N_19138);
and U24457 (N_24457,N_19759,N_17014);
nor U24458 (N_24458,N_16843,N_17396);
or U24459 (N_24459,N_17768,N_19997);
nor U24460 (N_24460,N_19424,N_15593);
nor U24461 (N_24461,N_19910,N_15459);
and U24462 (N_24462,N_18543,N_16693);
and U24463 (N_24463,N_16879,N_16001);
nand U24464 (N_24464,N_16282,N_17217);
nand U24465 (N_24465,N_15258,N_19775);
nand U24466 (N_24466,N_18429,N_15784);
xor U24467 (N_24467,N_15354,N_16354);
nor U24468 (N_24468,N_17190,N_15175);
xor U24469 (N_24469,N_15840,N_17860);
xnor U24470 (N_24470,N_18410,N_19935);
nand U24471 (N_24471,N_15182,N_19419);
nor U24472 (N_24472,N_18265,N_16653);
nand U24473 (N_24473,N_18772,N_18961);
xor U24474 (N_24474,N_19816,N_16450);
xnor U24475 (N_24475,N_19696,N_16251);
nor U24476 (N_24476,N_18990,N_16778);
xnor U24477 (N_24477,N_16431,N_17354);
and U24478 (N_24478,N_17620,N_17342);
nand U24479 (N_24479,N_17813,N_19474);
xor U24480 (N_24480,N_15865,N_18468);
nor U24481 (N_24481,N_19971,N_16562);
xnor U24482 (N_24482,N_18471,N_17769);
xnor U24483 (N_24483,N_17248,N_17365);
or U24484 (N_24484,N_18499,N_17223);
xnor U24485 (N_24485,N_17965,N_19708);
xor U24486 (N_24486,N_19387,N_17011);
nand U24487 (N_24487,N_15965,N_17570);
nor U24488 (N_24488,N_17470,N_18776);
or U24489 (N_24489,N_17829,N_19988);
nor U24490 (N_24490,N_18244,N_15940);
xnor U24491 (N_24491,N_17821,N_16374);
nor U24492 (N_24492,N_19932,N_16257);
xor U24493 (N_24493,N_17602,N_18822);
nor U24494 (N_24494,N_16683,N_19164);
or U24495 (N_24495,N_19220,N_15726);
nor U24496 (N_24496,N_16927,N_15630);
xor U24497 (N_24497,N_15257,N_15397);
or U24498 (N_24498,N_17236,N_16518);
and U24499 (N_24499,N_15094,N_15962);
or U24500 (N_24500,N_16226,N_17213);
and U24501 (N_24501,N_18344,N_18168);
nand U24502 (N_24502,N_17434,N_18321);
xor U24503 (N_24503,N_18251,N_15869);
and U24504 (N_24504,N_15672,N_15037);
and U24505 (N_24505,N_15948,N_16930);
or U24506 (N_24506,N_15324,N_15960);
or U24507 (N_24507,N_16897,N_18438);
and U24508 (N_24508,N_18975,N_19430);
xor U24509 (N_24509,N_16431,N_18741);
xor U24510 (N_24510,N_16172,N_19220);
xnor U24511 (N_24511,N_19261,N_18559);
xnor U24512 (N_24512,N_17343,N_19131);
nor U24513 (N_24513,N_16412,N_19143);
nand U24514 (N_24514,N_18408,N_19720);
or U24515 (N_24515,N_18380,N_15619);
and U24516 (N_24516,N_17724,N_17559);
nor U24517 (N_24517,N_17235,N_15515);
or U24518 (N_24518,N_16955,N_15234);
or U24519 (N_24519,N_16582,N_16273);
or U24520 (N_24520,N_19489,N_18886);
or U24521 (N_24521,N_16894,N_17197);
xnor U24522 (N_24522,N_15906,N_19295);
nor U24523 (N_24523,N_18992,N_18853);
xnor U24524 (N_24524,N_18233,N_16764);
or U24525 (N_24525,N_17874,N_16662);
and U24526 (N_24526,N_19546,N_17851);
nor U24527 (N_24527,N_19410,N_17251);
or U24528 (N_24528,N_15300,N_18387);
nor U24529 (N_24529,N_18861,N_18358);
or U24530 (N_24530,N_16445,N_18281);
and U24531 (N_24531,N_18382,N_16091);
and U24532 (N_24532,N_18136,N_17544);
xnor U24533 (N_24533,N_19269,N_18047);
nor U24534 (N_24534,N_16586,N_15477);
and U24535 (N_24535,N_15615,N_17510);
nand U24536 (N_24536,N_19034,N_16793);
xnor U24537 (N_24537,N_17776,N_18611);
and U24538 (N_24538,N_19989,N_17598);
nand U24539 (N_24539,N_17127,N_17508);
nor U24540 (N_24540,N_19006,N_15673);
or U24541 (N_24541,N_16768,N_16224);
or U24542 (N_24542,N_16323,N_17343);
and U24543 (N_24543,N_19580,N_17499);
xnor U24544 (N_24544,N_16987,N_17592);
xor U24545 (N_24545,N_18854,N_16751);
xor U24546 (N_24546,N_18668,N_17394);
and U24547 (N_24547,N_17472,N_15867);
or U24548 (N_24548,N_17453,N_18942);
or U24549 (N_24549,N_19517,N_16534);
nand U24550 (N_24550,N_16833,N_15064);
nor U24551 (N_24551,N_18330,N_15343);
xor U24552 (N_24552,N_15452,N_15638);
or U24553 (N_24553,N_17101,N_15278);
and U24554 (N_24554,N_15033,N_19346);
or U24555 (N_24555,N_19597,N_19610);
nor U24556 (N_24556,N_18492,N_16234);
xnor U24557 (N_24557,N_16868,N_15332);
xnor U24558 (N_24558,N_15119,N_16828);
nor U24559 (N_24559,N_18427,N_19445);
nand U24560 (N_24560,N_16045,N_18094);
xor U24561 (N_24561,N_19668,N_17607);
nand U24562 (N_24562,N_18531,N_15799);
nor U24563 (N_24563,N_18052,N_19484);
and U24564 (N_24564,N_19355,N_16754);
xor U24565 (N_24565,N_16392,N_19442);
and U24566 (N_24566,N_17478,N_16345);
xnor U24567 (N_24567,N_19282,N_19946);
and U24568 (N_24568,N_15042,N_16246);
or U24569 (N_24569,N_16591,N_18559);
xor U24570 (N_24570,N_19397,N_18713);
and U24571 (N_24571,N_19386,N_19184);
or U24572 (N_24572,N_15127,N_18271);
xor U24573 (N_24573,N_16376,N_19921);
nor U24574 (N_24574,N_17277,N_18101);
nor U24575 (N_24575,N_17464,N_18213);
or U24576 (N_24576,N_15002,N_15274);
nor U24577 (N_24577,N_15884,N_18303);
and U24578 (N_24578,N_19982,N_19703);
and U24579 (N_24579,N_19111,N_19072);
or U24580 (N_24580,N_19323,N_16129);
and U24581 (N_24581,N_19067,N_19942);
nor U24582 (N_24582,N_18004,N_19876);
and U24583 (N_24583,N_19156,N_18675);
or U24584 (N_24584,N_16980,N_18083);
and U24585 (N_24585,N_15313,N_17144);
nor U24586 (N_24586,N_15841,N_19382);
or U24587 (N_24587,N_18952,N_19151);
and U24588 (N_24588,N_18718,N_18808);
nor U24589 (N_24589,N_19794,N_19196);
nand U24590 (N_24590,N_16365,N_16499);
nor U24591 (N_24591,N_19150,N_17822);
or U24592 (N_24592,N_17175,N_17625);
or U24593 (N_24593,N_16873,N_18483);
and U24594 (N_24594,N_19187,N_16559);
nor U24595 (N_24595,N_17157,N_16236);
or U24596 (N_24596,N_18563,N_17367);
nor U24597 (N_24597,N_16634,N_19899);
or U24598 (N_24598,N_19741,N_16063);
nand U24599 (N_24599,N_19817,N_17801);
nand U24600 (N_24600,N_16339,N_18086);
nor U24601 (N_24601,N_17039,N_19413);
nand U24602 (N_24602,N_16204,N_15276);
nor U24603 (N_24603,N_15154,N_18667);
nor U24604 (N_24604,N_17589,N_19082);
or U24605 (N_24605,N_18079,N_15358);
xnor U24606 (N_24606,N_18539,N_17793);
nand U24607 (N_24607,N_17194,N_16885);
xnor U24608 (N_24608,N_17545,N_19872);
nand U24609 (N_24609,N_17819,N_17351);
nor U24610 (N_24610,N_18623,N_19514);
xnor U24611 (N_24611,N_19884,N_17317);
or U24612 (N_24612,N_16198,N_18631);
xor U24613 (N_24613,N_17220,N_16924);
nor U24614 (N_24614,N_19912,N_18359);
nand U24615 (N_24615,N_18006,N_17813);
nand U24616 (N_24616,N_15296,N_15406);
or U24617 (N_24617,N_16424,N_15931);
nand U24618 (N_24618,N_16829,N_16569);
and U24619 (N_24619,N_17316,N_18173);
nor U24620 (N_24620,N_17445,N_17253);
nand U24621 (N_24621,N_16855,N_19332);
nor U24622 (N_24622,N_17835,N_15982);
or U24623 (N_24623,N_18406,N_15172);
and U24624 (N_24624,N_18307,N_19263);
nor U24625 (N_24625,N_16358,N_17770);
or U24626 (N_24626,N_19850,N_16722);
or U24627 (N_24627,N_18241,N_16468);
and U24628 (N_24628,N_16150,N_15096);
or U24629 (N_24629,N_17276,N_18292);
or U24630 (N_24630,N_17260,N_19310);
nor U24631 (N_24631,N_16676,N_17307);
xnor U24632 (N_24632,N_16929,N_16642);
and U24633 (N_24633,N_16927,N_15990);
nor U24634 (N_24634,N_18106,N_16155);
xor U24635 (N_24635,N_17543,N_17156);
or U24636 (N_24636,N_16332,N_16550);
nand U24637 (N_24637,N_17368,N_18913);
nand U24638 (N_24638,N_17337,N_15940);
xnor U24639 (N_24639,N_18042,N_15272);
or U24640 (N_24640,N_19240,N_15518);
and U24641 (N_24641,N_16415,N_17945);
or U24642 (N_24642,N_19718,N_15342);
nand U24643 (N_24643,N_15958,N_19109);
and U24644 (N_24644,N_15728,N_19432);
nand U24645 (N_24645,N_17909,N_17885);
nor U24646 (N_24646,N_18343,N_19729);
nor U24647 (N_24647,N_17151,N_15115);
and U24648 (N_24648,N_18525,N_15059);
nand U24649 (N_24649,N_16445,N_18138);
and U24650 (N_24650,N_18152,N_19595);
or U24651 (N_24651,N_19493,N_17396);
or U24652 (N_24652,N_15356,N_18891);
xor U24653 (N_24653,N_16152,N_16296);
xor U24654 (N_24654,N_17568,N_16276);
and U24655 (N_24655,N_17413,N_19695);
xor U24656 (N_24656,N_15504,N_17880);
and U24657 (N_24657,N_15778,N_17747);
or U24658 (N_24658,N_17801,N_18204);
xnor U24659 (N_24659,N_17277,N_18399);
or U24660 (N_24660,N_15280,N_18291);
nand U24661 (N_24661,N_16638,N_17449);
nor U24662 (N_24662,N_19317,N_18226);
xor U24663 (N_24663,N_19608,N_18284);
xor U24664 (N_24664,N_15895,N_19056);
and U24665 (N_24665,N_15920,N_19312);
or U24666 (N_24666,N_15184,N_19180);
and U24667 (N_24667,N_17848,N_16025);
xnor U24668 (N_24668,N_16087,N_17922);
nor U24669 (N_24669,N_17547,N_15020);
nand U24670 (N_24670,N_18853,N_15196);
or U24671 (N_24671,N_16775,N_16401);
xor U24672 (N_24672,N_17338,N_17306);
nor U24673 (N_24673,N_17438,N_15788);
xor U24674 (N_24674,N_18693,N_19085);
nand U24675 (N_24675,N_15800,N_19929);
nand U24676 (N_24676,N_18994,N_18497);
or U24677 (N_24677,N_18278,N_15848);
nand U24678 (N_24678,N_16853,N_17360);
nand U24679 (N_24679,N_19338,N_17948);
and U24680 (N_24680,N_16268,N_16864);
xnor U24681 (N_24681,N_19627,N_16223);
nand U24682 (N_24682,N_15712,N_16365);
and U24683 (N_24683,N_17846,N_19617);
nand U24684 (N_24684,N_18807,N_16788);
nand U24685 (N_24685,N_18370,N_18765);
and U24686 (N_24686,N_19470,N_17961);
or U24687 (N_24687,N_19697,N_15540);
xor U24688 (N_24688,N_15852,N_19206);
xor U24689 (N_24689,N_19382,N_15540);
or U24690 (N_24690,N_19175,N_19000);
nor U24691 (N_24691,N_17852,N_18764);
or U24692 (N_24692,N_16284,N_18447);
or U24693 (N_24693,N_15144,N_17447);
xnor U24694 (N_24694,N_17722,N_17758);
nor U24695 (N_24695,N_16994,N_17316);
or U24696 (N_24696,N_19391,N_16650);
and U24697 (N_24697,N_15344,N_16783);
or U24698 (N_24698,N_15034,N_19722);
nor U24699 (N_24699,N_17298,N_17842);
and U24700 (N_24700,N_19555,N_16006);
nor U24701 (N_24701,N_18762,N_16070);
or U24702 (N_24702,N_19215,N_17398);
nor U24703 (N_24703,N_19590,N_16328);
or U24704 (N_24704,N_17728,N_18055);
or U24705 (N_24705,N_15043,N_17581);
xnor U24706 (N_24706,N_15941,N_16230);
xnor U24707 (N_24707,N_19962,N_15920);
nor U24708 (N_24708,N_17655,N_17273);
nand U24709 (N_24709,N_16963,N_15380);
xor U24710 (N_24710,N_18987,N_18017);
nor U24711 (N_24711,N_16099,N_15665);
nand U24712 (N_24712,N_18948,N_19984);
nand U24713 (N_24713,N_15790,N_19718);
xnor U24714 (N_24714,N_15904,N_16636);
and U24715 (N_24715,N_18826,N_18611);
nand U24716 (N_24716,N_15486,N_19546);
nand U24717 (N_24717,N_16241,N_15955);
and U24718 (N_24718,N_16624,N_19995);
xor U24719 (N_24719,N_18626,N_15385);
nand U24720 (N_24720,N_17974,N_15118);
or U24721 (N_24721,N_17716,N_19915);
and U24722 (N_24722,N_18094,N_17078);
and U24723 (N_24723,N_16701,N_17442);
or U24724 (N_24724,N_19813,N_18367);
nor U24725 (N_24725,N_18076,N_17609);
xnor U24726 (N_24726,N_16806,N_17434);
and U24727 (N_24727,N_17339,N_17360);
nor U24728 (N_24728,N_18282,N_18313);
nand U24729 (N_24729,N_16597,N_16920);
nand U24730 (N_24730,N_15467,N_19219);
nor U24731 (N_24731,N_18792,N_18555);
xnor U24732 (N_24732,N_19663,N_17344);
xor U24733 (N_24733,N_15717,N_18261);
and U24734 (N_24734,N_18583,N_17889);
nand U24735 (N_24735,N_17342,N_18304);
or U24736 (N_24736,N_15877,N_18080);
or U24737 (N_24737,N_15889,N_16926);
and U24738 (N_24738,N_17873,N_18742);
or U24739 (N_24739,N_18512,N_16091);
nand U24740 (N_24740,N_16388,N_15470);
xnor U24741 (N_24741,N_15064,N_16182);
nor U24742 (N_24742,N_18299,N_19354);
or U24743 (N_24743,N_17401,N_18809);
xor U24744 (N_24744,N_15192,N_16759);
xor U24745 (N_24745,N_17778,N_16878);
xnor U24746 (N_24746,N_15141,N_19209);
or U24747 (N_24747,N_17618,N_15044);
nor U24748 (N_24748,N_15598,N_15975);
and U24749 (N_24749,N_16221,N_19255);
nand U24750 (N_24750,N_15249,N_16900);
nor U24751 (N_24751,N_16552,N_17464);
xnor U24752 (N_24752,N_18496,N_17849);
nor U24753 (N_24753,N_16546,N_18855);
and U24754 (N_24754,N_19882,N_18167);
nand U24755 (N_24755,N_18501,N_19491);
nand U24756 (N_24756,N_19857,N_17650);
xnor U24757 (N_24757,N_16724,N_18258);
xnor U24758 (N_24758,N_15202,N_16027);
nor U24759 (N_24759,N_16417,N_17921);
or U24760 (N_24760,N_19245,N_19522);
xnor U24761 (N_24761,N_16735,N_16282);
nand U24762 (N_24762,N_15473,N_17275);
or U24763 (N_24763,N_16150,N_18895);
xnor U24764 (N_24764,N_16355,N_18321);
xnor U24765 (N_24765,N_15563,N_16367);
nor U24766 (N_24766,N_18938,N_16547);
and U24767 (N_24767,N_17074,N_17459);
nor U24768 (N_24768,N_17928,N_16066);
and U24769 (N_24769,N_17248,N_16722);
or U24770 (N_24770,N_17529,N_17041);
and U24771 (N_24771,N_17690,N_17677);
nand U24772 (N_24772,N_18567,N_19837);
nand U24773 (N_24773,N_18077,N_15461);
and U24774 (N_24774,N_19031,N_16451);
or U24775 (N_24775,N_16069,N_19996);
or U24776 (N_24776,N_19574,N_17192);
nand U24777 (N_24777,N_15250,N_19215);
and U24778 (N_24778,N_16783,N_16933);
or U24779 (N_24779,N_15486,N_18460);
and U24780 (N_24780,N_15051,N_16980);
nand U24781 (N_24781,N_18056,N_19145);
nand U24782 (N_24782,N_18614,N_17596);
or U24783 (N_24783,N_17365,N_19487);
nor U24784 (N_24784,N_16818,N_18374);
xnor U24785 (N_24785,N_15617,N_15270);
and U24786 (N_24786,N_15255,N_15213);
nor U24787 (N_24787,N_15409,N_19097);
nand U24788 (N_24788,N_17319,N_18635);
nor U24789 (N_24789,N_16217,N_17053);
or U24790 (N_24790,N_18736,N_15790);
nor U24791 (N_24791,N_18743,N_18337);
or U24792 (N_24792,N_18867,N_18090);
or U24793 (N_24793,N_15853,N_17848);
and U24794 (N_24794,N_17975,N_15206);
xor U24795 (N_24795,N_15142,N_19067);
xor U24796 (N_24796,N_18137,N_17531);
or U24797 (N_24797,N_18455,N_16707);
nor U24798 (N_24798,N_16463,N_19176);
and U24799 (N_24799,N_17589,N_15498);
and U24800 (N_24800,N_15265,N_15666);
nor U24801 (N_24801,N_19630,N_19717);
nor U24802 (N_24802,N_19779,N_15094);
xnor U24803 (N_24803,N_16482,N_18394);
xor U24804 (N_24804,N_18087,N_19061);
xnor U24805 (N_24805,N_15734,N_17999);
and U24806 (N_24806,N_18874,N_16258);
or U24807 (N_24807,N_18634,N_15331);
and U24808 (N_24808,N_16721,N_17637);
or U24809 (N_24809,N_16761,N_16692);
and U24810 (N_24810,N_17406,N_18093);
and U24811 (N_24811,N_19295,N_16181);
nand U24812 (N_24812,N_16566,N_16513);
xor U24813 (N_24813,N_19405,N_16526);
and U24814 (N_24814,N_15212,N_17790);
or U24815 (N_24815,N_18259,N_17829);
nand U24816 (N_24816,N_15029,N_19742);
nand U24817 (N_24817,N_19691,N_17443);
nand U24818 (N_24818,N_18864,N_18984);
or U24819 (N_24819,N_19637,N_16935);
and U24820 (N_24820,N_18422,N_19715);
nor U24821 (N_24821,N_17755,N_18501);
and U24822 (N_24822,N_18193,N_17160);
nor U24823 (N_24823,N_16038,N_18818);
nand U24824 (N_24824,N_15069,N_16723);
nor U24825 (N_24825,N_16086,N_18843);
xor U24826 (N_24826,N_19255,N_18280);
nor U24827 (N_24827,N_16320,N_16747);
nor U24828 (N_24828,N_16004,N_17696);
xnor U24829 (N_24829,N_15944,N_18255);
xnor U24830 (N_24830,N_18038,N_18132);
nand U24831 (N_24831,N_15799,N_18930);
and U24832 (N_24832,N_16843,N_19996);
and U24833 (N_24833,N_17267,N_18839);
or U24834 (N_24834,N_18258,N_18510);
nand U24835 (N_24835,N_16812,N_15307);
nor U24836 (N_24836,N_19158,N_15405);
nand U24837 (N_24837,N_17601,N_15691);
or U24838 (N_24838,N_18455,N_16361);
nor U24839 (N_24839,N_19858,N_18651);
and U24840 (N_24840,N_19145,N_16980);
and U24841 (N_24841,N_17572,N_18247);
and U24842 (N_24842,N_19402,N_18849);
xor U24843 (N_24843,N_17574,N_18371);
and U24844 (N_24844,N_15554,N_15224);
nor U24845 (N_24845,N_19068,N_15866);
or U24846 (N_24846,N_17686,N_18157);
xnor U24847 (N_24847,N_18025,N_18736);
and U24848 (N_24848,N_18301,N_19466);
nor U24849 (N_24849,N_16419,N_15035);
nand U24850 (N_24850,N_17029,N_18109);
xor U24851 (N_24851,N_17105,N_18330);
or U24852 (N_24852,N_17619,N_18204);
and U24853 (N_24853,N_17001,N_18551);
xor U24854 (N_24854,N_18500,N_15689);
nor U24855 (N_24855,N_18496,N_19303);
and U24856 (N_24856,N_17256,N_19018);
nand U24857 (N_24857,N_19547,N_17727);
nor U24858 (N_24858,N_19451,N_15415);
or U24859 (N_24859,N_18528,N_19927);
and U24860 (N_24860,N_17167,N_19145);
and U24861 (N_24861,N_18351,N_17092);
nor U24862 (N_24862,N_17165,N_19078);
or U24863 (N_24863,N_17554,N_17558);
and U24864 (N_24864,N_16483,N_19669);
nand U24865 (N_24865,N_18681,N_18654);
xnor U24866 (N_24866,N_19905,N_18827);
nor U24867 (N_24867,N_19391,N_18077);
and U24868 (N_24868,N_15270,N_18157);
xor U24869 (N_24869,N_19078,N_18005);
nand U24870 (N_24870,N_19713,N_19788);
or U24871 (N_24871,N_19535,N_18622);
nand U24872 (N_24872,N_19828,N_18308);
xnor U24873 (N_24873,N_19900,N_16458);
and U24874 (N_24874,N_17589,N_16244);
and U24875 (N_24875,N_19820,N_17222);
nand U24876 (N_24876,N_19114,N_16858);
nor U24877 (N_24877,N_17944,N_17405);
or U24878 (N_24878,N_16763,N_18499);
xor U24879 (N_24879,N_16753,N_15961);
xnor U24880 (N_24880,N_18088,N_16972);
and U24881 (N_24881,N_18697,N_17505);
nor U24882 (N_24882,N_19862,N_16834);
nand U24883 (N_24883,N_17851,N_18615);
xnor U24884 (N_24884,N_19514,N_19093);
nand U24885 (N_24885,N_17488,N_17749);
or U24886 (N_24886,N_18654,N_19498);
and U24887 (N_24887,N_15792,N_17972);
or U24888 (N_24888,N_17289,N_16581);
xnor U24889 (N_24889,N_17721,N_17247);
and U24890 (N_24890,N_16311,N_15672);
nor U24891 (N_24891,N_17680,N_16223);
nand U24892 (N_24892,N_19524,N_18311);
nor U24893 (N_24893,N_16853,N_17597);
nand U24894 (N_24894,N_17252,N_17149);
or U24895 (N_24895,N_19780,N_16575);
nor U24896 (N_24896,N_16923,N_18799);
and U24897 (N_24897,N_15123,N_16582);
and U24898 (N_24898,N_19613,N_17701);
nor U24899 (N_24899,N_15592,N_18863);
xor U24900 (N_24900,N_19261,N_15432);
xnor U24901 (N_24901,N_16939,N_17804);
nor U24902 (N_24902,N_19364,N_18198);
nor U24903 (N_24903,N_19092,N_16496);
nand U24904 (N_24904,N_17210,N_15111);
nand U24905 (N_24905,N_16328,N_18754);
and U24906 (N_24906,N_15782,N_15430);
or U24907 (N_24907,N_17234,N_16645);
xor U24908 (N_24908,N_15738,N_19183);
or U24909 (N_24909,N_15859,N_19596);
and U24910 (N_24910,N_18393,N_16018);
and U24911 (N_24911,N_15112,N_17882);
nor U24912 (N_24912,N_16395,N_19935);
xnor U24913 (N_24913,N_16025,N_19774);
nand U24914 (N_24914,N_19255,N_16739);
xnor U24915 (N_24915,N_17823,N_18098);
nand U24916 (N_24916,N_15522,N_18923);
xnor U24917 (N_24917,N_18243,N_17700);
or U24918 (N_24918,N_17463,N_19613);
xor U24919 (N_24919,N_17996,N_18516);
and U24920 (N_24920,N_17183,N_15428);
nor U24921 (N_24921,N_17736,N_18269);
nand U24922 (N_24922,N_15793,N_17674);
nand U24923 (N_24923,N_17658,N_19818);
or U24924 (N_24924,N_15397,N_18786);
or U24925 (N_24925,N_16139,N_16401);
or U24926 (N_24926,N_18626,N_16743);
and U24927 (N_24927,N_17943,N_17830);
nor U24928 (N_24928,N_18345,N_19039);
or U24929 (N_24929,N_18614,N_15934);
or U24930 (N_24930,N_17726,N_17617);
and U24931 (N_24931,N_19709,N_18089);
or U24932 (N_24932,N_18714,N_16492);
xor U24933 (N_24933,N_17931,N_17093);
nand U24934 (N_24934,N_19926,N_17990);
and U24935 (N_24935,N_16227,N_16733);
or U24936 (N_24936,N_15406,N_19351);
or U24937 (N_24937,N_18474,N_19696);
nor U24938 (N_24938,N_16063,N_18003);
or U24939 (N_24939,N_17047,N_18287);
nor U24940 (N_24940,N_16807,N_15810);
nor U24941 (N_24941,N_15888,N_19048);
or U24942 (N_24942,N_19760,N_17540);
xor U24943 (N_24943,N_19949,N_19962);
or U24944 (N_24944,N_16672,N_19104);
and U24945 (N_24945,N_18866,N_16020);
xor U24946 (N_24946,N_19548,N_18697);
xnor U24947 (N_24947,N_18631,N_19360);
nand U24948 (N_24948,N_17111,N_18346);
nand U24949 (N_24949,N_17918,N_15726);
nand U24950 (N_24950,N_16636,N_18778);
and U24951 (N_24951,N_15374,N_19364);
or U24952 (N_24952,N_15619,N_15727);
or U24953 (N_24953,N_17669,N_16191);
xor U24954 (N_24954,N_16880,N_18641);
nand U24955 (N_24955,N_19199,N_17078);
or U24956 (N_24956,N_19133,N_19969);
nand U24957 (N_24957,N_18607,N_18031);
or U24958 (N_24958,N_17530,N_15043);
and U24959 (N_24959,N_16283,N_19594);
nor U24960 (N_24960,N_17273,N_19467);
xor U24961 (N_24961,N_15391,N_19359);
and U24962 (N_24962,N_19062,N_15742);
nand U24963 (N_24963,N_19853,N_18830);
xnor U24964 (N_24964,N_17515,N_15257);
or U24965 (N_24965,N_15990,N_17695);
and U24966 (N_24966,N_17203,N_15843);
or U24967 (N_24967,N_15043,N_16406);
nor U24968 (N_24968,N_16142,N_16794);
nor U24969 (N_24969,N_16985,N_18675);
or U24970 (N_24970,N_15783,N_15186);
nand U24971 (N_24971,N_19601,N_18412);
or U24972 (N_24972,N_16114,N_16413);
nand U24973 (N_24973,N_15558,N_18269);
and U24974 (N_24974,N_16138,N_15289);
nand U24975 (N_24975,N_17242,N_16440);
nor U24976 (N_24976,N_16791,N_18510);
or U24977 (N_24977,N_15486,N_16839);
nand U24978 (N_24978,N_18608,N_18657);
xor U24979 (N_24979,N_16891,N_17452);
nor U24980 (N_24980,N_19714,N_17958);
or U24981 (N_24981,N_16376,N_15442);
and U24982 (N_24982,N_15926,N_18151);
and U24983 (N_24983,N_16593,N_17315);
or U24984 (N_24984,N_18326,N_17080);
and U24985 (N_24985,N_19169,N_19830);
nand U24986 (N_24986,N_16228,N_17728);
nor U24987 (N_24987,N_15286,N_17678);
nand U24988 (N_24988,N_16189,N_18870);
nand U24989 (N_24989,N_15018,N_15892);
nand U24990 (N_24990,N_19913,N_18457);
nand U24991 (N_24991,N_19464,N_18236);
and U24992 (N_24992,N_17787,N_19168);
nor U24993 (N_24993,N_18791,N_15632);
and U24994 (N_24994,N_18995,N_15311);
or U24995 (N_24995,N_15048,N_17470);
xnor U24996 (N_24996,N_15582,N_19516);
nand U24997 (N_24997,N_16714,N_16870);
nor U24998 (N_24998,N_18512,N_16764);
nor U24999 (N_24999,N_16526,N_17521);
nor U25000 (N_25000,N_20994,N_20935);
and U25001 (N_25001,N_23267,N_23054);
and U25002 (N_25002,N_21978,N_24836);
nand U25003 (N_25003,N_22324,N_24810);
or U25004 (N_25004,N_23690,N_21448);
nor U25005 (N_25005,N_21636,N_22367);
nand U25006 (N_25006,N_20517,N_22695);
nor U25007 (N_25007,N_20125,N_24484);
nand U25008 (N_25008,N_20087,N_24863);
or U25009 (N_25009,N_20059,N_20986);
xor U25010 (N_25010,N_22764,N_21659);
and U25011 (N_25011,N_22122,N_22230);
xnor U25012 (N_25012,N_20069,N_23473);
nor U25013 (N_25013,N_24471,N_24828);
and U25014 (N_25014,N_21902,N_24573);
and U25015 (N_25015,N_20704,N_21337);
or U25016 (N_25016,N_22504,N_20411);
or U25017 (N_25017,N_24513,N_20270);
and U25018 (N_25018,N_22569,N_24441);
or U25019 (N_25019,N_22580,N_24604);
xor U25020 (N_25020,N_20688,N_20181);
or U25021 (N_25021,N_22941,N_23102);
xor U25022 (N_25022,N_21302,N_24503);
and U25023 (N_25023,N_21262,N_20304);
xor U25024 (N_25024,N_23308,N_24050);
xor U25025 (N_25025,N_20220,N_22732);
nor U25026 (N_25026,N_21343,N_22151);
and U25027 (N_25027,N_22886,N_24387);
nand U25028 (N_25028,N_21016,N_23363);
or U25029 (N_25029,N_24028,N_24495);
nand U25030 (N_25030,N_22359,N_20095);
xnor U25031 (N_25031,N_20658,N_21348);
xor U25032 (N_25032,N_23554,N_21300);
or U25033 (N_25033,N_23620,N_21486);
and U25034 (N_25034,N_23646,N_21241);
nor U25035 (N_25035,N_21610,N_21047);
xor U25036 (N_25036,N_20939,N_20330);
or U25037 (N_25037,N_24696,N_23896);
and U25038 (N_25038,N_22404,N_22068);
and U25039 (N_25039,N_21235,N_21614);
nor U25040 (N_25040,N_23552,N_21417);
and U25041 (N_25041,N_21298,N_22576);
nor U25042 (N_25042,N_23687,N_20674);
nand U25043 (N_25043,N_23080,N_22493);
nor U25044 (N_25044,N_20637,N_23963);
or U25045 (N_25045,N_20878,N_21115);
or U25046 (N_25046,N_20138,N_21576);
and U25047 (N_25047,N_23011,N_20989);
xor U25048 (N_25048,N_23085,N_24148);
nor U25049 (N_25049,N_23979,N_23885);
nand U25050 (N_25050,N_20022,N_22366);
and U25051 (N_25051,N_20905,N_21023);
nand U25052 (N_25052,N_24116,N_20626);
nor U25053 (N_25053,N_23674,N_20021);
or U25054 (N_25054,N_20166,N_22100);
nor U25055 (N_25055,N_21216,N_20106);
and U25056 (N_25056,N_23930,N_22831);
nand U25057 (N_25057,N_20974,N_24791);
or U25058 (N_25058,N_20332,N_21371);
and U25059 (N_25059,N_20787,N_20980);
nand U25060 (N_25060,N_22360,N_20911);
nor U25061 (N_25061,N_23764,N_23947);
or U25062 (N_25062,N_22268,N_20144);
nand U25063 (N_25063,N_24758,N_23573);
or U25064 (N_25064,N_24579,N_24572);
xor U25065 (N_25065,N_22310,N_20193);
nor U25066 (N_25066,N_23544,N_22046);
and U25067 (N_25067,N_20689,N_24602);
nand U25068 (N_25068,N_24133,N_23458);
and U25069 (N_25069,N_22832,N_23701);
and U25070 (N_25070,N_23974,N_21281);
or U25071 (N_25071,N_21911,N_21273);
and U25072 (N_25072,N_23400,N_23742);
nand U25073 (N_25073,N_20274,N_23647);
or U25074 (N_25074,N_24629,N_24085);
and U25075 (N_25075,N_24100,N_20005);
or U25076 (N_25076,N_23733,N_21315);
xnor U25077 (N_25077,N_21490,N_24187);
or U25078 (N_25078,N_20412,N_24247);
xor U25079 (N_25079,N_22036,N_21325);
nand U25080 (N_25080,N_20768,N_24694);
nor U25081 (N_25081,N_21035,N_22882);
nor U25082 (N_25082,N_23104,N_21907);
or U25083 (N_25083,N_21946,N_20417);
xnor U25084 (N_25084,N_23890,N_24515);
nor U25085 (N_25085,N_23664,N_22468);
nor U25086 (N_25086,N_20035,N_24794);
nor U25087 (N_25087,N_22388,N_21901);
or U25088 (N_25088,N_22307,N_20129);
and U25089 (N_25089,N_23234,N_23824);
and U25090 (N_25090,N_22419,N_20908);
or U25091 (N_25091,N_24506,N_23900);
and U25092 (N_25092,N_21590,N_21691);
or U25093 (N_25093,N_20132,N_23180);
or U25094 (N_25094,N_22803,N_23019);
nand U25095 (N_25095,N_20840,N_20795);
nor U25096 (N_25096,N_21118,N_21772);
and U25097 (N_25097,N_24257,N_23295);
and U25098 (N_25098,N_24974,N_21932);
xnor U25099 (N_25099,N_21701,N_22523);
or U25100 (N_25100,N_24033,N_20718);
nor U25101 (N_25101,N_23698,N_22117);
and U25102 (N_25102,N_21621,N_23848);
xor U25103 (N_25103,N_24114,N_24264);
or U25104 (N_25104,N_22913,N_23721);
or U25105 (N_25105,N_22920,N_24489);
nor U25106 (N_25106,N_22270,N_21012);
and U25107 (N_25107,N_20030,N_22782);
nand U25108 (N_25108,N_22078,N_22980);
xnor U25109 (N_25109,N_21387,N_22605);
and U25110 (N_25110,N_20057,N_21852);
nor U25111 (N_25111,N_24212,N_22612);
nand U25112 (N_25112,N_24473,N_21109);
nor U25113 (N_25113,N_24708,N_21170);
or U25114 (N_25114,N_20807,N_21287);
or U25115 (N_25115,N_23422,N_21479);
and U25116 (N_25116,N_21573,N_21842);
or U25117 (N_25117,N_24802,N_23536);
nand U25118 (N_25118,N_22047,N_20261);
nor U25119 (N_25119,N_20845,N_20459);
or U25120 (N_25120,N_21703,N_23177);
xor U25121 (N_25121,N_21788,N_20897);
xnor U25122 (N_25122,N_20173,N_24551);
nand U25123 (N_25123,N_22616,N_21120);
or U25124 (N_25124,N_23596,N_20821);
nor U25125 (N_25125,N_22045,N_20971);
and U25126 (N_25126,N_20063,N_24436);
xor U25127 (N_25127,N_24955,N_20977);
xnor U25128 (N_25128,N_21061,N_24452);
or U25129 (N_25129,N_22051,N_22173);
and U25130 (N_25130,N_23655,N_23432);
xnor U25131 (N_25131,N_24711,N_23315);
or U25132 (N_25132,N_24988,N_20844);
xnor U25133 (N_25133,N_22639,N_24526);
nor U25134 (N_25134,N_20931,N_23513);
nand U25135 (N_25135,N_21961,N_24223);
and U25136 (N_25136,N_20218,N_21195);
nand U25137 (N_25137,N_21081,N_22836);
or U25138 (N_25138,N_22509,N_22397);
and U25139 (N_25139,N_23794,N_24216);
xor U25140 (N_25140,N_22017,N_21964);
nor U25141 (N_25141,N_21285,N_20549);
and U25142 (N_25142,N_20210,N_20273);
nand U25143 (N_25143,N_22623,N_21526);
xnor U25144 (N_25144,N_20298,N_22148);
xnor U25145 (N_25145,N_24851,N_23172);
xor U25146 (N_25146,N_23442,N_20376);
or U25147 (N_25147,N_20347,N_23207);
xor U25148 (N_25148,N_22220,N_23089);
and U25149 (N_25149,N_21257,N_23944);
nand U25150 (N_25150,N_20820,N_22169);
and U25151 (N_25151,N_20419,N_23840);
nor U25152 (N_25152,N_24585,N_21729);
xnor U25153 (N_25153,N_21456,N_24472);
and U25154 (N_25154,N_24895,N_23476);
nor U25155 (N_25155,N_22327,N_20227);
and U25156 (N_25156,N_22300,N_21347);
or U25157 (N_25157,N_23053,N_22071);
or U25158 (N_25158,N_24314,N_21543);
and U25159 (N_25159,N_21191,N_20188);
and U25160 (N_25160,N_21757,N_24049);
xor U25161 (N_25161,N_24368,N_23364);
or U25162 (N_25162,N_23821,N_20355);
xor U25163 (N_25163,N_20136,N_23776);
xor U25164 (N_25164,N_22384,N_20748);
nor U25165 (N_25165,N_24860,N_22872);
nand U25166 (N_25166,N_23411,N_20165);
and U25167 (N_25167,N_23167,N_21826);
nor U25168 (N_25168,N_20353,N_23078);
or U25169 (N_25169,N_21463,N_23635);
and U25170 (N_25170,N_22290,N_21723);
nor U25171 (N_25171,N_20947,N_22058);
and U25172 (N_25172,N_23171,N_21710);
or U25173 (N_25173,N_21785,N_22698);
or U25174 (N_25174,N_21917,N_22842);
nor U25175 (N_25175,N_23908,N_20640);
nand U25176 (N_25176,N_22684,N_22067);
nor U25177 (N_25177,N_22183,N_24866);
nand U25178 (N_25178,N_22704,N_20803);
nor U25179 (N_25179,N_21279,N_23713);
or U25180 (N_25180,N_21680,N_20211);
and U25181 (N_25181,N_20917,N_20946);
and U25182 (N_25182,N_24105,N_22355);
or U25183 (N_25183,N_20096,N_22779);
nand U25184 (N_25184,N_23287,N_20371);
nand U25185 (N_25185,N_23791,N_21155);
nor U25186 (N_25186,N_24180,N_21679);
xnor U25187 (N_25187,N_23741,N_23107);
nor U25188 (N_25188,N_24514,N_23567);
or U25189 (N_25189,N_20103,N_22902);
nor U25190 (N_25190,N_20725,N_21572);
xor U25191 (N_25191,N_23205,N_21158);
or U25192 (N_25192,N_20405,N_24981);
nand U25193 (N_25193,N_22552,N_24734);
nor U25194 (N_25194,N_22675,N_22891);
and U25195 (N_25195,N_23136,N_20791);
or U25196 (N_25196,N_22970,N_24095);
nand U25197 (N_25197,N_23148,N_20629);
nor U25198 (N_25198,N_20806,N_20323);
xor U25199 (N_25199,N_22571,N_23328);
and U25200 (N_25200,N_21827,N_22524);
nor U25201 (N_25201,N_24904,N_24448);
nand U25202 (N_25202,N_20809,N_21513);
or U25203 (N_25203,N_24975,N_20583);
nand U25204 (N_25204,N_22876,N_21224);
nand U25205 (N_25205,N_21683,N_23566);
xnor U25206 (N_25206,N_20161,N_21042);
nand U25207 (N_25207,N_22107,N_22425);
nor U25208 (N_25208,N_23321,N_24193);
or U25209 (N_25209,N_20607,N_24470);
nand U25210 (N_25210,N_24244,N_20385);
or U25211 (N_25211,N_22720,N_23756);
nor U25212 (N_25212,N_23925,N_24214);
nor U25213 (N_25213,N_23852,N_22655);
nand U25214 (N_25214,N_21750,N_22127);
and U25215 (N_25215,N_21251,N_24437);
xor U25216 (N_25216,N_22305,N_23462);
nor U25217 (N_25217,N_24576,N_20730);
xor U25218 (N_25218,N_23448,N_22936);
nand U25219 (N_25219,N_24291,N_20217);
nand U25220 (N_25220,N_20951,N_20401);
or U25221 (N_25221,N_22554,N_21447);
or U25222 (N_25222,N_24205,N_20901);
xor U25223 (N_25223,N_22240,N_24619);
and U25224 (N_25224,N_23586,N_22507);
xnor U25225 (N_25225,N_22018,N_22700);
or U25226 (N_25226,N_21424,N_24039);
nor U25227 (N_25227,N_20428,N_24393);
or U25228 (N_25228,N_24467,N_21949);
xnor U25229 (N_25229,N_22968,N_22674);
or U25230 (N_25230,N_21642,N_24752);
and U25231 (N_25231,N_23895,N_23705);
xnor U25232 (N_25232,N_23553,N_24031);
nor U25233 (N_25233,N_20363,N_23203);
nand U25234 (N_25234,N_21160,N_21982);
and U25235 (N_25235,N_24537,N_24270);
nor U25236 (N_25236,N_21899,N_20922);
xnor U25237 (N_25237,N_20687,N_22263);
or U25238 (N_25238,N_24906,N_24451);
nor U25239 (N_25239,N_24654,N_20723);
nor U25240 (N_25240,N_22330,N_22905);
nor U25241 (N_25241,N_21277,N_24927);
or U25242 (N_25242,N_24840,N_22588);
nand U25243 (N_25243,N_20311,N_24635);
nand U25244 (N_25244,N_22662,N_21380);
or U25245 (N_25245,N_23893,N_21464);
nor U25246 (N_25246,N_20987,N_22432);
and U25247 (N_25247,N_22904,N_23359);
xnor U25248 (N_25248,N_22219,N_22877);
xor U25249 (N_25249,N_21968,N_24333);
xnor U25250 (N_25250,N_24219,N_24192);
nand U25251 (N_25251,N_22761,N_24692);
or U25252 (N_25252,N_20249,N_20387);
nor U25253 (N_25253,N_22140,N_21648);
nor U25254 (N_25254,N_24279,N_22465);
xor U25255 (N_25255,N_20201,N_20187);
nand U25256 (N_25256,N_22277,N_21039);
xnor U25257 (N_25257,N_24486,N_24309);
nor U25258 (N_25258,N_23455,N_21475);
or U25259 (N_25259,N_21428,N_23498);
nor U25260 (N_25260,N_23212,N_24406);
or U25261 (N_25261,N_20959,N_22486);
nand U25262 (N_25262,N_21769,N_21773);
xor U25263 (N_25263,N_20116,N_23605);
or U25264 (N_25264,N_23463,N_20686);
nor U25265 (N_25265,N_20744,N_22824);
nor U25266 (N_25266,N_24175,N_20071);
or U25267 (N_25267,N_20802,N_23788);
nand U25268 (N_25268,N_21064,N_21225);
nor U25269 (N_25269,N_21079,N_23940);
xor U25270 (N_25270,N_21328,N_21681);
nor U25271 (N_25271,N_21686,N_20715);
nand U25272 (N_25272,N_21167,N_24403);
or U25273 (N_25273,N_24815,N_21809);
nand U25274 (N_25274,N_24672,N_23681);
nand U25275 (N_25275,N_24855,N_24960);
nor U25276 (N_25276,N_21781,N_23629);
nand U25277 (N_25277,N_23636,N_23158);
or U25278 (N_25278,N_23032,N_23391);
nor U25279 (N_25279,N_23174,N_22925);
nor U25280 (N_25280,N_24494,N_21290);
nand U25281 (N_25281,N_24786,N_24479);
or U25282 (N_25282,N_23751,N_20084);
nor U25283 (N_25283,N_23082,N_24342);
and U25284 (N_25284,N_23518,N_23031);
or U25285 (N_25285,N_22025,N_20796);
xnor U25286 (N_25286,N_21406,N_23650);
xnor U25287 (N_25287,N_21364,N_20487);
nor U25288 (N_25288,N_24996,N_23704);
and U25289 (N_25289,N_20893,N_22400);
nand U25290 (N_25290,N_23255,N_24676);
and U25291 (N_25291,N_22563,N_21232);
xnor U25292 (N_25292,N_22682,N_23071);
nand U25293 (N_25293,N_24150,N_24656);
and U25294 (N_25294,N_22194,N_22545);
or U25295 (N_25295,N_22659,N_24638);
nand U25296 (N_25296,N_21792,N_20455);
nand U25297 (N_25297,N_22844,N_20507);
xnor U25298 (N_25298,N_21635,N_24593);
nand U25299 (N_25299,N_23841,N_21765);
and U25300 (N_25300,N_22296,N_20317);
nand U25301 (N_25301,N_21937,N_23619);
nor U25302 (N_25302,N_22441,N_22322);
nor U25303 (N_25303,N_20282,N_20781);
nor U25304 (N_25304,N_22907,N_23770);
xnor U25305 (N_25305,N_20690,N_24926);
or U25306 (N_25306,N_24699,N_24340);
xnor U25307 (N_25307,N_23490,N_22619);
or U25308 (N_25308,N_21779,N_20623);
or U25309 (N_25309,N_21414,N_23798);
nand U25310 (N_25310,N_21820,N_20346);
or U25311 (N_25311,N_23334,N_22497);
nand U25312 (N_25312,N_23094,N_22777);
nand U25313 (N_25313,N_20968,N_21024);
and U25314 (N_25314,N_22378,N_20183);
or U25315 (N_25315,N_21980,N_22729);
nand U25316 (N_25316,N_20012,N_20427);
xor U25317 (N_25317,N_22829,N_24425);
xnor U25318 (N_25318,N_23757,N_23860);
or U25319 (N_25319,N_21518,N_22899);
nor U25320 (N_25320,N_24907,N_21077);
or U25321 (N_25321,N_22666,N_21133);
nand U25322 (N_25322,N_20657,N_20247);
xnor U25323 (N_25323,N_22175,N_21892);
and U25324 (N_25324,N_20604,N_24686);
or U25325 (N_25325,N_20779,N_22395);
nand U25326 (N_25326,N_21976,N_22265);
or U25327 (N_25327,N_20856,N_22917);
or U25328 (N_25328,N_20615,N_24400);
or U25329 (N_25329,N_21677,N_22204);
or U25330 (N_25330,N_24390,N_24339);
nor U25331 (N_25331,N_23665,N_20386);
nor U25332 (N_25332,N_24036,N_22440);
or U25333 (N_25333,N_22304,N_23105);
and U25334 (N_25334,N_24940,N_23736);
and U25335 (N_25335,N_23472,N_22299);
and U25336 (N_25336,N_23575,N_21927);
nand U25337 (N_25337,N_21309,N_20720);
nor U25338 (N_25338,N_20822,N_21615);
nor U25339 (N_25339,N_20631,N_24128);
and U25340 (N_25340,N_23820,N_23335);
nand U25341 (N_25341,N_20635,N_20262);
or U25342 (N_25342,N_23165,N_22631);
or U25343 (N_25343,N_20900,N_24939);
xor U25344 (N_25344,N_24596,N_24261);
and U25345 (N_25345,N_22869,N_22850);
nand U25346 (N_25346,N_21091,N_23541);
nand U25347 (N_25347,N_22621,N_23590);
or U25348 (N_25348,N_23491,N_20921);
and U25349 (N_25349,N_23987,N_20976);
nor U25350 (N_25350,N_23469,N_24041);
nand U25351 (N_25351,N_20842,N_24803);
and U25352 (N_25352,N_22939,N_23426);
and U25353 (N_25353,N_20521,N_21541);
nand U25354 (N_25354,N_20027,N_24127);
nor U25355 (N_25355,N_20747,N_21914);
and U25356 (N_25356,N_24421,N_23096);
nor U25357 (N_25357,N_23600,N_21972);
nor U25358 (N_25358,N_24529,N_22577);
or U25359 (N_25359,N_21661,N_22722);
and U25360 (N_25360,N_22976,N_20799);
or U25361 (N_25361,N_23970,N_22137);
xor U25362 (N_25362,N_21471,N_21009);
and U25363 (N_25363,N_23955,N_21231);
nand U25364 (N_25364,N_24396,N_24383);
nand U25365 (N_25365,N_23399,N_24322);
or U25366 (N_25366,N_20267,N_22422);
nor U25367 (N_25367,N_23216,N_21366);
xnor U25368 (N_25368,N_24580,N_22634);
xnor U25369 (N_25369,N_22863,N_24482);
or U25370 (N_25370,N_23272,N_23823);
and U25371 (N_25371,N_24885,N_23403);
xor U25372 (N_25372,N_23773,N_23163);
nor U25373 (N_25373,N_21666,N_24905);
xnor U25374 (N_25374,N_23068,N_23059);
and U25375 (N_25375,N_22889,N_23014);
and U25376 (N_25376,N_23867,N_24051);
or U25377 (N_25377,N_20654,N_23217);
xnor U25378 (N_25378,N_21459,N_21105);
or U25379 (N_25379,N_24542,N_21736);
xnor U25380 (N_25380,N_24060,N_20404);
nor U25381 (N_25381,N_21146,N_24121);
or U25382 (N_25382,N_24704,N_20389);
and U25383 (N_25383,N_23286,N_23168);
nand U25384 (N_25384,N_21386,N_24918);
xnor U25385 (N_25385,N_24023,N_20710);
nor U25386 (N_25386,N_22311,N_24915);
xor U25387 (N_25387,N_24883,N_23959);
xnor U25388 (N_25388,N_21295,N_21189);
or U25389 (N_25389,N_23630,N_21956);
nand U25390 (N_25390,N_22945,N_24160);
or U25391 (N_25391,N_24350,N_22013);
or U25392 (N_25392,N_23352,N_21596);
nor U25393 (N_25393,N_24949,N_22021);
or U25394 (N_25394,N_20743,N_22312);
xor U25395 (N_25395,N_23606,N_22548);
nor U25396 (N_25396,N_20661,N_22993);
or U25397 (N_25397,N_23584,N_20260);
and U25398 (N_25398,N_20301,N_20912);
or U25399 (N_25399,N_24652,N_20630);
xnor U25400 (N_25400,N_24004,N_21876);
nand U25401 (N_25401,N_20051,N_22023);
and U25402 (N_25402,N_21575,N_22691);
xor U25403 (N_25403,N_23747,N_21017);
or U25404 (N_25404,N_21981,N_20393);
nand U25405 (N_25405,N_23478,N_20192);
or U25406 (N_25406,N_22543,N_23306);
nand U25407 (N_25407,N_22737,N_23792);
and U25408 (N_25408,N_21829,N_21056);
nor U25409 (N_25409,N_24736,N_22599);
nor U25410 (N_25410,N_23484,N_24225);
nor U25411 (N_25411,N_21715,N_22730);
nand U25412 (N_25412,N_24826,N_24417);
and U25413 (N_25413,N_20128,N_22342);
nand U25414 (N_25414,N_24544,N_21897);
and U25415 (N_25415,N_23159,N_23583);
or U25416 (N_25416,N_22049,N_20316);
xnor U25417 (N_25417,N_20546,N_21570);
xor U25418 (N_25418,N_22822,N_24062);
nor U25419 (N_25419,N_24032,N_21605);
nand U25420 (N_25420,N_23574,N_21755);
or U25421 (N_25421,N_21114,N_23560);
and U25422 (N_25422,N_22202,N_24871);
or U25423 (N_25423,N_21752,N_23467);
or U25424 (N_25424,N_20773,N_20866);
xor U25425 (N_25425,N_23931,N_21721);
nor U25426 (N_25426,N_23210,N_23886);
and U25427 (N_25427,N_21999,N_21181);
xnor U25428 (N_25428,N_23826,N_23097);
or U25429 (N_25429,N_21175,N_20761);
xnor U25430 (N_25430,N_22344,N_24058);
and U25431 (N_25431,N_21935,N_21149);
nand U25432 (N_25432,N_22630,N_20678);
xnor U25433 (N_25433,N_24674,N_21088);
nor U25434 (N_25434,N_24080,N_20381);
and U25435 (N_25435,N_22225,N_20099);
or U25436 (N_25436,N_20573,N_24562);
and U25437 (N_25437,N_21288,N_24832);
xnor U25438 (N_25438,N_23202,N_22211);
and U25439 (N_25439,N_23018,N_21254);
xor U25440 (N_25440,N_22736,N_23769);
xor U25441 (N_25441,N_21354,N_20642);
and U25442 (N_25442,N_20612,N_23221);
and U25443 (N_25443,N_23452,N_24052);
and U25444 (N_25444,N_22858,N_22583);
and U25445 (N_25445,N_22178,N_22145);
and U25446 (N_25446,N_24937,N_24936);
xor U25447 (N_25447,N_24115,N_20650);
nand U25448 (N_25448,N_23240,N_21293);
xor U25449 (N_25449,N_23504,N_21623);
and U25450 (N_25450,N_21319,N_22817);
and U25451 (N_25451,N_20756,N_24217);
nand U25452 (N_25452,N_20685,N_21962);
and U25453 (N_25453,N_23051,N_22170);
nor U25454 (N_25454,N_22910,N_24901);
xnor U25455 (N_25455,N_20365,N_24712);
nor U25456 (N_25456,N_24152,N_24881);
xor U25457 (N_25457,N_23693,N_23892);
or U25458 (N_25458,N_21408,N_24977);
nor U25459 (N_25459,N_22705,N_20558);
nor U25460 (N_25460,N_23889,N_24560);
nand U25461 (N_25461,N_20200,N_21898);
nor U25462 (N_25462,N_22288,N_24986);
or U25463 (N_25463,N_22476,N_22979);
xor U25464 (N_25464,N_24663,N_20266);
and U25465 (N_25465,N_22082,N_24136);
or U25466 (N_25466,N_20159,N_22244);
nor U25467 (N_25467,N_23119,N_22550);
and U25468 (N_25468,N_22671,N_22261);
nand U25469 (N_25469,N_22014,N_21494);
nand U25470 (N_25470,N_23098,N_23616);
nor U25471 (N_25471,N_21502,N_20118);
nand U25472 (N_25472,N_21230,N_20497);
xor U25473 (N_25473,N_24898,N_22624);
or U25474 (N_25474,N_24878,N_21430);
or U25475 (N_25475,N_21075,N_22938);
and U25476 (N_25476,N_21402,N_21461);
and U25477 (N_25477,N_24285,N_24600);
and U25478 (N_25478,N_21807,N_22937);
xnor U25479 (N_25479,N_21110,N_24296);
or U25480 (N_25480,N_20966,N_20212);
nor U25481 (N_25481,N_20684,N_22234);
or U25482 (N_25482,N_21021,N_24555);
nand U25483 (N_25483,N_22650,N_20094);
nand U25484 (N_25484,N_24994,N_24741);
xor U25485 (N_25485,N_20195,N_24188);
nor U25486 (N_25486,N_23494,N_23135);
and U25487 (N_25487,N_20157,N_24304);
or U25488 (N_25488,N_23589,N_22594);
xor U25489 (N_25489,N_24185,N_21588);
nand U25490 (N_25490,N_20204,N_21672);
nor U25491 (N_25491,N_21753,N_22535);
and U25492 (N_25492,N_24414,N_22444);
nor U25493 (N_25493,N_21244,N_20603);
nor U25494 (N_25494,N_20049,N_21801);
and U25495 (N_25495,N_20460,N_21909);
xor U25496 (N_25496,N_23145,N_24892);
nand U25497 (N_25497,N_21746,N_23881);
nand U25498 (N_25498,N_22991,N_22079);
or U25499 (N_25499,N_20356,N_21699);
xnor U25500 (N_25500,N_21587,N_21790);
nor U25501 (N_25501,N_21934,N_23656);
xor U25502 (N_25502,N_21549,N_22697);
nor U25503 (N_25503,N_24424,N_21162);
or U25504 (N_25504,N_23219,N_20322);
nor U25505 (N_25505,N_23157,N_20757);
and U25506 (N_25506,N_21069,N_24026);
or U25507 (N_25507,N_22407,N_24415);
nand U25508 (N_25508,N_20503,N_24299);
xor U25509 (N_25509,N_22423,N_21329);
xnor U25510 (N_25510,N_21289,N_20065);
nor U25511 (N_25511,N_24307,N_20421);
nor U25512 (N_25512,N_23508,N_23754);
or U25513 (N_25513,N_23444,N_20598);
nor U25514 (N_25514,N_20235,N_22514);
nor U25515 (N_25515,N_24197,N_21488);
or U25516 (N_25516,N_23417,N_23904);
and U25517 (N_25517,N_20526,N_20068);
or U25518 (N_25518,N_21510,N_22541);
nor U25519 (N_25519,N_24386,N_24790);
and U25520 (N_25520,N_22719,N_21274);
nand U25521 (N_25521,N_23184,N_21970);
nand U25522 (N_25522,N_21080,N_21201);
and U25523 (N_25523,N_22450,N_23419);
and U25524 (N_25524,N_23735,N_22284);
and U25525 (N_25525,N_23877,N_21483);
and U25526 (N_25526,N_23370,N_22880);
nor U25527 (N_25527,N_24689,N_21043);
xor U25528 (N_25528,N_20256,N_24787);
and U25529 (N_25529,N_20746,N_22667);
and U25530 (N_25530,N_20438,N_22977);
nor U25531 (N_25531,N_21583,N_22713);
or U25532 (N_25532,N_23060,N_21758);
nand U25533 (N_25533,N_23680,N_20646);
xor U25534 (N_25534,N_24983,N_21465);
and U25535 (N_25535,N_20375,N_23752);
nand U25536 (N_25536,N_24982,N_20940);
and U25537 (N_25537,N_22478,N_24716);
nor U25538 (N_25538,N_23280,N_21540);
xor U25539 (N_25539,N_23236,N_22377);
xnor U25540 (N_25540,N_20683,N_22164);
xor U25541 (N_25541,N_23785,N_21164);
and U25542 (N_25542,N_22857,N_22665);
nand U25543 (N_25543,N_24732,N_22163);
xor U25544 (N_25544,N_22092,N_23389);
xor U25545 (N_25545,N_21791,N_20932);
and U25546 (N_25546,N_24615,N_21737);
nor U25547 (N_25547,N_22767,N_23418);
nand U25548 (N_25548,N_24327,N_24076);
nor U25549 (N_25549,N_23720,N_21228);
and U25550 (N_25550,N_23563,N_22115);
nand U25551 (N_25551,N_20611,N_21407);
nor U25552 (N_25552,N_21147,N_22708);
and U25553 (N_25553,N_22686,N_23438);
nor U25554 (N_25554,N_23628,N_22930);
or U25555 (N_25555,N_21132,N_21626);
nor U25556 (N_25556,N_23948,N_23602);
and U25557 (N_25557,N_21558,N_20407);
and U25558 (N_25558,N_24070,N_21700);
xor U25559 (N_25559,N_24138,N_23117);
nor U25560 (N_25560,N_24108,N_20763);
xnor U25561 (N_25561,N_21552,N_24657);
nand U25562 (N_25562,N_24282,N_23651);
or U25563 (N_25563,N_24017,N_23313);
and U25564 (N_25564,N_23353,N_22837);
nor U25565 (N_25565,N_20066,N_20519);
nor U25566 (N_25566,N_22198,N_23750);
or U25567 (N_25567,N_22370,N_20712);
and U25568 (N_25568,N_20950,N_20910);
nor U25569 (N_25569,N_21959,N_20139);
or U25570 (N_25570,N_20297,N_21263);
or U25571 (N_25571,N_23654,N_22405);
nor U25572 (N_25572,N_24557,N_23692);
nor U25573 (N_25573,N_23555,N_21550);
nor U25574 (N_25574,N_22205,N_21682);
and U25575 (N_25575,N_22218,N_22843);
nor U25576 (N_25576,N_20520,N_20784);
nor U25577 (N_25577,N_20281,N_22518);
nor U25578 (N_25578,N_22053,N_23740);
xor U25579 (N_25579,N_20081,N_22389);
nor U25580 (N_25580,N_22273,N_23185);
or U25581 (N_25581,N_20543,N_21814);
nand U25582 (N_25582,N_20186,N_22804);
and U25583 (N_25583,N_21524,N_23300);
and U25584 (N_25584,N_24764,N_23347);
xor U25585 (N_25585,N_24829,N_23638);
nor U25586 (N_25586,N_23627,N_21186);
xnor U25587 (N_25587,N_20341,N_22297);
nor U25588 (N_25588,N_20168,N_24606);
and U25589 (N_25589,N_24626,N_20018);
and U25590 (N_25590,N_23365,N_22592);
nand U25591 (N_25591,N_22676,N_24673);
nand U25592 (N_25592,N_20537,N_22960);
or U25593 (N_25593,N_24776,N_21248);
nand U25594 (N_25594,N_21307,N_20064);
nand U25595 (N_25595,N_21770,N_22814);
nor U25596 (N_25596,N_22138,N_21546);
and U25597 (N_25597,N_21333,N_21242);
nand U25598 (N_25598,N_22019,N_22638);
nand U25599 (N_25599,N_22011,N_22349);
nor U25600 (N_25600,N_21974,N_23739);
nor U25601 (N_25601,N_23164,N_20735);
and U25602 (N_25602,N_21220,N_23305);
nor U25603 (N_25603,N_23249,N_24438);
or U25604 (N_25604,N_23983,N_20749);
nand U25605 (N_25605,N_22967,N_20858);
xnor U25606 (N_25606,N_21304,N_23252);
and U25607 (N_25607,N_23188,N_24252);
nand U25608 (N_25608,N_20502,N_21784);
nand U25609 (N_25609,N_23039,N_22040);
nand U25610 (N_25610,N_20524,N_22947);
or U25611 (N_25611,N_21733,N_20992);
xor U25612 (N_25612,N_22663,N_22658);
nor U25613 (N_25613,N_23243,N_22525);
nor U25614 (N_25614,N_22186,N_22136);
or U25615 (N_25615,N_20416,N_24143);
or U25616 (N_25616,N_23338,N_24380);
xnor U25617 (N_25617,N_23984,N_24037);
or U25618 (N_25618,N_24389,N_22506);
xnor U25619 (N_25619,N_24595,N_21799);
nand U25620 (N_25620,N_23304,N_22853);
nor U25621 (N_25621,N_20926,N_23292);
nand U25622 (N_25622,N_20137,N_22969);
nor U25623 (N_25623,N_20213,N_24512);
xor U25624 (N_25624,N_22193,N_22932);
nand U25625 (N_25625,N_24844,N_21537);
or U25626 (N_25626,N_22114,N_22868);
xnor U25627 (N_25627,N_20666,N_24543);
and U25628 (N_25628,N_23169,N_21966);
and U25629 (N_25629,N_20745,N_21768);
and U25630 (N_25630,N_24891,N_21943);
nor U25631 (N_25631,N_22848,N_23858);
and U25632 (N_25632,N_24215,N_22901);
nand U25633 (N_25633,N_20740,N_23006);
and U25634 (N_25634,N_23341,N_21306);
or U25635 (N_25635,N_22208,N_24335);
and U25636 (N_25636,N_22678,N_24980);
nor U25637 (N_25637,N_20367,N_20606);
nand U25638 (N_25638,N_22614,N_24372);
xor U25639 (N_25639,N_24343,N_22413);
or U25640 (N_25640,N_20221,N_22001);
and U25641 (N_25641,N_22027,N_21604);
nor U25642 (N_25642,N_20877,N_20983);
nor U25643 (N_25643,N_23784,N_20191);
nor U25644 (N_25644,N_23263,N_22070);
and U25645 (N_25645,N_22227,N_22443);
or U25646 (N_25646,N_24651,N_24224);
or U25647 (N_25647,N_22762,N_20883);
nand U25648 (N_25648,N_24948,N_20566);
or U25649 (N_25649,N_24728,N_21520);
or U25650 (N_25650,N_24107,N_21895);
and U25651 (N_25651,N_20268,N_23471);
nand U25652 (N_25652,N_21203,N_21505);
nor U25653 (N_25653,N_24235,N_22231);
or U25654 (N_25654,N_24524,N_24920);
or U25655 (N_25655,N_24043,N_20437);
nor U25656 (N_25656,N_24687,N_21098);
nand U25657 (N_25657,N_20290,N_23291);
and U25658 (N_25658,N_23303,N_22073);
or U25659 (N_25659,N_21891,N_21469);
xnor U25660 (N_25660,N_22459,N_21468);
nand U25661 (N_25661,N_24811,N_21390);
xor U25662 (N_25662,N_20060,N_20008);
and U25663 (N_25663,N_22611,N_21063);
nor U25664 (N_25664,N_22709,N_21345);
or U25665 (N_25665,N_23383,N_22086);
nor U25666 (N_25666,N_24293,N_22978);
xnor U25667 (N_25667,N_20206,N_23564);
or U25668 (N_25668,N_23851,N_20484);
or U25669 (N_25669,N_21812,N_21744);
and U25670 (N_25670,N_20945,N_24377);
nor U25671 (N_25671,N_22409,N_21633);
nand U25672 (N_25672,N_24492,N_22426);
xor U25673 (N_25673,N_22933,N_24118);
nand U25674 (N_25674,N_23131,N_20568);
nand U25675 (N_25675,N_24166,N_23141);
nand U25676 (N_25676,N_22015,N_21735);
nor U25677 (N_25677,N_20010,N_21443);
nor U25678 (N_25678,N_23774,N_21070);
or U25679 (N_25679,N_24226,N_24351);
and U25680 (N_25680,N_22152,N_21015);
xnor U25681 (N_25681,N_23749,N_21905);
and U25682 (N_25682,N_22951,N_23525);
and U25683 (N_25683,N_22806,N_22233);
and U25684 (N_25684,N_22020,N_21392);
nand U25685 (N_25685,N_22540,N_21159);
nor U25686 (N_25686,N_20007,N_20104);
or U25687 (N_25687,N_22989,N_21495);
nand U25688 (N_25688,N_23395,N_21771);
or U25689 (N_25689,N_21501,N_22654);
xor U25690 (N_25690,N_23481,N_24646);
nand U25691 (N_25691,N_23023,N_20360);
nor U25692 (N_25692,N_21986,N_21280);
or U25693 (N_25693,N_24642,N_22847);
and U25694 (N_25694,N_22412,N_24364);
and U25695 (N_25695,N_23108,N_21127);
and U25696 (N_25696,N_23916,N_21894);
xor U25697 (N_25697,N_21460,N_22123);
nand U25698 (N_25698,N_21997,N_23845);
nand U25699 (N_25699,N_20726,N_21850);
xor U25700 (N_25700,N_24722,N_22604);
nor U25701 (N_25701,N_20776,N_20232);
nand U25702 (N_25702,N_24101,N_23763);
nand U25703 (N_25703,N_24238,N_22885);
nand U25704 (N_25704,N_22402,N_20814);
or U25705 (N_25705,N_24363,N_22000);
xnor U25706 (N_25706,N_22710,N_22357);
nor U25707 (N_25707,N_23933,N_20088);
nor U25708 (N_25708,N_22010,N_24770);
or U25709 (N_25709,N_22321,N_24607);
and U25710 (N_25710,N_23331,N_24027);
xor U25711 (N_25711,N_23095,N_20619);
and U25712 (N_25712,N_22491,N_20728);
and U25713 (N_25713,N_23397,N_20870);
and U25714 (N_25714,N_21645,N_24319);
nand U25715 (N_25715,N_24772,N_24917);
nand U25716 (N_25716,N_20390,N_23819);
xor U25717 (N_25717,N_24852,N_21868);
nand U25718 (N_25718,N_22495,N_21859);
or U25719 (N_25719,N_24730,N_21156);
xor U25720 (N_25720,N_22317,N_22895);
or U25721 (N_25721,N_22394,N_22813);
nand U25722 (N_25722,N_20564,N_21984);
or U25723 (N_25723,N_24229,N_20599);
nand U25724 (N_25724,N_23310,N_23501);
nand U25725 (N_25725,N_24227,N_23568);
nor U25726 (N_25726,N_21432,N_23194);
nor U25727 (N_25727,N_20855,N_21848);
and U25728 (N_25728,N_21382,N_23453);
nor U25729 (N_25729,N_21515,N_22787);
and U25730 (N_25730,N_23711,N_23007);
nand U25731 (N_25731,N_20028,N_20176);
and U25732 (N_25732,N_22908,N_23775);
nand U25733 (N_25733,N_22551,N_20565);
nor U25734 (N_25734,N_23813,N_22446);
or U25735 (N_25735,N_24814,N_24785);
xnor U25736 (N_25736,N_22066,N_20047);
xnor U25737 (N_25737,N_24231,N_24502);
nand U25738 (N_25738,N_20350,N_23803);
and U25739 (N_25739,N_21171,N_22786);
nand U25740 (N_25740,N_23844,N_21419);
and U25741 (N_25741,N_24220,N_20216);
or U25742 (N_25742,N_21963,N_24963);
and U25743 (N_25743,N_21173,N_22098);
and U25744 (N_25744,N_22089,N_21884);
or U25745 (N_25745,N_21462,N_22095);
or U25746 (N_25746,N_24173,N_20377);
xor U25747 (N_25747,N_21074,N_23571);
and U25748 (N_25748,N_23220,N_23799);
or U25749 (N_25749,N_24877,N_21261);
and U25750 (N_25750,N_21396,N_24648);
xnor U25751 (N_25751,N_24098,N_22093);
nor U25752 (N_25752,N_23079,N_22085);
and U25753 (N_25753,N_20145,N_23339);
and U25754 (N_25754,N_20396,N_23012);
or U25755 (N_25755,N_22593,N_23561);
xnor U25756 (N_25756,N_23807,N_20527);
xnor U25757 (N_25757,N_20923,N_23715);
nor U25758 (N_25758,N_20622,N_24218);
or U25759 (N_25759,N_24976,N_22801);
and U25760 (N_25760,N_22091,N_24093);
or U25761 (N_25761,N_23723,N_22641);
xor U25762 (N_25762,N_24094,N_24887);
nand U25763 (N_25763,N_20578,N_23384);
xor U25764 (N_25764,N_22003,N_24658);
or U25765 (N_25765,N_20885,N_22354);
xnor U25766 (N_25766,N_20034,N_22097);
xor U25767 (N_25767,N_24067,N_23748);
nand U25768 (N_25768,N_24819,N_23612);
xnor U25769 (N_25769,N_23708,N_21165);
nor U25770 (N_25770,N_20525,N_24057);
and U25771 (N_25771,N_20205,N_24015);
xor U25772 (N_25772,N_24624,N_23991);
nor U25773 (N_25773,N_21996,N_23888);
nor U25774 (N_25774,N_20529,N_24903);
nor U25775 (N_25775,N_24659,N_23128);
and U25776 (N_25776,N_24102,N_22002);
or U25777 (N_25777,N_23482,N_20602);
xor U25778 (N_25778,N_24329,N_20097);
or U25779 (N_25779,N_22453,N_24888);
nand U25780 (N_25780,N_20692,N_20155);
nor U25781 (N_25781,N_21994,N_24206);
and U25782 (N_25782,N_23326,N_23649);
or U25783 (N_25783,N_21908,N_20609);
nor U25784 (N_25784,N_24581,N_21268);
xnor U25785 (N_25785,N_23546,N_20703);
nor U25786 (N_25786,N_22336,N_24404);
or U25787 (N_25787,N_23632,N_22797);
xnor U25788 (N_25788,N_20575,N_22192);
nor U25789 (N_25789,N_23282,N_21592);
or U25790 (N_25790,N_23624,N_20861);
xor U25791 (N_25791,N_20229,N_20724);
nand U25792 (N_25792,N_23714,N_24487);
nor U25793 (N_25793,N_20962,N_21922);
xnor U25794 (N_25794,N_24016,N_24348);
and U25795 (N_25795,N_21863,N_23761);
xnor U25796 (N_25796,N_22132,N_24099);
and U25797 (N_25797,N_21836,N_21767);
nor U25798 (N_25798,N_23170,N_21816);
and U25799 (N_25799,N_22293,N_24410);
and U25800 (N_25800,N_20464,N_21514);
nor U25801 (N_25801,N_24260,N_20303);
xnor U25802 (N_25802,N_22005,N_22226);
and U25803 (N_25803,N_24065,N_22534);
nand U25804 (N_25804,N_21593,N_21239);
and U25805 (N_25805,N_20043,N_21747);
nand U25806 (N_25806,N_20253,N_22982);
nand U25807 (N_25807,N_20248,N_23755);
or U25808 (N_25808,N_20440,N_23371);
and U25809 (N_25809,N_21497,N_21639);
and U25810 (N_25810,N_22726,N_20751);
or U25811 (N_25811,N_23686,N_23658);
nor U25812 (N_25812,N_22608,N_24455);
nor U25813 (N_25813,N_21182,N_21453);
nor U25814 (N_25814,N_22096,N_24913);
nor U25815 (N_25815,N_23778,N_24540);
xnor U25816 (N_25816,N_24800,N_20616);
xor U25817 (N_25817,N_23201,N_21822);
nor U25818 (N_25818,N_24630,N_20919);
xor U25819 (N_25819,N_22255,N_20454);
and U25820 (N_25820,N_24053,N_22759);
nor U25821 (N_25821,N_21793,N_23683);
and U25822 (N_25822,N_22505,N_20942);
nand U25823 (N_25823,N_20996,N_24969);
and U25824 (N_25824,N_24729,N_20557);
nand U25825 (N_25825,N_22485,N_23069);
and U25826 (N_25826,N_23042,N_20706);
nand U25827 (N_25827,N_23949,N_22635);
nand U25828 (N_25828,N_23958,N_22499);
nand U25829 (N_25829,N_22496,N_24306);
nor U25830 (N_25830,N_20015,N_20163);
nand U25831 (N_25831,N_22928,N_22781);
and U25832 (N_25832,N_24132,N_24934);
nand U25833 (N_25833,N_22530,N_22435);
nand U25834 (N_25834,N_20750,N_23228);
and U25835 (N_25835,N_20089,N_23519);
nand U25836 (N_25836,N_23869,N_24597);
nor U25837 (N_25837,N_23617,N_21296);
nand U25838 (N_25838,N_21803,N_20914);
and U25839 (N_25839,N_22083,N_24078);
nor U25840 (N_25840,N_23677,N_23659);
or U25841 (N_25841,N_23719,N_21872);
and U25842 (N_25842,N_22747,N_23298);
and U25843 (N_25843,N_24158,N_24822);
nand U25844 (N_25844,N_22381,N_21825);
xnor U25845 (N_25845,N_23239,N_24493);
xnor U25846 (N_25846,N_21153,N_21521);
xor U25847 (N_25847,N_22069,N_22442);
nor U25848 (N_25848,N_20960,N_22106);
and U25849 (N_25849,N_20569,N_23517);
nand U25850 (N_25850,N_24376,N_24831);
nand U25851 (N_25851,N_24003,N_21442);
xnor U25852 (N_25852,N_20032,N_20970);
nand U25853 (N_25853,N_20816,N_20760);
nand U25854 (N_25854,N_24995,N_23129);
nand U25855 (N_25855,N_21847,N_24263);
and U25856 (N_25856,N_24880,N_20567);
and U25857 (N_25857,N_23923,N_21594);
xnor U25858 (N_25858,N_24527,N_23530);
nand U25859 (N_25859,N_24818,N_20889);
and U25860 (N_25860,N_24541,N_21253);
or U25861 (N_25861,N_21356,N_22037);
xnor U25862 (N_25862,N_20857,N_22455);
xor U25863 (N_25863,N_23706,N_20729);
xor U25864 (N_25864,N_21048,N_22998);
or U25865 (N_25865,N_23302,N_20002);
and U25866 (N_25866,N_20277,N_21264);
or U25867 (N_25867,N_21689,N_24274);
or U25868 (N_25868,N_24523,N_23762);
and U25869 (N_25869,N_21215,N_21650);
xor U25870 (N_25870,N_23336,N_22896);
or U25871 (N_25871,N_24534,N_23929);
nor U25872 (N_25872,N_24181,N_21476);
or U25873 (N_25873,N_23248,N_24320);
or U25874 (N_25874,N_22555,N_21269);
nand U25875 (N_25875,N_20196,N_24256);
nand U25876 (N_25876,N_21104,N_24784);
nor U25877 (N_25877,N_24805,N_20156);
nor U25878 (N_25878,N_23868,N_23642);
nand U25879 (N_25879,N_24938,N_21841);
nor U25880 (N_25880,N_22615,N_23618);
nand U25881 (N_25881,N_23866,N_20969);
nor U25882 (N_25882,N_22579,N_23558);
nor U25883 (N_25883,N_21106,N_21503);
nor U25884 (N_25884,N_24516,N_23323);
nor U25885 (N_25885,N_20124,N_21987);
nor U25886 (N_25886,N_21741,N_21742);
or U25887 (N_25887,N_20587,N_22673);
or U25888 (N_25888,N_23832,N_21227);
and U25889 (N_25889,N_24644,N_20597);
or U25890 (N_25890,N_21399,N_24042);
and U25891 (N_25891,N_21873,N_24678);
or U25892 (N_25892,N_23855,N_21619);
or U25893 (N_25893,N_21940,N_22012);
and U25894 (N_25894,N_24884,N_20753);
or U25895 (N_25895,N_21995,N_23192);
nor U25896 (N_25896,N_21815,N_20676);
or U25897 (N_25897,N_23973,N_24627);
xnor U25898 (N_25898,N_24521,N_24925);
nor U25899 (N_25899,N_24733,N_23849);
nand U25900 (N_25900,N_23998,N_23905);
and U25901 (N_25901,N_24623,N_21355);
and U25902 (N_25902,N_21305,N_21924);
xnor U25903 (N_25903,N_21211,N_21643);
nor U25904 (N_25904,N_22339,N_23430);
nor U25905 (N_25905,N_20033,N_22916);
xnor U25906 (N_25906,N_23369,N_21671);
xor U25907 (N_25907,N_23535,N_22602);
nand U25908 (N_25908,N_23507,N_24952);
or U25909 (N_25909,N_20675,N_23256);
or U25910 (N_25910,N_21835,N_22888);
nand U25911 (N_25911,N_23124,N_20467);
nor U25912 (N_25912,N_24167,N_22306);
xnor U25913 (N_25913,N_23029,N_23503);
xnor U25914 (N_25914,N_21368,N_23522);
nand U25915 (N_25915,N_21324,N_21313);
nand U25916 (N_25916,N_20559,N_23045);
and U25917 (N_25917,N_23694,N_20766);
and U25918 (N_25918,N_23260,N_22189);
xor U25919 (N_25919,N_22934,N_23717);
nor U25920 (N_25920,N_24705,N_23645);
xnor U25921 (N_25921,N_21528,N_22846);
nor U25922 (N_25922,N_22873,N_24021);
nor U25923 (N_25923,N_23547,N_21933);
xor U25924 (N_25924,N_20009,N_24685);
nand U25925 (N_25925,N_21172,N_20943);
nand U25926 (N_25926,N_23809,N_20896);
nor U25927 (N_25927,N_20636,N_21378);
or U25928 (N_25928,N_24879,N_23731);
or U25929 (N_25929,N_21690,N_21693);
nor U25930 (N_25930,N_23333,N_23675);
nor U25931 (N_25931,N_22918,N_20638);
nor U25932 (N_25932,N_23375,N_23040);
nor U25933 (N_25933,N_20798,N_23515);
nand U25934 (N_25934,N_20279,N_20083);
or U25935 (N_25935,N_23842,N_20770);
nand U25936 (N_25936,N_21629,N_23034);
or U25937 (N_25937,N_22460,N_21896);
xnor U25938 (N_25938,N_21582,N_24923);
nand U25939 (N_25939,N_21886,N_23499);
and U25940 (N_25940,N_22785,N_21885);
nor U25941 (N_25941,N_20456,N_24972);
and U25942 (N_25942,N_21204,N_20130);
xor U25943 (N_25943,N_24824,N_21702);
xnor U25944 (N_25944,N_23972,N_22439);
xor U25945 (N_25945,N_21275,N_20052);
nor U25946 (N_25946,N_22721,N_20736);
nand U25947 (N_25947,N_23960,N_24442);
nor U25948 (N_25948,N_20516,N_24719);
xnor U25949 (N_25949,N_20511,N_24834);
and U25950 (N_25950,N_23912,N_23093);
nor U25951 (N_25951,N_22584,N_23818);
and U25952 (N_25952,N_21580,N_21395);
or U25953 (N_25953,N_21748,N_24675);
or U25954 (N_25954,N_23376,N_23075);
nor U25955 (N_25955,N_23829,N_21669);
nand U25956 (N_25956,N_20352,N_23643);
and U25957 (N_25957,N_24843,N_21103);
nand U25958 (N_25958,N_23539,N_21818);
nor U25959 (N_25959,N_20620,N_22451);
or U25960 (N_25960,N_23502,N_20869);
and U25961 (N_25961,N_23149,N_20532);
xnor U25962 (N_25962,N_21716,N_22723);
xor U25963 (N_25963,N_21845,N_23483);
and U25964 (N_25964,N_20148,N_24771);
nor U25965 (N_25965,N_24780,N_23449);
nor U25966 (N_25966,N_20506,N_24566);
nand U25967 (N_25967,N_20036,N_24849);
nand U25968 (N_25968,N_23008,N_24366);
nor U25969 (N_25969,N_22177,N_20056);
or U25970 (N_25970,N_24097,N_21210);
nor U25971 (N_25971,N_22798,N_22778);
nor U25972 (N_25972,N_22390,N_22826);
nand U25973 (N_25973,N_22914,N_22156);
or U25974 (N_25974,N_22477,N_20494);
and U25975 (N_25975,N_20890,N_22789);
or U25976 (N_25976,N_24315,N_24190);
or U25977 (N_25977,N_21890,N_20681);
nand U25978 (N_25978,N_21138,N_24552);
nor U25979 (N_25979,N_21992,N_21466);
or U25980 (N_25980,N_23110,N_20716);
xor U25981 (N_25981,N_21709,N_22161);
nor U25982 (N_25982,N_20933,N_23283);
and U25983 (N_25983,N_20208,N_21482);
and U25984 (N_25984,N_23917,N_24754);
and U25985 (N_25985,N_22958,N_20477);
nand U25986 (N_25986,N_20649,N_20378);
nor U25987 (N_25987,N_23480,N_21777);
and U25988 (N_25988,N_22690,N_20329);
nor U25989 (N_25989,N_24288,N_20383);
nand U25990 (N_25990,N_24454,N_24172);
or U25991 (N_25991,N_24924,N_22546);
nor U25992 (N_25992,N_20518,N_23850);
xor U25993 (N_25993,N_23937,N_21092);
nor U25994 (N_25994,N_22050,N_23670);
xnor U25995 (N_25995,N_22597,N_22190);
nand U25996 (N_25996,N_23003,N_23357);
and U25997 (N_25997,N_23978,N_23440);
and U25998 (N_25998,N_21266,N_22356);
and U25999 (N_25999,N_23247,N_20754);
xnor U26000 (N_26000,N_21731,N_24253);
or U26001 (N_26001,N_24536,N_22646);
or U26002 (N_26002,N_21252,N_22223);
nand U26003 (N_26003,N_20194,N_23597);
nand U26004 (N_26004,N_23587,N_23943);
nand U26005 (N_26005,N_21446,N_21794);
xnor U26006 (N_26006,N_21194,N_23130);
and U26007 (N_26007,N_23468,N_23865);
nand U26008 (N_26008,N_23951,N_24240);
and U26009 (N_26009,N_24075,N_22154);
xnor U26010 (N_26010,N_22434,N_23578);
or U26011 (N_26011,N_20801,N_20483);
nand U26012 (N_26012,N_24381,N_20984);
xor U26013 (N_26013,N_24869,N_22319);
or U26014 (N_26014,N_21036,N_22769);
nand U26015 (N_26015,N_21179,N_23786);
nor U26016 (N_26016,N_23175,N_20269);
nor U26017 (N_26017,N_22661,N_22617);
nand U26018 (N_26018,N_24632,N_21223);
xnor U26019 (N_26019,N_22259,N_23288);
nor U26020 (N_26020,N_20349,N_24483);
and U26021 (N_26021,N_20430,N_24498);
or U26022 (N_26022,N_23344,N_20415);
and U26023 (N_26023,N_24007,N_20535);
nor U26024 (N_26024,N_20498,N_20334);
or U26025 (N_26025,N_23309,N_23700);
and U26026 (N_26026,N_20853,N_24807);
xnor U26027 (N_26027,N_22679,N_22055);
and U26028 (N_26028,N_20595,N_24153);
nand U26029 (N_26029,N_22487,N_21196);
and U26030 (N_26030,N_21101,N_21010);
and U26031 (N_26031,N_24522,N_20244);
xor U26032 (N_26032,N_21844,N_21323);
and U26033 (N_26033,N_23941,N_21856);
or U26034 (N_26034,N_21373,N_21121);
nor U26035 (N_26035,N_20852,N_23907);
xnor U26036 (N_26036,N_24558,N_21119);
and U26037 (N_26037,N_23966,N_20702);
nor U26038 (N_26038,N_20954,N_20143);
or U26039 (N_26039,N_23543,N_22841);
and U26040 (N_26040,N_22200,N_23067);
nor U26041 (N_26041,N_23673,N_24010);
nand U26042 (N_26042,N_22492,N_20326);
nand U26043 (N_26043,N_24286,N_23406);
and U26044 (N_26044,N_22022,N_22498);
xor U26045 (N_26045,N_22228,N_21640);
nand U26046 (N_26046,N_21067,N_21874);
nand U26047 (N_26047,N_22986,N_24063);
nor U26048 (N_26048,N_21385,N_23257);
xor U26049 (N_26049,N_23134,N_22501);
or U26050 (N_26050,N_20433,N_21749);
nand U26051 (N_26051,N_23611,N_21928);
xor U26052 (N_26052,N_20046,N_20907);
nand U26053 (N_26053,N_23846,N_22110);
and U26054 (N_26054,N_23367,N_24653);
nand U26055 (N_26055,N_22254,N_23744);
nor U26056 (N_26056,N_22503,N_20114);
and U26057 (N_26057,N_24897,N_21157);
or U26058 (N_26058,N_23716,N_24886);
and U26059 (N_26059,N_20647,N_21774);
nand U26060 (N_26060,N_21651,N_21944);
and U26061 (N_26061,N_21455,N_24025);
nand U26062 (N_26062,N_24858,N_23827);
xnor U26063 (N_26063,N_22433,N_21499);
and U26064 (N_26064,N_21249,N_20785);
nand U26065 (N_26065,N_22398,N_22207);
xnor U26066 (N_26066,N_20872,N_24086);
nand U26067 (N_26067,N_20874,N_24269);
or U26068 (N_26068,N_23005,N_24317);
xnor U26069 (N_26069,N_23186,N_23634);
and U26070 (N_26070,N_24577,N_22510);
xor U26071 (N_26071,N_24999,N_21002);
xnor U26072 (N_26072,N_21030,N_21631);
nor U26073 (N_26073,N_21685,N_24959);
xnor U26074 (N_26074,N_21440,N_20040);
or U26075 (N_26075,N_22214,N_21154);
nand U26076 (N_26076,N_22056,N_23529);
or U26077 (N_26077,N_22340,N_20541);
nand U26078 (N_26078,N_24701,N_23588);
nor U26079 (N_26079,N_21357,N_23026);
xnor U26080 (N_26080,N_22135,N_21960);
or U26081 (N_26081,N_20509,N_21603);
nor U26082 (N_26082,N_22116,N_24480);
or U26083 (N_26083,N_20981,N_22792);
and U26084 (N_26084,N_24505,N_24827);
nor U26085 (N_26085,N_21169,N_21051);
xor U26086 (N_26086,N_20850,N_24151);
or U26087 (N_26087,N_23922,N_22150);
or U26088 (N_26088,N_21539,N_22609);
xor U26089 (N_26089,N_20648,N_22302);
xnor U26090 (N_26090,N_23621,N_23924);
nor U26091 (N_26091,N_20944,N_24628);
or U26092 (N_26092,N_21553,N_24550);
or U26093 (N_26093,N_23349,N_24456);
xnor U26094 (N_26094,N_24222,N_23676);
and U26095 (N_26095,N_20925,N_20677);
xor U26096 (N_26096,N_22484,N_20714);
and U26097 (N_26097,N_20285,N_24125);
nor U26098 (N_26098,N_20767,N_23196);
nor U26099 (N_26099,N_24731,N_22687);
and U26100 (N_26100,N_24990,N_22805);
and U26101 (N_26101,N_23162,N_24398);
nor U26102 (N_26102,N_22217,N_24777);
nor U26103 (N_26103,N_20388,N_23354);
or U26104 (N_26104,N_21134,N_21602);
and U26105 (N_26105,N_21206,N_24491);
or U26106 (N_26106,N_21318,N_24374);
and U26107 (N_26107,N_23594,N_23037);
xor U26108 (N_26108,N_23576,N_24889);
nor U26109 (N_26109,N_24056,N_21751);
xnor U26110 (N_26110,N_21798,N_22289);
nand U26111 (N_26111,N_21435,N_22931);
nand U26112 (N_26112,N_22415,N_24809);
xor U26113 (N_26113,N_23802,N_23464);
xor U26114 (N_26114,N_23077,N_20909);
or U26115 (N_26115,N_24801,N_20092);
xor U26116 (N_26116,N_20127,N_24013);
nor U26117 (N_26117,N_22464,N_20471);
xnor U26118 (N_26118,N_22809,N_23559);
nor U26119 (N_26119,N_23903,N_24046);
or U26120 (N_26120,N_21862,N_22557);
xnor U26121 (N_26121,N_21617,N_24164);
nand U26122 (N_26122,N_23771,N_24677);
and U26123 (N_26123,N_20793,N_21314);
or U26124 (N_26124,N_23439,N_20160);
and U26125 (N_26125,N_23155,N_20733);
xnor U26126 (N_26126,N_22463,N_22652);
xnor U26127 (N_26127,N_20691,N_20561);
and U26128 (N_26128,N_20058,N_20150);
nor U26129 (N_26129,N_24305,N_22802);
nand U26130 (N_26130,N_24700,N_23322);
or U26131 (N_26131,N_20293,N_22924);
nor U26132 (N_26132,N_23864,N_24103);
xor U26133 (N_26133,N_21879,N_22399);
xor U26134 (N_26134,N_24792,N_21046);
nand U26135 (N_26135,N_24428,N_20679);
xor U26136 (N_26136,N_23935,N_23810);
xor U26137 (N_26137,N_21865,N_24688);
nand U26138 (N_26138,N_20126,N_23254);
xor U26139 (N_26139,N_22840,N_21229);
xnor U26140 (N_26140,N_23401,N_23126);
nand U26141 (N_26141,N_24636,N_23737);
or U26142 (N_26142,N_20479,N_22335);
nand U26143 (N_26143,N_23825,N_22981);
and U26144 (N_26144,N_21126,N_21344);
nand U26145 (N_26145,N_21367,N_22222);
or U26146 (N_26146,N_21439,N_22935);
nor U26147 (N_26147,N_20466,N_20177);
and U26148 (N_26148,N_24744,N_23662);
xor U26149 (N_26149,N_21696,N_20851);
nand U26150 (N_26150,N_22346,N_23603);
xnor U26151 (N_26151,N_24129,N_20403);
xor U26152 (N_26152,N_21034,N_23797);
xnor U26153 (N_26153,N_21838,N_24055);
xnor U26154 (N_26154,N_21756,N_20903);
nand U26155 (N_26155,N_22770,N_22266);
and U26156 (N_26156,N_23434,N_24767);
nand U26157 (N_26157,N_23317,N_20169);
xor U26158 (N_26158,N_22915,N_22084);
or U26159 (N_26159,N_22209,N_23876);
or U26160 (N_26160,N_23238,N_20246);
nor U26161 (N_26161,N_22247,N_24248);
nor U26162 (N_26162,N_23114,N_21111);
nand U26163 (N_26163,N_23639,N_21571);
nor U26164 (N_26164,N_22744,N_20671);
and U26165 (N_26165,N_21782,N_23100);
nor U26166 (N_26166,N_21516,N_20711);
and U26167 (N_26167,N_20924,N_21931);
and U26168 (N_26168,N_24749,N_23640);
nand U26169 (N_26169,N_22041,N_24622);
and U26170 (N_26170,N_21317,N_22995);
nor U26171 (N_26171,N_22956,N_24496);
nand U26172 (N_26172,N_21137,N_23815);
and U26173 (N_26173,N_23857,N_20794);
and U26174 (N_26174,N_24429,N_21577);
and U26175 (N_26175,N_22607,N_24661);
nor U26176 (N_26176,N_22111,N_24074);
nand U26177 (N_26177,N_20288,N_24354);
nand U26178 (N_26178,N_22285,N_22065);
or U26179 (N_26179,N_20006,N_22315);
and U26180 (N_26180,N_21150,N_22418);
xor U26181 (N_26181,N_20577,N_21087);
xnor U26182 (N_26182,N_20764,N_23839);
xnor U26183 (N_26183,N_22807,N_23009);
xor U26184 (N_26184,N_23783,N_20617);
or U26185 (N_26185,N_20812,N_24778);
nor U26186 (N_26186,N_24616,N_20336);
nand U26187 (N_26187,N_21834,N_22892);
nor U26188 (N_26188,N_22212,N_24433);
and U26189 (N_26189,N_24817,N_24228);
or U26190 (N_26190,N_22626,N_23076);
and U26191 (N_26191,N_24476,N_21823);
xor U26192 (N_26192,N_20461,N_21561);
nor U26193 (N_26193,N_24258,N_21544);
and U26194 (N_26194,N_23526,N_21441);
nand U26195 (N_26195,N_20149,N_21436);
xnor U26196 (N_26196,N_24798,N_24045);
or U26197 (N_26197,N_21370,N_22795);
xor U26198 (N_26198,N_20472,N_23329);
nor U26199 (N_26199,N_21942,N_22707);
xor U26200 (N_26200,N_24945,N_24533);
nand U26201 (N_26201,N_21058,N_23609);
nand U26202 (N_26202,N_24145,N_23028);
xnor U26203 (N_26203,N_24242,N_21839);
xor U26204 (N_26204,N_22119,N_23660);
xnor U26205 (N_26205,N_23127,N_21449);
nand U26206 (N_26206,N_20624,N_23613);
or U26207 (N_26207,N_22187,N_24157);
nor U26208 (N_26208,N_21198,N_24953);
or U26209 (N_26209,N_23016,N_20310);
nor U26210 (N_26210,N_22923,N_23374);
nand U26211 (N_26211,N_20927,N_21320);
and U26212 (N_26212,N_23261,N_22866);
xor U26213 (N_26213,N_22077,N_23245);
nor U26214 (N_26214,N_22267,N_20886);
and U26215 (N_26215,N_22508,N_24266);
xor U26216 (N_26216,N_23301,N_21951);
nor U26217 (N_26217,N_20110,N_22291);
or U26218 (N_26218,N_22912,N_22029);
or U26219 (N_26219,N_23942,N_24788);
xnor U26220 (N_26220,N_22323,N_24588);
nor U26221 (N_26221,N_21945,N_24896);
nand U26222 (N_26222,N_21384,N_20345);
xor U26223 (N_26223,N_24401,N_22677);
and U26224 (N_26224,N_21340,N_21397);
and U26225 (N_26225,N_21952,N_22232);
or U26226 (N_26226,N_20324,N_21941);
nor U26227 (N_26227,N_22739,N_24357);
xnor U26228 (N_26228,N_24011,N_22474);
and U26229 (N_26229,N_21389,N_21647);
and U26230 (N_26230,N_22500,N_21238);
nor U26231 (N_26231,N_22333,N_23516);
xor U26232 (N_26232,N_24446,N_20402);
or U26233 (N_26233,N_20374,N_22681);
nand U26234 (N_26234,N_22983,N_20839);
nand U26235 (N_26235,N_22855,N_23396);
nor U26236 (N_26236,N_22038,N_24567);
or U26237 (N_26237,N_22517,N_22757);
and U26238 (N_26238,N_21451,N_20338);
nor U26239 (N_26239,N_20379,N_21649);
and U26240 (N_26240,N_20589,N_21005);
nor U26241 (N_26241,N_24481,N_22727);
or U26242 (N_26242,N_21129,N_23796);
nand U26243 (N_26243,N_21775,N_23542);
nor U26244 (N_26244,N_20991,N_24402);
or U26245 (N_26245,N_24292,N_21411);
nor U26246 (N_26246,N_23181,N_21166);
nor U26247 (N_26247,N_24379,N_21762);
xor U26248 (N_26248,N_22854,N_23492);
nand U26249 (N_26249,N_22246,N_22637);
xnor U26250 (N_26250,N_23420,N_24237);
and U26251 (N_26251,N_20458,N_24302);
xnor U26252 (N_26252,N_23269,N_22174);
xor U26253 (N_26253,N_23615,N_23910);
nand U26254 (N_26254,N_20026,N_22740);
or U26255 (N_26255,N_23488,N_20141);
nor U26256 (N_26256,N_20938,N_21620);
nand U26257 (N_26257,N_21766,N_21711);
or U26258 (N_26258,N_22772,N_23065);
nand U26259 (N_26259,N_24199,N_21316);
nor U26260 (N_26260,N_20593,N_22565);
xnor U26261 (N_26261,N_23327,N_23427);
xor U26262 (N_26262,N_20031,N_21485);
or U26263 (N_26263,N_22856,N_21342);
or U26264 (N_26264,N_21301,N_23150);
and U26265 (N_26265,N_24933,N_23994);
nor U26266 (N_26266,N_22436,N_21278);
nand U26267 (N_26267,N_21113,N_20435);
nand U26268 (N_26268,N_22196,N_23091);
nor U26269 (N_26269,N_23271,N_20394);
xnor U26270 (N_26270,N_20672,N_23856);
nor U26271 (N_26271,N_21212,N_24059);
or U26272 (N_26272,N_22570,N_23020);
nand U26273 (N_26273,N_23570,N_21125);
nand U26274 (N_26274,N_21888,N_20255);
or U26275 (N_26275,N_23533,N_23195);
or U26276 (N_26276,N_24141,N_24842);
nor U26277 (N_26277,N_24316,N_24928);
nor U26278 (N_26278,N_23198,N_24755);
nand U26279 (N_26279,N_20209,N_23265);
xor U26280 (N_26280,N_20633,N_24432);
xnor U26281 (N_26281,N_20928,N_20550);
nor U26282 (N_26282,N_22522,N_24942);
or U26283 (N_26283,N_22158,N_20879);
xnor U26284 (N_26284,N_21525,N_23689);
nand U26285 (N_26285,N_22600,N_24323);
xnor U26286 (N_26286,N_20772,N_21918);
nor U26287 (N_26287,N_23608,N_21925);
nand U26288 (N_26288,N_23225,N_20560);
nor U26289 (N_26289,N_22343,N_24142);
and U26290 (N_26290,N_24946,N_23883);
xnor U26291 (N_26291,N_20848,N_21116);
or U26292 (N_26292,N_21086,N_20420);
nor U26293 (N_26293,N_21638,N_21877);
nand U26294 (N_26294,N_22033,N_21547);
or U26295 (N_26295,N_23377,N_21973);
nand U26296 (N_26296,N_20547,N_21403);
or U26297 (N_26297,N_24126,N_20572);
or U26298 (N_26298,N_21031,N_24048);
or U26299 (N_26299,N_24856,N_21018);
and U26300 (N_26300,N_21117,N_22649);
and U26301 (N_26301,N_22734,N_22042);
xnor U26302 (N_26302,N_20447,N_20488);
nor U26303 (N_26303,N_20955,N_22758);
nor U26304 (N_26304,N_24113,N_23527);
and U26305 (N_26305,N_20392,N_24239);
nor U26306 (N_26306,N_23743,N_21102);
or U26307 (N_26307,N_21761,N_21335);
xnor U26308 (N_26308,N_23780,N_22295);
nand U26309 (N_26309,N_24964,N_22887);
and U26310 (N_26310,N_24773,N_24717);
or U26311 (N_26311,N_23139,N_24637);
or U26312 (N_26312,N_22985,N_20788);
xor U26313 (N_26313,N_22622,N_22996);
nand U26314 (N_26314,N_20463,N_20846);
and U26315 (N_26315,N_21983,N_24563);
nor U26316 (N_26316,N_20563,N_21145);
xor U26317 (N_26317,N_23314,N_20739);
and U26318 (N_26318,N_22075,N_20584);
and U26319 (N_26319,N_22533,N_24349);
or U26320 (N_26320,N_24670,N_23115);
xor U26321 (N_26321,N_23534,N_23429);
nor U26322 (N_26322,N_21969,N_21041);
or U26323 (N_26323,N_20588,N_23266);
and U26324 (N_26324,N_21606,N_21557);
or U26325 (N_26325,N_23398,N_21143);
nand U26326 (N_26326,N_20863,N_24511);
or U26327 (N_26327,N_22898,N_24549);
nor U26328 (N_26328,N_20695,N_23268);
and U26329 (N_26329,N_22521,N_22922);
or U26330 (N_26330,N_24440,N_20997);
and U26331 (N_26331,N_24609,N_24412);
xor U26332 (N_26332,N_21670,N_23120);
nor U26333 (N_26333,N_24775,N_20252);
nand U26334 (N_26334,N_24762,N_20373);
nand U26335 (N_26335,N_23348,N_24804);
nand U26336 (N_26336,N_21967,N_22748);
nor U26337 (N_26337,N_23918,N_20272);
nor U26338 (N_26338,N_21778,N_24159);
xnor U26339 (N_26339,N_23416,N_22147);
nand U26340 (N_26340,N_21352,N_21350);
xnor U26341 (N_26341,N_24556,N_23625);
nor U26342 (N_26342,N_21719,N_23793);
nand U26343 (N_26343,N_21427,N_22642);
xnor U26344 (N_26344,N_21535,N_22104);
nor U26345 (N_26345,N_21393,N_23766);
nand U26346 (N_26346,N_21270,N_20759);
and U26347 (N_26347,N_21450,N_23988);
xor U26348 (N_26348,N_23610,N_24034);
and U26349 (N_26349,N_23407,N_24813);
or U26350 (N_26350,N_22909,N_22210);
or U26351 (N_26351,N_23279,N_21500);
xor U26352 (N_26352,N_23622,N_24392);
xor U26353 (N_26353,N_24519,N_22818);
xnor U26354 (N_26354,N_20585,N_20215);
nand U26355 (N_26355,N_24477,N_22838);
or U26356 (N_26356,N_20223,N_22884);
nor U26357 (N_26357,N_22182,N_23532);
nand U26358 (N_26358,N_21207,N_22248);
nor U26359 (N_26359,N_22316,N_20696);
xnor U26360 (N_26360,N_22746,N_23604);
nand U26361 (N_26361,N_23938,N_21509);
nor U26362 (N_26362,N_21739,N_20399);
or U26363 (N_26363,N_23485,N_24594);
and U26364 (N_26364,N_21910,N_23957);
nor U26365 (N_26365,N_20871,N_24466);
or U26366 (N_26366,N_22008,N_21665);
nand U26367 (N_26367,N_22699,N_21338);
xnor U26368 (N_26368,N_23033,N_24170);
and U26369 (N_26369,N_24290,N_24006);
or U26370 (N_26370,N_21965,N_20534);
or U26371 (N_26371,N_23246,N_23337);
and U26372 (N_26372,N_24507,N_23691);
nor U26373 (N_26373,N_20409,N_22059);
nor U26374 (N_26374,N_24232,N_21044);
xor U26375 (N_26375,N_22424,N_22558);
and U26376 (N_26376,N_24584,N_22461);
and U26377 (N_26377,N_24535,N_23154);
nor U26378 (N_26378,N_23106,N_21083);
xor U26379 (N_26379,N_22636,N_22475);
nor U26380 (N_26380,N_22589,N_20964);
nand U26381 (N_26381,N_20982,N_22141);
and U26382 (N_26382,N_20308,N_20358);
nand U26383 (N_26383,N_21705,N_22990);
xnor U26384 (N_26384,N_20830,N_24985);
nor U26385 (N_26385,N_24510,N_21330);
xor U26386 (N_26386,N_22815,N_23208);
nand U26387 (N_26387,N_20719,N_21178);
and U26388 (N_26388,N_20314,N_21653);
and U26389 (N_26389,N_24748,N_22755);
nor U26390 (N_26390,N_23213,N_21532);
nor U26391 (N_26391,N_24610,N_23822);
or U26392 (N_26392,N_24735,N_22386);
xor U26393 (N_26393,N_20102,N_22410);
or U26394 (N_26394,N_24641,N_20039);
nor U26395 (N_26395,N_24369,N_23173);
and U26396 (N_26396,N_21597,N_21831);
and U26397 (N_26397,N_21808,N_23926);
nor U26398 (N_26398,N_21139,N_22113);
nor U26399 (N_26399,N_22099,N_24605);
nor U26400 (N_26400,N_23022,N_23277);
and U26401 (N_26401,N_24530,N_24726);
nand U26402 (N_26402,N_21720,N_24030);
nor U26403 (N_26403,N_21418,N_23830);
and U26404 (N_26404,N_20953,N_24738);
nor U26405 (N_26405,N_22490,N_22961);
and U26406 (N_26406,N_23276,N_22987);
or U26407 (N_26407,N_21764,N_20811);
nand U26408 (N_26408,N_24574,N_24111);
and U26409 (N_26409,N_24155,N_22643);
and U26410 (N_26410,N_20000,N_20233);
and U26411 (N_26411,N_23969,N_23226);
xnor U26412 (N_26412,N_20634,N_21662);
and U26413 (N_26413,N_20482,N_20682);
or U26414 (N_26414,N_23393,N_24962);
nand U26415 (N_26415,N_24598,N_21548);
or U26416 (N_26416,N_22294,N_21607);
nand U26417 (N_26417,N_21401,N_20755);
or U26418 (N_26418,N_23191,N_21555);
nand U26419 (N_26419,N_23294,N_24768);
nor U26420 (N_26420,N_20574,N_23421);
xor U26421 (N_26421,N_21975,N_21245);
nand U26422 (N_26422,N_21234,N_24104);
nor U26423 (N_26423,N_22358,N_21704);
and U26424 (N_26424,N_22364,N_21953);
nand U26425 (N_26425,N_24139,N_20406);
nor U26426 (N_26426,N_20621,N_22715);
and U26427 (N_26427,N_22325,N_24740);
nand U26428 (N_26428,N_20722,N_24665);
and U26429 (N_26429,N_20408,N_21904);
and U26430 (N_26430,N_22479,N_21020);
and U26431 (N_26431,N_23390,N_20610);
nand U26432 (N_26432,N_22606,N_24277);
and U26433 (N_26433,N_21259,N_21233);
nor U26434 (N_26434,N_20457,N_23661);
and U26435 (N_26435,N_20645,N_24453);
nand U26436 (N_26436,N_24018,N_22185);
nand U26437 (N_26437,N_24345,N_24385);
and U26438 (N_26438,N_24997,N_23901);
and U26439 (N_26439,N_24243,N_21033);
and U26440 (N_26440,N_21530,N_20841);
or U26441 (N_26441,N_22303,N_23779);
nor U26442 (N_26442,N_21800,N_22074);
and U26443 (N_26443,N_22959,N_22090);
or U26444 (N_26444,N_23146,N_20446);
nand U26445 (N_26445,N_20359,N_24233);
or U26446 (N_26446,N_23460,N_24820);
nor U26447 (N_26447,N_24312,N_21237);
and U26448 (N_26448,N_23805,N_22445);
nand U26449 (N_26449,N_20737,N_20017);
xnor U26450 (N_26450,N_22900,N_20245);
nor U26451 (N_26451,N_24156,N_22906);
and U26452 (N_26452,N_23461,N_20501);
nor U26453 (N_26453,N_20862,N_24209);
nand U26454 (N_26454,N_23509,N_24457);
nand U26455 (N_26455,N_22168,N_20061);
and U26456 (N_26456,N_21821,N_23551);
xor U26457 (N_26457,N_23413,N_23837);
nand U26458 (N_26458,N_20254,N_24478);
nor U26459 (N_26459,N_22203,N_24000);
and U26460 (N_26460,N_24796,N_20957);
xor U26461 (N_26461,N_20302,N_22320);
and U26462 (N_26462,N_23725,N_22683);
and U26463 (N_26463,N_22024,N_24799);
nand U26464 (N_26464,N_24706,N_22574);
or U26465 (N_26465,N_22260,N_21478);
xor U26466 (N_26466,N_22672,N_24019);
nand U26467 (N_26467,N_21174,N_20562);
nor U26468 (N_26468,N_23350,N_20054);
xnor U26469 (N_26469,N_24956,N_24912);
nand U26470 (N_26470,N_24532,N_22660);
and U26471 (N_26471,N_24603,N_22408);
or U26472 (N_26472,N_23863,N_21013);
or U26473 (N_26473,N_21903,N_23319);
xor U26474 (N_26474,N_21361,N_20708);
xor U26475 (N_26475,N_21988,N_20029);
or U26476 (N_26476,N_21722,N_23013);
nor U26477 (N_26477,N_20775,N_21493);
or U26478 (N_26478,N_24987,N_21618);
nor U26479 (N_26479,N_21840,N_24146);
or U26480 (N_26480,N_24245,N_20734);
nor U26481 (N_26481,N_23470,N_22994);
nand U26482 (N_26482,N_24993,N_23090);
nor U26483 (N_26483,N_20037,N_23593);
xor U26484 (N_26484,N_23056,N_23906);
nor U26485 (N_26485,N_23795,N_23441);
and U26486 (N_26486,N_21527,N_22275);
nand U26487 (N_26487,N_20831,N_21422);
xnor U26488 (N_26488,N_21192,N_23702);
nand U26489 (N_26489,N_21674,N_22954);
nand U26490 (N_26490,N_22754,N_24131);
nand U26491 (N_26491,N_22179,N_20961);
nor U26492 (N_26492,N_24747,N_24698);
xnor U26493 (N_26493,N_21855,N_24090);
nor U26494 (N_26494,N_24774,N_24497);
and U26495 (N_26495,N_22601,N_22520);
and U26496 (N_26496,N_20280,N_23814);
or U26497 (N_26497,N_21265,N_23870);
or U26498 (N_26498,N_23801,N_20618);
xor U26499 (N_26499,N_20038,N_24742);
or U26500 (N_26500,N_22375,N_20462);
or U26501 (N_26501,N_20230,N_21508);
nor U26502 (N_26502,N_22314,N_24262);
xor U26503 (N_26503,N_22867,N_20449);
or U26504 (N_26504,N_20465,N_21480);
nand U26505 (N_26505,N_22457,N_20048);
xor U26506 (N_26506,N_20865,N_21805);
nand U26507 (N_26507,N_21512,N_22108);
or U26508 (N_26508,N_21190,N_21763);
xor U26509 (N_26509,N_23985,N_24416);
or U26510 (N_26510,N_22057,N_22144);
and U26511 (N_26511,N_24707,N_24830);
or U26512 (N_26512,N_24501,N_20448);
nor U26513 (N_26513,N_23388,N_24324);
nor U26514 (N_26514,N_20956,N_21881);
or U26515 (N_26515,N_22007,N_24745);
nand U26516 (N_26516,N_23259,N_24469);
xor U26517 (N_26517,N_20895,N_23614);
xor U26518 (N_26518,N_24310,N_24763);
nor U26519 (N_26519,N_21628,N_24922);
nor U26520 (N_26520,N_20004,N_22062);
nand U26521 (N_26521,N_21326,N_22793);
nor U26522 (N_26522,N_20701,N_20536);
xnor U26523 (N_26523,N_20174,N_23450);
or U26524 (N_26524,N_24413,N_24591);
nor U26525 (N_26525,N_21993,N_21585);
nand U26526 (N_26526,N_22788,N_20432);
nor U26527 (N_26527,N_24449,N_24447);
nand U26528 (N_26528,N_20915,N_22153);
nor U26529 (N_26529,N_23230,N_23964);
or U26530 (N_26530,N_20453,N_23808);
nor U26531 (N_26531,N_22469,N_24617);
nor U26532 (N_26532,N_23873,N_22835);
nand U26533 (N_26533,N_21864,N_22942);
nand U26534 (N_26534,N_22766,N_20299);
nor U26535 (N_26535,N_23709,N_24208);
nand U26536 (N_26536,N_20512,N_24124);
nor U26537 (N_26537,N_23911,N_20296);
or U26538 (N_26538,N_24278,N_21082);
and U26539 (N_26539,N_23044,N_22365);
and U26540 (N_26540,N_20024,N_22350);
nand U26541 (N_26541,N_22800,N_21684);
or U26542 (N_26542,N_21707,N_22146);
nand U26543 (N_26543,N_24935,N_23111);
or U26544 (N_26544,N_24546,N_22725);
xor U26545 (N_26545,N_21740,N_20431);
nor U26546 (N_26546,N_24528,N_21331);
nand U26547 (N_26547,N_22120,N_20891);
xnor U26548 (N_26548,N_21795,N_20275);
nand U26549 (N_26549,N_22034,N_22973);
or U26550 (N_26550,N_20198,N_23986);
nand U26551 (N_26551,N_20100,N_21457);
nor U26552 (N_26552,N_24399,N_20514);
nand U26553 (N_26553,N_22352,N_20082);
or U26554 (N_26554,N_20632,N_21291);
nand U26555 (N_26555,N_24207,N_20318);
nor U26556 (N_26556,N_23451,N_21957);
xor U26557 (N_26557,N_23423,N_24195);
and U26558 (N_26558,N_21107,N_20859);
and U26559 (N_26559,N_22382,N_21025);
nand U26560 (N_26560,N_21728,N_23296);
nor U26561 (N_26561,N_22927,N_24710);
xor U26562 (N_26562,N_23404,N_20843);
or U26563 (N_26563,N_21341,N_23712);
and U26564 (N_26564,N_20320,N_22582);
nand U26565 (N_26565,N_21506,N_24909);
nand U26566 (N_26566,N_23241,N_22337);
or U26567 (N_26567,N_20551,N_23726);
nor U26568 (N_26568,N_23179,N_21880);
or U26569 (N_26569,N_22043,N_20372);
xnor U26570 (N_26570,N_22865,N_21819);
and U26571 (N_26571,N_22952,N_24079);
xnor U26572 (N_26572,N_23843,N_24490);
and U26573 (N_26573,N_20892,N_23118);
nand U26574 (N_26574,N_22331,N_24759);
and U26575 (N_26575,N_21420,N_22921);
xor U26576 (N_26576,N_24394,N_24553);
or U26577 (N_26577,N_23695,N_21811);
nor U26578 (N_26578,N_23746,N_21600);
or U26579 (N_26579,N_20436,N_23980);
xnor U26580 (N_26580,N_23099,N_22645);
and U26581 (N_26581,N_21529,N_22962);
and U26582 (N_26582,N_20656,N_20067);
nor U26583 (N_26583,N_24825,N_20790);
xnor U26584 (N_26584,N_21955,N_22278);
xnor U26585 (N_26585,N_20131,N_22280);
xor U26586 (N_26586,N_20478,N_22911);
nor U26587 (N_26587,N_22166,N_21837);
xnor U26588 (N_26588,N_22839,N_22347);
and U26589 (N_26589,N_22696,N_20826);
or U26590 (N_26590,N_21954,N_21011);
nand U26591 (N_26591,N_23872,N_20698);
xor U26592 (N_26592,N_22326,N_21507);
xor U26593 (N_26593,N_24570,N_23806);
nand U26594 (N_26594,N_23074,N_21989);
or U26595 (N_26595,N_23222,N_20276);
xor U26596 (N_26596,N_24647,N_22467);
nor U26597 (N_26597,N_20312,N_23244);
nor U26598 (N_26598,N_21599,N_20119);
nand U26599 (N_26599,N_21611,N_21511);
nand U26600 (N_26600,N_21920,N_24110);
nand U26601 (N_26601,N_23125,N_23199);
xor U26602 (N_26602,N_23859,N_20050);
and U26603 (N_26603,N_20797,N_22878);
and U26604 (N_26604,N_23320,N_23433);
nand U26605 (N_26605,N_24806,N_22026);
and U26606 (N_26606,N_24531,N_22567);
or U26607 (N_26607,N_21644,N_22249);
xor U26608 (N_26608,N_22258,N_21950);
xnor U26609 (N_26609,N_22997,N_20178);
or U26610 (N_26610,N_23190,N_21990);
xor U26611 (N_26611,N_22361,N_21991);
nand U26612 (N_26612,N_20328,N_24038);
xnor U26613 (N_26613,N_23800,N_23945);
nand U26614 (N_26614,N_22308,N_23879);
xnor U26615 (N_26615,N_20357,N_23153);
or U26616 (N_26616,N_21568,N_24418);
or U26617 (N_26617,N_24499,N_23685);
xnor U26618 (N_26618,N_23278,N_21817);
or U26619 (N_26619,N_20916,N_21977);
nand U26620 (N_26620,N_23550,N_24313);
nor U26621 (N_26621,N_21586,N_22416);
nor U26622 (N_26622,N_20993,N_20077);
nor U26623 (N_26623,N_24297,N_22252);
nor U26624 (N_26624,N_24182,N_20444);
nand U26625 (N_26625,N_24723,N_24303);
xnor U26626 (N_26626,N_20941,N_21936);
nand U26627 (N_26627,N_20384,N_20732);
nor U26628 (N_26628,N_23874,N_24200);
and U26629 (N_26629,N_22627,N_21883);
nand U26630 (N_26630,N_20780,N_22134);
or U26631 (N_26631,N_24360,N_20817);
and U26632 (N_26632,N_20485,N_23382);
xor U26633 (N_26633,N_22131,N_20782);
nand U26634 (N_26634,N_23123,N_23414);
nor U26635 (N_26635,N_20590,N_20999);
and U26636 (N_26636,N_23812,N_20339);
and U26637 (N_26637,N_23524,N_21272);
xor U26638 (N_26638,N_22526,N_21875);
xor U26639 (N_26639,N_24633,N_23765);
nor U26640 (N_26640,N_24365,N_22680);
nor U26641 (N_26641,N_22250,N_20265);
or U26642 (N_26642,N_24582,N_24761);
and U26643 (N_26643,N_23437,N_20287);
nand U26644 (N_26644,N_23027,N_21271);
nor U26645 (N_26645,N_21376,N_22919);
and U26646 (N_26646,N_24864,N_24355);
or U26647 (N_26647,N_23897,N_20237);
or U26648 (N_26648,N_21276,N_20493);
nand U26649 (N_26649,N_22264,N_23232);
or U26650 (N_26650,N_21467,N_22224);
and U26651 (N_26651,N_23531,N_21574);
nand U26652 (N_26652,N_23345,N_22159);
and U26653 (N_26653,N_20120,N_21040);
xor U26654 (N_26654,N_23760,N_21734);
nor U26655 (N_26655,N_22257,N_21660);
or U26656 (N_26656,N_20825,N_21202);
nand U26657 (N_26657,N_20425,N_24382);
nand U26658 (N_26658,N_21833,N_20182);
or U26659 (N_26659,N_23580,N_21123);
or U26660 (N_26660,N_22213,N_20370);
nand U26661 (N_26661,N_20400,N_21563);
or U26662 (N_26662,N_24929,N_23144);
and U26663 (N_26663,N_22794,N_24508);
nor U26664 (N_26664,N_21346,N_24268);
nand U26665 (N_26665,N_24645,N_24109);
nand U26666 (N_26666,N_24395,N_23753);
or U26667 (N_26667,N_22329,N_24681);
xnor U26668 (N_26668,N_20337,N_22701);
or U26669 (N_26669,N_24149,N_23112);
nor U26670 (N_26670,N_20777,N_21404);
xnor U26671 (N_26671,N_20264,N_24204);
nand U26672 (N_26672,N_21565,N_23999);
nand U26673 (N_26673,N_23684,N_23956);
nand U26674 (N_26674,N_20135,N_22820);
xnor U26675 (N_26675,N_20697,N_22180);
and U26676 (N_26676,N_21454,N_21929);
nand U26677 (N_26677,N_23121,N_24919);
xnor U26678 (N_26678,N_24462,N_20025);
and U26679 (N_26679,N_20225,N_24875);
xnor U26680 (N_26680,N_24273,N_21985);
nand U26681 (N_26681,N_24434,N_24271);
xnor U26682 (N_26682,N_24612,N_22964);
xor U26683 (N_26683,N_23847,N_23936);
and U26684 (N_26684,N_23358,N_23409);
xnor U26685 (N_26685,N_24854,N_22784);
xor U26686 (N_26686,N_21608,N_24203);
and U26687 (N_26687,N_22030,N_22064);
or U26688 (N_26688,N_21089,N_21745);
nand U26689 (N_26689,N_21096,N_23250);
xnor U26690 (N_26690,N_20819,N_23030);
xnor U26691 (N_26691,N_24081,N_24916);
xor U26692 (N_26692,N_20289,N_24861);
xnor U26693 (N_26693,N_23523,N_22374);
nor U26694 (N_26694,N_24873,N_20226);
nand U26695 (N_26695,N_23671,N_24589);
and U26696 (N_26696,N_24191,N_21410);
xnor U26697 (N_26697,N_23982,N_23176);
and U26698 (N_26698,N_20545,N_20146);
or U26699 (N_26699,N_21569,N_22406);
nor U26700 (N_26700,N_20752,N_21663);
xnor U26701 (N_26701,N_22688,N_24249);
nand U26702 (N_26702,N_22229,N_24005);
nor U26703 (N_26703,N_22768,N_20164);
xnor U26704 (N_26704,N_22870,N_22851);
or U26705 (N_26705,N_20197,N_24328);
xnor U26706 (N_26706,N_20452,N_22197);
nor U26707 (N_26707,N_24727,N_20271);
nor U26708 (N_26708,N_24251,N_20827);
nand U26709 (N_26709,N_22448,N_23599);
nand U26710 (N_26710,N_23920,N_23038);
or U26711 (N_26711,N_22741,N_24426);
or U26712 (N_26712,N_23231,N_24649);
nor U26713 (N_26713,N_24808,N_20833);
or U26714 (N_26714,N_20913,N_22515);
and U26715 (N_26715,N_23346,N_22472);
xor U26716 (N_26716,N_23505,N_20902);
or U26717 (N_26717,N_22553,N_24525);
and U26718 (N_26718,N_20533,N_22251);
or U26719 (N_26719,N_21094,N_21226);
nand U26720 (N_26720,N_23046,N_21726);
nand U26721 (N_26721,N_22783,N_22685);
nand U26722 (N_26722,N_22651,N_24867);
xor U26723 (N_26723,N_23486,N_21652);
nor U26724 (N_26724,N_24341,N_20523);
nand U26725 (N_26725,N_21434,N_22016);
nor U26726 (N_26726,N_20382,N_23284);
nand U26727 (N_26727,N_21218,N_22595);
nand U26728 (N_26728,N_20721,N_21008);
xnor U26729 (N_26729,N_23204,N_21760);
and U26730 (N_26730,N_21363,N_23898);
nor U26731 (N_26731,N_20085,N_23637);
xor U26732 (N_26732,N_21124,N_23696);
and U26733 (N_26733,N_20515,N_23002);
nor U26734 (N_26734,N_20652,N_22629);
nand U26735 (N_26735,N_24353,N_20199);
nand U26736 (N_26736,N_24713,N_24202);
or U26737 (N_26737,N_21930,N_22590);
and U26738 (N_26738,N_20655,N_20343);
or U26739 (N_26739,N_24009,N_23387);
xnor U26740 (N_26740,N_22431,N_23996);
or U26741 (N_26741,N_20693,N_23592);
nor U26742 (N_26742,N_24422,N_24439);
or U26743 (N_26743,N_20930,N_23062);
xor U26744 (N_26744,N_21375,N_23557);
or U26745 (N_26745,N_20664,N_24718);
nand U26746 (N_26746,N_24839,N_23623);
nand U26747 (N_26747,N_23214,N_23392);
nor U26748 (N_26748,N_20434,N_23047);
and U26749 (N_26749,N_24973,N_24545);
or U26750 (N_26750,N_24154,N_22591);
nand U26751 (N_26751,N_24384,N_21724);
or U26752 (N_26752,N_21377,N_22414);
nor U26753 (N_26753,N_20259,N_20837);
nor U26754 (N_26754,N_21496,N_24961);
nor U26755 (N_26755,N_24702,N_24944);
nor U26756 (N_26756,N_24337,N_21858);
nand U26757 (N_26757,N_22972,N_22984);
nor U26758 (N_26758,N_22519,N_24816);
or U26759 (N_26759,N_21676,N_22992);
nand U26760 (N_26760,N_23281,N_23697);
nor U26761 (N_26761,N_23836,N_21489);
nand U26762 (N_26762,N_21445,N_23758);
and U26763 (N_26763,N_23579,N_20142);
and U26764 (N_26764,N_23511,N_22458);
nand U26765 (N_26765,N_23081,N_20123);
nor U26766 (N_26766,N_20491,N_20397);
or U26767 (N_26767,N_22890,N_24538);
nand U26768 (N_26768,N_21026,N_23200);
or U26769 (N_26769,N_22044,N_24460);
nor U26770 (N_26770,N_21381,N_21613);
or U26771 (N_26771,N_23361,N_24853);
or U26772 (N_26772,N_22028,N_22124);
nor U26773 (N_26773,N_24254,N_24870);
nand U26774 (N_26774,N_24397,N_21504);
and U26775 (N_26775,N_20291,N_23990);
nor U26776 (N_26776,N_23024,N_23976);
or U26777 (N_26777,N_24930,N_21312);
and U26778 (N_26778,N_23443,N_23569);
and U26779 (N_26779,N_22060,N_22664);
xnor U26780 (N_26780,N_24407,N_24272);
and U26781 (N_26781,N_23224,N_22560);
or U26782 (N_26782,N_22669,N_20936);
nand U26783 (N_26783,N_22470,N_21519);
and U26784 (N_26784,N_21057,N_24210);
nand U26785 (N_26785,N_24669,N_20894);
nand U26786 (N_26786,N_21627,N_24375);
nor U26787 (N_26787,N_20486,N_22712);
xnor U26788 (N_26788,N_20849,N_22714);
nand U26789 (N_26789,N_20582,N_21832);
and U26790 (N_26790,N_20552,N_20538);
nor U26791 (N_26791,N_23122,N_22181);
or U26792 (N_26792,N_21001,N_24643);
nand U26793 (N_26793,N_20414,N_23161);
and U26794 (N_26794,N_20771,N_23066);
nand U26795 (N_26795,N_21725,N_21208);
or U26796 (N_26796,N_21282,N_20003);
xnor U26797 (N_26797,N_22353,N_21900);
xor U26798 (N_26798,N_20663,N_20601);
or U26799 (N_26799,N_23206,N_22963);
xor U26800 (N_26800,N_20228,N_22004);
nor U26801 (N_26801,N_22482,N_23745);
nand U26802 (N_26802,N_20470,N_20835);
xnor U26803 (N_26803,N_21697,N_24890);
and U26804 (N_26804,N_22849,N_24631);
or U26805 (N_26805,N_22466,N_20528);
and U26806 (N_26806,N_24461,N_22165);
or U26807 (N_26807,N_22199,N_22823);
and U26808 (N_26808,N_20625,N_21405);
nand U26809 (N_26809,N_22549,N_20076);
xor U26810 (N_26810,N_21554,N_20641);
nor U26811 (N_26811,N_22706,N_23952);
xor U26812 (N_26812,N_22883,N_24236);
or U26813 (N_26813,N_21022,N_23626);
or U26814 (N_26814,N_23209,N_23132);
nand U26815 (N_26815,N_20413,N_22373);
nand U26816 (N_26816,N_22819,N_23156);
or U26817 (N_26817,N_20854,N_24613);
or U26818 (N_26818,N_24756,N_21796);
or U26819 (N_26819,N_22598,N_20011);
nor U26820 (N_26820,N_23087,N_21654);
xnor U26821 (N_26821,N_21472,N_20158);
xnor U26822 (N_26822,N_21657,N_24465);
xnor U26823 (N_26823,N_22380,N_24992);
xor U26824 (N_26824,N_22454,N_24845);
and U26825 (N_26825,N_23223,N_23853);
xnor U26826 (N_26826,N_21438,N_22610);
nand U26827 (N_26827,N_20887,N_21517);
and U26828 (N_26828,N_23854,N_21128);
xnor U26829 (N_26829,N_20368,N_21053);
nand U26830 (N_26830,N_22171,N_23882);
or U26831 (N_26831,N_21308,N_20531);
and U26832 (N_26832,N_21256,N_24620);
nand U26833 (N_26833,N_24168,N_22348);
xnor U26834 (N_26834,N_23528,N_20023);
or U26835 (N_26835,N_23510,N_22032);
xnor U26836 (N_26836,N_21068,N_20700);
or U26837 (N_26837,N_20013,N_21786);
nor U26838 (N_26838,N_21452,N_22133);
or U26839 (N_26839,N_24795,N_20473);
xor U26840 (N_26840,N_24902,N_22539);
or U26841 (N_26841,N_24336,N_20490);
xor U26842 (N_26842,N_21947,N_24583);
xnor U26843 (N_26843,N_23138,N_20669);
or U26844 (N_26844,N_24431,N_24287);
or U26845 (N_26845,N_21830,N_22536);
xnor U26846 (N_26846,N_22206,N_21052);
or U26847 (N_26847,N_23036,N_20179);
and U26848 (N_26848,N_20670,N_20875);
or U26849 (N_26849,N_20542,N_20995);
nand U26850 (N_26850,N_23235,N_22790);
and U26851 (N_26851,N_22334,N_20581);
nand U26852 (N_26852,N_24565,N_23493);
xnor U26853 (N_26853,N_22094,N_22653);
or U26854 (N_26854,N_20555,N_20627);
nand U26855 (N_26855,N_20335,N_21236);
nand U26856 (N_26856,N_21255,N_21311);
nor U26857 (N_26857,N_23496,N_20239);
nand U26858 (N_26858,N_24346,N_22845);
xnor U26859 (N_26859,N_21130,N_20786);
xor U26860 (N_26860,N_23722,N_24753);
nor U26861 (N_26861,N_20727,N_23899);
and U26862 (N_26862,N_23790,N_20203);
nor U26863 (N_26863,N_20053,N_21678);
nand U26864 (N_26864,N_22531,N_21416);
or U26865 (N_26865,N_23311,N_24265);
and U26866 (N_26866,N_24106,N_23189);
or U26867 (N_26867,N_23838,N_23410);
or U26868 (N_26868,N_21000,N_22393);
or U26869 (N_26869,N_20286,N_23921);
nor U26870 (N_26870,N_22859,N_21090);
or U26871 (N_26871,N_21581,N_21813);
or U26872 (N_26872,N_22112,N_20778);
and U26873 (N_26873,N_23447,N_20219);
or U26874 (N_26874,N_24621,N_20860);
nor U26875 (N_26875,N_20445,N_22702);
or U26876 (N_26876,N_22810,N_21473);
or U26877 (N_26877,N_22753,N_24281);
nand U26878 (N_26878,N_20014,N_20608);
nand U26879 (N_26879,N_24468,N_23116);
nor U26880 (N_26880,N_22773,N_20117);
or U26881 (N_26881,N_23932,N_20929);
xnor U26882 (N_26882,N_20170,N_22121);
and U26883 (N_26883,N_24444,N_23343);
nor U26884 (N_26884,N_21374,N_24450);
xor U26885 (N_26885,N_20668,N_23166);
xnor U26886 (N_26886,N_23989,N_22052);
nand U26887 (N_26887,N_21369,N_24267);
and U26888 (N_26888,N_21867,N_22396);
or U26889 (N_26889,N_23251,N_23425);
nor U26890 (N_26890,N_24872,N_23113);
xnor U26891 (N_26891,N_23961,N_21545);
and U26892 (N_26892,N_20020,N_20258);
nand U26893 (N_26893,N_24488,N_22716);
nand U26894 (N_26894,N_24458,N_22162);
nand U26895 (N_26895,N_24174,N_23197);
nor U26896 (N_26896,N_21168,N_23878);
nand U26897 (N_26897,N_24587,N_24666);
or U26898 (N_26898,N_23477,N_21339);
nor U26899 (N_26899,N_22827,N_23152);
nor U26900 (N_26900,N_21327,N_20918);
nand U26901 (N_26901,N_22860,N_23734);
and U26902 (N_26902,N_24569,N_21423);
or U26903 (N_26903,N_20513,N_23565);
or U26904 (N_26904,N_24561,N_23965);
nand U26905 (N_26905,N_22430,N_23307);
xnor U26906 (N_26906,N_24921,N_24874);
nor U26907 (N_26907,N_20180,N_22791);
and U26908 (N_26908,N_22272,N_20398);
or U26909 (N_26909,N_22155,N_23738);
and U26910 (N_26910,N_20354,N_24144);
xnor U26911 (N_26911,N_22048,N_24430);
and U26912 (N_26912,N_20113,N_22578);
nand U26913 (N_26913,N_20090,N_23050);
nand U26914 (N_26914,N_20395,N_21135);
and U26915 (N_26915,N_20651,N_21714);
nor U26916 (N_26916,N_22694,N_20741);
nand U26917 (N_26917,N_24769,N_20325);
nand U26918 (N_26918,N_24178,N_20151);
and U26919 (N_26919,N_21797,N_22253);
and U26920 (N_26920,N_23218,N_22456);
nand U26921 (N_26921,N_21140,N_24941);
nand U26922 (N_26922,N_22618,N_24012);
nand U26923 (N_26923,N_22039,N_24475);
nor U26924 (N_26924,N_24077,N_22063);
nand U26925 (N_26925,N_23233,N_20147);
xor U26926 (N_26926,N_21014,N_23977);
or U26927 (N_26927,N_20263,N_23373);
xor U26928 (N_26928,N_24276,N_21055);
nand U26929 (N_26929,N_20644,N_23967);
nand U26930 (N_26930,N_22438,N_22080);
nand U26931 (N_26931,N_24838,N_22756);
nand U26932 (N_26932,N_21869,N_24459);
nand U26933 (N_26933,N_21297,N_22926);
nor U26934 (N_26934,N_22403,N_23914);
and U26935 (N_26935,N_22061,N_24781);
nor U26936 (N_26936,N_22081,N_23828);
or U26937 (N_26937,N_24184,N_20108);
nand U26938 (N_26938,N_21887,N_21601);
nor U26939 (N_26939,N_20475,N_20949);
and U26940 (N_26940,N_20504,N_21413);
and U26941 (N_26941,N_24835,N_21372);
nand U26942 (N_26942,N_24087,N_21219);
nand U26943 (N_26943,N_21551,N_23366);
nand U26944 (N_26944,N_23412,N_20508);
nand U26945 (N_26945,N_22281,N_23297);
and U26946 (N_26946,N_21531,N_23759);
and U26947 (N_26947,N_20838,N_20418);
xor U26948 (N_26948,N_24655,N_20238);
or U26949 (N_26949,N_24865,N_20899);
nor U26950 (N_26950,N_21853,N_24047);
and U26951 (N_26951,N_22561,N_20162);
and U26952 (N_26952,N_24951,N_20762);
nand U26953 (N_26953,N_24388,N_21429);
and U26954 (N_26954,N_22564,N_24554);
or U26955 (N_26955,N_24089,N_20443);
nand U26956 (N_26956,N_23992,N_21391);
nand U26957 (N_26957,N_23653,N_21637);
xnor U26958 (N_26958,N_23092,N_23312);
xor U26959 (N_26959,N_22862,N_24682);
xor U26960 (N_26960,N_23699,N_23913);
nor U26961 (N_26961,N_22974,N_22692);
xnor U26962 (N_26962,N_20344,N_22513);
or U26963 (N_26963,N_20544,N_20906);
nor U26964 (N_26964,N_24221,N_21609);
nor U26965 (N_26965,N_21152,N_22235);
nor U26966 (N_26966,N_21303,N_20112);
nor U26967 (N_26967,N_22948,N_20019);
nand U26968 (N_26968,N_24882,N_23057);
nand U26969 (N_26969,N_23229,N_24405);
nand U26970 (N_26970,N_23474,N_20172);
xor U26971 (N_26971,N_21854,N_20662);
xnor U26972 (N_26972,N_21477,N_20965);
and U26973 (N_26973,N_24371,N_22776);
and U26974 (N_26974,N_24812,N_22328);
nand U26975 (N_26975,N_23274,N_21076);
nor U26976 (N_26976,N_24931,N_22372);
or U26977 (N_26977,N_24608,N_21148);
nor U26978 (N_26978,N_22072,N_24575);
nor U26979 (N_26979,N_21562,N_24137);
nor U26980 (N_26980,N_24040,N_24547);
nor U26981 (N_26981,N_24275,N_20783);
nand U26982 (N_26982,N_20522,N_21200);
and U26983 (N_26983,N_23767,N_21732);
nand U26984 (N_26984,N_24664,N_22743);
and U26985 (N_26985,N_23436,N_22812);
and U26986 (N_26986,N_21415,N_23004);
nand U26987 (N_26987,N_24957,N_23549);
xor U26988 (N_26988,N_23043,N_23015);
nor U26989 (N_26989,N_22101,N_23072);
nor U26990 (N_26990,N_24330,N_21802);
nor U26991 (N_26991,N_22351,N_22172);
or U26992 (N_26992,N_20480,N_22276);
xor U26993 (N_26993,N_21579,N_24420);
xnor U26994 (N_26994,N_22332,N_24504);
xor U26995 (N_26995,N_21177,N_24176);
and U26996 (N_26996,N_23500,N_22950);
nor U26997 (N_26997,N_22447,N_24662);
nand U26998 (N_26998,N_22693,N_20295);
xor U26999 (N_26999,N_21007,N_24848);
or U27000 (N_27000,N_24797,N_21246);
xor U27001 (N_27001,N_24984,N_24419);
xnor U27002 (N_27002,N_23378,N_20105);
and U27003 (N_27003,N_23064,N_23768);
and U27004 (N_27004,N_23368,N_24737);
xor U27005 (N_27005,N_23688,N_22728);
nor U27006 (N_27006,N_22966,N_21321);
nand U27007 (N_27007,N_22894,N_21161);
nand U27008 (N_27008,N_22749,N_23293);
and U27009 (N_27009,N_20468,N_24066);
nor U27010 (N_27010,N_22944,N_23833);
nor U27011 (N_27011,N_23727,N_21979);
nand U27012 (N_27012,N_20800,N_20305);
nor U27013 (N_27013,N_21866,N_22562);
xor U27014 (N_27014,N_23521,N_24751);
or U27015 (N_27015,N_24321,N_21292);
and U27016 (N_27016,N_24318,N_24625);
nand U27017 (N_27017,N_24868,N_22731);
nand U27018 (N_27018,N_24084,N_20998);
nand U27019 (N_27019,N_23834,N_23730);
and U27020 (N_27020,N_21144,N_21578);
or U27021 (N_27021,N_20366,N_23591);
nand U27022 (N_27022,N_20667,N_24991);
nor U27023 (N_27023,N_24179,N_20171);
or U27024 (N_27024,N_22298,N_20973);
xnor U27025 (N_27025,N_23953,N_21938);
xor U27026 (N_27026,N_24862,N_22774);
or U27027 (N_27027,N_23073,N_23572);
xnor U27028 (N_27028,N_21388,N_24679);
nand U27029 (N_27029,N_21284,N_23495);
xor U27030 (N_27030,N_22532,N_22988);
nor U27031 (N_27031,N_21612,N_22401);
nand U27032 (N_27032,N_20202,N_20153);
xor U27033 (N_27033,N_23915,N_22613);
and U27034 (N_27034,N_21915,N_20985);
nand U27035 (N_27035,N_21567,N_24893);
and U27036 (N_27036,N_21655,N_24096);
nand U27037 (N_27037,N_24119,N_20348);
nand U27038 (N_27038,N_22828,N_22745);
nor U27039 (N_27039,N_23811,N_23061);
and U27040 (N_27040,N_21687,N_21913);
or U27041 (N_27041,N_22449,N_22237);
nand U27042 (N_27042,N_22816,N_24943);
or U27043 (N_27043,N_23884,N_20500);
or U27044 (N_27044,N_20882,N_20539);
nor U27045 (N_27045,N_20185,N_22241);
or U27046 (N_27046,N_22362,N_20184);
nand U27047 (N_27047,N_21754,N_20614);
xor U27048 (N_27048,N_20571,N_21097);
nand U27049 (N_27049,N_22689,N_22369);
nand U27050 (N_27050,N_21912,N_24338);
nor U27051 (N_27051,N_21804,N_21675);
xnor U27052 (N_27052,N_20847,N_23975);
nand U27053 (N_27053,N_24592,N_24073);
xor U27054 (N_27054,N_22215,N_23215);
nand U27055 (N_27055,N_21926,N_22566);
or U27056 (N_27056,N_23227,N_21240);
xnor U27057 (N_27057,N_23577,N_23372);
and U27058 (N_27058,N_24198,N_23537);
nand U27059 (N_27059,N_22760,N_21260);
nand U27060 (N_27060,N_20963,N_20810);
xor U27061 (N_27061,N_22427,N_23934);
nor U27062 (N_27062,N_23318,N_21131);
nand U27063 (N_27063,N_20823,N_21584);
and U27064 (N_27064,N_20380,N_23459);
xor U27065 (N_27065,N_23362,N_20643);
and U27066 (N_27066,N_24464,N_24967);
and U27067 (N_27067,N_20152,N_21437);
xor U27068 (N_27068,N_23928,N_21860);
nor U27069 (N_27069,N_22167,N_24130);
xor U27070 (N_27070,N_24054,N_21893);
xnor U27071 (N_27071,N_22556,N_21656);
or U27072 (N_27072,N_24088,N_20868);
or U27073 (N_27073,N_22338,N_22391);
nand U27074 (N_27074,N_22511,N_24122);
nand U27075 (N_27075,N_22437,N_23707);
and U27076 (N_27076,N_22188,N_22644);
nor U27077 (N_27077,N_23424,N_21073);
nor U27078 (N_27078,N_24671,N_21706);
or U27079 (N_27079,N_23000,N_21003);
or U27080 (N_27080,N_23431,N_21789);
and U27081 (N_27081,N_20240,N_20439);
nor U27082 (N_27082,N_24211,N_22452);
or U27083 (N_27083,N_20442,N_21362);
xnor U27084 (N_27084,N_20257,N_24068);
nand U27085 (N_27085,N_23001,N_24334);
xnor U27086 (N_27086,N_23772,N_21828);
or U27087 (N_27087,N_22129,N_24370);
xnor U27088 (N_27088,N_21258,N_22109);
nor U27089 (N_27089,N_20481,N_20774);
and U27090 (N_27090,N_20073,N_20107);
and U27091 (N_27091,N_22544,N_23142);
and U27092 (N_27092,N_22735,N_20553);
and U27093 (N_27093,N_23385,N_20224);
and U27094 (N_27094,N_23997,N_21939);
nor U27095 (N_27095,N_22031,N_20041);
nor U27096 (N_27096,N_24196,N_23025);
and U27097 (N_27097,N_23340,N_20653);
or U27098 (N_27098,N_21692,N_20450);
or U27099 (N_27099,N_22269,N_23520);
nand U27100 (N_27100,N_20294,N_20075);
nand U27101 (N_27101,N_21365,N_20423);
and U27102 (N_27102,N_22371,N_23211);
or U27103 (N_27103,N_22733,N_20292);
nand U27104 (N_27104,N_21299,N_22668);
or U27105 (N_27105,N_20190,N_22750);
nor U27106 (N_27106,N_20818,N_20639);
nand U27107 (N_27107,N_24715,N_24409);
or U27108 (N_27108,N_21857,N_20898);
nand U27109 (N_27109,N_21595,N_21824);
xnor U27110 (N_27110,N_21038,N_20044);
xor U27111 (N_27111,N_20062,N_20391);
nor U27112 (N_27112,N_21294,N_23143);
or U27113 (N_27113,N_20990,N_23035);
nor U27114 (N_27114,N_20832,N_22383);
and U27115 (N_27115,N_20306,N_24331);
or U27116 (N_27116,N_21921,N_20628);
nand U27117 (N_27117,N_20864,N_22633);
nor U27118 (N_27118,N_24162,N_22184);
and U27119 (N_27119,N_24358,N_20836);
xnor U27120 (N_27120,N_24255,N_24112);
xnor U27121 (N_27121,N_24356,N_22488);
nor U27122 (N_27122,N_24361,N_21906);
or U27123 (N_27123,N_24189,N_20496);
and U27124 (N_27124,N_23049,N_21688);
nor U27125 (N_27125,N_23540,N_22076);
xor U27126 (N_27126,N_24022,N_20072);
nor U27127 (N_27127,N_21049,N_24020);
and U27128 (N_27128,N_23902,N_24571);
and U27129 (N_27129,N_23405,N_23445);
and U27130 (N_27130,N_24295,N_22385);
or U27131 (N_27131,N_20086,N_24998);
or U27132 (N_27132,N_22283,N_21060);
nor U27133 (N_27133,N_20499,N_21470);
and U27134 (N_27134,N_23598,N_21093);
nand U27135 (N_27135,N_23160,N_24601);
nand U27136 (N_27136,N_22516,N_23887);
and U27137 (N_27137,N_22572,N_24284);
nand U27138 (N_27138,N_24782,N_22821);
nand U27139 (N_27139,N_21780,N_23787);
nor U27140 (N_27140,N_21759,N_23402);
or U27141 (N_27141,N_20769,N_21919);
or U27142 (N_27142,N_23010,N_24968);
nor U27143 (N_27143,N_21522,N_23667);
nand U27144 (N_27144,N_21141,N_22542);
xor U27145 (N_27145,N_24690,N_20115);
and U27146 (N_27146,N_22871,N_23875);
nand U27147 (N_27147,N_24301,N_23270);
nor U27148 (N_27148,N_21221,N_22483);
and U27149 (N_27149,N_24163,N_23668);
xor U27150 (N_27150,N_22243,N_20680);
or U27151 (N_27151,N_24161,N_24378);
nor U27152 (N_27152,N_21286,N_21112);
nand U27153 (N_27153,N_23140,N_22239);
or U27154 (N_27154,N_20016,N_24120);
nand U27155 (N_27155,N_20717,N_23446);
or U27156 (N_27156,N_22879,N_20474);
and U27157 (N_27157,N_22632,N_22221);
nor U27158 (N_27158,N_22765,N_24958);
and U27159 (N_27159,N_21624,N_22245);
and U27160 (N_27160,N_20888,N_23728);
and U27161 (N_27161,N_22481,N_24298);
nand U27162 (N_27162,N_22157,N_24899);
or U27163 (N_27163,N_20331,N_21332);
xor U27164 (N_27164,N_20231,N_24859);
xnor U27165 (N_27165,N_21188,N_24979);
nand U27166 (N_27166,N_23332,N_24373);
or U27167 (N_27167,N_23672,N_23548);
nor U27168 (N_27168,N_20805,N_22940);
and U27169 (N_27169,N_24234,N_22628);
xnor U27170 (N_27170,N_23506,N_24347);
nor U27171 (N_27171,N_24850,N_24311);
nand U27172 (N_27172,N_20492,N_24618);
nand U27173 (N_27173,N_22309,N_24914);
xnor U27174 (N_27174,N_24072,N_24590);
xnor U27175 (N_27175,N_24435,N_21616);
xnor U27176 (N_27176,N_21019,N_22006);
nor U27177 (N_27177,N_20694,N_20880);
nand U27178 (N_27178,N_21250,N_22191);
or U27179 (N_27179,N_21727,N_20765);
nor U27180 (N_27180,N_24391,N_20813);
nand U27181 (N_27181,N_20713,N_21358);
and U27182 (N_27182,N_20867,N_20098);
or U27183 (N_27183,N_21498,N_23351);
and U27184 (N_27184,N_21846,N_20140);
xnor U27185 (N_27185,N_24760,N_24002);
nor U27186 (N_27186,N_24518,N_23781);
nor U27187 (N_27187,N_20278,N_24443);
xnor U27188 (N_27188,N_21180,N_22763);
xor U27189 (N_27189,N_23633,N_24720);
xnor U27190 (N_27190,N_22149,N_23048);
xnor U27191 (N_27191,N_24061,N_20109);
xor U27192 (N_27192,N_20510,N_23290);
or U27193 (N_27193,N_24194,N_20321);
nor U27194 (N_27194,N_21409,N_23663);
nor U27195 (N_27195,N_22830,N_24071);
or U27196 (N_27196,N_21783,N_24783);
or U27197 (N_27197,N_20594,N_20613);
and U27198 (N_27198,N_22573,N_22527);
nor U27199 (N_27199,N_24300,N_24123);
nor U27200 (N_27200,N_24029,N_23178);
nor U27201 (N_27201,N_24965,N_21591);
xnor U27202 (N_27202,N_21971,N_21481);
or U27203 (N_27203,N_23088,N_21534);
nor U27204 (N_27204,N_21474,N_22318);
nor U27205 (N_27205,N_20591,N_24724);
nor U27206 (N_27206,N_22420,N_20091);
and U27207 (N_27207,N_22345,N_22421);
xnor U27208 (N_27208,N_21444,N_21359);
and U27209 (N_27209,N_24837,N_20101);
or U27210 (N_27210,N_24750,N_24714);
and U27211 (N_27211,N_21718,N_20738);
or U27212 (N_27212,N_24908,N_20742);
nand U27213 (N_27213,N_21646,N_24793);
nor U27214 (N_27214,N_20988,N_24746);
nor U27215 (N_27215,N_20319,N_23285);
nand U27216 (N_27216,N_20948,N_21187);
xnor U27217 (N_27217,N_22852,N_24857);
and U27218 (N_27218,N_24359,N_22429);
nor U27219 (N_27219,N_20586,N_20699);
nand U27220 (N_27220,N_23682,N_22279);
or U27221 (N_27221,N_22711,N_20476);
nand U27222 (N_27222,N_24427,N_20121);
nand U27223 (N_27223,N_21099,N_23789);
xnor U27224 (N_27224,N_22512,N_22596);
xnor U27225 (N_27225,N_22529,N_23063);
nor U27226 (N_27226,N_24947,N_24186);
xnor U27227 (N_27227,N_23187,N_22955);
nor U27228 (N_27228,N_20815,N_20451);
nor U27229 (N_27229,N_24064,N_23514);
and U27230 (N_27230,N_22313,N_24140);
or U27231 (N_27231,N_23487,N_20283);
nand U27232 (N_27232,N_20369,N_24703);
or U27233 (N_27233,N_23275,N_22796);
and U27234 (N_27234,N_22808,N_21542);
nand U27235 (N_27235,N_22088,N_24259);
nand U27236 (N_27236,N_23981,N_20362);
nand U27237 (N_27237,N_24614,N_20410);
nand U27238 (N_27238,N_24634,N_24823);
nand U27239 (N_27239,N_23831,N_22428);
xnor U27240 (N_27240,N_24721,N_20364);
nor U27241 (N_27241,N_22271,N_23950);
nor U27242 (N_27242,N_24445,N_21806);
xnor U27243 (N_27243,N_21197,N_24971);
xnor U27244 (N_27244,N_20934,N_21491);
nor U27245 (N_27245,N_23021,N_24092);
nand U27246 (N_27246,N_23968,N_23242);
nand U27247 (N_27247,N_21199,N_22201);
xor U27248 (N_27248,N_24463,N_24568);
xnor U27249 (N_27249,N_22287,N_20340);
or U27250 (N_27250,N_23582,N_20707);
xnor U27251 (N_27251,N_22286,N_24548);
nand U27252 (N_27252,N_22903,N_20937);
or U27253 (N_27253,N_20530,N_22825);
or U27254 (N_27254,N_24280,N_22657);
nand U27255 (N_27255,N_21078,N_23835);
or U27256 (N_27256,N_23394,N_21425);
xor U27257 (N_27257,N_21664,N_20250);
or U27258 (N_27258,N_21566,N_20351);
and U27259 (N_27259,N_24611,N_22811);
nand U27260 (N_27260,N_21484,N_24250);
and U27261 (N_27261,N_22975,N_24789);
nor U27262 (N_27262,N_20579,N_22363);
nand U27263 (N_27263,N_21810,N_23435);
nand U27264 (N_27264,N_21556,N_23919);
or U27265 (N_27265,N_20327,N_24559);
xor U27266 (N_27266,N_22301,N_22262);
and U27267 (N_27267,N_23710,N_21322);
nand U27268 (N_27268,N_21222,N_22833);
nor U27269 (N_27269,N_22411,N_22054);
or U27270 (N_27270,N_21630,N_23538);
nor U27271 (N_27271,N_23466,N_20659);
nand U27272 (N_27272,N_24008,N_22656);
nor U27273 (N_27273,N_24900,N_21247);
xnor U27274 (N_27274,N_20978,N_22568);
nor U27275 (N_27275,N_20789,N_22799);
xnor U27276 (N_27276,N_20441,N_21085);
and U27277 (N_27277,N_22559,N_20709);
nand U27278 (N_27278,N_24578,N_20580);
and U27279 (N_27279,N_21634,N_24691);
and U27280 (N_27280,N_23595,N_20422);
or U27281 (N_27281,N_23386,N_20554);
or U27282 (N_27282,N_22881,N_23086);
xnor U27283 (N_27283,N_23718,N_24683);
xnor U27284 (N_27284,N_20705,N_21394);
nand U27285 (N_27285,N_21176,N_21889);
and U27286 (N_27286,N_24325,N_23325);
and U27287 (N_27287,N_21923,N_21698);
xnor U27288 (N_27288,N_24680,N_21787);
nor U27289 (N_27289,N_21108,N_20079);
xnor U27290 (N_27290,N_22142,N_23103);
nand U27291 (N_27291,N_24294,N_24954);
nor U27292 (N_27292,N_23607,N_20979);
and U27293 (N_27293,N_22953,N_22103);
nand U27294 (N_27294,N_20361,N_23880);
xnor U27295 (N_27295,N_21398,N_21622);
xor U27296 (N_27296,N_22143,N_21217);
nand U27297 (N_27297,N_23253,N_22971);
or U27298 (N_27298,N_24599,N_22775);
nor U27299 (N_27299,N_24024,N_21851);
and U27300 (N_27300,N_24564,N_21214);
nor U27301 (N_27301,N_23258,N_22587);
nand U27302 (N_27302,N_20001,N_22585);
and U27303 (N_27303,N_24517,N_22897);
or U27304 (N_27304,N_23147,N_23109);
xnor U27305 (N_27305,N_22480,N_21412);
nand U27306 (N_27306,N_20080,N_21084);
or U27307 (N_27307,N_24169,N_22102);
xnor U27308 (N_27308,N_21029,N_20596);
and U27309 (N_27309,N_21184,N_20424);
xnor U27310 (N_27310,N_24241,N_24246);
or U27311 (N_27311,N_24847,N_21730);
or U27312 (N_27312,N_20154,N_23862);
nand U27313 (N_27313,N_20242,N_20469);
or U27314 (N_27314,N_23724,N_21560);
nor U27315 (N_27315,N_21536,N_23415);
and U27316 (N_27316,N_20505,N_23939);
or U27317 (N_27317,N_21163,N_24950);
nand U27318 (N_27318,N_24765,N_22874);
xor U27319 (N_27319,N_20070,N_20829);
and U27320 (N_27320,N_20834,N_24069);
or U27321 (N_27321,N_23379,N_21658);
xnor U27322 (N_27322,N_24684,N_20055);
and U27323 (N_27323,N_23356,N_21843);
or U27324 (N_27324,N_21559,N_21243);
or U27325 (N_27325,N_21267,N_21673);
and U27326 (N_27326,N_23017,N_24201);
nand U27327 (N_27327,N_22130,N_23652);
and U27328 (N_27328,N_22724,N_22128);
xor U27329 (N_27329,N_22368,N_22087);
or U27330 (N_27330,N_20824,N_21183);
nand U27331 (N_27331,N_23927,N_22387);
nand U27332 (N_27332,N_21353,N_21095);
nor U27333 (N_27333,N_22537,N_20236);
nand U27334 (N_27334,N_21625,N_24485);
nand U27335 (N_27335,N_24743,N_22009);
nor U27336 (N_27336,N_22861,N_21027);
nand U27337 (N_27337,N_20972,N_20078);
nand U27338 (N_27338,N_20731,N_23052);
and U27339 (N_27339,N_20904,N_21360);
nor U27340 (N_27340,N_22780,N_23562);
nor U27341 (N_27341,N_23133,N_23101);
xor U27342 (N_27342,N_24697,N_24308);
xor U27343 (N_27343,N_24709,N_24423);
nor U27344 (N_27344,N_22379,N_24520);
and U27345 (N_27345,N_23891,N_21059);
nor U27346 (N_27346,N_24083,N_23703);
xor U27347 (N_27347,N_21050,N_24134);
or U27348 (N_27348,N_20074,N_21538);
nand U27349 (N_27349,N_24932,N_21071);
xnor U27350 (N_27350,N_22236,N_22640);
nand U27351 (N_27351,N_22274,N_22489);
and U27352 (N_27352,N_21054,N_24183);
nand U27353 (N_27353,N_21632,N_20307);
or U27354 (N_27354,N_23264,N_22160);
nor U27355 (N_27355,N_22943,N_22256);
nand U27356 (N_27356,N_22647,N_22462);
and U27357 (N_27357,N_21433,N_22238);
or U27358 (N_27358,N_24035,N_20241);
or U27359 (N_27359,N_23732,N_23465);
or U27360 (N_27360,N_20884,N_23408);
nand U27361 (N_27361,N_22751,N_22742);
nand U27362 (N_27362,N_23475,N_20967);
and U27363 (N_27363,N_21694,N_20333);
xor U27364 (N_27364,N_23380,N_24213);
xnor U27365 (N_27365,N_20758,N_20605);
nor U27366 (N_27366,N_24821,N_22528);
xnor U27367 (N_27367,N_24082,N_23678);
or U27368 (N_27368,N_22216,N_21458);
xnor U27369 (N_27369,N_20222,N_20665);
nor U27370 (N_27370,N_20570,N_20122);
or U27371 (N_27371,N_23151,N_21193);
nand U27372 (N_27372,N_21878,N_20540);
nand U27373 (N_27373,N_21065,N_20133);
nand U27374 (N_27374,N_21717,N_21564);
and U27375 (N_27375,N_20342,N_24667);
xor U27376 (N_27376,N_21713,N_24500);
xnor U27377 (N_27377,N_21185,N_22471);
nand U27378 (N_27378,N_23262,N_23816);
or U27379 (N_27379,N_23183,N_21948);
xor U27380 (N_27380,N_21122,N_22957);
xnor U27381 (N_27381,N_23729,N_21641);
and U27382 (N_27382,N_23330,N_24846);
and U27383 (N_27383,N_23055,N_21136);
nor U27384 (N_27384,N_24171,N_21426);
xor U27385 (N_27385,N_24539,N_21695);
nor U27386 (N_27386,N_21310,N_20309);
nor U27387 (N_27387,N_20876,N_22620);
and U27388 (N_27388,N_22242,N_22834);
nor U27389 (N_27389,N_21589,N_23894);
nand U27390 (N_27390,N_23804,N_20920);
nand U27391 (N_27391,N_23381,N_22929);
nor U27392 (N_27392,N_24668,N_20495);
or U27393 (N_27393,N_21421,N_22717);
nand U27394 (N_27394,N_22771,N_24362);
xor U27395 (N_27395,N_21598,N_23909);
and U27396 (N_27396,N_23454,N_23817);
nor U27397 (N_27397,N_22893,N_22126);
and U27398 (N_27398,N_20042,N_22586);
nor U27399 (N_27399,N_23342,N_21487);
xnor U27400 (N_27400,N_24779,N_24411);
nand U27401 (N_27401,N_23456,N_23648);
nor U27402 (N_27402,N_24833,N_23299);
nor U27403 (N_27403,N_20134,N_21336);
and U27404 (N_27404,N_24230,N_22035);
or U27405 (N_27405,N_22341,N_21151);
and U27406 (N_27406,N_22965,N_21668);
or U27407 (N_27407,N_21062,N_20284);
xnor U27408 (N_27408,N_24725,N_20167);
and U27409 (N_27409,N_22502,N_22376);
xnor U27410 (N_27410,N_20576,N_22139);
nor U27411 (N_27411,N_23182,N_23669);
and U27412 (N_27412,N_20808,N_22538);
xnor U27413 (N_27413,N_21870,N_21882);
or U27414 (N_27414,N_22738,N_23084);
nand U27415 (N_27415,N_24147,N_23782);
nor U27416 (N_27416,N_23545,N_21958);
nand U27417 (N_27417,N_23995,N_24876);
and U27418 (N_27418,N_20243,N_23324);
xor U27419 (N_27419,N_22292,N_23993);
nor U27420 (N_27420,N_23273,N_20315);
nand U27421 (N_27421,N_23360,N_24408);
nand U27422 (N_27422,N_20234,N_24135);
or U27423 (N_27423,N_20804,N_24014);
nand U27424 (N_27424,N_23556,N_21205);
nor U27425 (N_27425,N_22195,N_20975);
nor U27426 (N_27426,N_22282,N_21283);
nand U27427 (N_27427,N_22575,N_22125);
xor U27428 (N_27428,N_21523,N_20600);
nand U27429 (N_27429,N_21916,N_22547);
nor U27430 (N_27430,N_24283,N_23070);
nand U27431 (N_27431,N_24177,N_24640);
nand U27432 (N_27432,N_24001,N_21142);
nand U27433 (N_27433,N_21045,N_24739);
and U27434 (N_27434,N_24344,N_24352);
nand U27435 (N_27435,N_24165,N_21667);
and U27436 (N_27436,N_23237,N_23457);
and U27437 (N_27437,N_24650,N_24911);
nand U27438 (N_27438,N_22417,N_20251);
and U27439 (N_27439,N_22752,N_23871);
nand U27440 (N_27440,N_21032,N_23644);
and U27441 (N_27441,N_21004,N_22176);
and U27442 (N_27442,N_21708,N_22118);
nand U27443 (N_27443,N_21213,N_21379);
nand U27444 (N_27444,N_24894,N_22949);
nor U27445 (N_27445,N_21738,N_23479);
and U27446 (N_27446,N_22473,N_24326);
or U27447 (N_27447,N_23666,N_24117);
and U27448 (N_27448,N_20175,N_23962);
or U27449 (N_27449,N_23289,N_24332);
xor U27450 (N_27450,N_22703,N_23861);
or U27451 (N_27451,N_21349,N_22875);
and U27452 (N_27452,N_21066,N_20556);
nand U27453 (N_27453,N_24989,N_21533);
nand U27454 (N_27454,N_20313,N_21400);
nor U27455 (N_27455,N_23041,N_21006);
and U27456 (N_27456,N_24509,N_23601);
nand U27457 (N_27457,N_21776,N_24841);
nand U27458 (N_27458,N_20207,N_23585);
nor U27459 (N_27459,N_21334,N_23083);
nor U27460 (N_27460,N_23581,N_23631);
and U27461 (N_27461,N_20958,N_23497);
xnor U27462 (N_27462,N_23058,N_24693);
and U27463 (N_27463,N_20881,N_20548);
nand U27464 (N_27464,N_21028,N_21998);
and U27465 (N_27465,N_20045,N_20426);
xnor U27466 (N_27466,N_24091,N_22999);
or U27467 (N_27467,N_24910,N_24639);
xnor U27468 (N_27468,N_22105,N_20189);
nand U27469 (N_27469,N_22648,N_20828);
and U27470 (N_27470,N_23641,N_21209);
nor U27471 (N_27471,N_24966,N_23489);
xnor U27472 (N_27472,N_20300,N_20111);
nand U27473 (N_27473,N_21712,N_24978);
xnor U27474 (N_27474,N_24970,N_22392);
nor U27475 (N_27475,N_22581,N_23946);
xor U27476 (N_27476,N_20792,N_24695);
nand U27477 (N_27477,N_23954,N_22625);
nor U27478 (N_27478,N_24044,N_23193);
and U27479 (N_27479,N_24757,N_24289);
nand U27480 (N_27480,N_23657,N_23316);
nor U27481 (N_27481,N_21431,N_22718);
or U27482 (N_27482,N_20093,N_22864);
nor U27483 (N_27483,N_21100,N_23679);
or U27484 (N_27484,N_22946,N_24367);
nand U27485 (N_27485,N_20952,N_20489);
and U27486 (N_27486,N_21072,N_23355);
nand U27487 (N_27487,N_20673,N_21492);
nor U27488 (N_27488,N_24474,N_23777);
nor U27489 (N_27489,N_23512,N_22670);
xor U27490 (N_27490,N_21871,N_20660);
xnor U27491 (N_27491,N_21861,N_21743);
xnor U27492 (N_27492,N_23137,N_20873);
or U27493 (N_27493,N_21849,N_22494);
or U27494 (N_27494,N_21037,N_24586);
xnor U27495 (N_27495,N_23971,N_21383);
nand U27496 (N_27496,N_20214,N_24766);
nand U27497 (N_27497,N_23428,N_20429);
xor U27498 (N_27498,N_24660,N_21351);
and U27499 (N_27499,N_22603,N_20592);
nor U27500 (N_27500,N_22002,N_20029);
nand U27501 (N_27501,N_20891,N_21308);
nor U27502 (N_27502,N_21847,N_22169);
nand U27503 (N_27503,N_24186,N_22423);
and U27504 (N_27504,N_23045,N_20614);
nand U27505 (N_27505,N_23269,N_23397);
xnor U27506 (N_27506,N_23981,N_20311);
nand U27507 (N_27507,N_22559,N_24565);
or U27508 (N_27508,N_20324,N_22417);
nor U27509 (N_27509,N_24810,N_20511);
xnor U27510 (N_27510,N_23341,N_22331);
nor U27511 (N_27511,N_24673,N_24449);
or U27512 (N_27512,N_23832,N_20539);
nor U27513 (N_27513,N_23821,N_23854);
and U27514 (N_27514,N_23619,N_24164);
and U27515 (N_27515,N_22321,N_23275);
nor U27516 (N_27516,N_23454,N_23694);
or U27517 (N_27517,N_24325,N_22816);
nand U27518 (N_27518,N_23320,N_21583);
or U27519 (N_27519,N_24238,N_20181);
xor U27520 (N_27520,N_23661,N_24298);
xor U27521 (N_27521,N_20600,N_23270);
and U27522 (N_27522,N_23335,N_21900);
nor U27523 (N_27523,N_23918,N_24829);
nor U27524 (N_27524,N_21713,N_24747);
xnor U27525 (N_27525,N_21665,N_23797);
nor U27526 (N_27526,N_22653,N_23054);
nand U27527 (N_27527,N_21210,N_20907);
xnor U27528 (N_27528,N_21082,N_23724);
xnor U27529 (N_27529,N_23673,N_24678);
xnor U27530 (N_27530,N_20593,N_21781);
nand U27531 (N_27531,N_22293,N_20067);
and U27532 (N_27532,N_21578,N_23586);
or U27533 (N_27533,N_20045,N_22662);
or U27534 (N_27534,N_24635,N_24155);
xor U27535 (N_27535,N_21311,N_20641);
and U27536 (N_27536,N_20373,N_22432);
nor U27537 (N_27537,N_24639,N_22213);
xor U27538 (N_27538,N_22198,N_22579);
nor U27539 (N_27539,N_21929,N_23086);
nor U27540 (N_27540,N_20075,N_20091);
and U27541 (N_27541,N_22806,N_21687);
or U27542 (N_27542,N_23294,N_24520);
xor U27543 (N_27543,N_23990,N_21912);
nand U27544 (N_27544,N_20126,N_21739);
xnor U27545 (N_27545,N_22242,N_24393);
nor U27546 (N_27546,N_22343,N_20474);
and U27547 (N_27547,N_24351,N_23309);
and U27548 (N_27548,N_23614,N_24277);
nand U27549 (N_27549,N_20754,N_21424);
nand U27550 (N_27550,N_20704,N_24150);
or U27551 (N_27551,N_23518,N_22800);
nor U27552 (N_27552,N_23132,N_24228);
and U27553 (N_27553,N_21857,N_22580);
xnor U27554 (N_27554,N_22919,N_20817);
nand U27555 (N_27555,N_21054,N_24621);
and U27556 (N_27556,N_20518,N_24188);
and U27557 (N_27557,N_22103,N_21559);
and U27558 (N_27558,N_21043,N_22545);
and U27559 (N_27559,N_23681,N_24796);
nor U27560 (N_27560,N_21672,N_23123);
nor U27561 (N_27561,N_20399,N_21304);
nand U27562 (N_27562,N_21088,N_21237);
and U27563 (N_27563,N_23139,N_20151);
or U27564 (N_27564,N_23309,N_22910);
and U27565 (N_27565,N_22493,N_21389);
nor U27566 (N_27566,N_23635,N_21477);
or U27567 (N_27567,N_20684,N_20346);
and U27568 (N_27568,N_23927,N_24669);
and U27569 (N_27569,N_22425,N_23072);
xnor U27570 (N_27570,N_24799,N_21643);
nor U27571 (N_27571,N_21721,N_22400);
or U27572 (N_27572,N_21426,N_23684);
and U27573 (N_27573,N_22911,N_21018);
nor U27574 (N_27574,N_20196,N_21283);
or U27575 (N_27575,N_21086,N_20760);
nor U27576 (N_27576,N_23272,N_23892);
nand U27577 (N_27577,N_21476,N_23112);
nor U27578 (N_27578,N_23677,N_20514);
or U27579 (N_27579,N_21145,N_22261);
xor U27580 (N_27580,N_22782,N_23408);
nor U27581 (N_27581,N_20487,N_21771);
xnor U27582 (N_27582,N_24115,N_24869);
and U27583 (N_27583,N_23653,N_24447);
and U27584 (N_27584,N_22054,N_23545);
or U27585 (N_27585,N_23993,N_23918);
or U27586 (N_27586,N_21125,N_21586);
and U27587 (N_27587,N_23859,N_20841);
xor U27588 (N_27588,N_21246,N_21252);
or U27589 (N_27589,N_21561,N_22873);
nor U27590 (N_27590,N_23591,N_20422);
xnor U27591 (N_27591,N_22075,N_24629);
or U27592 (N_27592,N_22033,N_22318);
or U27593 (N_27593,N_20721,N_21105);
or U27594 (N_27594,N_24094,N_22341);
or U27595 (N_27595,N_23817,N_22255);
nor U27596 (N_27596,N_22580,N_23706);
or U27597 (N_27597,N_22814,N_20132);
xor U27598 (N_27598,N_23589,N_24453);
nor U27599 (N_27599,N_20229,N_20493);
and U27600 (N_27600,N_24172,N_24559);
nor U27601 (N_27601,N_22871,N_24399);
nand U27602 (N_27602,N_24594,N_23034);
nor U27603 (N_27603,N_21167,N_20414);
nand U27604 (N_27604,N_24941,N_23267);
nand U27605 (N_27605,N_22708,N_24603);
or U27606 (N_27606,N_23949,N_20775);
nor U27607 (N_27607,N_20830,N_23005);
or U27608 (N_27608,N_23610,N_24941);
nor U27609 (N_27609,N_22995,N_23449);
or U27610 (N_27610,N_23240,N_21731);
xnor U27611 (N_27611,N_23945,N_21213);
or U27612 (N_27612,N_22301,N_24480);
nand U27613 (N_27613,N_21073,N_24462);
nand U27614 (N_27614,N_24477,N_22909);
xor U27615 (N_27615,N_23812,N_23878);
or U27616 (N_27616,N_20636,N_20526);
or U27617 (N_27617,N_20661,N_20093);
nor U27618 (N_27618,N_20999,N_21378);
nor U27619 (N_27619,N_22317,N_22786);
and U27620 (N_27620,N_21378,N_21083);
and U27621 (N_27621,N_22262,N_23696);
xor U27622 (N_27622,N_22573,N_22414);
or U27623 (N_27623,N_20226,N_21217);
or U27624 (N_27624,N_20812,N_24016);
nand U27625 (N_27625,N_21110,N_20552);
or U27626 (N_27626,N_24942,N_20855);
or U27627 (N_27627,N_20013,N_22550);
nand U27628 (N_27628,N_23674,N_21329);
or U27629 (N_27629,N_22832,N_20380);
nand U27630 (N_27630,N_24088,N_21042);
xor U27631 (N_27631,N_20270,N_20625);
or U27632 (N_27632,N_20596,N_23826);
or U27633 (N_27633,N_20995,N_20156);
or U27634 (N_27634,N_23804,N_21566);
xnor U27635 (N_27635,N_21606,N_22179);
or U27636 (N_27636,N_20318,N_24097);
or U27637 (N_27637,N_20989,N_23404);
or U27638 (N_27638,N_24591,N_20290);
nand U27639 (N_27639,N_22474,N_21155);
nand U27640 (N_27640,N_22390,N_24174);
nand U27641 (N_27641,N_20508,N_22328);
or U27642 (N_27642,N_24343,N_21391);
or U27643 (N_27643,N_21812,N_24947);
nand U27644 (N_27644,N_23444,N_24015);
nor U27645 (N_27645,N_24015,N_20446);
nor U27646 (N_27646,N_23078,N_20693);
and U27647 (N_27647,N_21618,N_21628);
and U27648 (N_27648,N_23975,N_22350);
xor U27649 (N_27649,N_21816,N_24183);
nor U27650 (N_27650,N_23836,N_24683);
nor U27651 (N_27651,N_24240,N_23468);
or U27652 (N_27652,N_20217,N_24160);
xor U27653 (N_27653,N_24752,N_20261);
nand U27654 (N_27654,N_20560,N_20412);
nor U27655 (N_27655,N_21539,N_22901);
xnor U27656 (N_27656,N_20171,N_21021);
or U27657 (N_27657,N_21476,N_20335);
nand U27658 (N_27658,N_22108,N_21311);
nand U27659 (N_27659,N_22321,N_20036);
xnor U27660 (N_27660,N_20465,N_24381);
and U27661 (N_27661,N_23172,N_24576);
or U27662 (N_27662,N_24230,N_24827);
nand U27663 (N_27663,N_21910,N_24295);
and U27664 (N_27664,N_20593,N_23104);
or U27665 (N_27665,N_22020,N_22871);
nand U27666 (N_27666,N_23622,N_23395);
nor U27667 (N_27667,N_24078,N_22654);
and U27668 (N_27668,N_21189,N_20773);
nand U27669 (N_27669,N_20136,N_23058);
or U27670 (N_27670,N_20321,N_22853);
and U27671 (N_27671,N_20539,N_20130);
or U27672 (N_27672,N_22389,N_21252);
nand U27673 (N_27673,N_21310,N_20399);
or U27674 (N_27674,N_22160,N_22920);
or U27675 (N_27675,N_21987,N_23423);
nor U27676 (N_27676,N_21221,N_23589);
or U27677 (N_27677,N_21978,N_20075);
xnor U27678 (N_27678,N_21644,N_21763);
xnor U27679 (N_27679,N_22887,N_23361);
and U27680 (N_27680,N_23865,N_21487);
or U27681 (N_27681,N_20812,N_22549);
nand U27682 (N_27682,N_22354,N_23470);
xor U27683 (N_27683,N_24806,N_24319);
xnor U27684 (N_27684,N_23172,N_24818);
nand U27685 (N_27685,N_22568,N_23455);
nand U27686 (N_27686,N_20927,N_21874);
nand U27687 (N_27687,N_24857,N_22121);
or U27688 (N_27688,N_21331,N_20250);
nand U27689 (N_27689,N_23281,N_21314);
or U27690 (N_27690,N_22949,N_23994);
nor U27691 (N_27691,N_22637,N_24564);
and U27692 (N_27692,N_24529,N_22939);
or U27693 (N_27693,N_22392,N_22355);
nand U27694 (N_27694,N_21755,N_21486);
xor U27695 (N_27695,N_22569,N_21794);
nand U27696 (N_27696,N_20601,N_24039);
nor U27697 (N_27697,N_23410,N_20133);
nor U27698 (N_27698,N_21903,N_24213);
nor U27699 (N_27699,N_23660,N_24144);
xor U27700 (N_27700,N_23902,N_22156);
nor U27701 (N_27701,N_23037,N_24238);
xor U27702 (N_27702,N_22979,N_23437);
nor U27703 (N_27703,N_23024,N_21642);
or U27704 (N_27704,N_20925,N_23328);
or U27705 (N_27705,N_22586,N_22487);
or U27706 (N_27706,N_21806,N_22555);
nand U27707 (N_27707,N_20302,N_21995);
nand U27708 (N_27708,N_23050,N_20225);
xnor U27709 (N_27709,N_22493,N_24246);
or U27710 (N_27710,N_22945,N_21598);
nor U27711 (N_27711,N_21159,N_21473);
xor U27712 (N_27712,N_21505,N_22598);
nor U27713 (N_27713,N_20599,N_21167);
and U27714 (N_27714,N_23927,N_23212);
xnor U27715 (N_27715,N_24383,N_20748);
and U27716 (N_27716,N_24661,N_22621);
and U27717 (N_27717,N_21115,N_23810);
nor U27718 (N_27718,N_20673,N_21113);
xnor U27719 (N_27719,N_20395,N_22727);
nand U27720 (N_27720,N_21171,N_21936);
and U27721 (N_27721,N_23431,N_23020);
xnor U27722 (N_27722,N_20713,N_20209);
xor U27723 (N_27723,N_20991,N_24936);
nand U27724 (N_27724,N_22016,N_20176);
nor U27725 (N_27725,N_21844,N_23453);
or U27726 (N_27726,N_21705,N_23659);
and U27727 (N_27727,N_24745,N_22330);
nor U27728 (N_27728,N_21802,N_23607);
xor U27729 (N_27729,N_24892,N_20241);
or U27730 (N_27730,N_20091,N_23000);
and U27731 (N_27731,N_21621,N_23476);
xor U27732 (N_27732,N_23386,N_22555);
or U27733 (N_27733,N_23702,N_22430);
and U27734 (N_27734,N_23476,N_21361);
nor U27735 (N_27735,N_24002,N_21727);
or U27736 (N_27736,N_24787,N_21906);
xor U27737 (N_27737,N_20089,N_22921);
or U27738 (N_27738,N_24173,N_22518);
nor U27739 (N_27739,N_21478,N_23305);
and U27740 (N_27740,N_20330,N_24311);
xnor U27741 (N_27741,N_21368,N_20565);
and U27742 (N_27742,N_23445,N_23953);
nor U27743 (N_27743,N_21677,N_24814);
xnor U27744 (N_27744,N_20857,N_21216);
nand U27745 (N_27745,N_20303,N_23602);
nor U27746 (N_27746,N_20995,N_21570);
or U27747 (N_27747,N_23392,N_20120);
xor U27748 (N_27748,N_23301,N_21033);
nor U27749 (N_27749,N_22151,N_23519);
nor U27750 (N_27750,N_20914,N_23141);
or U27751 (N_27751,N_21699,N_22602);
nand U27752 (N_27752,N_20724,N_20923);
and U27753 (N_27753,N_22666,N_23370);
nand U27754 (N_27754,N_21921,N_21964);
nor U27755 (N_27755,N_20377,N_20354);
xor U27756 (N_27756,N_23938,N_21641);
nor U27757 (N_27757,N_21133,N_20617);
and U27758 (N_27758,N_23093,N_21837);
or U27759 (N_27759,N_23344,N_21557);
and U27760 (N_27760,N_21977,N_20270);
and U27761 (N_27761,N_20773,N_22672);
and U27762 (N_27762,N_21875,N_23982);
nand U27763 (N_27763,N_24810,N_22975);
nor U27764 (N_27764,N_20835,N_20488);
nand U27765 (N_27765,N_22047,N_22583);
xnor U27766 (N_27766,N_21710,N_20766);
or U27767 (N_27767,N_23470,N_22881);
nand U27768 (N_27768,N_21921,N_21903);
nor U27769 (N_27769,N_24894,N_23754);
nor U27770 (N_27770,N_21143,N_22340);
nand U27771 (N_27771,N_20438,N_22180);
nor U27772 (N_27772,N_23398,N_21073);
and U27773 (N_27773,N_20222,N_20661);
nor U27774 (N_27774,N_23591,N_24086);
nand U27775 (N_27775,N_22727,N_24011);
xor U27776 (N_27776,N_21178,N_23339);
and U27777 (N_27777,N_21402,N_22287);
or U27778 (N_27778,N_20763,N_24754);
and U27779 (N_27779,N_22895,N_23052);
nor U27780 (N_27780,N_21082,N_20056);
nor U27781 (N_27781,N_20017,N_23741);
nand U27782 (N_27782,N_21877,N_24621);
nand U27783 (N_27783,N_21252,N_23363);
xor U27784 (N_27784,N_22872,N_20424);
xor U27785 (N_27785,N_21303,N_20017);
nor U27786 (N_27786,N_24685,N_21634);
nor U27787 (N_27787,N_21924,N_20745);
nor U27788 (N_27788,N_23417,N_20306);
nor U27789 (N_27789,N_20268,N_21339);
nor U27790 (N_27790,N_23262,N_20283);
xor U27791 (N_27791,N_24550,N_20851);
nand U27792 (N_27792,N_24529,N_22884);
or U27793 (N_27793,N_20051,N_24087);
and U27794 (N_27794,N_20960,N_21805);
xnor U27795 (N_27795,N_23542,N_24102);
and U27796 (N_27796,N_24783,N_22600);
or U27797 (N_27797,N_20124,N_23529);
or U27798 (N_27798,N_21914,N_23971);
nor U27799 (N_27799,N_24464,N_23340);
or U27800 (N_27800,N_23299,N_24087);
or U27801 (N_27801,N_24081,N_20560);
or U27802 (N_27802,N_20950,N_21982);
or U27803 (N_27803,N_21595,N_22444);
or U27804 (N_27804,N_24688,N_24353);
and U27805 (N_27805,N_21140,N_21295);
nand U27806 (N_27806,N_20129,N_21745);
nand U27807 (N_27807,N_20760,N_23059);
and U27808 (N_27808,N_24301,N_22781);
xnor U27809 (N_27809,N_24132,N_20436);
and U27810 (N_27810,N_22642,N_24482);
nor U27811 (N_27811,N_22136,N_20179);
xnor U27812 (N_27812,N_20745,N_24037);
and U27813 (N_27813,N_23944,N_22228);
xor U27814 (N_27814,N_24971,N_20047);
xor U27815 (N_27815,N_24148,N_23039);
xnor U27816 (N_27816,N_23722,N_20591);
nor U27817 (N_27817,N_20358,N_22176);
nor U27818 (N_27818,N_21981,N_20988);
xor U27819 (N_27819,N_21631,N_22128);
nand U27820 (N_27820,N_21621,N_21617);
xnor U27821 (N_27821,N_22045,N_21229);
or U27822 (N_27822,N_21355,N_23383);
xnor U27823 (N_27823,N_21758,N_23109);
and U27824 (N_27824,N_23286,N_24416);
nor U27825 (N_27825,N_23584,N_20890);
or U27826 (N_27826,N_20437,N_22587);
xnor U27827 (N_27827,N_20439,N_22898);
and U27828 (N_27828,N_21572,N_24567);
and U27829 (N_27829,N_22282,N_20039);
nor U27830 (N_27830,N_20490,N_23336);
nand U27831 (N_27831,N_23612,N_21499);
nor U27832 (N_27832,N_20548,N_20106);
xnor U27833 (N_27833,N_23377,N_23220);
nand U27834 (N_27834,N_21815,N_22464);
nand U27835 (N_27835,N_23568,N_21589);
and U27836 (N_27836,N_20502,N_21013);
and U27837 (N_27837,N_22018,N_24374);
nor U27838 (N_27838,N_21826,N_23840);
and U27839 (N_27839,N_20993,N_22862);
nand U27840 (N_27840,N_22660,N_23839);
nand U27841 (N_27841,N_21503,N_20908);
and U27842 (N_27842,N_21084,N_22374);
nand U27843 (N_27843,N_23549,N_23562);
nand U27844 (N_27844,N_22122,N_21417);
nand U27845 (N_27845,N_22156,N_24691);
or U27846 (N_27846,N_24193,N_23268);
or U27847 (N_27847,N_21114,N_23254);
nor U27848 (N_27848,N_20049,N_23148);
xnor U27849 (N_27849,N_21753,N_20839);
nor U27850 (N_27850,N_22083,N_20182);
xor U27851 (N_27851,N_22907,N_20553);
nor U27852 (N_27852,N_22103,N_22870);
nand U27853 (N_27853,N_21586,N_21954);
nand U27854 (N_27854,N_23108,N_21680);
or U27855 (N_27855,N_23368,N_21986);
xnor U27856 (N_27856,N_21172,N_21892);
or U27857 (N_27857,N_22141,N_20074);
or U27858 (N_27858,N_22865,N_23275);
xnor U27859 (N_27859,N_21229,N_22138);
and U27860 (N_27860,N_23324,N_20802);
and U27861 (N_27861,N_21854,N_20829);
nor U27862 (N_27862,N_22675,N_23422);
nor U27863 (N_27863,N_20690,N_21712);
nor U27864 (N_27864,N_23441,N_22335);
xnor U27865 (N_27865,N_23602,N_23925);
nand U27866 (N_27866,N_24222,N_21974);
and U27867 (N_27867,N_22139,N_22411);
or U27868 (N_27868,N_24017,N_24672);
nor U27869 (N_27869,N_22701,N_20708);
xor U27870 (N_27870,N_23409,N_24741);
xor U27871 (N_27871,N_21030,N_24055);
nor U27872 (N_27872,N_23650,N_20021);
and U27873 (N_27873,N_23680,N_24382);
nand U27874 (N_27874,N_22807,N_20053);
or U27875 (N_27875,N_23035,N_24714);
or U27876 (N_27876,N_22941,N_24077);
nand U27877 (N_27877,N_23509,N_23241);
xnor U27878 (N_27878,N_21420,N_20863);
and U27879 (N_27879,N_21165,N_22187);
or U27880 (N_27880,N_22407,N_21817);
or U27881 (N_27881,N_23907,N_20626);
or U27882 (N_27882,N_20759,N_21570);
xor U27883 (N_27883,N_21232,N_24879);
xor U27884 (N_27884,N_21414,N_23384);
or U27885 (N_27885,N_22223,N_24555);
and U27886 (N_27886,N_21301,N_23727);
and U27887 (N_27887,N_21910,N_23716);
nand U27888 (N_27888,N_22436,N_21601);
nor U27889 (N_27889,N_24541,N_22531);
xor U27890 (N_27890,N_21719,N_21557);
and U27891 (N_27891,N_21505,N_23301);
xor U27892 (N_27892,N_23885,N_22448);
nor U27893 (N_27893,N_23969,N_21709);
nand U27894 (N_27894,N_24828,N_23544);
and U27895 (N_27895,N_22794,N_22671);
and U27896 (N_27896,N_20614,N_23699);
nand U27897 (N_27897,N_22499,N_20446);
xor U27898 (N_27898,N_23908,N_24276);
and U27899 (N_27899,N_22433,N_22633);
xnor U27900 (N_27900,N_24522,N_23122);
xnor U27901 (N_27901,N_23942,N_21686);
nor U27902 (N_27902,N_21679,N_23567);
nor U27903 (N_27903,N_22353,N_21856);
nand U27904 (N_27904,N_24648,N_24497);
and U27905 (N_27905,N_21920,N_21392);
nor U27906 (N_27906,N_23937,N_21013);
xnor U27907 (N_27907,N_24948,N_20197);
and U27908 (N_27908,N_20743,N_24367);
or U27909 (N_27909,N_21270,N_23705);
nand U27910 (N_27910,N_24199,N_23541);
xnor U27911 (N_27911,N_22956,N_20541);
nand U27912 (N_27912,N_20210,N_21641);
xor U27913 (N_27913,N_22104,N_23847);
nor U27914 (N_27914,N_22484,N_21500);
xnor U27915 (N_27915,N_23721,N_23279);
or U27916 (N_27916,N_23321,N_20367);
nand U27917 (N_27917,N_24410,N_20168);
nand U27918 (N_27918,N_23771,N_23302);
nand U27919 (N_27919,N_22219,N_23779);
nor U27920 (N_27920,N_21090,N_20734);
and U27921 (N_27921,N_24004,N_23848);
and U27922 (N_27922,N_20075,N_20084);
and U27923 (N_27923,N_23697,N_22026);
and U27924 (N_27924,N_21041,N_20248);
and U27925 (N_27925,N_24877,N_22723);
xor U27926 (N_27926,N_21501,N_23291);
and U27927 (N_27927,N_22369,N_24544);
and U27928 (N_27928,N_21153,N_21185);
nand U27929 (N_27929,N_24934,N_20131);
and U27930 (N_27930,N_23155,N_24624);
nand U27931 (N_27931,N_23749,N_22116);
or U27932 (N_27932,N_20967,N_23919);
xor U27933 (N_27933,N_21909,N_20982);
or U27934 (N_27934,N_22436,N_22204);
and U27935 (N_27935,N_24640,N_23047);
nand U27936 (N_27936,N_24712,N_20971);
xnor U27937 (N_27937,N_20833,N_20910);
nand U27938 (N_27938,N_24336,N_22948);
xor U27939 (N_27939,N_23764,N_23870);
nand U27940 (N_27940,N_23604,N_20515);
nor U27941 (N_27941,N_24604,N_21523);
nor U27942 (N_27942,N_20557,N_21032);
nor U27943 (N_27943,N_22073,N_24269);
or U27944 (N_27944,N_22670,N_20981);
or U27945 (N_27945,N_24168,N_21762);
or U27946 (N_27946,N_23077,N_22843);
xnor U27947 (N_27947,N_23213,N_22511);
xor U27948 (N_27948,N_20636,N_22377);
nor U27949 (N_27949,N_20234,N_23897);
and U27950 (N_27950,N_22804,N_20354);
nand U27951 (N_27951,N_20449,N_22688);
nor U27952 (N_27952,N_21352,N_23463);
nor U27953 (N_27953,N_21684,N_21995);
or U27954 (N_27954,N_23531,N_21060);
xnor U27955 (N_27955,N_20118,N_22818);
and U27956 (N_27956,N_20842,N_22901);
nor U27957 (N_27957,N_20932,N_22621);
nand U27958 (N_27958,N_20802,N_23940);
or U27959 (N_27959,N_24360,N_24110);
or U27960 (N_27960,N_21884,N_20245);
xnor U27961 (N_27961,N_20975,N_24332);
nand U27962 (N_27962,N_21868,N_23503);
nand U27963 (N_27963,N_22500,N_21739);
and U27964 (N_27964,N_23959,N_21216);
or U27965 (N_27965,N_20983,N_24743);
nand U27966 (N_27966,N_20159,N_20928);
nand U27967 (N_27967,N_20206,N_22109);
nor U27968 (N_27968,N_20125,N_24530);
and U27969 (N_27969,N_23393,N_20794);
or U27970 (N_27970,N_23458,N_20121);
and U27971 (N_27971,N_22507,N_23757);
or U27972 (N_27972,N_23132,N_22236);
nand U27973 (N_27973,N_23777,N_23698);
or U27974 (N_27974,N_20047,N_20007);
nand U27975 (N_27975,N_20597,N_21191);
or U27976 (N_27976,N_24757,N_22363);
xnor U27977 (N_27977,N_21525,N_23143);
xor U27978 (N_27978,N_22356,N_24273);
xor U27979 (N_27979,N_23540,N_20671);
xnor U27980 (N_27980,N_21098,N_23042);
and U27981 (N_27981,N_22928,N_21392);
or U27982 (N_27982,N_21665,N_20227);
and U27983 (N_27983,N_20757,N_21833);
and U27984 (N_27984,N_22694,N_23849);
and U27985 (N_27985,N_20830,N_24141);
and U27986 (N_27986,N_24431,N_24688);
or U27987 (N_27987,N_21101,N_23950);
nand U27988 (N_27988,N_20825,N_20564);
or U27989 (N_27989,N_20148,N_24204);
xnor U27990 (N_27990,N_20638,N_23298);
or U27991 (N_27991,N_22338,N_24317);
nor U27992 (N_27992,N_21304,N_23894);
xor U27993 (N_27993,N_22335,N_21955);
and U27994 (N_27994,N_20227,N_20441);
and U27995 (N_27995,N_24615,N_23540);
nor U27996 (N_27996,N_20046,N_21101);
or U27997 (N_27997,N_24163,N_23272);
or U27998 (N_27998,N_21749,N_23466);
nand U27999 (N_27999,N_20593,N_24832);
xnor U28000 (N_28000,N_22578,N_24470);
nand U28001 (N_28001,N_23393,N_24071);
and U28002 (N_28002,N_24910,N_23658);
nand U28003 (N_28003,N_22361,N_23860);
xnor U28004 (N_28004,N_22656,N_21699);
and U28005 (N_28005,N_20486,N_21465);
nand U28006 (N_28006,N_22964,N_21854);
xor U28007 (N_28007,N_22283,N_21990);
nor U28008 (N_28008,N_22936,N_21212);
xor U28009 (N_28009,N_22221,N_20190);
or U28010 (N_28010,N_22890,N_23063);
nand U28011 (N_28011,N_23808,N_23213);
xnor U28012 (N_28012,N_22450,N_22809);
nor U28013 (N_28013,N_22644,N_22382);
nor U28014 (N_28014,N_22647,N_21051);
and U28015 (N_28015,N_24982,N_20424);
or U28016 (N_28016,N_21362,N_22770);
or U28017 (N_28017,N_24599,N_24734);
nand U28018 (N_28018,N_23905,N_24147);
and U28019 (N_28019,N_23915,N_20031);
or U28020 (N_28020,N_22784,N_22715);
xor U28021 (N_28021,N_23654,N_20418);
nor U28022 (N_28022,N_20387,N_20187);
or U28023 (N_28023,N_22012,N_21476);
xor U28024 (N_28024,N_20754,N_24088);
or U28025 (N_28025,N_24168,N_23472);
nor U28026 (N_28026,N_24430,N_20182);
nand U28027 (N_28027,N_22969,N_21923);
nor U28028 (N_28028,N_24721,N_23257);
nor U28029 (N_28029,N_22671,N_20662);
nor U28030 (N_28030,N_23875,N_23689);
and U28031 (N_28031,N_20347,N_24310);
xnor U28032 (N_28032,N_22775,N_23573);
xor U28033 (N_28033,N_20626,N_20413);
nand U28034 (N_28034,N_24267,N_20389);
nand U28035 (N_28035,N_21747,N_22037);
or U28036 (N_28036,N_20833,N_24140);
nor U28037 (N_28037,N_23875,N_21808);
xor U28038 (N_28038,N_20756,N_20212);
nand U28039 (N_28039,N_22440,N_24162);
xor U28040 (N_28040,N_21276,N_24113);
nor U28041 (N_28041,N_23791,N_21805);
and U28042 (N_28042,N_21365,N_20652);
nor U28043 (N_28043,N_20164,N_22438);
nand U28044 (N_28044,N_22007,N_20903);
or U28045 (N_28045,N_20256,N_24589);
or U28046 (N_28046,N_20122,N_21682);
and U28047 (N_28047,N_24318,N_23726);
xnor U28048 (N_28048,N_23654,N_23124);
and U28049 (N_28049,N_23807,N_24674);
nor U28050 (N_28050,N_24939,N_24024);
and U28051 (N_28051,N_23816,N_20768);
and U28052 (N_28052,N_21540,N_20985);
and U28053 (N_28053,N_24156,N_22949);
nor U28054 (N_28054,N_22962,N_21926);
nand U28055 (N_28055,N_23242,N_20040);
xor U28056 (N_28056,N_22315,N_22566);
and U28057 (N_28057,N_24985,N_20195);
xor U28058 (N_28058,N_24378,N_20251);
nor U28059 (N_28059,N_21576,N_23464);
nor U28060 (N_28060,N_23087,N_21937);
or U28061 (N_28061,N_22901,N_24336);
or U28062 (N_28062,N_22423,N_20433);
nor U28063 (N_28063,N_24427,N_21374);
or U28064 (N_28064,N_22459,N_23883);
nor U28065 (N_28065,N_20871,N_22402);
or U28066 (N_28066,N_24474,N_24695);
nor U28067 (N_28067,N_24293,N_20065);
xor U28068 (N_28068,N_23117,N_23594);
nor U28069 (N_28069,N_24652,N_24428);
xor U28070 (N_28070,N_24018,N_23215);
nor U28071 (N_28071,N_22121,N_23239);
nand U28072 (N_28072,N_22235,N_23480);
xor U28073 (N_28073,N_24759,N_22022);
and U28074 (N_28074,N_20130,N_20466);
nand U28075 (N_28075,N_20427,N_24286);
xnor U28076 (N_28076,N_24240,N_22674);
nand U28077 (N_28077,N_24549,N_24235);
nor U28078 (N_28078,N_24610,N_23028);
nor U28079 (N_28079,N_23070,N_21091);
nor U28080 (N_28080,N_24477,N_24991);
and U28081 (N_28081,N_22223,N_22413);
and U28082 (N_28082,N_23366,N_21263);
nand U28083 (N_28083,N_23827,N_20839);
nand U28084 (N_28084,N_24374,N_20291);
or U28085 (N_28085,N_23199,N_22675);
and U28086 (N_28086,N_24715,N_22470);
xor U28087 (N_28087,N_23491,N_23286);
or U28088 (N_28088,N_23694,N_22244);
xor U28089 (N_28089,N_20637,N_24448);
or U28090 (N_28090,N_23507,N_22466);
or U28091 (N_28091,N_24287,N_22886);
nor U28092 (N_28092,N_24592,N_22482);
xor U28093 (N_28093,N_23991,N_20996);
nand U28094 (N_28094,N_22783,N_20425);
nand U28095 (N_28095,N_21918,N_21754);
nand U28096 (N_28096,N_21027,N_23221);
nor U28097 (N_28097,N_22241,N_22183);
or U28098 (N_28098,N_23626,N_21742);
and U28099 (N_28099,N_24714,N_22318);
nor U28100 (N_28100,N_23102,N_24062);
nand U28101 (N_28101,N_24078,N_22590);
nor U28102 (N_28102,N_23144,N_24746);
xor U28103 (N_28103,N_22553,N_21956);
and U28104 (N_28104,N_24815,N_22619);
nand U28105 (N_28105,N_20488,N_21396);
nor U28106 (N_28106,N_23812,N_23880);
nor U28107 (N_28107,N_22811,N_24030);
nand U28108 (N_28108,N_23709,N_23119);
nand U28109 (N_28109,N_20539,N_23947);
nand U28110 (N_28110,N_24079,N_20446);
or U28111 (N_28111,N_21137,N_21485);
nand U28112 (N_28112,N_21293,N_21315);
nand U28113 (N_28113,N_20321,N_21096);
nand U28114 (N_28114,N_23190,N_21671);
nand U28115 (N_28115,N_21837,N_20737);
nand U28116 (N_28116,N_22886,N_24148);
nor U28117 (N_28117,N_23181,N_21483);
nand U28118 (N_28118,N_24660,N_20892);
xnor U28119 (N_28119,N_20648,N_20093);
and U28120 (N_28120,N_22147,N_23302);
xnor U28121 (N_28121,N_22954,N_21930);
nand U28122 (N_28122,N_20308,N_20421);
nand U28123 (N_28123,N_22738,N_20836);
or U28124 (N_28124,N_20157,N_22879);
nand U28125 (N_28125,N_20261,N_21773);
and U28126 (N_28126,N_24414,N_22731);
nor U28127 (N_28127,N_21737,N_24819);
or U28128 (N_28128,N_22085,N_20337);
nand U28129 (N_28129,N_24301,N_21289);
nand U28130 (N_28130,N_22933,N_21945);
or U28131 (N_28131,N_24595,N_20571);
and U28132 (N_28132,N_22679,N_23158);
or U28133 (N_28133,N_20790,N_20049);
xor U28134 (N_28134,N_24776,N_23415);
nand U28135 (N_28135,N_24065,N_23309);
or U28136 (N_28136,N_23842,N_23052);
nand U28137 (N_28137,N_21598,N_24431);
nor U28138 (N_28138,N_24344,N_23854);
xor U28139 (N_28139,N_22617,N_21954);
nand U28140 (N_28140,N_23044,N_24065);
nor U28141 (N_28141,N_24561,N_20873);
nand U28142 (N_28142,N_22723,N_22899);
nor U28143 (N_28143,N_21997,N_23575);
or U28144 (N_28144,N_22216,N_23526);
nand U28145 (N_28145,N_22509,N_20405);
and U28146 (N_28146,N_20499,N_23537);
nor U28147 (N_28147,N_21917,N_23012);
or U28148 (N_28148,N_21130,N_20646);
or U28149 (N_28149,N_24082,N_21078);
and U28150 (N_28150,N_24204,N_23788);
nor U28151 (N_28151,N_22500,N_22641);
nand U28152 (N_28152,N_21484,N_22420);
nor U28153 (N_28153,N_20720,N_23895);
xor U28154 (N_28154,N_24633,N_23380);
or U28155 (N_28155,N_21294,N_21910);
nor U28156 (N_28156,N_24554,N_24242);
nor U28157 (N_28157,N_20988,N_23238);
or U28158 (N_28158,N_23777,N_20847);
xor U28159 (N_28159,N_21213,N_24887);
or U28160 (N_28160,N_20939,N_22030);
and U28161 (N_28161,N_24025,N_24091);
nand U28162 (N_28162,N_20122,N_20981);
nor U28163 (N_28163,N_21439,N_24929);
or U28164 (N_28164,N_23531,N_21595);
xnor U28165 (N_28165,N_21183,N_24546);
and U28166 (N_28166,N_22570,N_20392);
and U28167 (N_28167,N_21272,N_23508);
nor U28168 (N_28168,N_20232,N_22070);
nand U28169 (N_28169,N_21223,N_20172);
nor U28170 (N_28170,N_22277,N_20019);
xor U28171 (N_28171,N_23840,N_21671);
nor U28172 (N_28172,N_20650,N_23151);
nor U28173 (N_28173,N_23126,N_23092);
or U28174 (N_28174,N_23535,N_24663);
nor U28175 (N_28175,N_20887,N_23733);
nor U28176 (N_28176,N_22917,N_24276);
xor U28177 (N_28177,N_21055,N_22673);
nor U28178 (N_28178,N_20478,N_20111);
xor U28179 (N_28179,N_23513,N_23495);
nor U28180 (N_28180,N_21025,N_23639);
nand U28181 (N_28181,N_24645,N_23918);
nand U28182 (N_28182,N_22927,N_22082);
nand U28183 (N_28183,N_21198,N_23996);
xor U28184 (N_28184,N_23744,N_22537);
xor U28185 (N_28185,N_21810,N_24004);
xor U28186 (N_28186,N_24036,N_22473);
or U28187 (N_28187,N_23123,N_20783);
nand U28188 (N_28188,N_22535,N_22294);
nor U28189 (N_28189,N_22929,N_21063);
or U28190 (N_28190,N_22118,N_24862);
nand U28191 (N_28191,N_21765,N_22197);
xnor U28192 (N_28192,N_24152,N_23083);
or U28193 (N_28193,N_24086,N_20923);
nor U28194 (N_28194,N_20392,N_22165);
nor U28195 (N_28195,N_21117,N_21112);
xnor U28196 (N_28196,N_21473,N_23755);
or U28197 (N_28197,N_22537,N_20733);
xnor U28198 (N_28198,N_22565,N_24645);
nand U28199 (N_28199,N_20914,N_24317);
and U28200 (N_28200,N_23589,N_23448);
nand U28201 (N_28201,N_24161,N_22036);
nand U28202 (N_28202,N_20829,N_21910);
nand U28203 (N_28203,N_23071,N_24578);
or U28204 (N_28204,N_21102,N_20092);
nand U28205 (N_28205,N_24259,N_20258);
xnor U28206 (N_28206,N_24911,N_23249);
and U28207 (N_28207,N_21380,N_21165);
nor U28208 (N_28208,N_22134,N_23021);
and U28209 (N_28209,N_20314,N_21337);
or U28210 (N_28210,N_22782,N_23870);
nand U28211 (N_28211,N_24195,N_22357);
nand U28212 (N_28212,N_24943,N_20510);
nand U28213 (N_28213,N_24959,N_21563);
xnor U28214 (N_28214,N_21986,N_24106);
nor U28215 (N_28215,N_21854,N_22089);
nand U28216 (N_28216,N_20422,N_21621);
nand U28217 (N_28217,N_21491,N_22344);
nor U28218 (N_28218,N_22719,N_22908);
xnor U28219 (N_28219,N_22378,N_24998);
nand U28220 (N_28220,N_24543,N_22382);
nand U28221 (N_28221,N_24260,N_23594);
xnor U28222 (N_28222,N_24432,N_23061);
xnor U28223 (N_28223,N_24707,N_20215);
xnor U28224 (N_28224,N_21884,N_20042);
nand U28225 (N_28225,N_20654,N_20622);
nor U28226 (N_28226,N_21145,N_20745);
nand U28227 (N_28227,N_21939,N_20931);
nor U28228 (N_28228,N_24571,N_21364);
nor U28229 (N_28229,N_22686,N_23862);
nand U28230 (N_28230,N_23588,N_20791);
and U28231 (N_28231,N_22189,N_20033);
xor U28232 (N_28232,N_21986,N_24846);
nand U28233 (N_28233,N_21855,N_20433);
or U28234 (N_28234,N_21137,N_23079);
xnor U28235 (N_28235,N_22925,N_21597);
nor U28236 (N_28236,N_24318,N_24687);
xnor U28237 (N_28237,N_20516,N_24705);
nand U28238 (N_28238,N_23697,N_24172);
nor U28239 (N_28239,N_24424,N_21130);
or U28240 (N_28240,N_21540,N_21096);
nand U28241 (N_28241,N_21927,N_20908);
and U28242 (N_28242,N_24383,N_22143);
nand U28243 (N_28243,N_21736,N_20822);
and U28244 (N_28244,N_22122,N_20853);
nor U28245 (N_28245,N_20868,N_21466);
and U28246 (N_28246,N_21104,N_20087);
and U28247 (N_28247,N_21097,N_20584);
nor U28248 (N_28248,N_22917,N_20072);
and U28249 (N_28249,N_23268,N_24968);
xnor U28250 (N_28250,N_21374,N_22473);
xor U28251 (N_28251,N_22561,N_20800);
xnor U28252 (N_28252,N_24479,N_22631);
nor U28253 (N_28253,N_23728,N_23630);
xor U28254 (N_28254,N_23442,N_24250);
xnor U28255 (N_28255,N_21032,N_20572);
or U28256 (N_28256,N_21893,N_24182);
xnor U28257 (N_28257,N_24950,N_21836);
xor U28258 (N_28258,N_21138,N_20356);
xnor U28259 (N_28259,N_20987,N_22727);
nor U28260 (N_28260,N_23855,N_22254);
xor U28261 (N_28261,N_20807,N_21044);
or U28262 (N_28262,N_21283,N_22418);
xnor U28263 (N_28263,N_21160,N_23538);
xor U28264 (N_28264,N_21360,N_22443);
and U28265 (N_28265,N_22496,N_21268);
or U28266 (N_28266,N_22973,N_23184);
nand U28267 (N_28267,N_22717,N_23630);
and U28268 (N_28268,N_22516,N_20026);
xor U28269 (N_28269,N_20992,N_21881);
xnor U28270 (N_28270,N_22009,N_23802);
and U28271 (N_28271,N_22512,N_21915);
or U28272 (N_28272,N_21378,N_24268);
and U28273 (N_28273,N_24970,N_24988);
nor U28274 (N_28274,N_22420,N_24637);
and U28275 (N_28275,N_22089,N_24049);
nor U28276 (N_28276,N_20277,N_23984);
nor U28277 (N_28277,N_21564,N_22060);
nand U28278 (N_28278,N_23863,N_23274);
xor U28279 (N_28279,N_22095,N_20958);
nand U28280 (N_28280,N_22278,N_21061);
or U28281 (N_28281,N_22122,N_23424);
or U28282 (N_28282,N_20748,N_21683);
nor U28283 (N_28283,N_24742,N_23149);
xor U28284 (N_28284,N_24711,N_20819);
or U28285 (N_28285,N_23803,N_20837);
xnor U28286 (N_28286,N_23265,N_24642);
nand U28287 (N_28287,N_20770,N_22523);
xor U28288 (N_28288,N_24330,N_21710);
xnor U28289 (N_28289,N_21806,N_21053);
or U28290 (N_28290,N_24220,N_24852);
nor U28291 (N_28291,N_24337,N_23349);
xor U28292 (N_28292,N_22178,N_23978);
nor U28293 (N_28293,N_21015,N_21422);
xnor U28294 (N_28294,N_22350,N_22940);
and U28295 (N_28295,N_21527,N_24259);
and U28296 (N_28296,N_23246,N_20104);
and U28297 (N_28297,N_21484,N_22124);
nor U28298 (N_28298,N_21627,N_20227);
xor U28299 (N_28299,N_23918,N_22365);
xnor U28300 (N_28300,N_22525,N_21027);
nor U28301 (N_28301,N_22455,N_20661);
nand U28302 (N_28302,N_20527,N_24950);
nor U28303 (N_28303,N_24386,N_22690);
or U28304 (N_28304,N_22433,N_22854);
and U28305 (N_28305,N_24044,N_21002);
nor U28306 (N_28306,N_22857,N_20234);
or U28307 (N_28307,N_24420,N_22814);
xor U28308 (N_28308,N_23468,N_23746);
or U28309 (N_28309,N_21837,N_20002);
xnor U28310 (N_28310,N_22146,N_22007);
or U28311 (N_28311,N_22823,N_20510);
and U28312 (N_28312,N_24200,N_20551);
nand U28313 (N_28313,N_23110,N_21969);
xnor U28314 (N_28314,N_22003,N_24183);
xnor U28315 (N_28315,N_24350,N_21869);
nor U28316 (N_28316,N_21343,N_24520);
nand U28317 (N_28317,N_24508,N_21360);
and U28318 (N_28318,N_24963,N_22242);
nand U28319 (N_28319,N_23753,N_21200);
nand U28320 (N_28320,N_24176,N_23699);
nand U28321 (N_28321,N_21690,N_22078);
nand U28322 (N_28322,N_24090,N_20211);
xnor U28323 (N_28323,N_21183,N_23994);
or U28324 (N_28324,N_23879,N_22481);
and U28325 (N_28325,N_20119,N_20866);
and U28326 (N_28326,N_24520,N_21335);
nor U28327 (N_28327,N_20420,N_22177);
nor U28328 (N_28328,N_20846,N_24716);
or U28329 (N_28329,N_24798,N_22277);
nor U28330 (N_28330,N_24524,N_24352);
xor U28331 (N_28331,N_24893,N_22881);
nor U28332 (N_28332,N_24011,N_21466);
nor U28333 (N_28333,N_24452,N_24155);
xnor U28334 (N_28334,N_23877,N_20032);
and U28335 (N_28335,N_22769,N_21954);
xor U28336 (N_28336,N_21758,N_21045);
xnor U28337 (N_28337,N_21857,N_20352);
nand U28338 (N_28338,N_24184,N_20299);
nand U28339 (N_28339,N_21118,N_23727);
xnor U28340 (N_28340,N_24530,N_23494);
nor U28341 (N_28341,N_22968,N_23893);
and U28342 (N_28342,N_21404,N_22095);
nand U28343 (N_28343,N_23193,N_24656);
or U28344 (N_28344,N_22145,N_21517);
nand U28345 (N_28345,N_24907,N_20914);
nand U28346 (N_28346,N_20568,N_20480);
and U28347 (N_28347,N_20552,N_20958);
or U28348 (N_28348,N_21016,N_21779);
and U28349 (N_28349,N_20922,N_22781);
or U28350 (N_28350,N_23803,N_24016);
and U28351 (N_28351,N_24054,N_23865);
nand U28352 (N_28352,N_20022,N_21505);
nor U28353 (N_28353,N_21297,N_22659);
or U28354 (N_28354,N_21527,N_20674);
nand U28355 (N_28355,N_24696,N_24340);
or U28356 (N_28356,N_20991,N_20397);
and U28357 (N_28357,N_23515,N_21889);
nor U28358 (N_28358,N_22246,N_23726);
and U28359 (N_28359,N_20157,N_21928);
nor U28360 (N_28360,N_22427,N_22723);
and U28361 (N_28361,N_22770,N_23739);
xor U28362 (N_28362,N_22976,N_24439);
nor U28363 (N_28363,N_22752,N_22984);
xnor U28364 (N_28364,N_21282,N_23872);
nor U28365 (N_28365,N_23850,N_23822);
xor U28366 (N_28366,N_21621,N_21916);
nand U28367 (N_28367,N_20520,N_21437);
nor U28368 (N_28368,N_21752,N_23736);
and U28369 (N_28369,N_22580,N_21704);
nand U28370 (N_28370,N_22514,N_21874);
nand U28371 (N_28371,N_20162,N_24450);
nor U28372 (N_28372,N_21894,N_24763);
nor U28373 (N_28373,N_23087,N_23003);
xor U28374 (N_28374,N_21059,N_23463);
or U28375 (N_28375,N_22528,N_24111);
xor U28376 (N_28376,N_20993,N_24325);
or U28377 (N_28377,N_24089,N_20825);
nand U28378 (N_28378,N_24642,N_24788);
nor U28379 (N_28379,N_20141,N_22620);
nor U28380 (N_28380,N_21976,N_21273);
xnor U28381 (N_28381,N_22345,N_21070);
and U28382 (N_28382,N_22706,N_20049);
or U28383 (N_28383,N_24657,N_21475);
nor U28384 (N_28384,N_24233,N_20273);
or U28385 (N_28385,N_20129,N_22267);
or U28386 (N_28386,N_21508,N_20403);
xnor U28387 (N_28387,N_24312,N_20851);
and U28388 (N_28388,N_21530,N_20043);
xnor U28389 (N_28389,N_22933,N_23288);
xor U28390 (N_28390,N_20072,N_20928);
and U28391 (N_28391,N_23213,N_22852);
nand U28392 (N_28392,N_24654,N_20230);
and U28393 (N_28393,N_21980,N_20308);
xor U28394 (N_28394,N_20242,N_22414);
nand U28395 (N_28395,N_24641,N_21927);
xnor U28396 (N_28396,N_24388,N_24868);
or U28397 (N_28397,N_24749,N_24464);
nand U28398 (N_28398,N_24843,N_21398);
and U28399 (N_28399,N_23715,N_24320);
nand U28400 (N_28400,N_22380,N_22731);
or U28401 (N_28401,N_20394,N_20164);
nand U28402 (N_28402,N_23529,N_21387);
nand U28403 (N_28403,N_20845,N_20136);
or U28404 (N_28404,N_21059,N_23587);
xor U28405 (N_28405,N_21646,N_23542);
nand U28406 (N_28406,N_24465,N_21427);
and U28407 (N_28407,N_20220,N_24956);
and U28408 (N_28408,N_20344,N_24494);
nand U28409 (N_28409,N_23103,N_20081);
or U28410 (N_28410,N_24117,N_22648);
xnor U28411 (N_28411,N_24153,N_24828);
or U28412 (N_28412,N_23205,N_22813);
nor U28413 (N_28413,N_22677,N_23415);
nor U28414 (N_28414,N_23547,N_22890);
or U28415 (N_28415,N_22823,N_23270);
or U28416 (N_28416,N_24507,N_24956);
nand U28417 (N_28417,N_24810,N_22208);
and U28418 (N_28418,N_24700,N_23879);
and U28419 (N_28419,N_24774,N_24081);
and U28420 (N_28420,N_23777,N_22827);
or U28421 (N_28421,N_21435,N_21666);
nor U28422 (N_28422,N_23044,N_21286);
nand U28423 (N_28423,N_22612,N_20576);
or U28424 (N_28424,N_22416,N_24818);
or U28425 (N_28425,N_22024,N_20977);
or U28426 (N_28426,N_24225,N_23199);
nand U28427 (N_28427,N_21156,N_21128);
nor U28428 (N_28428,N_21808,N_24010);
nand U28429 (N_28429,N_21097,N_24033);
or U28430 (N_28430,N_21365,N_23341);
nor U28431 (N_28431,N_20063,N_23063);
and U28432 (N_28432,N_20406,N_24018);
nor U28433 (N_28433,N_22430,N_21014);
or U28434 (N_28434,N_20102,N_21883);
nor U28435 (N_28435,N_24216,N_23344);
nor U28436 (N_28436,N_22760,N_20140);
and U28437 (N_28437,N_24973,N_21285);
xnor U28438 (N_28438,N_21194,N_21152);
xnor U28439 (N_28439,N_22277,N_24171);
and U28440 (N_28440,N_24122,N_24332);
and U28441 (N_28441,N_22766,N_23780);
xor U28442 (N_28442,N_20168,N_21346);
and U28443 (N_28443,N_22805,N_20294);
and U28444 (N_28444,N_20077,N_21963);
nand U28445 (N_28445,N_20991,N_20302);
nor U28446 (N_28446,N_23313,N_20450);
or U28447 (N_28447,N_22032,N_22745);
nor U28448 (N_28448,N_21939,N_24162);
nand U28449 (N_28449,N_20038,N_23702);
nand U28450 (N_28450,N_21986,N_22932);
xnor U28451 (N_28451,N_23389,N_20776);
nand U28452 (N_28452,N_22523,N_21153);
nor U28453 (N_28453,N_24009,N_21133);
or U28454 (N_28454,N_24374,N_20664);
nand U28455 (N_28455,N_20142,N_23161);
or U28456 (N_28456,N_23836,N_22589);
nor U28457 (N_28457,N_22617,N_24375);
nor U28458 (N_28458,N_23551,N_23497);
nand U28459 (N_28459,N_23086,N_22586);
nor U28460 (N_28460,N_22085,N_22059);
nand U28461 (N_28461,N_22547,N_23328);
xor U28462 (N_28462,N_22140,N_21874);
or U28463 (N_28463,N_24851,N_24438);
and U28464 (N_28464,N_22984,N_23759);
nand U28465 (N_28465,N_21997,N_21871);
or U28466 (N_28466,N_23216,N_24127);
nor U28467 (N_28467,N_21497,N_21397);
nor U28468 (N_28468,N_22799,N_24717);
nor U28469 (N_28469,N_21323,N_24078);
xor U28470 (N_28470,N_21782,N_20669);
nand U28471 (N_28471,N_21704,N_20004);
nor U28472 (N_28472,N_23444,N_20832);
nor U28473 (N_28473,N_20280,N_24085);
nor U28474 (N_28474,N_21693,N_21338);
xnor U28475 (N_28475,N_20448,N_22342);
nand U28476 (N_28476,N_24158,N_24375);
xnor U28477 (N_28477,N_23390,N_22904);
and U28478 (N_28478,N_22566,N_24480);
xor U28479 (N_28479,N_21359,N_24862);
and U28480 (N_28480,N_23932,N_23469);
nand U28481 (N_28481,N_21962,N_24728);
xnor U28482 (N_28482,N_22229,N_22643);
and U28483 (N_28483,N_21748,N_24762);
xnor U28484 (N_28484,N_24355,N_22832);
nand U28485 (N_28485,N_24688,N_20902);
xnor U28486 (N_28486,N_20088,N_20669);
nand U28487 (N_28487,N_24668,N_23673);
nand U28488 (N_28488,N_21464,N_23237);
or U28489 (N_28489,N_21963,N_24030);
and U28490 (N_28490,N_24045,N_23376);
nor U28491 (N_28491,N_24831,N_22895);
nor U28492 (N_28492,N_22925,N_24927);
nor U28493 (N_28493,N_21479,N_21448);
or U28494 (N_28494,N_22887,N_22893);
nand U28495 (N_28495,N_20245,N_21959);
or U28496 (N_28496,N_20813,N_24412);
or U28497 (N_28497,N_24985,N_20558);
or U28498 (N_28498,N_21570,N_24717);
or U28499 (N_28499,N_24504,N_24279);
or U28500 (N_28500,N_23863,N_22020);
or U28501 (N_28501,N_22152,N_24409);
nor U28502 (N_28502,N_24104,N_21201);
nand U28503 (N_28503,N_20109,N_20073);
or U28504 (N_28504,N_24723,N_21736);
nor U28505 (N_28505,N_21897,N_23633);
nand U28506 (N_28506,N_23029,N_22666);
xor U28507 (N_28507,N_24029,N_21719);
and U28508 (N_28508,N_23567,N_24840);
and U28509 (N_28509,N_24984,N_24362);
and U28510 (N_28510,N_23425,N_22106);
and U28511 (N_28511,N_23656,N_22777);
or U28512 (N_28512,N_22020,N_21347);
nor U28513 (N_28513,N_21566,N_23429);
xnor U28514 (N_28514,N_20904,N_21172);
and U28515 (N_28515,N_20628,N_24821);
and U28516 (N_28516,N_21013,N_24536);
nand U28517 (N_28517,N_20068,N_21545);
xor U28518 (N_28518,N_23506,N_20375);
and U28519 (N_28519,N_24527,N_24590);
or U28520 (N_28520,N_22853,N_21328);
or U28521 (N_28521,N_24138,N_24534);
nand U28522 (N_28522,N_21460,N_23786);
nor U28523 (N_28523,N_23849,N_24408);
xor U28524 (N_28524,N_20161,N_24165);
nor U28525 (N_28525,N_22907,N_20919);
nor U28526 (N_28526,N_20508,N_20118);
or U28527 (N_28527,N_20524,N_21294);
nor U28528 (N_28528,N_24608,N_21242);
nand U28529 (N_28529,N_22412,N_24090);
xnor U28530 (N_28530,N_21152,N_22308);
xnor U28531 (N_28531,N_22684,N_20118);
or U28532 (N_28532,N_24148,N_21288);
nand U28533 (N_28533,N_22569,N_22755);
nand U28534 (N_28534,N_22754,N_24101);
or U28535 (N_28535,N_24441,N_21988);
nor U28536 (N_28536,N_20527,N_23005);
or U28537 (N_28537,N_24572,N_23187);
or U28538 (N_28538,N_20859,N_24525);
nand U28539 (N_28539,N_23870,N_21171);
or U28540 (N_28540,N_24457,N_20862);
or U28541 (N_28541,N_23810,N_23881);
and U28542 (N_28542,N_22727,N_23602);
nor U28543 (N_28543,N_23788,N_21249);
and U28544 (N_28544,N_22300,N_20318);
nor U28545 (N_28545,N_22781,N_22863);
nor U28546 (N_28546,N_20273,N_23554);
or U28547 (N_28547,N_23045,N_22389);
xor U28548 (N_28548,N_21831,N_21751);
nor U28549 (N_28549,N_20267,N_21582);
nand U28550 (N_28550,N_23193,N_21708);
xor U28551 (N_28551,N_21666,N_20268);
nand U28552 (N_28552,N_24732,N_24479);
or U28553 (N_28553,N_23709,N_21312);
nand U28554 (N_28554,N_24580,N_20416);
nand U28555 (N_28555,N_24745,N_22784);
xor U28556 (N_28556,N_21978,N_23038);
and U28557 (N_28557,N_23959,N_24683);
nand U28558 (N_28558,N_23217,N_20923);
nor U28559 (N_28559,N_22308,N_23422);
or U28560 (N_28560,N_20250,N_24465);
nor U28561 (N_28561,N_24163,N_22328);
nand U28562 (N_28562,N_22325,N_24016);
or U28563 (N_28563,N_20740,N_23289);
and U28564 (N_28564,N_21184,N_21156);
nand U28565 (N_28565,N_21859,N_21178);
xnor U28566 (N_28566,N_22752,N_22536);
xor U28567 (N_28567,N_24070,N_21903);
or U28568 (N_28568,N_23713,N_20849);
or U28569 (N_28569,N_21801,N_22606);
or U28570 (N_28570,N_20999,N_20326);
nor U28571 (N_28571,N_22835,N_22774);
or U28572 (N_28572,N_21566,N_20923);
nand U28573 (N_28573,N_21617,N_20215);
nor U28574 (N_28574,N_23700,N_23597);
nor U28575 (N_28575,N_22636,N_21512);
nor U28576 (N_28576,N_20477,N_22036);
or U28577 (N_28577,N_22999,N_24758);
and U28578 (N_28578,N_23813,N_24100);
nand U28579 (N_28579,N_24754,N_20445);
xnor U28580 (N_28580,N_24733,N_24292);
nor U28581 (N_28581,N_24574,N_22708);
nand U28582 (N_28582,N_20121,N_23990);
nand U28583 (N_28583,N_20120,N_23805);
or U28584 (N_28584,N_21437,N_22532);
nand U28585 (N_28585,N_23540,N_23250);
nor U28586 (N_28586,N_22154,N_22417);
xor U28587 (N_28587,N_22908,N_20426);
xor U28588 (N_28588,N_21265,N_22178);
nand U28589 (N_28589,N_22200,N_24877);
nor U28590 (N_28590,N_23864,N_23497);
or U28591 (N_28591,N_22984,N_21317);
xor U28592 (N_28592,N_24297,N_20718);
and U28593 (N_28593,N_20957,N_22650);
and U28594 (N_28594,N_22864,N_21849);
and U28595 (N_28595,N_23035,N_21678);
nor U28596 (N_28596,N_20839,N_23274);
nand U28597 (N_28597,N_23671,N_21877);
or U28598 (N_28598,N_23058,N_20916);
and U28599 (N_28599,N_23785,N_20490);
nor U28600 (N_28600,N_22161,N_21118);
nor U28601 (N_28601,N_24931,N_22212);
nand U28602 (N_28602,N_22776,N_22015);
nand U28603 (N_28603,N_24601,N_21821);
or U28604 (N_28604,N_20624,N_21009);
and U28605 (N_28605,N_21752,N_21947);
xor U28606 (N_28606,N_21969,N_23108);
nand U28607 (N_28607,N_22611,N_21059);
nor U28608 (N_28608,N_22002,N_23860);
nand U28609 (N_28609,N_24591,N_22163);
nor U28610 (N_28610,N_23585,N_21726);
nor U28611 (N_28611,N_20188,N_20618);
nor U28612 (N_28612,N_22781,N_23065);
or U28613 (N_28613,N_23666,N_23470);
xor U28614 (N_28614,N_22016,N_21989);
and U28615 (N_28615,N_21897,N_24780);
or U28616 (N_28616,N_21796,N_22744);
xnor U28617 (N_28617,N_22097,N_24441);
xor U28618 (N_28618,N_23425,N_20126);
nor U28619 (N_28619,N_24829,N_21456);
and U28620 (N_28620,N_23817,N_21690);
nor U28621 (N_28621,N_21253,N_23127);
xnor U28622 (N_28622,N_23643,N_20262);
xor U28623 (N_28623,N_22771,N_24241);
nand U28624 (N_28624,N_24086,N_23987);
nand U28625 (N_28625,N_24930,N_24986);
or U28626 (N_28626,N_21609,N_21181);
nor U28627 (N_28627,N_20861,N_22518);
nor U28628 (N_28628,N_21819,N_20823);
nand U28629 (N_28629,N_22182,N_20476);
nor U28630 (N_28630,N_20179,N_21228);
and U28631 (N_28631,N_24658,N_24514);
and U28632 (N_28632,N_20628,N_24240);
nand U28633 (N_28633,N_23057,N_23006);
nand U28634 (N_28634,N_20501,N_20050);
nor U28635 (N_28635,N_23654,N_20611);
xnor U28636 (N_28636,N_21010,N_23869);
or U28637 (N_28637,N_20973,N_21640);
and U28638 (N_28638,N_21933,N_21547);
nand U28639 (N_28639,N_23773,N_24882);
xnor U28640 (N_28640,N_22855,N_23328);
and U28641 (N_28641,N_22672,N_24067);
xnor U28642 (N_28642,N_24047,N_24907);
or U28643 (N_28643,N_24905,N_22586);
nor U28644 (N_28644,N_21266,N_23431);
nor U28645 (N_28645,N_20205,N_22234);
and U28646 (N_28646,N_21066,N_24778);
xor U28647 (N_28647,N_23578,N_20903);
nand U28648 (N_28648,N_21920,N_22337);
nor U28649 (N_28649,N_23340,N_21762);
xnor U28650 (N_28650,N_22891,N_24811);
or U28651 (N_28651,N_23993,N_21270);
xor U28652 (N_28652,N_23570,N_23817);
xor U28653 (N_28653,N_22391,N_20578);
xnor U28654 (N_28654,N_24390,N_23654);
xnor U28655 (N_28655,N_21534,N_22084);
nand U28656 (N_28656,N_23703,N_22740);
or U28657 (N_28657,N_24394,N_24858);
nor U28658 (N_28658,N_23767,N_20539);
or U28659 (N_28659,N_23345,N_24437);
xor U28660 (N_28660,N_23525,N_22171);
nand U28661 (N_28661,N_22869,N_23360);
and U28662 (N_28662,N_23028,N_20226);
or U28663 (N_28663,N_23772,N_21159);
nor U28664 (N_28664,N_21268,N_21265);
or U28665 (N_28665,N_21989,N_20229);
nor U28666 (N_28666,N_20434,N_24599);
or U28667 (N_28667,N_23969,N_21959);
xor U28668 (N_28668,N_23476,N_21161);
nand U28669 (N_28669,N_22027,N_22901);
nor U28670 (N_28670,N_21312,N_22751);
nor U28671 (N_28671,N_23439,N_20452);
xnor U28672 (N_28672,N_20240,N_23874);
and U28673 (N_28673,N_20622,N_22182);
nand U28674 (N_28674,N_24119,N_24557);
or U28675 (N_28675,N_20765,N_24822);
xor U28676 (N_28676,N_20603,N_24235);
nor U28677 (N_28677,N_20754,N_21920);
xnor U28678 (N_28678,N_22452,N_20187);
or U28679 (N_28679,N_20254,N_23330);
nand U28680 (N_28680,N_20959,N_24926);
xnor U28681 (N_28681,N_21142,N_21738);
or U28682 (N_28682,N_23180,N_21956);
xnor U28683 (N_28683,N_20736,N_24931);
or U28684 (N_28684,N_24265,N_22002);
nand U28685 (N_28685,N_23720,N_20513);
nand U28686 (N_28686,N_24537,N_23578);
xnor U28687 (N_28687,N_21197,N_22416);
nor U28688 (N_28688,N_23348,N_23276);
nor U28689 (N_28689,N_21632,N_22320);
nand U28690 (N_28690,N_24369,N_21809);
or U28691 (N_28691,N_24638,N_24319);
nand U28692 (N_28692,N_20936,N_20966);
xor U28693 (N_28693,N_21780,N_21036);
nand U28694 (N_28694,N_22883,N_21747);
and U28695 (N_28695,N_20505,N_24105);
nor U28696 (N_28696,N_21056,N_21250);
nand U28697 (N_28697,N_24043,N_21109);
and U28698 (N_28698,N_23812,N_23867);
xor U28699 (N_28699,N_20497,N_23458);
and U28700 (N_28700,N_21390,N_23924);
or U28701 (N_28701,N_22869,N_22202);
nor U28702 (N_28702,N_20035,N_21567);
xor U28703 (N_28703,N_21708,N_22570);
or U28704 (N_28704,N_23900,N_24001);
xor U28705 (N_28705,N_21986,N_21023);
and U28706 (N_28706,N_24634,N_21103);
or U28707 (N_28707,N_21338,N_24035);
nor U28708 (N_28708,N_20653,N_23148);
nor U28709 (N_28709,N_20383,N_20946);
nand U28710 (N_28710,N_23188,N_23888);
or U28711 (N_28711,N_21192,N_23872);
and U28712 (N_28712,N_24782,N_21870);
or U28713 (N_28713,N_20062,N_23321);
nor U28714 (N_28714,N_22277,N_22893);
nand U28715 (N_28715,N_22901,N_21047);
and U28716 (N_28716,N_23777,N_21044);
and U28717 (N_28717,N_24615,N_21355);
xor U28718 (N_28718,N_22354,N_24131);
and U28719 (N_28719,N_24860,N_24163);
nand U28720 (N_28720,N_24477,N_20075);
and U28721 (N_28721,N_22769,N_22167);
nor U28722 (N_28722,N_20550,N_20503);
xor U28723 (N_28723,N_22085,N_22003);
nor U28724 (N_28724,N_24278,N_23285);
nor U28725 (N_28725,N_23064,N_20169);
nor U28726 (N_28726,N_20437,N_20877);
or U28727 (N_28727,N_24728,N_22670);
nor U28728 (N_28728,N_23617,N_22143);
or U28729 (N_28729,N_20027,N_24578);
or U28730 (N_28730,N_20702,N_20177);
and U28731 (N_28731,N_20079,N_23251);
or U28732 (N_28732,N_23355,N_20551);
or U28733 (N_28733,N_24557,N_21483);
or U28734 (N_28734,N_21501,N_24120);
xnor U28735 (N_28735,N_24927,N_23605);
and U28736 (N_28736,N_23928,N_24949);
nor U28737 (N_28737,N_22324,N_20214);
and U28738 (N_28738,N_24047,N_24667);
or U28739 (N_28739,N_24191,N_20360);
nor U28740 (N_28740,N_20845,N_20672);
xor U28741 (N_28741,N_22055,N_20130);
xor U28742 (N_28742,N_20463,N_20942);
or U28743 (N_28743,N_20159,N_21950);
xnor U28744 (N_28744,N_24286,N_24859);
and U28745 (N_28745,N_21460,N_24948);
and U28746 (N_28746,N_21923,N_21785);
or U28747 (N_28747,N_20849,N_23347);
and U28748 (N_28748,N_24135,N_24137);
nand U28749 (N_28749,N_24172,N_22583);
and U28750 (N_28750,N_23922,N_20872);
xnor U28751 (N_28751,N_20629,N_24590);
nor U28752 (N_28752,N_23918,N_24316);
nor U28753 (N_28753,N_22782,N_21656);
xnor U28754 (N_28754,N_22710,N_20073);
nor U28755 (N_28755,N_20452,N_20055);
nand U28756 (N_28756,N_23775,N_24800);
nor U28757 (N_28757,N_24002,N_22905);
nand U28758 (N_28758,N_24122,N_20619);
nor U28759 (N_28759,N_22357,N_21299);
nor U28760 (N_28760,N_23231,N_22973);
xnor U28761 (N_28761,N_20961,N_22704);
nand U28762 (N_28762,N_21049,N_21351);
nor U28763 (N_28763,N_24292,N_20696);
nor U28764 (N_28764,N_23621,N_22899);
and U28765 (N_28765,N_20992,N_21524);
nor U28766 (N_28766,N_23668,N_21218);
xnor U28767 (N_28767,N_20657,N_21966);
and U28768 (N_28768,N_21578,N_21867);
nor U28769 (N_28769,N_23890,N_23218);
nor U28770 (N_28770,N_22991,N_20145);
xor U28771 (N_28771,N_21617,N_20575);
and U28772 (N_28772,N_24363,N_21633);
nand U28773 (N_28773,N_24594,N_21948);
xnor U28774 (N_28774,N_24669,N_21558);
nor U28775 (N_28775,N_21003,N_24916);
nor U28776 (N_28776,N_20388,N_20533);
nor U28777 (N_28777,N_20490,N_21805);
nor U28778 (N_28778,N_22719,N_23618);
nor U28779 (N_28779,N_20218,N_21096);
or U28780 (N_28780,N_22824,N_21826);
or U28781 (N_28781,N_20317,N_22175);
or U28782 (N_28782,N_24615,N_20241);
or U28783 (N_28783,N_21740,N_24240);
and U28784 (N_28784,N_24078,N_20852);
and U28785 (N_28785,N_20267,N_21921);
nand U28786 (N_28786,N_22896,N_21421);
nand U28787 (N_28787,N_22941,N_20572);
or U28788 (N_28788,N_20041,N_21714);
xnor U28789 (N_28789,N_20435,N_20617);
nand U28790 (N_28790,N_21458,N_24643);
nor U28791 (N_28791,N_22133,N_22563);
nand U28792 (N_28792,N_21918,N_23037);
and U28793 (N_28793,N_23314,N_24002);
and U28794 (N_28794,N_23744,N_21356);
nor U28795 (N_28795,N_20701,N_21635);
or U28796 (N_28796,N_24086,N_23734);
nand U28797 (N_28797,N_23943,N_23059);
xnor U28798 (N_28798,N_24736,N_22964);
or U28799 (N_28799,N_23935,N_24954);
or U28800 (N_28800,N_23109,N_22675);
nor U28801 (N_28801,N_23331,N_20218);
nor U28802 (N_28802,N_22148,N_23249);
or U28803 (N_28803,N_23922,N_22600);
xnor U28804 (N_28804,N_22663,N_20175);
and U28805 (N_28805,N_21286,N_21129);
nand U28806 (N_28806,N_21287,N_21497);
nor U28807 (N_28807,N_21946,N_24722);
nor U28808 (N_28808,N_23497,N_23124);
or U28809 (N_28809,N_22616,N_24624);
nand U28810 (N_28810,N_22611,N_22224);
and U28811 (N_28811,N_23535,N_22476);
and U28812 (N_28812,N_24465,N_23098);
nand U28813 (N_28813,N_20244,N_21052);
nor U28814 (N_28814,N_23556,N_21030);
xnor U28815 (N_28815,N_21544,N_20165);
and U28816 (N_28816,N_20288,N_21747);
nor U28817 (N_28817,N_22744,N_24415);
and U28818 (N_28818,N_22689,N_23961);
nand U28819 (N_28819,N_23348,N_23260);
nor U28820 (N_28820,N_21122,N_23652);
nand U28821 (N_28821,N_22010,N_23472);
xor U28822 (N_28822,N_22510,N_21734);
xor U28823 (N_28823,N_24748,N_22353);
nand U28824 (N_28824,N_22676,N_24776);
nor U28825 (N_28825,N_22291,N_24522);
nor U28826 (N_28826,N_24904,N_24993);
xor U28827 (N_28827,N_20281,N_21139);
nand U28828 (N_28828,N_23123,N_20363);
and U28829 (N_28829,N_23419,N_21039);
and U28830 (N_28830,N_23549,N_22522);
nand U28831 (N_28831,N_21170,N_21323);
nand U28832 (N_28832,N_23092,N_23485);
xor U28833 (N_28833,N_21005,N_20147);
nor U28834 (N_28834,N_23907,N_21991);
or U28835 (N_28835,N_24952,N_23940);
nand U28836 (N_28836,N_23662,N_22102);
xor U28837 (N_28837,N_21525,N_20615);
nand U28838 (N_28838,N_24262,N_20975);
xor U28839 (N_28839,N_24981,N_23241);
and U28840 (N_28840,N_22215,N_22207);
nand U28841 (N_28841,N_23820,N_24670);
and U28842 (N_28842,N_21362,N_20110);
or U28843 (N_28843,N_23599,N_21119);
or U28844 (N_28844,N_22927,N_23215);
and U28845 (N_28845,N_20324,N_23027);
nand U28846 (N_28846,N_20713,N_23393);
nor U28847 (N_28847,N_20743,N_23474);
nand U28848 (N_28848,N_24988,N_24502);
xor U28849 (N_28849,N_21308,N_22717);
xnor U28850 (N_28850,N_20256,N_23757);
nor U28851 (N_28851,N_20085,N_22164);
or U28852 (N_28852,N_24563,N_22356);
and U28853 (N_28853,N_24111,N_24551);
nand U28854 (N_28854,N_21943,N_22598);
xor U28855 (N_28855,N_21282,N_23336);
nand U28856 (N_28856,N_21394,N_21322);
and U28857 (N_28857,N_22926,N_22762);
or U28858 (N_28858,N_21818,N_23267);
and U28859 (N_28859,N_23651,N_20642);
and U28860 (N_28860,N_20382,N_22591);
or U28861 (N_28861,N_22381,N_24814);
or U28862 (N_28862,N_21413,N_22596);
nand U28863 (N_28863,N_24424,N_20458);
and U28864 (N_28864,N_24562,N_24635);
or U28865 (N_28865,N_20572,N_20705);
nand U28866 (N_28866,N_24823,N_20409);
and U28867 (N_28867,N_20764,N_21142);
or U28868 (N_28868,N_20142,N_21590);
xnor U28869 (N_28869,N_22154,N_23469);
nand U28870 (N_28870,N_22708,N_20828);
nor U28871 (N_28871,N_22146,N_20719);
nand U28872 (N_28872,N_22764,N_20076);
nand U28873 (N_28873,N_21194,N_22143);
nor U28874 (N_28874,N_23585,N_21144);
and U28875 (N_28875,N_24801,N_21311);
or U28876 (N_28876,N_22469,N_21342);
nand U28877 (N_28877,N_23790,N_22536);
nand U28878 (N_28878,N_22703,N_22273);
or U28879 (N_28879,N_20737,N_20297);
nand U28880 (N_28880,N_21418,N_20934);
xnor U28881 (N_28881,N_21572,N_20969);
xnor U28882 (N_28882,N_20538,N_22914);
or U28883 (N_28883,N_23159,N_21920);
xnor U28884 (N_28884,N_21430,N_20806);
or U28885 (N_28885,N_24010,N_21210);
xnor U28886 (N_28886,N_23662,N_21909);
or U28887 (N_28887,N_22689,N_20098);
nor U28888 (N_28888,N_23788,N_21584);
xnor U28889 (N_28889,N_24421,N_24168);
nand U28890 (N_28890,N_23260,N_21674);
xnor U28891 (N_28891,N_21666,N_23677);
xnor U28892 (N_28892,N_20203,N_24031);
and U28893 (N_28893,N_24930,N_21190);
xor U28894 (N_28894,N_24634,N_22015);
or U28895 (N_28895,N_24999,N_20849);
and U28896 (N_28896,N_20553,N_23360);
xor U28897 (N_28897,N_23272,N_20693);
nand U28898 (N_28898,N_21119,N_21971);
xor U28899 (N_28899,N_20376,N_22096);
nand U28900 (N_28900,N_24318,N_23766);
or U28901 (N_28901,N_20348,N_20746);
nor U28902 (N_28902,N_23303,N_23834);
nand U28903 (N_28903,N_22594,N_20557);
nor U28904 (N_28904,N_22428,N_23798);
nor U28905 (N_28905,N_24412,N_20207);
or U28906 (N_28906,N_20015,N_21033);
and U28907 (N_28907,N_22089,N_20564);
xnor U28908 (N_28908,N_22815,N_20736);
xor U28909 (N_28909,N_21524,N_21588);
or U28910 (N_28910,N_24921,N_23156);
and U28911 (N_28911,N_24210,N_22455);
xnor U28912 (N_28912,N_21633,N_23560);
xnor U28913 (N_28913,N_20897,N_21912);
nor U28914 (N_28914,N_21281,N_22816);
or U28915 (N_28915,N_23563,N_22315);
xor U28916 (N_28916,N_20789,N_21250);
nor U28917 (N_28917,N_24961,N_22320);
nand U28918 (N_28918,N_24849,N_23309);
nor U28919 (N_28919,N_21111,N_22072);
or U28920 (N_28920,N_22257,N_20355);
xor U28921 (N_28921,N_20620,N_21284);
nor U28922 (N_28922,N_23979,N_23657);
xor U28923 (N_28923,N_21841,N_23526);
or U28924 (N_28924,N_20747,N_22658);
nor U28925 (N_28925,N_22818,N_24025);
nor U28926 (N_28926,N_22487,N_22006);
and U28927 (N_28927,N_21603,N_20382);
and U28928 (N_28928,N_21951,N_23273);
or U28929 (N_28929,N_23720,N_24393);
and U28930 (N_28930,N_24269,N_22842);
nand U28931 (N_28931,N_23711,N_22595);
nor U28932 (N_28932,N_23744,N_23186);
and U28933 (N_28933,N_22405,N_24885);
nor U28934 (N_28934,N_20903,N_20471);
nand U28935 (N_28935,N_21730,N_23636);
nor U28936 (N_28936,N_23094,N_22074);
and U28937 (N_28937,N_22355,N_22291);
nor U28938 (N_28938,N_21686,N_20061);
nor U28939 (N_28939,N_23421,N_24387);
or U28940 (N_28940,N_21538,N_22101);
nand U28941 (N_28941,N_20049,N_22082);
and U28942 (N_28942,N_24289,N_24731);
xnor U28943 (N_28943,N_20135,N_22952);
xor U28944 (N_28944,N_23956,N_22080);
and U28945 (N_28945,N_24720,N_23484);
nor U28946 (N_28946,N_23173,N_24234);
or U28947 (N_28947,N_21369,N_24686);
or U28948 (N_28948,N_21949,N_22258);
xor U28949 (N_28949,N_23358,N_21077);
nor U28950 (N_28950,N_24188,N_24613);
or U28951 (N_28951,N_23186,N_21517);
xnor U28952 (N_28952,N_22433,N_22843);
nor U28953 (N_28953,N_21741,N_22894);
nor U28954 (N_28954,N_20990,N_24573);
and U28955 (N_28955,N_20317,N_24591);
xor U28956 (N_28956,N_21879,N_24762);
xor U28957 (N_28957,N_24260,N_23220);
or U28958 (N_28958,N_21029,N_21263);
nand U28959 (N_28959,N_21434,N_23699);
nor U28960 (N_28960,N_23135,N_20434);
or U28961 (N_28961,N_21289,N_24853);
and U28962 (N_28962,N_24835,N_24464);
xnor U28963 (N_28963,N_24040,N_21814);
or U28964 (N_28964,N_20091,N_21527);
and U28965 (N_28965,N_21622,N_23930);
or U28966 (N_28966,N_21205,N_20926);
xnor U28967 (N_28967,N_22078,N_23507);
xnor U28968 (N_28968,N_22165,N_23428);
and U28969 (N_28969,N_24537,N_21410);
nand U28970 (N_28970,N_23399,N_22696);
or U28971 (N_28971,N_22912,N_24408);
xor U28972 (N_28972,N_24178,N_23241);
nand U28973 (N_28973,N_21574,N_20874);
nor U28974 (N_28974,N_22954,N_24046);
nor U28975 (N_28975,N_20418,N_22710);
nor U28976 (N_28976,N_20708,N_23081);
or U28977 (N_28977,N_22835,N_20831);
nand U28978 (N_28978,N_21630,N_24457);
and U28979 (N_28979,N_21948,N_23199);
xor U28980 (N_28980,N_24936,N_22701);
xnor U28981 (N_28981,N_24877,N_21771);
and U28982 (N_28982,N_22387,N_24969);
and U28983 (N_28983,N_20521,N_23505);
nand U28984 (N_28984,N_24541,N_24980);
nand U28985 (N_28985,N_20793,N_22594);
xor U28986 (N_28986,N_24572,N_24695);
nor U28987 (N_28987,N_22896,N_22634);
and U28988 (N_28988,N_22728,N_21683);
nand U28989 (N_28989,N_24403,N_23185);
nand U28990 (N_28990,N_21303,N_21627);
and U28991 (N_28991,N_20620,N_21201);
nand U28992 (N_28992,N_23165,N_23756);
xor U28993 (N_28993,N_23706,N_23771);
or U28994 (N_28994,N_20095,N_23261);
nand U28995 (N_28995,N_24144,N_23116);
nor U28996 (N_28996,N_21665,N_20161);
xor U28997 (N_28997,N_24580,N_22073);
nand U28998 (N_28998,N_23259,N_20468);
and U28999 (N_28999,N_24292,N_20957);
nor U29000 (N_29000,N_23411,N_21964);
xor U29001 (N_29001,N_20577,N_24515);
and U29002 (N_29002,N_22107,N_23079);
nor U29003 (N_29003,N_23090,N_21062);
or U29004 (N_29004,N_23640,N_20952);
and U29005 (N_29005,N_24482,N_22337);
nand U29006 (N_29006,N_21494,N_23997);
or U29007 (N_29007,N_22045,N_21717);
nand U29008 (N_29008,N_23492,N_23350);
or U29009 (N_29009,N_22534,N_21237);
xor U29010 (N_29010,N_21120,N_20817);
xnor U29011 (N_29011,N_22346,N_20536);
xnor U29012 (N_29012,N_23404,N_24065);
xor U29013 (N_29013,N_24370,N_20137);
and U29014 (N_29014,N_21274,N_21485);
xor U29015 (N_29015,N_21201,N_22956);
xnor U29016 (N_29016,N_21429,N_21517);
and U29017 (N_29017,N_21515,N_24196);
or U29018 (N_29018,N_21562,N_22319);
xor U29019 (N_29019,N_23485,N_23869);
or U29020 (N_29020,N_23857,N_23426);
or U29021 (N_29021,N_21906,N_20837);
nand U29022 (N_29022,N_21458,N_24694);
and U29023 (N_29023,N_22348,N_23732);
xnor U29024 (N_29024,N_22506,N_20833);
or U29025 (N_29025,N_22520,N_22352);
or U29026 (N_29026,N_20758,N_21065);
nor U29027 (N_29027,N_24677,N_22153);
nor U29028 (N_29028,N_21076,N_21646);
nor U29029 (N_29029,N_20699,N_23075);
nand U29030 (N_29030,N_24035,N_22239);
nor U29031 (N_29031,N_24453,N_24842);
xnor U29032 (N_29032,N_20087,N_20040);
and U29033 (N_29033,N_23820,N_20555);
nand U29034 (N_29034,N_20153,N_22955);
and U29035 (N_29035,N_21334,N_24805);
and U29036 (N_29036,N_24150,N_22013);
and U29037 (N_29037,N_20784,N_24985);
and U29038 (N_29038,N_23595,N_24934);
nor U29039 (N_29039,N_20788,N_23953);
and U29040 (N_29040,N_21697,N_24233);
or U29041 (N_29041,N_23267,N_21506);
or U29042 (N_29042,N_20743,N_22768);
nor U29043 (N_29043,N_20554,N_21218);
nor U29044 (N_29044,N_24714,N_22625);
nand U29045 (N_29045,N_23591,N_21565);
and U29046 (N_29046,N_22088,N_22142);
xor U29047 (N_29047,N_22263,N_20028);
nor U29048 (N_29048,N_21360,N_22463);
and U29049 (N_29049,N_20308,N_21826);
xor U29050 (N_29050,N_23488,N_24902);
or U29051 (N_29051,N_22958,N_23697);
and U29052 (N_29052,N_24167,N_23039);
xor U29053 (N_29053,N_24453,N_23610);
xnor U29054 (N_29054,N_24978,N_20829);
nor U29055 (N_29055,N_24798,N_21023);
or U29056 (N_29056,N_22225,N_22979);
or U29057 (N_29057,N_20406,N_24728);
xor U29058 (N_29058,N_23618,N_21023);
xnor U29059 (N_29059,N_23286,N_20935);
or U29060 (N_29060,N_22927,N_22722);
and U29061 (N_29061,N_21854,N_22558);
nand U29062 (N_29062,N_23441,N_21759);
and U29063 (N_29063,N_23136,N_23037);
nand U29064 (N_29064,N_20960,N_21125);
xor U29065 (N_29065,N_20340,N_21711);
xor U29066 (N_29066,N_24866,N_24792);
nor U29067 (N_29067,N_21692,N_20460);
xnor U29068 (N_29068,N_24259,N_20525);
and U29069 (N_29069,N_23516,N_22410);
nor U29070 (N_29070,N_20511,N_22178);
xnor U29071 (N_29071,N_24300,N_24514);
xor U29072 (N_29072,N_20544,N_22926);
and U29073 (N_29073,N_22493,N_24936);
xor U29074 (N_29074,N_21007,N_21173);
or U29075 (N_29075,N_24320,N_21060);
nand U29076 (N_29076,N_20186,N_24858);
or U29077 (N_29077,N_22775,N_23126);
nor U29078 (N_29078,N_21487,N_22608);
nor U29079 (N_29079,N_21064,N_21072);
nor U29080 (N_29080,N_21390,N_24460);
or U29081 (N_29081,N_22762,N_21961);
nor U29082 (N_29082,N_22361,N_23842);
or U29083 (N_29083,N_23137,N_24775);
nor U29084 (N_29084,N_20760,N_22387);
nand U29085 (N_29085,N_22767,N_23576);
or U29086 (N_29086,N_22284,N_20603);
and U29087 (N_29087,N_22473,N_22195);
or U29088 (N_29088,N_21283,N_24605);
xor U29089 (N_29089,N_23303,N_23285);
nand U29090 (N_29090,N_20383,N_21571);
nor U29091 (N_29091,N_24937,N_20942);
xor U29092 (N_29092,N_24622,N_21764);
nor U29093 (N_29093,N_22831,N_21824);
nor U29094 (N_29094,N_21992,N_22757);
nand U29095 (N_29095,N_21435,N_20708);
nand U29096 (N_29096,N_23976,N_20443);
or U29097 (N_29097,N_24904,N_21738);
nor U29098 (N_29098,N_20186,N_23799);
or U29099 (N_29099,N_21406,N_22403);
xnor U29100 (N_29100,N_20704,N_23487);
or U29101 (N_29101,N_24138,N_20861);
xnor U29102 (N_29102,N_22060,N_22649);
xnor U29103 (N_29103,N_22228,N_21545);
nor U29104 (N_29104,N_22872,N_22916);
xnor U29105 (N_29105,N_24919,N_20538);
xnor U29106 (N_29106,N_22573,N_24369);
and U29107 (N_29107,N_24523,N_20474);
and U29108 (N_29108,N_21260,N_20274);
xnor U29109 (N_29109,N_22697,N_23858);
nor U29110 (N_29110,N_20521,N_22885);
nand U29111 (N_29111,N_23676,N_20607);
nor U29112 (N_29112,N_21066,N_21437);
and U29113 (N_29113,N_24427,N_23448);
or U29114 (N_29114,N_20065,N_24137);
nand U29115 (N_29115,N_22523,N_21955);
nand U29116 (N_29116,N_21415,N_21864);
nand U29117 (N_29117,N_23088,N_21882);
xnor U29118 (N_29118,N_20006,N_23362);
xor U29119 (N_29119,N_20432,N_24175);
nor U29120 (N_29120,N_22718,N_24459);
or U29121 (N_29121,N_21647,N_22175);
nand U29122 (N_29122,N_21077,N_21583);
xor U29123 (N_29123,N_21174,N_21895);
xor U29124 (N_29124,N_24911,N_20269);
nand U29125 (N_29125,N_20018,N_24037);
nand U29126 (N_29126,N_23202,N_20877);
and U29127 (N_29127,N_24090,N_23357);
nor U29128 (N_29128,N_23701,N_20446);
nor U29129 (N_29129,N_22114,N_22861);
nand U29130 (N_29130,N_21168,N_23546);
and U29131 (N_29131,N_20425,N_21634);
and U29132 (N_29132,N_23779,N_20942);
or U29133 (N_29133,N_23735,N_22926);
and U29134 (N_29134,N_24237,N_24282);
and U29135 (N_29135,N_20649,N_24363);
and U29136 (N_29136,N_20248,N_24073);
or U29137 (N_29137,N_23844,N_24537);
nand U29138 (N_29138,N_22681,N_21733);
xor U29139 (N_29139,N_24686,N_22041);
nand U29140 (N_29140,N_24049,N_23259);
nor U29141 (N_29141,N_23481,N_20319);
and U29142 (N_29142,N_22782,N_23009);
xor U29143 (N_29143,N_22723,N_23870);
and U29144 (N_29144,N_22436,N_22138);
or U29145 (N_29145,N_20015,N_21856);
nor U29146 (N_29146,N_24495,N_22871);
or U29147 (N_29147,N_22439,N_20799);
or U29148 (N_29148,N_21726,N_21628);
and U29149 (N_29149,N_22829,N_21847);
or U29150 (N_29150,N_20662,N_22855);
nand U29151 (N_29151,N_21284,N_22976);
nor U29152 (N_29152,N_22224,N_20069);
or U29153 (N_29153,N_21789,N_24044);
xor U29154 (N_29154,N_23825,N_23740);
xnor U29155 (N_29155,N_24291,N_23748);
or U29156 (N_29156,N_21994,N_20506);
nor U29157 (N_29157,N_20770,N_20139);
xor U29158 (N_29158,N_23869,N_21718);
nor U29159 (N_29159,N_24581,N_21855);
or U29160 (N_29160,N_21802,N_21239);
and U29161 (N_29161,N_24469,N_20207);
and U29162 (N_29162,N_21088,N_21793);
nor U29163 (N_29163,N_24859,N_23094);
or U29164 (N_29164,N_22948,N_20486);
nand U29165 (N_29165,N_22693,N_23683);
and U29166 (N_29166,N_21528,N_22682);
or U29167 (N_29167,N_20689,N_23064);
nor U29168 (N_29168,N_20902,N_20943);
nand U29169 (N_29169,N_20088,N_20860);
xnor U29170 (N_29170,N_20426,N_22157);
xnor U29171 (N_29171,N_24180,N_22316);
xnor U29172 (N_29172,N_23569,N_23160);
xnor U29173 (N_29173,N_23902,N_24060);
xnor U29174 (N_29174,N_20753,N_23098);
nand U29175 (N_29175,N_24934,N_24887);
or U29176 (N_29176,N_24532,N_21899);
and U29177 (N_29177,N_24827,N_20426);
nand U29178 (N_29178,N_20085,N_21891);
or U29179 (N_29179,N_21027,N_23035);
nand U29180 (N_29180,N_24957,N_22655);
and U29181 (N_29181,N_20919,N_22342);
and U29182 (N_29182,N_20733,N_22829);
xor U29183 (N_29183,N_24372,N_21026);
nor U29184 (N_29184,N_21191,N_23476);
xnor U29185 (N_29185,N_21233,N_24629);
xor U29186 (N_29186,N_24367,N_22387);
nor U29187 (N_29187,N_20218,N_24301);
or U29188 (N_29188,N_22091,N_20762);
nand U29189 (N_29189,N_22561,N_23534);
or U29190 (N_29190,N_21311,N_22045);
nand U29191 (N_29191,N_23689,N_21363);
xor U29192 (N_29192,N_23560,N_21717);
xnor U29193 (N_29193,N_22090,N_23071);
and U29194 (N_29194,N_20885,N_24831);
nand U29195 (N_29195,N_20894,N_21839);
and U29196 (N_29196,N_20442,N_20969);
and U29197 (N_29197,N_22721,N_21691);
and U29198 (N_29198,N_22099,N_20432);
nor U29199 (N_29199,N_21369,N_21254);
nor U29200 (N_29200,N_23593,N_22678);
and U29201 (N_29201,N_21811,N_21432);
nor U29202 (N_29202,N_21526,N_21545);
nor U29203 (N_29203,N_20267,N_23897);
and U29204 (N_29204,N_22591,N_23971);
nor U29205 (N_29205,N_24824,N_22220);
nor U29206 (N_29206,N_24811,N_21818);
xnor U29207 (N_29207,N_22491,N_21651);
nor U29208 (N_29208,N_23347,N_23003);
nor U29209 (N_29209,N_23370,N_21489);
and U29210 (N_29210,N_22211,N_22254);
or U29211 (N_29211,N_23307,N_20716);
and U29212 (N_29212,N_21612,N_23499);
xnor U29213 (N_29213,N_24315,N_24939);
nor U29214 (N_29214,N_20422,N_22859);
nand U29215 (N_29215,N_21723,N_22101);
nor U29216 (N_29216,N_20152,N_21142);
nand U29217 (N_29217,N_20519,N_20845);
xor U29218 (N_29218,N_23037,N_23710);
or U29219 (N_29219,N_20924,N_22508);
nand U29220 (N_29220,N_23912,N_20246);
nor U29221 (N_29221,N_23265,N_20229);
nand U29222 (N_29222,N_22711,N_21313);
xor U29223 (N_29223,N_20606,N_20026);
nor U29224 (N_29224,N_24596,N_22526);
xor U29225 (N_29225,N_21403,N_23376);
or U29226 (N_29226,N_20888,N_23475);
and U29227 (N_29227,N_23078,N_24588);
xor U29228 (N_29228,N_20995,N_23602);
or U29229 (N_29229,N_24793,N_21846);
nor U29230 (N_29230,N_23587,N_22044);
and U29231 (N_29231,N_21915,N_22277);
or U29232 (N_29232,N_20176,N_20306);
nor U29233 (N_29233,N_21180,N_23707);
nor U29234 (N_29234,N_24649,N_24789);
nor U29235 (N_29235,N_23978,N_24499);
nor U29236 (N_29236,N_23826,N_22934);
xnor U29237 (N_29237,N_23902,N_21619);
or U29238 (N_29238,N_22569,N_23987);
and U29239 (N_29239,N_20318,N_24584);
xnor U29240 (N_29240,N_23739,N_21443);
xor U29241 (N_29241,N_23510,N_22439);
nor U29242 (N_29242,N_21811,N_23803);
xnor U29243 (N_29243,N_22915,N_20392);
xnor U29244 (N_29244,N_24079,N_23495);
xnor U29245 (N_29245,N_22992,N_21437);
nand U29246 (N_29246,N_22625,N_20093);
nor U29247 (N_29247,N_22992,N_21584);
and U29248 (N_29248,N_22750,N_21853);
nand U29249 (N_29249,N_23732,N_23934);
or U29250 (N_29250,N_21604,N_24992);
or U29251 (N_29251,N_21315,N_23831);
or U29252 (N_29252,N_20704,N_24406);
xor U29253 (N_29253,N_24034,N_22283);
nand U29254 (N_29254,N_22146,N_22079);
nand U29255 (N_29255,N_24320,N_21857);
nand U29256 (N_29256,N_24019,N_21019);
xnor U29257 (N_29257,N_22868,N_23125);
nor U29258 (N_29258,N_22622,N_24033);
xor U29259 (N_29259,N_22029,N_22892);
xor U29260 (N_29260,N_24334,N_22169);
and U29261 (N_29261,N_24706,N_21497);
or U29262 (N_29262,N_21672,N_22376);
xor U29263 (N_29263,N_23014,N_20549);
xnor U29264 (N_29264,N_20217,N_23946);
xor U29265 (N_29265,N_21300,N_22941);
nand U29266 (N_29266,N_20760,N_21066);
nand U29267 (N_29267,N_24459,N_22657);
or U29268 (N_29268,N_20750,N_20280);
xor U29269 (N_29269,N_21552,N_23158);
nand U29270 (N_29270,N_23556,N_22005);
nor U29271 (N_29271,N_22376,N_23254);
or U29272 (N_29272,N_23822,N_21802);
nor U29273 (N_29273,N_21624,N_23324);
or U29274 (N_29274,N_23625,N_22621);
xnor U29275 (N_29275,N_21379,N_20830);
nor U29276 (N_29276,N_21110,N_21909);
xor U29277 (N_29277,N_21627,N_22630);
nor U29278 (N_29278,N_20534,N_22682);
xnor U29279 (N_29279,N_20758,N_23080);
and U29280 (N_29280,N_20911,N_24200);
and U29281 (N_29281,N_23895,N_20290);
nand U29282 (N_29282,N_21522,N_24552);
xor U29283 (N_29283,N_21326,N_20423);
and U29284 (N_29284,N_24331,N_22052);
and U29285 (N_29285,N_21006,N_24380);
xor U29286 (N_29286,N_22098,N_21070);
xor U29287 (N_29287,N_21468,N_20125);
nand U29288 (N_29288,N_21763,N_22817);
and U29289 (N_29289,N_21932,N_20639);
or U29290 (N_29290,N_23392,N_24681);
xnor U29291 (N_29291,N_21277,N_20281);
nand U29292 (N_29292,N_20726,N_24345);
nor U29293 (N_29293,N_20930,N_20442);
xor U29294 (N_29294,N_21707,N_24308);
nor U29295 (N_29295,N_22737,N_23061);
nand U29296 (N_29296,N_23760,N_21586);
nand U29297 (N_29297,N_22968,N_23675);
xor U29298 (N_29298,N_21602,N_22943);
xnor U29299 (N_29299,N_24560,N_22927);
xor U29300 (N_29300,N_23607,N_22341);
nand U29301 (N_29301,N_22341,N_23455);
and U29302 (N_29302,N_20594,N_23659);
nor U29303 (N_29303,N_21319,N_20712);
xnor U29304 (N_29304,N_21618,N_22379);
and U29305 (N_29305,N_24363,N_20820);
and U29306 (N_29306,N_20686,N_24376);
or U29307 (N_29307,N_22473,N_23587);
nand U29308 (N_29308,N_20109,N_20851);
or U29309 (N_29309,N_21934,N_22630);
and U29310 (N_29310,N_24707,N_21739);
and U29311 (N_29311,N_21720,N_21941);
xnor U29312 (N_29312,N_21251,N_21866);
nor U29313 (N_29313,N_23316,N_22254);
nor U29314 (N_29314,N_24045,N_22869);
xor U29315 (N_29315,N_20363,N_22022);
nor U29316 (N_29316,N_20291,N_20211);
and U29317 (N_29317,N_20549,N_21856);
nand U29318 (N_29318,N_21980,N_24270);
and U29319 (N_29319,N_24933,N_24749);
xnor U29320 (N_29320,N_23771,N_22382);
nor U29321 (N_29321,N_24270,N_23554);
xor U29322 (N_29322,N_24517,N_20866);
xnor U29323 (N_29323,N_23176,N_23927);
nor U29324 (N_29324,N_20435,N_23924);
or U29325 (N_29325,N_20458,N_20231);
xor U29326 (N_29326,N_23340,N_21881);
and U29327 (N_29327,N_23951,N_23120);
xnor U29328 (N_29328,N_22418,N_23496);
nor U29329 (N_29329,N_21173,N_21432);
nand U29330 (N_29330,N_21550,N_20734);
xnor U29331 (N_29331,N_24348,N_20655);
or U29332 (N_29332,N_20695,N_21381);
nor U29333 (N_29333,N_24017,N_22596);
nand U29334 (N_29334,N_23816,N_23264);
nor U29335 (N_29335,N_24025,N_20125);
xnor U29336 (N_29336,N_24798,N_22297);
nand U29337 (N_29337,N_22000,N_21723);
xor U29338 (N_29338,N_24339,N_23282);
or U29339 (N_29339,N_23198,N_22459);
or U29340 (N_29340,N_20505,N_22424);
nor U29341 (N_29341,N_21757,N_20094);
nand U29342 (N_29342,N_24588,N_21571);
or U29343 (N_29343,N_23727,N_20046);
xnor U29344 (N_29344,N_20635,N_23781);
nand U29345 (N_29345,N_22687,N_20591);
xnor U29346 (N_29346,N_24221,N_22381);
or U29347 (N_29347,N_24062,N_23893);
or U29348 (N_29348,N_21926,N_23435);
or U29349 (N_29349,N_20244,N_23653);
and U29350 (N_29350,N_23077,N_23942);
nor U29351 (N_29351,N_22781,N_24876);
and U29352 (N_29352,N_22403,N_20591);
or U29353 (N_29353,N_22790,N_24501);
nand U29354 (N_29354,N_22990,N_20694);
or U29355 (N_29355,N_24220,N_23705);
nor U29356 (N_29356,N_22058,N_24277);
or U29357 (N_29357,N_20734,N_20815);
and U29358 (N_29358,N_21456,N_23697);
or U29359 (N_29359,N_24787,N_24897);
xnor U29360 (N_29360,N_22868,N_22042);
and U29361 (N_29361,N_24989,N_20953);
xor U29362 (N_29362,N_24790,N_24502);
nor U29363 (N_29363,N_21253,N_23484);
xor U29364 (N_29364,N_24552,N_21851);
and U29365 (N_29365,N_22979,N_20033);
xor U29366 (N_29366,N_24310,N_23498);
or U29367 (N_29367,N_20734,N_23785);
nand U29368 (N_29368,N_21240,N_24895);
and U29369 (N_29369,N_21216,N_22246);
or U29370 (N_29370,N_20206,N_23172);
nand U29371 (N_29371,N_20271,N_21198);
nor U29372 (N_29372,N_21480,N_23205);
and U29373 (N_29373,N_20684,N_22237);
xnor U29374 (N_29374,N_20737,N_22583);
nand U29375 (N_29375,N_21322,N_20598);
nand U29376 (N_29376,N_22876,N_20730);
xor U29377 (N_29377,N_23721,N_21192);
nand U29378 (N_29378,N_23009,N_20416);
or U29379 (N_29379,N_23425,N_22347);
nor U29380 (N_29380,N_22750,N_22198);
or U29381 (N_29381,N_22943,N_21350);
nand U29382 (N_29382,N_24211,N_23178);
and U29383 (N_29383,N_21135,N_21906);
nand U29384 (N_29384,N_24298,N_22206);
or U29385 (N_29385,N_21241,N_21667);
or U29386 (N_29386,N_24872,N_21783);
nand U29387 (N_29387,N_23849,N_24053);
nor U29388 (N_29388,N_21418,N_21132);
or U29389 (N_29389,N_22984,N_23342);
nor U29390 (N_29390,N_20587,N_21017);
and U29391 (N_29391,N_22983,N_24623);
or U29392 (N_29392,N_23433,N_22656);
or U29393 (N_29393,N_22269,N_23310);
or U29394 (N_29394,N_21256,N_21566);
nor U29395 (N_29395,N_21424,N_21654);
xnor U29396 (N_29396,N_22545,N_24337);
nand U29397 (N_29397,N_23024,N_24466);
nor U29398 (N_29398,N_23653,N_20626);
or U29399 (N_29399,N_20709,N_23717);
or U29400 (N_29400,N_22671,N_22910);
xnor U29401 (N_29401,N_24006,N_23650);
or U29402 (N_29402,N_22266,N_20061);
or U29403 (N_29403,N_22652,N_20789);
and U29404 (N_29404,N_22483,N_24724);
or U29405 (N_29405,N_22640,N_20715);
xor U29406 (N_29406,N_20849,N_21489);
xor U29407 (N_29407,N_20321,N_22832);
xor U29408 (N_29408,N_24329,N_24529);
and U29409 (N_29409,N_22419,N_21333);
nor U29410 (N_29410,N_22085,N_20131);
or U29411 (N_29411,N_21004,N_22995);
xnor U29412 (N_29412,N_23885,N_24256);
xor U29413 (N_29413,N_20466,N_22335);
nand U29414 (N_29414,N_22964,N_23508);
and U29415 (N_29415,N_22923,N_23607);
nand U29416 (N_29416,N_21524,N_21090);
nor U29417 (N_29417,N_20605,N_20374);
xnor U29418 (N_29418,N_22975,N_23114);
nand U29419 (N_29419,N_21352,N_24650);
and U29420 (N_29420,N_21865,N_21628);
nand U29421 (N_29421,N_21422,N_23033);
or U29422 (N_29422,N_20103,N_21414);
and U29423 (N_29423,N_23871,N_23089);
and U29424 (N_29424,N_23231,N_23202);
xor U29425 (N_29425,N_23731,N_22483);
nand U29426 (N_29426,N_24665,N_22470);
and U29427 (N_29427,N_20155,N_20183);
or U29428 (N_29428,N_23373,N_20673);
and U29429 (N_29429,N_23224,N_21112);
xnor U29430 (N_29430,N_22749,N_21617);
nand U29431 (N_29431,N_21451,N_24514);
and U29432 (N_29432,N_22337,N_23299);
or U29433 (N_29433,N_20547,N_21067);
and U29434 (N_29434,N_21087,N_22060);
nor U29435 (N_29435,N_22343,N_23812);
and U29436 (N_29436,N_24855,N_22003);
xnor U29437 (N_29437,N_23528,N_20256);
xnor U29438 (N_29438,N_20205,N_24637);
xor U29439 (N_29439,N_21667,N_23484);
or U29440 (N_29440,N_21906,N_24975);
xor U29441 (N_29441,N_22909,N_20778);
nand U29442 (N_29442,N_20424,N_20036);
xor U29443 (N_29443,N_22214,N_23906);
xnor U29444 (N_29444,N_21129,N_23358);
or U29445 (N_29445,N_22945,N_22534);
and U29446 (N_29446,N_22773,N_24198);
xor U29447 (N_29447,N_24105,N_20895);
or U29448 (N_29448,N_24077,N_21933);
nand U29449 (N_29449,N_22413,N_23802);
nor U29450 (N_29450,N_24524,N_23013);
xnor U29451 (N_29451,N_21306,N_22009);
nand U29452 (N_29452,N_20190,N_24578);
xnor U29453 (N_29453,N_22240,N_24980);
and U29454 (N_29454,N_20470,N_23980);
or U29455 (N_29455,N_22442,N_21880);
nor U29456 (N_29456,N_20127,N_23703);
nand U29457 (N_29457,N_22861,N_20640);
xor U29458 (N_29458,N_23291,N_22359);
xor U29459 (N_29459,N_21382,N_21643);
xnor U29460 (N_29460,N_20213,N_23542);
nand U29461 (N_29461,N_24659,N_23805);
nor U29462 (N_29462,N_24956,N_22036);
and U29463 (N_29463,N_21889,N_20162);
or U29464 (N_29464,N_24734,N_23411);
and U29465 (N_29465,N_24857,N_22063);
or U29466 (N_29466,N_20515,N_22635);
xor U29467 (N_29467,N_21752,N_24182);
xnor U29468 (N_29468,N_21439,N_23590);
and U29469 (N_29469,N_20430,N_23834);
or U29470 (N_29470,N_21351,N_23648);
xnor U29471 (N_29471,N_24150,N_23904);
nand U29472 (N_29472,N_23961,N_21593);
xor U29473 (N_29473,N_22108,N_20785);
nor U29474 (N_29474,N_22024,N_21610);
nand U29475 (N_29475,N_24946,N_20134);
nand U29476 (N_29476,N_24899,N_22740);
nand U29477 (N_29477,N_24626,N_21036);
and U29478 (N_29478,N_22989,N_23063);
xor U29479 (N_29479,N_20692,N_21268);
or U29480 (N_29480,N_20959,N_24360);
xor U29481 (N_29481,N_21871,N_21917);
xor U29482 (N_29482,N_24968,N_20810);
xor U29483 (N_29483,N_21868,N_21165);
nand U29484 (N_29484,N_23038,N_22257);
nor U29485 (N_29485,N_20397,N_20984);
nor U29486 (N_29486,N_23090,N_20345);
or U29487 (N_29487,N_21407,N_23781);
or U29488 (N_29488,N_20271,N_21946);
nand U29489 (N_29489,N_21557,N_20030);
or U29490 (N_29490,N_24171,N_20664);
or U29491 (N_29491,N_20638,N_22836);
xor U29492 (N_29492,N_24486,N_22545);
and U29493 (N_29493,N_22283,N_24598);
xor U29494 (N_29494,N_21142,N_24629);
or U29495 (N_29495,N_24124,N_21844);
and U29496 (N_29496,N_21349,N_24895);
and U29497 (N_29497,N_21299,N_24590);
and U29498 (N_29498,N_21249,N_21583);
nor U29499 (N_29499,N_21672,N_24503);
and U29500 (N_29500,N_24986,N_21300);
nor U29501 (N_29501,N_20510,N_22795);
nand U29502 (N_29502,N_20636,N_22936);
xnor U29503 (N_29503,N_24480,N_23888);
nand U29504 (N_29504,N_20222,N_21429);
or U29505 (N_29505,N_24380,N_23736);
nand U29506 (N_29506,N_22960,N_23009);
or U29507 (N_29507,N_21428,N_22374);
or U29508 (N_29508,N_23148,N_21495);
nand U29509 (N_29509,N_21593,N_22187);
nor U29510 (N_29510,N_21557,N_24049);
nor U29511 (N_29511,N_20113,N_23411);
or U29512 (N_29512,N_24959,N_21705);
nand U29513 (N_29513,N_23526,N_21024);
xnor U29514 (N_29514,N_24178,N_22797);
nand U29515 (N_29515,N_24253,N_21972);
xor U29516 (N_29516,N_20582,N_20193);
xnor U29517 (N_29517,N_23164,N_23801);
or U29518 (N_29518,N_21105,N_20604);
nand U29519 (N_29519,N_21198,N_23089);
nor U29520 (N_29520,N_22240,N_20477);
and U29521 (N_29521,N_23386,N_22272);
or U29522 (N_29522,N_21991,N_20499);
nand U29523 (N_29523,N_23747,N_23714);
and U29524 (N_29524,N_20779,N_23606);
nand U29525 (N_29525,N_20123,N_24000);
and U29526 (N_29526,N_20865,N_23646);
and U29527 (N_29527,N_21169,N_23434);
nor U29528 (N_29528,N_23008,N_24257);
nor U29529 (N_29529,N_24759,N_24407);
or U29530 (N_29530,N_23501,N_22866);
or U29531 (N_29531,N_24207,N_21517);
xnor U29532 (N_29532,N_23243,N_22278);
nor U29533 (N_29533,N_22069,N_24287);
nor U29534 (N_29534,N_23043,N_23988);
or U29535 (N_29535,N_20650,N_22735);
or U29536 (N_29536,N_23677,N_24658);
nor U29537 (N_29537,N_24399,N_23989);
or U29538 (N_29538,N_22187,N_23088);
xnor U29539 (N_29539,N_23614,N_21136);
and U29540 (N_29540,N_24685,N_24148);
nand U29541 (N_29541,N_24484,N_22851);
xor U29542 (N_29542,N_22309,N_21227);
or U29543 (N_29543,N_21988,N_22247);
nor U29544 (N_29544,N_24566,N_21043);
and U29545 (N_29545,N_24413,N_22236);
nor U29546 (N_29546,N_23907,N_21105);
and U29547 (N_29547,N_24518,N_24456);
nor U29548 (N_29548,N_23596,N_21870);
nor U29549 (N_29549,N_20069,N_22847);
nor U29550 (N_29550,N_23025,N_24839);
and U29551 (N_29551,N_20793,N_23826);
nand U29552 (N_29552,N_24132,N_24770);
nor U29553 (N_29553,N_24314,N_24224);
or U29554 (N_29554,N_20297,N_22555);
or U29555 (N_29555,N_23166,N_23876);
nor U29556 (N_29556,N_23165,N_21932);
nand U29557 (N_29557,N_23483,N_22525);
and U29558 (N_29558,N_22747,N_21683);
nand U29559 (N_29559,N_22313,N_23320);
xnor U29560 (N_29560,N_22887,N_21857);
nand U29561 (N_29561,N_21227,N_22959);
or U29562 (N_29562,N_23180,N_24129);
or U29563 (N_29563,N_21228,N_22800);
nor U29564 (N_29564,N_24092,N_22937);
xor U29565 (N_29565,N_20716,N_20625);
nand U29566 (N_29566,N_24037,N_22994);
and U29567 (N_29567,N_24886,N_22165);
nor U29568 (N_29568,N_24846,N_23227);
xnor U29569 (N_29569,N_24105,N_23437);
nand U29570 (N_29570,N_22878,N_20602);
or U29571 (N_29571,N_24467,N_22420);
nor U29572 (N_29572,N_23262,N_21736);
xor U29573 (N_29573,N_24807,N_20730);
nand U29574 (N_29574,N_21455,N_23162);
nand U29575 (N_29575,N_24791,N_22810);
nand U29576 (N_29576,N_24466,N_23209);
xnor U29577 (N_29577,N_20728,N_23428);
nand U29578 (N_29578,N_24564,N_21081);
and U29579 (N_29579,N_21140,N_24814);
nand U29580 (N_29580,N_20061,N_23088);
and U29581 (N_29581,N_24299,N_20903);
nor U29582 (N_29582,N_20622,N_21174);
or U29583 (N_29583,N_24096,N_24890);
nor U29584 (N_29584,N_24625,N_22149);
xnor U29585 (N_29585,N_24912,N_21331);
nand U29586 (N_29586,N_22377,N_20012);
or U29587 (N_29587,N_20615,N_22991);
nand U29588 (N_29588,N_20943,N_24810);
or U29589 (N_29589,N_23627,N_24202);
or U29590 (N_29590,N_21591,N_23572);
and U29591 (N_29591,N_20452,N_22293);
or U29592 (N_29592,N_21217,N_23830);
and U29593 (N_29593,N_23229,N_23990);
nand U29594 (N_29594,N_23117,N_24474);
nand U29595 (N_29595,N_21898,N_22324);
nor U29596 (N_29596,N_22370,N_24714);
nand U29597 (N_29597,N_24065,N_22512);
xnor U29598 (N_29598,N_24144,N_24405);
xnor U29599 (N_29599,N_20624,N_20441);
xnor U29600 (N_29600,N_21801,N_22159);
or U29601 (N_29601,N_24429,N_24512);
or U29602 (N_29602,N_24261,N_23305);
nand U29603 (N_29603,N_24669,N_21122);
and U29604 (N_29604,N_20755,N_22608);
nand U29605 (N_29605,N_20608,N_23822);
and U29606 (N_29606,N_23102,N_24321);
or U29607 (N_29607,N_20428,N_24451);
and U29608 (N_29608,N_22216,N_23630);
and U29609 (N_29609,N_24415,N_24553);
or U29610 (N_29610,N_21914,N_21225);
and U29611 (N_29611,N_20328,N_20349);
nor U29612 (N_29612,N_22591,N_23010);
nand U29613 (N_29613,N_23109,N_23113);
nand U29614 (N_29614,N_21062,N_22612);
or U29615 (N_29615,N_23596,N_23492);
and U29616 (N_29616,N_20878,N_20829);
or U29617 (N_29617,N_22360,N_20950);
nand U29618 (N_29618,N_23082,N_23859);
nand U29619 (N_29619,N_20638,N_21041);
xor U29620 (N_29620,N_20988,N_24147);
xnor U29621 (N_29621,N_22510,N_20609);
or U29622 (N_29622,N_22738,N_22170);
and U29623 (N_29623,N_20875,N_23215);
or U29624 (N_29624,N_24124,N_24818);
xnor U29625 (N_29625,N_24514,N_22771);
nor U29626 (N_29626,N_21719,N_24550);
or U29627 (N_29627,N_24315,N_23651);
or U29628 (N_29628,N_22793,N_24206);
and U29629 (N_29629,N_20235,N_20663);
and U29630 (N_29630,N_24051,N_23752);
or U29631 (N_29631,N_21843,N_21854);
nor U29632 (N_29632,N_24096,N_23915);
nand U29633 (N_29633,N_22522,N_20482);
or U29634 (N_29634,N_20554,N_22359);
and U29635 (N_29635,N_23364,N_23687);
and U29636 (N_29636,N_21609,N_20409);
or U29637 (N_29637,N_24698,N_24590);
xor U29638 (N_29638,N_20878,N_23500);
and U29639 (N_29639,N_20701,N_23235);
nand U29640 (N_29640,N_21975,N_20186);
nand U29641 (N_29641,N_23678,N_22918);
and U29642 (N_29642,N_21061,N_21683);
and U29643 (N_29643,N_23733,N_21155);
nor U29644 (N_29644,N_23531,N_22401);
xnor U29645 (N_29645,N_23193,N_24913);
nor U29646 (N_29646,N_22306,N_21547);
nor U29647 (N_29647,N_24160,N_24199);
and U29648 (N_29648,N_22939,N_20462);
xnor U29649 (N_29649,N_22531,N_23342);
nor U29650 (N_29650,N_22174,N_24019);
nor U29651 (N_29651,N_22500,N_21429);
nor U29652 (N_29652,N_22425,N_22820);
and U29653 (N_29653,N_22339,N_21436);
or U29654 (N_29654,N_21146,N_22886);
nor U29655 (N_29655,N_22924,N_23214);
nor U29656 (N_29656,N_24106,N_20362);
xor U29657 (N_29657,N_22443,N_21000);
nor U29658 (N_29658,N_24379,N_24643);
and U29659 (N_29659,N_24164,N_20807);
or U29660 (N_29660,N_20054,N_22998);
nand U29661 (N_29661,N_24612,N_22096);
and U29662 (N_29662,N_22030,N_20737);
or U29663 (N_29663,N_21361,N_23886);
nand U29664 (N_29664,N_22622,N_22770);
nand U29665 (N_29665,N_24199,N_20926);
or U29666 (N_29666,N_21238,N_20094);
nor U29667 (N_29667,N_20819,N_22348);
or U29668 (N_29668,N_22892,N_21869);
nor U29669 (N_29669,N_23821,N_22646);
nor U29670 (N_29670,N_24064,N_22303);
or U29671 (N_29671,N_21860,N_20744);
nand U29672 (N_29672,N_24130,N_21057);
nand U29673 (N_29673,N_21975,N_20030);
nor U29674 (N_29674,N_20796,N_23090);
nor U29675 (N_29675,N_22291,N_23001);
xor U29676 (N_29676,N_20543,N_21529);
nand U29677 (N_29677,N_24302,N_20452);
nor U29678 (N_29678,N_24058,N_20587);
and U29679 (N_29679,N_20395,N_22735);
nor U29680 (N_29680,N_23009,N_22632);
or U29681 (N_29681,N_21226,N_23339);
and U29682 (N_29682,N_22455,N_21814);
xnor U29683 (N_29683,N_20719,N_24562);
nand U29684 (N_29684,N_20803,N_24456);
and U29685 (N_29685,N_20677,N_24520);
xnor U29686 (N_29686,N_24753,N_23739);
nand U29687 (N_29687,N_23184,N_21858);
xnor U29688 (N_29688,N_21399,N_23739);
xor U29689 (N_29689,N_22125,N_22061);
nand U29690 (N_29690,N_23696,N_24698);
xnor U29691 (N_29691,N_20253,N_23122);
or U29692 (N_29692,N_22784,N_23630);
nand U29693 (N_29693,N_20556,N_24360);
nor U29694 (N_29694,N_21977,N_21181);
or U29695 (N_29695,N_24512,N_24520);
nor U29696 (N_29696,N_21978,N_23953);
and U29697 (N_29697,N_23076,N_21096);
and U29698 (N_29698,N_22126,N_22032);
or U29699 (N_29699,N_22102,N_23849);
nand U29700 (N_29700,N_23313,N_24942);
xor U29701 (N_29701,N_21125,N_22004);
or U29702 (N_29702,N_23516,N_23220);
or U29703 (N_29703,N_23752,N_20917);
or U29704 (N_29704,N_21769,N_22713);
xor U29705 (N_29705,N_23312,N_24003);
or U29706 (N_29706,N_24849,N_23716);
or U29707 (N_29707,N_23818,N_20146);
xor U29708 (N_29708,N_23731,N_22980);
nor U29709 (N_29709,N_22478,N_23189);
or U29710 (N_29710,N_22860,N_23541);
nand U29711 (N_29711,N_20739,N_22520);
nor U29712 (N_29712,N_20682,N_23998);
nor U29713 (N_29713,N_24176,N_21600);
xnor U29714 (N_29714,N_23361,N_20374);
nor U29715 (N_29715,N_23813,N_22969);
and U29716 (N_29716,N_21493,N_22610);
and U29717 (N_29717,N_24079,N_22048);
nand U29718 (N_29718,N_22512,N_22731);
or U29719 (N_29719,N_23585,N_23260);
nor U29720 (N_29720,N_24558,N_24535);
or U29721 (N_29721,N_21292,N_21932);
xor U29722 (N_29722,N_22943,N_24931);
nand U29723 (N_29723,N_20642,N_20200);
and U29724 (N_29724,N_22943,N_23271);
xnor U29725 (N_29725,N_21342,N_20762);
xor U29726 (N_29726,N_22138,N_22440);
nand U29727 (N_29727,N_24062,N_24807);
nor U29728 (N_29728,N_20230,N_20343);
nand U29729 (N_29729,N_23280,N_24006);
and U29730 (N_29730,N_22067,N_22527);
and U29731 (N_29731,N_21550,N_21598);
nand U29732 (N_29732,N_24718,N_22754);
nand U29733 (N_29733,N_20332,N_21623);
and U29734 (N_29734,N_21905,N_22334);
xnor U29735 (N_29735,N_21993,N_21779);
nand U29736 (N_29736,N_23563,N_24345);
nor U29737 (N_29737,N_23304,N_20350);
xor U29738 (N_29738,N_24674,N_22602);
xnor U29739 (N_29739,N_24282,N_20085);
and U29740 (N_29740,N_23970,N_24818);
xor U29741 (N_29741,N_21790,N_23946);
or U29742 (N_29742,N_21876,N_24534);
or U29743 (N_29743,N_20570,N_20487);
and U29744 (N_29744,N_22992,N_20830);
and U29745 (N_29745,N_24133,N_20790);
xnor U29746 (N_29746,N_23615,N_22464);
nor U29747 (N_29747,N_24845,N_20730);
and U29748 (N_29748,N_24547,N_23964);
nor U29749 (N_29749,N_22020,N_20413);
or U29750 (N_29750,N_21412,N_24142);
or U29751 (N_29751,N_22433,N_23229);
nor U29752 (N_29752,N_20677,N_23240);
nor U29753 (N_29753,N_20773,N_22141);
xnor U29754 (N_29754,N_20456,N_21832);
xnor U29755 (N_29755,N_20946,N_21784);
and U29756 (N_29756,N_21181,N_24472);
or U29757 (N_29757,N_24265,N_22007);
nand U29758 (N_29758,N_23591,N_24165);
xor U29759 (N_29759,N_24587,N_20765);
and U29760 (N_29760,N_23793,N_24940);
and U29761 (N_29761,N_23569,N_23152);
xnor U29762 (N_29762,N_24463,N_23284);
or U29763 (N_29763,N_23937,N_22571);
and U29764 (N_29764,N_23823,N_20380);
and U29765 (N_29765,N_21853,N_21127);
nor U29766 (N_29766,N_22186,N_21751);
and U29767 (N_29767,N_20965,N_22138);
nor U29768 (N_29768,N_20087,N_24460);
nand U29769 (N_29769,N_21960,N_20411);
nand U29770 (N_29770,N_24596,N_23032);
nor U29771 (N_29771,N_21906,N_23609);
nand U29772 (N_29772,N_21037,N_22064);
and U29773 (N_29773,N_23152,N_21126);
nand U29774 (N_29774,N_23734,N_24936);
xor U29775 (N_29775,N_21513,N_21545);
or U29776 (N_29776,N_20022,N_23387);
nor U29777 (N_29777,N_21772,N_20737);
nand U29778 (N_29778,N_23509,N_23428);
xor U29779 (N_29779,N_23498,N_21664);
xnor U29780 (N_29780,N_24433,N_22503);
or U29781 (N_29781,N_20205,N_20975);
nor U29782 (N_29782,N_21414,N_23137);
and U29783 (N_29783,N_20939,N_22378);
nor U29784 (N_29784,N_20859,N_22098);
xnor U29785 (N_29785,N_22439,N_22943);
nand U29786 (N_29786,N_24260,N_22215);
nand U29787 (N_29787,N_24046,N_23894);
and U29788 (N_29788,N_24087,N_23298);
nand U29789 (N_29789,N_20678,N_24048);
nor U29790 (N_29790,N_23000,N_24643);
xor U29791 (N_29791,N_21279,N_22132);
nand U29792 (N_29792,N_22349,N_22632);
xnor U29793 (N_29793,N_21107,N_22848);
xor U29794 (N_29794,N_22592,N_24365);
nand U29795 (N_29795,N_23940,N_21920);
nand U29796 (N_29796,N_24955,N_24120);
xnor U29797 (N_29797,N_23067,N_22836);
nor U29798 (N_29798,N_24069,N_23617);
or U29799 (N_29799,N_20291,N_24057);
nand U29800 (N_29800,N_21997,N_22285);
nand U29801 (N_29801,N_24071,N_22752);
nor U29802 (N_29802,N_20993,N_20326);
nand U29803 (N_29803,N_20478,N_21716);
and U29804 (N_29804,N_22605,N_23879);
xnor U29805 (N_29805,N_20799,N_22826);
nand U29806 (N_29806,N_20580,N_22444);
and U29807 (N_29807,N_24000,N_23621);
xor U29808 (N_29808,N_24061,N_23348);
or U29809 (N_29809,N_23384,N_22498);
and U29810 (N_29810,N_20238,N_24494);
or U29811 (N_29811,N_20608,N_23793);
and U29812 (N_29812,N_23149,N_20748);
nor U29813 (N_29813,N_20190,N_24445);
nand U29814 (N_29814,N_22935,N_20915);
or U29815 (N_29815,N_20797,N_23877);
or U29816 (N_29816,N_22247,N_21587);
xnor U29817 (N_29817,N_23389,N_24648);
xor U29818 (N_29818,N_23859,N_20322);
nor U29819 (N_29819,N_21848,N_22235);
or U29820 (N_29820,N_22603,N_21070);
and U29821 (N_29821,N_21669,N_21226);
or U29822 (N_29822,N_24702,N_20863);
or U29823 (N_29823,N_22413,N_22491);
or U29824 (N_29824,N_24422,N_22327);
xor U29825 (N_29825,N_24365,N_22093);
and U29826 (N_29826,N_20304,N_23028);
or U29827 (N_29827,N_23927,N_24606);
nand U29828 (N_29828,N_24800,N_21500);
xnor U29829 (N_29829,N_23264,N_23162);
and U29830 (N_29830,N_23909,N_21693);
nor U29831 (N_29831,N_20656,N_21052);
nand U29832 (N_29832,N_22427,N_24097);
or U29833 (N_29833,N_23617,N_21551);
nand U29834 (N_29834,N_20840,N_23361);
nand U29835 (N_29835,N_23994,N_24762);
nor U29836 (N_29836,N_21809,N_23666);
nor U29837 (N_29837,N_24724,N_20867);
and U29838 (N_29838,N_21694,N_21237);
nor U29839 (N_29839,N_23785,N_20301);
xnor U29840 (N_29840,N_20811,N_22103);
nand U29841 (N_29841,N_22122,N_20843);
or U29842 (N_29842,N_23683,N_22311);
nor U29843 (N_29843,N_24859,N_23927);
or U29844 (N_29844,N_20043,N_21659);
xnor U29845 (N_29845,N_22516,N_20138);
xnor U29846 (N_29846,N_20215,N_20497);
xnor U29847 (N_29847,N_22535,N_24355);
xnor U29848 (N_29848,N_20781,N_21572);
and U29849 (N_29849,N_23565,N_21360);
and U29850 (N_29850,N_22484,N_23773);
nand U29851 (N_29851,N_22286,N_24509);
xnor U29852 (N_29852,N_24744,N_24291);
or U29853 (N_29853,N_22135,N_22517);
or U29854 (N_29854,N_23445,N_24984);
xor U29855 (N_29855,N_20575,N_22672);
nor U29856 (N_29856,N_20161,N_22433);
nand U29857 (N_29857,N_24897,N_23309);
and U29858 (N_29858,N_21108,N_24012);
nor U29859 (N_29859,N_24006,N_21402);
nand U29860 (N_29860,N_20749,N_21716);
and U29861 (N_29861,N_22531,N_24020);
and U29862 (N_29862,N_24812,N_24977);
xnor U29863 (N_29863,N_22140,N_24367);
nor U29864 (N_29864,N_20462,N_20609);
or U29865 (N_29865,N_23637,N_20076);
and U29866 (N_29866,N_21444,N_20233);
and U29867 (N_29867,N_24742,N_22959);
nand U29868 (N_29868,N_24400,N_21304);
xor U29869 (N_29869,N_20780,N_20347);
and U29870 (N_29870,N_20194,N_24645);
nand U29871 (N_29871,N_23186,N_21890);
or U29872 (N_29872,N_22297,N_21432);
nand U29873 (N_29873,N_20332,N_20909);
nor U29874 (N_29874,N_22700,N_24596);
nand U29875 (N_29875,N_21002,N_24595);
nand U29876 (N_29876,N_21190,N_24109);
nand U29877 (N_29877,N_23490,N_24269);
xor U29878 (N_29878,N_21832,N_21748);
nand U29879 (N_29879,N_24037,N_23652);
xnor U29880 (N_29880,N_21482,N_21851);
or U29881 (N_29881,N_22808,N_21206);
nand U29882 (N_29882,N_21457,N_24782);
nor U29883 (N_29883,N_24350,N_24572);
and U29884 (N_29884,N_22985,N_21469);
nor U29885 (N_29885,N_23657,N_20030);
and U29886 (N_29886,N_22914,N_20956);
xor U29887 (N_29887,N_22633,N_22127);
nand U29888 (N_29888,N_21307,N_22941);
nor U29889 (N_29889,N_21051,N_22675);
nand U29890 (N_29890,N_23280,N_20876);
nand U29891 (N_29891,N_22335,N_23890);
xor U29892 (N_29892,N_24192,N_21151);
nor U29893 (N_29893,N_23651,N_23353);
xnor U29894 (N_29894,N_22523,N_24820);
xnor U29895 (N_29895,N_22801,N_22947);
and U29896 (N_29896,N_23071,N_20264);
nor U29897 (N_29897,N_22204,N_22368);
or U29898 (N_29898,N_20099,N_21644);
xnor U29899 (N_29899,N_23474,N_24499);
nand U29900 (N_29900,N_24874,N_24217);
nand U29901 (N_29901,N_20693,N_22855);
or U29902 (N_29902,N_24628,N_23213);
nor U29903 (N_29903,N_24709,N_24675);
nand U29904 (N_29904,N_20744,N_20589);
or U29905 (N_29905,N_22464,N_23222);
xnor U29906 (N_29906,N_21525,N_23595);
xor U29907 (N_29907,N_22482,N_20616);
nand U29908 (N_29908,N_22696,N_23823);
xnor U29909 (N_29909,N_24526,N_23668);
xor U29910 (N_29910,N_22885,N_22067);
xor U29911 (N_29911,N_23645,N_20475);
nor U29912 (N_29912,N_20725,N_23938);
and U29913 (N_29913,N_20589,N_24906);
or U29914 (N_29914,N_23895,N_21324);
nor U29915 (N_29915,N_21851,N_20629);
nor U29916 (N_29916,N_21591,N_20132);
nand U29917 (N_29917,N_23212,N_23717);
and U29918 (N_29918,N_22946,N_21553);
or U29919 (N_29919,N_23218,N_23952);
xor U29920 (N_29920,N_23327,N_22360);
or U29921 (N_29921,N_24123,N_21497);
and U29922 (N_29922,N_20266,N_21066);
or U29923 (N_29923,N_20879,N_24615);
and U29924 (N_29924,N_22696,N_21508);
nor U29925 (N_29925,N_23212,N_21378);
and U29926 (N_29926,N_23953,N_23206);
nor U29927 (N_29927,N_22711,N_22577);
and U29928 (N_29928,N_21733,N_22453);
nor U29929 (N_29929,N_21862,N_24312);
or U29930 (N_29930,N_22740,N_20969);
or U29931 (N_29931,N_23007,N_20253);
or U29932 (N_29932,N_20489,N_20298);
nor U29933 (N_29933,N_21637,N_24630);
or U29934 (N_29934,N_22712,N_20812);
or U29935 (N_29935,N_20185,N_22626);
xor U29936 (N_29936,N_23584,N_21770);
and U29937 (N_29937,N_23517,N_24427);
nor U29938 (N_29938,N_20138,N_20667);
xor U29939 (N_29939,N_22274,N_21117);
and U29940 (N_29940,N_22090,N_23289);
nor U29941 (N_29941,N_21682,N_22341);
xor U29942 (N_29942,N_21147,N_23117);
and U29943 (N_29943,N_23293,N_21993);
xor U29944 (N_29944,N_23091,N_20249);
nor U29945 (N_29945,N_22762,N_20865);
nand U29946 (N_29946,N_23084,N_24539);
nor U29947 (N_29947,N_20156,N_22964);
xor U29948 (N_29948,N_22027,N_23848);
nand U29949 (N_29949,N_23968,N_20330);
nor U29950 (N_29950,N_24976,N_21421);
nand U29951 (N_29951,N_23675,N_20129);
or U29952 (N_29952,N_22347,N_24427);
xor U29953 (N_29953,N_21015,N_20578);
and U29954 (N_29954,N_22208,N_22093);
and U29955 (N_29955,N_24118,N_24184);
and U29956 (N_29956,N_21864,N_21166);
nand U29957 (N_29957,N_20900,N_21652);
xor U29958 (N_29958,N_22412,N_20021);
or U29959 (N_29959,N_23340,N_21076);
or U29960 (N_29960,N_21673,N_21725);
xor U29961 (N_29961,N_22439,N_23185);
and U29962 (N_29962,N_21620,N_22589);
nand U29963 (N_29963,N_20407,N_21376);
and U29964 (N_29964,N_24912,N_22540);
nor U29965 (N_29965,N_23481,N_21614);
and U29966 (N_29966,N_22352,N_22052);
xor U29967 (N_29967,N_21587,N_21086);
nand U29968 (N_29968,N_21877,N_23546);
and U29969 (N_29969,N_23220,N_23061);
nand U29970 (N_29970,N_24416,N_21121);
nor U29971 (N_29971,N_24516,N_24693);
xnor U29972 (N_29972,N_20838,N_20100);
xnor U29973 (N_29973,N_21220,N_24884);
and U29974 (N_29974,N_22947,N_20535);
and U29975 (N_29975,N_22910,N_21534);
nand U29976 (N_29976,N_20811,N_20494);
or U29977 (N_29977,N_24293,N_21706);
and U29978 (N_29978,N_24250,N_21516);
nand U29979 (N_29979,N_24392,N_24343);
or U29980 (N_29980,N_21924,N_21837);
or U29981 (N_29981,N_21771,N_23063);
nor U29982 (N_29982,N_23790,N_21819);
xnor U29983 (N_29983,N_23669,N_24587);
nand U29984 (N_29984,N_21921,N_20649);
and U29985 (N_29985,N_23742,N_23833);
nand U29986 (N_29986,N_20192,N_21190);
or U29987 (N_29987,N_20727,N_20000);
nand U29988 (N_29988,N_24881,N_20319);
xor U29989 (N_29989,N_21056,N_23345);
nand U29990 (N_29990,N_23501,N_23682);
or U29991 (N_29991,N_21887,N_20920);
or U29992 (N_29992,N_24775,N_22577);
nand U29993 (N_29993,N_22112,N_22324);
and U29994 (N_29994,N_21377,N_23986);
xor U29995 (N_29995,N_22726,N_23224);
and U29996 (N_29996,N_23993,N_21742);
xor U29997 (N_29997,N_21259,N_21494);
nand U29998 (N_29998,N_24547,N_23883);
xor U29999 (N_29999,N_23591,N_24675);
nand UO_0 (O_0,N_28017,N_28284);
nor UO_1 (O_1,N_29540,N_28497);
and UO_2 (O_2,N_25043,N_27188);
and UO_3 (O_3,N_26179,N_28022);
nor UO_4 (O_4,N_27133,N_27371);
nor UO_5 (O_5,N_26467,N_26295);
xnor UO_6 (O_6,N_28160,N_26563);
nor UO_7 (O_7,N_27411,N_26226);
and UO_8 (O_8,N_27159,N_27297);
nor UO_9 (O_9,N_26067,N_25700);
nand UO_10 (O_10,N_27638,N_25209);
nand UO_11 (O_11,N_26427,N_28975);
xor UO_12 (O_12,N_27030,N_27458);
and UO_13 (O_13,N_29177,N_27864);
and UO_14 (O_14,N_28104,N_29628);
xor UO_15 (O_15,N_25438,N_27464);
nand UO_16 (O_16,N_29575,N_27034);
and UO_17 (O_17,N_25070,N_28925);
xnor UO_18 (O_18,N_28416,N_28588);
and UO_19 (O_19,N_25024,N_25973);
or UO_20 (O_20,N_26748,N_28279);
and UO_21 (O_21,N_27250,N_29156);
nor UO_22 (O_22,N_29245,N_27406);
xor UO_23 (O_23,N_25900,N_29512);
nor UO_24 (O_24,N_27685,N_25513);
and UO_25 (O_25,N_29425,N_28020);
and UO_26 (O_26,N_25254,N_29279);
or UO_27 (O_27,N_26499,N_26592);
and UO_28 (O_28,N_28651,N_25224);
nor UO_29 (O_29,N_29771,N_25793);
or UO_30 (O_30,N_26309,N_29986);
and UO_31 (O_31,N_27799,N_26985);
nor UO_32 (O_32,N_25594,N_25531);
nand UO_33 (O_33,N_25415,N_26365);
xnor UO_34 (O_34,N_28737,N_28903);
and UO_35 (O_35,N_29809,N_25441);
and UO_36 (O_36,N_27665,N_25033);
nand UO_37 (O_37,N_25901,N_27395);
nor UO_38 (O_38,N_26141,N_28624);
xor UO_39 (O_39,N_26659,N_25814);
and UO_40 (O_40,N_28287,N_27619);
nand UO_41 (O_41,N_27571,N_27357);
nor UO_42 (O_42,N_26548,N_25671);
nor UO_43 (O_43,N_28200,N_29980);
nand UO_44 (O_44,N_25970,N_26180);
and UO_45 (O_45,N_27251,N_27845);
or UO_46 (O_46,N_26899,N_26550);
nand UO_47 (O_47,N_28562,N_29769);
nand UO_48 (O_48,N_29542,N_27540);
xor UO_49 (O_49,N_28335,N_29858);
nand UO_50 (O_50,N_29555,N_29496);
and UO_51 (O_51,N_25612,N_27696);
and UO_52 (O_52,N_28576,N_28509);
nor UO_53 (O_53,N_26335,N_27436);
xnor UO_54 (O_54,N_25038,N_27239);
and UO_55 (O_55,N_26975,N_25191);
xnor UO_56 (O_56,N_29972,N_25950);
or UO_57 (O_57,N_28374,N_27616);
nand UO_58 (O_58,N_27027,N_28194);
nor UO_59 (O_59,N_26241,N_27330);
and UO_60 (O_60,N_27256,N_28776);
nand UO_61 (O_61,N_28628,N_27714);
nand UO_62 (O_62,N_26122,N_25064);
nand UO_63 (O_63,N_25027,N_26643);
and UO_64 (O_64,N_27545,N_25492);
nor UO_65 (O_65,N_29011,N_26133);
and UO_66 (O_66,N_25596,N_25889);
nand UO_67 (O_67,N_27683,N_29160);
or UO_68 (O_68,N_26394,N_25683);
nor UO_69 (O_69,N_29743,N_27876);
and UO_70 (O_70,N_25204,N_27315);
nor UO_71 (O_71,N_27544,N_27935);
xor UO_72 (O_72,N_27981,N_25633);
nor UO_73 (O_73,N_27636,N_28841);
or UO_74 (O_74,N_26282,N_26436);
or UO_75 (O_75,N_29451,N_26255);
xnor UO_76 (O_76,N_26676,N_28171);
nand UO_77 (O_77,N_27702,N_29982);
or UO_78 (O_78,N_27926,N_29065);
nand UO_79 (O_79,N_28074,N_25971);
and UO_80 (O_80,N_28041,N_25420);
xor UO_81 (O_81,N_26321,N_28260);
and UO_82 (O_82,N_25959,N_25097);
xor UO_83 (O_83,N_29926,N_28470);
xnor UO_84 (O_84,N_25249,N_28960);
nor UO_85 (O_85,N_29539,N_27018);
or UO_86 (O_86,N_25831,N_26755);
and UO_87 (O_87,N_26339,N_26784);
nand UO_88 (O_88,N_29404,N_26913);
and UO_89 (O_89,N_26936,N_25346);
xor UO_90 (O_90,N_25331,N_26840);
nand UO_91 (O_91,N_28752,N_26507);
xor UO_92 (O_92,N_29917,N_28662);
nand UO_93 (O_93,N_26732,N_29170);
and UO_94 (O_94,N_26838,N_27094);
nor UO_95 (O_95,N_27692,N_25977);
and UO_96 (O_96,N_27198,N_26198);
xor UO_97 (O_97,N_29835,N_26478);
and UO_98 (O_98,N_25516,N_27867);
xor UO_99 (O_99,N_28247,N_28135);
nand UO_100 (O_100,N_25945,N_29817);
nor UO_101 (O_101,N_28859,N_29311);
xor UO_102 (O_102,N_25680,N_26614);
or UO_103 (O_103,N_29352,N_25375);
nand UO_104 (O_104,N_28229,N_29762);
xnor UO_105 (O_105,N_29370,N_27815);
nand UO_106 (O_106,N_27091,N_28610);
and UO_107 (O_107,N_25867,N_29636);
nand UO_108 (O_108,N_27412,N_26223);
xor UO_109 (O_109,N_26170,N_26422);
nor UO_110 (O_110,N_28481,N_27106);
and UO_111 (O_111,N_28542,N_26195);
or UO_112 (O_112,N_26600,N_27704);
or UO_113 (O_113,N_26235,N_26617);
nor UO_114 (O_114,N_25910,N_27587);
or UO_115 (O_115,N_25741,N_28245);
and UO_116 (O_116,N_29253,N_28832);
nor UO_117 (O_117,N_25974,N_26930);
and UO_118 (O_118,N_26519,N_28646);
and UO_119 (O_119,N_28922,N_26257);
nand UO_120 (O_120,N_25282,N_26227);
nor UO_121 (O_121,N_26421,N_25177);
or UO_122 (O_122,N_25557,N_28653);
nand UO_123 (O_123,N_29999,N_26968);
xor UO_124 (O_124,N_26542,N_29675);
and UO_125 (O_125,N_28206,N_25001);
or UO_126 (O_126,N_27490,N_29784);
nor UO_127 (O_127,N_28661,N_26286);
xor UO_128 (O_128,N_29050,N_28429);
and UO_129 (O_129,N_26809,N_29484);
nand UO_130 (O_130,N_29880,N_26729);
or UO_131 (O_131,N_26385,N_28082);
xor UO_132 (O_132,N_25462,N_29647);
and UO_133 (O_133,N_28489,N_28120);
nand UO_134 (O_134,N_28549,N_29560);
nand UO_135 (O_135,N_26698,N_27614);
xnor UO_136 (O_136,N_26770,N_29992);
or UO_137 (O_137,N_28919,N_25887);
xor UO_138 (O_138,N_27370,N_28800);
or UO_139 (O_139,N_28574,N_28359);
nor UO_140 (O_140,N_28125,N_28191);
nand UO_141 (O_141,N_26292,N_29329);
nor UO_142 (O_142,N_29318,N_26854);
nand UO_143 (O_143,N_26582,N_26711);
xnor UO_144 (O_144,N_26124,N_27923);
xor UO_145 (O_145,N_29009,N_25181);
and UO_146 (O_146,N_26147,N_27611);
nand UO_147 (O_147,N_27374,N_25560);
nor UO_148 (O_148,N_27123,N_26783);
or UO_149 (O_149,N_25032,N_29386);
xor UO_150 (O_150,N_27800,N_26443);
nand UO_151 (O_151,N_26044,N_25935);
nand UO_152 (O_152,N_28762,N_25854);
nor UO_153 (O_153,N_27884,N_25886);
nand UO_154 (O_154,N_27069,N_27017);
or UO_155 (O_155,N_29483,N_25322);
and UO_156 (O_156,N_25387,N_27722);
nor UO_157 (O_157,N_28060,N_29796);
xor UO_158 (O_158,N_25692,N_28600);
xor UO_159 (O_159,N_29744,N_27546);
or UO_160 (O_160,N_26684,N_26782);
nor UO_161 (O_161,N_28122,N_25401);
and UO_162 (O_162,N_29543,N_27946);
or UO_163 (O_163,N_28031,N_27785);
and UO_164 (O_164,N_28274,N_26864);
and UO_165 (O_165,N_26991,N_28984);
xnor UO_166 (O_166,N_26739,N_27369);
nor UO_167 (O_167,N_27512,N_25156);
nor UO_168 (O_168,N_28598,N_27667);
nor UO_169 (O_169,N_27038,N_28615);
and UO_170 (O_170,N_27456,N_25685);
nand UO_171 (O_171,N_26173,N_27718);
nor UO_172 (O_172,N_25075,N_25555);
nand UO_173 (O_173,N_25273,N_28143);
xor UO_174 (O_174,N_29124,N_28913);
nand UO_175 (O_175,N_28201,N_27589);
nand UO_176 (O_176,N_28557,N_27332);
nor UO_177 (O_177,N_27457,N_25634);
nor UO_178 (O_178,N_28044,N_28230);
xor UO_179 (O_179,N_27103,N_29938);
nand UO_180 (O_180,N_28740,N_28926);
or UO_181 (O_181,N_29854,N_27608);
and UO_182 (O_182,N_25058,N_25303);
or UO_183 (O_183,N_25501,N_26746);
or UO_184 (O_184,N_25758,N_28699);
nor UO_185 (O_185,N_25173,N_26983);
nor UO_186 (O_186,N_29394,N_26182);
nand UO_187 (O_187,N_26845,N_29067);
xnor UO_188 (O_188,N_28650,N_25522);
nand UO_189 (O_189,N_28483,N_25771);
xor UO_190 (O_190,N_25658,N_26976);
xor UO_191 (O_191,N_26967,N_26069);
nor UO_192 (O_192,N_26792,N_28631);
xor UO_193 (O_193,N_26926,N_26724);
or UO_194 (O_194,N_28000,N_27590);
nand UO_195 (O_195,N_27713,N_29228);
or UO_196 (O_196,N_26814,N_26110);
nand UO_197 (O_197,N_25246,N_29461);
and UO_198 (O_198,N_25257,N_28540);
or UO_199 (O_199,N_28132,N_26259);
nor UO_200 (O_200,N_28681,N_27009);
nor UO_201 (O_201,N_25479,N_29391);
xnor UO_202 (O_202,N_27430,N_25100);
nor UO_203 (O_203,N_26709,N_27757);
or UO_204 (O_204,N_25983,N_26607);
and UO_205 (O_205,N_27707,N_26253);
or UO_206 (O_206,N_26004,N_28121);
and UO_207 (O_207,N_29884,N_27344);
xor UO_208 (O_208,N_27929,N_26588);
or UO_209 (O_209,N_26440,N_29805);
and UO_210 (O_210,N_26603,N_28073);
xor UO_211 (O_211,N_26777,N_26974);
xor UO_212 (O_212,N_29783,N_28952);
or UO_213 (O_213,N_26671,N_28528);
xor UO_214 (O_214,N_27189,N_29166);
xor UO_215 (O_215,N_29632,N_28158);
and UO_216 (O_216,N_29446,N_25351);
xor UO_217 (O_217,N_25539,N_29673);
and UO_218 (O_218,N_27631,N_25388);
and UO_219 (O_219,N_29105,N_27081);
and UO_220 (O_220,N_28847,N_25768);
or UO_221 (O_221,N_28730,N_27193);
or UO_222 (O_222,N_25980,N_28454);
or UO_223 (O_223,N_27674,N_27759);
or UO_224 (O_224,N_28683,N_27440);
xnor UO_225 (O_225,N_25819,N_29274);
or UO_226 (O_226,N_26722,N_25708);
nand UO_227 (O_227,N_27041,N_29458);
or UO_228 (O_228,N_25563,N_25454);
and UO_229 (O_229,N_25409,N_29314);
or UO_230 (O_230,N_29471,N_28317);
nor UO_231 (O_231,N_27957,N_27036);
or UO_232 (O_232,N_28879,N_28912);
and UO_233 (O_233,N_25229,N_26336);
and UO_234 (O_234,N_28395,N_27905);
xor UO_235 (O_235,N_27663,N_26756);
and UO_236 (O_236,N_25183,N_29466);
nand UO_237 (O_237,N_27160,N_26672);
nand UO_238 (O_238,N_27329,N_28695);
nand UO_239 (O_239,N_27225,N_26345);
nand UO_240 (O_240,N_26915,N_26776);
nor UO_241 (O_241,N_26728,N_28592);
xnor UO_242 (O_242,N_26002,N_28219);
and UO_243 (O_243,N_26549,N_26095);
nor UO_244 (O_244,N_27048,N_27422);
xor UO_245 (O_245,N_28867,N_26523);
or UO_246 (O_246,N_28711,N_27124);
or UO_247 (O_247,N_26795,N_29725);
xor UO_248 (O_248,N_26463,N_28364);
and UO_249 (O_249,N_25448,N_26202);
and UO_250 (O_250,N_25558,N_25028);
nand UO_251 (O_251,N_28726,N_25337);
xnor UO_252 (O_252,N_28788,N_26639);
nand UO_253 (O_253,N_29635,N_26948);
nor UO_254 (O_254,N_25523,N_25366);
or UO_255 (O_255,N_29094,N_28927);
and UO_256 (O_256,N_25996,N_28619);
nand UO_257 (O_257,N_29117,N_29367);
nor UO_258 (O_258,N_25083,N_29006);
nand UO_259 (O_259,N_27824,N_27285);
nand UO_260 (O_260,N_26708,N_26094);
xnor UO_261 (O_261,N_25564,N_26921);
or UO_262 (O_262,N_29293,N_25789);
xnor UO_263 (O_263,N_25638,N_27801);
and UO_264 (O_264,N_29180,N_25731);
xor UO_265 (O_265,N_29022,N_27355);
xnor UO_266 (O_266,N_29178,N_26396);
nand UO_267 (O_267,N_28732,N_28485);
and UO_268 (O_268,N_25088,N_29222);
and UO_269 (O_269,N_26749,N_27296);
nor UO_270 (O_270,N_28543,N_27210);
and UO_271 (O_271,N_28423,N_27382);
nor UO_272 (O_272,N_25650,N_28962);
and UO_273 (O_273,N_28982,N_26049);
nor UO_274 (O_274,N_26754,N_27971);
xnor UO_275 (O_275,N_27673,N_27945);
nor UO_276 (O_276,N_27183,N_29856);
and UO_277 (O_277,N_29573,N_25614);
xor UO_278 (O_278,N_28321,N_29075);
and UO_279 (O_279,N_27287,N_26406);
or UO_280 (O_280,N_28316,N_25251);
and UO_281 (O_281,N_27200,N_25013);
and UO_282 (O_282,N_27213,N_28837);
xor UO_283 (O_283,N_25002,N_27699);
and UO_284 (O_284,N_29915,N_28564);
or UO_285 (O_285,N_27166,N_25000);
nor UO_286 (O_286,N_25404,N_25572);
xor UO_287 (O_287,N_29307,N_27120);
nor UO_288 (O_288,N_28467,N_25076);
xor UO_289 (O_289,N_28178,N_29076);
and UO_290 (O_290,N_29593,N_26896);
or UO_291 (O_291,N_27465,N_25110);
and UO_292 (O_292,N_27359,N_27377);
and UO_293 (O_293,N_26943,N_27862);
nor UO_294 (O_294,N_25292,N_28917);
or UO_295 (O_295,N_27071,N_29128);
xnor UO_296 (O_296,N_26237,N_28996);
or UO_297 (O_297,N_28731,N_25504);
nand UO_298 (O_298,N_26876,N_27341);
and UO_299 (O_299,N_28633,N_29997);
nand UO_300 (O_300,N_25528,N_27844);
nand UO_301 (O_301,N_26250,N_26284);
xnor UO_302 (O_302,N_28197,N_27909);
xor UO_303 (O_303,N_25035,N_27684);
or UO_304 (O_304,N_28319,N_29069);
nor UO_305 (O_305,N_26111,N_28884);
nor UO_306 (O_306,N_26283,N_28465);
nand UO_307 (O_307,N_26252,N_26839);
nand UO_308 (O_308,N_29860,N_27102);
xnor UO_309 (O_309,N_27519,N_28340);
nor UO_310 (O_310,N_29712,N_27079);
or UO_311 (O_311,N_27230,N_27536);
or UO_312 (O_312,N_28812,N_28008);
nand UO_313 (O_313,N_28290,N_25606);
or UO_314 (O_314,N_27218,N_29697);
xor UO_315 (O_315,N_26668,N_27990);
nor UO_316 (O_316,N_29190,N_28707);
and UO_317 (O_317,N_25858,N_27237);
and UO_318 (O_318,N_29153,N_28873);
xnor UO_319 (O_319,N_29879,N_25837);
xnor UO_320 (O_320,N_26702,N_26922);
nor UO_321 (O_321,N_27535,N_26054);
nor UO_322 (O_322,N_26298,N_29183);
and UO_323 (O_323,N_29135,N_29761);
nor UO_324 (O_324,N_29102,N_29015);
nor UO_325 (O_325,N_27021,N_27754);
or UO_326 (O_326,N_28590,N_29832);
nor UO_327 (O_327,N_25948,N_26105);
xor UO_328 (O_328,N_25221,N_26885);
nor UO_329 (O_329,N_29481,N_25020);
and UO_330 (O_330,N_27158,N_29270);
and UO_331 (O_331,N_29513,N_29137);
and UO_332 (O_332,N_25139,N_28669);
xnor UO_333 (O_333,N_27523,N_29152);
nand UO_334 (O_334,N_26473,N_29621);
or UO_335 (O_335,N_27090,N_25905);
or UO_336 (O_336,N_28932,N_29230);
or UO_337 (O_337,N_27117,N_29336);
nand UO_338 (O_338,N_25413,N_26058);
or UO_339 (O_339,N_29072,N_26697);
nor UO_340 (O_340,N_29189,N_26305);
and UO_341 (O_341,N_27324,N_25823);
nor UO_342 (O_342,N_27394,N_29295);
nand UO_343 (O_343,N_28415,N_27605);
nand UO_344 (O_344,N_26497,N_27122);
nor UO_345 (O_345,N_29871,N_27861);
xor UO_346 (O_346,N_28571,N_26190);
nand UO_347 (O_347,N_28016,N_29384);
nor UO_348 (O_348,N_28830,N_28510);
or UO_349 (O_349,N_26844,N_28724);
and UO_350 (O_350,N_28626,N_25506);
nand UO_351 (O_351,N_26664,N_28751);
xnor UO_352 (O_352,N_25654,N_26175);
nor UO_353 (O_353,N_25082,N_28258);
and UO_354 (O_354,N_25389,N_26780);
nor UO_355 (O_355,N_25707,N_29099);
nand UO_356 (O_356,N_25616,N_26013);
nand UO_357 (O_357,N_28254,N_28898);
xnor UO_358 (O_358,N_26912,N_29694);
and UO_359 (O_359,N_27064,N_27109);
nand UO_360 (O_360,N_29289,N_25095);
nand UO_361 (O_361,N_25086,N_26458);
nor UO_362 (O_362,N_28768,N_27461);
nor UO_363 (O_363,N_25993,N_29488);
nor UO_364 (O_364,N_29755,N_27810);
nor UO_365 (O_365,N_29885,N_27248);
or UO_366 (O_366,N_25185,N_25481);
nand UO_367 (O_367,N_27553,N_25094);
nor UO_368 (O_368,N_27023,N_28114);
nand UO_369 (O_369,N_28580,N_26815);
and UO_370 (O_370,N_25987,N_28582);
or UO_371 (O_371,N_26152,N_26666);
and UO_372 (O_372,N_29339,N_27860);
xnor UO_373 (O_373,N_27467,N_25336);
nand UO_374 (O_374,N_26859,N_27451);
and UO_375 (O_375,N_29833,N_26744);
nor UO_376 (O_376,N_29998,N_25137);
and UO_377 (O_377,N_29603,N_27579);
xor UO_378 (O_378,N_25717,N_29489);
xnor UO_379 (O_379,N_29702,N_27555);
xor UO_380 (O_380,N_29836,N_27520);
or UO_381 (O_381,N_28746,N_28381);
or UO_382 (O_382,N_25126,N_26893);
nand UO_383 (O_383,N_28920,N_27984);
nor UO_384 (O_384,N_27044,N_28591);
and UO_385 (O_385,N_28660,N_29087);
xor UO_386 (O_386,N_28209,N_29609);
xnor UO_387 (O_387,N_28559,N_25856);
or UO_388 (O_388,N_29179,N_27675);
and UO_389 (O_389,N_28261,N_28622);
nor UO_390 (O_390,N_27443,N_29114);
and UO_391 (O_391,N_27477,N_25140);
and UO_392 (O_392,N_25681,N_25686);
nor UO_393 (O_393,N_25532,N_29366);
xor UO_394 (O_394,N_28028,N_25678);
nor UO_395 (O_395,N_28231,N_29460);
xnor UO_396 (O_396,N_29017,N_29748);
nor UO_397 (O_397,N_26430,N_29759);
and UO_398 (O_398,N_28336,N_29775);
nor UO_399 (O_399,N_26829,N_25483);
nor UO_400 (O_400,N_25966,N_28313);
nand UO_401 (O_401,N_25418,N_28393);
nand UO_402 (O_402,N_29400,N_28346);
nand UO_403 (O_403,N_27226,N_27319);
and UO_404 (O_404,N_27100,N_27776);
xor UO_405 (O_405,N_29732,N_26349);
nor UO_406 (O_406,N_26313,N_28307);
nor UO_407 (O_407,N_27110,N_28506);
nor UO_408 (O_408,N_28648,N_27507);
and UO_409 (O_409,N_27276,N_29368);
nand UO_410 (O_410,N_29263,N_25272);
nand UO_411 (O_411,N_28754,N_29150);
xor UO_412 (O_412,N_25426,N_27541);
nand UO_413 (O_413,N_26945,N_27660);
xnor UO_414 (O_414,N_26263,N_28502);
and UO_415 (O_415,N_25396,N_29000);
and UO_416 (O_416,N_27425,N_27356);
nand UO_417 (O_417,N_26794,N_27392);
xor UO_418 (O_418,N_27872,N_26387);
nor UO_419 (O_419,N_29202,N_29996);
nand UO_420 (O_420,N_28348,N_27416);
or UO_421 (O_421,N_26219,N_26453);
and UO_422 (O_422,N_25120,N_29966);
or UO_423 (O_423,N_29729,N_26460);
xor UO_424 (O_424,N_25308,N_25601);
xnor UO_425 (O_425,N_25761,N_29045);
or UO_426 (O_426,N_27615,N_29514);
or UO_427 (O_427,N_25157,N_27847);
nand UO_428 (O_428,N_27994,N_29953);
nand UO_429 (O_429,N_29167,N_25382);
nand UO_430 (O_430,N_27770,N_28672);
nand UO_431 (O_431,N_27354,N_29613);
and UO_432 (O_432,N_25459,N_26793);
xor UO_433 (O_433,N_29172,N_27893);
nand UO_434 (O_434,N_29049,N_27664);
xnor UO_435 (O_435,N_27538,N_25194);
or UO_436 (O_436,N_29850,N_27951);
nand UO_437 (O_437,N_27145,N_29639);
nor UO_438 (O_438,N_25862,N_29902);
nor UO_439 (O_439,N_26447,N_27715);
xnor UO_440 (O_440,N_26304,N_29056);
xor UO_441 (O_441,N_28055,N_27516);
xnor UO_442 (O_442,N_25115,N_25988);
nand UO_443 (O_443,N_27635,N_26125);
or UO_444 (O_444,N_25381,N_27599);
xor UO_445 (O_445,N_28164,N_26966);
xor UO_446 (O_446,N_27428,N_28471);
nor UO_447 (O_447,N_28086,N_28198);
nor UO_448 (O_448,N_26932,N_28593);
nand UO_449 (O_449,N_27679,N_26493);
xnor UO_450 (O_450,N_25453,N_29301);
and UO_451 (O_451,N_25992,N_26620);
xnor UO_452 (O_452,N_25424,N_28302);
and UO_453 (O_453,N_27934,N_27574);
xor UO_454 (O_454,N_25690,N_28161);
xor UO_455 (O_455,N_27559,N_27093);
xnor UO_456 (O_456,N_26310,N_27916);
xor UO_457 (O_457,N_26351,N_27940);
or UO_458 (O_458,N_28192,N_27077);
and UO_459 (O_459,N_29249,N_29242);
nand UO_460 (O_460,N_25764,N_29822);
xor UO_461 (O_461,N_26665,N_27281);
and UO_462 (O_462,N_29186,N_29260);
nor UO_463 (O_463,N_25072,N_25384);
or UO_464 (O_464,N_27409,N_26027);
and UO_465 (O_465,N_29674,N_26738);
and UO_466 (O_466,N_28692,N_26516);
xnor UO_467 (O_467,N_26290,N_29756);
xor UO_468 (O_468,N_26873,N_26890);
and UO_469 (O_469,N_25664,N_25329);
nor UO_470 (O_470,N_26568,N_28741);
nand UO_471 (O_471,N_27868,N_25933);
nand UO_472 (O_472,N_27504,N_27502);
xnor UO_473 (O_473,N_25160,N_28948);
nor UO_474 (O_474,N_29062,N_28461);
and UO_475 (O_475,N_28882,N_29371);
xor UO_476 (O_476,N_25928,N_28756);
nor UO_477 (O_477,N_26959,N_29215);
nor UO_478 (O_478,N_25326,N_26834);
xor UO_479 (O_479,N_25878,N_26374);
xnor UO_480 (O_480,N_25573,N_26802);
and UO_481 (O_481,N_25188,N_27883);
xor UO_482 (O_482,N_28684,N_26047);
xor UO_483 (O_483,N_28487,N_25269);
nand UO_484 (O_484,N_27136,N_27184);
nand UO_485 (O_485,N_25958,N_25080);
and UO_486 (O_486,N_26598,N_28456);
xnor UO_487 (O_487,N_29054,N_26832);
or UO_488 (O_488,N_26522,N_25569);
nor UO_489 (O_489,N_28596,N_27505);
and UO_490 (O_490,N_26630,N_29309);
nor UO_491 (O_491,N_29994,N_29584);
nand UO_492 (O_492,N_27643,N_27780);
or UO_493 (O_493,N_26515,N_26944);
and UO_494 (O_494,N_29332,N_25848);
or UO_495 (O_495,N_25073,N_26660);
nand UO_496 (O_496,N_26995,N_28366);
nand UO_497 (O_497,N_28150,N_26841);
nor UO_498 (O_498,N_27235,N_29291);
and UO_499 (O_499,N_27343,N_29343);
xnor UO_500 (O_500,N_25317,N_28545);
xor UO_501 (O_501,N_25212,N_29046);
nor UO_502 (O_502,N_25648,N_29456);
or UO_503 (O_503,N_27711,N_29088);
or UO_504 (O_504,N_27180,N_27806);
xor UO_505 (O_505,N_26622,N_25914);
nand UO_506 (O_506,N_27208,N_28805);
xor UO_507 (O_507,N_28180,N_28070);
nor UO_508 (O_508,N_26129,N_26391);
or UO_509 (O_509,N_28743,N_29767);
nor UO_510 (O_510,N_26655,N_29115);
nand UO_511 (O_511,N_25061,N_29376);
nand UO_512 (O_512,N_28609,N_25402);
xor UO_513 (O_513,N_29718,N_25197);
or UO_514 (O_514,N_26540,N_25223);
nor UO_515 (O_515,N_26470,N_29604);
nor UO_516 (O_516,N_28281,N_25148);
nor UO_517 (O_517,N_27263,N_27853);
nand UO_518 (O_518,N_29845,N_28351);
or UO_519 (O_519,N_28492,N_27890);
or UO_520 (O_520,N_28839,N_29701);
nand UO_521 (O_521,N_27275,N_28136);
or UO_522 (O_522,N_28778,N_25801);
or UO_523 (O_523,N_26725,N_25053);
nand UO_524 (O_524,N_26176,N_29933);
nand UO_525 (O_525,N_29793,N_26418);
and UO_526 (O_526,N_27266,N_25979);
xor UO_527 (O_527,N_26765,N_28371);
nor UO_528 (O_528,N_29853,N_25476);
and UO_529 (O_529,N_25796,N_29408);
and UO_530 (O_530,N_28782,N_26092);
xnor UO_531 (O_531,N_28248,N_28077);
and UO_532 (O_532,N_25877,N_25691);
or UO_533 (O_533,N_25328,N_25025);
nor UO_534 (O_534,N_25968,N_26713);
nand UO_535 (O_535,N_25163,N_27518);
nand UO_536 (O_536,N_25849,N_25376);
xor UO_537 (O_537,N_27846,N_27837);
and UO_538 (O_538,N_26957,N_27529);
and UO_539 (O_539,N_29134,N_29390);
nand UO_540 (O_540,N_28029,N_27289);
nand UO_541 (O_541,N_26040,N_28872);
xnor UO_542 (O_542,N_26505,N_26136);
or UO_543 (O_543,N_27243,N_28417);
and UO_544 (O_544,N_26730,N_28515);
xor UO_545 (O_545,N_27424,N_26014);
or UO_546 (O_546,N_29350,N_27626);
xor UO_547 (O_547,N_26449,N_27695);
xnor UO_548 (O_548,N_28498,N_27784);
xor UO_549 (O_549,N_27282,N_26327);
and UO_550 (O_550,N_25490,N_27294);
nor UO_551 (O_551,N_27569,N_26140);
or UO_552 (O_552,N_25833,N_29106);
and UO_553 (O_553,N_29717,N_28685);
xor UO_554 (O_554,N_26760,N_25365);
or UO_555 (O_555,N_26862,N_26016);
nor UO_556 (O_556,N_26685,N_29735);
or UO_557 (O_557,N_28057,N_28155);
xor UO_558 (O_558,N_25180,N_25561);
nand UO_559 (O_559,N_25631,N_28457);
or UO_560 (O_560,N_27125,N_29248);
or UO_561 (O_561,N_29764,N_25443);
or UO_562 (O_562,N_29437,N_29438);
nor UO_563 (O_563,N_29219,N_28146);
and UO_564 (O_564,N_25472,N_25884);
nor UO_565 (O_565,N_26168,N_28232);
and UO_566 (O_566,N_25762,N_26101);
or UO_567 (O_567,N_27524,N_28541);
or UO_568 (O_568,N_27610,N_28108);
and UO_569 (O_569,N_27305,N_26400);
nand UO_570 (O_570,N_25362,N_25334);
xnor UO_571 (O_571,N_28376,N_28696);
and UO_572 (O_572,N_26775,N_26414);
and UO_573 (O_573,N_25068,N_29497);
nor UO_574 (O_574,N_25545,N_25917);
nand UO_575 (O_575,N_26196,N_28403);
xor UO_576 (O_576,N_26192,N_27609);
and UO_577 (O_577,N_29205,N_25279);
nand UO_578 (O_578,N_29261,N_25739);
nor UO_579 (O_579,N_26098,N_25444);
nand UO_580 (O_580,N_27222,N_27493);
or UO_581 (O_581,N_28005,N_26874);
xnor UO_582 (O_582,N_26552,N_26112);
xnor UO_583 (O_583,N_28611,N_27140);
nand UO_584 (O_584,N_26380,N_27337);
nand UO_585 (O_585,N_25635,N_26590);
or UO_586 (O_586,N_25391,N_26599);
nand UO_587 (O_587,N_26267,N_29554);
or UO_588 (O_588,N_25986,N_29873);
or UO_589 (O_589,N_28329,N_25360);
and UO_590 (O_590,N_28480,N_26560);
nand UO_591 (O_591,N_25668,N_25162);
and UO_592 (O_592,N_27922,N_26997);
xor UO_593 (O_593,N_25855,N_26787);
or UO_594 (O_594,N_26682,N_27037);
xnor UO_595 (O_595,N_25009,N_26687);
or UO_596 (O_596,N_26177,N_25985);
and UO_597 (O_597,N_29428,N_28068);
or UO_598 (O_598,N_29815,N_27568);
and UO_599 (O_599,N_25335,N_25345);
nor UO_600 (O_600,N_26998,N_28654);
or UO_601 (O_601,N_27086,N_29654);
and UO_602 (O_602,N_29785,N_28392);
nand UO_603 (O_603,N_25751,N_28799);
or UO_604 (O_604,N_25795,N_26085);
nand UO_605 (O_605,N_29546,N_29276);
nor UO_606 (O_606,N_25484,N_28115);
nor UO_607 (O_607,N_25283,N_29830);
xor UO_608 (O_608,N_26881,N_27501);
xor UO_609 (O_609,N_29766,N_26018);
or UO_610 (O_610,N_27948,N_29631);
nor UO_611 (O_611,N_29977,N_28914);
xnor UO_612 (O_612,N_29173,N_27818);
xnor UO_613 (O_613,N_25008,N_29557);
nand UO_614 (O_614,N_26486,N_27814);
nor UO_615 (O_615,N_26119,N_25955);
nor UO_616 (O_616,N_29900,N_28061);
xnor UO_617 (O_617,N_26642,N_25466);
nand UO_618 (O_618,N_25258,N_26416);
nand UO_619 (O_619,N_28761,N_27530);
and UO_620 (O_620,N_27383,N_27085);
xor UO_621 (O_621,N_27959,N_29220);
xnor UO_622 (O_622,N_26823,N_25482);
nor UO_623 (O_623,N_28964,N_27972);
nand UO_624 (O_624,N_25294,N_26594);
nor UO_625 (O_625,N_28406,N_27481);
nand UO_626 (O_626,N_26323,N_29440);
nor UO_627 (O_627,N_25442,N_26376);
nor UO_628 (O_628,N_28512,N_25982);
or UO_629 (O_629,N_29116,N_29185);
or UO_630 (O_630,N_26626,N_26821);
or UO_631 (O_631,N_28658,N_27469);
nor UO_632 (O_632,N_28735,N_29216);
or UO_633 (O_633,N_27521,N_25244);
nand UO_634 (O_634,N_27393,N_25323);
nand UO_635 (O_635,N_26469,N_26662);
nand UO_636 (O_636,N_29950,N_28360);
nand UO_637 (O_637,N_27431,N_26410);
nor UO_638 (O_638,N_29812,N_29672);
and UO_639 (O_639,N_28630,N_29284);
nor UO_640 (O_640,N_29763,N_27185);
nor UO_641 (O_641,N_25480,N_29235);
xnor UO_642 (O_642,N_28802,N_26187);
nand UO_643 (O_643,N_29027,N_28099);
or UO_644 (O_644,N_29585,N_29282);
and UO_645 (O_645,N_27491,N_26311);
nor UO_646 (O_646,N_26317,N_25550);
or UO_647 (O_647,N_26940,N_25217);
and UO_648 (O_648,N_25458,N_29798);
and UO_649 (O_649,N_25791,N_26456);
xor UO_650 (O_650,N_27967,N_27762);
xnor UO_651 (O_651,N_27999,N_27895);
xor UO_652 (O_652,N_28306,N_27376);
nand UO_653 (O_653,N_25581,N_26958);
nor UO_654 (O_654,N_29740,N_29907);
and UO_655 (O_655,N_29503,N_27249);
nand UO_656 (O_656,N_27207,N_26273);
xnor UO_657 (O_657,N_27921,N_25364);
and UO_658 (O_658,N_26867,N_26907);
or UO_659 (O_659,N_29224,N_28856);
nor UO_660 (O_660,N_25805,N_29129);
or UO_661 (O_661,N_25417,N_29989);
or UO_662 (O_662,N_25296,N_27639);
nor UO_663 (O_663,N_27691,N_27385);
and UO_664 (O_664,N_28869,N_25135);
and UO_665 (O_665,N_27775,N_29958);
and UO_666 (O_666,N_26271,N_29144);
or UO_667 (O_667,N_26157,N_28438);
or UO_668 (O_668,N_26565,N_27258);
nand UO_669 (O_669,N_28401,N_28204);
nor UO_670 (O_670,N_28310,N_28218);
or UO_671 (O_671,N_25892,N_27052);
and UO_672 (O_672,N_29158,N_29644);
and UO_673 (O_673,N_27840,N_29341);
or UO_674 (O_674,N_25722,N_25339);
nor UO_675 (O_675,N_25994,N_25285);
xnor UO_676 (O_676,N_29952,N_28824);
and UO_677 (O_677,N_27557,N_29623);
xor UO_678 (O_678,N_25565,N_25562);
or UO_679 (O_679,N_28995,N_28988);
xor UO_680 (O_680,N_26099,N_26360);
and UO_681 (O_681,N_28827,N_26889);
nand UO_682 (O_682,N_25719,N_29565);
xnor UO_683 (O_683,N_26035,N_27484);
nand UO_684 (O_684,N_26143,N_25641);
nand UO_685 (O_685,N_27548,N_26358);
nand UO_686 (O_686,N_28468,N_28526);
nor UO_687 (O_687,N_27658,N_25216);
and UO_688 (O_688,N_26379,N_25997);
and UO_689 (O_689,N_26091,N_26167);
nand UO_690 (O_690,N_26640,N_27358);
and UO_691 (O_691,N_28686,N_27672);
and UO_692 (O_692,N_28049,N_27311);
and UO_693 (O_693,N_25976,N_29522);
nand UO_694 (O_694,N_26189,N_29002);
and UO_695 (O_695,N_26835,N_25399);
nand UO_696 (O_696,N_29090,N_25010);
xnor UO_697 (O_697,N_26397,N_25777);
or UO_698 (O_698,N_25757,N_26883);
nand UO_699 (O_699,N_29930,N_26901);
xnor UO_700 (O_700,N_28064,N_25250);
xnor UO_701 (O_701,N_28240,N_29161);
or UO_702 (O_702,N_28341,N_29434);
and UO_703 (O_703,N_25348,N_27751);
or UO_704 (O_704,N_25822,N_26923);
xnor UO_705 (O_705,N_25069,N_25559);
nor UO_706 (O_706,N_27384,N_26481);
nand UO_707 (O_707,N_27932,N_28142);
nor UO_708 (O_708,N_26804,N_28129);
xnor UO_709 (O_709,N_26584,N_29423);
xor UO_710 (O_710,N_25821,N_28162);
or UO_711 (O_711,N_29445,N_26624);
and UO_712 (O_712,N_28156,N_27816);
or UO_713 (O_713,N_26570,N_26046);
and UO_714 (O_714,N_26183,N_27901);
and UO_715 (O_715,N_25187,N_28195);
nand UO_716 (O_716,N_27462,N_25546);
and UO_717 (O_717,N_25609,N_27402);
or UO_718 (O_718,N_28644,N_29032);
nor UO_719 (O_719,N_28620,N_28807);
nor UO_720 (O_720,N_28058,N_28929);
xnor UO_721 (O_721,N_28076,N_29646);
xnor UO_722 (O_722,N_29578,N_26372);
or UO_723 (O_723,N_26382,N_28518);
and UO_724 (O_724,N_25597,N_26268);
or UO_725 (O_725,N_25679,N_29058);
and UO_726 (O_726,N_25727,N_26240);
nand UO_727 (O_727,N_27471,N_25149);
xor UO_728 (O_728,N_26266,N_29713);
nor UO_729 (O_729,N_27592,N_26020);
and UO_730 (O_730,N_25781,N_26482);
and UO_731 (O_731,N_29174,N_29469);
nor UO_732 (O_732,N_27224,N_29048);
nor UO_733 (O_733,N_29828,N_27760);
xnor UO_734 (O_734,N_29078,N_26079);
xor UO_735 (O_735,N_29956,N_27204);
or UO_736 (O_736,N_28389,N_28780);
and UO_737 (O_737,N_28634,N_26865);
nor UO_738 (O_738,N_25904,N_27177);
or UO_739 (O_739,N_27703,N_26393);
and UO_740 (O_740,N_25102,N_28004);
nand UO_741 (O_741,N_27716,N_25926);
nand UO_742 (O_742,N_28353,N_26296);
nand UO_743 (O_743,N_25699,N_28728);
and UO_744 (O_744,N_25603,N_27264);
nand UO_745 (O_745,N_28069,N_28792);
and UO_746 (O_746,N_27496,N_25753);
xor UO_747 (O_747,N_27552,N_26123);
xnor UO_748 (O_748,N_25760,N_29491);
nand UO_749 (O_749,N_28038,N_27657);
xor UO_750 (O_750,N_26597,N_27363);
and UO_751 (O_751,N_25245,N_26354);
and UO_752 (O_752,N_26619,N_28930);
nor UO_753 (O_753,N_27391,N_27678);
nand UO_754 (O_754,N_26205,N_27653);
xnor UO_755 (O_755,N_29657,N_28876);
nor UO_756 (O_756,N_25651,N_25219);
nand UO_757 (O_757,N_25624,N_29285);
or UO_758 (O_758,N_29409,N_25919);
and UO_759 (O_759,N_29728,N_25499);
xor UO_760 (O_760,N_25592,N_29250);
or UO_761 (O_761,N_27365,N_25735);
xnor UO_762 (O_762,N_28689,N_29937);
nor UO_763 (O_763,N_27809,N_27730);
or UO_764 (O_764,N_27708,N_29551);
or UO_765 (O_765,N_26343,N_26377);
and UO_766 (O_766,N_29501,N_25261);
or UO_767 (O_767,N_25780,N_29820);
nand UO_768 (O_768,N_25059,N_27455);
and UO_769 (O_769,N_27510,N_25215);
or UO_770 (O_770,N_25742,N_26531);
or UO_771 (O_771,N_26539,N_27234);
nor UO_772 (O_772,N_25723,N_28533);
and UO_773 (O_773,N_26138,N_28106);
or UO_774 (O_774,N_28174,N_25938);
or UO_775 (O_775,N_29226,N_29875);
xnor UO_776 (O_776,N_29210,N_29943);
or UO_777 (O_777,N_28719,N_26952);
nor UO_778 (O_778,N_25920,N_28271);
or UO_779 (O_779,N_27483,N_28535);
nor UO_780 (O_780,N_26333,N_27791);
nor UO_781 (O_781,N_26852,N_26217);
nand UO_782 (O_782,N_25371,N_25653);
or UO_783 (O_783,N_29424,N_25524);
nor UO_784 (O_784,N_26464,N_26256);
nor UO_785 (O_785,N_28822,N_25607);
and UO_786 (O_786,N_25514,N_27335);
xor UO_787 (O_787,N_29749,N_25433);
xnor UO_788 (O_788,N_25370,N_26494);
nand UO_789 (O_789,N_26949,N_26737);
xor UO_790 (O_790,N_26750,N_27680);
xor UO_791 (O_791,N_27745,N_28203);
nand UO_792 (O_792,N_27452,N_29092);
nor UO_793 (O_793,N_26090,N_26314);
or UO_794 (O_794,N_25610,N_25645);
and UO_795 (O_795,N_25128,N_27441);
nand UO_796 (O_796,N_27020,N_29541);
nor UO_797 (O_797,N_27897,N_26225);
nand UO_798 (O_798,N_26148,N_29719);
nand UO_799 (O_799,N_27700,N_27303);
nand UO_800 (O_800,N_27503,N_26524);
nand UO_801 (O_801,N_29599,N_25618);
and UO_802 (O_802,N_29891,N_29450);
or UO_803 (O_803,N_29316,N_28291);
or UO_804 (O_804,N_25736,N_25918);
xnor UO_805 (O_805,N_28575,N_28257);
or UO_806 (O_806,N_27634,N_26608);
nand UO_807 (O_807,N_27126,N_28112);
or UO_808 (O_808,N_26355,N_28586);
xor UO_809 (O_809,N_26887,N_29187);
or UO_810 (O_810,N_27931,N_25497);
or UO_811 (O_811,N_28954,N_27811);
or UO_812 (O_812,N_29797,N_25022);
nor UO_813 (O_813,N_26796,N_26228);
and UO_814 (O_814,N_26006,N_28478);
nor UO_815 (O_815,N_29310,N_27202);
nor UO_816 (O_816,N_25023,N_29876);
xor UO_817 (O_817,N_26121,N_26249);
nor UO_818 (O_818,N_29004,N_28091);
xor UO_819 (O_819,N_26925,N_28870);
or UO_820 (O_820,N_25324,N_25655);
xnor UO_821 (O_821,N_25556,N_25876);
nor UO_822 (O_822,N_28815,N_25014);
and UO_823 (O_823,N_26723,N_29942);
nand UO_824 (O_824,N_25309,N_28331);
xor UO_825 (O_825,N_29165,N_29754);
or UO_826 (O_826,N_28296,N_25380);
xnor UO_827 (O_827,N_28665,N_25451);
and UO_828 (O_828,N_26653,N_29120);
nand UO_829 (O_829,N_28133,N_27556);
nand UO_830 (O_830,N_29277,N_25657);
or UO_831 (O_831,N_27259,N_25827);
or UO_832 (O_832,N_26116,N_29143);
or UO_833 (O_833,N_27152,N_29670);
and UO_834 (O_834,N_26291,N_25705);
and UO_835 (O_835,N_29969,N_25505);
or UO_836 (O_836,N_28264,N_25575);
xnor UO_837 (O_837,N_26810,N_27401);
and UO_838 (O_838,N_25325,N_25225);
nor UO_839 (O_839,N_25912,N_26510);
nor UO_840 (O_840,N_28779,N_29119);
nor UO_841 (O_841,N_26233,N_26017);
and UO_842 (O_842,N_28220,N_27654);
or UO_843 (O_843,N_29864,N_27581);
nor UO_844 (O_844,N_25766,N_29727);
nand UO_845 (O_845,N_27982,N_25542);
nand UO_846 (O_846,N_29467,N_28972);
or UO_847 (O_847,N_25520,N_28190);
nor UO_848 (O_848,N_25407,N_27835);
or UO_849 (O_849,N_27220,N_28517);
or UO_850 (O_850,N_28736,N_26025);
and UO_851 (O_851,N_29903,N_25600);
nor UO_852 (O_852,N_25344,N_27310);
nand UO_853 (O_853,N_26052,N_26477);
nand UO_854 (O_854,N_25447,N_27301);
and UO_855 (O_855,N_29305,N_26371);
and UO_856 (O_856,N_25290,N_27676);
nor UO_857 (O_857,N_28697,N_29831);
nor UO_858 (O_858,N_27352,N_28556);
xor UO_859 (O_859,N_27686,N_28552);
xor UO_860 (O_860,N_29711,N_26924);
nand UO_861 (O_861,N_28581,N_25171);
or UO_862 (O_862,N_29855,N_25271);
nand UO_863 (O_863,N_26483,N_28771);
xnor UO_864 (O_864,N_29530,N_28983);
and UO_865 (O_865,N_28516,N_26155);
or UO_866 (O_866,N_27888,N_26281);
and UO_867 (O_867,N_29387,N_26606);
nor UO_868 (O_868,N_28418,N_29233);
nor UO_869 (O_869,N_28645,N_25019);
and UO_870 (O_870,N_28705,N_29237);
nand UO_871 (O_871,N_26086,N_28035);
xor UO_872 (O_872,N_27221,N_29147);
and UO_873 (O_873,N_27063,N_25167);
xor UO_874 (O_874,N_29605,N_26325);
nor UO_875 (O_875,N_25763,N_29923);
or UO_876 (O_876,N_26057,N_25989);
nand UO_877 (O_877,N_27973,N_27542);
nor UO_878 (O_878,N_26294,N_27163);
nor UO_879 (O_879,N_28318,N_25737);
nor UO_880 (O_880,N_25253,N_29095);
or UO_881 (O_881,N_29296,N_25755);
or UO_882 (O_882,N_27706,N_29133);
nand UO_883 (O_883,N_25270,N_28391);
nand UO_884 (O_884,N_27293,N_26933);
or UO_885 (O_885,N_25908,N_29535);
xor UO_886 (O_886,N_28090,N_27309);
xor UO_887 (O_887,N_29693,N_28817);
or UO_888 (O_888,N_28409,N_25353);
nor UO_889 (O_889,N_26126,N_26605);
nor UO_890 (O_890,N_25773,N_27029);
nand UO_891 (O_891,N_28010,N_28124);
and UO_892 (O_892,N_28969,N_25021);
nor UO_893 (O_893,N_27271,N_27836);
or UO_894 (O_894,N_28720,N_29415);
nand UO_895 (O_895,N_25909,N_25547);
nand UO_896 (O_896,N_28739,N_26089);
or UO_897 (O_897,N_29246,N_26096);
xnor UO_898 (O_898,N_25810,N_29396);
nand UO_899 (O_899,N_25903,N_26512);
nor UO_900 (O_900,N_28636,N_26692);
or UO_901 (O_901,N_28893,N_26726);
nand UO_902 (O_902,N_27015,N_26870);
or UO_903 (O_903,N_26171,N_25065);
xnor UO_904 (O_904,N_25495,N_26452);
xnor UO_905 (O_905,N_26127,N_28093);
nor UO_906 (O_906,N_27632,N_29217);
or UO_907 (O_907,N_27171,N_25885);
and UO_908 (O_908,N_28087,N_28789);
xnor UO_909 (O_909,N_29698,N_27480);
or UO_910 (O_910,N_27591,N_28617);
or UO_911 (O_911,N_28021,N_27952);
or UO_912 (O_912,N_25293,N_29606);
nor UO_913 (O_913,N_28127,N_28095);
nand UO_914 (O_914,N_25169,N_28790);
nor UO_915 (O_915,N_26102,N_29566);
xnor UO_916 (O_916,N_27116,N_26408);
and UO_917 (O_917,N_28379,N_28921);
xor UO_918 (O_918,N_28034,N_26454);
nor UO_919 (O_919,N_25626,N_25423);
xor UO_920 (O_920,N_28173,N_26444);
nand UO_921 (O_921,N_27414,N_29103);
or UO_922 (O_922,N_26654,N_27139);
or UO_923 (O_923,N_28659,N_29123);
nand UO_924 (O_924,N_29600,N_26434);
or UO_925 (O_925,N_27260,N_25085);
nor UO_926 (O_926,N_25101,N_26849);
nand UO_927 (O_927,N_28137,N_27114);
nor UO_928 (O_928,N_26533,N_28043);
and UO_929 (O_929,N_29436,N_27802);
or UO_930 (O_930,N_29112,N_27405);
and UO_931 (O_931,N_27005,N_27105);
and UO_932 (O_932,N_28947,N_26627);
xnor UO_933 (O_933,N_25871,N_27701);
or UO_934 (O_934,N_27273,N_27642);
xor UO_935 (O_935,N_29447,N_29346);
nor UO_936 (O_936,N_29844,N_28186);
xnor UO_937 (O_937,N_28836,N_29517);
nor UO_938 (O_938,N_28878,N_27924);
or UO_939 (O_939,N_28324,N_28902);
xnor UO_940 (O_940,N_28119,N_27974);
xor UO_941 (O_941,N_27325,N_28801);
or UO_942 (O_942,N_29730,N_26947);
xor UO_943 (O_943,N_28618,N_25701);
xnor UO_944 (O_944,N_29323,N_26131);
nor UO_945 (O_945,N_26404,N_28579);
and UO_946 (O_946,N_29649,N_26541);
nor UO_947 (O_947,N_29556,N_27526);
nor UO_948 (O_948,N_26162,N_27306);
or UO_949 (O_949,N_27562,N_25262);
xnor UO_950 (O_950,N_27157,N_28488);
or UO_951 (O_951,N_29947,N_25850);
and UO_952 (O_952,N_28315,N_26789);
nor UO_953 (O_953,N_26751,N_25310);
and UO_954 (O_954,N_27131,N_27334);
nor UO_955 (O_955,N_28259,N_28712);
xor UO_956 (O_956,N_27944,N_27709);
nor UO_957 (O_957,N_29411,N_25779);
nor UO_958 (O_958,N_25636,N_26554);
xor UO_959 (O_959,N_28987,N_27367);
and UO_960 (O_960,N_28252,N_27227);
nor UO_961 (O_961,N_28139,N_27317);
or UO_962 (O_962,N_29463,N_29683);
nand UO_963 (O_963,N_28312,N_26905);
xnor UO_964 (O_964,N_26234,N_26229);
nor UO_965 (O_965,N_27765,N_27950);
and UO_966 (O_966,N_25352,N_28985);
xor UO_967 (O_967,N_26022,N_27238);
xnor UO_968 (O_968,N_27466,N_25544);
nor UO_969 (O_969,N_29696,N_29159);
nand UO_970 (O_970,N_25642,N_27095);
and UO_971 (O_971,N_26368,N_25682);
nand UO_972 (O_972,N_27807,N_25284);
and UO_973 (O_973,N_26461,N_27348);
xnor UO_974 (O_974,N_28880,N_25667);
and UO_975 (O_975,N_28363,N_26318);
nor UO_976 (O_976,N_29733,N_27886);
or UO_977 (O_977,N_29036,N_25321);
nor UO_978 (O_978,N_28772,N_28846);
or UO_979 (O_979,N_27059,N_27936);
xnor UO_980 (O_980,N_28380,N_25785);
xnor UO_981 (O_981,N_29397,N_25586);
nor UO_982 (O_982,N_27920,N_29035);
nand UO_983 (O_983,N_26688,N_25591);
and UO_984 (O_984,N_25693,N_27141);
xor UO_985 (O_985,N_28639,N_27379);
nand UO_986 (O_986,N_28503,N_28145);
nor UO_987 (O_987,N_27439,N_27572);
xor UO_988 (O_988,N_28484,N_29229);
nor UO_989 (O_989,N_28455,N_29225);
xor UO_990 (O_990,N_25697,N_27578);
and UO_991 (O_991,N_27941,N_29101);
or UO_992 (O_992,N_25718,N_28716);
nand UO_993 (O_993,N_27112,N_27232);
or UO_994 (O_994,N_29898,N_26384);
xnor UO_995 (O_995,N_29089,N_27143);
and UO_996 (O_996,N_26287,N_29882);
and UO_997 (O_997,N_28613,N_26819);
xnor UO_998 (O_998,N_26395,N_26347);
xnor UO_999 (O_999,N_29736,N_27148);
and UO_1000 (O_1000,N_29778,N_26596);
or UO_1001 (O_1001,N_26093,N_27115);
xor UO_1002 (O_1002,N_26348,N_25548);
xnor UO_1003 (O_1003,N_28899,N_27006);
or UO_1004 (O_1004,N_27689,N_27026);
or UO_1005 (O_1005,N_27927,N_28019);
or UO_1006 (O_1006,N_25412,N_29622);
or UO_1007 (O_1007,N_27789,N_27975);
and UO_1008 (O_1008,N_26994,N_28670);
nand UO_1009 (O_1009,N_29633,N_28785);
or UO_1010 (O_1010,N_26041,N_25280);
xor UO_1011 (O_1011,N_29405,N_26674);
or UO_1012 (O_1012,N_25239,N_27150);
nand UO_1013 (O_1013,N_27003,N_29399);
or UO_1014 (O_1014,N_26135,N_27101);
nand UO_1015 (O_1015,N_27318,N_25783);
nand UO_1016 (O_1016,N_25732,N_29678);
or UO_1017 (O_1017,N_26402,N_29984);
nor UO_1018 (O_1018,N_25242,N_27511);
nand UO_1019 (O_1019,N_29921,N_27597);
nor UO_1020 (O_1020,N_28980,N_25570);
nand UO_1021 (O_1021,N_26875,N_26269);
or UO_1022 (O_1022,N_27375,N_27274);
xnor UO_1023 (O_1023,N_25782,N_29625);
or UO_1024 (O_1024,N_26489,N_29122);
xor UO_1025 (O_1025,N_27362,N_28326);
nor UO_1026 (O_1026,N_29283,N_28272);
nor UO_1027 (O_1027,N_28704,N_26083);
xnor UO_1028 (O_1028,N_29025,N_26978);
and UO_1029 (O_1029,N_26683,N_26258);
and UO_1030 (O_1030,N_27915,N_29801);
nand UO_1031 (O_1031,N_28765,N_29684);
xor UO_1032 (O_1032,N_25184,N_27168);
xnor UO_1033 (O_1033,N_29008,N_29130);
and UO_1034 (O_1034,N_28026,N_29382);
and UO_1035 (O_1035,N_29206,N_26191);
nor UO_1036 (O_1036,N_28548,N_29714);
or UO_1037 (O_1037,N_28784,N_29723);
nand UO_1038 (O_1038,N_29378,N_28831);
and UO_1039 (O_1039,N_28285,N_28508);
and UO_1040 (O_1040,N_27988,N_27042);
nand UO_1041 (O_1041,N_28795,N_27595);
nand UO_1042 (O_1042,N_29380,N_29799);
or UO_1043 (O_1043,N_29974,N_28039);
nand UO_1044 (O_1044,N_27201,N_26062);
nor UO_1045 (O_1045,N_25951,N_25468);
nor UO_1046 (O_1046,N_26942,N_28993);
xnor UO_1047 (O_1047,N_27821,N_28094);
nor UO_1048 (O_1048,N_26232,N_29861);
nor UO_1049 (O_1049,N_27292,N_29944);
xnor UO_1050 (O_1050,N_26130,N_25902);
and UO_1051 (O_1051,N_27498,N_28117);
and UO_1052 (O_1052,N_28890,N_28623);
nand UO_1053 (O_1053,N_29629,N_29849);
or UO_1054 (O_1054,N_29645,N_29176);
nand UO_1055 (O_1055,N_28233,N_29581);
xor UO_1056 (O_1056,N_29716,N_25536);
or UO_1057 (O_1057,N_28011,N_27278);
or UO_1058 (O_1058,N_29968,N_27825);
or UO_1059 (O_1059,N_29610,N_28023);
xnor UO_1060 (O_1060,N_26609,N_27805);
nand UO_1061 (O_1061,N_29792,N_28956);
nand UO_1062 (O_1062,N_25145,N_29164);
xnor UO_1063 (O_1063,N_25605,N_29193);
xnor UO_1064 (O_1064,N_25113,N_26633);
nor UO_1065 (O_1065,N_28003,N_26551);
nor UO_1066 (O_1066,N_27242,N_25602);
and UO_1067 (O_1067,N_25288,N_29666);
nor UO_1068 (O_1068,N_26822,N_25820);
nand UO_1069 (O_1069,N_28794,N_25830);
nor UO_1070 (O_1070,N_26689,N_25984);
or UO_1071 (O_1071,N_26586,N_25182);
xor UO_1072 (O_1072,N_26577,N_26847);
or UO_1073 (O_1073,N_27345,N_25026);
xnor UO_1074 (O_1074,N_27049,N_25613);
xor UO_1075 (O_1075,N_26307,N_25425);
xor UO_1076 (O_1076,N_29679,N_27795);
or UO_1077 (O_1077,N_26670,N_25117);
nand UO_1078 (O_1078,N_29544,N_29407);
xnor UO_1079 (O_1079,N_29963,N_26743);
and UO_1080 (O_1080,N_25368,N_28747);
xnor UO_1081 (O_1081,N_26036,N_28214);
or UO_1082 (O_1082,N_25790,N_26537);
or UO_1083 (O_1083,N_29641,N_27381);
and UO_1084 (O_1084,N_28565,N_29618);
nor UO_1085 (O_1085,N_25007,N_28092);
and UO_1086 (O_1086,N_28521,N_27621);
nor UO_1087 (O_1087,N_25314,N_29617);
nor UO_1088 (O_1088,N_28123,N_29118);
nand UO_1089 (O_1089,N_29085,N_29312);
xor UO_1090 (O_1090,N_25278,N_27035);
or UO_1091 (O_1091,N_26446,N_26070);
xor UO_1092 (O_1092,N_28666,N_26207);
or UO_1093 (O_1093,N_26361,N_28141);
or UO_1094 (O_1094,N_29427,N_29973);
and UO_1095 (O_1095,N_28529,N_29750);
and UO_1096 (O_1096,N_29583,N_27460);
nand UO_1097 (O_1097,N_25846,N_28464);
xnor UO_1098 (O_1098,N_28301,N_29881);
nand UO_1099 (O_1099,N_25628,N_27797);
nand UO_1100 (O_1100,N_28262,N_29269);
or UO_1101 (O_1101,N_29302,N_29079);
xor UO_1102 (O_1102,N_28961,N_26128);
xor UO_1103 (O_1103,N_28809,N_28957);
xnor UO_1104 (O_1104,N_26735,N_26591);
nor UO_1105 (O_1105,N_29200,N_25263);
xnor UO_1106 (O_1106,N_25277,N_25857);
nand UO_1107 (O_1107,N_28777,N_26984);
xnor UO_1108 (O_1108,N_27588,N_28682);
nand UO_1109 (O_1109,N_25990,N_28370);
nand UO_1110 (O_1110,N_26951,N_28906);
nor UO_1111 (O_1111,N_27447,N_29433);
nor UO_1112 (O_1112,N_29526,N_27937);
or UO_1113 (O_1113,N_25241,N_26145);
nor UO_1114 (O_1114,N_26209,N_25897);
xnor UO_1115 (O_1115,N_28322,N_28333);
nor UO_1116 (O_1116,N_25111,N_28688);
nand UO_1117 (O_1117,N_28244,N_27474);
nand UO_1118 (O_1118,N_29388,N_26346);
nand UO_1119 (O_1119,N_26736,N_25947);
nor UO_1120 (O_1120,N_26843,N_26694);
nand UO_1121 (O_1121,N_26417,N_26064);
and UO_1122 (O_1122,N_26919,N_27648);
or UO_1123 (O_1123,N_26312,N_26747);
xnor UO_1124 (O_1124,N_29677,N_27043);
or UO_1125 (O_1125,N_26558,N_27199);
xnor UO_1126 (O_1126,N_26788,N_25911);
and UO_1127 (O_1127,N_27396,N_26693);
xor UO_1128 (O_1128,N_29426,N_27047);
and UO_1129 (O_1129,N_28584,N_25078);
and UO_1130 (O_1130,N_29417,N_25584);
nor UO_1131 (O_1131,N_27268,N_26761);
or UO_1132 (O_1132,N_28297,N_28051);
and UO_1133 (O_1133,N_28923,N_28523);
and UO_1134 (O_1134,N_29091,N_29708);
nand UO_1135 (O_1135,N_28632,N_27134);
and UO_1136 (O_1136,N_28531,N_29470);
or UO_1137 (O_1137,N_26103,N_29634);
and UO_1138 (O_1138,N_27328,N_27786);
and UO_1139 (O_1139,N_27075,N_26576);
and UO_1140 (O_1140,N_29278,N_29653);
xnor UO_1141 (O_1141,N_28368,N_28989);
xor UO_1142 (O_1142,N_26696,N_27891);
xnor UO_1143 (O_1143,N_28246,N_28491);
or UO_1144 (O_1144,N_25327,N_26352);
nand UO_1145 (O_1145,N_26535,N_28447);
xor UO_1146 (O_1146,N_28612,N_28183);
and UO_1147 (O_1147,N_26681,N_27848);
and UO_1148 (O_1148,N_29211,N_27410);
xnor UO_1149 (O_1149,N_29640,N_29569);
xor UO_1150 (O_1150,N_25227,N_28625);
and UO_1151 (O_1151,N_29287,N_27793);
nand UO_1152 (O_1152,N_25806,N_26502);
xnor UO_1153 (O_1153,N_28434,N_29360);
or UO_1154 (O_1154,N_28054,N_28442);
and UO_1155 (O_1155,N_27803,N_25179);
nand UO_1156 (O_1156,N_29545,N_25711);
and UO_1157 (O_1157,N_29480,N_29502);
nand UO_1158 (O_1158,N_28294,N_28181);
and UO_1159 (O_1159,N_29791,N_29671);
and UO_1160 (O_1160,N_27724,N_25804);
xor UO_1161 (O_1161,N_28169,N_26636);
xor UO_1162 (O_1162,N_28338,N_28001);
nand UO_1163 (O_1163,N_25390,N_28766);
xnor UO_1164 (O_1164,N_25434,N_27833);
and UO_1165 (O_1165,N_29925,N_27567);
nor UO_1166 (O_1166,N_26242,N_27252);
or UO_1167 (O_1167,N_28691,N_27403);
or UO_1168 (O_1168,N_28723,N_25622);
and UO_1169 (O_1169,N_28798,N_26326);
nand UO_1170 (O_1170,N_26695,N_25047);
and UO_1171 (O_1171,N_27729,N_29315);
and UO_1172 (O_1172,N_27766,N_27088);
and UO_1173 (O_1173,N_27746,N_26927);
or UO_1174 (O_1174,N_27720,N_26514);
or UO_1175 (O_1175,N_29163,N_25661);
or UO_1176 (O_1176,N_28757,N_28910);
nand UO_1177 (O_1177,N_27280,N_27637);
nor UO_1178 (O_1178,N_26363,N_26139);
nor UO_1179 (O_1179,N_29383,N_29726);
and UO_1180 (O_1180,N_29570,N_27969);
nor UO_1181 (O_1181,N_29319,N_29531);
xnor UO_1182 (O_1182,N_25131,N_25899);
or UO_1183 (O_1183,N_27272,N_26329);
xor UO_1184 (O_1184,N_25750,N_29924);
xor UO_1185 (O_1185,N_26109,N_28889);
and UO_1186 (O_1186,N_26007,N_29231);
nand UO_1187 (O_1187,N_29909,N_26733);
nand UO_1188 (O_1188,N_29449,N_25787);
nor UO_1189 (O_1189,N_25373,N_27794);
nand UO_1190 (O_1190,N_29406,N_25432);
nand UO_1191 (O_1191,N_29747,N_29097);
nor UO_1192 (O_1192,N_25312,N_29330);
or UO_1193 (O_1193,N_26753,N_25341);
nor UO_1194 (O_1194,N_29911,N_29598);
nor UO_1195 (O_1195,N_26763,N_27128);
nor UO_1196 (O_1196,N_26280,N_29468);
and UO_1197 (O_1197,N_25231,N_27857);
or UO_1198 (O_1198,N_26506,N_28286);
and UO_1199 (O_1199,N_28796,N_27882);
or UO_1200 (O_1200,N_25330,N_29886);
xnor UO_1201 (O_1201,N_25503,N_28828);
nand UO_1202 (O_1202,N_27099,N_29136);
and UO_1203 (O_1203,N_29110,N_29435);
xnor UO_1204 (O_1204,N_29962,N_25864);
xor UO_1205 (O_1205,N_27655,N_28934);
nand UO_1206 (O_1206,N_29847,N_28479);
xnor UO_1207 (O_1207,N_27151,N_25875);
nor UO_1208 (O_1208,N_26742,N_28793);
nand UO_1209 (O_1209,N_29661,N_28694);
and UO_1210 (O_1210,N_27773,N_25091);
nor UO_1211 (O_1211,N_27993,N_25898);
or UO_1212 (O_1212,N_25623,N_25342);
and UO_1213 (O_1213,N_27181,N_29663);
nor UO_1214 (O_1214,N_27433,N_29547);
or UO_1215 (O_1215,N_26042,N_26445);
xor UO_1216 (O_1216,N_28311,N_29342);
and UO_1217 (O_1217,N_25883,N_27061);
and UO_1218 (O_1218,N_26911,N_25549);
or UO_1219 (O_1219,N_29191,N_26931);
or UO_1220 (O_1220,N_29558,N_27783);
nand UO_1221 (O_1221,N_26289,N_28978);
nor UO_1222 (O_1222,N_25944,N_29983);
or UO_1223 (O_1223,N_29182,N_28477);
or UO_1224 (O_1224,N_29298,N_27000);
or UO_1225 (O_1225,N_27925,N_26401);
or UO_1226 (O_1226,N_29892,N_26680);
and UO_1227 (O_1227,N_27641,N_28388);
nor UO_1228 (O_1228,N_25233,N_29052);
or UO_1229 (O_1229,N_26337,N_25940);
or UO_1230 (O_1230,N_26285,N_29331);
nor UO_1231 (O_1231,N_26556,N_25121);
nand UO_1232 (O_1232,N_27978,N_26818);
xnor UO_1233 (O_1233,N_28269,N_25234);
or UO_1234 (O_1234,N_28791,N_28235);
xor UO_1235 (O_1235,N_29699,N_29444);
nand UO_1236 (O_1236,N_28621,N_29651);
nand UO_1237 (O_1237,N_28361,N_26442);
nand UO_1238 (O_1238,N_27531,N_26043);
nand UO_1239 (O_1239,N_29901,N_29813);
or UO_1240 (O_1240,N_27351,N_25583);
nand UO_1241 (O_1241,N_27419,N_29734);
or UO_1242 (O_1242,N_29472,N_25372);
nand UO_1243 (O_1243,N_29991,N_28826);
nand UO_1244 (O_1244,N_26181,N_25725);
nand UO_1245 (O_1245,N_26868,N_25712);
nor UO_1246 (O_1246,N_25888,N_29642);
and UO_1247 (O_1247,N_25132,N_29389);
and UO_1248 (O_1248,N_27788,N_28189);
xnor UO_1249 (O_1249,N_25202,N_29232);
nor UO_1250 (O_1250,N_26411,N_29919);
nor UO_1251 (O_1251,N_29132,N_25709);
nand UO_1252 (O_1252,N_28385,N_27829);
and UO_1253 (O_1253,N_28273,N_27752);
nand UO_1254 (O_1254,N_29922,N_26165);
nor UO_1255 (O_1255,N_27463,N_25896);
xnor UO_1256 (O_1256,N_29704,N_26424);
or UO_1257 (O_1257,N_29800,N_28446);
nor UO_1258 (O_1258,N_26946,N_27885);
nand UO_1259 (O_1259,N_28819,N_27333);
nand UO_1260 (O_1260,N_25627,N_25107);
nand UO_1261 (O_1261,N_28036,N_28764);
and UO_1262 (O_1262,N_28749,N_26824);
xnor UO_1263 (O_1263,N_26767,N_26645);
nand UO_1264 (O_1264,N_29913,N_27421);
nor UO_1265 (O_1265,N_27622,N_27098);
and UO_1266 (O_1266,N_27832,N_27321);
nand UO_1267 (O_1267,N_29550,N_29271);
nand UO_1268 (O_1268,N_25543,N_26357);
xor UO_1269 (O_1269,N_29753,N_25630);
xnor UO_1270 (O_1270,N_29615,N_27488);
nand UO_1271 (O_1271,N_28177,N_29014);
or UO_1272 (O_1272,N_26805,N_29139);
nand UO_1273 (O_1273,N_29044,N_25016);
xor UO_1274 (O_1274,N_29738,N_28100);
nor UO_1275 (O_1275,N_25198,N_29476);
nor UO_1276 (O_1276,N_27583,N_28002);
nand UO_1277 (O_1277,N_28678,N_28511);
and UO_1278 (O_1278,N_28974,N_28495);
nand UO_1279 (O_1279,N_28268,N_28866);
xnor UO_1280 (O_1280,N_27563,N_25287);
and UO_1281 (O_1281,N_26332,N_28377);
or UO_1282 (O_1282,N_26886,N_28727);
xor UO_1283 (O_1283,N_29223,N_27777);
or UO_1284 (O_1284,N_27176,N_26658);
or UO_1285 (O_1285,N_29013,N_25238);
xnor UO_1286 (O_1286,N_29257,N_28475);
nand UO_1287 (O_1287,N_25383,N_28851);
nand UO_1288 (O_1288,N_26270,N_26472);
xor UO_1289 (O_1289,N_25060,N_27933);
nand UO_1290 (O_1290,N_27564,N_28444);
nor UO_1291 (O_1291,N_27943,N_26910);
nor UO_1292 (O_1292,N_28563,N_27024);
and UO_1293 (O_1293,N_27624,N_27577);
and UO_1294 (O_1294,N_29304,N_27279);
or UO_1295 (O_1295,N_28706,N_27870);
xnor UO_1296 (O_1296,N_25941,N_29244);
nand UO_1297 (O_1297,N_27739,N_27366);
nor UO_1298 (O_1298,N_28422,N_26107);
and UO_1299 (O_1299,N_29374,N_28825);
nand UO_1300 (O_1300,N_28675,N_26378);
nand UO_1301 (O_1301,N_28176,N_25192);
nand UO_1302 (O_1302,N_27107,N_28895);
and UO_1303 (O_1303,N_25190,N_28387);
or UO_1304 (O_1304,N_29510,N_27364);
xor UO_1305 (O_1305,N_27865,N_26615);
nor UO_1306 (O_1306,N_26066,N_27054);
and UO_1307 (O_1307,N_25930,N_28887);
xnor UO_1308 (O_1308,N_26579,N_25208);
and UO_1309 (O_1309,N_25469,N_26920);
and UO_1310 (O_1310,N_27186,N_29209);
nand UO_1311 (O_1311,N_29337,N_26474);
or UO_1312 (O_1312,N_29240,N_28713);
or UO_1313 (O_1313,N_27690,N_25084);
nor UO_1314 (O_1314,N_25127,N_25786);
or UO_1315 (O_1315,N_28138,N_26657);
nor UO_1316 (O_1316,N_27118,N_25519);
and UO_1317 (O_1317,N_27649,N_28608);
nand UO_1318 (O_1318,N_25172,N_28342);
xnor UO_1319 (O_1319,N_28405,N_26437);
and UO_1320 (O_1320,N_26856,N_28400);
nor UO_1321 (O_1321,N_25201,N_28701);
or UO_1322 (O_1322,N_27554,N_26667);
nor UO_1323 (O_1323,N_25553,N_27389);
or UO_1324 (O_1324,N_26861,N_29024);
xnor UO_1325 (O_1325,N_25813,N_25005);
nor UO_1326 (O_1326,N_28238,N_25052);
xor UO_1327 (O_1327,N_28781,N_26065);
nor UO_1328 (O_1328,N_26431,N_28275);
nor UO_1329 (O_1329,N_25205,N_27790);
nor UO_1330 (O_1330,N_28532,N_29500);
or UO_1331 (O_1331,N_27913,N_29047);
or UO_1332 (O_1332,N_27822,N_26707);
and UO_1333 (O_1333,N_26860,N_26786);
xnor UO_1334 (O_1334,N_25754,N_29959);
and UO_1335 (O_1335,N_25500,N_27191);
nand UO_1336 (O_1336,N_27147,N_26953);
xor UO_1337 (O_1337,N_28007,N_26078);
nor UO_1338 (O_1338,N_25535,N_28105);
nand UO_1339 (O_1339,N_29506,N_27426);
xor UO_1340 (O_1340,N_29857,N_25133);
and UO_1341 (O_1341,N_29899,N_28052);
and UO_1342 (O_1342,N_26137,N_28823);
nor UO_1343 (O_1343,N_29452,N_28803);
nand UO_1344 (O_1344,N_27983,N_28172);
nand UO_1345 (O_1345,N_28835,N_28088);
and UO_1346 (O_1346,N_27532,N_25440);
or UO_1347 (O_1347,N_28597,N_29739);
or UO_1348 (O_1348,N_26222,N_29781);
or UO_1349 (O_1349,N_26097,N_26218);
and UO_1350 (O_1350,N_26543,N_26194);
or UO_1351 (O_1351,N_27958,N_26438);
or UO_1352 (O_1352,N_25045,N_27244);
and UO_1353 (O_1353,N_26260,N_29010);
xnor UO_1354 (O_1354,N_25703,N_26455);
nand UO_1355 (O_1355,N_26160,N_28759);
xor UO_1356 (O_1356,N_26023,N_25457);
nand UO_1357 (O_1357,N_29802,N_27144);
nor UO_1358 (O_1358,N_28320,N_29568);
nand UO_1359 (O_1359,N_29321,N_29064);
xnor UO_1360 (O_1360,N_26820,N_25125);
or UO_1361 (O_1361,N_29904,N_25096);
or UO_1362 (O_1362,N_26029,N_27040);
nor UO_1363 (O_1363,N_28419,N_28047);
nand UO_1364 (O_1364,N_29108,N_28212);
nand UO_1365 (O_1365,N_29111,N_27323);
nand UO_1366 (O_1366,N_26038,N_28655);
or UO_1367 (O_1367,N_25942,N_27053);
nand UO_1368 (O_1368,N_29486,N_25138);
and UO_1369 (O_1369,N_28357,N_29462);
nand UO_1370 (O_1370,N_28128,N_28522);
nor UO_1371 (O_1371,N_29591,N_28024);
nand UO_1372 (O_1372,N_25534,N_26026);
or UO_1373 (O_1373,N_27985,N_26475);
nor UO_1374 (O_1374,N_27302,N_26144);
nor UO_1375 (O_1375,N_27349,N_25621);
xor UO_1376 (O_1376,N_28452,N_27448);
or UO_1377 (O_1377,N_25408,N_26517);
or UO_1378 (O_1378,N_25203,N_25429);
xor UO_1379 (O_1379,N_26161,N_28525);
xnor UO_1380 (O_1380,N_27741,N_27558);
nand UO_1381 (O_1381,N_25077,N_27565);
nand UO_1382 (O_1382,N_26631,N_25445);
and UO_1383 (O_1383,N_28411,N_25090);
or UO_1384 (O_1384,N_27339,N_25206);
and UO_1385 (O_1385,N_29021,N_28421);
xor UO_1386 (O_1386,N_26479,N_25012);
or UO_1387 (O_1387,N_26053,N_26963);
nand UO_1388 (O_1388,N_26741,N_27764);
or UO_1389 (O_1389,N_26254,N_28863);
xnor UO_1390 (O_1390,N_27513,N_29572);
nand UO_1391 (O_1391,N_29537,N_29825);
nor UO_1392 (O_1392,N_25316,N_25403);
nor UO_1393 (O_1393,N_29521,N_26511);
or UO_1394 (O_1394,N_28671,N_28293);
nor UO_1395 (O_1395,N_29780,N_25772);
nor UO_1396 (O_1396,N_26215,N_26265);
nor UO_1397 (O_1397,N_27378,N_26734);
nor UO_1398 (O_1398,N_26245,N_26717);
nor UO_1399 (O_1399,N_25649,N_27705);
nor UO_1400 (O_1400,N_27104,N_25839);
or UO_1401 (O_1401,N_27543,N_29929);
nor UO_1402 (O_1402,N_27874,N_27894);
nor UO_1403 (O_1403,N_26021,N_28018);
or UO_1404 (O_1404,N_27347,N_27593);
or UO_1405 (O_1405,N_26034,N_27904);
and UO_1406 (O_1406,N_28025,N_26989);
xor UO_1407 (O_1407,N_26459,N_26451);
or UO_1408 (O_1408,N_29883,N_28963);
and UO_1409 (O_1409,N_25720,N_26331);
xnor UO_1410 (O_1410,N_26938,N_29081);
nor UO_1411 (O_1411,N_27879,N_29808);
nand UO_1412 (O_1412,N_29676,N_25213);
nor UO_1413 (O_1413,N_26399,N_26230);
and UO_1414 (O_1414,N_26525,N_27604);
xor UO_1415 (O_1415,N_25579,N_26048);
and UO_1416 (O_1416,N_28973,N_29349);
nor UO_1417 (O_1417,N_26651,N_26781);
xor UO_1418 (O_1418,N_26572,N_28369);
and UO_1419 (O_1419,N_25104,N_29429);
and UO_1420 (O_1420,N_26293,N_25029);
xnor UO_1421 (O_1421,N_27625,N_25915);
nor UO_1422 (O_1422,N_28992,N_28566);
nor UO_1423 (O_1423,N_28067,N_27368);
xor UO_1424 (O_1424,N_25414,N_27087);
nor UO_1425 (O_1425,N_25611,N_25333);
and UO_1426 (O_1426,N_29601,N_25834);
nor UO_1427 (O_1427,N_29418,N_25836);
and UO_1428 (O_1428,N_28216,N_25835);
nand UO_1429 (O_1429,N_25710,N_25734);
nand UO_1430 (O_1430,N_26297,N_26970);
nor UO_1431 (O_1431,N_26521,N_29333);
nand UO_1432 (O_1432,N_29142,N_25297);
nand UO_1433 (O_1433,N_27736,N_25694);
xnor UO_1434 (O_1434,N_29121,N_29620);
nand UO_1435 (O_1435,N_29934,N_25210);
and UO_1436 (O_1436,N_28435,N_27550);
and UO_1437 (O_1437,N_28131,N_26538);
and UO_1438 (O_1438,N_29786,N_27019);
or UO_1439 (O_1439,N_26015,N_28638);
nand UO_1440 (O_1440,N_29985,N_25747);
nand UO_1441 (O_1441,N_27960,N_28555);
and UO_1442 (O_1442,N_27896,N_27843);
xor UO_1443 (O_1443,N_25922,N_25475);
nand UO_1444 (O_1444,N_25222,N_27073);
nand UO_1445 (O_1445,N_28840,N_26353);
and UO_1446 (O_1446,N_27056,N_28179);
nand UO_1447 (O_1447,N_27113,N_29243);
xor UO_1448 (O_1448,N_26197,N_26629);
and UO_1449 (O_1449,N_25473,N_26184);
xor UO_1450 (O_1450,N_26366,N_25050);
nand UO_1451 (O_1451,N_29774,N_29442);
xnor UO_1452 (O_1452,N_25116,N_29737);
nand UO_1453 (O_1453,N_27919,N_25477);
or UO_1454 (O_1454,N_27768,N_27854);
nand UO_1455 (O_1455,N_28908,N_28641);
nand UO_1456 (O_1456,N_25625,N_27723);
nor UO_1457 (O_1457,N_28937,N_27606);
or UO_1458 (O_1458,N_26977,N_28854);
xor UO_1459 (O_1459,N_25695,N_28810);
nor UO_1460 (O_1460,N_27828,N_29268);
or UO_1461 (O_1461,N_26303,N_26465);
and UO_1462 (O_1462,N_25471,N_25042);
nand UO_1463 (O_1463,N_28949,N_28157);
xnor UO_1464 (O_1464,N_29098,N_27601);
nand UO_1465 (O_1465,N_28725,N_25300);
nand UO_1466 (O_1466,N_26797,N_28283);
xor UO_1467 (O_1467,N_29412,N_26869);
and UO_1468 (O_1468,N_29688,N_29768);
nand UO_1469 (O_1469,N_27500,N_28277);
xnor UO_1470 (O_1470,N_28110,N_25392);
and UO_1471 (O_1471,N_28979,N_27586);
or UO_1472 (O_1472,N_29335,N_28829);
nand UO_1473 (O_1473,N_26248,N_29976);
and UO_1474 (O_1474,N_29355,N_27121);
nor UO_1475 (O_1475,N_28399,N_26830);
xor UO_1476 (O_1476,N_26863,N_25105);
nor UO_1477 (O_1477,N_27169,N_25411);
nand UO_1478 (O_1478,N_25478,N_28227);
and UO_1479 (O_1479,N_26842,N_26037);
xnor UO_1480 (O_1480,N_25040,N_29154);
or UO_1481 (O_1481,N_25807,N_28877);
nor UO_1482 (O_1482,N_25792,N_29627);
and UO_1483 (O_1483,N_25427,N_26108);
or UO_1484 (O_1484,N_25079,N_28188);
and UO_1485 (O_1485,N_28474,N_28627);
or UO_1486 (O_1486,N_27742,N_28550);
and UO_1487 (O_1487,N_26405,N_26392);
nand UO_1488 (O_1488,N_27437,N_25243);
nand UO_1489 (O_1489,N_28770,N_28205);
nand UO_1490 (O_1490,N_27007,N_25260);
and UO_1491 (O_1491,N_28504,N_25460);
nor UO_1492 (O_1492,N_25428,N_26705);
nand UO_1493 (O_1493,N_26224,N_28078);
nand UO_1494 (O_1494,N_27434,N_27001);
and UO_1495 (O_1495,N_26074,N_26564);
xnor UO_1496 (O_1496,N_26625,N_29608);
xnor UO_1497 (O_1497,N_25721,N_28459);
and UO_1498 (O_1498,N_27710,N_29188);
nand UO_1499 (O_1499,N_29906,N_29795);
and UO_1500 (O_1500,N_27841,N_29643);
nor UO_1501 (O_1501,N_29574,N_28849);
or UO_1502 (O_1502,N_26638,N_29100);
nor UO_1503 (O_1503,N_29709,N_29422);
nor UO_1504 (O_1504,N_26199,N_25087);
nand UO_1505 (O_1505,N_28938,N_29971);
and UO_1506 (O_1506,N_26491,N_29478);
nand UO_1507 (O_1507,N_27726,N_28208);
nand UO_1508 (O_1508,N_28473,N_29393);
and UO_1509 (O_1509,N_27525,N_25775);
nand UO_1510 (O_1510,N_27475,N_25598);
and UO_1511 (O_1511,N_25527,N_28490);
xnor UO_1512 (O_1512,N_26990,N_26001);
or UO_1513 (O_1513,N_29788,N_28999);
xnor UO_1514 (O_1514,N_27342,N_29381);
and UO_1515 (O_1515,N_27399,N_27733);
nand UO_1516 (O_1516,N_29687,N_26104);
nor UO_1517 (O_1517,N_27902,N_28875);
nand UO_1518 (O_1518,N_26338,N_25393);
or UO_1519 (O_1519,N_25494,N_26132);
or UO_1520 (O_1520,N_29012,N_26439);
xnor UO_1521 (O_1521,N_27659,N_28441);
or UO_1522 (O_1522,N_29055,N_26828);
nor UO_1523 (O_1523,N_25832,N_29914);
or UO_1524 (O_1524,N_28886,N_28436);
or UO_1525 (O_1525,N_28561,N_28437);
or UO_1526 (O_1526,N_26364,N_25146);
nor UO_1527 (O_1527,N_28460,N_25788);
nor UO_1528 (O_1528,N_25726,N_27939);
nand UO_1529 (O_1529,N_27167,N_27066);
xor UO_1530 (O_1530,N_28270,N_25842);
nor UO_1531 (O_1531,N_28236,N_29731);
nor UO_1532 (O_1532,N_26082,N_25358);
or UO_1533 (O_1533,N_27300,N_27194);
nor UO_1534 (O_1534,N_27076,N_29630);
nor UO_1535 (O_1535,N_27528,N_28986);
or UO_1536 (O_1536,N_25812,N_27987);
nor UO_1537 (O_1537,N_29834,N_26871);
nor UO_1538 (O_1538,N_26117,N_27065);
nor UO_1539 (O_1539,N_27892,N_25868);
or UO_1540 (O_1540,N_29168,N_25340);
or UO_1541 (O_1541,N_26003,N_25152);
nor UO_1542 (O_1542,N_25151,N_29473);
or UO_1543 (O_1543,N_25039,N_25593);
and UO_1544 (O_1544,N_28356,N_28767);
nand UO_1545 (O_1545,N_26779,N_26895);
nand UO_1546 (O_1546,N_29018,N_27108);
and UO_1547 (O_1547,N_26727,N_29889);
or UO_1548 (O_1548,N_25696,N_28045);
nand UO_1549 (O_1549,N_26407,N_27725);
and UO_1550 (O_1550,N_29254,N_26433);
or UO_1551 (O_1551,N_25530,N_26833);
xnor UO_1552 (O_1552,N_28211,N_29945);
or UO_1553 (O_1553,N_25872,N_25256);
nand UO_1554 (O_1554,N_29867,N_25264);
nand UO_1555 (O_1555,N_25143,N_25688);
xnor UO_1556 (O_1556,N_29571,N_27413);
xor UO_1557 (O_1557,N_26166,N_27253);
xnor UO_1558 (O_1558,N_26485,N_28193);
nor UO_1559 (O_1559,N_28959,N_29548);
nor UO_1560 (O_1560,N_28744,N_27514);
xor UO_1561 (O_1561,N_28852,N_29037);
xnor UO_1562 (O_1562,N_25589,N_25529);
nand UO_1563 (O_1563,N_27908,N_27164);
or UO_1564 (O_1564,N_28493,N_27551);
and UO_1565 (O_1565,N_26669,N_25706);
or UO_1566 (O_1566,N_29611,N_26468);
or UO_1567 (O_1567,N_26580,N_26562);
or UO_1568 (O_1568,N_27671,N_29207);
and UO_1569 (O_1569,N_27607,N_25196);
or UO_1570 (O_1570,N_26721,N_27487);
nor UO_1571 (O_1571,N_29212,N_25103);
or UO_1572 (O_1572,N_28383,N_29151);
or UO_1573 (O_1573,N_27057,N_28159);
nand UO_1574 (O_1574,N_27454,N_26801);
nor UO_1575 (O_1575,N_28113,N_25357);
and UO_1576 (O_1576,N_28834,N_27887);
and UO_1577 (O_1577,N_27255,N_26762);
xnor UO_1578 (O_1578,N_28722,N_26610);
nor UO_1579 (O_1579,N_26370,N_26208);
nor UO_1580 (O_1580,N_26811,N_27269);
and UO_1581 (O_1581,N_25784,N_28647);
xnor UO_1582 (O_1582,N_26678,N_25236);
xor UO_1583 (O_1583,N_29848,N_29724);
and UO_1584 (O_1584,N_28845,N_26955);
or UO_1585 (O_1585,N_28448,N_27459);
nor UO_1586 (O_1586,N_27771,N_27834);
and UO_1587 (O_1587,N_25967,N_26172);
or UO_1588 (O_1588,N_29770,N_25961);
or UO_1589 (O_1589,N_29063,N_28629);
nand UO_1590 (O_1590,N_25936,N_28885);
nand UO_1591 (O_1591,N_25765,N_27211);
or UO_1592 (O_1592,N_27976,N_26529);
and UO_1593 (O_1593,N_29839,N_27267);
or UO_1594 (O_1594,N_25195,N_26150);
or UO_1595 (O_1595,N_29241,N_26185);
nor UO_1596 (O_1596,N_26758,N_27435);
xnor UO_1597 (O_1597,N_28116,N_27429);
or UO_1598 (O_1598,N_27859,N_28614);
and UO_1599 (O_1599,N_26880,N_26791);
nand UO_1600 (O_1600,N_26566,N_27613);
xnor UO_1601 (O_1601,N_28330,N_25698);
xnor UO_1602 (O_1602,N_26712,N_25554);
and UO_1603 (O_1603,N_25677,N_28808);
or UO_1604 (O_1604,N_28102,N_26996);
or UO_1605 (O_1605,N_29941,N_28328);
xor UO_1606 (O_1606,N_26593,N_25112);
or UO_1607 (O_1607,N_27721,N_25576);
or UO_1608 (O_1608,N_27002,N_25108);
or UO_1609 (O_1609,N_28527,N_27942);
nor UO_1610 (O_1610,N_27561,N_25419);
xor UO_1611 (O_1611,N_25374,N_26879);
nor UO_1612 (O_1612,N_29961,N_27796);
nor UO_1613 (O_1613,N_28850,N_29507);
nand UO_1614 (O_1614,N_25949,N_27576);
nor UO_1615 (O_1615,N_26239,N_25369);
nand UO_1616 (O_1616,N_26928,N_29662);
nor UO_1617 (O_1617,N_27778,N_29410);
and UO_1618 (O_1618,N_28184,N_27603);
nor UO_1619 (O_1619,N_29668,N_27866);
or UO_1620 (O_1620,N_28554,N_25400);
nand UO_1621 (O_1621,N_29395,N_27022);
nand UO_1622 (O_1622,N_28865,N_26567);
nor UO_1623 (O_1623,N_28323,N_27961);
or UO_1624 (O_1624,N_26441,N_27233);
nor UO_1625 (O_1625,N_28298,N_27445);
xor UO_1626 (O_1626,N_26087,N_26808);
xor UO_1627 (O_1627,N_28750,N_28998);
or UO_1628 (O_1628,N_28698,N_25295);
and UO_1629 (O_1629,N_25525,N_27130);
nand UO_1630 (O_1630,N_29910,N_29420);
nor UO_1631 (O_1631,N_26518,N_29826);
and UO_1632 (O_1632,N_25604,N_26381);
xor UO_1633 (O_1633,N_27647,N_29970);
and UO_1634 (O_1634,N_29453,N_26457);
and UO_1635 (O_1635,N_29487,N_28151);
nand UO_1636 (O_1636,N_25794,N_27515);
nor UO_1637 (O_1637,N_26359,N_25991);
xnor UO_1638 (O_1638,N_25954,N_26221);
or UO_1639 (O_1639,N_29681,N_25620);
or UO_1640 (O_1640,N_27468,N_25756);
nor UO_1641 (O_1641,N_27313,N_25200);
or UO_1642 (O_1642,N_27137,N_25689);
and UO_1643 (O_1643,N_27307,N_26080);
and UO_1644 (O_1644,N_25847,N_29954);
xnor UO_1645 (O_1645,N_26634,N_29007);
and UO_1646 (O_1646,N_29077,N_27898);
nand UO_1647 (O_1647,N_27083,N_27486);
xor UO_1648 (O_1648,N_27992,N_28967);
and UO_1649 (O_1649,N_25063,N_29377);
or UO_1650 (O_1650,N_25998,N_29949);
and UO_1651 (O_1651,N_25860,N_28888);
xnor UO_1652 (O_1652,N_29448,N_25153);
xnor UO_1653 (O_1653,N_29807,N_27438);
nor UO_1654 (O_1654,N_27820,N_26024);
nor UO_1655 (O_1655,N_26030,N_26649);
or UO_1656 (O_1656,N_28656,N_28012);
xnor UO_1657 (O_1657,N_25746,N_26700);
nand UO_1658 (O_1658,N_26320,N_26673);
or UO_1659 (O_1659,N_26918,N_26853);
nand UO_1660 (O_1660,N_28263,N_25824);
xnor UO_1661 (O_1661,N_27400,N_25890);
xor UO_1662 (O_1662,N_25574,N_25464);
nand UO_1663 (O_1663,N_28243,N_29213);
nor UO_1664 (O_1664,N_28458,N_26993);
or UO_1665 (O_1665,N_28546,N_26134);
nor UO_1666 (O_1666,N_27740,N_25166);
xor UO_1667 (O_1667,N_25489,N_26011);
xor UO_1668 (O_1668,N_26900,N_28753);
xor UO_1669 (O_1669,N_26557,N_25517);
and UO_1670 (O_1670,N_29364,N_27450);
and UO_1671 (O_1671,N_25165,N_26855);
nor UO_1672 (O_1672,N_27966,N_28056);
or UO_1673 (O_1673,N_26999,N_25676);
nor UO_1674 (O_1674,N_28071,N_29490);
xor UO_1675 (O_1675,N_29685,N_27295);
xnor UO_1676 (O_1676,N_28339,N_26279);
and UO_1677 (O_1677,N_25291,N_27240);
nor UO_1678 (O_1678,N_26618,N_25338);
xor UO_1679 (O_1679,N_29978,N_28560);
or UO_1680 (O_1680,N_27219,N_27173);
nor UO_1681 (O_1681,N_25881,N_25587);
xor UO_1682 (O_1682,N_27774,N_29862);
xnor UO_1683 (O_1683,N_27998,N_27142);
nor UO_1684 (O_1684,N_26826,N_25879);
nand UO_1685 (O_1685,N_29931,N_29201);
and UO_1686 (O_1686,N_27013,N_28742);
nand UO_1687 (O_1687,N_26604,N_25030);
or UO_1688 (O_1688,N_26415,N_25714);
xnor UO_1689 (O_1689,N_28314,N_28853);
and UO_1690 (O_1690,N_29369,N_27584);
nor UO_1691 (O_1691,N_29893,N_26908);
or UO_1692 (O_1692,N_29872,N_25929);
nor UO_1693 (O_1693,N_27417,N_26450);
nand UO_1694 (O_1694,N_28578,N_28855);
nand UO_1695 (O_1695,N_27889,N_29715);
or UO_1696 (O_1696,N_26858,N_25672);
or UO_1697 (O_1697,N_29782,N_28786);
xor UO_1698 (O_1698,N_25894,N_25130);
and UO_1699 (O_1699,N_29814,N_29595);
nand UO_1700 (O_1700,N_29325,N_28997);
nor UO_1701 (O_1701,N_25218,N_25062);
and UO_1702 (O_1702,N_29587,N_29259);
nor UO_1703 (O_1703,N_25669,N_28407);
or UO_1704 (O_1704,N_28367,N_28006);
or UO_1705 (O_1705,N_26316,N_28748);
xor UO_1706 (O_1706,N_28253,N_28251);
or UO_1707 (O_1707,N_26817,N_25715);
xor UO_1708 (O_1708,N_28637,N_26142);
xnor UO_1709 (O_1709,N_25037,N_25092);
and UO_1710 (O_1710,N_27372,N_27407);
xor UO_1711 (O_1711,N_27772,N_28848);
and UO_1712 (O_1712,N_26060,N_29181);
and UO_1713 (O_1713,N_26652,N_28942);
nor UO_1714 (O_1714,N_26764,N_29439);
and UO_1715 (O_1715,N_26055,N_26719);
nor UO_1716 (O_1716,N_26383,N_25474);
or UO_1717 (O_1717,N_28345,N_29482);
nand UO_1718 (O_1718,N_26388,N_29869);
nand UO_1719 (O_1719,N_25054,N_28225);
or UO_1720 (O_1720,N_29794,N_27497);
xor UO_1721 (O_1721,N_26420,N_27432);
or UO_1722 (O_1722,N_25305,N_27331);
and UO_1723 (O_1723,N_29365,N_28773);
nand UO_1724 (O_1724,N_27880,N_28871);
and UO_1725 (O_1725,N_29040,N_29043);
nor UO_1726 (O_1726,N_26063,N_26328);
and UO_1727 (O_1727,N_27989,N_27161);
or UO_1728 (O_1728,N_29060,N_29772);
nand UO_1729 (O_1729,N_28496,N_27537);
xnor UO_1730 (O_1730,N_29023,N_26613);
nand UO_1731 (O_1731,N_25119,N_27804);
nor UO_1732 (O_1732,N_29140,N_29096);
and UO_1733 (O_1733,N_26892,N_28668);
and UO_1734 (O_1734,N_25422,N_27283);
and UO_1735 (O_1735,N_27570,N_27877);
or UO_1736 (O_1736,N_28965,N_28945);
nand UO_1737 (O_1737,N_29955,N_28103);
nor UO_1738 (O_1738,N_28050,N_25662);
nor UO_1739 (O_1739,N_26903,N_27156);
nand UO_1740 (O_1740,N_28797,N_26585);
xor UO_1741 (O_1741,N_26965,N_26403);
xor UO_1742 (O_1742,N_26759,N_28168);
nor UO_1743 (O_1743,N_27340,N_25286);
nand UO_1744 (O_1744,N_25496,N_25803);
nor UO_1745 (O_1745,N_27449,N_28292);
nand UO_1746 (O_1746,N_28375,N_29061);
or UO_1747 (O_1747,N_25176,N_26581);
nor UO_1748 (O_1748,N_27155,N_28505);
nand UO_1749 (O_1749,N_27918,N_25313);
or UO_1750 (O_1750,N_28042,N_28680);
nor UO_1751 (O_1751,N_27336,N_28994);
nand UO_1752 (O_1752,N_29529,N_29149);
xor UO_1753 (O_1753,N_27646,N_27900);
or UO_1754 (O_1754,N_25071,N_26009);
xnor UO_1755 (O_1755,N_27304,N_27585);
xnor UO_1756 (O_1756,N_26530,N_29803);
xor UO_1757 (O_1757,N_29362,N_29592);
xnor UO_1758 (O_1758,N_25585,N_28896);
and UO_1759 (O_1759,N_26012,N_26897);
nor UO_1760 (O_1760,N_27360,N_26589);
nor UO_1761 (O_1761,N_26745,N_29870);
and UO_1762 (O_1762,N_28501,N_27212);
and UO_1763 (O_1763,N_26201,N_26487);
or UO_1764 (O_1764,N_28187,N_28048);
nand UO_1765 (O_1765,N_29935,N_29549);
nand UO_1766 (O_1766,N_25350,N_25446);
xor UO_1767 (O_1767,N_26324,N_27172);
nand UO_1768 (O_1768,N_25540,N_28858);
nand UO_1769 (O_1769,N_29534,N_26740);
and UO_1770 (O_1770,N_29757,N_28821);
or UO_1771 (O_1771,N_28881,N_27698);
xnor UO_1772 (O_1772,N_29308,N_25265);
or UO_1773 (O_1773,N_27954,N_29523);
nand UO_1774 (O_1774,N_27747,N_26969);
nand UO_1775 (O_1775,N_26825,N_27738);
or UO_1776 (O_1776,N_29345,N_28334);
nor UO_1777 (O_1777,N_25845,N_28472);
nand UO_1778 (O_1778,N_25512,N_29197);
and UO_1779 (O_1779,N_25800,N_29208);
and UO_1780 (O_1780,N_29964,N_27485);
nor UO_1781 (O_1781,N_25267,N_29811);
or UO_1782 (O_1782,N_27517,N_27028);
or UO_1783 (O_1783,N_27187,N_27645);
and UO_1784 (O_1784,N_29752,N_27265);
nand UO_1785 (O_1785,N_26526,N_29863);
or UO_1786 (O_1786,N_29262,N_27388);
nand UO_1787 (O_1787,N_28386,N_25663);
and UO_1788 (O_1788,N_28950,N_29824);
nor UO_1789 (O_1789,N_28390,N_25865);
and UO_1790 (O_1790,N_29234,N_28860);
nand UO_1791 (O_1791,N_29218,N_29199);
xnor UO_1792 (O_1792,N_27962,N_27623);
nand UO_1793 (O_1793,N_29741,N_26504);
nand UO_1794 (O_1794,N_27262,N_27734);
nand UO_1795 (O_1795,N_26807,N_27058);
nand UO_1796 (O_1796,N_25394,N_26077);
nand UO_1797 (O_1797,N_25880,N_27755);
or UO_1798 (O_1798,N_29841,N_28538);
nor UO_1799 (O_1799,N_29026,N_27955);
nor UO_1800 (O_1800,N_25818,N_28649);
and UO_1801 (O_1801,N_27327,N_27767);
or UO_1802 (O_1802,N_28991,N_26106);
nand UO_1803 (O_1803,N_27986,N_29589);
xor UO_1804 (O_1804,N_29751,N_29664);
or UO_1805 (O_1805,N_29637,N_25237);
nor UO_1806 (O_1806,N_28951,N_29401);
nor UO_1807 (O_1807,N_25124,N_25728);
nor UO_1808 (O_1808,N_28708,N_28977);
or UO_1809 (O_1809,N_27427,N_28282);
and UO_1810 (O_1810,N_27408,N_28990);
or UO_1811 (O_1811,N_29495,N_29327);
xnor UO_1812 (O_1812,N_26375,N_27697);
xor UO_1813 (O_1813,N_25937,N_29039);
or UO_1814 (O_1814,N_28883,N_27712);
and UO_1815 (O_1815,N_29525,N_27949);
nand UO_1816 (O_1816,N_27228,N_26720);
xnor UO_1817 (O_1817,N_29347,N_29141);
nor UO_1818 (O_1818,N_29066,N_28572);
nand UO_1819 (O_1819,N_29169,N_29912);
or UO_1820 (O_1820,N_25159,N_29351);
and UO_1821 (O_1821,N_27472,N_27580);
nand UO_1822 (O_1822,N_26846,N_26251);
and UO_1823 (O_1823,N_26987,N_25673);
nor UO_1824 (O_1824,N_25268,N_26275);
nor UO_1825 (O_1825,N_26193,N_28537);
or UO_1826 (O_1826,N_29392,N_26272);
xnor UO_1827 (O_1827,N_26238,N_25004);
and UO_1828 (O_1828,N_25702,N_28358);
nand UO_1829 (O_1829,N_25150,N_28931);
xnor UO_1830 (O_1830,N_29125,N_25743);
and UO_1831 (O_1831,N_29607,N_28687);
nor UO_1832 (O_1832,N_27217,N_26350);
xor UO_1833 (O_1833,N_27650,N_28449);
nand UO_1834 (O_1834,N_25640,N_28519);
or UO_1835 (O_1835,N_25590,N_29987);
nand UO_1836 (O_1836,N_25498,N_25081);
or UO_1837 (O_1837,N_25907,N_29940);
xor UO_1838 (O_1838,N_27346,N_28009);
nand UO_1839 (O_1839,N_27965,N_26587);
nor UO_1840 (O_1840,N_25656,N_27045);
and UO_1841 (O_1841,N_28081,N_26950);
nand UO_1842 (O_1842,N_28944,N_25089);
or UO_1843 (O_1843,N_25931,N_25036);
nand UO_1844 (O_1844,N_27782,N_27298);
or UO_1845 (O_1845,N_26914,N_29357);
nor UO_1846 (O_1846,N_29993,N_25347);
and UO_1847 (O_1847,N_28303,N_27246);
and UO_1848 (O_1848,N_26100,N_25207);
xor UO_1849 (O_1849,N_27165,N_27930);
nor UO_1850 (O_1850,N_26299,N_25684);
nand UO_1851 (O_1851,N_28745,N_25798);
nor UO_1852 (O_1852,N_25456,N_25158);
xnor UO_1853 (O_1853,N_26785,N_29359);
nand UO_1854 (O_1854,N_29403,N_25916);
nand UO_1855 (O_1855,N_27917,N_28607);
or UO_1856 (O_1856,N_25816,N_27731);
and UO_1857 (O_1857,N_27566,N_27670);
or UO_1858 (O_1858,N_28199,N_25235);
nor UO_1859 (O_1859,N_25298,N_28015);
nand UO_1860 (O_1860,N_25455,N_29527);
xnor UO_1861 (O_1861,N_29031,N_27749);
xor UO_1862 (O_1862,N_28818,N_25541);
nand UO_1863 (O_1863,N_25363,N_28362);
xor UO_1864 (O_1864,N_29338,N_26490);
nor UO_1865 (O_1865,N_28063,N_26929);
nor UO_1866 (O_1866,N_28289,N_29528);
or UO_1867 (O_1867,N_27856,N_26988);
and UO_1868 (O_1868,N_27995,N_27012);
xnor UO_1869 (O_1869,N_28709,N_29559);
and UO_1870 (O_1870,N_25046,N_27792);
xnor UO_1871 (O_1871,N_27494,N_27291);
or UO_1872 (O_1872,N_26710,N_26583);
or UO_1873 (O_1873,N_29354,N_25962);
or UO_1874 (O_1874,N_29660,N_28911);
nor UO_1875 (O_1875,N_29951,N_28469);
nand UO_1876 (O_1876,N_28382,N_28806);
nor UO_1877 (O_1877,N_26772,N_27813);
or UO_1878 (O_1878,N_26553,N_28109);
nand UO_1879 (O_1879,N_26902,N_29465);
or UO_1880 (O_1880,N_27787,N_29432);
nand UO_1881 (O_1881,N_25164,N_27582);
nand UO_1882 (O_1882,N_25659,N_28892);
nand UO_1883 (O_1883,N_25925,N_25906);
nand UO_1884 (O_1884,N_27728,N_29290);
nor UO_1885 (O_1885,N_28971,N_29038);
and UO_1886 (O_1886,N_29127,N_29563);
or UO_1887 (O_1887,N_27170,N_26650);
or UO_1888 (O_1888,N_25999,N_26425);
nand UO_1889 (O_1889,N_26616,N_25617);
nor UO_1890 (O_1890,N_29198,N_28663);
nor UO_1891 (O_1891,N_26056,N_27046);
and UO_1892 (O_1892,N_25675,N_26373);
or UO_1893 (O_1893,N_26288,N_25632);
nand UO_1894 (O_1894,N_29596,N_28864);
nor UO_1895 (O_1895,N_25355,N_25670);
and UO_1896 (O_1896,N_29457,N_29960);
xnor UO_1897 (O_1897,N_29113,N_25367);
nand UO_1898 (O_1898,N_28718,N_25057);
xor UO_1899 (O_1899,N_26813,N_26448);
nand UO_1900 (O_1900,N_27146,N_25122);
xnor UO_1901 (O_1901,N_27241,N_28569);
and UO_1902 (O_1902,N_28874,N_25247);
xor UO_1903 (O_1903,N_25299,N_25729);
or UO_1904 (O_1904,N_27004,N_29313);
nor UO_1905 (O_1905,N_28278,N_27594);
nand UO_1906 (O_1906,N_25799,N_28966);
or UO_1907 (O_1907,N_28897,N_29656);
xor UO_1908 (O_1908,N_25599,N_29590);
nand UO_1909 (O_1909,N_29192,N_25502);
nand UO_1910 (O_1910,N_25189,N_25142);
xnor UO_1911 (O_1911,N_27506,N_27779);
nor UO_1912 (O_1912,N_29988,N_25421);
or UO_1913 (O_1913,N_29019,N_29455);
xor UO_1914 (O_1914,N_26005,N_26508);
or UO_1915 (O_1915,N_25003,N_26413);
or UO_1916 (O_1916,N_25228,N_27380);
or UO_1917 (O_1917,N_26340,N_27206);
and UO_1918 (O_1918,N_25537,N_25666);
xor UO_1919 (O_1919,N_27991,N_28894);
nand UO_1920 (O_1920,N_27270,N_29742);
or UO_1921 (O_1921,N_28804,N_29918);
and UO_1922 (O_1922,N_29504,N_25687);
and UO_1923 (O_1923,N_28221,N_29247);
or UO_1924 (O_1924,N_29859,N_28861);
nor UO_1925 (O_1925,N_27288,N_29033);
nor UO_1926 (O_1926,N_27644,N_29042);
xnor UO_1927 (O_1927,N_29932,N_29552);
or UO_1928 (O_1928,N_26766,N_27781);
nor UO_1929 (O_1929,N_25639,N_29580);
nand UO_1930 (O_1930,N_27446,N_26536);
xnor UO_1931 (O_1931,N_28250,N_25566);
nand UO_1932 (O_1932,N_28587,N_28677);
and UO_1933 (O_1933,N_29536,N_27737);
xor UO_1934 (O_1934,N_29238,N_29745);
nand UO_1935 (O_1935,N_28602,N_27869);
nor UO_1936 (O_1936,N_27996,N_26206);
nand UO_1937 (O_1937,N_28946,N_27640);
nand UO_1938 (O_1938,N_29868,N_29773);
nand UO_1939 (O_1939,N_27033,N_27871);
or UO_1940 (O_1940,N_28833,N_26039);
or UO_1941 (O_1941,N_27055,N_29692);
and UO_1942 (O_1942,N_29562,N_28242);
xnor UO_1943 (O_1943,N_26872,N_29838);
xnor UO_1944 (O_1944,N_27875,N_25507);
and UO_1945 (O_1945,N_29255,N_26916);
nand UO_1946 (O_1946,N_27549,N_29843);
nor UO_1947 (O_1947,N_26204,N_29059);
xnor UO_1948 (O_1948,N_29146,N_28486);
nand UO_1949 (O_1949,N_28842,N_27858);
or UO_1950 (O_1950,N_26476,N_26611);
xor UO_1951 (O_1951,N_29686,N_28152);
xor UO_1952 (O_1952,N_29272,N_26010);
or UO_1953 (O_1953,N_26575,N_29505);
nor UO_1954 (O_1954,N_26799,N_29195);
or UO_1955 (O_1955,N_26595,N_28223);
and UO_1956 (O_1956,N_27831,N_28820);
and UO_1957 (O_1957,N_25289,N_28787);
nor UO_1958 (O_1958,N_25578,N_27195);
nor UO_1959 (O_1959,N_29908,N_26432);
xor UO_1960 (O_1960,N_26906,N_29057);
and UO_1961 (O_1961,N_29511,N_29576);
nor UO_1962 (O_1962,N_25161,N_25398);
or UO_1963 (O_1963,N_26973,N_27060);
and UO_1964 (O_1964,N_27997,N_28308);
or UO_1965 (O_1965,N_28304,N_25430);
or UO_1966 (O_1966,N_28085,N_29720);
and UO_1967 (O_1967,N_29475,N_29126);
or UO_1968 (O_1968,N_28904,N_27127);
or UO_1969 (O_1969,N_28300,N_27509);
xnor UO_1970 (O_1970,N_29703,N_25893);
nand UO_1971 (O_1971,N_28589,N_28738);
or UO_1972 (O_1972,N_28544,N_29669);
or UO_1973 (O_1973,N_26691,N_27629);
nand UO_1974 (O_1974,N_29840,N_28933);
and UO_1975 (O_1975,N_25275,N_26574);
nor UO_1976 (O_1976,N_25230,N_25332);
nor UO_1977 (O_1977,N_27223,N_25733);
and UO_1978 (O_1978,N_26306,N_29896);
or UO_1979 (O_1979,N_28427,N_29995);
and UO_1980 (O_1980,N_28337,N_29107);
xor UO_1981 (O_1981,N_25643,N_25306);
and UO_1982 (O_1982,N_26752,N_27473);
nand UO_1983 (O_1983,N_25406,N_29441);
nand UO_1984 (O_1984,N_28096,N_25882);
nand UO_1985 (O_1985,N_28305,N_25567);
or UO_1986 (O_1986,N_28536,N_28372);
nand UO_1987 (O_1987,N_25170,N_27881);
or UO_1988 (O_1988,N_25452,N_25552);
or UO_1989 (O_1989,N_29353,N_28567);
xor UO_1990 (O_1990,N_27489,N_26369);
xnor UO_1991 (O_1991,N_28568,N_28118);
and UO_1992 (O_1992,N_28027,N_28276);
xor UO_1993 (O_1993,N_26544,N_26315);
nor UO_1994 (O_1994,N_29251,N_27153);
or UO_1995 (O_1995,N_29819,N_29344);
xnor UO_1996 (O_1996,N_25467,N_29939);
or UO_1997 (O_1997,N_29358,N_26716);
xnor UO_1998 (O_1998,N_26941,N_26769);
nand UO_1999 (O_1999,N_29155,N_29454);
nand UO_2000 (O_2000,N_29821,N_28426);
nand UO_2001 (O_2001,N_26663,N_28843);
nor UO_2002 (O_2002,N_28175,N_29068);
and UO_2003 (O_2003,N_25952,N_28354);
xnor UO_2004 (O_2004,N_25981,N_28916);
nor UO_2005 (O_2005,N_26146,N_25304);
xnor UO_2006 (O_2006,N_27756,N_25748);
xnor UO_2007 (O_2007,N_25051,N_26342);
xor UO_2008 (O_2008,N_29300,N_28482);
nand UO_2009 (O_2009,N_29652,N_25252);
nand UO_2010 (O_2010,N_25356,N_27068);
and UO_2011 (O_2011,N_28594,N_27633);
or UO_2012 (O_2012,N_27082,N_27322);
nor UO_2013 (O_2013,N_29286,N_26236);
nor UO_2014 (O_2014,N_25248,N_28976);
nor UO_2015 (O_2015,N_27314,N_27404);
xor UO_2016 (O_2016,N_27533,N_29363);
xnor UO_2017 (O_2017,N_25488,N_27014);
nor UO_2018 (O_2018,N_27666,N_26435);
and UO_2019 (O_2019,N_26806,N_27527);
nor UO_2020 (O_2020,N_26278,N_27928);
nand UO_2021 (O_2021,N_28941,N_26488);
or UO_2022 (O_2022,N_27769,N_29084);
and UO_2023 (O_2023,N_27261,N_25232);
nor UO_2024 (O_2024,N_28097,N_29053);
or UO_2025 (O_2025,N_29612,N_26898);
nor UO_2026 (O_2026,N_26151,N_29171);
nor UO_2027 (O_2027,N_28443,N_26261);
nand UO_2028 (O_2028,N_28163,N_26701);
nand UO_2029 (O_2029,N_27681,N_27178);
nor UO_2030 (O_2030,N_28046,N_28414);
nand UO_2031 (O_2031,N_27744,N_25307);
or UO_2032 (O_2032,N_27284,N_26498);
nor UO_2033 (O_2033,N_26072,N_28838);
or UO_2034 (O_2034,N_25521,N_26981);
nor UO_2035 (O_2035,N_25044,N_28241);
xor UO_2036 (O_2036,N_26644,N_28606);
nand UO_2037 (O_2037,N_26632,N_29842);
or UO_2038 (O_2038,N_27661,N_26386);
xnor UO_2039 (O_2039,N_28299,N_29334);
or UO_2040 (O_2040,N_29204,N_25652);
and UO_2041 (O_2041,N_28577,N_26081);
or UO_2042 (O_2042,N_26019,N_28222);
and UO_2043 (O_2043,N_27179,N_28907);
nor UO_2044 (O_2044,N_29990,N_26188);
nor UO_2045 (O_2045,N_25018,N_28530);
xor UO_2046 (O_2046,N_29145,N_27032);
xnor UO_2047 (O_2047,N_27350,N_29148);
nand UO_2048 (O_2048,N_29348,N_29659);
and UO_2049 (O_2049,N_29804,N_29479);
and UO_2050 (O_2050,N_25410,N_27763);
or UO_2051 (O_2051,N_27677,N_27162);
and UO_2052 (O_2052,N_29477,N_27693);
and UO_2053 (O_2053,N_27418,N_29340);
and UO_2054 (O_2054,N_28690,N_28758);
or UO_2055 (O_2055,N_27873,N_27010);
or UO_2056 (O_2056,N_29494,N_25240);
and UO_2057 (O_2057,N_29758,N_26061);
xnor UO_2058 (O_2058,N_25226,N_29080);
nor UO_2059 (O_2059,N_28167,N_25716);
nor UO_2060 (O_2060,N_29082,N_26954);
nand UO_2061 (O_2061,N_29373,N_29789);
and UO_2062 (O_2062,N_27906,N_25863);
nand UO_2063 (O_2063,N_26774,N_26703);
xnor UO_2064 (O_2064,N_28811,N_27257);
and UO_2065 (O_2065,N_27863,N_28033);
and UO_2066 (O_2066,N_27316,N_25852);
or UO_2067 (O_2067,N_27688,N_29602);
xnor UO_2068 (O_2068,N_27051,N_26008);
nand UO_2069 (O_2069,N_25386,N_28037);
xor UO_2070 (O_2070,N_25932,N_28652);
xor UO_2071 (O_2071,N_25470,N_26527);
or UO_2072 (O_2072,N_25526,N_26210);
and UO_2073 (O_2073,N_27938,N_28280);
xor UO_2074 (O_2074,N_26214,N_26884);
or UO_2075 (O_2075,N_27651,N_29667);
nor UO_2076 (O_2076,N_25843,N_29109);
nand UO_2077 (O_2077,N_26917,N_27070);
nand UO_2078 (O_2078,N_29196,N_26850);
nand UO_2079 (O_2079,N_28373,N_28398);
nor UO_2080 (O_2080,N_29776,N_27522);
and UO_2081 (O_2081,N_27508,N_27442);
nand UO_2082 (O_2082,N_26714,N_25463);
nor UO_2083 (O_2083,N_25129,N_27132);
or UO_2084 (O_2084,N_25778,N_28182);
xnor UO_2085 (O_2085,N_28514,N_29051);
nor UO_2086 (O_2086,N_28013,N_29203);
xor UO_2087 (O_2087,N_27149,N_29965);
nand UO_2088 (O_2088,N_27326,N_27470);
and UO_2089 (O_2089,N_27373,N_27420);
and UO_2090 (O_2090,N_28349,N_28755);
or UO_2091 (O_2091,N_26836,N_26492);
nand UO_2092 (O_2092,N_26154,N_27495);
or UO_2093 (O_2093,N_26790,N_29299);
nand UO_2094 (O_2094,N_25776,N_29459);
and UO_2095 (O_2095,N_27482,N_27129);
and UO_2096 (O_2096,N_28717,N_26484);
nor UO_2097 (O_2097,N_25055,N_26757);
xnor UO_2098 (O_2098,N_28062,N_28053);
or UO_2099 (O_2099,N_28111,N_25437);
nor UO_2100 (O_2100,N_29264,N_27979);
or UO_2101 (O_2101,N_27492,N_29499);
nand UO_2102 (O_2102,N_25571,N_26602);
nand UO_2103 (O_2103,N_25435,N_27980);
or UO_2104 (O_2104,N_28404,N_28107);
xor UO_2105 (O_2105,N_29887,N_25518);
xor UO_2106 (O_2106,N_28905,N_29582);
or UO_2107 (O_2107,N_26866,N_26059);
nor UO_2108 (O_2108,N_25829,N_26547);
xor UO_2109 (O_2109,N_26322,N_27111);
nand UO_2110 (O_2110,N_28943,N_26715);
nand UO_2111 (O_2111,N_27652,N_25913);
xor UO_2112 (O_2112,N_27852,N_27398);
or UO_2113 (O_2113,N_26934,N_25730);
or UO_2114 (O_2114,N_28343,N_27687);
nand UO_2115 (O_2115,N_29372,N_27914);
xor UO_2116 (O_2116,N_25752,N_28430);
and UO_2117 (O_2117,N_29852,N_27669);
and UO_2118 (O_2118,N_28210,N_25647);
nand UO_2119 (O_2119,N_29890,N_29413);
and UO_2120 (O_2120,N_28674,N_28202);
and UO_2121 (O_2121,N_25315,N_26980);
or UO_2122 (O_2122,N_27627,N_27209);
nor UO_2123 (O_2123,N_26243,N_29464);
nand UO_2124 (O_2124,N_28224,N_29520);
xor UO_2125 (O_2125,N_29878,N_28673);
and UO_2126 (O_2126,N_29981,N_28098);
or UO_2127 (O_2127,N_28463,N_27386);
or UO_2128 (O_2128,N_26330,N_25343);
nor UO_2129 (O_2129,N_25141,N_28635);
and UO_2130 (O_2130,N_29041,N_28507);
nor UO_2131 (O_2131,N_28476,N_26084);
and UO_2132 (O_2132,N_27499,N_25595);
xor UO_2133 (O_2133,N_26800,N_27415);
and UO_2134 (O_2134,N_27338,N_26211);
or UO_2135 (O_2135,N_29016,N_28676);
nand UO_2136 (O_2136,N_28585,N_25665);
or UO_2137 (O_2137,N_28703,N_25155);
nor UO_2138 (O_2138,N_29414,N_26686);
nor UO_2139 (O_2139,N_26174,N_26308);
nand UO_2140 (O_2140,N_28288,N_25960);
nor UO_2141 (O_2141,N_25629,N_28763);
and UO_2142 (O_2142,N_28970,N_28309);
nand UO_2143 (O_2143,N_29020,N_29655);
nor UO_2144 (O_2144,N_29029,N_28327);
nor UO_2145 (O_2145,N_27215,N_27390);
and UO_2146 (O_2146,N_26971,N_29823);
nand UO_2147 (O_2147,N_25874,N_25533);
or UO_2148 (O_2148,N_27236,N_26051);
or UO_2149 (O_2149,N_27839,N_27361);
or UO_2150 (O_2150,N_28410,N_28595);
and UO_2151 (O_2151,N_28513,N_25485);
nor UO_2152 (O_2152,N_25397,N_28891);
or UO_2153 (O_2153,N_29398,N_27229);
or UO_2154 (O_2154,N_25274,N_25034);
or UO_2155 (O_2155,N_28350,N_28462);
nor UO_2156 (O_2156,N_26500,N_29638);
nand UO_2157 (O_2157,N_29322,N_29691);
nor UO_2158 (O_2158,N_28075,N_26648);
and UO_2159 (O_2159,N_25869,N_27719);
or UO_2160 (O_2160,N_29846,N_25840);
or UO_2161 (O_2161,N_28445,N_26878);
nor UO_2162 (O_2162,N_29586,N_25377);
nand UO_2163 (O_2163,N_29816,N_26877);
nand UO_2164 (O_2164,N_28237,N_28915);
nand UO_2165 (O_2165,N_29281,N_27247);
nor UO_2166 (O_2166,N_28072,N_28939);
xnor UO_2167 (O_2167,N_28213,N_26466);
or UO_2168 (O_2168,N_28814,N_28267);
or UO_2169 (O_2169,N_27231,N_26831);
xnor UO_2170 (O_2170,N_26561,N_28453);
xnor UO_2171 (O_2171,N_26032,N_25759);
xor UO_2172 (O_2172,N_29690,N_27277);
and UO_2173 (O_2173,N_25199,N_26419);
nand UO_2174 (O_2174,N_28144,N_26704);
xor UO_2175 (O_2175,N_25965,N_27743);
or UO_2176 (O_2176,N_25011,N_28130);
nor UO_2177 (O_2177,N_29515,N_28030);
nand UO_2178 (O_2178,N_26276,N_29658);
or UO_2179 (O_2179,N_29138,N_29104);
and UO_2180 (O_2180,N_26578,N_28397);
and UO_2181 (O_2181,N_29328,N_28603);
and UO_2182 (O_2182,N_27308,N_28083);
and UO_2183 (O_2183,N_26212,N_28365);
or UO_2184 (O_2184,N_25048,N_27761);
nor UO_2185 (O_2185,N_28428,N_29927);
and UO_2186 (O_2186,N_29936,N_28166);
and UO_2187 (O_2187,N_25744,N_26972);
xnor UO_2188 (O_2188,N_29421,N_25093);
xnor UO_2189 (O_2189,N_29524,N_25767);
nand UO_2190 (O_2190,N_26612,N_29485);
or UO_2191 (O_2191,N_28909,N_29894);
or UO_2192 (O_2192,N_28140,N_29837);
or UO_2193 (O_2193,N_25921,N_27899);
or UO_2194 (O_2194,N_25508,N_25175);
nor UO_2195 (O_2195,N_27823,N_29003);
nand UO_2196 (O_2196,N_26471,N_25031);
xor UO_2197 (O_2197,N_27182,N_25515);
nor UO_2198 (O_2198,N_25214,N_27387);
or UO_2199 (O_2199,N_27192,N_29443);
and UO_2200 (O_2200,N_29034,N_26300);
nand UO_2201 (O_2201,N_28769,N_29806);
and UO_2202 (O_2202,N_25774,N_27617);
nor UO_2203 (O_2203,N_28955,N_29948);
or UO_2204 (O_2204,N_28643,N_26956);
or UO_2205 (O_2205,N_28084,N_28775);
or UO_2206 (O_2206,N_27956,N_26882);
and UO_2207 (O_2207,N_27050,N_26894);
nand UO_2208 (O_2208,N_25106,N_25266);
nor UO_2209 (O_2209,N_29402,N_26246);
nand UO_2210 (O_2210,N_29070,N_27039);
and UO_2211 (O_2211,N_28558,N_28408);
nor UO_2212 (O_2212,N_29597,N_29700);
xnor UO_2213 (O_2213,N_27798,N_27190);
nor UO_2214 (O_2214,N_25817,N_26390);
xor UO_2215 (O_2215,N_29157,N_27842);
or UO_2216 (O_2216,N_25853,N_27539);
or UO_2217 (O_2217,N_28733,N_28700);
xnor UO_2218 (O_2218,N_27668,N_29616);
nand UO_2219 (O_2219,N_26277,N_25704);
and UO_2220 (O_2220,N_26773,N_26573);
xor UO_2221 (O_2221,N_25851,N_25964);
and UO_2222 (O_2222,N_27727,N_26962);
nand UO_2223 (O_2223,N_25439,N_25431);
and UO_2224 (O_2224,N_27819,N_29706);
or UO_2225 (O_2225,N_28217,N_28605);
nand UO_2226 (O_2226,N_26909,N_27878);
nor UO_2227 (O_2227,N_25416,N_26050);
nor UO_2228 (O_2228,N_29866,N_29356);
xor UO_2229 (O_2229,N_26904,N_25318);
and UO_2230 (O_2230,N_27573,N_25956);
xnor UO_2231 (O_2231,N_29385,N_25660);
nor UO_2232 (O_2232,N_27855,N_29916);
and UO_2233 (O_2233,N_26164,N_26501);
and UO_2234 (O_2234,N_27453,N_27476);
nor UO_2235 (O_2235,N_27197,N_29175);
nand UO_2236 (O_2236,N_28249,N_25395);
or UO_2237 (O_2237,N_26076,N_28154);
or UO_2238 (O_2238,N_29689,N_26203);
nor UO_2239 (O_2239,N_26816,N_27827);
nor UO_2240 (O_2240,N_25193,N_28816);
or UO_2241 (O_2241,N_27912,N_29001);
nand UO_2242 (O_2242,N_28032,N_29946);
nand UO_2243 (O_2243,N_28014,N_25099);
or UO_2244 (O_2244,N_25975,N_25861);
or UO_2245 (O_2245,N_26812,N_27600);
and UO_2246 (O_2246,N_28953,N_27214);
xor UO_2247 (O_2247,N_29865,N_26409);
nor UO_2248 (O_2248,N_26186,N_28384);
and UO_2249 (O_2249,N_28900,N_29294);
nor UO_2250 (O_2250,N_28715,N_25738);
xor UO_2251 (O_2251,N_26231,N_26635);
nor UO_2252 (O_2252,N_29682,N_25838);
xor UO_2253 (O_2253,N_29967,N_29317);
or UO_2254 (O_2254,N_29851,N_26158);
and UO_2255 (O_2255,N_29071,N_28234);
nor UO_2256 (O_2256,N_25147,N_29818);
xor UO_2257 (O_2257,N_28332,N_29252);
and UO_2258 (O_2258,N_28940,N_27203);
and UO_2259 (O_2259,N_26028,N_26656);
xnor UO_2260 (O_2260,N_29292,N_28040);
nand UO_2261 (O_2261,N_28868,N_28583);
nor UO_2262 (O_2262,N_25770,N_29236);
or UO_2263 (O_2263,N_26731,N_25259);
and UO_2264 (O_2264,N_27353,N_28080);
or UO_2265 (O_2265,N_27812,N_25588);
xor UO_2266 (O_2266,N_28642,N_25939);
xnor UO_2267 (O_2267,N_27618,N_29184);
nor UO_2268 (O_2268,N_29074,N_26213);
or UO_2269 (O_2269,N_28256,N_29288);
xnor UO_2270 (O_2270,N_26075,N_29624);
and UO_2271 (O_2271,N_26302,N_25946);
or UO_2272 (O_2272,N_25487,N_27135);
xnor UO_2273 (O_2273,N_26389,N_28547);
xor UO_2274 (O_2274,N_27299,N_26274);
and UO_2275 (O_2275,N_29787,N_28667);
xor UO_2276 (O_2276,N_25740,N_29790);
and UO_2277 (O_2277,N_26961,N_25074);
xor UO_2278 (O_2278,N_25067,N_25041);
nor UO_2279 (O_2279,N_26495,N_28813);
and UO_2280 (O_2280,N_27290,N_29779);
and UO_2281 (O_2281,N_28432,N_29746);
xor UO_2282 (O_2282,N_25844,N_28412);
and UO_2283 (O_2283,N_29533,N_25802);
nand UO_2284 (O_2284,N_27008,N_26937);
xnor UO_2285 (O_2285,N_25674,N_28958);
and UO_2286 (O_2286,N_25815,N_29594);
or UO_2287 (O_2287,N_27397,N_25580);
nor UO_2288 (O_2288,N_27612,N_27154);
nor UO_2289 (O_2289,N_29614,N_28935);
nor UO_2290 (O_2290,N_28413,N_27830);
nor UO_2291 (O_2291,N_26334,N_28431);
nand UO_2292 (O_2292,N_29273,N_25957);
xor UO_2293 (O_2293,N_29361,N_26690);
or UO_2294 (O_2294,N_26344,N_25749);
nand UO_2295 (O_2295,N_27444,N_29194);
nand UO_2296 (O_2296,N_28347,N_29538);
nand UO_2297 (O_2297,N_26045,N_26200);
and UO_2298 (O_2298,N_28196,N_27656);
nand UO_2299 (O_2299,N_25808,N_28170);
or UO_2300 (O_2300,N_25644,N_28901);
nor UO_2301 (O_2301,N_26033,N_28539);
nor UO_2302 (O_2302,N_25015,N_29320);
or UO_2303 (O_2303,N_28228,N_26398);
nor UO_2304 (O_2304,N_28968,N_29431);
nor UO_2305 (O_2305,N_28059,N_28433);
nand UO_2306 (O_2306,N_27968,N_26071);
or UO_2307 (O_2307,N_27320,N_29874);
nor UO_2308 (O_2308,N_28640,N_27067);
and UO_2309 (O_2309,N_28215,N_25615);
nor UO_2310 (O_2310,N_28425,N_28402);
and UO_2311 (O_2311,N_25582,N_26356);
or UO_2312 (O_2312,N_25405,N_27694);
or UO_2313 (O_2313,N_28207,N_25841);
or UO_2314 (O_2314,N_29030,N_26120);
xnor UO_2315 (O_2315,N_29297,N_25809);
xor UO_2316 (O_2316,N_25969,N_26216);
or UO_2317 (O_2317,N_28494,N_26068);
xnor UO_2318 (O_2318,N_28451,N_29239);
or UO_2319 (O_2319,N_29707,N_25724);
xnor UO_2320 (O_2320,N_26114,N_26992);
nor UO_2321 (O_2321,N_26771,N_25510);
nand UO_2322 (O_2322,N_26545,N_25825);
nand UO_2323 (O_2323,N_25509,N_29275);
xor UO_2324 (O_2324,N_28325,N_25186);
and UO_2325 (O_2325,N_27286,N_27717);
and UO_2326 (O_2326,N_26428,N_27750);
xnor UO_2327 (O_2327,N_25866,N_28520);
nand UO_2328 (O_2328,N_29619,N_28424);
nor UO_2329 (O_2329,N_28551,N_27423);
or UO_2330 (O_2330,N_27074,N_26675);
xor UO_2331 (O_2331,N_29777,N_28065);
nand UO_2332 (O_2332,N_26520,N_25178);
nand UO_2333 (O_2333,N_26163,N_25136);
nor UO_2334 (O_2334,N_26247,N_26778);
xnor UO_2335 (O_2335,N_29532,N_26156);
or UO_2336 (O_2336,N_25354,N_26000);
xor UO_2337 (O_2337,N_28679,N_29665);
nand UO_2338 (O_2338,N_26621,N_25379);
and UO_2339 (O_2339,N_25449,N_28126);
or UO_2340 (O_2340,N_25311,N_29561);
nand UO_2341 (O_2341,N_29979,N_26220);
and UO_2342 (O_2342,N_27560,N_26661);
or UO_2343 (O_2343,N_29710,N_29810);
nand UO_2344 (O_2344,N_26244,N_29162);
and UO_2345 (O_2345,N_28134,N_28239);
nor UO_2346 (O_2346,N_25828,N_25551);
nor UO_2347 (O_2347,N_25109,N_26429);
nand UO_2348 (O_2348,N_26509,N_29028);
nor UO_2349 (O_2349,N_26827,N_28396);
nor UO_2350 (O_2350,N_26341,N_26601);
nor UO_2351 (O_2351,N_28355,N_25995);
xor UO_2352 (O_2352,N_27732,N_28928);
and UO_2353 (O_2353,N_26679,N_26426);
nand UO_2354 (O_2354,N_27817,N_29765);
xnor UO_2355 (O_2355,N_25924,N_26423);
and UO_2356 (O_2356,N_29258,N_25319);
nor UO_2357 (O_2357,N_25450,N_25174);
xnor UO_2358 (O_2358,N_28149,N_26503);
nand UO_2359 (O_2359,N_26534,N_28936);
nor UO_2360 (O_2360,N_28604,N_29086);
nor UO_2361 (O_2361,N_25123,N_25797);
nor UO_2362 (O_2362,N_25637,N_25281);
or UO_2363 (O_2363,N_26623,N_25134);
nor UO_2364 (O_2364,N_29280,N_29266);
and UO_2365 (O_2365,N_28714,N_29214);
xnor UO_2366 (O_2366,N_26513,N_25745);
and UO_2367 (O_2367,N_26159,N_25923);
xnor UO_2368 (O_2368,N_26031,N_25276);
nor UO_2369 (O_2369,N_25895,N_28616);
xor UO_2370 (O_2370,N_29695,N_27245);
xor UO_2371 (O_2371,N_28601,N_25870);
or UO_2372 (O_2372,N_27953,N_28573);
xnor UO_2373 (O_2373,N_25811,N_27851);
nor UO_2374 (O_2374,N_29877,N_28862);
and UO_2375 (O_2375,N_28702,N_25066);
nor UO_2376 (O_2376,N_28352,N_27479);
nor UO_2377 (O_2377,N_26569,N_26559);
nor UO_2378 (O_2378,N_29579,N_28089);
nor UO_2379 (O_2379,N_26319,N_28499);
and UO_2380 (O_2380,N_29375,N_26647);
nor UO_2381 (O_2381,N_28844,N_26848);
xor UO_2382 (O_2382,N_27748,N_27078);
and UO_2383 (O_2383,N_25978,N_25320);
nand UO_2384 (O_2384,N_29516,N_28147);
nor UO_2385 (O_2385,N_26939,N_28440);
or UO_2386 (O_2386,N_26851,N_29829);
nand UO_2387 (O_2387,N_27205,N_26964);
or UO_2388 (O_2388,N_26532,N_27758);
nand UO_2389 (O_2389,N_29957,N_29928);
nand UO_2390 (O_2390,N_27947,N_27970);
nor UO_2391 (O_2391,N_29416,N_29567);
nand UO_2392 (O_2392,N_26571,N_28857);
nand UO_2393 (O_2393,N_26153,N_29680);
nand UO_2394 (O_2394,N_29518,N_26982);
nor UO_2395 (O_2395,N_29897,N_26986);
nand UO_2396 (O_2396,N_25144,N_27089);
nor UO_2397 (O_2397,N_26073,N_25963);
and UO_2398 (O_2398,N_27092,N_28760);
or UO_2399 (O_2399,N_29705,N_28185);
nor UO_2400 (O_2400,N_29326,N_28570);
nand UO_2401 (O_2401,N_25436,N_27826);
and UO_2402 (O_2402,N_28918,N_29267);
and UO_2403 (O_2403,N_26718,N_26960);
xnor UO_2404 (O_2404,N_27025,N_27910);
xor UO_2405 (O_2405,N_26677,N_25859);
xor UO_2406 (O_2406,N_27216,N_28420);
or UO_2407 (O_2407,N_27312,N_26935);
nand UO_2408 (O_2408,N_27735,N_27964);
nand UO_2409 (O_2409,N_25017,N_28534);
xnor UO_2410 (O_2410,N_27838,N_25465);
nand UO_2411 (O_2411,N_29430,N_26546);
xnor UO_2412 (O_2412,N_28101,N_27596);
xnor UO_2413 (O_2413,N_27254,N_27175);
nor UO_2414 (O_2414,N_25538,N_28295);
and UO_2415 (O_2415,N_26301,N_26367);
nor UO_2416 (O_2416,N_25301,N_25577);
and UO_2417 (O_2417,N_29303,N_25168);
nor UO_2418 (O_2418,N_27138,N_26641);
or UO_2419 (O_2419,N_25154,N_29888);
xor UO_2420 (O_2420,N_26113,N_26264);
nand UO_2421 (O_2421,N_29083,N_29760);
or UO_2422 (O_2422,N_27808,N_26706);
or UO_2423 (O_2423,N_27534,N_25114);
nand UO_2424 (O_2424,N_29508,N_25378);
nand UO_2425 (O_2425,N_26496,N_29493);
nand UO_2426 (O_2426,N_27084,N_25359);
or UO_2427 (O_2427,N_28924,N_26262);
nor UO_2428 (O_2428,N_29722,N_29920);
nor UO_2429 (O_2429,N_28599,N_25891);
or UO_2430 (O_2430,N_28466,N_29379);
nand UO_2431 (O_2431,N_26768,N_26115);
nand UO_2432 (O_2432,N_29588,N_28500);
or UO_2433 (O_2433,N_26169,N_29895);
nor UO_2434 (O_2434,N_25769,N_26837);
and UO_2435 (O_2435,N_29648,N_25491);
nor UO_2436 (O_2436,N_27174,N_25255);
and UO_2437 (O_2437,N_25098,N_26412);
nor UO_2438 (O_2438,N_25461,N_27602);
nor UO_2439 (O_2439,N_28079,N_29221);
nand UO_2440 (O_2440,N_27911,N_25953);
nor UO_2441 (O_2441,N_29519,N_25056);
or UO_2442 (O_2442,N_26362,N_29093);
nor UO_2443 (O_2443,N_29265,N_27963);
and UO_2444 (O_2444,N_28693,N_26555);
xnor UO_2445 (O_2445,N_26149,N_27620);
xnor UO_2446 (O_2446,N_27097,N_29564);
nand UO_2447 (O_2447,N_26891,N_27977);
and UO_2448 (O_2448,N_28066,N_29419);
xnor UO_2449 (O_2449,N_27753,N_29227);
nand UO_2450 (O_2450,N_27575,N_25943);
xor UO_2451 (O_2451,N_27903,N_29509);
and UO_2452 (O_2452,N_27011,N_25511);
nand UO_2453 (O_2453,N_27062,N_27628);
or UO_2454 (O_2454,N_28783,N_27850);
or UO_2455 (O_2455,N_25972,N_26088);
xor UO_2456 (O_2456,N_29073,N_26462);
nand UO_2457 (O_2457,N_28165,N_29005);
xor UO_2458 (O_2458,N_26979,N_26803);
nand UO_2459 (O_2459,N_25927,N_26646);
xor UO_2460 (O_2460,N_28148,N_27072);
xnor UO_2461 (O_2461,N_26699,N_26637);
xor UO_2462 (O_2462,N_29492,N_28524);
nand UO_2463 (O_2463,N_28265,N_25873);
nor UO_2464 (O_2464,N_28664,N_28450);
nor UO_2465 (O_2465,N_28266,N_25349);
nor UO_2466 (O_2466,N_28439,N_26118);
xor UO_2467 (O_2467,N_25302,N_26628);
xor UO_2468 (O_2468,N_27547,N_29131);
and UO_2469 (O_2469,N_29498,N_29474);
and UO_2470 (O_2470,N_27630,N_28378);
and UO_2471 (O_2471,N_29975,N_26798);
nor UO_2472 (O_2472,N_29827,N_25118);
xor UO_2473 (O_2473,N_28729,N_28774);
xor UO_2474 (O_2474,N_27119,N_28153);
and UO_2475 (O_2475,N_25006,N_27598);
xor UO_2476 (O_2476,N_25049,N_29626);
and UO_2477 (O_2477,N_27682,N_25361);
nor UO_2478 (O_2478,N_26480,N_28721);
or UO_2479 (O_2479,N_25826,N_28394);
xor UO_2480 (O_2480,N_25211,N_27662);
nand UO_2481 (O_2481,N_29553,N_25493);
nand UO_2482 (O_2482,N_28344,N_28255);
or UO_2483 (O_2483,N_25713,N_27907);
xor UO_2484 (O_2484,N_25608,N_27849);
xor UO_2485 (O_2485,N_25934,N_29306);
or UO_2486 (O_2486,N_29905,N_27031);
nand UO_2487 (O_2487,N_28226,N_25220);
nand UO_2488 (O_2488,N_29256,N_25385);
and UO_2489 (O_2489,N_28981,N_29577);
xnor UO_2490 (O_2490,N_26888,N_29721);
nand UO_2491 (O_2491,N_29324,N_27478);
nand UO_2492 (O_2492,N_28553,N_27096);
or UO_2493 (O_2493,N_26178,N_25568);
nand UO_2494 (O_2494,N_27196,N_27080);
and UO_2495 (O_2495,N_28710,N_28734);
or UO_2496 (O_2496,N_25646,N_27016);
and UO_2497 (O_2497,N_26857,N_26528);
nor UO_2498 (O_2498,N_29650,N_25619);
or UO_2499 (O_2499,N_28657,N_25486);
xor UO_2500 (O_2500,N_29893,N_25974);
nor UO_2501 (O_2501,N_28808,N_29921);
nor UO_2502 (O_2502,N_25281,N_26561);
nand UO_2503 (O_2503,N_27428,N_26918);
and UO_2504 (O_2504,N_25515,N_29562);
nor UO_2505 (O_2505,N_26440,N_29479);
and UO_2506 (O_2506,N_28270,N_28502);
nand UO_2507 (O_2507,N_28283,N_26681);
nor UO_2508 (O_2508,N_26841,N_26240);
and UO_2509 (O_2509,N_26641,N_25008);
or UO_2510 (O_2510,N_29684,N_26036);
nor UO_2511 (O_2511,N_27926,N_29858);
and UO_2512 (O_2512,N_27310,N_28325);
or UO_2513 (O_2513,N_28124,N_25852);
xnor UO_2514 (O_2514,N_29312,N_26616);
nand UO_2515 (O_2515,N_27365,N_26050);
and UO_2516 (O_2516,N_29048,N_26612);
nor UO_2517 (O_2517,N_28339,N_25547);
nand UO_2518 (O_2518,N_27960,N_27044);
xor UO_2519 (O_2519,N_27382,N_28614);
nand UO_2520 (O_2520,N_27715,N_26152);
and UO_2521 (O_2521,N_26183,N_27561);
xnor UO_2522 (O_2522,N_28805,N_26926);
or UO_2523 (O_2523,N_29650,N_25461);
xnor UO_2524 (O_2524,N_29973,N_25704);
xor UO_2525 (O_2525,N_28748,N_26159);
xor UO_2526 (O_2526,N_28289,N_28904);
nand UO_2527 (O_2527,N_29092,N_25078);
and UO_2528 (O_2528,N_25383,N_26050);
nand UO_2529 (O_2529,N_28598,N_26864);
nor UO_2530 (O_2530,N_25803,N_29608);
nor UO_2531 (O_2531,N_26257,N_26632);
and UO_2532 (O_2532,N_25420,N_26390);
and UO_2533 (O_2533,N_29160,N_27862);
nor UO_2534 (O_2534,N_28031,N_28781);
nand UO_2535 (O_2535,N_29514,N_28953);
and UO_2536 (O_2536,N_29277,N_26253);
and UO_2537 (O_2537,N_27628,N_26161);
xor UO_2538 (O_2538,N_28665,N_29486);
and UO_2539 (O_2539,N_25695,N_26537);
nor UO_2540 (O_2540,N_26195,N_29392);
and UO_2541 (O_2541,N_28189,N_29593);
and UO_2542 (O_2542,N_27965,N_27196);
xor UO_2543 (O_2543,N_27764,N_26414);
and UO_2544 (O_2544,N_28492,N_27968);
or UO_2545 (O_2545,N_28973,N_25972);
nand UO_2546 (O_2546,N_25657,N_28069);
and UO_2547 (O_2547,N_25385,N_27080);
and UO_2548 (O_2548,N_29676,N_26391);
xnor UO_2549 (O_2549,N_26584,N_25085);
and UO_2550 (O_2550,N_25690,N_29283);
and UO_2551 (O_2551,N_28012,N_26082);
xnor UO_2552 (O_2552,N_29751,N_29161);
xnor UO_2553 (O_2553,N_27416,N_25171);
nor UO_2554 (O_2554,N_29537,N_27428);
nor UO_2555 (O_2555,N_28656,N_26236);
xnor UO_2556 (O_2556,N_28746,N_25920);
nor UO_2557 (O_2557,N_26803,N_27372);
nor UO_2558 (O_2558,N_26915,N_26267);
and UO_2559 (O_2559,N_29761,N_27279);
or UO_2560 (O_2560,N_27733,N_27456);
nor UO_2561 (O_2561,N_28166,N_27818);
xor UO_2562 (O_2562,N_25773,N_25421);
xor UO_2563 (O_2563,N_25509,N_28740);
and UO_2564 (O_2564,N_27231,N_28953);
and UO_2565 (O_2565,N_29904,N_28093);
xnor UO_2566 (O_2566,N_26009,N_28592);
and UO_2567 (O_2567,N_26534,N_29172);
xnor UO_2568 (O_2568,N_26523,N_25578);
and UO_2569 (O_2569,N_25927,N_27137);
and UO_2570 (O_2570,N_25801,N_26751);
xor UO_2571 (O_2571,N_28575,N_25036);
nand UO_2572 (O_2572,N_25788,N_26963);
or UO_2573 (O_2573,N_27603,N_26875);
nor UO_2574 (O_2574,N_25061,N_25825);
xor UO_2575 (O_2575,N_25556,N_26457);
or UO_2576 (O_2576,N_26054,N_28660);
nand UO_2577 (O_2577,N_27200,N_29363);
or UO_2578 (O_2578,N_26619,N_28338);
nand UO_2579 (O_2579,N_27710,N_27647);
nand UO_2580 (O_2580,N_29220,N_26584);
or UO_2581 (O_2581,N_29227,N_26702);
nor UO_2582 (O_2582,N_26206,N_28728);
nor UO_2583 (O_2583,N_25432,N_28903);
nand UO_2584 (O_2584,N_28236,N_26724);
xor UO_2585 (O_2585,N_26030,N_27909);
xor UO_2586 (O_2586,N_27291,N_29934);
and UO_2587 (O_2587,N_25415,N_29824);
xor UO_2588 (O_2588,N_28684,N_25564);
nand UO_2589 (O_2589,N_26804,N_27669);
or UO_2590 (O_2590,N_29205,N_27618);
nand UO_2591 (O_2591,N_29361,N_25319);
and UO_2592 (O_2592,N_25115,N_27678);
nand UO_2593 (O_2593,N_28832,N_28540);
and UO_2594 (O_2594,N_28996,N_27548);
and UO_2595 (O_2595,N_27861,N_28840);
nor UO_2596 (O_2596,N_26295,N_26507);
and UO_2597 (O_2597,N_26920,N_26772);
xnor UO_2598 (O_2598,N_25729,N_25331);
and UO_2599 (O_2599,N_29971,N_29714);
nor UO_2600 (O_2600,N_28484,N_27981);
nor UO_2601 (O_2601,N_25580,N_26032);
nand UO_2602 (O_2602,N_29514,N_25120);
nand UO_2603 (O_2603,N_25247,N_28113);
xor UO_2604 (O_2604,N_26132,N_25637);
and UO_2605 (O_2605,N_28263,N_26580);
xor UO_2606 (O_2606,N_29026,N_26058);
or UO_2607 (O_2607,N_28654,N_26522);
nor UO_2608 (O_2608,N_25854,N_25002);
nand UO_2609 (O_2609,N_25380,N_28395);
nand UO_2610 (O_2610,N_28621,N_28389);
and UO_2611 (O_2611,N_26128,N_25049);
xor UO_2612 (O_2612,N_28470,N_26453);
and UO_2613 (O_2613,N_27846,N_26251);
xor UO_2614 (O_2614,N_26373,N_27548);
and UO_2615 (O_2615,N_27968,N_27017);
or UO_2616 (O_2616,N_26947,N_25131);
xor UO_2617 (O_2617,N_28552,N_26420);
or UO_2618 (O_2618,N_29546,N_27704);
xnor UO_2619 (O_2619,N_29382,N_29094);
xor UO_2620 (O_2620,N_26040,N_29496);
nand UO_2621 (O_2621,N_27369,N_25647);
and UO_2622 (O_2622,N_28239,N_27359);
and UO_2623 (O_2623,N_28487,N_25420);
nor UO_2624 (O_2624,N_28365,N_27511);
xnor UO_2625 (O_2625,N_26088,N_26095);
nand UO_2626 (O_2626,N_26607,N_29316);
nor UO_2627 (O_2627,N_28766,N_28528);
xor UO_2628 (O_2628,N_26445,N_25362);
or UO_2629 (O_2629,N_27420,N_25595);
xnor UO_2630 (O_2630,N_25783,N_29599);
nor UO_2631 (O_2631,N_29774,N_28316);
or UO_2632 (O_2632,N_27914,N_28102);
nor UO_2633 (O_2633,N_29064,N_28613);
xor UO_2634 (O_2634,N_27918,N_25618);
nor UO_2635 (O_2635,N_25780,N_29067);
and UO_2636 (O_2636,N_27237,N_26133);
xnor UO_2637 (O_2637,N_25911,N_27030);
nand UO_2638 (O_2638,N_26706,N_25466);
or UO_2639 (O_2639,N_29708,N_27619);
and UO_2640 (O_2640,N_26423,N_29347);
nand UO_2641 (O_2641,N_25938,N_29776);
and UO_2642 (O_2642,N_26148,N_29156);
and UO_2643 (O_2643,N_25989,N_25058);
nor UO_2644 (O_2644,N_29910,N_28662);
or UO_2645 (O_2645,N_26375,N_27840);
or UO_2646 (O_2646,N_27318,N_29387);
xor UO_2647 (O_2647,N_25506,N_27662);
and UO_2648 (O_2648,N_25584,N_29070);
and UO_2649 (O_2649,N_25071,N_28512);
xnor UO_2650 (O_2650,N_29150,N_26584);
or UO_2651 (O_2651,N_29056,N_27307);
nand UO_2652 (O_2652,N_29187,N_26203);
and UO_2653 (O_2653,N_29040,N_28098);
nor UO_2654 (O_2654,N_26183,N_29833);
and UO_2655 (O_2655,N_26973,N_28661);
xor UO_2656 (O_2656,N_26658,N_25916);
nor UO_2657 (O_2657,N_26055,N_29499);
nand UO_2658 (O_2658,N_28676,N_25415);
and UO_2659 (O_2659,N_26966,N_26061);
or UO_2660 (O_2660,N_27762,N_27831);
xor UO_2661 (O_2661,N_27545,N_25863);
xnor UO_2662 (O_2662,N_26558,N_28790);
nor UO_2663 (O_2663,N_25879,N_27406);
xnor UO_2664 (O_2664,N_25888,N_29293);
xor UO_2665 (O_2665,N_28074,N_26268);
nand UO_2666 (O_2666,N_28113,N_29441);
or UO_2667 (O_2667,N_27251,N_28219);
nor UO_2668 (O_2668,N_27260,N_29276);
and UO_2669 (O_2669,N_26264,N_27644);
nor UO_2670 (O_2670,N_27235,N_26096);
xnor UO_2671 (O_2671,N_28576,N_27856);
and UO_2672 (O_2672,N_29191,N_26263);
nor UO_2673 (O_2673,N_26514,N_25226);
nand UO_2674 (O_2674,N_29556,N_25921);
xor UO_2675 (O_2675,N_28790,N_29438);
nand UO_2676 (O_2676,N_25694,N_27468);
or UO_2677 (O_2677,N_28948,N_29381);
nor UO_2678 (O_2678,N_26811,N_27237);
nand UO_2679 (O_2679,N_26571,N_25822);
and UO_2680 (O_2680,N_28982,N_25686);
and UO_2681 (O_2681,N_29542,N_28937);
or UO_2682 (O_2682,N_26043,N_28150);
or UO_2683 (O_2683,N_28142,N_26118);
nand UO_2684 (O_2684,N_26588,N_29326);
or UO_2685 (O_2685,N_25490,N_28754);
and UO_2686 (O_2686,N_26816,N_25959);
or UO_2687 (O_2687,N_29823,N_29317);
nor UO_2688 (O_2688,N_25495,N_29724);
or UO_2689 (O_2689,N_28734,N_29836);
or UO_2690 (O_2690,N_27581,N_28920);
and UO_2691 (O_2691,N_29669,N_25280);
xnor UO_2692 (O_2692,N_29611,N_25957);
nand UO_2693 (O_2693,N_26091,N_28572);
xnor UO_2694 (O_2694,N_26356,N_26178);
or UO_2695 (O_2695,N_27644,N_26046);
nor UO_2696 (O_2696,N_28258,N_26630);
nor UO_2697 (O_2697,N_29294,N_26842);
xor UO_2698 (O_2698,N_27748,N_28671);
nand UO_2699 (O_2699,N_25613,N_29254);
nand UO_2700 (O_2700,N_28320,N_25697);
xnor UO_2701 (O_2701,N_28573,N_28984);
and UO_2702 (O_2702,N_29536,N_29300);
or UO_2703 (O_2703,N_27346,N_26944);
xnor UO_2704 (O_2704,N_26432,N_29572);
nand UO_2705 (O_2705,N_26678,N_26599);
or UO_2706 (O_2706,N_27730,N_27203);
xor UO_2707 (O_2707,N_29126,N_28091);
and UO_2708 (O_2708,N_28853,N_29394);
and UO_2709 (O_2709,N_27059,N_26633);
and UO_2710 (O_2710,N_26255,N_26668);
nand UO_2711 (O_2711,N_29154,N_27363);
xnor UO_2712 (O_2712,N_26420,N_26648);
nand UO_2713 (O_2713,N_26696,N_28003);
xor UO_2714 (O_2714,N_28870,N_25019);
xnor UO_2715 (O_2715,N_25706,N_25638);
or UO_2716 (O_2716,N_25871,N_29058);
nor UO_2717 (O_2717,N_27660,N_26200);
and UO_2718 (O_2718,N_26425,N_27073);
xnor UO_2719 (O_2719,N_29441,N_29541);
and UO_2720 (O_2720,N_29108,N_25795);
nor UO_2721 (O_2721,N_25171,N_25800);
or UO_2722 (O_2722,N_28852,N_26599);
xnor UO_2723 (O_2723,N_27807,N_28867);
or UO_2724 (O_2724,N_29911,N_27818);
nand UO_2725 (O_2725,N_29593,N_26910);
and UO_2726 (O_2726,N_25901,N_29332);
and UO_2727 (O_2727,N_27025,N_25156);
and UO_2728 (O_2728,N_25532,N_28057);
nand UO_2729 (O_2729,N_28301,N_26646);
or UO_2730 (O_2730,N_29080,N_27276);
and UO_2731 (O_2731,N_29668,N_28449);
xor UO_2732 (O_2732,N_25172,N_27009);
and UO_2733 (O_2733,N_27768,N_25999);
nor UO_2734 (O_2734,N_25495,N_29566);
nor UO_2735 (O_2735,N_29501,N_25502);
nor UO_2736 (O_2736,N_27499,N_29345);
xnor UO_2737 (O_2737,N_29722,N_26962);
nand UO_2738 (O_2738,N_25794,N_28458);
and UO_2739 (O_2739,N_29239,N_25855);
nor UO_2740 (O_2740,N_26834,N_25433);
nand UO_2741 (O_2741,N_28437,N_29062);
and UO_2742 (O_2742,N_28569,N_27383);
nand UO_2743 (O_2743,N_26986,N_26701);
or UO_2744 (O_2744,N_25774,N_29700);
and UO_2745 (O_2745,N_26640,N_29359);
nand UO_2746 (O_2746,N_25788,N_28502);
nor UO_2747 (O_2747,N_29060,N_29661);
or UO_2748 (O_2748,N_29931,N_25379);
nand UO_2749 (O_2749,N_29878,N_26918);
or UO_2750 (O_2750,N_29852,N_29740);
nand UO_2751 (O_2751,N_27623,N_26305);
and UO_2752 (O_2752,N_28285,N_28507);
or UO_2753 (O_2753,N_29322,N_28835);
xnor UO_2754 (O_2754,N_26380,N_28755);
and UO_2755 (O_2755,N_28271,N_29437);
nor UO_2756 (O_2756,N_27223,N_28684);
or UO_2757 (O_2757,N_29447,N_28945);
or UO_2758 (O_2758,N_28567,N_28508);
or UO_2759 (O_2759,N_25628,N_26302);
xor UO_2760 (O_2760,N_29175,N_29724);
nand UO_2761 (O_2761,N_29194,N_27856);
nand UO_2762 (O_2762,N_26026,N_27680);
and UO_2763 (O_2763,N_29552,N_26054);
nor UO_2764 (O_2764,N_27798,N_26335);
nand UO_2765 (O_2765,N_29713,N_29240);
nor UO_2766 (O_2766,N_29289,N_26893);
nor UO_2767 (O_2767,N_29739,N_27225);
xor UO_2768 (O_2768,N_25321,N_27993);
nand UO_2769 (O_2769,N_25746,N_27744);
xor UO_2770 (O_2770,N_28699,N_27392);
nor UO_2771 (O_2771,N_25968,N_29424);
nand UO_2772 (O_2772,N_25459,N_28495);
xnor UO_2773 (O_2773,N_25103,N_27222);
nand UO_2774 (O_2774,N_25531,N_28999);
nor UO_2775 (O_2775,N_29567,N_27676);
or UO_2776 (O_2776,N_29830,N_29465);
and UO_2777 (O_2777,N_28452,N_28489);
nand UO_2778 (O_2778,N_29155,N_28539);
xor UO_2779 (O_2779,N_29567,N_28320);
nor UO_2780 (O_2780,N_26043,N_28836);
and UO_2781 (O_2781,N_28476,N_28939);
nand UO_2782 (O_2782,N_25251,N_27526);
nor UO_2783 (O_2783,N_26685,N_28676);
and UO_2784 (O_2784,N_27654,N_29560);
nand UO_2785 (O_2785,N_25702,N_26220);
or UO_2786 (O_2786,N_28826,N_29273);
and UO_2787 (O_2787,N_26337,N_27238);
xor UO_2788 (O_2788,N_29039,N_28860);
nor UO_2789 (O_2789,N_27451,N_27281);
nand UO_2790 (O_2790,N_28413,N_28007);
nand UO_2791 (O_2791,N_29034,N_29388);
nand UO_2792 (O_2792,N_29806,N_28208);
nor UO_2793 (O_2793,N_27004,N_25546);
nand UO_2794 (O_2794,N_26684,N_27133);
or UO_2795 (O_2795,N_25102,N_28146);
and UO_2796 (O_2796,N_26897,N_27285);
nor UO_2797 (O_2797,N_25494,N_25924);
and UO_2798 (O_2798,N_27067,N_27722);
or UO_2799 (O_2799,N_29903,N_28988);
nand UO_2800 (O_2800,N_25529,N_28876);
nor UO_2801 (O_2801,N_28823,N_27595);
nor UO_2802 (O_2802,N_29962,N_27134);
or UO_2803 (O_2803,N_26249,N_28412);
nand UO_2804 (O_2804,N_29079,N_26093);
or UO_2805 (O_2805,N_25936,N_26070);
nand UO_2806 (O_2806,N_29398,N_26359);
xnor UO_2807 (O_2807,N_28458,N_27625);
and UO_2808 (O_2808,N_25001,N_26374);
xor UO_2809 (O_2809,N_25084,N_29644);
nor UO_2810 (O_2810,N_28863,N_29363);
or UO_2811 (O_2811,N_27527,N_27036);
or UO_2812 (O_2812,N_28452,N_27977);
or UO_2813 (O_2813,N_27025,N_28629);
nor UO_2814 (O_2814,N_25589,N_27809);
xnor UO_2815 (O_2815,N_25054,N_29644);
and UO_2816 (O_2816,N_28230,N_28118);
or UO_2817 (O_2817,N_26744,N_27410);
or UO_2818 (O_2818,N_25128,N_29849);
and UO_2819 (O_2819,N_26437,N_25724);
xor UO_2820 (O_2820,N_26481,N_26626);
and UO_2821 (O_2821,N_29460,N_25460);
nor UO_2822 (O_2822,N_29600,N_25625);
or UO_2823 (O_2823,N_25317,N_25815);
xnor UO_2824 (O_2824,N_25777,N_25614);
nor UO_2825 (O_2825,N_29577,N_29688);
xor UO_2826 (O_2826,N_26923,N_26921);
nand UO_2827 (O_2827,N_25909,N_27098);
nor UO_2828 (O_2828,N_27343,N_29908);
nand UO_2829 (O_2829,N_27827,N_26427);
and UO_2830 (O_2830,N_25496,N_27063);
or UO_2831 (O_2831,N_29620,N_29334);
and UO_2832 (O_2832,N_27231,N_25116);
nand UO_2833 (O_2833,N_25995,N_27983);
xor UO_2834 (O_2834,N_26578,N_27964);
and UO_2835 (O_2835,N_25993,N_27868);
or UO_2836 (O_2836,N_25087,N_29624);
and UO_2837 (O_2837,N_26623,N_28475);
nand UO_2838 (O_2838,N_29408,N_26137);
nand UO_2839 (O_2839,N_27313,N_29208);
or UO_2840 (O_2840,N_27918,N_26333);
and UO_2841 (O_2841,N_26017,N_26907);
nor UO_2842 (O_2842,N_25996,N_28886);
nor UO_2843 (O_2843,N_26577,N_26651);
and UO_2844 (O_2844,N_27805,N_26101);
nand UO_2845 (O_2845,N_29130,N_26394);
xnor UO_2846 (O_2846,N_28595,N_28470);
or UO_2847 (O_2847,N_29581,N_27679);
nand UO_2848 (O_2848,N_26840,N_28294);
and UO_2849 (O_2849,N_29290,N_25675);
and UO_2850 (O_2850,N_26715,N_29573);
or UO_2851 (O_2851,N_25598,N_27652);
and UO_2852 (O_2852,N_27487,N_28540);
xnor UO_2853 (O_2853,N_26968,N_25493);
xnor UO_2854 (O_2854,N_25427,N_25950);
nand UO_2855 (O_2855,N_25093,N_27513);
and UO_2856 (O_2856,N_25084,N_27498);
xor UO_2857 (O_2857,N_26532,N_26462);
or UO_2858 (O_2858,N_25802,N_29539);
nand UO_2859 (O_2859,N_27892,N_26882);
nor UO_2860 (O_2860,N_29002,N_27480);
and UO_2861 (O_2861,N_29891,N_27342);
or UO_2862 (O_2862,N_25058,N_28463);
nor UO_2863 (O_2863,N_26733,N_29476);
nor UO_2864 (O_2864,N_28394,N_28345);
xor UO_2865 (O_2865,N_29806,N_28059);
or UO_2866 (O_2866,N_25212,N_27642);
nand UO_2867 (O_2867,N_26853,N_28011);
nor UO_2868 (O_2868,N_27626,N_28208);
xnor UO_2869 (O_2869,N_29606,N_26466);
nand UO_2870 (O_2870,N_25106,N_28256);
nand UO_2871 (O_2871,N_28385,N_27862);
xnor UO_2872 (O_2872,N_27968,N_26522);
or UO_2873 (O_2873,N_29505,N_29545);
or UO_2874 (O_2874,N_26434,N_28726);
or UO_2875 (O_2875,N_26865,N_26077);
and UO_2876 (O_2876,N_29393,N_25918);
nor UO_2877 (O_2877,N_27050,N_25127);
nand UO_2878 (O_2878,N_29042,N_26507);
nand UO_2879 (O_2879,N_27917,N_25611);
and UO_2880 (O_2880,N_25786,N_27103);
xnor UO_2881 (O_2881,N_29401,N_27212);
nor UO_2882 (O_2882,N_25406,N_29207);
and UO_2883 (O_2883,N_26659,N_28787);
nand UO_2884 (O_2884,N_29636,N_27730);
or UO_2885 (O_2885,N_27655,N_27837);
nand UO_2886 (O_2886,N_25202,N_29387);
xor UO_2887 (O_2887,N_29628,N_27136);
or UO_2888 (O_2888,N_29340,N_25377);
nor UO_2889 (O_2889,N_28037,N_27014);
nand UO_2890 (O_2890,N_27126,N_27035);
or UO_2891 (O_2891,N_28927,N_29107);
nand UO_2892 (O_2892,N_28362,N_28397);
and UO_2893 (O_2893,N_28120,N_27392);
nor UO_2894 (O_2894,N_27792,N_26636);
nand UO_2895 (O_2895,N_25164,N_29900);
xnor UO_2896 (O_2896,N_25399,N_28476);
or UO_2897 (O_2897,N_25260,N_25041);
xor UO_2898 (O_2898,N_27045,N_25281);
xor UO_2899 (O_2899,N_25564,N_28408);
xnor UO_2900 (O_2900,N_29730,N_25397);
nand UO_2901 (O_2901,N_28132,N_29955);
nand UO_2902 (O_2902,N_26461,N_28200);
xor UO_2903 (O_2903,N_28268,N_28707);
xor UO_2904 (O_2904,N_29494,N_26980);
xor UO_2905 (O_2905,N_27921,N_27158);
xnor UO_2906 (O_2906,N_27431,N_28396);
xor UO_2907 (O_2907,N_27617,N_25131);
nor UO_2908 (O_2908,N_26994,N_25097);
and UO_2909 (O_2909,N_26991,N_27650);
nor UO_2910 (O_2910,N_27517,N_26723);
xnor UO_2911 (O_2911,N_29716,N_26553);
nor UO_2912 (O_2912,N_25960,N_25197);
and UO_2913 (O_2913,N_29142,N_25707);
xnor UO_2914 (O_2914,N_25749,N_27949);
or UO_2915 (O_2915,N_28412,N_29467);
or UO_2916 (O_2916,N_28902,N_26944);
nand UO_2917 (O_2917,N_25257,N_28979);
and UO_2918 (O_2918,N_29242,N_29349);
xor UO_2919 (O_2919,N_26739,N_29882);
nor UO_2920 (O_2920,N_29308,N_27304);
nor UO_2921 (O_2921,N_27422,N_25300);
and UO_2922 (O_2922,N_26295,N_29702);
and UO_2923 (O_2923,N_25380,N_28480);
xnor UO_2924 (O_2924,N_29363,N_25430);
or UO_2925 (O_2925,N_28278,N_25818);
or UO_2926 (O_2926,N_25964,N_27962);
and UO_2927 (O_2927,N_26952,N_28339);
and UO_2928 (O_2928,N_29963,N_27758);
nand UO_2929 (O_2929,N_29796,N_28680);
nand UO_2930 (O_2930,N_28571,N_26276);
xnor UO_2931 (O_2931,N_29120,N_26018);
or UO_2932 (O_2932,N_28381,N_28670);
nor UO_2933 (O_2933,N_28407,N_25535);
xnor UO_2934 (O_2934,N_27366,N_27242);
xnor UO_2935 (O_2935,N_25910,N_25706);
nor UO_2936 (O_2936,N_26488,N_25637);
xor UO_2937 (O_2937,N_29528,N_29797);
nor UO_2938 (O_2938,N_28426,N_29925);
xnor UO_2939 (O_2939,N_28177,N_26531);
xnor UO_2940 (O_2940,N_29756,N_28032);
nor UO_2941 (O_2941,N_26173,N_29454);
nand UO_2942 (O_2942,N_25312,N_26928);
and UO_2943 (O_2943,N_26462,N_26591);
nor UO_2944 (O_2944,N_26642,N_27034);
nor UO_2945 (O_2945,N_26988,N_29565);
xor UO_2946 (O_2946,N_29789,N_26434);
nor UO_2947 (O_2947,N_26475,N_26607);
or UO_2948 (O_2948,N_25483,N_29122);
xor UO_2949 (O_2949,N_27245,N_28863);
and UO_2950 (O_2950,N_29498,N_27152);
xnor UO_2951 (O_2951,N_27280,N_29277);
and UO_2952 (O_2952,N_28176,N_27342);
xor UO_2953 (O_2953,N_29213,N_26481);
xnor UO_2954 (O_2954,N_28838,N_26510);
and UO_2955 (O_2955,N_25270,N_29532);
or UO_2956 (O_2956,N_26157,N_25430);
nor UO_2957 (O_2957,N_27236,N_25861);
xnor UO_2958 (O_2958,N_26170,N_27836);
nor UO_2959 (O_2959,N_26006,N_26180);
nor UO_2960 (O_2960,N_26508,N_28459);
nand UO_2961 (O_2961,N_28529,N_27653);
nor UO_2962 (O_2962,N_29947,N_28439);
or UO_2963 (O_2963,N_25881,N_28433);
and UO_2964 (O_2964,N_28851,N_29859);
xnor UO_2965 (O_2965,N_26817,N_25208);
xor UO_2966 (O_2966,N_29847,N_25593);
or UO_2967 (O_2967,N_25255,N_25270);
nand UO_2968 (O_2968,N_27269,N_28992);
or UO_2969 (O_2969,N_25431,N_29891);
nand UO_2970 (O_2970,N_27848,N_29997);
nor UO_2971 (O_2971,N_26695,N_29911);
nand UO_2972 (O_2972,N_28502,N_27565);
nor UO_2973 (O_2973,N_26317,N_26371);
or UO_2974 (O_2974,N_27417,N_27745);
or UO_2975 (O_2975,N_26806,N_25714);
nand UO_2976 (O_2976,N_26416,N_27756);
nor UO_2977 (O_2977,N_26004,N_29318);
nor UO_2978 (O_2978,N_27756,N_28538);
xnor UO_2979 (O_2979,N_25209,N_27809);
or UO_2980 (O_2980,N_25895,N_28948);
nand UO_2981 (O_2981,N_29314,N_28988);
xor UO_2982 (O_2982,N_27191,N_26419);
nor UO_2983 (O_2983,N_26250,N_29202);
or UO_2984 (O_2984,N_28245,N_28698);
nand UO_2985 (O_2985,N_27915,N_29990);
xnor UO_2986 (O_2986,N_29945,N_28024);
nor UO_2987 (O_2987,N_29245,N_29735);
or UO_2988 (O_2988,N_28172,N_29755);
nor UO_2989 (O_2989,N_28519,N_25807);
xnor UO_2990 (O_2990,N_27595,N_25836);
and UO_2991 (O_2991,N_28236,N_25069);
and UO_2992 (O_2992,N_29362,N_28812);
and UO_2993 (O_2993,N_27752,N_29509);
nand UO_2994 (O_2994,N_27596,N_26402);
nand UO_2995 (O_2995,N_29941,N_26034);
xor UO_2996 (O_2996,N_29449,N_29498);
nor UO_2997 (O_2997,N_26568,N_28025);
and UO_2998 (O_2998,N_29594,N_25514);
and UO_2999 (O_2999,N_28784,N_27918);
or UO_3000 (O_3000,N_26140,N_29806);
nand UO_3001 (O_3001,N_25926,N_29107);
xnor UO_3002 (O_3002,N_29869,N_28481);
xnor UO_3003 (O_3003,N_26178,N_27165);
nor UO_3004 (O_3004,N_26671,N_28655);
nor UO_3005 (O_3005,N_26896,N_26391);
and UO_3006 (O_3006,N_25281,N_28070);
or UO_3007 (O_3007,N_27177,N_25803);
or UO_3008 (O_3008,N_27099,N_26293);
or UO_3009 (O_3009,N_25685,N_25724);
xor UO_3010 (O_3010,N_25450,N_26671);
xor UO_3011 (O_3011,N_28123,N_27087);
and UO_3012 (O_3012,N_27110,N_26362);
nand UO_3013 (O_3013,N_25610,N_26668);
and UO_3014 (O_3014,N_27784,N_28681);
and UO_3015 (O_3015,N_29483,N_27399);
or UO_3016 (O_3016,N_29766,N_27146);
and UO_3017 (O_3017,N_27233,N_26466);
nand UO_3018 (O_3018,N_28827,N_26836);
or UO_3019 (O_3019,N_27764,N_25177);
and UO_3020 (O_3020,N_25588,N_26013);
or UO_3021 (O_3021,N_25116,N_27600);
xnor UO_3022 (O_3022,N_26687,N_29290);
or UO_3023 (O_3023,N_27849,N_27369);
and UO_3024 (O_3024,N_25911,N_25971);
or UO_3025 (O_3025,N_28192,N_28513);
xor UO_3026 (O_3026,N_26230,N_28011);
or UO_3027 (O_3027,N_27475,N_26538);
nand UO_3028 (O_3028,N_29502,N_26330);
and UO_3029 (O_3029,N_29399,N_29867);
nor UO_3030 (O_3030,N_28966,N_26879);
nand UO_3031 (O_3031,N_28036,N_29153);
and UO_3032 (O_3032,N_26865,N_29308);
nand UO_3033 (O_3033,N_27143,N_27939);
or UO_3034 (O_3034,N_29714,N_26177);
and UO_3035 (O_3035,N_27631,N_26078);
or UO_3036 (O_3036,N_27866,N_27371);
xor UO_3037 (O_3037,N_29684,N_25735);
or UO_3038 (O_3038,N_25258,N_28201);
nor UO_3039 (O_3039,N_28314,N_28526);
or UO_3040 (O_3040,N_26136,N_29880);
and UO_3041 (O_3041,N_25625,N_25810);
and UO_3042 (O_3042,N_28287,N_27472);
nand UO_3043 (O_3043,N_26485,N_26736);
xor UO_3044 (O_3044,N_29470,N_29746);
nand UO_3045 (O_3045,N_26309,N_25216);
xor UO_3046 (O_3046,N_26131,N_25438);
nand UO_3047 (O_3047,N_27395,N_29574);
xnor UO_3048 (O_3048,N_29709,N_29807);
nand UO_3049 (O_3049,N_26130,N_29924);
nor UO_3050 (O_3050,N_26261,N_29739);
nand UO_3051 (O_3051,N_25046,N_27699);
xnor UO_3052 (O_3052,N_25974,N_28137);
xnor UO_3053 (O_3053,N_29687,N_28731);
nor UO_3054 (O_3054,N_27084,N_27705);
nand UO_3055 (O_3055,N_26084,N_25036);
nand UO_3056 (O_3056,N_29758,N_28266);
nor UO_3057 (O_3057,N_26046,N_25546);
nor UO_3058 (O_3058,N_25432,N_25884);
and UO_3059 (O_3059,N_26683,N_27360);
or UO_3060 (O_3060,N_29916,N_26466);
xor UO_3061 (O_3061,N_25992,N_29412);
or UO_3062 (O_3062,N_29735,N_25048);
and UO_3063 (O_3063,N_29587,N_25144);
nor UO_3064 (O_3064,N_25867,N_29140);
nor UO_3065 (O_3065,N_26581,N_28721);
nor UO_3066 (O_3066,N_28465,N_25648);
or UO_3067 (O_3067,N_29489,N_26492);
or UO_3068 (O_3068,N_26792,N_28435);
or UO_3069 (O_3069,N_29624,N_28658);
xnor UO_3070 (O_3070,N_28315,N_25484);
xor UO_3071 (O_3071,N_27773,N_25437);
nand UO_3072 (O_3072,N_28477,N_29812);
or UO_3073 (O_3073,N_25815,N_27224);
and UO_3074 (O_3074,N_25560,N_28464);
or UO_3075 (O_3075,N_26049,N_27560);
xnor UO_3076 (O_3076,N_26543,N_28854);
nor UO_3077 (O_3077,N_26252,N_25891);
and UO_3078 (O_3078,N_26115,N_25854);
nand UO_3079 (O_3079,N_27779,N_29137);
nand UO_3080 (O_3080,N_28195,N_26012);
xnor UO_3081 (O_3081,N_27088,N_28065);
nor UO_3082 (O_3082,N_28333,N_26864);
xnor UO_3083 (O_3083,N_27275,N_26810);
nand UO_3084 (O_3084,N_28277,N_25139);
nand UO_3085 (O_3085,N_28091,N_28679);
xor UO_3086 (O_3086,N_25033,N_26382);
and UO_3087 (O_3087,N_27144,N_25288);
nor UO_3088 (O_3088,N_29836,N_25062);
nor UO_3089 (O_3089,N_28469,N_26153);
nor UO_3090 (O_3090,N_26231,N_28359);
xor UO_3091 (O_3091,N_26321,N_26230);
or UO_3092 (O_3092,N_29349,N_29789);
and UO_3093 (O_3093,N_28407,N_28480);
nor UO_3094 (O_3094,N_29210,N_29525);
and UO_3095 (O_3095,N_26180,N_29520);
and UO_3096 (O_3096,N_27371,N_25026);
xor UO_3097 (O_3097,N_29051,N_28271);
nand UO_3098 (O_3098,N_25649,N_28442);
nand UO_3099 (O_3099,N_28306,N_27479);
nor UO_3100 (O_3100,N_25451,N_29617);
or UO_3101 (O_3101,N_26771,N_26102);
nand UO_3102 (O_3102,N_29317,N_27855);
nand UO_3103 (O_3103,N_25035,N_26921);
nand UO_3104 (O_3104,N_26738,N_29456);
or UO_3105 (O_3105,N_28064,N_28231);
nand UO_3106 (O_3106,N_25518,N_28708);
nor UO_3107 (O_3107,N_29909,N_25038);
nand UO_3108 (O_3108,N_27447,N_25326);
nor UO_3109 (O_3109,N_29769,N_29405);
xor UO_3110 (O_3110,N_25598,N_26512);
xor UO_3111 (O_3111,N_29735,N_25822);
and UO_3112 (O_3112,N_27930,N_27667);
or UO_3113 (O_3113,N_26384,N_27190);
nor UO_3114 (O_3114,N_25536,N_29660);
and UO_3115 (O_3115,N_25663,N_27349);
and UO_3116 (O_3116,N_29915,N_26071);
and UO_3117 (O_3117,N_26430,N_29814);
xor UO_3118 (O_3118,N_25217,N_26157);
nor UO_3119 (O_3119,N_27291,N_25028);
nor UO_3120 (O_3120,N_26729,N_28979);
and UO_3121 (O_3121,N_25322,N_26726);
or UO_3122 (O_3122,N_29952,N_29846);
and UO_3123 (O_3123,N_28080,N_27994);
nand UO_3124 (O_3124,N_25996,N_25349);
xnor UO_3125 (O_3125,N_26837,N_25861);
or UO_3126 (O_3126,N_26687,N_28369);
nor UO_3127 (O_3127,N_29501,N_25955);
xnor UO_3128 (O_3128,N_29986,N_27623);
nand UO_3129 (O_3129,N_26093,N_27692);
or UO_3130 (O_3130,N_25880,N_27730);
nor UO_3131 (O_3131,N_26262,N_26635);
nand UO_3132 (O_3132,N_28928,N_28651);
xor UO_3133 (O_3133,N_26139,N_27110);
nand UO_3134 (O_3134,N_29715,N_25087);
and UO_3135 (O_3135,N_27219,N_25387);
and UO_3136 (O_3136,N_28490,N_26877);
or UO_3137 (O_3137,N_27708,N_27873);
xor UO_3138 (O_3138,N_28654,N_25134);
nand UO_3139 (O_3139,N_25867,N_25219);
xor UO_3140 (O_3140,N_27514,N_28128);
nor UO_3141 (O_3141,N_28400,N_26995);
xnor UO_3142 (O_3142,N_27228,N_25849);
nor UO_3143 (O_3143,N_28402,N_27209);
nand UO_3144 (O_3144,N_28170,N_28590);
or UO_3145 (O_3145,N_27283,N_27113);
xnor UO_3146 (O_3146,N_28535,N_28458);
nor UO_3147 (O_3147,N_26053,N_28269);
nor UO_3148 (O_3148,N_26070,N_28337);
or UO_3149 (O_3149,N_26600,N_26843);
or UO_3150 (O_3150,N_26088,N_26738);
or UO_3151 (O_3151,N_28331,N_27563);
nand UO_3152 (O_3152,N_27142,N_29136);
and UO_3153 (O_3153,N_26948,N_29472);
xor UO_3154 (O_3154,N_26789,N_29640);
and UO_3155 (O_3155,N_27954,N_27622);
xor UO_3156 (O_3156,N_28357,N_25550);
xnor UO_3157 (O_3157,N_26782,N_29755);
xnor UO_3158 (O_3158,N_26430,N_25396);
nand UO_3159 (O_3159,N_28521,N_27103);
xnor UO_3160 (O_3160,N_28378,N_27906);
or UO_3161 (O_3161,N_26957,N_25793);
and UO_3162 (O_3162,N_28536,N_25798);
and UO_3163 (O_3163,N_28819,N_27290);
or UO_3164 (O_3164,N_26792,N_27074);
and UO_3165 (O_3165,N_27507,N_27581);
nand UO_3166 (O_3166,N_26807,N_29544);
nor UO_3167 (O_3167,N_26799,N_29936);
and UO_3168 (O_3168,N_26227,N_29598);
nand UO_3169 (O_3169,N_29373,N_26726);
nand UO_3170 (O_3170,N_25440,N_28388);
nor UO_3171 (O_3171,N_28524,N_27042);
nand UO_3172 (O_3172,N_25056,N_25349);
or UO_3173 (O_3173,N_28709,N_27431);
and UO_3174 (O_3174,N_25082,N_28430);
xor UO_3175 (O_3175,N_29016,N_29258);
or UO_3176 (O_3176,N_26936,N_25873);
and UO_3177 (O_3177,N_27642,N_25178);
nor UO_3178 (O_3178,N_29993,N_29232);
xnor UO_3179 (O_3179,N_27912,N_27330);
nand UO_3180 (O_3180,N_28370,N_29953);
nand UO_3181 (O_3181,N_29108,N_29513);
nor UO_3182 (O_3182,N_29643,N_29473);
and UO_3183 (O_3183,N_27388,N_27521);
nor UO_3184 (O_3184,N_26039,N_28711);
nand UO_3185 (O_3185,N_26900,N_28930);
or UO_3186 (O_3186,N_29570,N_25858);
or UO_3187 (O_3187,N_26222,N_25694);
nor UO_3188 (O_3188,N_28520,N_26824);
xor UO_3189 (O_3189,N_27872,N_28566);
or UO_3190 (O_3190,N_28391,N_29477);
nand UO_3191 (O_3191,N_26972,N_26927);
nor UO_3192 (O_3192,N_29257,N_28926);
nand UO_3193 (O_3193,N_28412,N_26132);
nand UO_3194 (O_3194,N_29012,N_27794);
xor UO_3195 (O_3195,N_27455,N_26243);
nand UO_3196 (O_3196,N_29407,N_25697);
nand UO_3197 (O_3197,N_27151,N_26604);
nand UO_3198 (O_3198,N_25210,N_26326);
nand UO_3199 (O_3199,N_25575,N_29159);
or UO_3200 (O_3200,N_29685,N_28871);
or UO_3201 (O_3201,N_29813,N_26515);
nor UO_3202 (O_3202,N_26010,N_27536);
nor UO_3203 (O_3203,N_26598,N_27053);
xor UO_3204 (O_3204,N_29056,N_27883);
nand UO_3205 (O_3205,N_25241,N_27697);
xnor UO_3206 (O_3206,N_28170,N_26794);
or UO_3207 (O_3207,N_25375,N_27410);
nand UO_3208 (O_3208,N_27098,N_27720);
nor UO_3209 (O_3209,N_26322,N_25893);
or UO_3210 (O_3210,N_25789,N_26340);
nor UO_3211 (O_3211,N_28938,N_26344);
and UO_3212 (O_3212,N_28104,N_28102);
or UO_3213 (O_3213,N_27361,N_29010);
nor UO_3214 (O_3214,N_28533,N_29934);
and UO_3215 (O_3215,N_26808,N_28833);
nor UO_3216 (O_3216,N_29945,N_28061);
nand UO_3217 (O_3217,N_29228,N_29770);
xor UO_3218 (O_3218,N_27513,N_25424);
nand UO_3219 (O_3219,N_28515,N_26436);
and UO_3220 (O_3220,N_27100,N_26265);
nand UO_3221 (O_3221,N_28480,N_29017);
or UO_3222 (O_3222,N_29329,N_28543);
nor UO_3223 (O_3223,N_25409,N_27809);
and UO_3224 (O_3224,N_26846,N_26235);
and UO_3225 (O_3225,N_28284,N_26414);
or UO_3226 (O_3226,N_25627,N_26475);
and UO_3227 (O_3227,N_28883,N_25488);
nand UO_3228 (O_3228,N_29188,N_28849);
nand UO_3229 (O_3229,N_25823,N_27680);
nand UO_3230 (O_3230,N_26684,N_27646);
nor UO_3231 (O_3231,N_29413,N_28889);
or UO_3232 (O_3232,N_28387,N_27859);
nor UO_3233 (O_3233,N_27734,N_29102);
nand UO_3234 (O_3234,N_27172,N_28387);
nor UO_3235 (O_3235,N_29931,N_26553);
and UO_3236 (O_3236,N_27609,N_26378);
and UO_3237 (O_3237,N_25197,N_27262);
nand UO_3238 (O_3238,N_27234,N_29752);
nor UO_3239 (O_3239,N_25547,N_27612);
xnor UO_3240 (O_3240,N_26296,N_27287);
or UO_3241 (O_3241,N_29069,N_28764);
xor UO_3242 (O_3242,N_27681,N_27805);
and UO_3243 (O_3243,N_26576,N_28679);
nor UO_3244 (O_3244,N_27738,N_27275);
nand UO_3245 (O_3245,N_25390,N_26498);
xnor UO_3246 (O_3246,N_25827,N_29465);
xnor UO_3247 (O_3247,N_28654,N_28276);
nand UO_3248 (O_3248,N_26036,N_26405);
and UO_3249 (O_3249,N_27396,N_25628);
or UO_3250 (O_3250,N_28676,N_25115);
xnor UO_3251 (O_3251,N_25444,N_27144);
and UO_3252 (O_3252,N_27375,N_26210);
nand UO_3253 (O_3253,N_26147,N_26528);
nand UO_3254 (O_3254,N_27892,N_29881);
xor UO_3255 (O_3255,N_27254,N_25235);
nor UO_3256 (O_3256,N_29381,N_26853);
xnor UO_3257 (O_3257,N_27520,N_25257);
or UO_3258 (O_3258,N_25663,N_28563);
and UO_3259 (O_3259,N_28277,N_29974);
nand UO_3260 (O_3260,N_27760,N_27528);
nand UO_3261 (O_3261,N_27765,N_27638);
xnor UO_3262 (O_3262,N_28277,N_27828);
or UO_3263 (O_3263,N_27221,N_29261);
nor UO_3264 (O_3264,N_25713,N_26587);
or UO_3265 (O_3265,N_26796,N_25485);
or UO_3266 (O_3266,N_28803,N_27315);
xor UO_3267 (O_3267,N_28375,N_29250);
nand UO_3268 (O_3268,N_25438,N_29004);
xor UO_3269 (O_3269,N_25623,N_29755);
or UO_3270 (O_3270,N_27251,N_25848);
or UO_3271 (O_3271,N_28765,N_28845);
xor UO_3272 (O_3272,N_28333,N_29890);
and UO_3273 (O_3273,N_25681,N_28118);
nand UO_3274 (O_3274,N_29899,N_27906);
nand UO_3275 (O_3275,N_26679,N_29052);
xor UO_3276 (O_3276,N_25078,N_27548);
and UO_3277 (O_3277,N_25473,N_27096);
and UO_3278 (O_3278,N_29572,N_26648);
nand UO_3279 (O_3279,N_29204,N_26746);
nand UO_3280 (O_3280,N_28683,N_27311);
and UO_3281 (O_3281,N_26236,N_29012);
xnor UO_3282 (O_3282,N_25508,N_27589);
nor UO_3283 (O_3283,N_28646,N_27718);
or UO_3284 (O_3284,N_25690,N_28326);
nor UO_3285 (O_3285,N_29632,N_28921);
xor UO_3286 (O_3286,N_29790,N_25213);
nand UO_3287 (O_3287,N_29051,N_26967);
nand UO_3288 (O_3288,N_28785,N_29854);
xor UO_3289 (O_3289,N_25186,N_29599);
nand UO_3290 (O_3290,N_27974,N_27236);
xor UO_3291 (O_3291,N_28994,N_25115);
nand UO_3292 (O_3292,N_27880,N_28322);
or UO_3293 (O_3293,N_26195,N_26729);
nand UO_3294 (O_3294,N_27358,N_29885);
and UO_3295 (O_3295,N_29263,N_28500);
nand UO_3296 (O_3296,N_25412,N_28079);
nand UO_3297 (O_3297,N_26951,N_26729);
and UO_3298 (O_3298,N_29336,N_25348);
nand UO_3299 (O_3299,N_28701,N_25345);
and UO_3300 (O_3300,N_29236,N_26589);
and UO_3301 (O_3301,N_26432,N_29319);
xor UO_3302 (O_3302,N_26364,N_28603);
or UO_3303 (O_3303,N_29843,N_28881);
nand UO_3304 (O_3304,N_28685,N_26772);
nor UO_3305 (O_3305,N_25377,N_26253);
xnor UO_3306 (O_3306,N_27914,N_26770);
nor UO_3307 (O_3307,N_29552,N_29192);
nand UO_3308 (O_3308,N_26283,N_25256);
or UO_3309 (O_3309,N_29811,N_28049);
xor UO_3310 (O_3310,N_29572,N_29127);
nor UO_3311 (O_3311,N_27331,N_26023);
xor UO_3312 (O_3312,N_29019,N_27708);
or UO_3313 (O_3313,N_29953,N_29058);
nor UO_3314 (O_3314,N_25689,N_25342);
and UO_3315 (O_3315,N_29026,N_25696);
and UO_3316 (O_3316,N_25925,N_29659);
and UO_3317 (O_3317,N_29815,N_26481);
or UO_3318 (O_3318,N_29295,N_27274);
nand UO_3319 (O_3319,N_26671,N_29500);
nand UO_3320 (O_3320,N_28177,N_26951);
or UO_3321 (O_3321,N_28797,N_26822);
nand UO_3322 (O_3322,N_29539,N_28642);
or UO_3323 (O_3323,N_25750,N_29953);
and UO_3324 (O_3324,N_25273,N_29007);
nor UO_3325 (O_3325,N_25596,N_26582);
and UO_3326 (O_3326,N_26514,N_29916);
xnor UO_3327 (O_3327,N_27013,N_28098);
nand UO_3328 (O_3328,N_25541,N_26431);
or UO_3329 (O_3329,N_26685,N_26899);
nor UO_3330 (O_3330,N_29755,N_27917);
nand UO_3331 (O_3331,N_26592,N_26620);
and UO_3332 (O_3332,N_28206,N_27873);
or UO_3333 (O_3333,N_25894,N_25717);
xor UO_3334 (O_3334,N_29850,N_29258);
nand UO_3335 (O_3335,N_25256,N_26112);
and UO_3336 (O_3336,N_26365,N_28275);
or UO_3337 (O_3337,N_26821,N_26510);
nor UO_3338 (O_3338,N_27640,N_28321);
and UO_3339 (O_3339,N_26974,N_25964);
and UO_3340 (O_3340,N_26388,N_25444);
nor UO_3341 (O_3341,N_26224,N_27249);
nand UO_3342 (O_3342,N_25972,N_28047);
xor UO_3343 (O_3343,N_25242,N_26317);
and UO_3344 (O_3344,N_28515,N_26561);
nor UO_3345 (O_3345,N_27946,N_29704);
nand UO_3346 (O_3346,N_27655,N_26059);
or UO_3347 (O_3347,N_26157,N_28623);
or UO_3348 (O_3348,N_28684,N_25716);
nand UO_3349 (O_3349,N_29502,N_26679);
or UO_3350 (O_3350,N_25424,N_25678);
nor UO_3351 (O_3351,N_28651,N_25281);
xor UO_3352 (O_3352,N_25147,N_29792);
xnor UO_3353 (O_3353,N_25853,N_28388);
xnor UO_3354 (O_3354,N_29784,N_25019);
nor UO_3355 (O_3355,N_29226,N_29441);
xor UO_3356 (O_3356,N_25347,N_29009);
and UO_3357 (O_3357,N_29457,N_28631);
nor UO_3358 (O_3358,N_27496,N_25477);
or UO_3359 (O_3359,N_25362,N_28209);
nor UO_3360 (O_3360,N_29650,N_29501);
nor UO_3361 (O_3361,N_25363,N_28230);
or UO_3362 (O_3362,N_27508,N_27680);
or UO_3363 (O_3363,N_29054,N_27793);
or UO_3364 (O_3364,N_27413,N_27877);
xor UO_3365 (O_3365,N_25216,N_25113);
nor UO_3366 (O_3366,N_29996,N_26570);
and UO_3367 (O_3367,N_25719,N_29938);
or UO_3368 (O_3368,N_28708,N_25379);
nand UO_3369 (O_3369,N_27858,N_26500);
or UO_3370 (O_3370,N_26309,N_27372);
and UO_3371 (O_3371,N_26180,N_27898);
nor UO_3372 (O_3372,N_28774,N_29389);
or UO_3373 (O_3373,N_25810,N_26661);
xnor UO_3374 (O_3374,N_25081,N_26988);
xnor UO_3375 (O_3375,N_28731,N_27274);
or UO_3376 (O_3376,N_28548,N_27828);
and UO_3377 (O_3377,N_26283,N_27051);
and UO_3378 (O_3378,N_25416,N_28171);
xor UO_3379 (O_3379,N_26191,N_29562);
nor UO_3380 (O_3380,N_26463,N_25958);
nand UO_3381 (O_3381,N_26375,N_28505);
and UO_3382 (O_3382,N_25499,N_25468);
nand UO_3383 (O_3383,N_28467,N_27786);
nand UO_3384 (O_3384,N_28333,N_25038);
nand UO_3385 (O_3385,N_28049,N_29459);
and UO_3386 (O_3386,N_25278,N_29012);
nor UO_3387 (O_3387,N_28090,N_26401);
xor UO_3388 (O_3388,N_25966,N_29206);
or UO_3389 (O_3389,N_28407,N_29211);
and UO_3390 (O_3390,N_25960,N_27813);
or UO_3391 (O_3391,N_29627,N_25770);
nand UO_3392 (O_3392,N_27227,N_27451);
xnor UO_3393 (O_3393,N_27222,N_29202);
and UO_3394 (O_3394,N_26767,N_26136);
nor UO_3395 (O_3395,N_27780,N_28741);
xor UO_3396 (O_3396,N_26252,N_28773);
or UO_3397 (O_3397,N_27689,N_27814);
or UO_3398 (O_3398,N_26893,N_25414);
and UO_3399 (O_3399,N_28504,N_25274);
xor UO_3400 (O_3400,N_27486,N_26362);
xor UO_3401 (O_3401,N_26439,N_28603);
xnor UO_3402 (O_3402,N_27968,N_28706);
xor UO_3403 (O_3403,N_27877,N_28294);
xnor UO_3404 (O_3404,N_27858,N_25667);
xor UO_3405 (O_3405,N_26974,N_29989);
nor UO_3406 (O_3406,N_28763,N_29073);
and UO_3407 (O_3407,N_28046,N_28301);
and UO_3408 (O_3408,N_26716,N_25557);
and UO_3409 (O_3409,N_29235,N_27239);
nor UO_3410 (O_3410,N_25105,N_29189);
nand UO_3411 (O_3411,N_25385,N_26135);
and UO_3412 (O_3412,N_26284,N_26024);
nand UO_3413 (O_3413,N_29927,N_26598);
or UO_3414 (O_3414,N_27129,N_25551);
nor UO_3415 (O_3415,N_25986,N_28360);
nor UO_3416 (O_3416,N_27878,N_27674);
xor UO_3417 (O_3417,N_28549,N_27936);
nand UO_3418 (O_3418,N_26224,N_27114);
and UO_3419 (O_3419,N_29554,N_27954);
nor UO_3420 (O_3420,N_29201,N_29355);
and UO_3421 (O_3421,N_28500,N_25532);
nor UO_3422 (O_3422,N_27181,N_26229);
nand UO_3423 (O_3423,N_27482,N_26113);
or UO_3424 (O_3424,N_26676,N_28422);
xor UO_3425 (O_3425,N_29513,N_27545);
or UO_3426 (O_3426,N_29579,N_26963);
nand UO_3427 (O_3427,N_28102,N_29568);
and UO_3428 (O_3428,N_28537,N_28039);
nand UO_3429 (O_3429,N_26483,N_26120);
and UO_3430 (O_3430,N_28377,N_29673);
nor UO_3431 (O_3431,N_28504,N_28438);
or UO_3432 (O_3432,N_29719,N_27671);
or UO_3433 (O_3433,N_27346,N_27158);
and UO_3434 (O_3434,N_25695,N_28889);
xor UO_3435 (O_3435,N_29623,N_29642);
or UO_3436 (O_3436,N_25513,N_28210);
nand UO_3437 (O_3437,N_28362,N_28327);
nand UO_3438 (O_3438,N_28536,N_27414);
nor UO_3439 (O_3439,N_27338,N_28184);
nand UO_3440 (O_3440,N_29294,N_26141);
nor UO_3441 (O_3441,N_28756,N_29474);
nand UO_3442 (O_3442,N_26661,N_27329);
and UO_3443 (O_3443,N_26469,N_29809);
nor UO_3444 (O_3444,N_28516,N_28699);
and UO_3445 (O_3445,N_27475,N_26679);
xnor UO_3446 (O_3446,N_27360,N_27283);
and UO_3447 (O_3447,N_29472,N_29573);
or UO_3448 (O_3448,N_25476,N_28262);
nor UO_3449 (O_3449,N_27005,N_28641);
and UO_3450 (O_3450,N_25344,N_26478);
nor UO_3451 (O_3451,N_29825,N_26176);
and UO_3452 (O_3452,N_25903,N_26047);
or UO_3453 (O_3453,N_28011,N_26007);
nand UO_3454 (O_3454,N_28064,N_26700);
nand UO_3455 (O_3455,N_28616,N_27643);
nor UO_3456 (O_3456,N_27084,N_29239);
nand UO_3457 (O_3457,N_29778,N_29962);
nor UO_3458 (O_3458,N_25953,N_27385);
and UO_3459 (O_3459,N_26731,N_27430);
and UO_3460 (O_3460,N_26784,N_26780);
and UO_3461 (O_3461,N_28103,N_26183);
or UO_3462 (O_3462,N_26315,N_25651);
nand UO_3463 (O_3463,N_28616,N_28207);
and UO_3464 (O_3464,N_29064,N_28091);
xor UO_3465 (O_3465,N_27910,N_28923);
nand UO_3466 (O_3466,N_28001,N_29002);
xnor UO_3467 (O_3467,N_26956,N_29015);
or UO_3468 (O_3468,N_28382,N_26214);
xnor UO_3469 (O_3469,N_27521,N_27335);
and UO_3470 (O_3470,N_26496,N_28688);
or UO_3471 (O_3471,N_25814,N_26658);
and UO_3472 (O_3472,N_26030,N_26377);
xnor UO_3473 (O_3473,N_29912,N_28305);
xor UO_3474 (O_3474,N_27198,N_29922);
nand UO_3475 (O_3475,N_26141,N_25209);
nand UO_3476 (O_3476,N_27076,N_28947);
and UO_3477 (O_3477,N_26961,N_28850);
and UO_3478 (O_3478,N_26633,N_25160);
nor UO_3479 (O_3479,N_29432,N_27413);
nand UO_3480 (O_3480,N_25727,N_25225);
nand UO_3481 (O_3481,N_29951,N_29425);
nor UO_3482 (O_3482,N_29609,N_29687);
xor UO_3483 (O_3483,N_27967,N_28090);
xor UO_3484 (O_3484,N_27157,N_29461);
and UO_3485 (O_3485,N_27393,N_29303);
nand UO_3486 (O_3486,N_27479,N_26320);
or UO_3487 (O_3487,N_25547,N_27147);
nor UO_3488 (O_3488,N_28349,N_26240);
or UO_3489 (O_3489,N_27543,N_27072);
nand UO_3490 (O_3490,N_28539,N_28524);
nand UO_3491 (O_3491,N_27539,N_25158);
or UO_3492 (O_3492,N_26862,N_27489);
xnor UO_3493 (O_3493,N_29993,N_28424);
or UO_3494 (O_3494,N_29743,N_28344);
xor UO_3495 (O_3495,N_26923,N_27145);
and UO_3496 (O_3496,N_29148,N_26790);
or UO_3497 (O_3497,N_29978,N_25869);
or UO_3498 (O_3498,N_29973,N_25904);
nor UO_3499 (O_3499,N_25693,N_29142);
endmodule