module basic_1000_10000_1500_10_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_270,In_935);
and U1 (N_1,In_622,In_415);
xnor U2 (N_2,In_90,In_842);
or U3 (N_3,In_604,In_649);
nor U4 (N_4,In_891,In_992);
nand U5 (N_5,In_541,In_943);
and U6 (N_6,In_662,In_688);
or U7 (N_7,In_754,In_776);
and U8 (N_8,In_819,In_998);
nand U9 (N_9,In_826,In_99);
nor U10 (N_10,In_860,In_446);
nor U11 (N_11,In_534,In_200);
nand U12 (N_12,In_879,In_613);
or U13 (N_13,In_997,In_991);
and U14 (N_14,In_75,In_671);
or U15 (N_15,In_91,In_118);
or U16 (N_16,In_920,In_564);
nor U17 (N_17,In_193,In_761);
nor U18 (N_18,In_885,In_771);
nor U19 (N_19,In_650,In_570);
and U20 (N_20,In_692,In_971);
or U21 (N_21,In_938,In_871);
and U22 (N_22,In_146,In_31);
and U23 (N_23,In_503,In_52);
nor U24 (N_24,In_736,In_957);
nand U25 (N_25,In_184,In_724);
nor U26 (N_26,In_419,In_80);
and U27 (N_27,In_71,In_441);
and U28 (N_28,In_960,In_257);
and U29 (N_29,In_693,In_51);
nand U30 (N_30,In_939,In_358);
nand U31 (N_31,In_332,In_827);
nand U32 (N_32,In_985,In_634);
nor U33 (N_33,In_691,In_142);
nor U34 (N_34,In_195,In_492);
nor U35 (N_35,In_896,In_149);
nor U36 (N_36,In_866,In_449);
and U37 (N_37,In_235,In_422);
and U38 (N_38,In_134,In_460);
and U39 (N_39,In_489,In_473);
nand U40 (N_40,In_224,In_397);
nand U41 (N_41,In_966,In_1);
and U42 (N_42,In_493,In_379);
or U43 (N_43,In_350,In_354);
or U44 (N_44,In_97,In_309);
nor U45 (N_45,In_181,In_645);
xnor U46 (N_46,In_176,In_208);
nor U47 (N_47,In_294,In_221);
nor U48 (N_48,In_57,In_199);
nor U49 (N_49,In_814,In_426);
and U50 (N_50,In_642,In_108);
or U51 (N_51,In_417,In_868);
and U52 (N_52,In_687,In_924);
nand U53 (N_53,In_73,In_822);
nand U54 (N_54,In_403,In_793);
and U55 (N_55,In_166,In_324);
and U56 (N_56,In_796,In_88);
nor U57 (N_57,In_631,In_274);
and U58 (N_58,In_690,In_594);
nand U59 (N_59,In_467,In_735);
and U60 (N_60,In_777,In_204);
or U61 (N_61,In_383,In_949);
nand U62 (N_62,In_770,In_303);
nor U63 (N_63,In_722,In_584);
or U64 (N_64,In_798,In_404);
or U65 (N_65,In_187,In_188);
nor U66 (N_66,In_501,In_3);
or U67 (N_67,In_664,In_384);
or U68 (N_68,In_268,In_792);
and U69 (N_69,In_869,In_472);
nor U70 (N_70,In_53,In_569);
or U71 (N_71,In_875,In_563);
and U72 (N_72,In_86,In_699);
nor U73 (N_73,In_409,In_810);
and U74 (N_74,In_277,In_716);
nor U75 (N_75,In_136,In_767);
nor U76 (N_76,In_157,In_6);
nand U77 (N_77,In_256,In_505);
xnor U78 (N_78,In_946,In_447);
nor U79 (N_79,In_682,In_972);
or U80 (N_80,In_8,In_261);
or U81 (N_81,In_228,In_612);
nand U82 (N_82,In_683,In_729);
nand U83 (N_83,In_273,In_525);
xnor U84 (N_84,In_704,In_260);
nor U85 (N_85,In_910,In_956);
nor U86 (N_86,In_799,In_583);
or U87 (N_87,In_129,In_490);
nand U88 (N_88,In_881,In_849);
and U89 (N_89,In_22,In_476);
and U90 (N_90,In_837,In_829);
and U91 (N_91,In_929,In_848);
and U92 (N_92,In_605,In_194);
nor U93 (N_93,In_341,In_661);
nor U94 (N_94,In_5,In_844);
and U95 (N_95,In_406,In_281);
or U96 (N_96,In_524,In_74);
or U97 (N_97,In_428,In_934);
nand U98 (N_98,In_655,In_601);
nor U99 (N_99,In_918,In_70);
and U100 (N_100,In_227,In_701);
nor U101 (N_101,In_271,In_486);
nand U102 (N_102,In_387,In_615);
nor U103 (N_103,In_940,In_122);
or U104 (N_104,In_82,In_515);
or U105 (N_105,In_626,In_775);
nor U106 (N_106,In_909,In_343);
or U107 (N_107,In_393,In_470);
nand U108 (N_108,In_301,In_313);
or U109 (N_109,In_630,In_319);
or U110 (N_110,In_340,In_161);
or U111 (N_111,In_49,In_894);
nor U112 (N_112,In_215,In_2);
nor U113 (N_113,In_884,In_41);
and U114 (N_114,In_714,In_171);
nor U115 (N_115,In_272,In_100);
or U116 (N_116,In_368,In_300);
nand U117 (N_117,In_201,In_238);
and U118 (N_118,In_405,In_61);
nand U119 (N_119,In_533,In_255);
and U120 (N_120,In_400,In_527);
nand U121 (N_121,In_648,In_247);
or U122 (N_122,In_308,In_592);
nand U123 (N_123,In_835,In_903);
and U124 (N_124,In_652,In_180);
and U125 (N_125,In_321,In_932);
nor U126 (N_126,In_820,In_876);
nand U127 (N_127,In_115,In_382);
nand U128 (N_128,In_755,In_568);
and U129 (N_129,In_520,In_902);
and U130 (N_130,In_590,In_953);
nor U131 (N_131,In_958,In_922);
nand U132 (N_132,In_380,In_983);
or U133 (N_133,In_596,In_475);
and U134 (N_134,In_111,In_65);
and U135 (N_135,In_951,In_213);
and U136 (N_136,In_591,In_32);
nand U137 (N_137,In_870,In_504);
and U138 (N_138,In_514,In_617);
or U139 (N_139,In_899,In_364);
nand U140 (N_140,In_55,In_192);
nand U141 (N_141,In_289,In_401);
or U142 (N_142,In_474,In_721);
nand U143 (N_143,In_363,In_167);
nand U144 (N_144,In_346,In_252);
nor U145 (N_145,In_865,In_571);
or U146 (N_146,In_597,In_141);
nor U147 (N_147,In_17,In_128);
nand U148 (N_148,In_395,In_450);
nand U149 (N_149,In_600,In_12);
nand U150 (N_150,In_962,In_995);
and U151 (N_151,In_984,In_703);
nand U152 (N_152,In_542,In_937);
nor U153 (N_153,In_39,In_312);
and U154 (N_154,In_185,In_680);
or U155 (N_155,In_314,In_916);
nand U156 (N_156,In_190,In_68);
and U157 (N_157,In_954,In_496);
nand U158 (N_158,In_981,In_518);
and U159 (N_159,In_310,In_381);
nor U160 (N_160,In_242,In_811);
or U161 (N_161,In_707,In_970);
nand U162 (N_162,In_732,In_582);
and U163 (N_163,In_912,In_521);
nand U164 (N_164,In_36,In_152);
and U165 (N_165,In_355,In_500);
or U166 (N_166,In_429,In_34);
nor U167 (N_167,In_926,In_338);
nor U168 (N_168,In_548,In_240);
nor U169 (N_169,In_751,In_480);
nand U170 (N_170,In_170,In_697);
nor U171 (N_171,In_280,In_616);
nor U172 (N_172,In_538,In_366);
and U173 (N_173,In_567,In_788);
and U174 (N_174,In_673,In_126);
or U175 (N_175,In_580,In_156);
nand U176 (N_176,In_928,In_336);
and U177 (N_177,In_132,In_353);
and U178 (N_178,In_745,In_702);
nor U179 (N_179,In_435,In_378);
nor U180 (N_180,In_620,In_110);
or U181 (N_181,In_425,In_197);
or U182 (N_182,In_494,In_24);
and U183 (N_183,In_765,In_320);
and U184 (N_184,In_973,In_396);
or U185 (N_185,In_809,In_431);
or U186 (N_186,In_11,In_974);
and U187 (N_187,In_328,In_807);
nor U188 (N_188,In_365,In_887);
or U189 (N_189,In_511,In_952);
and U190 (N_190,In_20,In_16);
nor U191 (N_191,In_667,In_69);
nand U192 (N_192,In_644,In_98);
nand U193 (N_193,In_479,In_506);
or U194 (N_194,In_588,In_81);
nor U195 (N_195,In_394,In_677);
nor U196 (N_196,In_84,In_519);
and U197 (N_197,In_163,In_333);
or U198 (N_198,In_746,In_442);
nor U199 (N_199,In_219,In_815);
nand U200 (N_200,In_672,In_639);
and U201 (N_201,In_824,In_674);
nor U202 (N_202,In_982,In_609);
nor U203 (N_203,In_357,In_174);
or U204 (N_204,In_877,In_857);
and U205 (N_205,In_237,In_517);
nand U206 (N_206,In_230,In_436);
nand U207 (N_207,In_941,In_434);
and U208 (N_208,In_818,In_968);
and U209 (N_209,In_959,In_444);
or U210 (N_210,In_539,In_742);
nand U211 (N_211,In_558,In_872);
nor U212 (N_212,In_63,In_205);
nor U213 (N_213,In_112,In_990);
or U214 (N_214,In_48,In_172);
nand U215 (N_215,In_522,In_689);
or U216 (N_216,In_102,In_978);
xnor U217 (N_217,In_318,In_882);
xnor U218 (N_218,In_169,In_483);
and U219 (N_219,In_821,In_706);
nand U220 (N_220,In_298,In_653);
xor U221 (N_221,In_345,In_220);
or U222 (N_222,In_456,In_577);
or U223 (N_223,In_113,In_635);
xor U224 (N_224,In_813,In_606);
nand U225 (N_225,In_440,In_585);
nand U226 (N_226,In_787,In_627);
nand U227 (N_227,In_684,In_445);
and U228 (N_228,In_944,In_131);
nor U229 (N_229,In_150,In_737);
nand U230 (N_230,In_337,In_963);
and U231 (N_231,In_402,In_399);
and U232 (N_232,In_443,In_930);
nand U233 (N_233,In_840,In_833);
nor U234 (N_234,In_715,In_720);
nor U235 (N_235,In_743,In_608);
xor U236 (N_236,In_651,In_694);
nor U237 (N_237,In_209,In_351);
or U238 (N_238,In_484,In_727);
nand U239 (N_239,In_532,In_372);
or U240 (N_240,In_549,In_222);
nor U241 (N_241,In_893,In_104);
and U242 (N_242,In_589,In_778);
or U243 (N_243,In_178,In_873);
and U244 (N_244,In_806,In_322);
or U245 (N_245,In_800,In_375);
or U246 (N_246,In_471,In_225);
nor U247 (N_247,In_744,In_66);
or U248 (N_248,In_660,In_462);
nor U249 (N_249,In_752,In_578);
nand U250 (N_250,In_481,In_618);
nor U251 (N_251,In_54,In_976);
nand U252 (N_252,In_987,In_214);
or U253 (N_253,In_72,In_67);
or U254 (N_254,In_843,In_389);
nor U255 (N_255,In_579,In_390);
or U256 (N_256,In_823,In_839);
or U257 (N_257,In_845,In_643);
or U258 (N_258,In_923,In_279);
or U259 (N_259,In_695,In_854);
nand U260 (N_260,In_797,In_760);
nor U261 (N_261,In_241,In_349);
or U262 (N_262,In_994,In_741);
nand U263 (N_263,In_153,In_565);
nand U264 (N_264,In_151,In_679);
and U265 (N_265,In_581,In_698);
nor U266 (N_266,In_143,In_795);
or U267 (N_267,In_125,In_638);
xnor U268 (N_268,In_251,In_529);
nand U269 (N_269,In_250,In_874);
or U270 (N_270,In_211,In_226);
nand U271 (N_271,In_105,In_657);
and U272 (N_272,In_244,In_287);
and U273 (N_273,In_77,In_947);
or U274 (N_274,In_304,In_43);
nand U275 (N_275,In_14,In_423);
and U276 (N_276,In_847,In_785);
nand U277 (N_277,In_619,In_196);
or U278 (N_278,In_544,In_836);
or U279 (N_279,In_636,In_283);
and U280 (N_280,In_359,In_905);
nor U281 (N_281,In_710,In_794);
nand U282 (N_282,In_834,In_326);
nand U283 (N_283,In_637,In_790);
or U284 (N_284,In_323,In_83);
nand U285 (N_285,In_369,In_79);
or U286 (N_286,In_44,In_708);
or U287 (N_287,In_421,In_25);
and U288 (N_288,In_654,In_121);
and U289 (N_289,In_623,In_545);
and U290 (N_290,In_621,In_551);
and U291 (N_291,In_282,In_468);
or U292 (N_292,In_407,In_413);
nand U293 (N_293,In_92,In_898);
or U294 (N_294,In_726,In_915);
or U295 (N_295,In_124,In_640);
or U296 (N_296,In_772,In_576);
and U297 (N_297,In_461,In_713);
nor U298 (N_298,In_669,In_663);
and U299 (N_299,In_371,In_878);
nor U300 (N_300,In_988,In_477);
and U301 (N_301,In_160,In_676);
nor U302 (N_302,In_408,In_327);
nor U303 (N_303,In_719,In_769);
nor U304 (N_304,In_668,In_602);
and U305 (N_305,In_278,In_78);
and U306 (N_306,In_948,In_348);
or U307 (N_307,In_967,In_851);
and U308 (N_308,In_598,In_816);
and U309 (N_309,In_202,In_925);
and U310 (N_310,In_259,In_89);
and U311 (N_311,In_502,In_610);
nor U312 (N_312,In_895,In_158);
and U313 (N_313,In_19,In_537);
or U314 (N_314,In_262,In_398);
nand U315 (N_315,In_284,In_198);
nor U316 (N_316,In_979,In_675);
or U317 (N_317,In_803,In_183);
and U318 (N_318,In_147,In_94);
and U319 (N_319,In_46,In_718);
nand U320 (N_320,In_290,In_186);
or U321 (N_321,In_802,In_317);
nor U322 (N_322,In_921,In_783);
and U323 (N_323,In_904,In_164);
and U324 (N_324,In_632,In_0);
nor U325 (N_325,In_485,In_452);
nor U326 (N_326,In_488,In_254);
nand U327 (N_327,In_498,In_412);
or U328 (N_328,In_764,In_416);
or U329 (N_329,In_233,In_325);
and U330 (N_330,In_248,In_206);
or U331 (N_331,In_120,In_852);
and U332 (N_332,In_999,In_886);
and U333 (N_333,In_392,In_919);
nor U334 (N_334,In_464,In_831);
nor U335 (N_335,In_173,In_311);
and U336 (N_336,In_572,In_45);
and U337 (N_337,In_784,In_825);
nor U338 (N_338,In_344,In_103);
and U339 (N_339,In_29,In_977);
and U340 (N_340,In_10,In_774);
and U341 (N_341,In_253,In_299);
nor U342 (N_342,In_739,In_629);
or U343 (N_343,In_291,In_931);
and U344 (N_344,In_352,In_42);
and U345 (N_345,In_9,In_838);
nand U346 (N_346,In_560,In_58);
nand U347 (N_347,In_587,In_853);
or U348 (N_348,In_993,In_207);
nor U349 (N_349,In_374,In_900);
or U350 (N_350,In_457,In_267);
nor U351 (N_351,In_154,In_388);
nor U352 (N_352,In_21,In_499);
and U353 (N_353,In_850,In_574);
xor U354 (N_354,In_817,In_658);
nand U355 (N_355,In_93,In_748);
or U356 (N_356,In_546,In_463);
and U357 (N_357,In_917,In_296);
or U358 (N_358,In_859,In_437);
nand U359 (N_359,In_607,In_276);
or U360 (N_360,In_696,In_555);
and U361 (N_361,In_801,In_562);
nand U362 (N_362,In_730,In_482);
nand U363 (N_363,In_458,In_897);
and U364 (N_364,In_681,In_779);
and U365 (N_365,In_234,In_27);
nor U366 (N_366,In_773,In_554);
or U367 (N_367,In_35,In_625);
nor U368 (N_368,In_137,In_526);
nand U369 (N_369,In_263,In_245);
or U370 (N_370,In_135,In_360);
nand U371 (N_371,In_433,In_556);
and U372 (N_372,In_367,In_933);
nand U373 (N_373,In_535,In_711);
or U374 (N_374,In_832,In_530);
or U375 (N_375,In_911,In_804);
and U376 (N_376,In_189,In_969);
and U377 (N_377,In_411,In_808);
and U378 (N_378,In_536,In_666);
or U379 (N_379,In_624,In_685);
and U380 (N_380,In_339,In_410);
nand U381 (N_381,In_561,In_759);
or U382 (N_382,In_763,In_386);
nand U383 (N_383,In_614,In_497);
or U384 (N_384,In_717,In_782);
nand U385 (N_385,In_523,In_232);
or U386 (N_386,In_989,In_531);
and U387 (N_387,In_47,In_709);
or U388 (N_388,In_37,In_864);
or U389 (N_389,In_603,In_586);
or U390 (N_390,In_249,In_306);
and U391 (N_391,In_439,In_453);
nor U392 (N_392,In_76,In_686);
nand U393 (N_393,In_553,In_216);
nor U394 (N_394,In_647,In_95);
nand U395 (N_395,In_334,In_780);
and U396 (N_396,In_659,In_302);
nand U397 (N_397,In_316,In_335);
nand U398 (N_398,In_758,In_391);
or U399 (N_399,In_965,In_862);
nand U400 (N_400,In_950,In_427);
or U401 (N_401,In_906,In_107);
nand U402 (N_402,In_60,In_145);
xor U403 (N_403,In_293,In_509);
nand U404 (N_404,In_18,In_996);
nand U405 (N_405,In_628,In_239);
nor U406 (N_406,In_64,In_414);
or U407 (N_407,In_753,In_890);
nor U408 (N_408,In_980,In_218);
or U409 (N_409,In_101,In_889);
and U410 (N_410,In_33,In_15);
or U411 (N_411,In_469,In_880);
and U412 (N_412,In_528,In_510);
and U413 (N_413,In_179,In_913);
or U414 (N_414,In_362,In_907);
nand U415 (N_415,In_786,In_678);
and U416 (N_416,In_212,In_559);
and U417 (N_417,In_448,In_789);
and U418 (N_418,In_656,In_805);
nor U419 (N_419,In_705,In_127);
and U420 (N_420,In_231,In_119);
or U421 (N_421,In_28,In_841);
nand U422 (N_422,In_85,In_144);
or U423 (N_423,In_747,In_750);
or U424 (N_424,In_665,In_513);
nor U425 (N_425,In_114,In_130);
or U426 (N_426,In_550,In_466);
nor U427 (N_427,In_182,In_858);
nor U428 (N_428,In_438,In_432);
or U429 (N_429,In_593,In_243);
nand U430 (N_430,In_740,In_385);
or U431 (N_431,In_516,In_430);
or U432 (N_432,In_908,In_376);
xor U433 (N_433,In_236,In_139);
nand U434 (N_434,In_945,In_4);
and U435 (N_435,In_62,In_23);
or U436 (N_436,In_955,In_56);
and U437 (N_437,In_573,In_749);
xor U438 (N_438,In_633,In_96);
and U439 (N_439,In_356,In_269);
or U440 (N_440,In_830,In_13);
nor U441 (N_441,In_964,In_264);
or U442 (N_442,In_491,In_454);
nand U443 (N_443,In_26,In_566);
nand U444 (N_444,In_140,In_495);
xnor U445 (N_445,In_733,In_768);
or U446 (N_446,In_246,In_275);
nor U447 (N_447,In_599,In_210);
and U448 (N_448,In_641,In_540);
nand U449 (N_449,In_942,In_861);
or U450 (N_450,In_30,In_914);
and U451 (N_451,In_165,In_725);
nand U452 (N_452,In_670,In_883);
nand U453 (N_453,In_40,In_305);
or U454 (N_454,In_288,In_508);
and U455 (N_455,In_138,In_38);
or U456 (N_456,In_459,In_455);
and U457 (N_457,In_59,In_856);
or U458 (N_458,In_543,In_168);
nor U459 (N_459,In_285,In_828);
xor U460 (N_460,In_106,In_888);
xnor U461 (N_461,In_812,In_901);
nor U462 (N_462,In_155,In_738);
nand U463 (N_463,In_756,In_266);
or U464 (N_464,In_217,In_791);
nor U465 (N_465,In_229,In_418);
nand U466 (N_466,In_175,In_731);
and U467 (N_467,In_191,In_420);
or U468 (N_468,In_611,In_292);
or U469 (N_469,In_50,In_370);
and U470 (N_470,In_162,In_297);
or U471 (N_471,In_757,In_867);
and U472 (N_472,In_347,In_557);
nor U473 (N_473,In_986,In_116);
and U474 (N_474,In_133,In_159);
nor U475 (N_475,In_148,In_424);
nand U476 (N_476,In_330,In_286);
nand U477 (N_477,In_377,In_512);
nor U478 (N_478,In_465,In_487);
nand U479 (N_479,In_203,In_547);
or U480 (N_480,In_258,In_961);
nand U481 (N_481,In_863,In_373);
or U482 (N_482,In_307,In_451);
and U483 (N_483,In_846,In_728);
or U484 (N_484,In_329,In_762);
or U485 (N_485,In_7,In_361);
nor U486 (N_486,In_712,In_87);
nand U487 (N_487,In_855,In_700);
nand U488 (N_488,In_936,In_507);
nand U489 (N_489,In_646,In_295);
and U490 (N_490,In_975,In_342);
nor U491 (N_491,In_331,In_123);
or U492 (N_492,In_892,In_177);
or U493 (N_493,In_109,In_552);
nor U494 (N_494,In_315,In_223);
xor U495 (N_495,In_766,In_478);
and U496 (N_496,In_723,In_265);
nor U497 (N_497,In_595,In_781);
or U498 (N_498,In_927,In_575);
or U499 (N_499,In_117,In_734);
or U500 (N_500,In_166,In_195);
nand U501 (N_501,In_209,In_330);
nor U502 (N_502,In_496,In_802);
or U503 (N_503,In_533,In_575);
and U504 (N_504,In_892,In_644);
or U505 (N_505,In_515,In_665);
and U506 (N_506,In_398,In_387);
or U507 (N_507,In_412,In_905);
nand U508 (N_508,In_176,In_526);
or U509 (N_509,In_753,In_431);
and U510 (N_510,In_893,In_347);
or U511 (N_511,In_47,In_147);
nand U512 (N_512,In_903,In_556);
or U513 (N_513,In_103,In_907);
nor U514 (N_514,In_56,In_440);
xor U515 (N_515,In_934,In_154);
and U516 (N_516,In_223,In_620);
nor U517 (N_517,In_389,In_508);
nor U518 (N_518,In_533,In_931);
and U519 (N_519,In_492,In_615);
or U520 (N_520,In_695,In_146);
xor U521 (N_521,In_988,In_764);
nand U522 (N_522,In_487,In_642);
xnor U523 (N_523,In_126,In_160);
nor U524 (N_524,In_719,In_239);
nand U525 (N_525,In_179,In_560);
or U526 (N_526,In_218,In_549);
nand U527 (N_527,In_293,In_194);
nor U528 (N_528,In_873,In_447);
nand U529 (N_529,In_717,In_507);
and U530 (N_530,In_680,In_353);
and U531 (N_531,In_255,In_466);
or U532 (N_532,In_548,In_796);
or U533 (N_533,In_449,In_976);
nand U534 (N_534,In_878,In_649);
and U535 (N_535,In_583,In_748);
and U536 (N_536,In_606,In_10);
nand U537 (N_537,In_484,In_302);
and U538 (N_538,In_422,In_774);
nand U539 (N_539,In_541,In_793);
or U540 (N_540,In_693,In_614);
or U541 (N_541,In_139,In_620);
nand U542 (N_542,In_723,In_341);
and U543 (N_543,In_397,In_821);
and U544 (N_544,In_99,In_795);
or U545 (N_545,In_761,In_503);
or U546 (N_546,In_546,In_982);
and U547 (N_547,In_77,In_310);
nor U548 (N_548,In_39,In_145);
xor U549 (N_549,In_110,In_210);
and U550 (N_550,In_553,In_401);
xnor U551 (N_551,In_764,In_626);
nor U552 (N_552,In_749,In_766);
nor U553 (N_553,In_624,In_466);
or U554 (N_554,In_738,In_489);
nand U555 (N_555,In_485,In_840);
and U556 (N_556,In_783,In_833);
and U557 (N_557,In_841,In_352);
xor U558 (N_558,In_650,In_779);
or U559 (N_559,In_505,In_794);
and U560 (N_560,In_282,In_708);
nor U561 (N_561,In_167,In_674);
nor U562 (N_562,In_11,In_616);
nor U563 (N_563,In_928,In_598);
or U564 (N_564,In_496,In_210);
or U565 (N_565,In_243,In_234);
nor U566 (N_566,In_872,In_583);
or U567 (N_567,In_495,In_249);
or U568 (N_568,In_367,In_688);
and U569 (N_569,In_641,In_0);
and U570 (N_570,In_57,In_821);
nand U571 (N_571,In_669,In_314);
and U572 (N_572,In_902,In_443);
and U573 (N_573,In_23,In_676);
and U574 (N_574,In_860,In_47);
or U575 (N_575,In_852,In_718);
and U576 (N_576,In_777,In_370);
nand U577 (N_577,In_51,In_717);
and U578 (N_578,In_170,In_898);
or U579 (N_579,In_957,In_834);
and U580 (N_580,In_886,In_605);
or U581 (N_581,In_564,In_169);
nand U582 (N_582,In_387,In_181);
nand U583 (N_583,In_508,In_920);
or U584 (N_584,In_564,In_94);
and U585 (N_585,In_322,In_229);
or U586 (N_586,In_531,In_683);
nand U587 (N_587,In_483,In_823);
xnor U588 (N_588,In_348,In_43);
nand U589 (N_589,In_50,In_522);
nor U590 (N_590,In_448,In_455);
nor U591 (N_591,In_754,In_295);
and U592 (N_592,In_112,In_485);
nand U593 (N_593,In_234,In_4);
nand U594 (N_594,In_83,In_362);
or U595 (N_595,In_180,In_193);
and U596 (N_596,In_706,In_979);
nand U597 (N_597,In_81,In_718);
nand U598 (N_598,In_829,In_358);
nor U599 (N_599,In_122,In_767);
nand U600 (N_600,In_412,In_648);
xor U601 (N_601,In_537,In_861);
or U602 (N_602,In_501,In_423);
nand U603 (N_603,In_11,In_443);
nor U604 (N_604,In_997,In_564);
or U605 (N_605,In_718,In_977);
or U606 (N_606,In_75,In_806);
nand U607 (N_607,In_861,In_607);
nand U608 (N_608,In_288,In_821);
and U609 (N_609,In_640,In_271);
or U610 (N_610,In_139,In_102);
or U611 (N_611,In_900,In_715);
nand U612 (N_612,In_549,In_927);
nor U613 (N_613,In_204,In_744);
or U614 (N_614,In_856,In_931);
and U615 (N_615,In_934,In_532);
nand U616 (N_616,In_160,In_497);
or U617 (N_617,In_52,In_443);
or U618 (N_618,In_126,In_696);
or U619 (N_619,In_573,In_360);
nor U620 (N_620,In_105,In_157);
nand U621 (N_621,In_492,In_838);
nand U622 (N_622,In_851,In_763);
nor U623 (N_623,In_284,In_792);
nor U624 (N_624,In_41,In_990);
nand U625 (N_625,In_194,In_591);
xor U626 (N_626,In_519,In_849);
and U627 (N_627,In_659,In_216);
and U628 (N_628,In_309,In_100);
or U629 (N_629,In_787,In_392);
nand U630 (N_630,In_407,In_962);
and U631 (N_631,In_639,In_418);
nand U632 (N_632,In_465,In_12);
and U633 (N_633,In_438,In_509);
nand U634 (N_634,In_473,In_950);
nand U635 (N_635,In_354,In_771);
or U636 (N_636,In_591,In_184);
and U637 (N_637,In_572,In_373);
nand U638 (N_638,In_410,In_175);
or U639 (N_639,In_766,In_433);
nand U640 (N_640,In_467,In_92);
and U641 (N_641,In_606,In_244);
nor U642 (N_642,In_369,In_794);
nand U643 (N_643,In_181,In_43);
and U644 (N_644,In_984,In_432);
and U645 (N_645,In_869,In_886);
nand U646 (N_646,In_13,In_630);
nor U647 (N_647,In_838,In_930);
and U648 (N_648,In_50,In_330);
nor U649 (N_649,In_645,In_295);
and U650 (N_650,In_7,In_924);
and U651 (N_651,In_997,In_359);
and U652 (N_652,In_710,In_974);
or U653 (N_653,In_914,In_684);
and U654 (N_654,In_608,In_901);
nor U655 (N_655,In_559,In_853);
or U656 (N_656,In_878,In_58);
nor U657 (N_657,In_935,In_1);
nand U658 (N_658,In_943,In_336);
nand U659 (N_659,In_865,In_416);
nor U660 (N_660,In_30,In_317);
xnor U661 (N_661,In_154,In_616);
nor U662 (N_662,In_230,In_434);
and U663 (N_663,In_564,In_397);
nor U664 (N_664,In_866,In_639);
nor U665 (N_665,In_680,In_261);
or U666 (N_666,In_520,In_360);
nand U667 (N_667,In_527,In_915);
and U668 (N_668,In_337,In_114);
nand U669 (N_669,In_122,In_598);
or U670 (N_670,In_443,In_698);
or U671 (N_671,In_184,In_394);
xnor U672 (N_672,In_126,In_333);
or U673 (N_673,In_831,In_628);
nand U674 (N_674,In_554,In_371);
nor U675 (N_675,In_314,In_335);
nand U676 (N_676,In_200,In_487);
nor U677 (N_677,In_935,In_936);
or U678 (N_678,In_260,In_110);
and U679 (N_679,In_128,In_845);
nand U680 (N_680,In_461,In_627);
nor U681 (N_681,In_84,In_858);
and U682 (N_682,In_691,In_376);
nor U683 (N_683,In_923,In_543);
or U684 (N_684,In_610,In_725);
nand U685 (N_685,In_155,In_998);
or U686 (N_686,In_344,In_301);
or U687 (N_687,In_500,In_380);
and U688 (N_688,In_497,In_394);
nand U689 (N_689,In_464,In_186);
and U690 (N_690,In_73,In_273);
and U691 (N_691,In_506,In_726);
nor U692 (N_692,In_949,In_345);
and U693 (N_693,In_908,In_803);
nand U694 (N_694,In_888,In_528);
and U695 (N_695,In_715,In_925);
nand U696 (N_696,In_198,In_127);
and U697 (N_697,In_809,In_748);
and U698 (N_698,In_611,In_501);
nand U699 (N_699,In_79,In_154);
nand U700 (N_700,In_780,In_940);
and U701 (N_701,In_767,In_467);
and U702 (N_702,In_37,In_322);
nor U703 (N_703,In_582,In_196);
or U704 (N_704,In_96,In_192);
nand U705 (N_705,In_472,In_635);
nand U706 (N_706,In_850,In_641);
nand U707 (N_707,In_424,In_245);
or U708 (N_708,In_715,In_861);
xor U709 (N_709,In_303,In_736);
nor U710 (N_710,In_325,In_997);
or U711 (N_711,In_712,In_935);
nor U712 (N_712,In_631,In_953);
nand U713 (N_713,In_456,In_779);
and U714 (N_714,In_347,In_123);
or U715 (N_715,In_77,In_897);
nand U716 (N_716,In_71,In_430);
and U717 (N_717,In_908,In_706);
or U718 (N_718,In_784,In_435);
nand U719 (N_719,In_234,In_861);
nor U720 (N_720,In_776,In_463);
nor U721 (N_721,In_70,In_889);
and U722 (N_722,In_403,In_181);
or U723 (N_723,In_273,In_785);
nor U724 (N_724,In_46,In_513);
nor U725 (N_725,In_15,In_709);
nand U726 (N_726,In_570,In_136);
nor U727 (N_727,In_957,In_625);
and U728 (N_728,In_2,In_556);
or U729 (N_729,In_861,In_54);
nor U730 (N_730,In_80,In_674);
nor U731 (N_731,In_556,In_825);
and U732 (N_732,In_524,In_924);
or U733 (N_733,In_426,In_663);
nor U734 (N_734,In_404,In_744);
and U735 (N_735,In_421,In_328);
nand U736 (N_736,In_181,In_746);
or U737 (N_737,In_229,In_570);
or U738 (N_738,In_286,In_484);
and U739 (N_739,In_443,In_656);
and U740 (N_740,In_509,In_782);
nand U741 (N_741,In_575,In_461);
nand U742 (N_742,In_329,In_544);
nor U743 (N_743,In_764,In_189);
and U744 (N_744,In_943,In_281);
nor U745 (N_745,In_296,In_246);
or U746 (N_746,In_746,In_486);
and U747 (N_747,In_251,In_860);
nor U748 (N_748,In_445,In_690);
nor U749 (N_749,In_8,In_228);
or U750 (N_750,In_947,In_979);
nand U751 (N_751,In_208,In_414);
nand U752 (N_752,In_584,In_781);
and U753 (N_753,In_867,In_901);
nor U754 (N_754,In_627,In_591);
nand U755 (N_755,In_496,In_349);
nor U756 (N_756,In_822,In_525);
and U757 (N_757,In_157,In_531);
or U758 (N_758,In_641,In_392);
and U759 (N_759,In_833,In_516);
or U760 (N_760,In_803,In_911);
or U761 (N_761,In_303,In_306);
and U762 (N_762,In_323,In_243);
and U763 (N_763,In_985,In_249);
nand U764 (N_764,In_215,In_204);
nand U765 (N_765,In_435,In_512);
nor U766 (N_766,In_522,In_654);
nor U767 (N_767,In_924,In_531);
nor U768 (N_768,In_771,In_478);
and U769 (N_769,In_401,In_313);
nor U770 (N_770,In_769,In_896);
nor U771 (N_771,In_654,In_418);
nor U772 (N_772,In_946,In_38);
and U773 (N_773,In_314,In_251);
or U774 (N_774,In_295,In_710);
and U775 (N_775,In_562,In_967);
nand U776 (N_776,In_91,In_895);
and U777 (N_777,In_137,In_813);
nand U778 (N_778,In_842,In_981);
and U779 (N_779,In_719,In_149);
nor U780 (N_780,In_18,In_667);
nor U781 (N_781,In_588,In_565);
nor U782 (N_782,In_984,In_125);
or U783 (N_783,In_476,In_242);
nor U784 (N_784,In_606,In_608);
nor U785 (N_785,In_143,In_579);
and U786 (N_786,In_771,In_882);
nand U787 (N_787,In_302,In_734);
nor U788 (N_788,In_240,In_434);
and U789 (N_789,In_414,In_286);
or U790 (N_790,In_113,In_229);
nor U791 (N_791,In_696,In_120);
or U792 (N_792,In_375,In_504);
or U793 (N_793,In_445,In_17);
and U794 (N_794,In_915,In_4);
nor U795 (N_795,In_377,In_13);
nand U796 (N_796,In_957,In_399);
and U797 (N_797,In_248,In_303);
nand U798 (N_798,In_868,In_511);
nand U799 (N_799,In_460,In_227);
nor U800 (N_800,In_135,In_129);
nand U801 (N_801,In_718,In_878);
nand U802 (N_802,In_324,In_0);
nor U803 (N_803,In_759,In_649);
and U804 (N_804,In_881,In_871);
and U805 (N_805,In_644,In_451);
and U806 (N_806,In_85,In_847);
or U807 (N_807,In_570,In_459);
nor U808 (N_808,In_788,In_725);
and U809 (N_809,In_297,In_181);
nand U810 (N_810,In_307,In_156);
nor U811 (N_811,In_710,In_85);
and U812 (N_812,In_263,In_241);
nor U813 (N_813,In_706,In_300);
or U814 (N_814,In_248,In_953);
or U815 (N_815,In_336,In_342);
nor U816 (N_816,In_833,In_768);
nand U817 (N_817,In_260,In_115);
nand U818 (N_818,In_290,In_945);
nor U819 (N_819,In_107,In_29);
nand U820 (N_820,In_593,In_863);
and U821 (N_821,In_349,In_314);
xor U822 (N_822,In_757,In_144);
and U823 (N_823,In_670,In_880);
nor U824 (N_824,In_389,In_322);
and U825 (N_825,In_757,In_241);
or U826 (N_826,In_543,In_475);
nand U827 (N_827,In_481,In_635);
or U828 (N_828,In_102,In_551);
and U829 (N_829,In_693,In_202);
and U830 (N_830,In_516,In_925);
and U831 (N_831,In_477,In_207);
or U832 (N_832,In_142,In_441);
or U833 (N_833,In_424,In_182);
nand U834 (N_834,In_204,In_268);
nand U835 (N_835,In_594,In_495);
and U836 (N_836,In_45,In_620);
or U837 (N_837,In_662,In_497);
nand U838 (N_838,In_658,In_853);
nand U839 (N_839,In_988,In_873);
nand U840 (N_840,In_458,In_85);
nor U841 (N_841,In_604,In_879);
nand U842 (N_842,In_6,In_14);
and U843 (N_843,In_837,In_556);
xnor U844 (N_844,In_572,In_749);
nor U845 (N_845,In_428,In_58);
nand U846 (N_846,In_127,In_903);
nor U847 (N_847,In_561,In_75);
nor U848 (N_848,In_673,In_273);
nor U849 (N_849,In_628,In_840);
nor U850 (N_850,In_749,In_992);
nor U851 (N_851,In_926,In_111);
and U852 (N_852,In_268,In_380);
nor U853 (N_853,In_217,In_208);
or U854 (N_854,In_678,In_777);
nand U855 (N_855,In_31,In_557);
nor U856 (N_856,In_716,In_216);
and U857 (N_857,In_708,In_690);
and U858 (N_858,In_722,In_787);
and U859 (N_859,In_530,In_535);
nor U860 (N_860,In_832,In_211);
nand U861 (N_861,In_110,In_279);
nand U862 (N_862,In_97,In_712);
and U863 (N_863,In_548,In_375);
and U864 (N_864,In_165,In_133);
nor U865 (N_865,In_698,In_631);
and U866 (N_866,In_902,In_880);
xnor U867 (N_867,In_316,In_909);
and U868 (N_868,In_20,In_726);
or U869 (N_869,In_749,In_386);
and U870 (N_870,In_743,In_952);
and U871 (N_871,In_447,In_338);
or U872 (N_872,In_503,In_197);
and U873 (N_873,In_243,In_959);
and U874 (N_874,In_957,In_201);
or U875 (N_875,In_281,In_95);
nor U876 (N_876,In_845,In_256);
or U877 (N_877,In_196,In_261);
and U878 (N_878,In_984,In_613);
and U879 (N_879,In_517,In_982);
or U880 (N_880,In_404,In_389);
nor U881 (N_881,In_277,In_0);
nor U882 (N_882,In_569,In_75);
nand U883 (N_883,In_663,In_368);
nor U884 (N_884,In_622,In_821);
or U885 (N_885,In_994,In_594);
nor U886 (N_886,In_957,In_77);
and U887 (N_887,In_711,In_387);
or U888 (N_888,In_912,In_181);
and U889 (N_889,In_709,In_140);
and U890 (N_890,In_840,In_184);
and U891 (N_891,In_5,In_117);
and U892 (N_892,In_369,In_490);
nor U893 (N_893,In_788,In_995);
nor U894 (N_894,In_702,In_527);
nand U895 (N_895,In_964,In_762);
nand U896 (N_896,In_453,In_470);
or U897 (N_897,In_883,In_710);
and U898 (N_898,In_494,In_933);
nor U899 (N_899,In_876,In_575);
or U900 (N_900,In_653,In_660);
nor U901 (N_901,In_424,In_39);
and U902 (N_902,In_637,In_57);
nand U903 (N_903,In_488,In_578);
and U904 (N_904,In_240,In_570);
xnor U905 (N_905,In_224,In_418);
nand U906 (N_906,In_878,In_952);
nand U907 (N_907,In_866,In_313);
nand U908 (N_908,In_752,In_634);
and U909 (N_909,In_721,In_495);
or U910 (N_910,In_800,In_806);
nor U911 (N_911,In_509,In_827);
and U912 (N_912,In_4,In_780);
and U913 (N_913,In_371,In_432);
and U914 (N_914,In_403,In_975);
nor U915 (N_915,In_239,In_224);
and U916 (N_916,In_514,In_513);
or U917 (N_917,In_583,In_650);
nor U918 (N_918,In_29,In_589);
or U919 (N_919,In_997,In_862);
xor U920 (N_920,In_362,In_481);
nand U921 (N_921,In_401,In_951);
nor U922 (N_922,In_321,In_675);
nand U923 (N_923,In_322,In_462);
or U924 (N_924,In_181,In_5);
nand U925 (N_925,In_652,In_86);
or U926 (N_926,In_160,In_62);
nand U927 (N_927,In_272,In_647);
or U928 (N_928,In_156,In_841);
and U929 (N_929,In_365,In_989);
and U930 (N_930,In_903,In_427);
nand U931 (N_931,In_930,In_154);
and U932 (N_932,In_967,In_757);
and U933 (N_933,In_16,In_806);
nor U934 (N_934,In_327,In_569);
nor U935 (N_935,In_324,In_503);
nand U936 (N_936,In_118,In_242);
or U937 (N_937,In_920,In_52);
and U938 (N_938,In_721,In_346);
and U939 (N_939,In_610,In_814);
nand U940 (N_940,In_697,In_869);
and U941 (N_941,In_165,In_42);
nand U942 (N_942,In_949,In_470);
nand U943 (N_943,In_292,In_873);
and U944 (N_944,In_670,In_231);
nor U945 (N_945,In_486,In_39);
and U946 (N_946,In_165,In_706);
nand U947 (N_947,In_435,In_64);
or U948 (N_948,In_143,In_168);
and U949 (N_949,In_63,In_423);
and U950 (N_950,In_149,In_148);
and U951 (N_951,In_227,In_173);
nor U952 (N_952,In_473,In_351);
nand U953 (N_953,In_27,In_106);
and U954 (N_954,In_26,In_874);
and U955 (N_955,In_691,In_126);
and U956 (N_956,In_933,In_623);
nand U957 (N_957,In_479,In_577);
nand U958 (N_958,In_760,In_529);
nor U959 (N_959,In_959,In_188);
xnor U960 (N_960,In_461,In_579);
and U961 (N_961,In_183,In_61);
and U962 (N_962,In_345,In_230);
or U963 (N_963,In_992,In_694);
and U964 (N_964,In_884,In_81);
or U965 (N_965,In_116,In_170);
and U966 (N_966,In_790,In_66);
and U967 (N_967,In_121,In_574);
nor U968 (N_968,In_987,In_801);
nand U969 (N_969,In_780,In_523);
and U970 (N_970,In_711,In_617);
nand U971 (N_971,In_879,In_64);
or U972 (N_972,In_683,In_844);
or U973 (N_973,In_460,In_382);
and U974 (N_974,In_657,In_601);
nor U975 (N_975,In_967,In_841);
or U976 (N_976,In_764,In_192);
and U977 (N_977,In_913,In_878);
or U978 (N_978,In_581,In_6);
and U979 (N_979,In_282,In_749);
or U980 (N_980,In_503,In_632);
nor U981 (N_981,In_90,In_796);
and U982 (N_982,In_293,In_247);
or U983 (N_983,In_275,In_72);
or U984 (N_984,In_353,In_665);
and U985 (N_985,In_759,In_281);
or U986 (N_986,In_370,In_270);
and U987 (N_987,In_227,In_568);
nand U988 (N_988,In_624,In_62);
nand U989 (N_989,In_57,In_388);
xor U990 (N_990,In_945,In_254);
and U991 (N_991,In_692,In_78);
nor U992 (N_992,In_358,In_737);
and U993 (N_993,In_120,In_763);
and U994 (N_994,In_104,In_433);
nor U995 (N_995,In_159,In_901);
or U996 (N_996,In_379,In_534);
nand U997 (N_997,In_252,In_967);
nand U998 (N_998,In_87,In_171);
or U999 (N_999,In_895,In_770);
nand U1000 (N_1000,N_515,N_209);
nor U1001 (N_1001,N_85,N_21);
nor U1002 (N_1002,N_348,N_0);
nand U1003 (N_1003,N_216,N_736);
or U1004 (N_1004,N_935,N_851);
and U1005 (N_1005,N_501,N_39);
nor U1006 (N_1006,N_932,N_127);
nand U1007 (N_1007,N_861,N_247);
nor U1008 (N_1008,N_810,N_176);
nand U1009 (N_1009,N_997,N_218);
and U1010 (N_1010,N_587,N_337);
nand U1011 (N_1011,N_600,N_390);
nor U1012 (N_1012,N_959,N_947);
nand U1013 (N_1013,N_219,N_112);
and U1014 (N_1014,N_551,N_150);
and U1015 (N_1015,N_760,N_86);
and U1016 (N_1016,N_36,N_647);
or U1017 (N_1017,N_771,N_584);
xnor U1018 (N_1018,N_184,N_89);
or U1019 (N_1019,N_537,N_929);
and U1020 (N_1020,N_152,N_496);
nand U1021 (N_1021,N_333,N_78);
or U1022 (N_1022,N_80,N_814);
nand U1023 (N_1023,N_875,N_548);
or U1024 (N_1024,N_714,N_31);
nand U1025 (N_1025,N_938,N_290);
nand U1026 (N_1026,N_778,N_463);
nand U1027 (N_1027,N_344,N_960);
nor U1028 (N_1028,N_481,N_255);
nand U1029 (N_1029,N_583,N_962);
or U1030 (N_1030,N_822,N_759);
nand U1031 (N_1031,N_111,N_448);
and U1032 (N_1032,N_624,N_241);
and U1033 (N_1033,N_968,N_418);
or U1034 (N_1034,N_664,N_104);
and U1035 (N_1035,N_79,N_285);
or U1036 (N_1036,N_202,N_565);
or U1037 (N_1037,N_301,N_883);
nand U1038 (N_1038,N_137,N_697);
nor U1039 (N_1039,N_735,N_471);
and U1040 (N_1040,N_453,N_803);
nand U1041 (N_1041,N_821,N_941);
and U1042 (N_1042,N_748,N_654);
nor U1043 (N_1043,N_722,N_110);
nand U1044 (N_1044,N_68,N_130);
and U1045 (N_1045,N_939,N_377);
or U1046 (N_1046,N_563,N_543);
nand U1047 (N_1047,N_914,N_281);
or U1048 (N_1048,N_553,N_222);
or U1049 (N_1049,N_922,N_944);
nand U1050 (N_1050,N_456,N_532);
nor U1051 (N_1051,N_863,N_884);
nor U1052 (N_1052,N_250,N_720);
nor U1053 (N_1053,N_592,N_383);
nand U1054 (N_1054,N_887,N_574);
or U1055 (N_1055,N_829,N_106);
and U1056 (N_1056,N_895,N_562);
xor U1057 (N_1057,N_375,N_120);
nand U1058 (N_1058,N_906,N_610);
nand U1059 (N_1059,N_890,N_510);
and U1060 (N_1060,N_267,N_159);
and U1061 (N_1061,N_846,N_332);
and U1062 (N_1062,N_633,N_279);
or U1063 (N_1063,N_916,N_564);
and U1064 (N_1064,N_168,N_165);
or U1065 (N_1065,N_276,N_527);
or U1066 (N_1066,N_589,N_685);
and U1067 (N_1067,N_995,N_561);
nand U1068 (N_1068,N_619,N_528);
and U1069 (N_1069,N_64,N_795);
nor U1070 (N_1070,N_825,N_94);
or U1071 (N_1071,N_368,N_950);
nor U1072 (N_1072,N_193,N_384);
nand U1073 (N_1073,N_793,N_369);
nand U1074 (N_1074,N_6,N_292);
nor U1075 (N_1075,N_965,N_200);
nor U1076 (N_1076,N_310,N_792);
nand U1077 (N_1077,N_27,N_198);
nand U1078 (N_1078,N_770,N_540);
nor U1079 (N_1079,N_151,N_12);
or U1080 (N_1080,N_177,N_430);
or U1081 (N_1081,N_275,N_262);
and U1082 (N_1082,N_270,N_781);
nor U1083 (N_1083,N_840,N_167);
nor U1084 (N_1084,N_409,N_180);
or U1085 (N_1085,N_831,N_924);
nor U1086 (N_1086,N_314,N_539);
nand U1087 (N_1087,N_242,N_323);
nor U1088 (N_1088,N_772,N_755);
nor U1089 (N_1089,N_309,N_33);
nand U1090 (N_1090,N_316,N_625);
nor U1091 (N_1091,N_598,N_918);
or U1092 (N_1092,N_889,N_674);
or U1093 (N_1093,N_227,N_91);
or U1094 (N_1094,N_737,N_236);
nor U1095 (N_1095,N_656,N_252);
or U1096 (N_1096,N_53,N_980);
and U1097 (N_1097,N_148,N_7);
nand U1098 (N_1098,N_261,N_100);
or U1099 (N_1099,N_933,N_170);
or U1100 (N_1100,N_635,N_949);
and U1101 (N_1101,N_660,N_166);
nor U1102 (N_1102,N_305,N_313);
nand U1103 (N_1103,N_204,N_853);
nand U1104 (N_1104,N_596,N_511);
nor U1105 (N_1105,N_730,N_491);
or U1106 (N_1106,N_293,N_899);
nand U1107 (N_1107,N_238,N_132);
or U1108 (N_1108,N_212,N_901);
nor U1109 (N_1109,N_860,N_682);
nand U1110 (N_1110,N_81,N_15);
or U1111 (N_1111,N_766,N_83);
nand U1112 (N_1112,N_666,N_359);
or U1113 (N_1113,N_670,N_604);
and U1114 (N_1114,N_70,N_497);
or U1115 (N_1115,N_3,N_639);
or U1116 (N_1116,N_535,N_63);
and U1117 (N_1117,N_44,N_577);
and U1118 (N_1118,N_109,N_740);
and U1119 (N_1119,N_458,N_345);
and U1120 (N_1120,N_277,N_459);
nand U1121 (N_1121,N_580,N_67);
or U1122 (N_1122,N_894,N_213);
nand U1123 (N_1123,N_17,N_582);
and U1124 (N_1124,N_628,N_547);
nor U1125 (N_1125,N_122,N_665);
and U1126 (N_1126,N_61,N_597);
nor U1127 (N_1127,N_379,N_174);
and U1128 (N_1128,N_963,N_489);
or U1129 (N_1129,N_723,N_676);
nor U1130 (N_1130,N_975,N_672);
or U1131 (N_1131,N_392,N_542);
nand U1132 (N_1132,N_964,N_342);
nor U1133 (N_1133,N_444,N_928);
nand U1134 (N_1134,N_178,N_357);
and U1135 (N_1135,N_645,N_23);
or U1136 (N_1136,N_857,N_492);
nand U1137 (N_1137,N_273,N_677);
and U1138 (N_1138,N_620,N_335);
and U1139 (N_1139,N_762,N_438);
and U1140 (N_1140,N_441,N_678);
or U1141 (N_1141,N_671,N_451);
nand U1142 (N_1142,N_526,N_49);
nor U1143 (N_1143,N_284,N_160);
nand U1144 (N_1144,N_5,N_60);
nand U1145 (N_1145,N_35,N_454);
and U1146 (N_1146,N_787,N_719);
and U1147 (N_1147,N_721,N_668);
or U1148 (N_1148,N_606,N_338);
nand U1149 (N_1149,N_50,N_278);
nor U1150 (N_1150,N_406,N_773);
nor U1151 (N_1151,N_791,N_559);
nor U1152 (N_1152,N_864,N_123);
nor U1153 (N_1153,N_657,N_217);
nand U1154 (N_1154,N_783,N_321);
nand U1155 (N_1155,N_426,N_758);
and U1156 (N_1156,N_673,N_162);
nand U1157 (N_1157,N_298,N_402);
or U1158 (N_1158,N_847,N_228);
nor U1159 (N_1159,N_374,N_419);
nor U1160 (N_1160,N_994,N_818);
xor U1161 (N_1161,N_744,N_991);
nand U1162 (N_1162,N_591,N_424);
or U1163 (N_1163,N_993,N_832);
xnor U1164 (N_1164,N_196,N_627);
or U1165 (N_1165,N_530,N_414);
nor U1166 (N_1166,N_294,N_182);
and U1167 (N_1167,N_513,N_552);
nand U1168 (N_1168,N_893,N_943);
or U1169 (N_1169,N_412,N_520);
nor U1170 (N_1170,N_769,N_362);
nand U1171 (N_1171,N_128,N_696);
nand U1172 (N_1172,N_339,N_990);
and U1173 (N_1173,N_912,N_692);
nand U1174 (N_1174,N_806,N_880);
nor U1175 (N_1175,N_705,N_571);
nor U1176 (N_1176,N_554,N_920);
nand U1177 (N_1177,N_40,N_655);
nor U1178 (N_1178,N_907,N_784);
and U1179 (N_1179,N_304,N_979);
nand U1180 (N_1180,N_869,N_891);
and U1181 (N_1181,N_917,N_74);
and U1182 (N_1182,N_19,N_486);
or U1183 (N_1183,N_650,N_560);
nand U1184 (N_1184,N_585,N_649);
and U1185 (N_1185,N_897,N_833);
nand U1186 (N_1186,N_229,N_779);
or U1187 (N_1187,N_157,N_545);
and U1188 (N_1188,N_147,N_190);
nand U1189 (N_1189,N_312,N_428);
xnor U1190 (N_1190,N_488,N_955);
and U1191 (N_1191,N_601,N_62);
xnor U1192 (N_1192,N_476,N_487);
nand U1193 (N_1193,N_900,N_119);
nand U1194 (N_1194,N_498,N_318);
nand U1195 (N_1195,N_181,N_808);
and U1196 (N_1196,N_461,N_282);
or U1197 (N_1197,N_156,N_14);
or U1198 (N_1198,N_37,N_504);
or U1199 (N_1199,N_616,N_9);
and U1200 (N_1200,N_11,N_754);
nor U1201 (N_1201,N_927,N_794);
or U1202 (N_1202,N_24,N_16);
nor U1203 (N_1203,N_474,N_734);
nand U1204 (N_1204,N_214,N_437);
nand U1205 (N_1205,N_509,N_324);
or U1206 (N_1206,N_455,N_88);
nand U1207 (N_1207,N_425,N_707);
and U1208 (N_1208,N_191,N_500);
nor U1209 (N_1209,N_823,N_984);
and U1210 (N_1210,N_667,N_612);
nor U1211 (N_1211,N_838,N_34);
nand U1212 (N_1212,N_113,N_925);
nor U1213 (N_1213,N_370,N_519);
nor U1214 (N_1214,N_394,N_179);
xnor U1215 (N_1215,N_593,N_4);
nor U1216 (N_1216,N_470,N_490);
nor U1217 (N_1217,N_629,N_199);
nand U1218 (N_1218,N_796,N_764);
and U1219 (N_1219,N_765,N_435);
nand U1220 (N_1220,N_381,N_642);
nor U1221 (N_1221,N_133,N_231);
nand U1222 (N_1222,N_709,N_237);
or U1223 (N_1223,N_55,N_988);
and U1224 (N_1224,N_364,N_852);
nor U1225 (N_1225,N_187,N_856);
nor U1226 (N_1226,N_114,N_817);
nand U1227 (N_1227,N_144,N_274);
or U1228 (N_1228,N_983,N_878);
nand U1229 (N_1229,N_103,N_42);
nor U1230 (N_1230,N_961,N_420);
nor U1231 (N_1231,N_566,N_82);
nor U1232 (N_1232,N_615,N_630);
or U1233 (N_1233,N_839,N_834);
nor U1234 (N_1234,N_328,N_84);
or U1235 (N_1235,N_439,N_373);
nand U1236 (N_1236,N_235,N_475);
nand U1237 (N_1237,N_725,N_651);
nor U1238 (N_1238,N_269,N_715);
xor U1239 (N_1239,N_266,N_595);
nor U1240 (N_1240,N_976,N_608);
nand U1241 (N_1241,N_395,N_549);
nand U1242 (N_1242,N_265,N_815);
and U1243 (N_1243,N_41,N_399);
and U1244 (N_1244,N_909,N_46);
or U1245 (N_1245,N_322,N_751);
nor U1246 (N_1246,N_32,N_77);
and U1247 (N_1247,N_978,N_879);
or U1248 (N_1248,N_538,N_805);
nand U1249 (N_1249,N_18,N_675);
or U1250 (N_1250,N_465,N_248);
and U1251 (N_1251,N_87,N_798);
nor U1252 (N_1252,N_609,N_807);
nor U1253 (N_1253,N_20,N_249);
nor U1254 (N_1254,N_172,N_524);
nand U1255 (N_1255,N_816,N_69);
nand U1256 (N_1256,N_643,N_516);
or U1257 (N_1257,N_578,N_403);
nand U1258 (N_1258,N_862,N_320);
and U1259 (N_1259,N_923,N_361);
or U1260 (N_1260,N_686,N_733);
and U1261 (N_1261,N_135,N_712);
nand U1262 (N_1262,N_349,N_391);
and U1263 (N_1263,N_786,N_529);
and U1264 (N_1264,N_175,N_155);
and U1265 (N_1265,N_969,N_65);
nor U1266 (N_1266,N_108,N_299);
nand U1267 (N_1267,N_306,N_54);
or U1268 (N_1268,N_953,N_272);
and U1269 (N_1269,N_812,N_71);
nor U1270 (N_1270,N_347,N_908);
nor U1271 (N_1271,N_747,N_346);
nand U1272 (N_1272,N_905,N_681);
nand U1273 (N_1273,N_809,N_43);
or U1274 (N_1274,N_605,N_703);
and U1275 (N_1275,N_830,N_802);
and U1276 (N_1276,N_291,N_257);
nor U1277 (N_1277,N_124,N_843);
nor U1278 (N_1278,N_367,N_945);
and U1279 (N_1279,N_508,N_75);
or U1280 (N_1280,N_462,N_544);
or U1281 (N_1281,N_371,N_505);
nand U1282 (N_1282,N_205,N_97);
or U1283 (N_1283,N_244,N_940);
nand U1284 (N_1284,N_776,N_96);
nor U1285 (N_1285,N_763,N_996);
nor U1286 (N_1286,N_930,N_724);
nor U1287 (N_1287,N_26,N_886);
and U1288 (N_1288,N_404,N_360);
nand U1289 (N_1289,N_57,N_824);
nand U1290 (N_1290,N_263,N_317);
and U1291 (N_1291,N_297,N_844);
nor U1292 (N_1292,N_226,N_141);
nor U1293 (N_1293,N_289,N_1);
or U1294 (N_1294,N_753,N_708);
and U1295 (N_1295,N_107,N_479);
nand U1296 (N_1296,N_576,N_203);
nor U1297 (N_1297,N_201,N_325);
nor U1298 (N_1298,N_457,N_607);
nand U1299 (N_1299,N_621,N_623);
nand U1300 (N_1300,N_240,N_259);
or U1301 (N_1301,N_573,N_870);
nor U1302 (N_1302,N_389,N_485);
and U1303 (N_1303,N_48,N_836);
or U1304 (N_1304,N_308,N_503);
xnor U1305 (N_1305,N_183,N_173);
or U1306 (N_1306,N_892,N_998);
or U1307 (N_1307,N_466,N_447);
nand U1308 (N_1308,N_385,N_931);
nor U1309 (N_1309,N_101,N_326);
and U1310 (N_1310,N_121,N_102);
and U1311 (N_1311,N_659,N_850);
nand U1312 (N_1312,N_827,N_286);
or U1313 (N_1313,N_154,N_260);
nand U1314 (N_1314,N_613,N_690);
nand U1315 (N_1315,N_253,N_365);
nand U1316 (N_1316,N_602,N_207);
and U1317 (N_1317,N_729,N_431);
nor U1318 (N_1318,N_334,N_855);
xor U1319 (N_1319,N_521,N_256);
and U1320 (N_1320,N_713,N_268);
or U1321 (N_1321,N_866,N_845);
or U1322 (N_1322,N_728,N_954);
and U1323 (N_1323,N_429,N_688);
nand U1324 (N_1324,N_820,N_98);
nor U1325 (N_1325,N_568,N_987);
and U1326 (N_1326,N_220,N_469);
and U1327 (N_1327,N_254,N_415);
nand U1328 (N_1328,N_710,N_859);
or U1329 (N_1329,N_958,N_319);
nand U1330 (N_1330,N_327,N_115);
xor U1331 (N_1331,N_484,N_731);
xor U1332 (N_1332,N_417,N_694);
and U1333 (N_1333,N_433,N_258);
nor U1334 (N_1334,N_646,N_185);
nor U1335 (N_1335,N_421,N_788);
and U1336 (N_1336,N_494,N_502);
nand U1337 (N_1337,N_295,N_726);
nand U1338 (N_1338,N_507,N_210);
nand U1339 (N_1339,N_105,N_467);
nor U1340 (N_1340,N_142,N_874);
and U1341 (N_1341,N_397,N_689);
or U1342 (N_1342,N_631,N_398);
nor U1343 (N_1343,N_658,N_464);
or U1344 (N_1344,N_768,N_340);
and U1345 (N_1345,N_331,N_234);
nor U1346 (N_1346,N_283,N_999);
and U1347 (N_1347,N_449,N_926);
or U1348 (N_1348,N_881,N_767);
nor U1349 (N_1349,N_303,N_716);
and U1350 (N_1350,N_611,N_38);
or U1351 (N_1351,N_693,N_662);
nand U1352 (N_1352,N_30,N_329);
nand U1353 (N_1353,N_974,N_911);
nor U1354 (N_1354,N_223,N_849);
and U1355 (N_1355,N_330,N_443);
nand U1356 (N_1356,N_867,N_718);
and U1357 (N_1357,N_136,N_985);
or U1358 (N_1358,N_432,N_550);
or U1359 (N_1359,N_982,N_557);
or U1360 (N_1360,N_95,N_761);
nand U1361 (N_1361,N_915,N_622);
xor U1362 (N_1362,N_819,N_921);
or U1363 (N_1363,N_970,N_59);
or U1364 (N_1364,N_942,N_232);
nand U1365 (N_1365,N_904,N_756);
or U1366 (N_1366,N_478,N_572);
or U1367 (N_1367,N_460,N_653);
or U1368 (N_1368,N_145,N_396);
or U1369 (N_1369,N_757,N_790);
or U1370 (N_1370,N_189,N_13);
or U1371 (N_1371,N_10,N_25);
and U1372 (N_1372,N_221,N_353);
or U1373 (N_1373,N_981,N_966);
nand U1374 (N_1374,N_58,N_702);
or U1375 (N_1375,N_506,N_738);
nand U1376 (N_1376,N_813,N_743);
nand U1377 (N_1377,N_679,N_871);
nand U1378 (N_1378,N_967,N_599);
or U1379 (N_1379,N_948,N_876);
nor U1380 (N_1380,N_872,N_296);
nand U1381 (N_1381,N_684,N_410);
nand U1382 (N_1382,N_896,N_742);
nor U1383 (N_1383,N_90,N_636);
and U1384 (N_1384,N_780,N_416);
nand U1385 (N_1385,N_868,N_302);
and U1386 (N_1386,N_775,N_700);
xnor U1387 (N_1387,N_423,N_422);
or U1388 (N_1388,N_804,N_163);
or U1389 (N_1389,N_118,N_411);
and U1390 (N_1390,N_72,N_581);
nand U1391 (N_1391,N_143,N_146);
and U1392 (N_1392,N_746,N_356);
or U1393 (N_1393,N_233,N_352);
and U1394 (N_1394,N_835,N_211);
nor U1395 (N_1395,N_919,N_687);
nand U1396 (N_1396,N_197,N_752);
nand U1397 (N_1397,N_669,N_797);
nor U1398 (N_1398,N_518,N_663);
or U1399 (N_1399,N_785,N_315);
nand U1400 (N_1400,N_590,N_531);
nand U1401 (N_1401,N_140,N_188);
nor U1402 (N_1402,N_363,N_243);
nand U1403 (N_1403,N_388,N_826);
nand U1404 (N_1404,N_271,N_382);
nor U1405 (N_1405,N_408,N_556);
and U1406 (N_1406,N_401,N_480);
or U1407 (N_1407,N_129,N_898);
nand U1408 (N_1408,N_986,N_957);
nor U1409 (N_1409,N_450,N_732);
nor U1410 (N_1410,N_380,N_691);
nor U1411 (N_1411,N_902,N_701);
nor U1412 (N_1412,N_588,N_56);
nor U1413 (N_1413,N_186,N_885);
nand U1414 (N_1414,N_311,N_386);
or U1415 (N_1415,N_873,N_376);
or U1416 (N_1416,N_52,N_956);
or U1417 (N_1417,N_536,N_164);
nand U1418 (N_1418,N_704,N_533);
nor U1419 (N_1419,N_224,N_372);
and U1420 (N_1420,N_575,N_644);
and U1421 (N_1421,N_171,N_387);
or U1422 (N_1422,N_76,N_517);
and U1423 (N_1423,N_711,N_638);
or U1424 (N_1424,N_245,N_215);
nor U1425 (N_1425,N_632,N_225);
xor U1426 (N_1426,N_618,N_614);
nand U1427 (N_1427,N_727,N_251);
nand U1428 (N_1428,N_882,N_92);
or U1429 (N_1429,N_8,N_512);
and U1430 (N_1430,N_51,N_579);
and U1431 (N_1431,N_440,N_499);
xor U1432 (N_1432,N_208,N_483);
nand U1433 (N_1433,N_280,N_99);
and U1434 (N_1434,N_749,N_351);
and U1435 (N_1435,N_626,N_680);
or U1436 (N_1436,N_195,N_93);
nand U1437 (N_1437,N_343,N_811);
and U1438 (N_1438,N_641,N_782);
nand U1439 (N_1439,N_22,N_2);
and U1440 (N_1440,N_230,N_445);
nand U1441 (N_1441,N_523,N_698);
or U1442 (N_1442,N_366,N_652);
or U1443 (N_1443,N_446,N_750);
nor U1444 (N_1444,N_937,N_161);
or U1445 (N_1445,N_888,N_946);
nand U1446 (N_1446,N_973,N_570);
or U1447 (N_1447,N_405,N_264);
and U1448 (N_1448,N_468,N_706);
nand U1449 (N_1449,N_989,N_800);
and U1450 (N_1450,N_848,N_413);
nor U1451 (N_1451,N_45,N_47);
nand U1452 (N_1452,N_126,N_522);
nand U1453 (N_1453,N_858,N_717);
or U1454 (N_1454,N_452,N_407);
xnor U1455 (N_1455,N_586,N_534);
nand U1456 (N_1456,N_567,N_546);
xnor U1457 (N_1457,N_648,N_865);
nand U1458 (N_1458,N_117,N_436);
nand U1459 (N_1459,N_910,N_837);
nor U1460 (N_1460,N_741,N_493);
or U1461 (N_1461,N_28,N_358);
and U1462 (N_1462,N_169,N_473);
or U1463 (N_1463,N_341,N_393);
nor U1464 (N_1464,N_854,N_477);
nor U1465 (N_1465,N_801,N_246);
nor U1466 (N_1466,N_434,N_541);
nand U1467 (N_1467,N_634,N_952);
nor U1468 (N_1468,N_350,N_913);
nor U1469 (N_1469,N_934,N_951);
and U1470 (N_1470,N_699,N_482);
and U1471 (N_1471,N_73,N_971);
and U1472 (N_1472,N_287,N_355);
or U1473 (N_1473,N_400,N_695);
nand U1474 (N_1474,N_640,N_29);
and U1475 (N_1475,N_936,N_514);
nand U1476 (N_1476,N_354,N_828);
nand U1477 (N_1477,N_977,N_789);
nand U1478 (N_1478,N_116,N_139);
nor U1479 (N_1479,N_558,N_525);
xnor U1480 (N_1480,N_134,N_972);
nor U1481 (N_1481,N_774,N_66);
or U1482 (N_1482,N_745,N_877);
nand U1483 (N_1483,N_495,N_131);
nand U1484 (N_1484,N_661,N_603);
nor U1485 (N_1485,N_442,N_192);
or U1486 (N_1486,N_799,N_206);
or U1487 (N_1487,N_239,N_992);
or U1488 (N_1488,N_841,N_125);
nand U1489 (N_1489,N_138,N_739);
and U1490 (N_1490,N_617,N_555);
nor U1491 (N_1491,N_153,N_637);
nand U1492 (N_1492,N_288,N_842);
and U1493 (N_1493,N_683,N_336);
nor U1494 (N_1494,N_427,N_149);
nor U1495 (N_1495,N_158,N_194);
nand U1496 (N_1496,N_307,N_903);
nand U1497 (N_1497,N_777,N_378);
and U1498 (N_1498,N_569,N_300);
nor U1499 (N_1499,N_594,N_472);
or U1500 (N_1500,N_474,N_578);
nor U1501 (N_1501,N_918,N_99);
nand U1502 (N_1502,N_783,N_542);
or U1503 (N_1503,N_785,N_25);
or U1504 (N_1504,N_398,N_592);
and U1505 (N_1505,N_588,N_565);
nand U1506 (N_1506,N_496,N_814);
or U1507 (N_1507,N_700,N_500);
or U1508 (N_1508,N_786,N_419);
nand U1509 (N_1509,N_167,N_894);
nand U1510 (N_1510,N_470,N_946);
nor U1511 (N_1511,N_429,N_357);
or U1512 (N_1512,N_357,N_963);
and U1513 (N_1513,N_208,N_286);
nor U1514 (N_1514,N_791,N_437);
and U1515 (N_1515,N_216,N_201);
and U1516 (N_1516,N_647,N_279);
and U1517 (N_1517,N_859,N_345);
or U1518 (N_1518,N_671,N_160);
nor U1519 (N_1519,N_289,N_429);
nor U1520 (N_1520,N_844,N_988);
nor U1521 (N_1521,N_989,N_651);
or U1522 (N_1522,N_263,N_493);
nand U1523 (N_1523,N_760,N_366);
nor U1524 (N_1524,N_944,N_205);
nor U1525 (N_1525,N_602,N_915);
xor U1526 (N_1526,N_783,N_395);
or U1527 (N_1527,N_83,N_155);
and U1528 (N_1528,N_407,N_586);
nand U1529 (N_1529,N_314,N_249);
and U1530 (N_1530,N_390,N_710);
nor U1531 (N_1531,N_399,N_699);
nor U1532 (N_1532,N_786,N_793);
nand U1533 (N_1533,N_586,N_89);
or U1534 (N_1534,N_521,N_785);
and U1535 (N_1535,N_354,N_59);
nor U1536 (N_1536,N_602,N_899);
or U1537 (N_1537,N_445,N_101);
or U1538 (N_1538,N_235,N_155);
nor U1539 (N_1539,N_80,N_288);
nand U1540 (N_1540,N_382,N_740);
nor U1541 (N_1541,N_669,N_924);
nor U1542 (N_1542,N_413,N_760);
nand U1543 (N_1543,N_934,N_812);
and U1544 (N_1544,N_264,N_388);
and U1545 (N_1545,N_314,N_487);
or U1546 (N_1546,N_811,N_385);
nand U1547 (N_1547,N_959,N_372);
nor U1548 (N_1548,N_658,N_665);
nand U1549 (N_1549,N_392,N_708);
or U1550 (N_1550,N_470,N_686);
xor U1551 (N_1551,N_290,N_111);
nand U1552 (N_1552,N_55,N_220);
nand U1553 (N_1553,N_93,N_62);
or U1554 (N_1554,N_633,N_934);
or U1555 (N_1555,N_422,N_329);
and U1556 (N_1556,N_168,N_517);
or U1557 (N_1557,N_265,N_399);
nor U1558 (N_1558,N_709,N_149);
nand U1559 (N_1559,N_673,N_78);
or U1560 (N_1560,N_287,N_935);
nor U1561 (N_1561,N_431,N_459);
or U1562 (N_1562,N_497,N_37);
or U1563 (N_1563,N_525,N_490);
nor U1564 (N_1564,N_106,N_18);
nor U1565 (N_1565,N_857,N_902);
and U1566 (N_1566,N_759,N_587);
nand U1567 (N_1567,N_69,N_767);
and U1568 (N_1568,N_485,N_530);
or U1569 (N_1569,N_553,N_307);
or U1570 (N_1570,N_813,N_60);
or U1571 (N_1571,N_378,N_18);
and U1572 (N_1572,N_597,N_183);
and U1573 (N_1573,N_994,N_310);
or U1574 (N_1574,N_526,N_827);
and U1575 (N_1575,N_582,N_126);
xnor U1576 (N_1576,N_485,N_942);
and U1577 (N_1577,N_660,N_517);
nand U1578 (N_1578,N_509,N_932);
or U1579 (N_1579,N_693,N_863);
nand U1580 (N_1580,N_472,N_675);
nor U1581 (N_1581,N_530,N_459);
nand U1582 (N_1582,N_70,N_263);
nor U1583 (N_1583,N_599,N_687);
and U1584 (N_1584,N_554,N_208);
and U1585 (N_1585,N_709,N_75);
or U1586 (N_1586,N_37,N_138);
or U1587 (N_1587,N_827,N_501);
nand U1588 (N_1588,N_969,N_925);
nor U1589 (N_1589,N_725,N_288);
or U1590 (N_1590,N_689,N_188);
nor U1591 (N_1591,N_736,N_920);
xor U1592 (N_1592,N_348,N_344);
and U1593 (N_1593,N_589,N_694);
nand U1594 (N_1594,N_673,N_629);
nor U1595 (N_1595,N_869,N_963);
and U1596 (N_1596,N_580,N_186);
and U1597 (N_1597,N_881,N_302);
nand U1598 (N_1598,N_353,N_422);
nor U1599 (N_1599,N_458,N_362);
nor U1600 (N_1600,N_365,N_22);
nor U1601 (N_1601,N_34,N_684);
nand U1602 (N_1602,N_135,N_403);
nor U1603 (N_1603,N_41,N_954);
and U1604 (N_1604,N_953,N_238);
nand U1605 (N_1605,N_62,N_119);
nor U1606 (N_1606,N_570,N_118);
nand U1607 (N_1607,N_519,N_741);
and U1608 (N_1608,N_832,N_437);
and U1609 (N_1609,N_589,N_235);
nor U1610 (N_1610,N_901,N_668);
or U1611 (N_1611,N_894,N_625);
or U1612 (N_1612,N_4,N_74);
nor U1613 (N_1613,N_788,N_179);
or U1614 (N_1614,N_891,N_452);
nand U1615 (N_1615,N_633,N_311);
and U1616 (N_1616,N_397,N_807);
nor U1617 (N_1617,N_621,N_369);
and U1618 (N_1618,N_422,N_299);
or U1619 (N_1619,N_669,N_877);
and U1620 (N_1620,N_381,N_290);
nor U1621 (N_1621,N_375,N_459);
or U1622 (N_1622,N_167,N_169);
or U1623 (N_1623,N_631,N_743);
or U1624 (N_1624,N_632,N_750);
xor U1625 (N_1625,N_576,N_581);
or U1626 (N_1626,N_945,N_312);
or U1627 (N_1627,N_922,N_852);
nand U1628 (N_1628,N_486,N_400);
nand U1629 (N_1629,N_217,N_880);
and U1630 (N_1630,N_71,N_503);
nand U1631 (N_1631,N_22,N_223);
or U1632 (N_1632,N_673,N_787);
nor U1633 (N_1633,N_251,N_157);
and U1634 (N_1634,N_960,N_945);
and U1635 (N_1635,N_744,N_56);
nor U1636 (N_1636,N_72,N_875);
or U1637 (N_1637,N_855,N_157);
or U1638 (N_1638,N_142,N_903);
or U1639 (N_1639,N_971,N_893);
nand U1640 (N_1640,N_680,N_173);
or U1641 (N_1641,N_718,N_505);
or U1642 (N_1642,N_139,N_295);
nor U1643 (N_1643,N_561,N_88);
nor U1644 (N_1644,N_680,N_341);
and U1645 (N_1645,N_11,N_846);
or U1646 (N_1646,N_419,N_239);
nand U1647 (N_1647,N_597,N_261);
and U1648 (N_1648,N_659,N_58);
and U1649 (N_1649,N_235,N_792);
or U1650 (N_1650,N_528,N_683);
and U1651 (N_1651,N_970,N_221);
nor U1652 (N_1652,N_349,N_477);
and U1653 (N_1653,N_682,N_350);
and U1654 (N_1654,N_824,N_927);
nand U1655 (N_1655,N_410,N_963);
nor U1656 (N_1656,N_706,N_827);
nor U1657 (N_1657,N_654,N_117);
nand U1658 (N_1658,N_924,N_749);
xor U1659 (N_1659,N_908,N_837);
or U1660 (N_1660,N_249,N_523);
nand U1661 (N_1661,N_295,N_815);
nor U1662 (N_1662,N_278,N_323);
or U1663 (N_1663,N_353,N_702);
nand U1664 (N_1664,N_818,N_806);
nand U1665 (N_1665,N_366,N_490);
nor U1666 (N_1666,N_280,N_408);
or U1667 (N_1667,N_846,N_642);
and U1668 (N_1668,N_534,N_536);
and U1669 (N_1669,N_471,N_235);
nand U1670 (N_1670,N_363,N_624);
and U1671 (N_1671,N_608,N_585);
nor U1672 (N_1672,N_83,N_18);
or U1673 (N_1673,N_709,N_30);
nor U1674 (N_1674,N_998,N_740);
and U1675 (N_1675,N_776,N_685);
and U1676 (N_1676,N_185,N_579);
nor U1677 (N_1677,N_590,N_538);
or U1678 (N_1678,N_329,N_166);
or U1679 (N_1679,N_876,N_674);
and U1680 (N_1680,N_589,N_289);
nand U1681 (N_1681,N_390,N_801);
nor U1682 (N_1682,N_394,N_769);
and U1683 (N_1683,N_143,N_486);
or U1684 (N_1684,N_875,N_844);
nand U1685 (N_1685,N_516,N_686);
and U1686 (N_1686,N_989,N_109);
nor U1687 (N_1687,N_557,N_498);
or U1688 (N_1688,N_854,N_856);
nand U1689 (N_1689,N_190,N_674);
nor U1690 (N_1690,N_724,N_586);
and U1691 (N_1691,N_163,N_741);
nor U1692 (N_1692,N_721,N_161);
nand U1693 (N_1693,N_10,N_329);
nand U1694 (N_1694,N_62,N_28);
nor U1695 (N_1695,N_992,N_245);
nand U1696 (N_1696,N_996,N_872);
nand U1697 (N_1697,N_423,N_119);
and U1698 (N_1698,N_47,N_507);
or U1699 (N_1699,N_559,N_528);
or U1700 (N_1700,N_73,N_734);
nor U1701 (N_1701,N_682,N_230);
nor U1702 (N_1702,N_904,N_495);
or U1703 (N_1703,N_469,N_156);
nor U1704 (N_1704,N_288,N_317);
and U1705 (N_1705,N_317,N_398);
nor U1706 (N_1706,N_332,N_632);
nor U1707 (N_1707,N_318,N_304);
nor U1708 (N_1708,N_247,N_239);
nor U1709 (N_1709,N_377,N_589);
nand U1710 (N_1710,N_213,N_774);
and U1711 (N_1711,N_180,N_223);
or U1712 (N_1712,N_845,N_263);
nor U1713 (N_1713,N_43,N_884);
xnor U1714 (N_1714,N_230,N_131);
or U1715 (N_1715,N_548,N_838);
nand U1716 (N_1716,N_519,N_910);
or U1717 (N_1717,N_496,N_151);
or U1718 (N_1718,N_77,N_812);
and U1719 (N_1719,N_402,N_786);
and U1720 (N_1720,N_599,N_296);
and U1721 (N_1721,N_431,N_366);
nor U1722 (N_1722,N_677,N_606);
and U1723 (N_1723,N_757,N_561);
or U1724 (N_1724,N_759,N_245);
nor U1725 (N_1725,N_201,N_679);
nor U1726 (N_1726,N_886,N_512);
or U1727 (N_1727,N_328,N_876);
or U1728 (N_1728,N_605,N_1);
or U1729 (N_1729,N_451,N_476);
nand U1730 (N_1730,N_286,N_523);
or U1731 (N_1731,N_904,N_466);
nor U1732 (N_1732,N_7,N_191);
and U1733 (N_1733,N_407,N_693);
and U1734 (N_1734,N_276,N_827);
or U1735 (N_1735,N_861,N_675);
and U1736 (N_1736,N_734,N_764);
nand U1737 (N_1737,N_115,N_97);
or U1738 (N_1738,N_236,N_560);
nor U1739 (N_1739,N_918,N_164);
nor U1740 (N_1740,N_798,N_241);
nand U1741 (N_1741,N_536,N_370);
or U1742 (N_1742,N_822,N_446);
or U1743 (N_1743,N_491,N_773);
and U1744 (N_1744,N_283,N_362);
nor U1745 (N_1745,N_789,N_475);
nor U1746 (N_1746,N_119,N_40);
nand U1747 (N_1747,N_656,N_835);
and U1748 (N_1748,N_179,N_580);
and U1749 (N_1749,N_673,N_495);
nor U1750 (N_1750,N_988,N_931);
or U1751 (N_1751,N_260,N_404);
and U1752 (N_1752,N_53,N_341);
nor U1753 (N_1753,N_222,N_198);
or U1754 (N_1754,N_159,N_117);
and U1755 (N_1755,N_462,N_491);
nand U1756 (N_1756,N_42,N_299);
nor U1757 (N_1757,N_101,N_525);
and U1758 (N_1758,N_829,N_52);
nand U1759 (N_1759,N_801,N_216);
and U1760 (N_1760,N_267,N_621);
and U1761 (N_1761,N_169,N_814);
nand U1762 (N_1762,N_681,N_875);
and U1763 (N_1763,N_323,N_689);
and U1764 (N_1764,N_235,N_271);
nor U1765 (N_1765,N_924,N_903);
nor U1766 (N_1766,N_108,N_505);
nor U1767 (N_1767,N_779,N_439);
nor U1768 (N_1768,N_984,N_958);
and U1769 (N_1769,N_413,N_690);
nor U1770 (N_1770,N_760,N_578);
and U1771 (N_1771,N_942,N_143);
nand U1772 (N_1772,N_557,N_899);
nor U1773 (N_1773,N_625,N_339);
or U1774 (N_1774,N_216,N_638);
nand U1775 (N_1775,N_887,N_299);
or U1776 (N_1776,N_572,N_836);
or U1777 (N_1777,N_423,N_208);
and U1778 (N_1778,N_328,N_203);
and U1779 (N_1779,N_55,N_327);
or U1780 (N_1780,N_351,N_698);
nor U1781 (N_1781,N_187,N_324);
nor U1782 (N_1782,N_589,N_842);
nand U1783 (N_1783,N_351,N_607);
xnor U1784 (N_1784,N_788,N_132);
or U1785 (N_1785,N_649,N_471);
nor U1786 (N_1786,N_253,N_70);
and U1787 (N_1787,N_867,N_636);
nor U1788 (N_1788,N_534,N_26);
nor U1789 (N_1789,N_108,N_3);
and U1790 (N_1790,N_234,N_550);
or U1791 (N_1791,N_948,N_804);
or U1792 (N_1792,N_189,N_230);
nor U1793 (N_1793,N_781,N_52);
and U1794 (N_1794,N_664,N_577);
and U1795 (N_1795,N_973,N_550);
nand U1796 (N_1796,N_596,N_637);
or U1797 (N_1797,N_284,N_807);
and U1798 (N_1798,N_974,N_955);
nor U1799 (N_1799,N_730,N_379);
or U1800 (N_1800,N_210,N_851);
and U1801 (N_1801,N_15,N_208);
or U1802 (N_1802,N_317,N_482);
nor U1803 (N_1803,N_937,N_125);
xor U1804 (N_1804,N_670,N_786);
xnor U1805 (N_1805,N_880,N_728);
and U1806 (N_1806,N_991,N_114);
and U1807 (N_1807,N_274,N_771);
and U1808 (N_1808,N_279,N_10);
xnor U1809 (N_1809,N_822,N_205);
nor U1810 (N_1810,N_161,N_563);
nand U1811 (N_1811,N_66,N_695);
and U1812 (N_1812,N_73,N_801);
nand U1813 (N_1813,N_639,N_436);
and U1814 (N_1814,N_495,N_161);
or U1815 (N_1815,N_36,N_478);
nand U1816 (N_1816,N_158,N_506);
nor U1817 (N_1817,N_44,N_99);
and U1818 (N_1818,N_205,N_207);
nand U1819 (N_1819,N_171,N_856);
or U1820 (N_1820,N_469,N_261);
or U1821 (N_1821,N_92,N_538);
and U1822 (N_1822,N_425,N_71);
and U1823 (N_1823,N_122,N_519);
nand U1824 (N_1824,N_935,N_291);
or U1825 (N_1825,N_552,N_28);
and U1826 (N_1826,N_406,N_742);
and U1827 (N_1827,N_29,N_44);
nor U1828 (N_1828,N_358,N_983);
nand U1829 (N_1829,N_602,N_30);
nand U1830 (N_1830,N_606,N_799);
or U1831 (N_1831,N_752,N_847);
or U1832 (N_1832,N_370,N_234);
nor U1833 (N_1833,N_987,N_365);
nor U1834 (N_1834,N_304,N_388);
and U1835 (N_1835,N_474,N_183);
or U1836 (N_1836,N_715,N_413);
nand U1837 (N_1837,N_944,N_640);
nand U1838 (N_1838,N_108,N_838);
nand U1839 (N_1839,N_154,N_544);
and U1840 (N_1840,N_563,N_15);
nor U1841 (N_1841,N_716,N_523);
or U1842 (N_1842,N_123,N_454);
nand U1843 (N_1843,N_679,N_652);
or U1844 (N_1844,N_130,N_886);
nor U1845 (N_1845,N_939,N_761);
and U1846 (N_1846,N_911,N_627);
or U1847 (N_1847,N_140,N_973);
nor U1848 (N_1848,N_329,N_668);
nor U1849 (N_1849,N_299,N_143);
and U1850 (N_1850,N_62,N_917);
or U1851 (N_1851,N_160,N_775);
or U1852 (N_1852,N_526,N_29);
or U1853 (N_1853,N_766,N_619);
or U1854 (N_1854,N_798,N_504);
nand U1855 (N_1855,N_619,N_71);
and U1856 (N_1856,N_820,N_214);
nor U1857 (N_1857,N_594,N_932);
nand U1858 (N_1858,N_339,N_85);
nand U1859 (N_1859,N_350,N_718);
nor U1860 (N_1860,N_643,N_628);
nor U1861 (N_1861,N_36,N_638);
or U1862 (N_1862,N_179,N_617);
nand U1863 (N_1863,N_908,N_286);
nand U1864 (N_1864,N_730,N_426);
xnor U1865 (N_1865,N_448,N_893);
and U1866 (N_1866,N_135,N_330);
and U1867 (N_1867,N_940,N_874);
nor U1868 (N_1868,N_250,N_781);
and U1869 (N_1869,N_626,N_731);
nand U1870 (N_1870,N_211,N_415);
and U1871 (N_1871,N_479,N_838);
nand U1872 (N_1872,N_871,N_281);
nand U1873 (N_1873,N_619,N_659);
nand U1874 (N_1874,N_921,N_24);
nand U1875 (N_1875,N_389,N_710);
nor U1876 (N_1876,N_370,N_856);
nor U1877 (N_1877,N_836,N_446);
or U1878 (N_1878,N_57,N_761);
nand U1879 (N_1879,N_123,N_757);
nor U1880 (N_1880,N_84,N_33);
and U1881 (N_1881,N_552,N_712);
nand U1882 (N_1882,N_55,N_664);
nand U1883 (N_1883,N_181,N_646);
or U1884 (N_1884,N_997,N_35);
and U1885 (N_1885,N_483,N_599);
nor U1886 (N_1886,N_517,N_372);
nand U1887 (N_1887,N_509,N_881);
nand U1888 (N_1888,N_809,N_550);
and U1889 (N_1889,N_913,N_223);
or U1890 (N_1890,N_740,N_795);
or U1891 (N_1891,N_209,N_842);
nor U1892 (N_1892,N_532,N_562);
or U1893 (N_1893,N_812,N_316);
or U1894 (N_1894,N_422,N_99);
nor U1895 (N_1895,N_81,N_963);
nand U1896 (N_1896,N_791,N_224);
and U1897 (N_1897,N_983,N_443);
or U1898 (N_1898,N_747,N_26);
or U1899 (N_1899,N_834,N_9);
or U1900 (N_1900,N_26,N_696);
and U1901 (N_1901,N_697,N_487);
nor U1902 (N_1902,N_390,N_384);
nor U1903 (N_1903,N_294,N_81);
nor U1904 (N_1904,N_516,N_501);
nand U1905 (N_1905,N_575,N_914);
nand U1906 (N_1906,N_681,N_407);
nand U1907 (N_1907,N_917,N_514);
nor U1908 (N_1908,N_335,N_406);
nor U1909 (N_1909,N_793,N_323);
or U1910 (N_1910,N_571,N_584);
nor U1911 (N_1911,N_594,N_695);
or U1912 (N_1912,N_603,N_879);
or U1913 (N_1913,N_59,N_85);
and U1914 (N_1914,N_520,N_480);
nor U1915 (N_1915,N_634,N_949);
and U1916 (N_1916,N_424,N_988);
nand U1917 (N_1917,N_15,N_928);
nand U1918 (N_1918,N_377,N_673);
nor U1919 (N_1919,N_900,N_572);
xor U1920 (N_1920,N_276,N_493);
and U1921 (N_1921,N_662,N_490);
and U1922 (N_1922,N_562,N_346);
nand U1923 (N_1923,N_486,N_925);
or U1924 (N_1924,N_935,N_711);
and U1925 (N_1925,N_982,N_26);
and U1926 (N_1926,N_570,N_891);
and U1927 (N_1927,N_810,N_701);
nor U1928 (N_1928,N_560,N_605);
or U1929 (N_1929,N_967,N_57);
or U1930 (N_1930,N_231,N_157);
nor U1931 (N_1931,N_405,N_946);
or U1932 (N_1932,N_102,N_288);
or U1933 (N_1933,N_143,N_952);
nor U1934 (N_1934,N_107,N_166);
nor U1935 (N_1935,N_485,N_359);
or U1936 (N_1936,N_734,N_55);
or U1937 (N_1937,N_20,N_279);
and U1938 (N_1938,N_557,N_318);
nor U1939 (N_1939,N_55,N_452);
and U1940 (N_1940,N_150,N_74);
nor U1941 (N_1941,N_397,N_521);
or U1942 (N_1942,N_213,N_184);
or U1943 (N_1943,N_282,N_783);
and U1944 (N_1944,N_632,N_282);
nand U1945 (N_1945,N_261,N_57);
and U1946 (N_1946,N_216,N_832);
nand U1947 (N_1947,N_736,N_571);
and U1948 (N_1948,N_457,N_309);
nor U1949 (N_1949,N_6,N_284);
nor U1950 (N_1950,N_431,N_553);
nand U1951 (N_1951,N_231,N_960);
xor U1952 (N_1952,N_773,N_870);
or U1953 (N_1953,N_179,N_969);
or U1954 (N_1954,N_511,N_772);
and U1955 (N_1955,N_259,N_131);
or U1956 (N_1956,N_422,N_963);
or U1957 (N_1957,N_583,N_740);
nand U1958 (N_1958,N_840,N_409);
nand U1959 (N_1959,N_868,N_446);
nor U1960 (N_1960,N_632,N_237);
xor U1961 (N_1961,N_134,N_593);
nor U1962 (N_1962,N_535,N_704);
nor U1963 (N_1963,N_43,N_758);
nand U1964 (N_1964,N_119,N_398);
or U1965 (N_1965,N_521,N_591);
nand U1966 (N_1966,N_207,N_50);
nor U1967 (N_1967,N_469,N_162);
or U1968 (N_1968,N_539,N_493);
or U1969 (N_1969,N_658,N_229);
and U1970 (N_1970,N_366,N_559);
and U1971 (N_1971,N_569,N_384);
or U1972 (N_1972,N_898,N_32);
and U1973 (N_1973,N_640,N_47);
nor U1974 (N_1974,N_306,N_291);
nor U1975 (N_1975,N_679,N_641);
and U1976 (N_1976,N_342,N_526);
nor U1977 (N_1977,N_143,N_897);
xor U1978 (N_1978,N_806,N_691);
and U1979 (N_1979,N_34,N_851);
xor U1980 (N_1980,N_132,N_154);
nor U1981 (N_1981,N_226,N_34);
or U1982 (N_1982,N_515,N_975);
or U1983 (N_1983,N_141,N_290);
and U1984 (N_1984,N_335,N_396);
or U1985 (N_1985,N_100,N_399);
or U1986 (N_1986,N_670,N_622);
or U1987 (N_1987,N_234,N_686);
nor U1988 (N_1988,N_857,N_364);
nor U1989 (N_1989,N_409,N_500);
nand U1990 (N_1990,N_441,N_267);
or U1991 (N_1991,N_698,N_665);
nor U1992 (N_1992,N_398,N_261);
and U1993 (N_1993,N_861,N_126);
and U1994 (N_1994,N_35,N_652);
nand U1995 (N_1995,N_189,N_829);
nand U1996 (N_1996,N_371,N_614);
and U1997 (N_1997,N_827,N_584);
nor U1998 (N_1998,N_492,N_417);
nand U1999 (N_1999,N_389,N_15);
or U2000 (N_2000,N_1720,N_1552);
and U2001 (N_2001,N_1220,N_1511);
or U2002 (N_2002,N_1319,N_1615);
and U2003 (N_2003,N_1087,N_1467);
and U2004 (N_2004,N_1704,N_1716);
or U2005 (N_2005,N_1415,N_1584);
nor U2006 (N_2006,N_1572,N_1287);
nor U2007 (N_2007,N_1862,N_1362);
and U2008 (N_2008,N_1192,N_1271);
or U2009 (N_2009,N_1603,N_1509);
and U2010 (N_2010,N_1128,N_1930);
or U2011 (N_2011,N_1005,N_1018);
and U2012 (N_2012,N_1682,N_1080);
and U2013 (N_2013,N_1693,N_1420);
or U2014 (N_2014,N_1184,N_1485);
or U2015 (N_2015,N_1217,N_1673);
or U2016 (N_2016,N_1946,N_1084);
nand U2017 (N_2017,N_1134,N_1886);
or U2018 (N_2018,N_1563,N_1317);
nor U2019 (N_2019,N_1487,N_1230);
nor U2020 (N_2020,N_1522,N_1195);
or U2021 (N_2021,N_1438,N_1761);
and U2022 (N_2022,N_1428,N_1390);
and U2023 (N_2023,N_1360,N_1273);
nand U2024 (N_2024,N_1719,N_1728);
and U2025 (N_2025,N_1993,N_1754);
or U2026 (N_2026,N_1674,N_1888);
and U2027 (N_2027,N_1133,N_1560);
and U2028 (N_2028,N_1729,N_1205);
or U2029 (N_2029,N_1568,N_1636);
or U2030 (N_2030,N_1666,N_1864);
nor U2031 (N_2031,N_1879,N_1002);
and U2032 (N_2032,N_1742,N_1277);
nand U2033 (N_2033,N_1710,N_1947);
or U2034 (N_2034,N_1773,N_1974);
or U2035 (N_2035,N_1508,N_1379);
nor U2036 (N_2036,N_1727,N_1743);
and U2037 (N_2037,N_1770,N_1429);
or U2038 (N_2038,N_1979,N_1178);
nand U2039 (N_2039,N_1246,N_1451);
or U2040 (N_2040,N_1296,N_1654);
nand U2041 (N_2041,N_1017,N_1997);
nor U2042 (N_2042,N_1288,N_1469);
nor U2043 (N_2043,N_1397,N_1531);
nand U2044 (N_2044,N_1374,N_1035);
or U2045 (N_2045,N_1836,N_1763);
or U2046 (N_2046,N_1818,N_1122);
nor U2047 (N_2047,N_1387,N_1493);
nand U2048 (N_2048,N_1088,N_1829);
and U2049 (N_2049,N_1593,N_1585);
nor U2050 (N_2050,N_1521,N_1067);
and U2051 (N_2051,N_1938,N_1834);
nand U2052 (N_2052,N_1648,N_1866);
nor U2053 (N_2053,N_1100,N_1331);
nor U2054 (N_2054,N_1903,N_1341);
or U2055 (N_2055,N_1305,N_1247);
and U2056 (N_2056,N_1403,N_1858);
nor U2057 (N_2057,N_1587,N_1077);
or U2058 (N_2058,N_1262,N_1882);
nor U2059 (N_2059,N_1985,N_1433);
or U2060 (N_2060,N_1984,N_1890);
or U2061 (N_2061,N_1547,N_1242);
nand U2062 (N_2062,N_1964,N_1263);
nor U2063 (N_2063,N_1426,N_1855);
nand U2064 (N_2064,N_1434,N_1109);
or U2065 (N_2065,N_1101,N_1118);
and U2066 (N_2066,N_1701,N_1012);
nand U2067 (N_2067,N_1141,N_1571);
or U2068 (N_2068,N_1057,N_1942);
nor U2069 (N_2069,N_1735,N_1611);
or U2070 (N_2070,N_1801,N_1838);
nor U2071 (N_2071,N_1145,N_1095);
or U2072 (N_2072,N_1744,N_1339);
nor U2073 (N_2073,N_1807,N_1457);
and U2074 (N_2074,N_1904,N_1896);
or U2075 (N_2075,N_1258,N_1028);
and U2076 (N_2076,N_1090,N_1776);
nand U2077 (N_2077,N_1690,N_1800);
nor U2078 (N_2078,N_1089,N_1392);
and U2079 (N_2079,N_1453,N_1958);
nor U2080 (N_2080,N_1162,N_1261);
nand U2081 (N_2081,N_1049,N_1034);
nand U2082 (N_2082,N_1638,N_1445);
or U2083 (N_2083,N_1234,N_1083);
and U2084 (N_2084,N_1169,N_1285);
and U2085 (N_2085,N_1959,N_1977);
nand U2086 (N_2086,N_1340,N_1127);
and U2087 (N_2087,N_1476,N_1675);
or U2088 (N_2088,N_1739,N_1972);
and U2089 (N_2089,N_1065,N_1950);
and U2090 (N_2090,N_1383,N_1414);
nand U2091 (N_2091,N_1146,N_1410);
and U2092 (N_2092,N_1595,N_1692);
and U2093 (N_2093,N_1185,N_1538);
and U2094 (N_2094,N_1001,N_1197);
nor U2095 (N_2095,N_1000,N_1700);
or U2096 (N_2096,N_1495,N_1062);
and U2097 (N_2097,N_1499,N_1767);
or U2098 (N_2098,N_1986,N_1021);
or U2099 (N_2099,N_1071,N_1315);
nor U2100 (N_2100,N_1981,N_1111);
and U2101 (N_2101,N_1507,N_1871);
xnor U2102 (N_2102,N_1150,N_1207);
or U2103 (N_2103,N_1074,N_1782);
or U2104 (N_2104,N_1009,N_1799);
and U2105 (N_2105,N_1458,N_1978);
nor U2106 (N_2106,N_1004,N_1789);
nand U2107 (N_2107,N_1470,N_1435);
or U2108 (N_2108,N_1644,N_1759);
and U2109 (N_2109,N_1119,N_1771);
and U2110 (N_2110,N_1527,N_1699);
nor U2111 (N_2111,N_1050,N_1618);
or U2112 (N_2112,N_1494,N_1282);
nand U2113 (N_2113,N_1885,N_1833);
nand U2114 (N_2114,N_1188,N_1766);
nand U2115 (N_2115,N_1899,N_1884);
or U2116 (N_2116,N_1738,N_1055);
and U2117 (N_2117,N_1289,N_1252);
or U2118 (N_2118,N_1955,N_1629);
or U2119 (N_2119,N_1244,N_1301);
and U2120 (N_2120,N_1819,N_1165);
or U2121 (N_2121,N_1039,N_1424);
and U2122 (N_2122,N_1350,N_1160);
xor U2123 (N_2123,N_1381,N_1279);
and U2124 (N_2124,N_1854,N_1052);
nor U2125 (N_2125,N_1321,N_1248);
nor U2126 (N_2126,N_1837,N_1411);
nor U2127 (N_2127,N_1852,N_1757);
xor U2128 (N_2128,N_1148,N_1902);
nor U2129 (N_2129,N_1781,N_1956);
and U2130 (N_2130,N_1733,N_1907);
and U2131 (N_2131,N_1877,N_1870);
and U2132 (N_2132,N_1402,N_1616);
nor U2133 (N_2133,N_1174,N_1559);
nor U2134 (N_2134,N_1219,N_1345);
and U2135 (N_2135,N_1968,N_1103);
nor U2136 (N_2136,N_1524,N_1580);
nor U2137 (N_2137,N_1689,N_1490);
or U2138 (N_2138,N_1688,N_1259);
or U2139 (N_2139,N_1928,N_1056);
and U2140 (N_2140,N_1546,N_1177);
nor U2141 (N_2141,N_1276,N_1250);
and U2142 (N_2142,N_1382,N_1681);
nand U2143 (N_2143,N_1123,N_1007);
or U2144 (N_2144,N_1971,N_1752);
xor U2145 (N_2145,N_1164,N_1224);
or U2146 (N_2146,N_1663,N_1365);
nand U2147 (N_2147,N_1199,N_1917);
and U2148 (N_2148,N_1655,N_1810);
or U2149 (N_2149,N_1008,N_1992);
or U2150 (N_2150,N_1783,N_1504);
nor U2151 (N_2151,N_1935,N_1816);
nand U2152 (N_2152,N_1714,N_1600);
or U2153 (N_2153,N_1614,N_1367);
nor U2154 (N_2154,N_1839,N_1962);
nor U2155 (N_2155,N_1751,N_1466);
nor U2156 (N_2156,N_1144,N_1375);
nand U2157 (N_2157,N_1280,N_1054);
or U2158 (N_2158,N_1577,N_1401);
nor U2159 (N_2159,N_1058,N_1172);
and U2160 (N_2160,N_1064,N_1436);
or U2161 (N_2161,N_1033,N_1266);
nor U2162 (N_2162,N_1235,N_1159);
nor U2163 (N_2163,N_1722,N_1721);
nand U2164 (N_2164,N_1606,N_1740);
or U2165 (N_2165,N_1086,N_1599);
nor U2166 (N_2166,N_1386,N_1564);
nor U2167 (N_2167,N_1389,N_1846);
and U2168 (N_2168,N_1437,N_1463);
nor U2169 (N_2169,N_1683,N_1821);
xnor U2170 (N_2170,N_1417,N_1669);
and U2171 (N_2171,N_1473,N_1677);
and U2172 (N_2172,N_1963,N_1468);
and U2173 (N_2173,N_1803,N_1501);
and U2174 (N_2174,N_1941,N_1894);
nor U2175 (N_2175,N_1910,N_1322);
or U2176 (N_2176,N_1607,N_1349);
nand U2177 (N_2177,N_1909,N_1010);
and U2178 (N_2178,N_1412,N_1787);
nor U2179 (N_2179,N_1561,N_1991);
nand U2180 (N_2180,N_1650,N_1135);
or U2181 (N_2181,N_1432,N_1358);
or U2182 (N_2182,N_1822,N_1544);
and U2183 (N_2183,N_1925,N_1982);
or U2184 (N_2184,N_1209,N_1488);
nand U2185 (N_2185,N_1645,N_1724);
and U2186 (N_2186,N_1861,N_1758);
and U2187 (N_2187,N_1059,N_1756);
nor U2188 (N_2188,N_1204,N_1863);
nand U2189 (N_2189,N_1883,N_1845);
nor U2190 (N_2190,N_1210,N_1867);
nand U2191 (N_2191,N_1260,N_1460);
nor U2192 (N_2192,N_1642,N_1193);
or U2193 (N_2193,N_1191,N_1046);
or U2194 (N_2194,N_1398,N_1915);
or U2195 (N_2195,N_1302,N_1347);
nor U2196 (N_2196,N_1656,N_1368);
nor U2197 (N_2197,N_1667,N_1170);
or U2198 (N_2198,N_1422,N_1404);
nand U2199 (N_2199,N_1328,N_1525);
or U2200 (N_2200,N_1372,N_1811);
nand U2201 (N_2201,N_1400,N_1332);
nor U2202 (N_2202,N_1036,N_1736);
or U2203 (N_2203,N_1659,N_1329);
and U2204 (N_2204,N_1407,N_1256);
nand U2205 (N_2205,N_1881,N_1900);
and U2206 (N_2206,N_1717,N_1932);
nor U2207 (N_2207,N_1019,N_1316);
or U2208 (N_2208,N_1897,N_1954);
xnor U2209 (N_2209,N_1920,N_1312);
and U2210 (N_2210,N_1214,N_1860);
or U2211 (N_2211,N_1856,N_1774);
nor U2212 (N_2212,N_1623,N_1691);
and U2213 (N_2213,N_1586,N_1254);
nor U2214 (N_2214,N_1233,N_1857);
and U2215 (N_2215,N_1944,N_1427);
or U2216 (N_2216,N_1551,N_1483);
or U2217 (N_2217,N_1226,N_1653);
nor U2218 (N_2218,N_1988,N_1706);
and U2219 (N_2219,N_1750,N_1045);
nor U2220 (N_2220,N_1377,N_1306);
nand U2221 (N_2221,N_1394,N_1069);
nand U2222 (N_2222,N_1778,N_1446);
nor U2223 (N_2223,N_1300,N_1290);
nand U2224 (N_2224,N_1835,N_1041);
nor U2225 (N_2225,N_1269,N_1530);
and U2226 (N_2226,N_1622,N_1698);
nand U2227 (N_2227,N_1576,N_1718);
nand U2228 (N_2228,N_1557,N_1303);
and U2229 (N_2229,N_1536,N_1047);
or U2230 (N_2230,N_1384,N_1694);
or U2231 (N_2231,N_1307,N_1697);
nor U2232 (N_2232,N_1393,N_1117);
or U2233 (N_2233,N_1548,N_1291);
or U2234 (N_2234,N_1628,N_1765);
nor U2235 (N_2235,N_1933,N_1926);
or U2236 (N_2236,N_1042,N_1106);
xnor U2237 (N_2237,N_1936,N_1541);
or U2238 (N_2238,N_1450,N_1474);
and U2239 (N_2239,N_1558,N_1980);
nor U2240 (N_2240,N_1640,N_1998);
nor U2241 (N_2241,N_1486,N_1519);
nand U2242 (N_2242,N_1156,N_1797);
or U2243 (N_2243,N_1634,N_1173);
and U2244 (N_2244,N_1566,N_1874);
nor U2245 (N_2245,N_1887,N_1796);
nand U2246 (N_2246,N_1131,N_1939);
and U2247 (N_2247,N_1327,N_1705);
nand U2248 (N_2248,N_1355,N_1597);
or U2249 (N_2249,N_1180,N_1196);
or U2250 (N_2250,N_1989,N_1092);
nand U2251 (N_2251,N_1299,N_1533);
or U2252 (N_2252,N_1503,N_1832);
nand U2253 (N_2253,N_1711,N_1575);
nand U2254 (N_2254,N_1155,N_1598);
nor U2255 (N_2255,N_1114,N_1702);
nand U2256 (N_2256,N_1555,N_1421);
and U2257 (N_2257,N_1996,N_1684);
nor U2258 (N_2258,N_1658,N_1831);
nor U2259 (N_2259,N_1218,N_1625);
and U2260 (N_2260,N_1308,N_1070);
nor U2261 (N_2261,N_1462,N_1513);
or U2262 (N_2262,N_1491,N_1713);
xor U2263 (N_2263,N_1409,N_1051);
and U2264 (N_2264,N_1278,N_1171);
nand U2265 (N_2265,N_1583,N_1512);
or U2266 (N_2266,N_1072,N_1413);
nand U2267 (N_2267,N_1613,N_1608);
and U2268 (N_2268,N_1784,N_1430);
or U2269 (N_2269,N_1082,N_1573);
or U2270 (N_2270,N_1353,N_1708);
or U2271 (N_2271,N_1594,N_1553);
and U2272 (N_2272,N_1528,N_1651);
xnor U2273 (N_2273,N_1755,N_1342);
or U2274 (N_2274,N_1543,N_1175);
or U2275 (N_2275,N_1239,N_1138);
nand U2276 (N_2276,N_1610,N_1994);
nand U2277 (N_2277,N_1779,N_1027);
or U2278 (N_2278,N_1823,N_1324);
nand U2279 (N_2279,N_1359,N_1022);
and U2280 (N_2280,N_1805,N_1186);
and U2281 (N_2281,N_1023,N_1380);
and U2282 (N_2282,N_1652,N_1777);
nand U2283 (N_2283,N_1813,N_1356);
nand U2284 (N_2284,N_1228,N_1880);
or U2285 (N_2285,N_1116,N_1085);
nand U2286 (N_2286,N_1630,N_1498);
nand U2287 (N_2287,N_1662,N_1147);
and U2288 (N_2288,N_1927,N_1098);
nor U2289 (N_2289,N_1514,N_1987);
and U2290 (N_2290,N_1253,N_1703);
or U2291 (N_2291,N_1102,N_1323);
and U2292 (N_2292,N_1951,N_1515);
nand U2293 (N_2293,N_1672,N_1040);
nor U2294 (N_2294,N_1802,N_1901);
or U2295 (N_2295,N_1820,N_1922);
nand U2296 (N_2296,N_1746,N_1304);
and U2297 (N_2297,N_1479,N_1747);
or U2298 (N_2298,N_1416,N_1053);
or U2299 (N_2299,N_1913,N_1107);
or U2300 (N_2300,N_1668,N_1431);
nor U2301 (N_2301,N_1827,N_1297);
nor U2302 (N_2302,N_1764,N_1167);
xor U2303 (N_2303,N_1824,N_1310);
and U2304 (N_2304,N_1960,N_1320);
nor U2305 (N_2305,N_1068,N_1908);
or U2306 (N_2306,N_1461,N_1352);
and U2307 (N_2307,N_1791,N_1423);
nor U2308 (N_2308,N_1931,N_1136);
nand U2309 (N_2309,N_1670,N_1617);
xor U2310 (N_2310,N_1482,N_1200);
nor U2311 (N_2311,N_1646,N_1198);
nor U2312 (N_2312,N_1181,N_1545);
nand U2313 (N_2313,N_1293,N_1361);
or U2314 (N_2314,N_1337,N_1325);
and U2315 (N_2315,N_1274,N_1484);
nand U2316 (N_2316,N_1370,N_1723);
nor U2317 (N_2317,N_1741,N_1549);
nor U2318 (N_2318,N_1853,N_1505);
and U2319 (N_2319,N_1369,N_1604);
nand U2320 (N_2320,N_1840,N_1825);
or U2321 (N_2321,N_1183,N_1364);
and U2322 (N_2322,N_1808,N_1357);
and U2323 (N_2323,N_1194,N_1179);
nand U2324 (N_2324,N_1227,N_1343);
nor U2325 (N_2325,N_1612,N_1999);
nor U2326 (N_2326,N_1455,N_1680);
nor U2327 (N_2327,N_1591,N_1649);
nor U2328 (N_2328,N_1556,N_1624);
and U2329 (N_2329,N_1500,N_1581);
nand U2330 (N_2330,N_1489,N_1024);
and U2331 (N_2331,N_1665,N_1385);
nand U2332 (N_2332,N_1471,N_1526);
nor U2333 (N_2333,N_1295,N_1121);
nor U2334 (N_2334,N_1578,N_1523);
nand U2335 (N_2335,N_1872,N_1182);
nand U2336 (N_2336,N_1454,N_1923);
or U2337 (N_2337,N_1081,N_1775);
nand U2338 (N_2338,N_1934,N_1211);
or U2339 (N_2339,N_1075,N_1443);
or U2340 (N_2340,N_1678,N_1094);
or U2341 (N_2341,N_1129,N_1590);
and U2342 (N_2342,N_1709,N_1730);
xnor U2343 (N_2343,N_1213,N_1497);
and U2344 (N_2344,N_1143,N_1025);
and U2345 (N_2345,N_1333,N_1240);
nor U2346 (N_2346,N_1264,N_1496);
nand U2347 (N_2347,N_1091,N_1238);
nand U2348 (N_2348,N_1298,N_1158);
and U2349 (N_2349,N_1124,N_1110);
nor U2350 (N_2350,N_1952,N_1208);
nor U2351 (N_2351,N_1187,N_1848);
or U2352 (N_2352,N_1283,N_1793);
and U2353 (N_2353,N_1875,N_1762);
nor U2354 (N_2354,N_1176,N_1976);
nand U2355 (N_2355,N_1570,N_1395);
and U2356 (N_2356,N_1929,N_1973);
or U2357 (N_2357,N_1995,N_1620);
nor U2358 (N_2358,N_1786,N_1626);
nor U2359 (N_2359,N_1236,N_1265);
nor U2360 (N_2360,N_1229,N_1679);
nand U2361 (N_2361,N_1945,N_1037);
and U2362 (N_2362,N_1419,N_1806);
nor U2363 (N_2363,N_1975,N_1970);
nand U2364 (N_2364,N_1869,N_1532);
and U2365 (N_2365,N_1865,N_1804);
nor U2366 (N_2366,N_1452,N_1949);
nand U2367 (N_2367,N_1520,N_1873);
nor U2368 (N_2368,N_1707,N_1516);
or U2369 (N_2369,N_1475,N_1275);
and U2370 (N_2370,N_1480,N_1567);
and U2371 (N_2371,N_1647,N_1030);
and U2372 (N_2372,N_1911,N_1366);
nand U2373 (N_2373,N_1753,N_1163);
and U2374 (N_2374,N_1592,N_1768);
or U2375 (N_2375,N_1812,N_1011);
nor U2376 (N_2376,N_1660,N_1565);
nand U2377 (N_2377,N_1554,N_1601);
nand U2378 (N_2378,N_1602,N_1061);
or U2379 (N_2379,N_1940,N_1363);
or U2380 (N_2380,N_1579,N_1769);
or U2381 (N_2381,N_1937,N_1957);
nand U2382 (N_2382,N_1044,N_1948);
or U2383 (N_2383,N_1732,N_1425);
or U2384 (N_2384,N_1225,N_1168);
xor U2385 (N_2385,N_1893,N_1965);
nor U2386 (N_2386,N_1686,N_1916);
or U2387 (N_2387,N_1311,N_1715);
nor U2388 (N_2388,N_1898,N_1760);
or U2389 (N_2389,N_1631,N_1841);
nor U2390 (N_2390,N_1267,N_1335);
or U2391 (N_2391,N_1780,N_1843);
or U2392 (N_2392,N_1309,N_1478);
nand U2393 (N_2393,N_1657,N_1126);
nor U2394 (N_2394,N_1232,N_1859);
nand U2395 (N_2395,N_1222,N_1596);
nor U2396 (N_2396,N_1517,N_1712);
nand U2397 (N_2397,N_1346,N_1063);
or U2398 (N_2398,N_1849,N_1099);
and U2399 (N_2399,N_1790,N_1286);
or U2400 (N_2400,N_1635,N_1073);
nand U2401 (N_2401,N_1826,N_1272);
or U2402 (N_2402,N_1731,N_1270);
and U2403 (N_2403,N_1231,N_1815);
or U2404 (N_2404,N_1969,N_1621);
nor U2405 (N_2405,N_1465,N_1078);
nand U2406 (N_2406,N_1619,N_1223);
or U2407 (N_2407,N_1444,N_1016);
nand U2408 (N_2408,N_1396,N_1060);
and U2409 (N_2409,N_1878,N_1202);
and U2410 (N_2410,N_1892,N_1048);
and U2411 (N_2411,N_1643,N_1405);
nand U2412 (N_2412,N_1842,N_1664);
or U2413 (N_2413,N_1149,N_1237);
nand U2414 (N_2414,N_1013,N_1535);
or U2415 (N_2415,N_1391,N_1464);
xnor U2416 (N_2416,N_1502,N_1919);
xor U2417 (N_2417,N_1026,N_1406);
nand U2418 (N_2418,N_1518,N_1772);
nor U2419 (N_2419,N_1967,N_1685);
or U2420 (N_2420,N_1540,N_1850);
xnor U2421 (N_2421,N_1953,N_1550);
nor U2422 (N_2422,N_1216,N_1157);
or U2423 (N_2423,N_1140,N_1921);
and U2424 (N_2424,N_1354,N_1661);
or U2425 (N_2425,N_1506,N_1448);
or U2426 (N_2426,N_1043,N_1924);
or U2427 (N_2427,N_1817,N_1847);
nand U2428 (N_2428,N_1142,N_1990);
nand U2429 (N_2429,N_1785,N_1492);
or U2430 (N_2430,N_1113,N_1441);
nand U2431 (N_2431,N_1137,N_1014);
nand U2432 (N_2432,N_1459,N_1809);
nor U2433 (N_2433,N_1828,N_1268);
nor U2434 (N_2434,N_1189,N_1221);
nand U2435 (N_2435,N_1130,N_1408);
nand U2436 (N_2436,N_1108,N_1726);
or U2437 (N_2437,N_1418,N_1895);
nor U2438 (N_2438,N_1243,N_1257);
and U2439 (N_2439,N_1203,N_1868);
or U2440 (N_2440,N_1294,N_1605);
or U2441 (N_2441,N_1112,N_1079);
nor U2442 (N_2442,N_1093,N_1115);
and U2443 (N_2443,N_1206,N_1912);
nor U2444 (N_2444,N_1687,N_1439);
and U2445 (N_2445,N_1249,N_1748);
nand U2446 (N_2446,N_1166,N_1695);
or U2447 (N_2447,N_1537,N_1914);
nand U2448 (N_2448,N_1348,N_1440);
or U2449 (N_2449,N_1830,N_1152);
and U2450 (N_2450,N_1006,N_1639);
and U2451 (N_2451,N_1105,N_1003);
nand U2452 (N_2452,N_1966,N_1031);
nand U2453 (N_2453,N_1338,N_1139);
and U2454 (N_2454,N_1632,N_1529);
nor U2455 (N_2455,N_1905,N_1983);
nand U2456 (N_2456,N_1097,N_1794);
and U2457 (N_2457,N_1943,N_1589);
and U2458 (N_2458,N_1313,N_1745);
nand U2459 (N_2459,N_1734,N_1344);
xnor U2460 (N_2460,N_1334,N_1671);
nor U2461 (N_2461,N_1190,N_1676);
nand U2462 (N_2462,N_1038,N_1637);
nand U2463 (N_2463,N_1918,N_1889);
nand U2464 (N_2464,N_1281,N_1542);
nor U2465 (N_2465,N_1373,N_1201);
xnor U2466 (N_2466,N_1104,N_1245);
nand U2467 (N_2467,N_1376,N_1456);
nand U2468 (N_2468,N_1292,N_1442);
nand U2469 (N_2469,N_1569,N_1020);
nor U2470 (N_2470,N_1153,N_1284);
and U2471 (N_2471,N_1609,N_1961);
or U2472 (N_2472,N_1151,N_1330);
nand U2473 (N_2473,N_1212,N_1627);
and U2474 (N_2474,N_1472,N_1795);
nor U2475 (N_2475,N_1633,N_1029);
nor U2476 (N_2476,N_1582,N_1539);
nor U2477 (N_2477,N_1725,N_1326);
and U2478 (N_2478,N_1066,N_1255);
and U2479 (N_2479,N_1096,N_1574);
and U2480 (N_2480,N_1314,N_1562);
and U2481 (N_2481,N_1477,N_1481);
nand U2482 (N_2482,N_1318,N_1588);
nand U2483 (N_2483,N_1125,N_1534);
and U2484 (N_2484,N_1015,N_1851);
nor U2485 (N_2485,N_1891,N_1120);
nand U2486 (N_2486,N_1696,N_1351);
or U2487 (N_2487,N_1076,N_1749);
and U2488 (N_2488,N_1641,N_1032);
nor U2489 (N_2489,N_1132,N_1906);
and U2490 (N_2490,N_1371,N_1844);
nand U2491 (N_2491,N_1161,N_1449);
or U2492 (N_2492,N_1447,N_1792);
xor U2493 (N_2493,N_1388,N_1737);
or U2494 (N_2494,N_1788,N_1251);
nand U2495 (N_2495,N_1399,N_1510);
nor U2496 (N_2496,N_1798,N_1154);
nor U2497 (N_2497,N_1241,N_1876);
nand U2498 (N_2498,N_1215,N_1378);
nor U2499 (N_2499,N_1336,N_1814);
xor U2500 (N_2500,N_1332,N_1518);
and U2501 (N_2501,N_1767,N_1034);
nor U2502 (N_2502,N_1264,N_1563);
nand U2503 (N_2503,N_1708,N_1983);
and U2504 (N_2504,N_1417,N_1269);
or U2505 (N_2505,N_1708,N_1502);
nor U2506 (N_2506,N_1814,N_1500);
and U2507 (N_2507,N_1274,N_1731);
and U2508 (N_2508,N_1813,N_1319);
and U2509 (N_2509,N_1328,N_1217);
nand U2510 (N_2510,N_1907,N_1688);
and U2511 (N_2511,N_1955,N_1863);
or U2512 (N_2512,N_1191,N_1115);
and U2513 (N_2513,N_1731,N_1909);
and U2514 (N_2514,N_1151,N_1919);
nor U2515 (N_2515,N_1223,N_1072);
and U2516 (N_2516,N_1255,N_1983);
or U2517 (N_2517,N_1623,N_1099);
or U2518 (N_2518,N_1250,N_1151);
nand U2519 (N_2519,N_1288,N_1714);
nor U2520 (N_2520,N_1778,N_1426);
and U2521 (N_2521,N_1368,N_1564);
or U2522 (N_2522,N_1899,N_1977);
and U2523 (N_2523,N_1051,N_1641);
and U2524 (N_2524,N_1271,N_1278);
xor U2525 (N_2525,N_1528,N_1439);
nor U2526 (N_2526,N_1970,N_1335);
nand U2527 (N_2527,N_1613,N_1006);
nand U2528 (N_2528,N_1044,N_1576);
and U2529 (N_2529,N_1688,N_1374);
nor U2530 (N_2530,N_1482,N_1640);
nand U2531 (N_2531,N_1536,N_1270);
nor U2532 (N_2532,N_1582,N_1124);
or U2533 (N_2533,N_1124,N_1566);
xor U2534 (N_2534,N_1435,N_1209);
and U2535 (N_2535,N_1324,N_1914);
or U2536 (N_2536,N_1392,N_1963);
and U2537 (N_2537,N_1077,N_1691);
and U2538 (N_2538,N_1549,N_1381);
nor U2539 (N_2539,N_1083,N_1091);
and U2540 (N_2540,N_1698,N_1082);
nand U2541 (N_2541,N_1565,N_1771);
nor U2542 (N_2542,N_1084,N_1350);
and U2543 (N_2543,N_1129,N_1840);
or U2544 (N_2544,N_1181,N_1492);
nand U2545 (N_2545,N_1921,N_1440);
xor U2546 (N_2546,N_1513,N_1010);
xnor U2547 (N_2547,N_1202,N_1300);
or U2548 (N_2548,N_1857,N_1434);
and U2549 (N_2549,N_1130,N_1596);
nor U2550 (N_2550,N_1243,N_1502);
nor U2551 (N_2551,N_1751,N_1947);
and U2552 (N_2552,N_1522,N_1667);
nor U2553 (N_2553,N_1443,N_1490);
or U2554 (N_2554,N_1236,N_1477);
nor U2555 (N_2555,N_1957,N_1110);
nor U2556 (N_2556,N_1832,N_1377);
nor U2557 (N_2557,N_1331,N_1024);
nand U2558 (N_2558,N_1263,N_1732);
and U2559 (N_2559,N_1608,N_1876);
and U2560 (N_2560,N_1705,N_1218);
nor U2561 (N_2561,N_1192,N_1098);
or U2562 (N_2562,N_1382,N_1187);
and U2563 (N_2563,N_1291,N_1287);
nand U2564 (N_2564,N_1742,N_1051);
and U2565 (N_2565,N_1746,N_1677);
or U2566 (N_2566,N_1840,N_1218);
nand U2567 (N_2567,N_1110,N_1359);
nand U2568 (N_2568,N_1078,N_1501);
nand U2569 (N_2569,N_1238,N_1665);
nor U2570 (N_2570,N_1075,N_1335);
or U2571 (N_2571,N_1313,N_1551);
nor U2572 (N_2572,N_1575,N_1142);
nand U2573 (N_2573,N_1017,N_1524);
nand U2574 (N_2574,N_1794,N_1791);
and U2575 (N_2575,N_1220,N_1606);
nand U2576 (N_2576,N_1341,N_1093);
or U2577 (N_2577,N_1513,N_1023);
nand U2578 (N_2578,N_1559,N_1953);
and U2579 (N_2579,N_1517,N_1335);
nor U2580 (N_2580,N_1854,N_1522);
nor U2581 (N_2581,N_1979,N_1596);
nor U2582 (N_2582,N_1106,N_1905);
nor U2583 (N_2583,N_1875,N_1805);
nor U2584 (N_2584,N_1320,N_1023);
nor U2585 (N_2585,N_1261,N_1349);
or U2586 (N_2586,N_1902,N_1336);
and U2587 (N_2587,N_1792,N_1035);
or U2588 (N_2588,N_1630,N_1890);
and U2589 (N_2589,N_1891,N_1321);
nor U2590 (N_2590,N_1470,N_1263);
or U2591 (N_2591,N_1204,N_1208);
or U2592 (N_2592,N_1997,N_1470);
xor U2593 (N_2593,N_1595,N_1693);
nor U2594 (N_2594,N_1457,N_1391);
or U2595 (N_2595,N_1906,N_1095);
nor U2596 (N_2596,N_1411,N_1634);
xor U2597 (N_2597,N_1111,N_1524);
nand U2598 (N_2598,N_1368,N_1261);
nand U2599 (N_2599,N_1648,N_1047);
nand U2600 (N_2600,N_1845,N_1533);
nor U2601 (N_2601,N_1066,N_1173);
nand U2602 (N_2602,N_1994,N_1753);
nand U2603 (N_2603,N_1386,N_1488);
or U2604 (N_2604,N_1299,N_1931);
and U2605 (N_2605,N_1666,N_1748);
and U2606 (N_2606,N_1136,N_1972);
and U2607 (N_2607,N_1384,N_1630);
nor U2608 (N_2608,N_1682,N_1690);
nand U2609 (N_2609,N_1124,N_1422);
nor U2610 (N_2610,N_1060,N_1508);
nor U2611 (N_2611,N_1511,N_1141);
or U2612 (N_2612,N_1869,N_1458);
or U2613 (N_2613,N_1216,N_1337);
nor U2614 (N_2614,N_1191,N_1693);
and U2615 (N_2615,N_1824,N_1816);
and U2616 (N_2616,N_1584,N_1350);
nor U2617 (N_2617,N_1772,N_1264);
nor U2618 (N_2618,N_1076,N_1570);
and U2619 (N_2619,N_1395,N_1268);
and U2620 (N_2620,N_1270,N_1758);
nand U2621 (N_2621,N_1114,N_1808);
and U2622 (N_2622,N_1275,N_1391);
nand U2623 (N_2623,N_1533,N_1557);
nor U2624 (N_2624,N_1380,N_1033);
xnor U2625 (N_2625,N_1824,N_1716);
nor U2626 (N_2626,N_1448,N_1781);
nand U2627 (N_2627,N_1421,N_1837);
xnor U2628 (N_2628,N_1950,N_1457);
nor U2629 (N_2629,N_1272,N_1592);
nor U2630 (N_2630,N_1592,N_1917);
and U2631 (N_2631,N_1000,N_1718);
or U2632 (N_2632,N_1576,N_1666);
nand U2633 (N_2633,N_1647,N_1768);
or U2634 (N_2634,N_1681,N_1062);
or U2635 (N_2635,N_1971,N_1390);
nand U2636 (N_2636,N_1429,N_1581);
nor U2637 (N_2637,N_1745,N_1991);
xor U2638 (N_2638,N_1797,N_1245);
or U2639 (N_2639,N_1698,N_1863);
nor U2640 (N_2640,N_1112,N_1054);
nor U2641 (N_2641,N_1113,N_1152);
or U2642 (N_2642,N_1781,N_1916);
nor U2643 (N_2643,N_1828,N_1826);
nand U2644 (N_2644,N_1522,N_1366);
and U2645 (N_2645,N_1459,N_1906);
and U2646 (N_2646,N_1166,N_1767);
and U2647 (N_2647,N_1119,N_1068);
and U2648 (N_2648,N_1492,N_1920);
xor U2649 (N_2649,N_1523,N_1120);
nand U2650 (N_2650,N_1756,N_1610);
and U2651 (N_2651,N_1726,N_1620);
nor U2652 (N_2652,N_1665,N_1440);
and U2653 (N_2653,N_1642,N_1482);
or U2654 (N_2654,N_1911,N_1305);
and U2655 (N_2655,N_1608,N_1094);
or U2656 (N_2656,N_1027,N_1920);
or U2657 (N_2657,N_1836,N_1129);
or U2658 (N_2658,N_1752,N_1410);
nand U2659 (N_2659,N_1935,N_1107);
nand U2660 (N_2660,N_1595,N_1218);
and U2661 (N_2661,N_1743,N_1730);
nand U2662 (N_2662,N_1504,N_1192);
and U2663 (N_2663,N_1870,N_1560);
and U2664 (N_2664,N_1962,N_1419);
and U2665 (N_2665,N_1098,N_1901);
nor U2666 (N_2666,N_1311,N_1710);
nand U2667 (N_2667,N_1924,N_1234);
nand U2668 (N_2668,N_1904,N_1456);
nor U2669 (N_2669,N_1456,N_1678);
nor U2670 (N_2670,N_1112,N_1206);
nand U2671 (N_2671,N_1255,N_1126);
and U2672 (N_2672,N_1686,N_1407);
and U2673 (N_2673,N_1852,N_1088);
or U2674 (N_2674,N_1622,N_1957);
or U2675 (N_2675,N_1148,N_1843);
and U2676 (N_2676,N_1655,N_1633);
and U2677 (N_2677,N_1001,N_1209);
nand U2678 (N_2678,N_1955,N_1378);
nor U2679 (N_2679,N_1838,N_1150);
nor U2680 (N_2680,N_1611,N_1336);
nor U2681 (N_2681,N_1296,N_1720);
nor U2682 (N_2682,N_1352,N_1746);
or U2683 (N_2683,N_1493,N_1029);
nand U2684 (N_2684,N_1207,N_1293);
nand U2685 (N_2685,N_1775,N_1038);
or U2686 (N_2686,N_1229,N_1736);
nor U2687 (N_2687,N_1453,N_1639);
and U2688 (N_2688,N_1270,N_1601);
nand U2689 (N_2689,N_1704,N_1719);
and U2690 (N_2690,N_1834,N_1962);
or U2691 (N_2691,N_1661,N_1634);
nand U2692 (N_2692,N_1786,N_1920);
nand U2693 (N_2693,N_1828,N_1118);
and U2694 (N_2694,N_1340,N_1207);
nand U2695 (N_2695,N_1069,N_1868);
nand U2696 (N_2696,N_1216,N_1591);
nor U2697 (N_2697,N_1214,N_1007);
and U2698 (N_2698,N_1417,N_1951);
nand U2699 (N_2699,N_1718,N_1956);
and U2700 (N_2700,N_1401,N_1750);
or U2701 (N_2701,N_1129,N_1101);
nand U2702 (N_2702,N_1629,N_1178);
or U2703 (N_2703,N_1530,N_1792);
nor U2704 (N_2704,N_1807,N_1798);
nor U2705 (N_2705,N_1211,N_1009);
and U2706 (N_2706,N_1876,N_1294);
or U2707 (N_2707,N_1552,N_1705);
and U2708 (N_2708,N_1607,N_1402);
nor U2709 (N_2709,N_1302,N_1686);
nand U2710 (N_2710,N_1018,N_1188);
or U2711 (N_2711,N_1489,N_1219);
and U2712 (N_2712,N_1523,N_1700);
nor U2713 (N_2713,N_1308,N_1598);
or U2714 (N_2714,N_1352,N_1549);
or U2715 (N_2715,N_1954,N_1652);
and U2716 (N_2716,N_1604,N_1794);
or U2717 (N_2717,N_1800,N_1909);
nor U2718 (N_2718,N_1650,N_1943);
nor U2719 (N_2719,N_1693,N_1944);
or U2720 (N_2720,N_1894,N_1182);
or U2721 (N_2721,N_1953,N_1893);
or U2722 (N_2722,N_1003,N_1442);
or U2723 (N_2723,N_1969,N_1439);
and U2724 (N_2724,N_1771,N_1818);
or U2725 (N_2725,N_1332,N_1306);
or U2726 (N_2726,N_1649,N_1655);
or U2727 (N_2727,N_1750,N_1478);
nand U2728 (N_2728,N_1848,N_1671);
nand U2729 (N_2729,N_1237,N_1463);
xnor U2730 (N_2730,N_1943,N_1378);
nor U2731 (N_2731,N_1949,N_1578);
or U2732 (N_2732,N_1931,N_1449);
nor U2733 (N_2733,N_1995,N_1395);
nand U2734 (N_2734,N_1478,N_1738);
nand U2735 (N_2735,N_1616,N_1134);
and U2736 (N_2736,N_1553,N_1747);
and U2737 (N_2737,N_1778,N_1976);
nor U2738 (N_2738,N_1877,N_1284);
nand U2739 (N_2739,N_1168,N_1673);
nand U2740 (N_2740,N_1213,N_1609);
nor U2741 (N_2741,N_1768,N_1116);
and U2742 (N_2742,N_1715,N_1211);
nand U2743 (N_2743,N_1271,N_1041);
nor U2744 (N_2744,N_1569,N_1000);
nand U2745 (N_2745,N_1818,N_1057);
nor U2746 (N_2746,N_1560,N_1556);
nand U2747 (N_2747,N_1130,N_1797);
and U2748 (N_2748,N_1528,N_1359);
and U2749 (N_2749,N_1369,N_1352);
nand U2750 (N_2750,N_1880,N_1830);
xor U2751 (N_2751,N_1807,N_1114);
nor U2752 (N_2752,N_1821,N_1718);
nand U2753 (N_2753,N_1235,N_1738);
and U2754 (N_2754,N_1884,N_1243);
and U2755 (N_2755,N_1672,N_1419);
nand U2756 (N_2756,N_1838,N_1466);
and U2757 (N_2757,N_1209,N_1433);
nand U2758 (N_2758,N_1911,N_1913);
or U2759 (N_2759,N_1755,N_1540);
and U2760 (N_2760,N_1266,N_1678);
nor U2761 (N_2761,N_1720,N_1619);
nand U2762 (N_2762,N_1525,N_1994);
or U2763 (N_2763,N_1711,N_1966);
or U2764 (N_2764,N_1762,N_1689);
and U2765 (N_2765,N_1791,N_1440);
nand U2766 (N_2766,N_1913,N_1822);
nand U2767 (N_2767,N_1671,N_1720);
nor U2768 (N_2768,N_1495,N_1004);
nand U2769 (N_2769,N_1339,N_1020);
xnor U2770 (N_2770,N_1788,N_1402);
nor U2771 (N_2771,N_1513,N_1022);
and U2772 (N_2772,N_1304,N_1382);
or U2773 (N_2773,N_1483,N_1407);
nor U2774 (N_2774,N_1874,N_1216);
nand U2775 (N_2775,N_1932,N_1867);
and U2776 (N_2776,N_1468,N_1234);
or U2777 (N_2777,N_1049,N_1704);
and U2778 (N_2778,N_1234,N_1481);
and U2779 (N_2779,N_1530,N_1962);
nor U2780 (N_2780,N_1222,N_1084);
nor U2781 (N_2781,N_1741,N_1384);
and U2782 (N_2782,N_1281,N_1940);
nor U2783 (N_2783,N_1037,N_1637);
nand U2784 (N_2784,N_1160,N_1909);
or U2785 (N_2785,N_1492,N_1552);
or U2786 (N_2786,N_1788,N_1645);
and U2787 (N_2787,N_1486,N_1084);
and U2788 (N_2788,N_1156,N_1096);
xor U2789 (N_2789,N_1611,N_1058);
or U2790 (N_2790,N_1809,N_1835);
nand U2791 (N_2791,N_1844,N_1597);
nor U2792 (N_2792,N_1172,N_1537);
nand U2793 (N_2793,N_1754,N_1400);
xnor U2794 (N_2794,N_1018,N_1958);
and U2795 (N_2795,N_1895,N_1062);
nor U2796 (N_2796,N_1188,N_1232);
nand U2797 (N_2797,N_1313,N_1441);
nand U2798 (N_2798,N_1500,N_1005);
nand U2799 (N_2799,N_1239,N_1365);
nor U2800 (N_2800,N_1291,N_1038);
and U2801 (N_2801,N_1315,N_1091);
or U2802 (N_2802,N_1276,N_1500);
nor U2803 (N_2803,N_1372,N_1384);
nand U2804 (N_2804,N_1753,N_1649);
nor U2805 (N_2805,N_1532,N_1797);
or U2806 (N_2806,N_1310,N_1815);
and U2807 (N_2807,N_1573,N_1299);
nor U2808 (N_2808,N_1186,N_1732);
or U2809 (N_2809,N_1746,N_1088);
and U2810 (N_2810,N_1880,N_1431);
and U2811 (N_2811,N_1116,N_1123);
and U2812 (N_2812,N_1513,N_1331);
nor U2813 (N_2813,N_1984,N_1086);
or U2814 (N_2814,N_1894,N_1102);
nand U2815 (N_2815,N_1205,N_1696);
nor U2816 (N_2816,N_1744,N_1561);
nand U2817 (N_2817,N_1677,N_1038);
and U2818 (N_2818,N_1595,N_1520);
and U2819 (N_2819,N_1655,N_1501);
or U2820 (N_2820,N_1616,N_1489);
nand U2821 (N_2821,N_1475,N_1481);
and U2822 (N_2822,N_1725,N_1144);
nor U2823 (N_2823,N_1847,N_1891);
nor U2824 (N_2824,N_1784,N_1578);
nand U2825 (N_2825,N_1835,N_1444);
and U2826 (N_2826,N_1438,N_1836);
or U2827 (N_2827,N_1862,N_1143);
nor U2828 (N_2828,N_1386,N_1271);
or U2829 (N_2829,N_1185,N_1358);
and U2830 (N_2830,N_1207,N_1818);
nand U2831 (N_2831,N_1927,N_1060);
nand U2832 (N_2832,N_1807,N_1500);
and U2833 (N_2833,N_1558,N_1855);
and U2834 (N_2834,N_1704,N_1068);
xor U2835 (N_2835,N_1443,N_1227);
and U2836 (N_2836,N_1305,N_1778);
nand U2837 (N_2837,N_1353,N_1964);
nor U2838 (N_2838,N_1609,N_1292);
and U2839 (N_2839,N_1511,N_1209);
and U2840 (N_2840,N_1734,N_1487);
nor U2841 (N_2841,N_1925,N_1515);
and U2842 (N_2842,N_1026,N_1131);
and U2843 (N_2843,N_1625,N_1765);
nor U2844 (N_2844,N_1981,N_1316);
and U2845 (N_2845,N_1290,N_1738);
nand U2846 (N_2846,N_1910,N_1384);
and U2847 (N_2847,N_1711,N_1946);
nand U2848 (N_2848,N_1746,N_1482);
nor U2849 (N_2849,N_1732,N_1812);
and U2850 (N_2850,N_1875,N_1906);
or U2851 (N_2851,N_1164,N_1132);
nand U2852 (N_2852,N_1874,N_1478);
or U2853 (N_2853,N_1895,N_1658);
and U2854 (N_2854,N_1053,N_1149);
and U2855 (N_2855,N_1284,N_1733);
and U2856 (N_2856,N_1488,N_1204);
nor U2857 (N_2857,N_1734,N_1532);
nand U2858 (N_2858,N_1986,N_1311);
nor U2859 (N_2859,N_1739,N_1168);
and U2860 (N_2860,N_1697,N_1213);
or U2861 (N_2861,N_1500,N_1218);
and U2862 (N_2862,N_1290,N_1253);
or U2863 (N_2863,N_1801,N_1379);
or U2864 (N_2864,N_1805,N_1332);
and U2865 (N_2865,N_1835,N_1090);
or U2866 (N_2866,N_1932,N_1716);
and U2867 (N_2867,N_1045,N_1023);
and U2868 (N_2868,N_1976,N_1908);
or U2869 (N_2869,N_1211,N_1675);
xor U2870 (N_2870,N_1383,N_1571);
nor U2871 (N_2871,N_1937,N_1118);
nand U2872 (N_2872,N_1877,N_1912);
and U2873 (N_2873,N_1000,N_1684);
and U2874 (N_2874,N_1352,N_1015);
and U2875 (N_2875,N_1520,N_1565);
nand U2876 (N_2876,N_1502,N_1771);
nand U2877 (N_2877,N_1464,N_1298);
nor U2878 (N_2878,N_1927,N_1168);
and U2879 (N_2879,N_1212,N_1233);
and U2880 (N_2880,N_1567,N_1348);
nand U2881 (N_2881,N_1325,N_1043);
and U2882 (N_2882,N_1800,N_1333);
nor U2883 (N_2883,N_1661,N_1257);
nor U2884 (N_2884,N_1886,N_1584);
and U2885 (N_2885,N_1688,N_1875);
or U2886 (N_2886,N_1013,N_1616);
and U2887 (N_2887,N_1799,N_1765);
nor U2888 (N_2888,N_1690,N_1777);
nand U2889 (N_2889,N_1028,N_1910);
and U2890 (N_2890,N_1030,N_1673);
nand U2891 (N_2891,N_1961,N_1873);
nand U2892 (N_2892,N_1998,N_1806);
xnor U2893 (N_2893,N_1658,N_1107);
xor U2894 (N_2894,N_1422,N_1669);
nor U2895 (N_2895,N_1870,N_1466);
nand U2896 (N_2896,N_1044,N_1577);
nor U2897 (N_2897,N_1617,N_1704);
nor U2898 (N_2898,N_1719,N_1278);
or U2899 (N_2899,N_1244,N_1716);
or U2900 (N_2900,N_1831,N_1576);
nor U2901 (N_2901,N_1787,N_1221);
nor U2902 (N_2902,N_1511,N_1276);
and U2903 (N_2903,N_1159,N_1182);
nand U2904 (N_2904,N_1407,N_1420);
or U2905 (N_2905,N_1830,N_1728);
and U2906 (N_2906,N_1200,N_1656);
nor U2907 (N_2907,N_1924,N_1034);
nor U2908 (N_2908,N_1547,N_1031);
nor U2909 (N_2909,N_1129,N_1876);
nor U2910 (N_2910,N_1398,N_1636);
nor U2911 (N_2911,N_1151,N_1263);
nor U2912 (N_2912,N_1495,N_1737);
and U2913 (N_2913,N_1596,N_1870);
nor U2914 (N_2914,N_1375,N_1854);
nor U2915 (N_2915,N_1334,N_1973);
nor U2916 (N_2916,N_1019,N_1081);
or U2917 (N_2917,N_1694,N_1165);
nor U2918 (N_2918,N_1349,N_1425);
nand U2919 (N_2919,N_1168,N_1120);
nand U2920 (N_2920,N_1580,N_1544);
or U2921 (N_2921,N_1797,N_1106);
nand U2922 (N_2922,N_1604,N_1282);
nand U2923 (N_2923,N_1013,N_1957);
xnor U2924 (N_2924,N_1945,N_1145);
nor U2925 (N_2925,N_1357,N_1775);
or U2926 (N_2926,N_1462,N_1443);
nand U2927 (N_2927,N_1319,N_1651);
and U2928 (N_2928,N_1322,N_1887);
and U2929 (N_2929,N_1239,N_1159);
or U2930 (N_2930,N_1427,N_1214);
nor U2931 (N_2931,N_1475,N_1066);
and U2932 (N_2932,N_1286,N_1388);
nor U2933 (N_2933,N_1898,N_1253);
nand U2934 (N_2934,N_1784,N_1807);
nand U2935 (N_2935,N_1187,N_1352);
nand U2936 (N_2936,N_1722,N_1389);
nand U2937 (N_2937,N_1826,N_1114);
and U2938 (N_2938,N_1838,N_1235);
or U2939 (N_2939,N_1704,N_1050);
and U2940 (N_2940,N_1190,N_1919);
or U2941 (N_2941,N_1018,N_1392);
and U2942 (N_2942,N_1349,N_1374);
nand U2943 (N_2943,N_1231,N_1340);
or U2944 (N_2944,N_1700,N_1934);
nand U2945 (N_2945,N_1537,N_1085);
nand U2946 (N_2946,N_1854,N_1645);
or U2947 (N_2947,N_1156,N_1307);
and U2948 (N_2948,N_1775,N_1145);
xor U2949 (N_2949,N_1853,N_1461);
and U2950 (N_2950,N_1754,N_1307);
or U2951 (N_2951,N_1384,N_1138);
nor U2952 (N_2952,N_1866,N_1925);
or U2953 (N_2953,N_1160,N_1689);
nand U2954 (N_2954,N_1358,N_1527);
nor U2955 (N_2955,N_1661,N_1532);
nand U2956 (N_2956,N_1997,N_1455);
nor U2957 (N_2957,N_1326,N_1864);
nor U2958 (N_2958,N_1405,N_1691);
and U2959 (N_2959,N_1085,N_1107);
and U2960 (N_2960,N_1237,N_1460);
or U2961 (N_2961,N_1682,N_1368);
nand U2962 (N_2962,N_1640,N_1973);
or U2963 (N_2963,N_1406,N_1280);
nand U2964 (N_2964,N_1728,N_1311);
nand U2965 (N_2965,N_1114,N_1205);
xor U2966 (N_2966,N_1956,N_1294);
nand U2967 (N_2967,N_1786,N_1142);
and U2968 (N_2968,N_1663,N_1625);
nand U2969 (N_2969,N_1050,N_1378);
and U2970 (N_2970,N_1401,N_1188);
nor U2971 (N_2971,N_1133,N_1763);
or U2972 (N_2972,N_1358,N_1940);
and U2973 (N_2973,N_1429,N_1118);
nor U2974 (N_2974,N_1269,N_1505);
nor U2975 (N_2975,N_1922,N_1021);
nand U2976 (N_2976,N_1623,N_1697);
or U2977 (N_2977,N_1106,N_1087);
or U2978 (N_2978,N_1654,N_1866);
and U2979 (N_2979,N_1403,N_1803);
nor U2980 (N_2980,N_1760,N_1173);
nand U2981 (N_2981,N_1272,N_1021);
nor U2982 (N_2982,N_1841,N_1312);
or U2983 (N_2983,N_1992,N_1932);
or U2984 (N_2984,N_1735,N_1945);
nand U2985 (N_2985,N_1441,N_1214);
and U2986 (N_2986,N_1685,N_1879);
nand U2987 (N_2987,N_1437,N_1232);
nand U2988 (N_2988,N_1851,N_1027);
nand U2989 (N_2989,N_1128,N_1182);
and U2990 (N_2990,N_1172,N_1715);
nand U2991 (N_2991,N_1785,N_1390);
nor U2992 (N_2992,N_1621,N_1952);
nor U2993 (N_2993,N_1187,N_1304);
nand U2994 (N_2994,N_1051,N_1072);
nand U2995 (N_2995,N_1862,N_1923);
nand U2996 (N_2996,N_1929,N_1046);
nor U2997 (N_2997,N_1872,N_1476);
or U2998 (N_2998,N_1311,N_1317);
and U2999 (N_2999,N_1687,N_1187);
and U3000 (N_3000,N_2684,N_2956);
and U3001 (N_3001,N_2365,N_2428);
nand U3002 (N_3002,N_2071,N_2023);
nand U3003 (N_3003,N_2567,N_2368);
nor U3004 (N_3004,N_2402,N_2622);
nand U3005 (N_3005,N_2735,N_2372);
nor U3006 (N_3006,N_2135,N_2155);
or U3007 (N_3007,N_2092,N_2668);
or U3008 (N_3008,N_2916,N_2286);
nor U3009 (N_3009,N_2929,N_2305);
nand U3010 (N_3010,N_2460,N_2193);
or U3011 (N_3011,N_2435,N_2664);
and U3012 (N_3012,N_2142,N_2274);
or U3013 (N_3013,N_2782,N_2583);
and U3014 (N_3014,N_2827,N_2679);
or U3015 (N_3015,N_2288,N_2014);
nand U3016 (N_3016,N_2983,N_2663);
nor U3017 (N_3017,N_2579,N_2808);
and U3018 (N_3018,N_2661,N_2870);
and U3019 (N_3019,N_2855,N_2660);
nand U3020 (N_3020,N_2657,N_2382);
nor U3021 (N_3021,N_2619,N_2159);
nand U3022 (N_3022,N_2090,N_2882);
nand U3023 (N_3023,N_2708,N_2821);
and U3024 (N_3024,N_2207,N_2917);
nor U3025 (N_3025,N_2051,N_2409);
nand U3026 (N_3026,N_2358,N_2872);
and U3027 (N_3027,N_2322,N_2411);
nor U3028 (N_3028,N_2762,N_2127);
or U3029 (N_3029,N_2361,N_2292);
and U3030 (N_3030,N_2601,N_2438);
nand U3031 (N_3031,N_2978,N_2050);
or U3032 (N_3032,N_2718,N_2323);
nand U3033 (N_3033,N_2891,N_2444);
and U3034 (N_3034,N_2055,N_2338);
and U3035 (N_3035,N_2743,N_2859);
nand U3036 (N_3036,N_2784,N_2229);
and U3037 (N_3037,N_2283,N_2775);
nand U3038 (N_3038,N_2058,N_2613);
nand U3039 (N_3039,N_2732,N_2678);
nor U3040 (N_3040,N_2451,N_2764);
xor U3041 (N_3041,N_2133,N_2144);
nor U3042 (N_3042,N_2550,N_2353);
xnor U3043 (N_3043,N_2319,N_2608);
or U3044 (N_3044,N_2041,N_2632);
nor U3045 (N_3045,N_2290,N_2406);
and U3046 (N_3046,N_2976,N_2988);
or U3047 (N_3047,N_2046,N_2880);
nand U3048 (N_3048,N_2896,N_2443);
and U3049 (N_3049,N_2836,N_2560);
nor U3050 (N_3050,N_2250,N_2065);
or U3051 (N_3051,N_2226,N_2310);
nand U3052 (N_3052,N_2778,N_2659);
or U3053 (N_3053,N_2815,N_2355);
and U3054 (N_3054,N_2677,N_2273);
nor U3055 (N_3055,N_2883,N_2333);
and U3056 (N_3056,N_2697,N_2706);
nor U3057 (N_3057,N_2696,N_2154);
nand U3058 (N_3058,N_2963,N_2504);
nand U3059 (N_3059,N_2424,N_2729);
nor U3060 (N_3060,N_2432,N_2776);
or U3061 (N_3061,N_2826,N_2833);
and U3062 (N_3062,N_2492,N_2884);
or U3063 (N_3063,N_2793,N_2466);
xor U3064 (N_3064,N_2630,N_2328);
and U3065 (N_3065,N_2379,N_2397);
nand U3066 (N_3066,N_2792,N_2446);
nand U3067 (N_3067,N_2434,N_2957);
nand U3068 (N_3068,N_2119,N_2543);
nor U3069 (N_3069,N_2810,N_2096);
and U3070 (N_3070,N_2057,N_2961);
nand U3071 (N_3071,N_2938,N_2255);
xor U3072 (N_3072,N_2923,N_2126);
or U3073 (N_3073,N_2238,N_2997);
nor U3074 (N_3074,N_2172,N_2831);
xnor U3075 (N_3075,N_2332,N_2813);
and U3076 (N_3076,N_2337,N_2575);
or U3077 (N_3077,N_2723,N_2299);
or U3078 (N_3078,N_2503,N_2053);
or U3079 (N_3079,N_2124,N_2311);
nor U3080 (N_3080,N_2116,N_2376);
nand U3081 (N_3081,N_2289,N_2812);
nand U3082 (N_3082,N_2941,N_2202);
or U3083 (N_3083,N_2750,N_2436);
nand U3084 (N_3084,N_2807,N_2072);
nand U3085 (N_3085,N_2141,N_2561);
nor U3086 (N_3086,N_2099,N_2847);
or U3087 (N_3087,N_2794,N_2535);
nor U3088 (N_3088,N_2441,N_2069);
or U3089 (N_3089,N_2029,N_2393);
nor U3090 (N_3090,N_2469,N_2738);
or U3091 (N_3091,N_2841,N_2817);
nand U3092 (N_3092,N_2722,N_2703);
nand U3093 (N_3093,N_2673,N_2828);
nor U3094 (N_3094,N_2086,N_2080);
or U3095 (N_3095,N_2910,N_2030);
or U3096 (N_3096,N_2167,N_2903);
nor U3097 (N_3097,N_2911,N_2758);
or U3098 (N_3098,N_2962,N_2400);
and U3099 (N_3099,N_2721,N_2196);
or U3100 (N_3100,N_2905,N_2129);
or U3101 (N_3101,N_2048,N_2313);
xnor U3102 (N_3102,N_2582,N_2125);
nand U3103 (N_3103,N_2330,N_2110);
and U3104 (N_3104,N_2858,N_2034);
or U3105 (N_3105,N_2741,N_2624);
and U3106 (N_3106,N_2060,N_2078);
nand U3107 (N_3107,N_2385,N_2166);
nor U3108 (N_3108,N_2066,N_2993);
and U3109 (N_3109,N_2416,N_2730);
and U3110 (N_3110,N_2000,N_2147);
and U3111 (N_3111,N_2566,N_2887);
nand U3112 (N_3112,N_2075,N_2820);
or U3113 (N_3113,N_2405,N_2208);
and U3114 (N_3114,N_2426,N_2982);
or U3115 (N_3115,N_2596,N_2533);
nand U3116 (N_3116,N_2984,N_2349);
and U3117 (N_3117,N_2079,N_2979);
or U3118 (N_3118,N_2518,N_2981);
or U3119 (N_3119,N_2942,N_2248);
or U3120 (N_3120,N_2879,N_2398);
nand U3121 (N_3121,N_2669,N_2958);
nor U3122 (N_3122,N_2001,N_2590);
and U3123 (N_3123,N_2136,N_2482);
or U3124 (N_3124,N_2570,N_2939);
nand U3125 (N_3125,N_2783,N_2946);
nand U3126 (N_3126,N_2893,N_2263);
or U3127 (N_3127,N_2035,N_2595);
nor U3128 (N_3128,N_2731,N_2915);
and U3129 (N_3129,N_2878,N_2187);
or U3130 (N_3130,N_2597,N_2199);
nand U3131 (N_3131,N_2763,N_2890);
nor U3132 (N_3132,N_2969,N_2170);
nand U3133 (N_3133,N_2948,N_2399);
or U3134 (N_3134,N_2727,N_2264);
xnor U3135 (N_3135,N_2391,N_2851);
and U3136 (N_3136,N_2656,N_2056);
and U3137 (N_3137,N_2759,N_2483);
or U3138 (N_3138,N_2370,N_2968);
and U3139 (N_3139,N_2375,N_2213);
or U3140 (N_3140,N_2487,N_2371);
and U3141 (N_3141,N_2239,N_2746);
or U3142 (N_3142,N_2865,N_2928);
or U3143 (N_3143,N_2157,N_2485);
or U3144 (N_3144,N_2307,N_2484);
and U3145 (N_3145,N_2612,N_2599);
and U3146 (N_3146,N_2991,N_2236);
nand U3147 (N_3147,N_2621,N_2117);
nand U3148 (N_3148,N_2242,N_2529);
nor U3149 (N_3149,N_2388,N_2037);
nand U3150 (N_3150,N_2574,N_2645);
or U3151 (N_3151,N_2798,N_2137);
nand U3152 (N_3152,N_2874,N_2546);
and U3153 (N_3153,N_2654,N_2083);
and U3154 (N_3154,N_2070,N_2260);
or U3155 (N_3155,N_2181,N_2182);
nor U3156 (N_3156,N_2510,N_2293);
or U3157 (N_3157,N_2052,N_2009);
nand U3158 (N_3158,N_2369,N_2519);
xnor U3159 (N_3159,N_2633,N_2251);
nor U3160 (N_3160,N_2838,N_2216);
nand U3161 (N_3161,N_2085,N_2790);
nor U3162 (N_3162,N_2284,N_2131);
nand U3163 (N_3163,N_2118,N_2024);
nor U3164 (N_3164,N_2215,N_2285);
and U3165 (N_3165,N_2606,N_2555);
nor U3166 (N_3166,N_2960,N_2860);
and U3167 (N_3167,N_2713,N_2985);
nor U3168 (N_3168,N_2572,N_2246);
nand U3169 (N_3169,N_2294,N_2287);
nand U3170 (N_3170,N_2699,N_2747);
and U3171 (N_3171,N_2588,N_2927);
or U3172 (N_3172,N_2521,N_2105);
nand U3173 (N_3173,N_2598,N_2839);
and U3174 (N_3174,N_2909,N_2809);
nand U3175 (N_3175,N_2276,N_2094);
and U3176 (N_3176,N_2930,N_2044);
nor U3177 (N_3177,N_2427,N_2611);
nor U3178 (N_3178,N_2600,N_2770);
and U3179 (N_3179,N_2327,N_2183);
and U3180 (N_3180,N_2501,N_2220);
nor U3181 (N_3181,N_2002,N_2087);
or U3182 (N_3182,N_2692,N_2174);
or U3183 (N_3183,N_2651,N_2152);
and U3184 (N_3184,N_2016,N_2043);
and U3185 (N_3185,N_2298,N_2728);
or U3186 (N_3186,N_2212,N_2556);
nor U3187 (N_3187,N_2457,N_2945);
or U3188 (N_3188,N_2218,N_2077);
nand U3189 (N_3189,N_2108,N_2547);
nor U3190 (N_3190,N_2716,N_2655);
and U3191 (N_3191,N_2495,N_2694);
nand U3192 (N_3192,N_2201,N_2774);
and U3193 (N_3193,N_2734,N_2303);
or U3194 (N_3194,N_2326,N_2455);
nand U3195 (N_3195,N_2297,N_2875);
and U3196 (N_3196,N_2950,N_2832);
xnor U3197 (N_3197,N_2671,N_2146);
nand U3198 (N_3198,N_2953,N_2502);
nor U3199 (N_3199,N_2081,N_2394);
or U3200 (N_3200,N_2802,N_2824);
nor U3201 (N_3201,N_2966,N_2279);
xnor U3202 (N_3202,N_2499,N_2450);
nand U3203 (N_3203,N_2410,N_2433);
or U3204 (N_3204,N_2805,N_2816);
or U3205 (N_3205,N_2688,N_2063);
or U3206 (N_3206,N_2190,N_2038);
nor U3207 (N_3207,N_2104,N_2800);
and U3208 (N_3208,N_2717,N_2359);
and U3209 (N_3209,N_2474,N_2390);
or U3210 (N_3210,N_2581,N_2940);
and U3211 (N_3211,N_2804,N_2591);
or U3212 (N_3212,N_2753,N_2021);
and U3213 (N_3213,N_2362,N_2791);
or U3214 (N_3214,N_2088,N_2974);
and U3215 (N_3215,N_2908,N_2015);
nand U3216 (N_3216,N_2225,N_2098);
nand U3217 (N_3217,N_2013,N_2578);
and U3218 (N_3218,N_2366,N_2524);
nor U3219 (N_3219,N_2569,N_2760);
nor U3220 (N_3220,N_2670,N_2799);
and U3221 (N_3221,N_2835,N_2165);
or U3222 (N_3222,N_2711,N_2430);
nor U3223 (N_3223,N_2489,N_2736);
or U3224 (N_3224,N_2840,N_2562);
and U3225 (N_3225,N_2228,N_2414);
nor U3226 (N_3226,N_2068,N_2959);
nand U3227 (N_3227,N_2237,N_2467);
nor U3228 (N_3228,N_2440,N_2522);
and U3229 (N_3229,N_2245,N_2089);
or U3230 (N_3230,N_2766,N_2350);
xor U3231 (N_3231,N_2607,N_2772);
nor U3232 (N_3232,N_2857,N_2179);
nand U3233 (N_3233,N_2342,N_2554);
or U3234 (N_3234,N_2465,N_2230);
nor U3235 (N_3235,N_2257,N_2500);
or U3236 (N_3236,N_2885,N_2160);
nand U3237 (N_3237,N_2262,N_2490);
xnor U3238 (N_3238,N_2845,N_2740);
or U3239 (N_3239,N_2296,N_2918);
or U3240 (N_3240,N_2819,N_2040);
and U3241 (N_3241,N_2949,N_2944);
or U3242 (N_3242,N_2223,N_2877);
and U3243 (N_3243,N_2867,N_2437);
nor U3244 (N_3244,N_2291,N_2061);
nor U3245 (N_3245,N_2360,N_2091);
or U3246 (N_3246,N_2986,N_2453);
nand U3247 (N_3247,N_2520,N_2275);
and U3248 (N_3248,N_2445,N_2317);
nor U3249 (N_3249,N_2200,N_2054);
nor U3250 (N_3250,N_2609,N_2989);
nand U3251 (N_3251,N_2203,N_2266);
nand U3252 (N_3252,N_2925,N_2616);
or U3253 (N_3253,N_2169,N_2922);
nor U3254 (N_3254,N_2536,N_2488);
and U3255 (N_3255,N_2900,N_2271);
or U3256 (N_3256,N_2111,N_2639);
nand U3257 (N_3257,N_2640,N_2647);
nor U3258 (N_3258,N_2897,N_2509);
or U3259 (N_3259,N_2109,N_2047);
nor U3260 (N_3260,N_2464,N_2823);
nand U3261 (N_3261,N_2803,N_2980);
and U3262 (N_3262,N_2121,N_2478);
nand U3263 (N_3263,N_2408,N_2497);
nor U3264 (N_3264,N_2892,N_2295);
and U3265 (N_3265,N_2100,N_2022);
nand U3266 (N_3266,N_2646,N_2304);
nor U3267 (N_3267,N_2834,N_2249);
and U3268 (N_3268,N_2666,N_2280);
or U3269 (N_3269,N_2964,N_2848);
and U3270 (N_3270,N_2593,N_2937);
or U3271 (N_3271,N_2904,N_2592);
or U3272 (N_3272,N_2649,N_2545);
or U3273 (N_3273,N_2321,N_2475);
nor U3274 (N_3274,N_2348,N_2525);
or U3275 (N_3275,N_2779,N_2143);
nor U3276 (N_3276,N_2972,N_2395);
nand U3277 (N_3277,N_2683,N_2818);
and U3278 (N_3278,N_2936,N_2352);
or U3279 (N_3279,N_2914,N_2797);
or U3280 (N_3280,N_2148,N_2565);
or U3281 (N_3281,N_2415,N_2019);
and U3282 (N_3282,N_2843,N_2615);
nand U3283 (N_3283,N_2439,N_2259);
and U3284 (N_3284,N_2744,N_2132);
nand U3285 (N_3285,N_2977,N_2045);
and U3286 (N_3286,N_2346,N_2773);
nand U3287 (N_3287,N_2335,N_2527);
and U3288 (N_3288,N_2955,N_2448);
nor U3289 (N_3289,N_2505,N_2244);
nor U3290 (N_3290,N_2171,N_2139);
or U3291 (N_3291,N_2685,N_2681);
and U3292 (N_3292,N_2343,N_2067);
nand U3293 (N_3293,N_2301,N_2856);
nor U3294 (N_3294,N_2373,N_2752);
and U3295 (N_3295,N_2853,N_2272);
nand U3296 (N_3296,N_2906,N_2462);
or U3297 (N_3297,N_2617,N_2888);
or U3298 (N_3298,N_2185,N_2998);
and U3299 (N_3299,N_2481,N_2999);
or U3300 (N_3300,N_2227,N_2454);
and U3301 (N_3301,N_2219,N_2552);
xor U3302 (N_3302,N_2195,N_2217);
nand U3303 (N_3303,N_2221,N_2894);
nor U3304 (N_3304,N_2757,N_2042);
or U3305 (N_3305,N_2324,N_2967);
nand U3306 (N_3306,N_2261,N_2281);
nand U3307 (N_3307,N_2913,N_2755);
nand U3308 (N_3308,N_2702,N_2205);
xnor U3309 (N_3309,N_2383,N_2719);
nor U3310 (N_3310,N_2107,N_2267);
nor U3311 (N_3311,N_2122,N_2175);
and U3312 (N_3312,N_2233,N_2517);
or U3313 (N_3313,N_2496,N_2479);
and U3314 (N_3314,N_2407,N_2541);
nor U3315 (N_3315,N_2341,N_2252);
nor U3316 (N_3316,N_2354,N_2866);
or U3317 (N_3317,N_2173,N_2682);
and U3318 (N_3318,N_2951,N_2846);
nand U3319 (N_3319,N_2318,N_2025);
nand U3320 (N_3320,N_2302,N_2602);
nor U3321 (N_3321,N_2667,N_2452);
or U3322 (N_3322,N_2074,N_2036);
and U3323 (N_3323,N_2198,N_2745);
or U3324 (N_3324,N_2557,N_2367);
nand U3325 (N_3325,N_2629,N_2258);
nand U3326 (N_3326,N_2020,N_2336);
nand U3327 (N_3327,N_2114,N_2636);
or U3328 (N_3328,N_2282,N_2975);
and U3329 (N_3329,N_2234,N_2192);
nor U3330 (N_3330,N_2447,N_2027);
and U3331 (N_3331,N_2902,N_2003);
nor U3332 (N_3332,N_2516,N_2850);
and U3333 (N_3333,N_2480,N_2811);
and U3334 (N_3334,N_2005,N_2351);
and U3335 (N_3335,N_2970,N_2584);
nor U3336 (N_3336,N_2780,N_2726);
and U3337 (N_3337,N_2634,N_2638);
nor U3338 (N_3338,N_2564,N_2101);
and U3339 (N_3339,N_2339,N_2162);
xnor U3340 (N_3340,N_2429,N_2994);
nor U3341 (N_3341,N_2103,N_2700);
or U3342 (N_3342,N_2308,N_2754);
nand U3343 (N_3343,N_2268,N_2854);
and U3344 (N_3344,N_2680,N_2720);
nand U3345 (N_3345,N_2990,N_2537);
nand U3346 (N_3346,N_2786,N_2625);
nand U3347 (N_3347,N_2392,N_2620);
nor U3348 (N_3348,N_2577,N_2788);
nor U3349 (N_3349,N_2231,N_2912);
nor U3350 (N_3350,N_2269,N_2331);
and U3351 (N_3351,N_2222,N_2418);
nor U3352 (N_3352,N_2423,N_2039);
and U3353 (N_3353,N_2387,N_2907);
nand U3354 (N_3354,N_2586,N_2540);
xor U3355 (N_3355,N_2931,N_2476);
or U3356 (N_3356,N_2364,N_2689);
nand U3357 (N_3357,N_2120,N_2184);
nor U3358 (N_3358,N_2232,N_2442);
nor U3359 (N_3359,N_2357,N_2344);
nand U3360 (N_3360,N_2761,N_2589);
nand U3361 (N_3361,N_2210,N_2587);
nand U3362 (N_3362,N_2176,N_2926);
and U3363 (N_3363,N_2064,N_2412);
or U3364 (N_3364,N_2345,N_2549);
nand U3365 (N_3365,N_2559,N_2377);
nand U3366 (N_3366,N_2168,N_2924);
or U3367 (N_3367,N_2224,N_2254);
nand U3368 (N_3368,N_2277,N_2511);
or U3369 (N_3369,N_2386,N_2463);
nor U3370 (N_3370,N_2539,N_2449);
nand U3371 (N_3371,N_2158,N_2420);
nand U3372 (N_3372,N_2695,N_2115);
nor U3373 (N_3373,N_2523,N_2724);
or U3374 (N_3374,N_2073,N_2186);
nor U3375 (N_3375,N_2189,N_2710);
or U3376 (N_3376,N_2919,N_2513);
nand U3377 (N_3377,N_2471,N_2725);
nor U3378 (N_3378,N_2008,N_2707);
nor U3379 (N_3379,N_2934,N_2102);
nand U3380 (N_3380,N_2140,N_2691);
or U3381 (N_3381,N_2243,N_2932);
or U3382 (N_3382,N_2571,N_2806);
nand U3383 (N_3383,N_2526,N_2401);
nor U3384 (N_3384,N_2861,N_2751);
nand U3385 (N_3385,N_2614,N_2658);
xnor U3386 (N_3386,N_2568,N_2765);
or U3387 (N_3387,N_2194,N_2781);
nand U3388 (N_3388,N_2486,N_2204);
or U3389 (N_3389,N_2756,N_2873);
and U3390 (N_3390,N_2749,N_2796);
or U3391 (N_3391,N_2704,N_2844);
or U3392 (N_3392,N_2610,N_2422);
and U3393 (N_3393,N_2188,N_2895);
nor U3394 (N_3394,N_2363,N_2635);
nand U3395 (N_3395,N_2130,N_2177);
nand U3396 (N_3396,N_2106,N_2863);
and U3397 (N_3397,N_2652,N_2748);
nor U3398 (N_3398,N_2012,N_2507);
nor U3399 (N_3399,N_2028,N_2628);
nand U3400 (N_3400,N_2240,N_2709);
nand U3401 (N_3401,N_2082,N_2627);
or U3402 (N_3402,N_2653,N_2306);
nor U3403 (N_3403,N_2605,N_2933);
nor U3404 (N_3404,N_2211,N_2769);
or U3405 (N_3405,N_2494,N_2134);
and U3406 (N_3406,N_2742,N_2417);
nor U3407 (N_3407,N_2714,N_2553);
nor U3408 (N_3408,N_2603,N_2626);
nor U3409 (N_3409,N_2899,N_2876);
or U3410 (N_3410,N_2693,N_2995);
or U3411 (N_3411,N_2270,N_2643);
and U3412 (N_3412,N_2825,N_2644);
and U3413 (N_3413,N_2347,N_2973);
nor U3414 (N_3414,N_2325,N_2642);
or U3415 (N_3415,N_2686,N_2690);
and U3416 (N_3416,N_2795,N_2675);
or U3417 (N_3417,N_2178,N_2952);
or U3418 (N_3418,N_2687,N_2315);
or U3419 (N_3419,N_2701,N_2007);
and U3420 (N_3420,N_2886,N_2316);
nand U3421 (N_3421,N_2739,N_2381);
nor U3422 (N_3422,N_2868,N_2580);
or U3423 (N_3423,N_2265,N_2456);
nand U3424 (N_3424,N_2864,N_2425);
or U3425 (N_3425,N_2163,N_2623);
nor U3426 (N_3426,N_2789,N_2340);
or U3427 (N_3427,N_2197,N_2421);
nor U3428 (N_3428,N_2996,N_2881);
nand U3429 (N_3429,N_2641,N_2594);
or U3430 (N_3430,N_2389,N_2151);
and U3431 (N_3431,N_2538,N_2247);
nor U3432 (N_3432,N_2241,N_2512);
nand U3433 (N_3433,N_2631,N_2128);
or U3434 (N_3434,N_2309,N_2206);
or U3435 (N_3435,N_2563,N_2384);
or U3436 (N_3436,N_2472,N_2737);
xor U3437 (N_3437,N_2650,N_2777);
and U3438 (N_3438,N_2093,N_2076);
nand U3439 (N_3439,N_2935,N_2180);
nand U3440 (N_3440,N_2698,N_2059);
nand U3441 (N_3441,N_2062,N_2123);
and U3442 (N_3442,N_2508,N_2149);
and U3443 (N_3443,N_2901,N_2558);
xnor U3444 (N_3444,N_2862,N_2032);
and U3445 (N_3445,N_2604,N_2733);
or U3446 (N_3446,N_2712,N_2477);
nor U3447 (N_3447,N_2871,N_2459);
and U3448 (N_3448,N_2461,N_2506);
and U3449 (N_3449,N_2842,N_2637);
nand U3450 (N_3450,N_2150,N_2889);
and U3451 (N_3451,N_2648,N_2113);
or U3452 (N_3452,N_2514,N_2822);
nand U3453 (N_3453,N_2404,N_2837);
and U3454 (N_3454,N_2097,N_2965);
nand U3455 (N_3455,N_2209,N_2235);
and U3456 (N_3456,N_2665,N_2705);
or U3457 (N_3457,N_2491,N_2314);
or U3458 (N_3458,N_2530,N_2715);
or U3459 (N_3459,N_2145,N_2576);
and U3460 (N_3460,N_2403,N_2138);
nor U3461 (N_3461,N_2084,N_2771);
or U3462 (N_3462,N_2768,N_2413);
nor U3463 (N_3463,N_2214,N_2662);
or U3464 (N_3464,N_2814,N_2787);
or U3465 (N_3465,N_2112,N_2618);
or U3466 (N_3466,N_2548,N_2920);
or U3467 (N_3467,N_2468,N_2829);
xnor U3468 (N_3468,N_2921,N_2396);
and U3469 (N_3469,N_2031,N_2528);
and U3470 (N_3470,N_2544,N_2943);
nor U3471 (N_3471,N_2672,N_2191);
or U3472 (N_3472,N_2992,N_2542);
and U3473 (N_3473,N_2849,N_2164);
or U3474 (N_3474,N_2515,N_2676);
nand U3475 (N_3475,N_2334,N_2531);
nand U3476 (N_3476,N_2498,N_2532);
or U3477 (N_3477,N_2987,N_2473);
and U3478 (N_3478,N_2898,N_2018);
and U3479 (N_3479,N_2006,N_2049);
and U3480 (N_3480,N_2374,N_2329);
nand U3481 (N_3481,N_2801,N_2278);
or U3482 (N_3482,N_2431,N_2026);
or U3483 (N_3483,N_2551,N_2017);
nand U3484 (N_3484,N_2033,N_2095);
or U3485 (N_3485,N_2852,N_2971);
nand U3486 (N_3486,N_2674,N_2378);
or U3487 (N_3487,N_2320,N_2954);
or U3488 (N_3488,N_2253,N_2011);
and U3489 (N_3489,N_2470,N_2419);
nor U3490 (N_3490,N_2010,N_2534);
and U3491 (N_3491,N_2947,N_2767);
and U3492 (N_3492,N_2869,N_2458);
or U3493 (N_3493,N_2573,N_2585);
and U3494 (N_3494,N_2161,N_2830);
or U3495 (N_3495,N_2356,N_2256);
and U3496 (N_3496,N_2156,N_2312);
nor U3497 (N_3497,N_2004,N_2493);
nand U3498 (N_3498,N_2380,N_2300);
and U3499 (N_3499,N_2153,N_2785);
or U3500 (N_3500,N_2311,N_2211);
and U3501 (N_3501,N_2403,N_2035);
nand U3502 (N_3502,N_2422,N_2228);
or U3503 (N_3503,N_2442,N_2810);
nand U3504 (N_3504,N_2329,N_2633);
and U3505 (N_3505,N_2847,N_2158);
nor U3506 (N_3506,N_2043,N_2881);
nor U3507 (N_3507,N_2266,N_2401);
nand U3508 (N_3508,N_2598,N_2844);
and U3509 (N_3509,N_2551,N_2207);
or U3510 (N_3510,N_2745,N_2186);
nor U3511 (N_3511,N_2316,N_2375);
nor U3512 (N_3512,N_2550,N_2501);
and U3513 (N_3513,N_2162,N_2381);
and U3514 (N_3514,N_2447,N_2077);
nor U3515 (N_3515,N_2521,N_2396);
nor U3516 (N_3516,N_2182,N_2034);
or U3517 (N_3517,N_2908,N_2959);
nor U3518 (N_3518,N_2587,N_2714);
nor U3519 (N_3519,N_2894,N_2089);
nand U3520 (N_3520,N_2643,N_2075);
and U3521 (N_3521,N_2395,N_2351);
nor U3522 (N_3522,N_2293,N_2468);
nand U3523 (N_3523,N_2173,N_2984);
and U3524 (N_3524,N_2503,N_2626);
and U3525 (N_3525,N_2265,N_2425);
or U3526 (N_3526,N_2147,N_2148);
nand U3527 (N_3527,N_2854,N_2185);
or U3528 (N_3528,N_2359,N_2272);
and U3529 (N_3529,N_2326,N_2238);
nor U3530 (N_3530,N_2851,N_2884);
nand U3531 (N_3531,N_2546,N_2864);
nor U3532 (N_3532,N_2481,N_2920);
nand U3533 (N_3533,N_2796,N_2530);
nand U3534 (N_3534,N_2426,N_2648);
or U3535 (N_3535,N_2738,N_2951);
nor U3536 (N_3536,N_2359,N_2905);
nand U3537 (N_3537,N_2675,N_2026);
or U3538 (N_3538,N_2863,N_2841);
and U3539 (N_3539,N_2510,N_2344);
and U3540 (N_3540,N_2069,N_2821);
and U3541 (N_3541,N_2099,N_2957);
nor U3542 (N_3542,N_2289,N_2232);
and U3543 (N_3543,N_2617,N_2000);
or U3544 (N_3544,N_2505,N_2606);
or U3545 (N_3545,N_2194,N_2976);
and U3546 (N_3546,N_2957,N_2414);
xor U3547 (N_3547,N_2147,N_2245);
and U3548 (N_3548,N_2173,N_2224);
nor U3549 (N_3549,N_2504,N_2776);
and U3550 (N_3550,N_2330,N_2988);
and U3551 (N_3551,N_2442,N_2003);
nor U3552 (N_3552,N_2192,N_2751);
or U3553 (N_3553,N_2618,N_2030);
nand U3554 (N_3554,N_2379,N_2889);
nor U3555 (N_3555,N_2092,N_2170);
nor U3556 (N_3556,N_2101,N_2717);
nand U3557 (N_3557,N_2487,N_2879);
or U3558 (N_3558,N_2463,N_2424);
and U3559 (N_3559,N_2067,N_2286);
nor U3560 (N_3560,N_2382,N_2920);
or U3561 (N_3561,N_2270,N_2818);
nor U3562 (N_3562,N_2111,N_2949);
or U3563 (N_3563,N_2616,N_2670);
and U3564 (N_3564,N_2390,N_2931);
or U3565 (N_3565,N_2297,N_2335);
and U3566 (N_3566,N_2217,N_2477);
or U3567 (N_3567,N_2429,N_2637);
nor U3568 (N_3568,N_2201,N_2384);
or U3569 (N_3569,N_2707,N_2274);
nand U3570 (N_3570,N_2951,N_2831);
and U3571 (N_3571,N_2020,N_2532);
nand U3572 (N_3572,N_2776,N_2019);
or U3573 (N_3573,N_2522,N_2363);
and U3574 (N_3574,N_2310,N_2718);
and U3575 (N_3575,N_2760,N_2554);
nor U3576 (N_3576,N_2854,N_2480);
nand U3577 (N_3577,N_2693,N_2958);
and U3578 (N_3578,N_2015,N_2044);
nand U3579 (N_3579,N_2994,N_2559);
and U3580 (N_3580,N_2057,N_2591);
nand U3581 (N_3581,N_2564,N_2044);
nand U3582 (N_3582,N_2422,N_2517);
or U3583 (N_3583,N_2275,N_2622);
or U3584 (N_3584,N_2196,N_2212);
nand U3585 (N_3585,N_2179,N_2243);
nand U3586 (N_3586,N_2077,N_2471);
nor U3587 (N_3587,N_2015,N_2748);
and U3588 (N_3588,N_2435,N_2179);
nand U3589 (N_3589,N_2042,N_2592);
or U3590 (N_3590,N_2015,N_2510);
or U3591 (N_3591,N_2637,N_2873);
nand U3592 (N_3592,N_2205,N_2512);
nand U3593 (N_3593,N_2299,N_2173);
or U3594 (N_3594,N_2509,N_2077);
and U3595 (N_3595,N_2049,N_2712);
nand U3596 (N_3596,N_2314,N_2636);
and U3597 (N_3597,N_2461,N_2469);
nand U3598 (N_3598,N_2342,N_2453);
nand U3599 (N_3599,N_2251,N_2223);
nand U3600 (N_3600,N_2168,N_2899);
or U3601 (N_3601,N_2897,N_2475);
or U3602 (N_3602,N_2452,N_2378);
and U3603 (N_3603,N_2747,N_2547);
nand U3604 (N_3604,N_2851,N_2772);
and U3605 (N_3605,N_2207,N_2977);
or U3606 (N_3606,N_2920,N_2164);
and U3607 (N_3607,N_2643,N_2194);
nor U3608 (N_3608,N_2466,N_2278);
or U3609 (N_3609,N_2080,N_2491);
nor U3610 (N_3610,N_2274,N_2696);
and U3611 (N_3611,N_2757,N_2423);
and U3612 (N_3612,N_2222,N_2033);
nand U3613 (N_3613,N_2978,N_2663);
nand U3614 (N_3614,N_2853,N_2543);
nand U3615 (N_3615,N_2426,N_2659);
nor U3616 (N_3616,N_2971,N_2309);
nand U3617 (N_3617,N_2080,N_2746);
nor U3618 (N_3618,N_2781,N_2672);
or U3619 (N_3619,N_2081,N_2902);
nor U3620 (N_3620,N_2034,N_2468);
or U3621 (N_3621,N_2687,N_2667);
nand U3622 (N_3622,N_2106,N_2528);
nand U3623 (N_3623,N_2022,N_2827);
or U3624 (N_3624,N_2134,N_2069);
nor U3625 (N_3625,N_2119,N_2070);
nor U3626 (N_3626,N_2042,N_2579);
nand U3627 (N_3627,N_2997,N_2893);
and U3628 (N_3628,N_2124,N_2904);
or U3629 (N_3629,N_2533,N_2167);
or U3630 (N_3630,N_2816,N_2429);
nand U3631 (N_3631,N_2705,N_2362);
or U3632 (N_3632,N_2925,N_2019);
nor U3633 (N_3633,N_2043,N_2738);
and U3634 (N_3634,N_2838,N_2303);
and U3635 (N_3635,N_2694,N_2389);
and U3636 (N_3636,N_2430,N_2134);
and U3637 (N_3637,N_2518,N_2389);
nor U3638 (N_3638,N_2521,N_2366);
or U3639 (N_3639,N_2841,N_2143);
nor U3640 (N_3640,N_2966,N_2602);
nor U3641 (N_3641,N_2859,N_2158);
nand U3642 (N_3642,N_2245,N_2686);
or U3643 (N_3643,N_2359,N_2398);
or U3644 (N_3644,N_2080,N_2831);
and U3645 (N_3645,N_2269,N_2349);
nand U3646 (N_3646,N_2450,N_2228);
xor U3647 (N_3647,N_2241,N_2915);
nand U3648 (N_3648,N_2658,N_2749);
or U3649 (N_3649,N_2443,N_2495);
or U3650 (N_3650,N_2678,N_2887);
nand U3651 (N_3651,N_2018,N_2551);
or U3652 (N_3652,N_2811,N_2616);
nand U3653 (N_3653,N_2370,N_2759);
nor U3654 (N_3654,N_2294,N_2766);
nor U3655 (N_3655,N_2587,N_2149);
and U3656 (N_3656,N_2005,N_2203);
and U3657 (N_3657,N_2275,N_2526);
and U3658 (N_3658,N_2242,N_2092);
or U3659 (N_3659,N_2145,N_2151);
nand U3660 (N_3660,N_2107,N_2490);
and U3661 (N_3661,N_2938,N_2598);
or U3662 (N_3662,N_2613,N_2896);
nor U3663 (N_3663,N_2639,N_2303);
xor U3664 (N_3664,N_2303,N_2093);
xor U3665 (N_3665,N_2339,N_2239);
nand U3666 (N_3666,N_2888,N_2513);
or U3667 (N_3667,N_2351,N_2250);
nor U3668 (N_3668,N_2261,N_2576);
nand U3669 (N_3669,N_2820,N_2475);
and U3670 (N_3670,N_2399,N_2075);
and U3671 (N_3671,N_2133,N_2235);
or U3672 (N_3672,N_2885,N_2642);
nand U3673 (N_3673,N_2889,N_2977);
and U3674 (N_3674,N_2336,N_2225);
nor U3675 (N_3675,N_2756,N_2646);
nor U3676 (N_3676,N_2704,N_2248);
or U3677 (N_3677,N_2758,N_2815);
nor U3678 (N_3678,N_2350,N_2661);
nor U3679 (N_3679,N_2741,N_2921);
nand U3680 (N_3680,N_2273,N_2476);
xnor U3681 (N_3681,N_2866,N_2651);
nand U3682 (N_3682,N_2918,N_2357);
and U3683 (N_3683,N_2932,N_2663);
and U3684 (N_3684,N_2455,N_2739);
nor U3685 (N_3685,N_2549,N_2386);
or U3686 (N_3686,N_2499,N_2072);
nand U3687 (N_3687,N_2044,N_2216);
nor U3688 (N_3688,N_2643,N_2906);
nand U3689 (N_3689,N_2322,N_2474);
nand U3690 (N_3690,N_2346,N_2897);
nor U3691 (N_3691,N_2895,N_2027);
nor U3692 (N_3692,N_2050,N_2560);
nand U3693 (N_3693,N_2935,N_2923);
or U3694 (N_3694,N_2664,N_2136);
nor U3695 (N_3695,N_2418,N_2904);
or U3696 (N_3696,N_2278,N_2249);
nand U3697 (N_3697,N_2310,N_2744);
nand U3698 (N_3698,N_2673,N_2207);
nand U3699 (N_3699,N_2707,N_2250);
or U3700 (N_3700,N_2928,N_2705);
or U3701 (N_3701,N_2678,N_2348);
nand U3702 (N_3702,N_2061,N_2718);
or U3703 (N_3703,N_2441,N_2305);
nor U3704 (N_3704,N_2636,N_2401);
nand U3705 (N_3705,N_2472,N_2682);
nand U3706 (N_3706,N_2458,N_2313);
nor U3707 (N_3707,N_2748,N_2850);
and U3708 (N_3708,N_2445,N_2993);
nand U3709 (N_3709,N_2347,N_2720);
or U3710 (N_3710,N_2892,N_2792);
and U3711 (N_3711,N_2716,N_2670);
nor U3712 (N_3712,N_2738,N_2662);
and U3713 (N_3713,N_2214,N_2443);
or U3714 (N_3714,N_2382,N_2955);
nand U3715 (N_3715,N_2379,N_2708);
nand U3716 (N_3716,N_2740,N_2441);
nor U3717 (N_3717,N_2850,N_2913);
nand U3718 (N_3718,N_2464,N_2184);
xnor U3719 (N_3719,N_2936,N_2276);
or U3720 (N_3720,N_2837,N_2672);
and U3721 (N_3721,N_2253,N_2427);
nand U3722 (N_3722,N_2880,N_2611);
nand U3723 (N_3723,N_2214,N_2653);
and U3724 (N_3724,N_2328,N_2561);
and U3725 (N_3725,N_2640,N_2957);
nand U3726 (N_3726,N_2790,N_2781);
nand U3727 (N_3727,N_2186,N_2764);
nor U3728 (N_3728,N_2317,N_2930);
and U3729 (N_3729,N_2811,N_2256);
and U3730 (N_3730,N_2918,N_2217);
nor U3731 (N_3731,N_2256,N_2521);
or U3732 (N_3732,N_2213,N_2583);
nand U3733 (N_3733,N_2782,N_2999);
or U3734 (N_3734,N_2172,N_2051);
or U3735 (N_3735,N_2682,N_2296);
or U3736 (N_3736,N_2847,N_2368);
and U3737 (N_3737,N_2443,N_2647);
and U3738 (N_3738,N_2541,N_2654);
nand U3739 (N_3739,N_2883,N_2595);
or U3740 (N_3740,N_2141,N_2562);
nor U3741 (N_3741,N_2745,N_2971);
nand U3742 (N_3742,N_2075,N_2806);
or U3743 (N_3743,N_2717,N_2299);
nor U3744 (N_3744,N_2125,N_2084);
or U3745 (N_3745,N_2588,N_2933);
or U3746 (N_3746,N_2456,N_2161);
nand U3747 (N_3747,N_2026,N_2062);
or U3748 (N_3748,N_2354,N_2878);
nor U3749 (N_3749,N_2201,N_2318);
nand U3750 (N_3750,N_2826,N_2798);
and U3751 (N_3751,N_2124,N_2680);
or U3752 (N_3752,N_2620,N_2917);
or U3753 (N_3753,N_2334,N_2660);
nor U3754 (N_3754,N_2806,N_2463);
nand U3755 (N_3755,N_2111,N_2945);
or U3756 (N_3756,N_2639,N_2004);
nand U3757 (N_3757,N_2825,N_2509);
nand U3758 (N_3758,N_2920,N_2642);
and U3759 (N_3759,N_2765,N_2770);
nand U3760 (N_3760,N_2897,N_2842);
nand U3761 (N_3761,N_2897,N_2496);
or U3762 (N_3762,N_2248,N_2116);
and U3763 (N_3763,N_2378,N_2984);
nor U3764 (N_3764,N_2490,N_2693);
xor U3765 (N_3765,N_2044,N_2297);
nor U3766 (N_3766,N_2914,N_2624);
nand U3767 (N_3767,N_2979,N_2133);
nand U3768 (N_3768,N_2574,N_2342);
or U3769 (N_3769,N_2842,N_2923);
nor U3770 (N_3770,N_2238,N_2303);
or U3771 (N_3771,N_2109,N_2782);
and U3772 (N_3772,N_2205,N_2745);
and U3773 (N_3773,N_2777,N_2898);
nand U3774 (N_3774,N_2391,N_2151);
and U3775 (N_3775,N_2723,N_2041);
and U3776 (N_3776,N_2569,N_2044);
and U3777 (N_3777,N_2048,N_2885);
or U3778 (N_3778,N_2755,N_2443);
nor U3779 (N_3779,N_2970,N_2409);
and U3780 (N_3780,N_2622,N_2242);
nand U3781 (N_3781,N_2302,N_2737);
nand U3782 (N_3782,N_2331,N_2284);
nand U3783 (N_3783,N_2216,N_2152);
or U3784 (N_3784,N_2893,N_2722);
nor U3785 (N_3785,N_2122,N_2121);
or U3786 (N_3786,N_2320,N_2630);
and U3787 (N_3787,N_2823,N_2620);
or U3788 (N_3788,N_2640,N_2696);
nand U3789 (N_3789,N_2990,N_2702);
and U3790 (N_3790,N_2488,N_2746);
and U3791 (N_3791,N_2311,N_2158);
xor U3792 (N_3792,N_2304,N_2766);
and U3793 (N_3793,N_2718,N_2438);
or U3794 (N_3794,N_2547,N_2083);
and U3795 (N_3795,N_2029,N_2480);
nand U3796 (N_3796,N_2731,N_2019);
and U3797 (N_3797,N_2109,N_2600);
and U3798 (N_3798,N_2192,N_2345);
nand U3799 (N_3799,N_2157,N_2862);
or U3800 (N_3800,N_2181,N_2934);
and U3801 (N_3801,N_2560,N_2381);
or U3802 (N_3802,N_2886,N_2139);
nor U3803 (N_3803,N_2779,N_2595);
nor U3804 (N_3804,N_2162,N_2206);
nor U3805 (N_3805,N_2309,N_2579);
nand U3806 (N_3806,N_2827,N_2184);
and U3807 (N_3807,N_2425,N_2089);
xor U3808 (N_3808,N_2560,N_2569);
and U3809 (N_3809,N_2746,N_2235);
or U3810 (N_3810,N_2815,N_2503);
and U3811 (N_3811,N_2599,N_2506);
and U3812 (N_3812,N_2650,N_2060);
nand U3813 (N_3813,N_2900,N_2798);
nand U3814 (N_3814,N_2648,N_2202);
nand U3815 (N_3815,N_2010,N_2198);
nand U3816 (N_3816,N_2139,N_2375);
and U3817 (N_3817,N_2786,N_2449);
or U3818 (N_3818,N_2553,N_2333);
or U3819 (N_3819,N_2267,N_2241);
or U3820 (N_3820,N_2600,N_2097);
or U3821 (N_3821,N_2173,N_2270);
nand U3822 (N_3822,N_2034,N_2603);
nand U3823 (N_3823,N_2628,N_2888);
nor U3824 (N_3824,N_2117,N_2649);
or U3825 (N_3825,N_2290,N_2356);
and U3826 (N_3826,N_2455,N_2420);
or U3827 (N_3827,N_2438,N_2040);
or U3828 (N_3828,N_2752,N_2084);
or U3829 (N_3829,N_2942,N_2039);
nor U3830 (N_3830,N_2821,N_2744);
or U3831 (N_3831,N_2531,N_2935);
and U3832 (N_3832,N_2040,N_2593);
nor U3833 (N_3833,N_2935,N_2670);
nor U3834 (N_3834,N_2709,N_2834);
nand U3835 (N_3835,N_2798,N_2002);
nor U3836 (N_3836,N_2121,N_2020);
and U3837 (N_3837,N_2299,N_2414);
nand U3838 (N_3838,N_2161,N_2851);
and U3839 (N_3839,N_2490,N_2301);
xor U3840 (N_3840,N_2861,N_2590);
and U3841 (N_3841,N_2594,N_2926);
and U3842 (N_3842,N_2184,N_2351);
or U3843 (N_3843,N_2202,N_2112);
nor U3844 (N_3844,N_2723,N_2466);
or U3845 (N_3845,N_2325,N_2251);
or U3846 (N_3846,N_2687,N_2679);
nand U3847 (N_3847,N_2987,N_2649);
nor U3848 (N_3848,N_2431,N_2971);
nor U3849 (N_3849,N_2527,N_2245);
and U3850 (N_3850,N_2747,N_2099);
and U3851 (N_3851,N_2357,N_2371);
or U3852 (N_3852,N_2399,N_2204);
or U3853 (N_3853,N_2540,N_2308);
and U3854 (N_3854,N_2207,N_2961);
and U3855 (N_3855,N_2540,N_2176);
nor U3856 (N_3856,N_2191,N_2639);
nand U3857 (N_3857,N_2681,N_2095);
and U3858 (N_3858,N_2735,N_2470);
nand U3859 (N_3859,N_2866,N_2085);
nor U3860 (N_3860,N_2662,N_2084);
or U3861 (N_3861,N_2132,N_2413);
or U3862 (N_3862,N_2608,N_2874);
or U3863 (N_3863,N_2622,N_2156);
and U3864 (N_3864,N_2900,N_2876);
xnor U3865 (N_3865,N_2191,N_2134);
nor U3866 (N_3866,N_2688,N_2288);
nor U3867 (N_3867,N_2025,N_2661);
nor U3868 (N_3868,N_2238,N_2036);
nor U3869 (N_3869,N_2574,N_2945);
xnor U3870 (N_3870,N_2927,N_2164);
or U3871 (N_3871,N_2809,N_2094);
and U3872 (N_3872,N_2410,N_2251);
nand U3873 (N_3873,N_2248,N_2709);
nor U3874 (N_3874,N_2042,N_2072);
nand U3875 (N_3875,N_2466,N_2626);
or U3876 (N_3876,N_2879,N_2090);
or U3877 (N_3877,N_2145,N_2603);
or U3878 (N_3878,N_2411,N_2038);
nor U3879 (N_3879,N_2934,N_2776);
and U3880 (N_3880,N_2091,N_2361);
and U3881 (N_3881,N_2133,N_2039);
nand U3882 (N_3882,N_2123,N_2423);
and U3883 (N_3883,N_2629,N_2750);
or U3884 (N_3884,N_2900,N_2459);
nor U3885 (N_3885,N_2211,N_2275);
nand U3886 (N_3886,N_2935,N_2247);
or U3887 (N_3887,N_2006,N_2694);
nor U3888 (N_3888,N_2164,N_2377);
nor U3889 (N_3889,N_2801,N_2299);
or U3890 (N_3890,N_2433,N_2213);
xnor U3891 (N_3891,N_2487,N_2771);
or U3892 (N_3892,N_2094,N_2406);
and U3893 (N_3893,N_2514,N_2460);
and U3894 (N_3894,N_2098,N_2003);
nand U3895 (N_3895,N_2973,N_2354);
and U3896 (N_3896,N_2790,N_2732);
nor U3897 (N_3897,N_2188,N_2759);
or U3898 (N_3898,N_2791,N_2025);
nor U3899 (N_3899,N_2593,N_2925);
and U3900 (N_3900,N_2385,N_2939);
nand U3901 (N_3901,N_2839,N_2713);
and U3902 (N_3902,N_2863,N_2188);
and U3903 (N_3903,N_2221,N_2690);
and U3904 (N_3904,N_2793,N_2514);
nor U3905 (N_3905,N_2202,N_2888);
and U3906 (N_3906,N_2688,N_2163);
xnor U3907 (N_3907,N_2894,N_2045);
or U3908 (N_3908,N_2499,N_2057);
or U3909 (N_3909,N_2930,N_2833);
xnor U3910 (N_3910,N_2068,N_2867);
nand U3911 (N_3911,N_2383,N_2982);
and U3912 (N_3912,N_2258,N_2938);
and U3913 (N_3913,N_2359,N_2287);
nor U3914 (N_3914,N_2887,N_2962);
xor U3915 (N_3915,N_2512,N_2284);
and U3916 (N_3916,N_2309,N_2708);
nand U3917 (N_3917,N_2961,N_2152);
and U3918 (N_3918,N_2238,N_2790);
nor U3919 (N_3919,N_2608,N_2988);
xor U3920 (N_3920,N_2851,N_2241);
nand U3921 (N_3921,N_2254,N_2594);
or U3922 (N_3922,N_2075,N_2489);
nor U3923 (N_3923,N_2115,N_2819);
and U3924 (N_3924,N_2706,N_2640);
xnor U3925 (N_3925,N_2817,N_2093);
and U3926 (N_3926,N_2640,N_2364);
or U3927 (N_3927,N_2220,N_2354);
nor U3928 (N_3928,N_2310,N_2597);
nor U3929 (N_3929,N_2386,N_2688);
nand U3930 (N_3930,N_2140,N_2714);
or U3931 (N_3931,N_2659,N_2044);
or U3932 (N_3932,N_2795,N_2824);
nand U3933 (N_3933,N_2789,N_2256);
nor U3934 (N_3934,N_2448,N_2487);
nand U3935 (N_3935,N_2066,N_2950);
or U3936 (N_3936,N_2221,N_2679);
nand U3937 (N_3937,N_2432,N_2598);
or U3938 (N_3938,N_2295,N_2155);
nor U3939 (N_3939,N_2307,N_2446);
or U3940 (N_3940,N_2189,N_2417);
nand U3941 (N_3941,N_2579,N_2910);
xnor U3942 (N_3942,N_2620,N_2787);
nand U3943 (N_3943,N_2264,N_2635);
nor U3944 (N_3944,N_2706,N_2936);
or U3945 (N_3945,N_2178,N_2633);
nor U3946 (N_3946,N_2102,N_2263);
and U3947 (N_3947,N_2022,N_2120);
or U3948 (N_3948,N_2348,N_2093);
nor U3949 (N_3949,N_2320,N_2570);
nor U3950 (N_3950,N_2259,N_2247);
or U3951 (N_3951,N_2212,N_2703);
nor U3952 (N_3952,N_2592,N_2137);
nor U3953 (N_3953,N_2157,N_2533);
or U3954 (N_3954,N_2216,N_2794);
nand U3955 (N_3955,N_2583,N_2081);
nor U3956 (N_3956,N_2325,N_2490);
and U3957 (N_3957,N_2653,N_2057);
and U3958 (N_3958,N_2137,N_2118);
and U3959 (N_3959,N_2012,N_2692);
nand U3960 (N_3960,N_2529,N_2030);
nand U3961 (N_3961,N_2225,N_2398);
and U3962 (N_3962,N_2479,N_2976);
or U3963 (N_3963,N_2692,N_2903);
nand U3964 (N_3964,N_2968,N_2939);
or U3965 (N_3965,N_2234,N_2486);
nand U3966 (N_3966,N_2738,N_2371);
nor U3967 (N_3967,N_2171,N_2468);
or U3968 (N_3968,N_2448,N_2989);
nor U3969 (N_3969,N_2444,N_2701);
nor U3970 (N_3970,N_2320,N_2499);
nor U3971 (N_3971,N_2599,N_2687);
or U3972 (N_3972,N_2078,N_2332);
nor U3973 (N_3973,N_2164,N_2724);
nor U3974 (N_3974,N_2809,N_2067);
nor U3975 (N_3975,N_2002,N_2258);
or U3976 (N_3976,N_2655,N_2759);
nand U3977 (N_3977,N_2394,N_2815);
nand U3978 (N_3978,N_2354,N_2716);
nand U3979 (N_3979,N_2091,N_2924);
or U3980 (N_3980,N_2305,N_2330);
nand U3981 (N_3981,N_2986,N_2047);
nand U3982 (N_3982,N_2655,N_2731);
nand U3983 (N_3983,N_2106,N_2029);
nand U3984 (N_3984,N_2532,N_2135);
or U3985 (N_3985,N_2264,N_2590);
nor U3986 (N_3986,N_2186,N_2890);
and U3987 (N_3987,N_2300,N_2937);
nor U3988 (N_3988,N_2574,N_2830);
or U3989 (N_3989,N_2441,N_2566);
nand U3990 (N_3990,N_2920,N_2175);
nand U3991 (N_3991,N_2581,N_2762);
and U3992 (N_3992,N_2907,N_2665);
nand U3993 (N_3993,N_2652,N_2645);
and U3994 (N_3994,N_2126,N_2152);
or U3995 (N_3995,N_2761,N_2960);
nand U3996 (N_3996,N_2328,N_2779);
nor U3997 (N_3997,N_2245,N_2960);
nand U3998 (N_3998,N_2808,N_2782);
or U3999 (N_3999,N_2623,N_2781);
and U4000 (N_4000,N_3084,N_3058);
nand U4001 (N_4001,N_3898,N_3694);
and U4002 (N_4002,N_3813,N_3165);
and U4003 (N_4003,N_3782,N_3386);
xor U4004 (N_4004,N_3465,N_3932);
and U4005 (N_4005,N_3013,N_3558);
nor U4006 (N_4006,N_3327,N_3766);
and U4007 (N_4007,N_3841,N_3969);
or U4008 (N_4008,N_3296,N_3714);
nand U4009 (N_4009,N_3721,N_3475);
nand U4010 (N_4010,N_3651,N_3306);
or U4011 (N_4011,N_3248,N_3147);
or U4012 (N_4012,N_3685,N_3307);
nand U4013 (N_4013,N_3647,N_3487);
and U4014 (N_4014,N_3679,N_3463);
or U4015 (N_4015,N_3482,N_3047);
and U4016 (N_4016,N_3895,N_3676);
xnor U4017 (N_4017,N_3731,N_3748);
and U4018 (N_4018,N_3590,N_3967);
or U4019 (N_4019,N_3501,N_3508);
nor U4020 (N_4020,N_3717,N_3314);
nand U4021 (N_4021,N_3191,N_3571);
nand U4022 (N_4022,N_3597,N_3493);
nand U4023 (N_4023,N_3411,N_3078);
nor U4024 (N_4024,N_3933,N_3010);
or U4025 (N_4025,N_3071,N_3308);
xnor U4026 (N_4026,N_3427,N_3228);
nand U4027 (N_4027,N_3613,N_3910);
nand U4028 (N_4028,N_3509,N_3915);
nand U4029 (N_4029,N_3178,N_3189);
nor U4030 (N_4030,N_3018,N_3061);
or U4031 (N_4031,N_3123,N_3213);
or U4032 (N_4032,N_3658,N_3513);
or U4033 (N_4033,N_3347,N_3890);
nand U4034 (N_4034,N_3335,N_3575);
and U4035 (N_4035,N_3741,N_3941);
and U4036 (N_4036,N_3049,N_3008);
and U4037 (N_4037,N_3469,N_3989);
nand U4038 (N_4038,N_3311,N_3626);
xor U4039 (N_4039,N_3938,N_3863);
nor U4040 (N_4040,N_3510,N_3461);
or U4041 (N_4041,N_3977,N_3958);
or U4042 (N_4042,N_3615,N_3838);
and U4043 (N_4043,N_3081,N_3170);
nand U4044 (N_4044,N_3065,N_3090);
or U4045 (N_4045,N_3979,N_3420);
nor U4046 (N_4046,N_3003,N_3075);
nand U4047 (N_4047,N_3210,N_3288);
nor U4048 (N_4048,N_3168,N_3323);
nand U4049 (N_4049,N_3947,N_3569);
and U4050 (N_4050,N_3784,N_3754);
and U4051 (N_4051,N_3552,N_3579);
nand U4052 (N_4052,N_3543,N_3177);
or U4053 (N_4053,N_3230,N_3141);
nor U4054 (N_4054,N_3423,N_3856);
and U4055 (N_4055,N_3542,N_3346);
nand U4056 (N_4056,N_3609,N_3183);
or U4057 (N_4057,N_3974,N_3749);
or U4058 (N_4058,N_3247,N_3871);
nor U4059 (N_4059,N_3945,N_3586);
nand U4060 (N_4060,N_3892,N_3269);
nand U4061 (N_4061,N_3968,N_3527);
nor U4062 (N_4062,N_3556,N_3879);
and U4063 (N_4063,N_3039,N_3512);
or U4064 (N_4064,N_3176,N_3921);
or U4065 (N_4065,N_3711,N_3403);
nor U4066 (N_4066,N_3514,N_3037);
nand U4067 (N_4067,N_3117,N_3948);
and U4068 (N_4068,N_3523,N_3873);
xor U4069 (N_4069,N_3393,N_3254);
or U4070 (N_4070,N_3935,N_3361);
nor U4071 (N_4071,N_3855,N_3916);
nand U4072 (N_4072,N_3100,N_3404);
nor U4073 (N_4073,N_3310,N_3326);
or U4074 (N_4074,N_3499,N_3623);
and U4075 (N_4075,N_3229,N_3359);
nand U4076 (N_4076,N_3919,N_3011);
nand U4077 (N_4077,N_3930,N_3038);
nor U4078 (N_4078,N_3407,N_3662);
nor U4079 (N_4079,N_3900,N_3923);
nand U4080 (N_4080,N_3860,N_3004);
nor U4081 (N_4081,N_3829,N_3161);
nor U4082 (N_4082,N_3080,N_3878);
nand U4083 (N_4083,N_3864,N_3857);
nor U4084 (N_4084,N_3196,N_3681);
or U4085 (N_4085,N_3019,N_3724);
and U4086 (N_4086,N_3054,N_3344);
and U4087 (N_4087,N_3227,N_3283);
nor U4088 (N_4088,N_3445,N_3048);
nand U4089 (N_4089,N_3752,N_3688);
and U4090 (N_4090,N_3596,N_3431);
nand U4091 (N_4091,N_3650,N_3972);
and U4092 (N_4092,N_3174,N_3005);
and U4093 (N_4093,N_3204,N_3495);
and U4094 (N_4094,N_3128,N_3264);
nor U4095 (N_4095,N_3365,N_3743);
or U4096 (N_4096,N_3554,N_3888);
nand U4097 (N_4097,N_3608,N_3056);
nor U4098 (N_4098,N_3663,N_3492);
and U4099 (N_4099,N_3628,N_3937);
or U4100 (N_4100,N_3524,N_3810);
or U4101 (N_4101,N_3237,N_3985);
nor U4102 (N_4102,N_3376,N_3113);
nand U4103 (N_4103,N_3153,N_3506);
nor U4104 (N_4104,N_3066,N_3118);
nor U4105 (N_4105,N_3238,N_3925);
xnor U4106 (N_4106,N_3295,N_3397);
nor U4107 (N_4107,N_3671,N_3400);
and U4108 (N_4108,N_3374,N_3821);
or U4109 (N_4109,N_3394,N_3106);
nor U4110 (N_4110,N_3631,N_3127);
nor U4111 (N_4111,N_3576,N_3203);
or U4112 (N_4112,N_3819,N_3618);
xnor U4113 (N_4113,N_3740,N_3601);
nand U4114 (N_4114,N_3534,N_3126);
or U4115 (N_4115,N_3162,N_3978);
and U4116 (N_4116,N_3578,N_3529);
nand U4117 (N_4117,N_3886,N_3073);
nand U4118 (N_4118,N_3466,N_3755);
or U4119 (N_4119,N_3836,N_3927);
nor U4120 (N_4120,N_3040,N_3520);
nor U4121 (N_4121,N_3758,N_3866);
and U4122 (N_4122,N_3336,N_3707);
and U4123 (N_4123,N_3896,N_3846);
nand U4124 (N_4124,N_3151,N_3515);
nor U4125 (N_4125,N_3762,N_3622);
nor U4126 (N_4126,N_3158,N_3555);
and U4127 (N_4127,N_3472,N_3239);
nand U4128 (N_4128,N_3635,N_3322);
or U4129 (N_4129,N_3425,N_3481);
nand U4130 (N_4130,N_3187,N_3715);
nor U4131 (N_4131,N_3774,N_3457);
nor U4132 (N_4132,N_3190,N_3259);
and U4133 (N_4133,N_3442,N_3253);
and U4134 (N_4134,N_3994,N_3451);
and U4135 (N_4135,N_3192,N_3936);
or U4136 (N_4136,N_3250,N_3928);
and U4137 (N_4137,N_3258,N_3876);
nor U4138 (N_4138,N_3496,N_3324);
and U4139 (N_4139,N_3991,N_3175);
nand U4140 (N_4140,N_3562,N_3124);
or U4141 (N_4141,N_3353,N_3212);
and U4142 (N_4142,N_3450,N_3318);
nor U4143 (N_4143,N_3889,N_3998);
nor U4144 (N_4144,N_3130,N_3231);
nand U4145 (N_4145,N_3728,N_3949);
nand U4146 (N_4146,N_3242,N_3806);
and U4147 (N_4147,N_3030,N_3447);
or U4148 (N_4148,N_3435,N_3154);
nand U4149 (N_4149,N_3918,N_3455);
and U4150 (N_4150,N_3086,N_3036);
or U4151 (N_4151,N_3682,N_3800);
and U4152 (N_4152,N_3480,N_3497);
or U4153 (N_4153,N_3379,N_3788);
or U4154 (N_4154,N_3720,N_3845);
nand U4155 (N_4155,N_3697,N_3104);
or U4156 (N_4156,N_3537,N_3870);
nand U4157 (N_4157,N_3753,N_3587);
or U4158 (N_4158,N_3517,N_3216);
nor U4159 (N_4159,N_3677,N_3751);
and U4160 (N_4160,N_3279,N_3026);
or U4161 (N_4161,N_3186,N_3364);
nor U4162 (N_4162,N_3391,N_3068);
or U4163 (N_4163,N_3559,N_3822);
and U4164 (N_4164,N_3478,N_3414);
and U4165 (N_4165,N_3840,N_3598);
nand U4166 (N_4166,N_3275,N_3453);
or U4167 (N_4167,N_3611,N_3419);
xor U4168 (N_4168,N_3332,N_3815);
nor U4169 (N_4169,N_3144,N_3869);
and U4170 (N_4170,N_3438,N_3057);
and U4171 (N_4171,N_3592,N_3799);
and U4172 (N_4172,N_3826,N_3468);
or U4173 (N_4173,N_3486,N_3901);
or U4174 (N_4174,N_3903,N_3444);
nor U4175 (N_4175,N_3764,N_3756);
nand U4176 (N_4176,N_3727,N_3792);
nand U4177 (N_4177,N_3834,N_3603);
and U4178 (N_4178,N_3348,N_3265);
nor U4179 (N_4179,N_3546,N_3441);
nand U4180 (N_4180,N_3612,N_3827);
nand U4181 (N_4181,N_3767,N_3287);
nor U4182 (N_4182,N_3561,N_3368);
nand U4183 (N_4183,N_3640,N_3820);
nor U4184 (N_4184,N_3331,N_3433);
and U4185 (N_4185,N_3255,N_3405);
or U4186 (N_4186,N_3745,N_3140);
or U4187 (N_4187,N_3732,N_3730);
nor U4188 (N_4188,N_3415,N_3260);
and U4189 (N_4189,N_3350,N_3803);
nor U4190 (N_4190,N_3645,N_3459);
nand U4191 (N_4191,N_3595,N_3408);
nand U4192 (N_4192,N_3341,N_3023);
nor U4193 (N_4193,N_3528,N_3675);
nand U4194 (N_4194,N_3135,N_3725);
nand U4195 (N_4195,N_3678,N_3354);
nor U4196 (N_4196,N_3027,N_3297);
nand U4197 (N_4197,N_3891,N_3665);
xnor U4198 (N_4198,N_3470,N_3795);
nor U4199 (N_4199,N_3567,N_3772);
nand U4200 (N_4200,N_3851,N_3990);
xnor U4201 (N_4201,N_3853,N_3179);
and U4202 (N_4202,N_3533,N_3961);
or U4203 (N_4203,N_3302,N_3103);
nor U4204 (N_4204,N_3156,N_3125);
nand U4205 (N_4205,N_3548,N_3723);
or U4206 (N_4206,N_3074,N_3001);
and U4207 (N_4207,N_3050,N_3245);
nand U4208 (N_4208,N_3842,N_3808);
or U4209 (N_4209,N_3538,N_3959);
nor U4210 (N_4210,N_3121,N_3096);
or U4211 (N_4211,N_3389,N_3739);
or U4212 (N_4212,N_3284,N_3416);
and U4213 (N_4213,N_3807,N_3794);
and U4214 (N_4214,N_3747,N_3594);
or U4215 (N_4215,N_3219,N_3164);
and U4216 (N_4216,N_3695,N_3002);
nor U4217 (N_4217,N_3600,N_3865);
nand U4218 (N_4218,N_3252,N_3584);
nand U4219 (N_4219,N_3356,N_3309);
xor U4220 (N_4220,N_3518,N_3837);
or U4221 (N_4221,N_3588,N_3396);
and U4222 (N_4222,N_3046,N_3022);
nor U4223 (N_4223,N_3181,N_3966);
and U4224 (N_4224,N_3913,N_3217);
nor U4225 (N_4225,N_3021,N_3885);
nor U4226 (N_4226,N_3012,N_3377);
or U4227 (N_4227,N_3098,N_3102);
and U4228 (N_4228,N_3312,N_3363);
or U4229 (N_4229,N_3484,N_3271);
nand U4230 (N_4230,N_3643,N_3236);
nor U4231 (N_4231,N_3564,N_3041);
nand U4232 (N_4232,N_3340,N_3964);
or U4233 (N_4233,N_3184,N_3105);
nor U4234 (N_4234,N_3642,N_3796);
nor U4235 (N_4235,N_3610,N_3536);
nand U4236 (N_4236,N_3654,N_3693);
or U4237 (N_4237,N_3883,N_3244);
and U4238 (N_4238,N_3067,N_3850);
and U4239 (N_4239,N_3372,N_3630);
and U4240 (N_4240,N_3462,N_3063);
nand U4241 (N_4241,N_3490,N_3540);
or U4242 (N_4242,N_3769,N_3568);
nand U4243 (N_4243,N_3224,N_3294);
nand U4244 (N_4244,N_3045,N_3059);
nor U4245 (N_4245,N_3222,N_3342);
nor U4246 (N_4246,N_3549,N_3976);
and U4247 (N_4247,N_3395,N_3718);
nand U4248 (N_4248,N_3273,N_3726);
and U4249 (N_4249,N_3494,N_3163);
nor U4250 (N_4250,N_3648,N_3198);
nand U4251 (N_4251,N_3778,N_3735);
or U4252 (N_4252,N_3914,N_3383);
or U4253 (N_4253,N_3378,N_3032);
nor U4254 (N_4254,N_3634,N_3706);
or U4255 (N_4255,N_3182,N_3235);
nand U4256 (N_4256,N_3384,N_3303);
nand U4257 (N_4257,N_3737,N_3894);
nor U4258 (N_4258,N_3020,N_3722);
nor U4259 (N_4259,N_3290,N_3240);
or U4260 (N_4260,N_3861,N_3070);
nand U4261 (N_4261,N_3315,N_3401);
or U4262 (N_4262,N_3452,N_3924);
and U4263 (N_4263,N_3076,N_3996);
nor U4264 (N_4264,N_3884,N_3009);
and U4265 (N_4265,N_3757,N_3926);
nor U4266 (N_4266,N_3031,N_3101);
nand U4267 (N_4267,N_3355,N_3114);
or U4268 (N_4268,N_3744,N_3907);
nand U4269 (N_4269,N_3984,N_3698);
or U4270 (N_4270,N_3607,N_3893);
nor U4271 (N_4271,N_3300,N_3025);
nand U4272 (N_4272,N_3828,N_3357);
xnor U4273 (N_4273,N_3491,N_3656);
and U4274 (N_4274,N_3006,N_3809);
nor U4275 (N_4275,N_3670,N_3370);
and U4276 (N_4276,N_3565,N_3768);
nand U4277 (N_4277,N_3188,N_3051);
or U4278 (N_4278,N_3691,N_3360);
or U4279 (N_4279,N_3708,N_3793);
nand U4280 (N_4280,N_3316,N_3781);
nand U4281 (N_4281,N_3385,N_3358);
nor U4282 (N_4282,N_3818,N_3251);
nand U4283 (N_4283,N_3659,N_3897);
nor U4284 (N_4284,N_3215,N_3166);
xnor U4285 (N_4285,N_3146,N_3970);
or U4286 (N_4286,N_3313,N_3811);
nand U4287 (N_4287,N_3077,N_3805);
nor U4288 (N_4288,N_3193,N_3646);
nor U4289 (N_4289,N_3773,N_3485);
or U4290 (N_4290,N_3133,N_3798);
or U4291 (N_4291,N_3145,N_3167);
or U4292 (N_4292,N_3952,N_3729);
nand U4293 (N_4293,N_3330,N_3432);
and U4294 (N_4294,N_3232,N_3657);
or U4295 (N_4295,N_3489,N_3017);
or U4296 (N_4296,N_3687,N_3097);
or U4297 (N_4297,N_3507,N_3881);
nand U4298 (N_4298,N_3713,N_3849);
and U4299 (N_4299,N_3987,N_3911);
and U4300 (N_4300,N_3566,N_3142);
nor U4301 (N_4301,N_3424,N_3007);
and U4302 (N_4302,N_3701,N_3931);
or U4303 (N_4303,N_3877,N_3940);
and U4304 (N_4304,N_3553,N_3993);
or U4305 (N_4305,N_3627,N_3243);
nand U4306 (N_4306,N_3093,N_3522);
or U4307 (N_4307,N_3624,N_3477);
or U4308 (N_4308,N_3434,N_3333);
and U4309 (N_4309,N_3488,N_3843);
and U4310 (N_4310,N_3476,N_3334);
or U4311 (N_4311,N_3995,N_3234);
nor U4312 (N_4312,N_3418,N_3015);
and U4313 (N_4313,N_3814,N_3734);
and U4314 (N_4314,N_3787,N_3282);
nand U4315 (N_4315,N_3632,N_3044);
and U4316 (N_4316,N_3636,N_3351);
nor U4317 (N_4317,N_3917,N_3625);
and U4318 (N_4318,N_3317,N_3502);
nor U4319 (N_4319,N_3859,N_3443);
or U4320 (N_4320,N_3249,N_3220);
nor U4321 (N_4321,N_3973,N_3109);
nand U4322 (N_4322,N_3581,N_3352);
nor U4323 (N_4323,N_3412,N_3115);
or U4324 (N_4324,N_3205,N_3209);
and U4325 (N_4325,N_3131,N_3053);
nand U4326 (N_4326,N_3362,N_3211);
or U4327 (N_4327,N_3942,N_3902);
or U4328 (N_4328,N_3573,N_3652);
and U4329 (N_4329,N_3226,N_3899);
and U4330 (N_4330,N_3338,N_3110);
and U4331 (N_4331,N_3844,N_3399);
and U4332 (N_4332,N_3912,N_3583);
nor U4333 (N_4333,N_3329,N_3906);
and U4334 (N_4334,N_3272,N_3882);
nand U4335 (N_4335,N_3771,N_3129);
nand U4336 (N_4336,N_3975,N_3464);
or U4337 (N_4337,N_3526,N_3847);
nand U4338 (N_4338,N_3684,N_3206);
nand U4339 (N_4339,N_3505,N_3421);
or U4340 (N_4340,N_3939,N_3950);
nand U4341 (N_4341,N_3388,N_3137);
nand U4342 (N_4342,N_3957,N_3664);
or U4343 (N_4343,N_3270,N_3208);
nor U4344 (N_4344,N_3256,N_3280);
or U4345 (N_4345,N_3325,N_3577);
nor U4346 (N_4346,N_3817,N_3835);
nor U4347 (N_4347,N_3298,N_3742);
or U4348 (N_4348,N_3667,N_3980);
nand U4349 (N_4349,N_3560,N_3500);
xor U4350 (N_4350,N_3875,N_3458);
or U4351 (N_4351,N_3276,N_3172);
and U4352 (N_4352,N_3381,N_3511);
nand U4353 (N_4353,N_3880,N_3981);
nand U4354 (N_4354,N_3572,N_3733);
or U4355 (N_4355,N_3922,N_3719);
nor U4356 (N_4356,N_3825,N_3088);
or U4357 (N_4357,N_3199,N_3159);
or U4358 (N_4358,N_3417,N_3079);
or U4359 (N_4359,N_3152,N_3690);
or U4360 (N_4360,N_3997,N_3904);
and U4361 (N_4361,N_3149,N_3956);
and U4362 (N_4362,N_3321,N_3644);
and U4363 (N_4363,N_3095,N_3551);
or U4364 (N_4364,N_3083,N_3532);
nor U4365 (N_4365,N_3868,N_3233);
or U4366 (N_4366,N_3136,N_3965);
nor U4367 (N_4367,N_3770,N_3483);
and U4368 (N_4368,N_3962,N_3872);
xnor U4369 (N_4369,N_3703,N_3301);
or U4370 (N_4370,N_3413,N_3519);
and U4371 (N_4371,N_3789,N_3402);
nand U4372 (N_4372,N_3390,N_3563);
and U4373 (N_4373,N_3446,N_3775);
nor U4374 (N_4374,N_3448,N_3591);
or U4375 (N_4375,N_3014,N_3689);
nor U4376 (N_4376,N_3779,N_3620);
nand U4377 (N_4377,N_3160,N_3440);
nor U4378 (N_4378,N_3171,N_3069);
or U4379 (N_4379,N_3791,N_3197);
xor U4380 (N_4380,N_3954,N_3200);
or U4381 (N_4381,N_3557,N_3367);
nand U4382 (N_4382,N_3530,N_3305);
nor U4383 (N_4383,N_3429,N_3736);
nand U4384 (N_4384,N_3746,N_3261);
nor U4385 (N_4385,N_3143,N_3262);
nor U4386 (N_4386,N_3138,N_3328);
and U4387 (N_4387,N_3674,N_3833);
nor U4388 (N_4388,N_3366,N_3293);
nand U4389 (N_4389,N_3139,N_3765);
and U4390 (N_4390,N_3202,N_3375);
or U4391 (N_4391,N_3278,N_3862);
nand U4392 (N_4392,N_3373,N_3241);
xor U4393 (N_4393,N_3060,N_3428);
nand U4394 (N_4394,N_3544,N_3369);
nor U4395 (N_4395,N_3908,N_3426);
or U4396 (N_4396,N_3982,N_3042);
and U4397 (N_4397,N_3029,N_3812);
or U4398 (N_4398,N_3503,N_3602);
nor U4399 (N_4399,N_3092,N_3382);
and U4400 (N_4400,N_3763,N_3132);
and U4401 (N_4401,N_3525,N_3207);
nor U4402 (N_4402,N_3951,N_3673);
and U4403 (N_4403,N_3195,N_3797);
or U4404 (N_4404,N_3712,N_3804);
nor U4405 (N_4405,N_3194,N_3541);
and U4406 (N_4406,N_3286,N_3830);
nor U4407 (N_4407,N_3479,N_3289);
nor U4408 (N_4408,N_3122,N_3593);
nand U4409 (N_4409,N_3638,N_3672);
nor U4410 (N_4410,N_3988,N_3831);
and U4411 (N_4411,N_3649,N_3705);
nand U4412 (N_4412,N_3055,N_3460);
nand U4413 (N_4413,N_3535,N_3641);
or U4414 (N_4414,N_3218,N_3946);
or U4415 (N_4415,N_3802,N_3043);
nand U4416 (N_4416,N_3823,N_3173);
or U4417 (N_4417,N_3589,N_3983);
and U4418 (N_4418,N_3380,N_3574);
nand U4419 (N_4419,N_3692,N_3449);
and U4420 (N_4420,N_3606,N_3339);
xor U4421 (N_4421,N_3150,N_3999);
and U4422 (N_4422,N_3867,N_3225);
nand U4423 (N_4423,N_3436,N_3454);
or U4424 (N_4424,N_3016,N_3304);
or U4425 (N_4425,N_3082,N_3201);
and U4426 (N_4426,N_3277,N_3274);
nand U4427 (N_4427,N_3858,N_3848);
nand U4428 (N_4428,N_3091,N_3089);
and U4429 (N_4429,N_3474,N_3680);
or U4430 (N_4430,N_3221,N_3854);
xnor U4431 (N_4431,N_3874,N_3666);
or U4432 (N_4432,N_3920,N_3299);
nand U4433 (N_4433,N_3157,N_3349);
nand U4434 (N_4434,N_3521,N_3406);
nor U4435 (N_4435,N_3852,N_3467);
nand U4436 (N_4436,N_3545,N_3909);
and U4437 (N_4437,N_3887,N_3777);
and U4438 (N_4438,N_3409,N_3944);
nand U4439 (N_4439,N_3292,N_3437);
xnor U4440 (N_4440,N_3824,N_3761);
nor U4441 (N_4441,N_3345,N_3619);
nor U4442 (N_4442,N_3291,N_3780);
nand U4443 (N_4443,N_3704,N_3085);
nor U4444 (N_4444,N_3320,N_3816);
or U4445 (N_4445,N_3257,N_3072);
and U4446 (N_4446,N_3268,N_3637);
nand U4447 (N_4447,N_3439,N_3738);
or U4448 (N_4448,N_3547,N_3783);
nor U4449 (N_4449,N_3832,N_3786);
and U4450 (N_4450,N_3034,N_3702);
or U4451 (N_4451,N_3599,N_3052);
nand U4452 (N_4452,N_3653,N_3992);
and U4453 (N_4453,N_3108,N_3148);
or U4454 (N_4454,N_3929,N_3953);
and U4455 (N_4455,N_3986,N_3617);
nand U4456 (N_4456,N_3760,N_3516);
and U4457 (N_4457,N_3683,N_3539);
or U4458 (N_4458,N_3621,N_3614);
and U4459 (N_4459,N_3639,N_3759);
or U4460 (N_4460,N_3776,N_3629);
nor U4461 (N_4461,N_3319,N_3686);
nor U4462 (N_4462,N_3116,N_3422);
nand U4463 (N_4463,N_3266,N_3582);
nand U4464 (N_4464,N_3223,N_3585);
nand U4465 (N_4465,N_3267,N_3668);
nand U4466 (N_4466,N_3387,N_3471);
and U4467 (N_4467,N_3633,N_3000);
or U4468 (N_4468,N_3696,N_3430);
and U4469 (N_4469,N_3398,N_3661);
or U4470 (N_4470,N_3963,N_3099);
nand U4471 (N_4471,N_3246,N_3710);
nor U4472 (N_4472,N_3111,N_3033);
and U4473 (N_4473,N_3655,N_3960);
nand U4474 (N_4474,N_3498,N_3028);
nand U4475 (N_4475,N_3185,N_3580);
or U4476 (N_4476,N_3371,N_3155);
and U4477 (N_4477,N_3660,N_3699);
and U4478 (N_4478,N_3616,N_3112);
nand U4479 (N_4479,N_3955,N_3550);
and U4480 (N_4480,N_3281,N_3790);
nand U4481 (N_4481,N_3107,N_3905);
nor U4482 (N_4482,N_3971,N_3180);
xor U4483 (N_4483,N_3024,N_3669);
xnor U4484 (N_4484,N_3750,N_3570);
nand U4485 (N_4485,N_3943,N_3801);
nand U4486 (N_4486,N_3263,N_3473);
or U4487 (N_4487,N_3716,N_3035);
nor U4488 (N_4488,N_3214,N_3531);
or U4489 (N_4489,N_3785,N_3062);
and U4490 (N_4490,N_3839,N_3709);
nor U4491 (N_4491,N_3410,N_3094);
and U4492 (N_4492,N_3087,N_3343);
nand U4493 (N_4493,N_3064,N_3285);
nand U4494 (N_4494,N_3119,N_3700);
nand U4495 (N_4495,N_3934,N_3337);
and U4496 (N_4496,N_3605,N_3504);
xnor U4497 (N_4497,N_3456,N_3134);
or U4498 (N_4498,N_3169,N_3120);
and U4499 (N_4499,N_3604,N_3392);
or U4500 (N_4500,N_3489,N_3131);
nand U4501 (N_4501,N_3914,N_3501);
nand U4502 (N_4502,N_3324,N_3522);
nand U4503 (N_4503,N_3329,N_3746);
xnor U4504 (N_4504,N_3768,N_3353);
nand U4505 (N_4505,N_3168,N_3712);
or U4506 (N_4506,N_3792,N_3721);
nand U4507 (N_4507,N_3699,N_3820);
or U4508 (N_4508,N_3397,N_3681);
and U4509 (N_4509,N_3957,N_3055);
nand U4510 (N_4510,N_3672,N_3957);
nor U4511 (N_4511,N_3679,N_3054);
nand U4512 (N_4512,N_3094,N_3535);
nand U4513 (N_4513,N_3701,N_3680);
xor U4514 (N_4514,N_3071,N_3212);
and U4515 (N_4515,N_3377,N_3893);
or U4516 (N_4516,N_3216,N_3620);
nand U4517 (N_4517,N_3764,N_3527);
and U4518 (N_4518,N_3882,N_3374);
and U4519 (N_4519,N_3418,N_3464);
nand U4520 (N_4520,N_3794,N_3429);
or U4521 (N_4521,N_3330,N_3409);
xor U4522 (N_4522,N_3992,N_3710);
nor U4523 (N_4523,N_3107,N_3645);
nor U4524 (N_4524,N_3552,N_3307);
nand U4525 (N_4525,N_3201,N_3061);
xnor U4526 (N_4526,N_3860,N_3965);
nand U4527 (N_4527,N_3408,N_3964);
and U4528 (N_4528,N_3798,N_3850);
or U4529 (N_4529,N_3845,N_3903);
and U4530 (N_4530,N_3755,N_3229);
nand U4531 (N_4531,N_3013,N_3213);
or U4532 (N_4532,N_3318,N_3798);
nand U4533 (N_4533,N_3327,N_3341);
or U4534 (N_4534,N_3025,N_3944);
nor U4535 (N_4535,N_3570,N_3384);
nand U4536 (N_4536,N_3544,N_3518);
nor U4537 (N_4537,N_3660,N_3240);
nor U4538 (N_4538,N_3771,N_3785);
and U4539 (N_4539,N_3917,N_3730);
nor U4540 (N_4540,N_3025,N_3479);
nor U4541 (N_4541,N_3878,N_3211);
and U4542 (N_4542,N_3968,N_3029);
or U4543 (N_4543,N_3851,N_3647);
nor U4544 (N_4544,N_3696,N_3335);
and U4545 (N_4545,N_3800,N_3665);
nand U4546 (N_4546,N_3966,N_3401);
nand U4547 (N_4547,N_3189,N_3134);
and U4548 (N_4548,N_3955,N_3272);
or U4549 (N_4549,N_3546,N_3996);
nand U4550 (N_4550,N_3834,N_3632);
or U4551 (N_4551,N_3103,N_3692);
or U4552 (N_4552,N_3366,N_3405);
and U4553 (N_4553,N_3418,N_3100);
or U4554 (N_4554,N_3259,N_3252);
and U4555 (N_4555,N_3990,N_3009);
nor U4556 (N_4556,N_3603,N_3213);
nand U4557 (N_4557,N_3869,N_3312);
and U4558 (N_4558,N_3202,N_3768);
and U4559 (N_4559,N_3486,N_3717);
and U4560 (N_4560,N_3493,N_3720);
or U4561 (N_4561,N_3490,N_3593);
nor U4562 (N_4562,N_3884,N_3551);
nand U4563 (N_4563,N_3800,N_3013);
nor U4564 (N_4564,N_3641,N_3927);
or U4565 (N_4565,N_3680,N_3805);
nor U4566 (N_4566,N_3845,N_3640);
or U4567 (N_4567,N_3134,N_3702);
nand U4568 (N_4568,N_3688,N_3757);
and U4569 (N_4569,N_3773,N_3402);
and U4570 (N_4570,N_3601,N_3651);
nand U4571 (N_4571,N_3218,N_3390);
or U4572 (N_4572,N_3073,N_3867);
nand U4573 (N_4573,N_3997,N_3778);
or U4574 (N_4574,N_3134,N_3697);
nand U4575 (N_4575,N_3805,N_3237);
or U4576 (N_4576,N_3770,N_3897);
and U4577 (N_4577,N_3591,N_3034);
nor U4578 (N_4578,N_3255,N_3743);
and U4579 (N_4579,N_3427,N_3660);
nand U4580 (N_4580,N_3367,N_3186);
and U4581 (N_4581,N_3311,N_3377);
or U4582 (N_4582,N_3546,N_3371);
and U4583 (N_4583,N_3241,N_3051);
and U4584 (N_4584,N_3794,N_3132);
nor U4585 (N_4585,N_3856,N_3336);
xor U4586 (N_4586,N_3286,N_3816);
nand U4587 (N_4587,N_3099,N_3922);
nor U4588 (N_4588,N_3158,N_3247);
and U4589 (N_4589,N_3707,N_3263);
xor U4590 (N_4590,N_3842,N_3077);
or U4591 (N_4591,N_3631,N_3647);
nor U4592 (N_4592,N_3147,N_3294);
or U4593 (N_4593,N_3644,N_3817);
nand U4594 (N_4594,N_3502,N_3872);
or U4595 (N_4595,N_3263,N_3371);
and U4596 (N_4596,N_3525,N_3014);
and U4597 (N_4597,N_3842,N_3580);
nor U4598 (N_4598,N_3073,N_3950);
nand U4599 (N_4599,N_3070,N_3349);
nand U4600 (N_4600,N_3263,N_3294);
nor U4601 (N_4601,N_3975,N_3370);
nor U4602 (N_4602,N_3029,N_3745);
nor U4603 (N_4603,N_3869,N_3387);
or U4604 (N_4604,N_3986,N_3213);
and U4605 (N_4605,N_3876,N_3438);
or U4606 (N_4606,N_3391,N_3699);
nor U4607 (N_4607,N_3553,N_3864);
and U4608 (N_4608,N_3183,N_3897);
and U4609 (N_4609,N_3841,N_3328);
nor U4610 (N_4610,N_3878,N_3056);
nor U4611 (N_4611,N_3452,N_3509);
or U4612 (N_4612,N_3717,N_3268);
and U4613 (N_4613,N_3983,N_3238);
nor U4614 (N_4614,N_3285,N_3378);
and U4615 (N_4615,N_3871,N_3677);
nand U4616 (N_4616,N_3665,N_3859);
or U4617 (N_4617,N_3703,N_3116);
and U4618 (N_4618,N_3938,N_3591);
nand U4619 (N_4619,N_3856,N_3753);
nor U4620 (N_4620,N_3086,N_3178);
and U4621 (N_4621,N_3253,N_3205);
and U4622 (N_4622,N_3666,N_3635);
and U4623 (N_4623,N_3014,N_3703);
nor U4624 (N_4624,N_3560,N_3813);
nand U4625 (N_4625,N_3635,N_3599);
or U4626 (N_4626,N_3501,N_3863);
and U4627 (N_4627,N_3974,N_3103);
and U4628 (N_4628,N_3971,N_3187);
xor U4629 (N_4629,N_3650,N_3774);
nor U4630 (N_4630,N_3975,N_3112);
and U4631 (N_4631,N_3733,N_3994);
nand U4632 (N_4632,N_3679,N_3291);
xnor U4633 (N_4633,N_3410,N_3688);
and U4634 (N_4634,N_3430,N_3892);
nor U4635 (N_4635,N_3471,N_3202);
nand U4636 (N_4636,N_3348,N_3251);
and U4637 (N_4637,N_3190,N_3722);
or U4638 (N_4638,N_3197,N_3639);
nor U4639 (N_4639,N_3421,N_3033);
nor U4640 (N_4640,N_3815,N_3119);
nor U4641 (N_4641,N_3258,N_3232);
nand U4642 (N_4642,N_3908,N_3235);
or U4643 (N_4643,N_3864,N_3861);
nor U4644 (N_4644,N_3104,N_3456);
nand U4645 (N_4645,N_3472,N_3258);
nand U4646 (N_4646,N_3432,N_3084);
or U4647 (N_4647,N_3264,N_3740);
xnor U4648 (N_4648,N_3081,N_3888);
nor U4649 (N_4649,N_3155,N_3409);
nor U4650 (N_4650,N_3065,N_3973);
and U4651 (N_4651,N_3015,N_3462);
nand U4652 (N_4652,N_3337,N_3267);
nand U4653 (N_4653,N_3816,N_3053);
and U4654 (N_4654,N_3107,N_3007);
and U4655 (N_4655,N_3826,N_3231);
nor U4656 (N_4656,N_3769,N_3375);
nor U4657 (N_4657,N_3895,N_3181);
nand U4658 (N_4658,N_3672,N_3586);
or U4659 (N_4659,N_3993,N_3723);
nand U4660 (N_4660,N_3748,N_3170);
nand U4661 (N_4661,N_3379,N_3257);
or U4662 (N_4662,N_3907,N_3165);
or U4663 (N_4663,N_3673,N_3002);
or U4664 (N_4664,N_3233,N_3874);
and U4665 (N_4665,N_3524,N_3101);
and U4666 (N_4666,N_3729,N_3219);
xor U4667 (N_4667,N_3468,N_3957);
or U4668 (N_4668,N_3626,N_3378);
or U4669 (N_4669,N_3506,N_3231);
and U4670 (N_4670,N_3381,N_3964);
and U4671 (N_4671,N_3496,N_3243);
nand U4672 (N_4672,N_3482,N_3918);
nor U4673 (N_4673,N_3450,N_3803);
nand U4674 (N_4674,N_3284,N_3457);
nand U4675 (N_4675,N_3498,N_3784);
nand U4676 (N_4676,N_3245,N_3258);
nand U4677 (N_4677,N_3244,N_3017);
nor U4678 (N_4678,N_3640,N_3620);
nor U4679 (N_4679,N_3116,N_3500);
or U4680 (N_4680,N_3236,N_3035);
nand U4681 (N_4681,N_3623,N_3982);
and U4682 (N_4682,N_3728,N_3507);
and U4683 (N_4683,N_3446,N_3616);
nand U4684 (N_4684,N_3823,N_3228);
xnor U4685 (N_4685,N_3710,N_3389);
and U4686 (N_4686,N_3899,N_3171);
and U4687 (N_4687,N_3684,N_3098);
nand U4688 (N_4688,N_3066,N_3242);
nand U4689 (N_4689,N_3536,N_3768);
and U4690 (N_4690,N_3725,N_3261);
and U4691 (N_4691,N_3819,N_3456);
nor U4692 (N_4692,N_3093,N_3939);
nor U4693 (N_4693,N_3555,N_3059);
nor U4694 (N_4694,N_3150,N_3962);
and U4695 (N_4695,N_3250,N_3293);
and U4696 (N_4696,N_3489,N_3370);
nor U4697 (N_4697,N_3040,N_3592);
or U4698 (N_4698,N_3705,N_3344);
nand U4699 (N_4699,N_3957,N_3652);
xnor U4700 (N_4700,N_3757,N_3202);
or U4701 (N_4701,N_3971,N_3066);
nor U4702 (N_4702,N_3972,N_3589);
and U4703 (N_4703,N_3064,N_3535);
nor U4704 (N_4704,N_3803,N_3263);
xor U4705 (N_4705,N_3253,N_3108);
and U4706 (N_4706,N_3653,N_3009);
or U4707 (N_4707,N_3098,N_3276);
and U4708 (N_4708,N_3350,N_3493);
nor U4709 (N_4709,N_3999,N_3208);
and U4710 (N_4710,N_3393,N_3395);
nand U4711 (N_4711,N_3890,N_3933);
and U4712 (N_4712,N_3881,N_3139);
or U4713 (N_4713,N_3964,N_3773);
or U4714 (N_4714,N_3721,N_3559);
nor U4715 (N_4715,N_3889,N_3309);
xnor U4716 (N_4716,N_3003,N_3705);
nand U4717 (N_4717,N_3217,N_3296);
nor U4718 (N_4718,N_3822,N_3201);
nor U4719 (N_4719,N_3136,N_3098);
nand U4720 (N_4720,N_3926,N_3137);
nor U4721 (N_4721,N_3501,N_3904);
nand U4722 (N_4722,N_3382,N_3254);
xnor U4723 (N_4723,N_3004,N_3217);
nor U4724 (N_4724,N_3131,N_3949);
nor U4725 (N_4725,N_3528,N_3113);
and U4726 (N_4726,N_3568,N_3339);
or U4727 (N_4727,N_3953,N_3541);
nor U4728 (N_4728,N_3006,N_3217);
nand U4729 (N_4729,N_3875,N_3717);
and U4730 (N_4730,N_3663,N_3681);
and U4731 (N_4731,N_3502,N_3963);
or U4732 (N_4732,N_3777,N_3421);
and U4733 (N_4733,N_3598,N_3843);
nor U4734 (N_4734,N_3132,N_3979);
nand U4735 (N_4735,N_3169,N_3869);
or U4736 (N_4736,N_3931,N_3782);
nor U4737 (N_4737,N_3577,N_3010);
xnor U4738 (N_4738,N_3967,N_3729);
nor U4739 (N_4739,N_3308,N_3781);
and U4740 (N_4740,N_3391,N_3441);
and U4741 (N_4741,N_3097,N_3889);
nand U4742 (N_4742,N_3270,N_3432);
and U4743 (N_4743,N_3648,N_3321);
nor U4744 (N_4744,N_3475,N_3309);
nand U4745 (N_4745,N_3938,N_3840);
or U4746 (N_4746,N_3370,N_3913);
or U4747 (N_4747,N_3045,N_3651);
or U4748 (N_4748,N_3156,N_3084);
nand U4749 (N_4749,N_3319,N_3553);
nand U4750 (N_4750,N_3943,N_3596);
nand U4751 (N_4751,N_3792,N_3580);
or U4752 (N_4752,N_3319,N_3977);
nand U4753 (N_4753,N_3851,N_3152);
nor U4754 (N_4754,N_3879,N_3856);
and U4755 (N_4755,N_3174,N_3831);
nor U4756 (N_4756,N_3575,N_3398);
nor U4757 (N_4757,N_3643,N_3003);
xnor U4758 (N_4758,N_3943,N_3646);
nor U4759 (N_4759,N_3361,N_3354);
nand U4760 (N_4760,N_3926,N_3758);
nor U4761 (N_4761,N_3870,N_3762);
and U4762 (N_4762,N_3008,N_3547);
nor U4763 (N_4763,N_3198,N_3941);
and U4764 (N_4764,N_3698,N_3989);
nor U4765 (N_4765,N_3017,N_3271);
and U4766 (N_4766,N_3395,N_3091);
and U4767 (N_4767,N_3160,N_3159);
and U4768 (N_4768,N_3670,N_3893);
or U4769 (N_4769,N_3472,N_3884);
and U4770 (N_4770,N_3507,N_3522);
nand U4771 (N_4771,N_3942,N_3425);
nand U4772 (N_4772,N_3080,N_3127);
or U4773 (N_4773,N_3478,N_3869);
nor U4774 (N_4774,N_3448,N_3671);
nand U4775 (N_4775,N_3392,N_3536);
and U4776 (N_4776,N_3534,N_3154);
nor U4777 (N_4777,N_3914,N_3395);
and U4778 (N_4778,N_3434,N_3560);
or U4779 (N_4779,N_3271,N_3768);
nand U4780 (N_4780,N_3407,N_3055);
or U4781 (N_4781,N_3100,N_3698);
and U4782 (N_4782,N_3476,N_3985);
and U4783 (N_4783,N_3817,N_3295);
nand U4784 (N_4784,N_3484,N_3406);
or U4785 (N_4785,N_3759,N_3670);
and U4786 (N_4786,N_3153,N_3885);
nor U4787 (N_4787,N_3988,N_3918);
nand U4788 (N_4788,N_3878,N_3091);
nand U4789 (N_4789,N_3525,N_3647);
or U4790 (N_4790,N_3018,N_3319);
or U4791 (N_4791,N_3708,N_3350);
and U4792 (N_4792,N_3792,N_3550);
nor U4793 (N_4793,N_3705,N_3113);
or U4794 (N_4794,N_3198,N_3073);
and U4795 (N_4795,N_3352,N_3276);
nand U4796 (N_4796,N_3370,N_3378);
and U4797 (N_4797,N_3306,N_3162);
nand U4798 (N_4798,N_3990,N_3299);
nand U4799 (N_4799,N_3989,N_3515);
or U4800 (N_4800,N_3684,N_3956);
nor U4801 (N_4801,N_3600,N_3087);
and U4802 (N_4802,N_3074,N_3662);
and U4803 (N_4803,N_3040,N_3311);
nand U4804 (N_4804,N_3073,N_3625);
or U4805 (N_4805,N_3944,N_3091);
nor U4806 (N_4806,N_3703,N_3243);
nand U4807 (N_4807,N_3370,N_3497);
and U4808 (N_4808,N_3951,N_3509);
xor U4809 (N_4809,N_3825,N_3058);
nand U4810 (N_4810,N_3823,N_3408);
and U4811 (N_4811,N_3816,N_3515);
and U4812 (N_4812,N_3155,N_3642);
or U4813 (N_4813,N_3275,N_3324);
and U4814 (N_4814,N_3995,N_3605);
xnor U4815 (N_4815,N_3656,N_3263);
nor U4816 (N_4816,N_3271,N_3074);
and U4817 (N_4817,N_3058,N_3286);
nor U4818 (N_4818,N_3226,N_3426);
and U4819 (N_4819,N_3643,N_3466);
or U4820 (N_4820,N_3609,N_3596);
or U4821 (N_4821,N_3277,N_3901);
nand U4822 (N_4822,N_3761,N_3440);
nor U4823 (N_4823,N_3749,N_3772);
xor U4824 (N_4824,N_3252,N_3040);
and U4825 (N_4825,N_3197,N_3735);
and U4826 (N_4826,N_3646,N_3797);
nand U4827 (N_4827,N_3094,N_3563);
and U4828 (N_4828,N_3324,N_3610);
nand U4829 (N_4829,N_3864,N_3777);
or U4830 (N_4830,N_3362,N_3659);
nand U4831 (N_4831,N_3370,N_3724);
and U4832 (N_4832,N_3516,N_3251);
and U4833 (N_4833,N_3403,N_3183);
nand U4834 (N_4834,N_3412,N_3844);
nor U4835 (N_4835,N_3413,N_3518);
and U4836 (N_4836,N_3288,N_3253);
or U4837 (N_4837,N_3403,N_3099);
xor U4838 (N_4838,N_3131,N_3476);
nor U4839 (N_4839,N_3259,N_3693);
nand U4840 (N_4840,N_3861,N_3741);
and U4841 (N_4841,N_3611,N_3137);
nand U4842 (N_4842,N_3146,N_3567);
nor U4843 (N_4843,N_3495,N_3097);
nand U4844 (N_4844,N_3255,N_3565);
nor U4845 (N_4845,N_3545,N_3953);
nor U4846 (N_4846,N_3188,N_3969);
nor U4847 (N_4847,N_3658,N_3978);
and U4848 (N_4848,N_3079,N_3620);
nor U4849 (N_4849,N_3573,N_3491);
and U4850 (N_4850,N_3558,N_3694);
nor U4851 (N_4851,N_3318,N_3996);
nor U4852 (N_4852,N_3576,N_3985);
and U4853 (N_4853,N_3034,N_3230);
and U4854 (N_4854,N_3103,N_3414);
and U4855 (N_4855,N_3426,N_3900);
nor U4856 (N_4856,N_3649,N_3678);
and U4857 (N_4857,N_3240,N_3428);
and U4858 (N_4858,N_3526,N_3688);
or U4859 (N_4859,N_3554,N_3631);
and U4860 (N_4860,N_3330,N_3136);
and U4861 (N_4861,N_3544,N_3765);
and U4862 (N_4862,N_3142,N_3857);
nand U4863 (N_4863,N_3885,N_3911);
or U4864 (N_4864,N_3253,N_3181);
nor U4865 (N_4865,N_3035,N_3629);
xnor U4866 (N_4866,N_3874,N_3893);
nand U4867 (N_4867,N_3086,N_3755);
nand U4868 (N_4868,N_3579,N_3782);
xor U4869 (N_4869,N_3542,N_3094);
nand U4870 (N_4870,N_3433,N_3386);
nand U4871 (N_4871,N_3204,N_3466);
or U4872 (N_4872,N_3134,N_3931);
nor U4873 (N_4873,N_3208,N_3466);
nor U4874 (N_4874,N_3920,N_3718);
and U4875 (N_4875,N_3093,N_3748);
nand U4876 (N_4876,N_3263,N_3590);
nor U4877 (N_4877,N_3328,N_3570);
or U4878 (N_4878,N_3599,N_3549);
or U4879 (N_4879,N_3838,N_3429);
or U4880 (N_4880,N_3427,N_3962);
nand U4881 (N_4881,N_3162,N_3563);
or U4882 (N_4882,N_3246,N_3160);
nand U4883 (N_4883,N_3001,N_3560);
or U4884 (N_4884,N_3793,N_3951);
or U4885 (N_4885,N_3939,N_3422);
xnor U4886 (N_4886,N_3189,N_3480);
nor U4887 (N_4887,N_3993,N_3036);
nand U4888 (N_4888,N_3014,N_3760);
or U4889 (N_4889,N_3608,N_3565);
or U4890 (N_4890,N_3382,N_3411);
nor U4891 (N_4891,N_3028,N_3119);
nor U4892 (N_4892,N_3160,N_3950);
nor U4893 (N_4893,N_3442,N_3633);
or U4894 (N_4894,N_3596,N_3754);
or U4895 (N_4895,N_3085,N_3767);
nor U4896 (N_4896,N_3035,N_3164);
or U4897 (N_4897,N_3374,N_3309);
or U4898 (N_4898,N_3507,N_3645);
or U4899 (N_4899,N_3804,N_3615);
nor U4900 (N_4900,N_3646,N_3601);
and U4901 (N_4901,N_3253,N_3020);
nand U4902 (N_4902,N_3426,N_3413);
or U4903 (N_4903,N_3945,N_3441);
nor U4904 (N_4904,N_3444,N_3831);
nand U4905 (N_4905,N_3865,N_3583);
nor U4906 (N_4906,N_3894,N_3830);
nand U4907 (N_4907,N_3691,N_3378);
nor U4908 (N_4908,N_3952,N_3175);
nor U4909 (N_4909,N_3896,N_3455);
or U4910 (N_4910,N_3703,N_3654);
nand U4911 (N_4911,N_3677,N_3861);
nor U4912 (N_4912,N_3087,N_3656);
nor U4913 (N_4913,N_3403,N_3011);
nor U4914 (N_4914,N_3507,N_3257);
or U4915 (N_4915,N_3981,N_3445);
or U4916 (N_4916,N_3120,N_3657);
nor U4917 (N_4917,N_3333,N_3706);
nand U4918 (N_4918,N_3095,N_3854);
nand U4919 (N_4919,N_3751,N_3177);
nor U4920 (N_4920,N_3868,N_3157);
or U4921 (N_4921,N_3706,N_3289);
nand U4922 (N_4922,N_3147,N_3999);
nand U4923 (N_4923,N_3855,N_3668);
nor U4924 (N_4924,N_3889,N_3311);
nor U4925 (N_4925,N_3996,N_3801);
nand U4926 (N_4926,N_3405,N_3597);
or U4927 (N_4927,N_3891,N_3679);
or U4928 (N_4928,N_3555,N_3896);
nand U4929 (N_4929,N_3438,N_3644);
or U4930 (N_4930,N_3791,N_3248);
nand U4931 (N_4931,N_3655,N_3387);
or U4932 (N_4932,N_3780,N_3389);
or U4933 (N_4933,N_3728,N_3047);
nand U4934 (N_4934,N_3494,N_3715);
or U4935 (N_4935,N_3670,N_3896);
nor U4936 (N_4936,N_3446,N_3176);
nor U4937 (N_4937,N_3403,N_3859);
nand U4938 (N_4938,N_3156,N_3949);
nor U4939 (N_4939,N_3742,N_3686);
or U4940 (N_4940,N_3082,N_3685);
and U4941 (N_4941,N_3873,N_3434);
and U4942 (N_4942,N_3811,N_3822);
xnor U4943 (N_4943,N_3857,N_3917);
nor U4944 (N_4944,N_3097,N_3506);
nand U4945 (N_4945,N_3100,N_3816);
and U4946 (N_4946,N_3607,N_3686);
xor U4947 (N_4947,N_3311,N_3967);
nor U4948 (N_4948,N_3406,N_3552);
or U4949 (N_4949,N_3458,N_3876);
nand U4950 (N_4950,N_3407,N_3863);
nor U4951 (N_4951,N_3769,N_3893);
and U4952 (N_4952,N_3968,N_3268);
nor U4953 (N_4953,N_3839,N_3598);
or U4954 (N_4954,N_3693,N_3111);
nor U4955 (N_4955,N_3258,N_3051);
nand U4956 (N_4956,N_3822,N_3548);
and U4957 (N_4957,N_3543,N_3041);
nor U4958 (N_4958,N_3205,N_3005);
nand U4959 (N_4959,N_3489,N_3728);
or U4960 (N_4960,N_3585,N_3628);
nor U4961 (N_4961,N_3546,N_3216);
or U4962 (N_4962,N_3668,N_3786);
or U4963 (N_4963,N_3614,N_3479);
nor U4964 (N_4964,N_3325,N_3372);
and U4965 (N_4965,N_3487,N_3260);
nand U4966 (N_4966,N_3423,N_3901);
nor U4967 (N_4967,N_3890,N_3454);
and U4968 (N_4968,N_3432,N_3393);
nand U4969 (N_4969,N_3121,N_3574);
nand U4970 (N_4970,N_3771,N_3533);
and U4971 (N_4971,N_3687,N_3211);
or U4972 (N_4972,N_3425,N_3483);
or U4973 (N_4973,N_3123,N_3675);
nor U4974 (N_4974,N_3652,N_3807);
nor U4975 (N_4975,N_3543,N_3423);
nor U4976 (N_4976,N_3239,N_3853);
nor U4977 (N_4977,N_3288,N_3165);
nor U4978 (N_4978,N_3174,N_3062);
nand U4979 (N_4979,N_3120,N_3042);
and U4980 (N_4980,N_3310,N_3047);
or U4981 (N_4981,N_3059,N_3901);
and U4982 (N_4982,N_3863,N_3921);
and U4983 (N_4983,N_3372,N_3629);
nor U4984 (N_4984,N_3435,N_3106);
nor U4985 (N_4985,N_3733,N_3041);
and U4986 (N_4986,N_3780,N_3422);
or U4987 (N_4987,N_3161,N_3020);
or U4988 (N_4988,N_3548,N_3308);
and U4989 (N_4989,N_3358,N_3060);
nand U4990 (N_4990,N_3919,N_3281);
or U4991 (N_4991,N_3286,N_3146);
nor U4992 (N_4992,N_3824,N_3462);
nand U4993 (N_4993,N_3644,N_3554);
nor U4994 (N_4994,N_3770,N_3596);
nand U4995 (N_4995,N_3796,N_3535);
nor U4996 (N_4996,N_3114,N_3761);
nand U4997 (N_4997,N_3684,N_3574);
nor U4998 (N_4998,N_3755,N_3260);
nand U4999 (N_4999,N_3616,N_3117);
and U5000 (N_5000,N_4934,N_4478);
or U5001 (N_5001,N_4458,N_4674);
and U5002 (N_5002,N_4499,N_4994);
or U5003 (N_5003,N_4689,N_4266);
and U5004 (N_5004,N_4643,N_4144);
nand U5005 (N_5005,N_4972,N_4541);
nor U5006 (N_5006,N_4318,N_4650);
nand U5007 (N_5007,N_4671,N_4420);
nand U5008 (N_5008,N_4071,N_4929);
or U5009 (N_5009,N_4641,N_4280);
xnor U5010 (N_5010,N_4157,N_4899);
or U5011 (N_5011,N_4917,N_4717);
nor U5012 (N_5012,N_4102,N_4881);
or U5013 (N_5013,N_4007,N_4315);
and U5014 (N_5014,N_4445,N_4508);
or U5015 (N_5015,N_4634,N_4750);
nor U5016 (N_5016,N_4698,N_4060);
or U5017 (N_5017,N_4401,N_4854);
or U5018 (N_5018,N_4673,N_4466);
or U5019 (N_5019,N_4287,N_4675);
and U5020 (N_5020,N_4614,N_4774);
nand U5021 (N_5021,N_4577,N_4137);
or U5022 (N_5022,N_4148,N_4164);
nand U5023 (N_5023,N_4762,N_4555);
nand U5024 (N_5024,N_4801,N_4307);
nand U5025 (N_5025,N_4023,N_4233);
and U5026 (N_5026,N_4243,N_4291);
nand U5027 (N_5027,N_4691,N_4259);
nor U5028 (N_5028,N_4639,N_4656);
nand U5029 (N_5029,N_4716,N_4727);
nor U5030 (N_5030,N_4904,N_4652);
nand U5031 (N_5031,N_4820,N_4601);
and U5032 (N_5032,N_4185,N_4624);
nor U5033 (N_5033,N_4228,N_4591);
and U5034 (N_5034,N_4193,N_4200);
nor U5035 (N_5035,N_4524,N_4590);
and U5036 (N_5036,N_4719,N_4460);
or U5037 (N_5037,N_4404,N_4018);
nand U5038 (N_5038,N_4299,N_4089);
nor U5039 (N_5039,N_4501,N_4270);
nand U5040 (N_5040,N_4553,N_4787);
and U5041 (N_5041,N_4852,N_4968);
nand U5042 (N_5042,N_4066,N_4284);
or U5043 (N_5043,N_4003,N_4245);
nand U5044 (N_5044,N_4609,N_4300);
and U5045 (N_5045,N_4561,N_4026);
nor U5046 (N_5046,N_4676,N_4921);
or U5047 (N_5047,N_4608,N_4181);
or U5048 (N_5048,N_4989,N_4394);
and U5049 (N_5049,N_4120,N_4531);
nor U5050 (N_5050,N_4850,N_4887);
or U5051 (N_5051,N_4145,N_4818);
nor U5052 (N_5052,N_4579,N_4724);
or U5053 (N_5053,N_4596,N_4668);
nor U5054 (N_5054,N_4140,N_4384);
or U5055 (N_5055,N_4187,N_4309);
or U5056 (N_5056,N_4283,N_4685);
and U5057 (N_5057,N_4570,N_4225);
nand U5058 (N_5058,N_4482,N_4679);
nor U5059 (N_5059,N_4433,N_4680);
nor U5060 (N_5060,N_4910,N_4043);
and U5061 (N_5061,N_4976,N_4024);
and U5062 (N_5062,N_4021,N_4097);
nor U5063 (N_5063,N_4012,N_4017);
nor U5064 (N_5064,N_4099,N_4034);
nor U5065 (N_5065,N_4432,N_4763);
or U5066 (N_5066,N_4841,N_4327);
nor U5067 (N_5067,N_4878,N_4532);
nand U5068 (N_5068,N_4045,N_4036);
nor U5069 (N_5069,N_4441,N_4585);
nand U5070 (N_5070,N_4895,N_4058);
nand U5071 (N_5071,N_4785,N_4449);
nor U5072 (N_5072,N_4303,N_4336);
or U5073 (N_5073,N_4706,N_4476);
or U5074 (N_5074,N_4825,N_4006);
or U5075 (N_5075,N_4324,N_4901);
and U5076 (N_5076,N_4958,N_4106);
or U5077 (N_5077,N_4393,N_4790);
or U5078 (N_5078,N_4313,N_4397);
or U5079 (N_5079,N_4985,N_4273);
or U5080 (N_5080,N_4407,N_4931);
nand U5081 (N_5081,N_4953,N_4741);
or U5082 (N_5082,N_4169,N_4661);
and U5083 (N_5083,N_4234,N_4778);
or U5084 (N_5084,N_4897,N_4281);
nor U5085 (N_5085,N_4389,N_4035);
and U5086 (N_5086,N_4042,N_4430);
nand U5087 (N_5087,N_4849,N_4578);
and U5088 (N_5088,N_4311,N_4756);
or U5089 (N_5089,N_4919,N_4347);
and U5090 (N_5090,N_4992,N_4076);
and U5091 (N_5091,N_4167,N_4419);
nand U5092 (N_5092,N_4703,N_4831);
and U5093 (N_5093,N_4814,N_4943);
or U5094 (N_5094,N_4571,N_4429);
and U5095 (N_5095,N_4371,N_4344);
nand U5096 (N_5096,N_4782,N_4382);
nand U5097 (N_5097,N_4049,N_4216);
and U5098 (N_5098,N_4132,N_4957);
nor U5099 (N_5099,N_4542,N_4948);
or U5100 (N_5100,N_4069,N_4847);
nand U5101 (N_5101,N_4484,N_4129);
or U5102 (N_5102,N_4644,N_4447);
and U5103 (N_5103,N_4241,N_4010);
and U5104 (N_5104,N_4208,N_4052);
and U5105 (N_5105,N_4437,N_4543);
nor U5106 (N_5106,N_4098,N_4892);
and U5107 (N_5107,N_4960,N_4272);
nand U5108 (N_5108,N_4363,N_4584);
or U5109 (N_5109,N_4574,N_4016);
nor U5110 (N_5110,N_4902,N_4114);
or U5111 (N_5111,N_4222,N_4837);
nor U5112 (N_5112,N_4062,N_4728);
nor U5113 (N_5113,N_4298,N_4343);
and U5114 (N_5114,N_4710,N_4462);
nor U5115 (N_5115,N_4775,N_4356);
or U5116 (N_5116,N_4421,N_4961);
nor U5117 (N_5117,N_4398,N_4970);
nand U5118 (N_5118,N_4323,N_4658);
nor U5119 (N_5119,N_4130,N_4285);
and U5120 (N_5120,N_4370,N_4978);
nor U5121 (N_5121,N_4510,N_4143);
nor U5122 (N_5122,N_4033,N_4088);
nor U5123 (N_5123,N_4802,N_4768);
and U5124 (N_5124,N_4512,N_4304);
nand U5125 (N_5125,N_4594,N_4330);
and U5126 (N_5126,N_4452,N_4568);
nand U5127 (N_5127,N_4166,N_4723);
nor U5128 (N_5128,N_4294,N_4070);
and U5129 (N_5129,N_4456,N_4626);
or U5130 (N_5130,N_4424,N_4411);
nor U5131 (N_5131,N_4332,N_4136);
or U5132 (N_5132,N_4823,N_4075);
nor U5133 (N_5133,N_4400,N_4883);
nor U5134 (N_5134,N_4128,N_4359);
nor U5135 (N_5135,N_4108,N_4158);
or U5136 (N_5136,N_4950,N_4240);
and U5137 (N_5137,N_4282,N_4882);
or U5138 (N_5138,N_4889,N_4559);
or U5139 (N_5139,N_4677,N_4645);
nor U5140 (N_5140,N_4780,N_4073);
or U5141 (N_5141,N_4403,N_4699);
nand U5142 (N_5142,N_4564,N_4939);
or U5143 (N_5143,N_4156,N_4467);
nor U5144 (N_5144,N_4325,N_4615);
or U5145 (N_5145,N_4443,N_4886);
and U5146 (N_5146,N_4457,N_4842);
and U5147 (N_5147,N_4969,N_4736);
and U5148 (N_5148,N_4048,N_4995);
nor U5149 (N_5149,N_4163,N_4505);
or U5150 (N_5150,N_4821,N_4804);
nor U5151 (N_5151,N_4230,N_4172);
or U5152 (N_5152,N_4981,N_4759);
nor U5153 (N_5153,N_4235,N_4515);
nand U5154 (N_5154,N_4681,N_4538);
and U5155 (N_5155,N_4471,N_4748);
and U5156 (N_5156,N_4700,N_4492);
and U5157 (N_5157,N_4204,N_4544);
and U5158 (N_5158,N_4173,N_4548);
nor U5159 (N_5159,N_4552,N_4556);
nand U5160 (N_5160,N_4226,N_4357);
xor U5161 (N_5161,N_4168,N_4055);
nor U5162 (N_5162,N_4253,N_4781);
or U5163 (N_5163,N_4868,N_4388);
nor U5164 (N_5164,N_4117,N_4182);
nand U5165 (N_5165,N_4051,N_4855);
and U5166 (N_5166,N_4924,N_4310);
and U5167 (N_5167,N_4268,N_4326);
nand U5168 (N_5168,N_4227,N_4001);
or U5169 (N_5169,N_4251,N_4475);
and U5170 (N_5170,N_4378,N_4722);
or U5171 (N_5171,N_4490,N_4670);
and U5172 (N_5172,N_4582,N_4399);
nor U5173 (N_5173,N_4059,N_4891);
or U5174 (N_5174,N_4973,N_4730);
nand U5175 (N_5175,N_4489,N_4613);
nand U5176 (N_5176,N_4341,N_4005);
or U5177 (N_5177,N_4755,N_4198);
nand U5178 (N_5178,N_4472,N_4528);
or U5179 (N_5179,N_4745,N_4610);
nand U5180 (N_5180,N_4342,N_4880);
nand U5181 (N_5181,N_4836,N_4301);
and U5182 (N_5182,N_4025,N_4905);
nand U5183 (N_5183,N_4545,N_4547);
and U5184 (N_5184,N_4374,N_4599);
or U5185 (N_5185,N_4362,N_4426);
or U5186 (N_5186,N_4293,N_4534);
nor U5187 (N_5187,N_4121,N_4250);
nand U5188 (N_5188,N_4971,N_4800);
nor U5189 (N_5189,N_4927,N_4573);
and U5190 (N_5190,N_4754,N_4219);
or U5191 (N_5191,N_4779,N_4705);
or U5192 (N_5192,N_4997,N_4815);
nor U5193 (N_5193,N_4757,N_4211);
or U5194 (N_5194,N_4870,N_4348);
or U5195 (N_5195,N_4367,N_4739);
and U5196 (N_5196,N_4205,N_4737);
nor U5197 (N_5197,N_4575,N_4199);
nor U5198 (N_5198,N_4838,N_4857);
nand U5199 (N_5199,N_4869,N_4258);
and U5200 (N_5200,N_4920,N_4056);
or U5201 (N_5201,N_4470,N_4597);
nand U5202 (N_5202,N_4189,N_4663);
nand U5203 (N_5203,N_4942,N_4795);
or U5204 (N_5204,N_4580,N_4805);
or U5205 (N_5205,N_4461,N_4642);
nor U5206 (N_5206,N_4149,N_4637);
or U5207 (N_5207,N_4183,N_4949);
and U5208 (N_5208,N_4122,N_4749);
xnor U5209 (N_5209,N_4376,N_4925);
or U5210 (N_5210,N_4212,N_4050);
and U5211 (N_5211,N_4146,N_4161);
and U5212 (N_5212,N_4718,N_4331);
nand U5213 (N_5213,N_4751,N_4828);
and U5214 (N_5214,N_4366,N_4684);
nand U5215 (N_5215,N_4278,N_4087);
nor U5216 (N_5216,N_4909,N_4708);
nand U5217 (N_5217,N_4289,N_4526);
nand U5218 (N_5218,N_4983,N_4618);
nand U5219 (N_5219,N_4474,N_4141);
and U5220 (N_5220,N_4714,N_4834);
nor U5221 (N_5221,N_4203,N_4525);
and U5222 (N_5222,N_4977,N_4192);
and U5223 (N_5223,N_4179,N_4853);
nand U5224 (N_5224,N_4635,N_4306);
nor U5225 (N_5225,N_4621,N_4220);
and U5226 (N_5226,N_4349,N_4100);
and U5227 (N_5227,N_4529,N_4712);
nor U5228 (N_5228,N_4697,N_4119);
or U5229 (N_5229,N_4620,N_4940);
or U5230 (N_5230,N_4254,N_4410);
nand U5231 (N_5231,N_4798,N_4535);
nor U5232 (N_5232,N_4096,N_4091);
nand U5233 (N_5233,N_4554,N_4789);
or U5234 (N_5234,N_4009,N_4065);
nor U5235 (N_5235,N_4436,N_4105);
nand U5236 (N_5236,N_4987,N_4930);
nand U5237 (N_5237,N_4090,N_4540);
and U5238 (N_5238,N_4979,N_4455);
nor U5239 (N_5239,N_4412,N_4369);
xnor U5240 (N_5240,N_4874,N_4409);
nor U5241 (N_5241,N_4380,N_4171);
and U5242 (N_5242,N_4623,N_4980);
or U5243 (N_5243,N_4742,N_4257);
nor U5244 (N_5244,N_4990,N_4765);
or U5245 (N_5245,N_4771,N_4562);
nor U5246 (N_5246,N_4083,N_4358);
or U5247 (N_5247,N_4817,N_4080);
and U5248 (N_5248,N_4277,N_4845);
or U5249 (N_5249,N_4127,N_4735);
nand U5250 (N_5250,N_4947,N_4239);
or U5251 (N_5251,N_4416,N_4279);
and U5252 (N_5252,N_4488,N_4955);
nand U5253 (N_5253,N_4851,N_4893);
nand U5254 (N_5254,N_4162,N_4170);
and U5255 (N_5255,N_4201,N_4507);
and U5256 (N_5256,N_4709,N_4236);
and U5257 (N_5257,N_4876,N_4190);
and U5258 (N_5258,N_4695,N_4061);
nor U5259 (N_5259,N_4118,N_4064);
nand U5260 (N_5260,N_4493,N_4711);
and U5261 (N_5261,N_4896,N_4464);
or U5262 (N_5262,N_4391,N_4937);
and U5263 (N_5263,N_4605,N_4788);
and U5264 (N_5264,N_4068,N_4022);
nor U5265 (N_5265,N_4669,N_4646);
nor U5266 (N_5266,N_4686,N_4606);
nor U5267 (N_5267,N_4693,N_4224);
nor U5268 (N_5268,N_4338,N_4648);
and U5269 (N_5269,N_4588,N_4827);
nor U5270 (N_5270,N_4898,N_4862);
nor U5271 (N_5271,N_4858,N_4209);
and U5272 (N_5272,N_4133,N_4352);
nand U5273 (N_5273,N_4856,N_4350);
and U5274 (N_5274,N_4151,N_4633);
and U5275 (N_5275,N_4560,N_4191);
nand U5276 (N_5276,N_4473,N_4746);
and U5277 (N_5277,N_4498,N_4696);
nor U5278 (N_5278,N_4687,N_4095);
or U5279 (N_5279,N_4664,N_4451);
or U5280 (N_5280,N_4549,N_4469);
nor U5281 (N_5281,N_4809,N_4627);
and U5282 (N_5282,N_4672,N_4666);
and U5283 (N_5283,N_4335,N_4491);
and U5284 (N_5284,N_4938,N_4513);
and U5285 (N_5285,N_4082,N_4986);
or U5286 (N_5286,N_4832,N_4423);
and U5287 (N_5287,N_4678,N_4002);
nand U5288 (N_5288,N_4395,N_4569);
nand U5289 (N_5289,N_4629,N_4998);
or U5290 (N_5290,N_4587,N_4365);
nand U5291 (N_5291,N_4337,N_4288);
or U5292 (N_5292,N_4607,N_4622);
and U5293 (N_5293,N_4113,N_4843);
nand U5294 (N_5294,N_4126,N_4632);
and U5295 (N_5295,N_4086,N_4966);
nand U5296 (N_5296,N_4769,N_4996);
nor U5297 (N_5297,N_4178,N_4028);
or U5298 (N_5298,N_4519,N_4640);
and U5299 (N_5299,N_4504,N_4131);
nor U5300 (N_5300,N_4517,N_4654);
nor U5301 (N_5301,N_4165,N_4551);
nor U5302 (N_5302,N_4000,N_4900);
and U5303 (N_5303,N_4506,N_4109);
or U5304 (N_5304,N_4791,N_4019);
or U5305 (N_5305,N_4319,N_4450);
and U5306 (N_5306,N_4244,N_4916);
nor U5307 (N_5307,N_4184,N_4030);
nor U5308 (N_5308,N_4913,N_4773);
or U5309 (N_5309,N_4074,N_4683);
and U5310 (N_5310,N_4636,N_4922);
or U5311 (N_5311,N_4353,N_4057);
nor U5312 (N_5312,N_4381,N_4269);
and U5313 (N_5313,N_4238,N_4999);
or U5314 (N_5314,N_4085,N_4772);
nor U5315 (N_5315,N_4351,N_4767);
nor U5316 (N_5316,N_4142,N_4803);
or U5317 (N_5317,N_4232,N_4271);
nor U5318 (N_5318,N_4667,N_4612);
nor U5319 (N_5319,N_4333,N_4446);
or U5320 (N_5320,N_4072,N_4125);
xor U5321 (N_5321,N_4725,N_4103);
or U5322 (N_5322,N_4392,N_4890);
nand U5323 (N_5323,N_4732,N_4766);
nand U5324 (N_5324,N_4954,N_4425);
nand U5325 (N_5325,N_4593,N_4387);
nand U5326 (N_5326,N_4566,N_4565);
nor U5327 (N_5327,N_4385,N_4720);
and U5328 (N_5328,N_4375,N_4242);
and U5329 (N_5329,N_4077,N_4427);
and U5330 (N_5330,N_4885,N_4214);
nand U5331 (N_5331,N_4194,N_4263);
nor U5332 (N_5332,N_4483,N_4213);
xnor U5333 (N_5333,N_4134,N_4459);
or U5334 (N_5334,N_4340,N_4796);
or U5335 (N_5335,N_4063,N_4274);
and U5336 (N_5336,N_4797,N_4093);
nor U5337 (N_5337,N_4041,N_4334);
or U5338 (N_5338,N_4558,N_4744);
and U5339 (N_5339,N_4522,N_4255);
nor U5340 (N_5340,N_4320,N_4631);
nand U5341 (N_5341,N_4414,N_4864);
nor U5342 (N_5342,N_4112,N_4625);
or U5343 (N_5343,N_4908,N_4665);
and U5344 (N_5344,N_4946,N_4249);
nand U5345 (N_5345,N_4733,N_4047);
nand U5346 (N_5346,N_4811,N_4463);
and U5347 (N_5347,N_4413,N_4296);
nand U5348 (N_5348,N_4229,N_4701);
nand U5349 (N_5349,N_4933,N_4509);
nand U5350 (N_5350,N_4563,N_4328);
nor U5351 (N_5351,N_4321,N_4431);
and U5352 (N_5352,N_4941,N_4111);
and U5353 (N_5353,N_4595,N_4521);
or U5354 (N_5354,N_4871,N_4314);
nor U5355 (N_5355,N_4477,N_4967);
and U5356 (N_5356,N_4223,N_4956);
nor U5357 (N_5357,N_4884,N_4479);
and U5358 (N_5358,N_4993,N_4260);
or U5359 (N_5359,N_4152,N_4760);
nand U5360 (N_5360,N_4914,N_4013);
or U5361 (N_5361,N_4747,N_4794);
or U5362 (N_5362,N_4107,N_4485);
nand U5363 (N_5363,N_4888,N_4039);
and U5364 (N_5364,N_4758,N_4453);
and U5365 (N_5365,N_4176,N_4014);
and U5366 (N_5366,N_4497,N_4417);
nand U5367 (N_5367,N_4777,N_4386);
nand U5368 (N_5368,N_4786,N_4576);
and U5369 (N_5369,N_4500,N_4752);
or U5370 (N_5370,N_4308,N_4067);
and U5371 (N_5371,N_4824,N_4405);
nor U5372 (N_5372,N_4731,N_4935);
and U5373 (N_5373,N_4963,N_4206);
or U5374 (N_5374,N_4428,N_4835);
or U5375 (N_5375,N_4761,N_4812);
nor U5376 (N_5376,N_4784,N_4770);
nor U5377 (N_5377,N_4740,N_4139);
and U5378 (N_5378,N_4846,N_4523);
and U5379 (N_5379,N_4516,N_4662);
nor U5380 (N_5380,N_4355,N_4264);
nor U5381 (N_5381,N_4813,N_4177);
nand U5382 (N_5382,N_4647,N_4422);
nand U5383 (N_5383,N_4926,N_4015);
xor U5384 (N_5384,N_4975,N_4550);
or U5385 (N_5385,N_4207,N_4912);
nand U5386 (N_5386,N_4792,N_4377);
xor U5387 (N_5387,N_4682,N_4936);
and U5388 (N_5388,N_4322,N_4514);
nand U5389 (N_5389,N_4372,N_4600);
nand U5390 (N_5390,N_4415,N_4038);
nor U5391 (N_5391,N_4434,N_4844);
and U5392 (N_5392,N_4903,N_4444);
nor U5393 (N_5393,N_4833,N_4196);
nand U5394 (N_5394,N_4197,N_4974);
and U5395 (N_5395,N_4879,N_4275);
or U5396 (N_5396,N_4029,N_4503);
or U5397 (N_5397,N_4031,N_4572);
or U5398 (N_5398,N_4810,N_4267);
nor U5399 (N_5399,N_4402,N_4964);
nand U5400 (N_5400,N_4704,N_4383);
and U5401 (N_5401,N_4611,N_4872);
nor U5402 (N_5402,N_4546,N_4753);
nand U5403 (N_5403,N_4040,N_4866);
nand U5404 (N_5404,N_4262,N_4442);
nand U5405 (N_5405,N_4175,N_4875);
or U5406 (N_5406,N_4502,N_4628);
nand U5407 (N_5407,N_4329,N_4160);
nor U5408 (N_5408,N_4435,N_4092);
and U5409 (N_5409,N_4616,N_4944);
nand U5410 (N_5410,N_4603,N_4602);
or U5411 (N_5411,N_4297,N_4799);
nand U5412 (N_5412,N_4008,N_4237);
or U5413 (N_5413,N_4486,N_4032);
and U5414 (N_5414,N_4657,N_4027);
or U5415 (N_5415,N_4583,N_4246);
or U5416 (N_5416,N_4292,N_4959);
nand U5417 (N_5417,N_4218,N_4923);
and U5418 (N_5418,N_4991,N_4217);
nand U5419 (N_5419,N_4202,N_4361);
or U5420 (N_5420,N_4807,N_4406);
or U5421 (N_5421,N_4454,N_4653);
and U5422 (N_5422,N_4079,N_4907);
and U5423 (N_5423,N_4764,N_4848);
and U5424 (N_5424,N_4982,N_4830);
nand U5425 (N_5425,N_4911,N_4586);
and U5426 (N_5426,N_4418,N_4918);
and U5427 (N_5427,N_4396,N_4153);
nor U5428 (N_5428,N_4638,N_4465);
or U5429 (N_5429,N_4829,N_4592);
nand U5430 (N_5430,N_4373,N_4873);
and U5431 (N_5431,N_4533,N_4617);
or U5432 (N_5432,N_4688,N_4276);
and U5433 (N_5433,N_4520,N_4734);
or U5434 (N_5434,N_4527,N_4537);
and U5435 (N_5435,N_4702,N_4364);
nor U5436 (N_5436,N_4715,N_4690);
and U5437 (N_5437,N_4776,N_4988);
or U5438 (N_5438,N_4115,N_4044);
and U5439 (N_5439,N_4379,N_4619);
and U5440 (N_5440,N_4174,N_4440);
nor U5441 (N_5441,N_4630,N_4054);
xnor U5442 (N_5442,N_4078,N_4494);
and U5443 (N_5443,N_4819,N_4004);
and U5444 (N_5444,N_4826,N_4110);
nor U5445 (N_5445,N_4726,N_4894);
nor U5446 (N_5446,N_4286,N_4481);
or U5447 (N_5447,N_4861,N_4339);
or U5448 (N_5448,N_4536,N_4053);
or U5449 (N_5449,N_4020,N_4877);
nand U5450 (N_5450,N_4155,N_4101);
nand U5451 (N_5451,N_4604,N_4438);
nand U5452 (N_5452,N_4915,N_4081);
nor U5453 (N_5453,N_4738,N_4660);
nor U5454 (N_5454,N_4743,N_4951);
and U5455 (N_5455,N_4159,N_4317);
or U5456 (N_5456,N_4721,N_4928);
and U5457 (N_5457,N_4123,N_4651);
nand U5458 (N_5458,N_4195,N_4539);
or U5459 (N_5459,N_4659,N_4104);
and U5460 (N_5460,N_4840,N_4487);
nor U5461 (N_5461,N_4408,N_4302);
or U5462 (N_5462,N_4859,N_4084);
and U5463 (N_5463,N_4511,N_4816);
nand U5464 (N_5464,N_4215,N_4793);
and U5465 (N_5465,N_4124,N_4295);
or U5466 (N_5466,N_4713,N_4147);
nor U5467 (N_5467,N_4368,N_4808);
nand U5468 (N_5468,N_4305,N_4860);
xnor U5469 (N_5469,N_4037,N_4354);
and U5470 (N_5470,N_4655,N_4865);
nand U5471 (N_5471,N_4448,N_4248);
nor U5472 (N_5472,N_4011,N_4729);
and U5473 (N_5473,N_4186,N_4390);
nor U5474 (N_5474,N_4984,N_4231);
nor U5475 (N_5475,N_4116,N_4962);
nor U5476 (N_5476,N_4518,N_4707);
and U5477 (N_5477,N_4138,N_4530);
and U5478 (N_5478,N_4210,N_4135);
nor U5479 (N_5479,N_4598,N_4221);
nand U5480 (N_5480,N_4046,N_4094);
and U5481 (N_5481,N_4863,N_4290);
nand U5482 (N_5482,N_4247,N_4265);
nor U5483 (N_5483,N_4154,N_4346);
and U5484 (N_5484,N_4806,N_4312);
nand U5485 (N_5485,N_4932,N_4252);
nand U5486 (N_5486,N_4649,N_4906);
or U5487 (N_5487,N_4867,N_4581);
nor U5488 (N_5488,N_4945,N_4692);
nand U5489 (N_5489,N_4783,N_4589);
or U5490 (N_5490,N_4965,N_4345);
and U5491 (N_5491,N_4495,N_4439);
and U5492 (N_5492,N_4694,N_4261);
nor U5493 (N_5493,N_4180,N_4468);
nor U5494 (N_5494,N_4188,N_4360);
and U5495 (N_5495,N_4839,N_4567);
nand U5496 (N_5496,N_4496,N_4480);
nand U5497 (N_5497,N_4256,N_4822);
nor U5498 (N_5498,N_4952,N_4316);
nand U5499 (N_5499,N_4150,N_4557);
xor U5500 (N_5500,N_4901,N_4480);
and U5501 (N_5501,N_4191,N_4146);
or U5502 (N_5502,N_4640,N_4714);
nor U5503 (N_5503,N_4868,N_4618);
nor U5504 (N_5504,N_4659,N_4358);
nand U5505 (N_5505,N_4406,N_4139);
and U5506 (N_5506,N_4704,N_4443);
or U5507 (N_5507,N_4403,N_4728);
nand U5508 (N_5508,N_4468,N_4695);
or U5509 (N_5509,N_4274,N_4580);
nor U5510 (N_5510,N_4652,N_4584);
nor U5511 (N_5511,N_4210,N_4829);
nand U5512 (N_5512,N_4835,N_4920);
nand U5513 (N_5513,N_4627,N_4741);
nor U5514 (N_5514,N_4917,N_4300);
or U5515 (N_5515,N_4899,N_4035);
nand U5516 (N_5516,N_4929,N_4167);
or U5517 (N_5517,N_4051,N_4696);
or U5518 (N_5518,N_4729,N_4067);
nor U5519 (N_5519,N_4389,N_4805);
nor U5520 (N_5520,N_4967,N_4953);
nor U5521 (N_5521,N_4440,N_4979);
or U5522 (N_5522,N_4730,N_4595);
and U5523 (N_5523,N_4884,N_4074);
nand U5524 (N_5524,N_4299,N_4527);
nand U5525 (N_5525,N_4562,N_4668);
nor U5526 (N_5526,N_4296,N_4300);
nor U5527 (N_5527,N_4699,N_4050);
or U5528 (N_5528,N_4083,N_4459);
nand U5529 (N_5529,N_4539,N_4674);
xor U5530 (N_5530,N_4520,N_4262);
nor U5531 (N_5531,N_4860,N_4617);
nand U5532 (N_5532,N_4059,N_4262);
nor U5533 (N_5533,N_4837,N_4492);
nor U5534 (N_5534,N_4376,N_4080);
and U5535 (N_5535,N_4148,N_4632);
and U5536 (N_5536,N_4099,N_4178);
nand U5537 (N_5537,N_4941,N_4680);
or U5538 (N_5538,N_4616,N_4461);
nand U5539 (N_5539,N_4754,N_4813);
xnor U5540 (N_5540,N_4716,N_4237);
or U5541 (N_5541,N_4007,N_4056);
nor U5542 (N_5542,N_4559,N_4579);
nand U5543 (N_5543,N_4166,N_4826);
and U5544 (N_5544,N_4970,N_4014);
or U5545 (N_5545,N_4608,N_4711);
nor U5546 (N_5546,N_4149,N_4456);
or U5547 (N_5547,N_4285,N_4153);
or U5548 (N_5548,N_4552,N_4125);
or U5549 (N_5549,N_4918,N_4826);
nor U5550 (N_5550,N_4726,N_4651);
and U5551 (N_5551,N_4748,N_4758);
nor U5552 (N_5552,N_4984,N_4126);
and U5553 (N_5553,N_4294,N_4243);
or U5554 (N_5554,N_4475,N_4158);
nand U5555 (N_5555,N_4016,N_4854);
and U5556 (N_5556,N_4136,N_4362);
and U5557 (N_5557,N_4298,N_4245);
nand U5558 (N_5558,N_4343,N_4048);
and U5559 (N_5559,N_4673,N_4133);
and U5560 (N_5560,N_4983,N_4534);
and U5561 (N_5561,N_4332,N_4315);
and U5562 (N_5562,N_4803,N_4405);
nor U5563 (N_5563,N_4236,N_4925);
or U5564 (N_5564,N_4569,N_4845);
nor U5565 (N_5565,N_4746,N_4968);
nor U5566 (N_5566,N_4312,N_4066);
and U5567 (N_5567,N_4276,N_4375);
nor U5568 (N_5568,N_4590,N_4985);
nand U5569 (N_5569,N_4930,N_4707);
nand U5570 (N_5570,N_4409,N_4276);
and U5571 (N_5571,N_4839,N_4691);
nand U5572 (N_5572,N_4624,N_4603);
nor U5573 (N_5573,N_4030,N_4527);
nand U5574 (N_5574,N_4724,N_4389);
or U5575 (N_5575,N_4052,N_4138);
nor U5576 (N_5576,N_4164,N_4027);
nor U5577 (N_5577,N_4264,N_4804);
and U5578 (N_5578,N_4732,N_4857);
xor U5579 (N_5579,N_4578,N_4775);
and U5580 (N_5580,N_4113,N_4141);
nand U5581 (N_5581,N_4524,N_4678);
nand U5582 (N_5582,N_4551,N_4756);
nor U5583 (N_5583,N_4566,N_4221);
nand U5584 (N_5584,N_4051,N_4980);
nand U5585 (N_5585,N_4779,N_4616);
or U5586 (N_5586,N_4331,N_4736);
nor U5587 (N_5587,N_4490,N_4778);
nor U5588 (N_5588,N_4620,N_4928);
nor U5589 (N_5589,N_4062,N_4972);
nand U5590 (N_5590,N_4274,N_4640);
nor U5591 (N_5591,N_4137,N_4980);
nand U5592 (N_5592,N_4866,N_4737);
and U5593 (N_5593,N_4503,N_4518);
nor U5594 (N_5594,N_4598,N_4111);
nor U5595 (N_5595,N_4760,N_4344);
nor U5596 (N_5596,N_4430,N_4696);
nor U5597 (N_5597,N_4830,N_4675);
and U5598 (N_5598,N_4937,N_4306);
nor U5599 (N_5599,N_4867,N_4156);
or U5600 (N_5600,N_4906,N_4749);
nor U5601 (N_5601,N_4382,N_4442);
and U5602 (N_5602,N_4218,N_4325);
or U5603 (N_5603,N_4468,N_4136);
or U5604 (N_5604,N_4580,N_4160);
xnor U5605 (N_5605,N_4885,N_4524);
and U5606 (N_5606,N_4224,N_4036);
nand U5607 (N_5607,N_4672,N_4559);
or U5608 (N_5608,N_4337,N_4943);
nor U5609 (N_5609,N_4862,N_4899);
and U5610 (N_5610,N_4247,N_4916);
nand U5611 (N_5611,N_4274,N_4880);
nor U5612 (N_5612,N_4732,N_4576);
or U5613 (N_5613,N_4113,N_4571);
and U5614 (N_5614,N_4922,N_4685);
nand U5615 (N_5615,N_4350,N_4656);
nand U5616 (N_5616,N_4625,N_4278);
nor U5617 (N_5617,N_4611,N_4411);
or U5618 (N_5618,N_4709,N_4035);
or U5619 (N_5619,N_4222,N_4873);
nor U5620 (N_5620,N_4062,N_4891);
or U5621 (N_5621,N_4341,N_4112);
and U5622 (N_5622,N_4988,N_4163);
nor U5623 (N_5623,N_4038,N_4570);
xnor U5624 (N_5624,N_4029,N_4232);
or U5625 (N_5625,N_4316,N_4442);
and U5626 (N_5626,N_4863,N_4746);
nand U5627 (N_5627,N_4507,N_4827);
or U5628 (N_5628,N_4693,N_4763);
and U5629 (N_5629,N_4086,N_4996);
nor U5630 (N_5630,N_4493,N_4917);
or U5631 (N_5631,N_4994,N_4903);
nand U5632 (N_5632,N_4359,N_4858);
and U5633 (N_5633,N_4506,N_4487);
or U5634 (N_5634,N_4298,N_4334);
nand U5635 (N_5635,N_4718,N_4036);
nor U5636 (N_5636,N_4320,N_4959);
and U5637 (N_5637,N_4736,N_4735);
nand U5638 (N_5638,N_4098,N_4837);
or U5639 (N_5639,N_4151,N_4923);
and U5640 (N_5640,N_4737,N_4919);
or U5641 (N_5641,N_4141,N_4625);
nand U5642 (N_5642,N_4133,N_4954);
or U5643 (N_5643,N_4680,N_4035);
or U5644 (N_5644,N_4517,N_4667);
and U5645 (N_5645,N_4028,N_4814);
nand U5646 (N_5646,N_4352,N_4402);
nand U5647 (N_5647,N_4201,N_4506);
nand U5648 (N_5648,N_4866,N_4137);
or U5649 (N_5649,N_4575,N_4139);
nor U5650 (N_5650,N_4261,N_4247);
nor U5651 (N_5651,N_4297,N_4501);
or U5652 (N_5652,N_4834,N_4183);
nand U5653 (N_5653,N_4629,N_4570);
nor U5654 (N_5654,N_4965,N_4422);
or U5655 (N_5655,N_4956,N_4754);
nand U5656 (N_5656,N_4936,N_4090);
and U5657 (N_5657,N_4103,N_4192);
or U5658 (N_5658,N_4653,N_4460);
nor U5659 (N_5659,N_4102,N_4445);
nor U5660 (N_5660,N_4018,N_4889);
nand U5661 (N_5661,N_4193,N_4757);
and U5662 (N_5662,N_4910,N_4159);
nand U5663 (N_5663,N_4372,N_4783);
nand U5664 (N_5664,N_4094,N_4760);
and U5665 (N_5665,N_4051,N_4393);
nand U5666 (N_5666,N_4842,N_4408);
or U5667 (N_5667,N_4610,N_4526);
or U5668 (N_5668,N_4280,N_4579);
nor U5669 (N_5669,N_4135,N_4741);
and U5670 (N_5670,N_4916,N_4989);
or U5671 (N_5671,N_4267,N_4991);
nand U5672 (N_5672,N_4641,N_4245);
and U5673 (N_5673,N_4691,N_4936);
and U5674 (N_5674,N_4359,N_4505);
nand U5675 (N_5675,N_4442,N_4735);
nand U5676 (N_5676,N_4172,N_4353);
and U5677 (N_5677,N_4643,N_4688);
nor U5678 (N_5678,N_4250,N_4216);
or U5679 (N_5679,N_4084,N_4396);
and U5680 (N_5680,N_4592,N_4053);
and U5681 (N_5681,N_4831,N_4476);
and U5682 (N_5682,N_4914,N_4265);
nor U5683 (N_5683,N_4937,N_4707);
or U5684 (N_5684,N_4672,N_4532);
nor U5685 (N_5685,N_4201,N_4569);
and U5686 (N_5686,N_4041,N_4074);
nand U5687 (N_5687,N_4710,N_4125);
and U5688 (N_5688,N_4189,N_4071);
nand U5689 (N_5689,N_4815,N_4638);
or U5690 (N_5690,N_4080,N_4722);
or U5691 (N_5691,N_4315,N_4258);
or U5692 (N_5692,N_4319,N_4388);
or U5693 (N_5693,N_4311,N_4095);
nor U5694 (N_5694,N_4041,N_4594);
or U5695 (N_5695,N_4641,N_4982);
or U5696 (N_5696,N_4064,N_4032);
nor U5697 (N_5697,N_4852,N_4683);
nor U5698 (N_5698,N_4693,N_4564);
nand U5699 (N_5699,N_4922,N_4073);
nand U5700 (N_5700,N_4814,N_4791);
nor U5701 (N_5701,N_4448,N_4886);
nand U5702 (N_5702,N_4126,N_4070);
and U5703 (N_5703,N_4892,N_4229);
or U5704 (N_5704,N_4531,N_4772);
and U5705 (N_5705,N_4654,N_4878);
nor U5706 (N_5706,N_4831,N_4300);
or U5707 (N_5707,N_4376,N_4817);
nor U5708 (N_5708,N_4101,N_4160);
and U5709 (N_5709,N_4815,N_4385);
and U5710 (N_5710,N_4666,N_4547);
and U5711 (N_5711,N_4351,N_4150);
and U5712 (N_5712,N_4540,N_4408);
nand U5713 (N_5713,N_4275,N_4246);
or U5714 (N_5714,N_4574,N_4758);
nand U5715 (N_5715,N_4300,N_4534);
nor U5716 (N_5716,N_4642,N_4601);
or U5717 (N_5717,N_4439,N_4840);
and U5718 (N_5718,N_4674,N_4534);
nand U5719 (N_5719,N_4220,N_4419);
or U5720 (N_5720,N_4899,N_4083);
nor U5721 (N_5721,N_4335,N_4237);
nor U5722 (N_5722,N_4676,N_4455);
nor U5723 (N_5723,N_4913,N_4600);
or U5724 (N_5724,N_4153,N_4360);
nand U5725 (N_5725,N_4714,N_4590);
or U5726 (N_5726,N_4587,N_4546);
nand U5727 (N_5727,N_4642,N_4790);
nand U5728 (N_5728,N_4388,N_4569);
or U5729 (N_5729,N_4362,N_4245);
or U5730 (N_5730,N_4029,N_4977);
nand U5731 (N_5731,N_4678,N_4299);
nand U5732 (N_5732,N_4706,N_4803);
nor U5733 (N_5733,N_4494,N_4418);
nor U5734 (N_5734,N_4788,N_4621);
and U5735 (N_5735,N_4054,N_4375);
or U5736 (N_5736,N_4092,N_4106);
nand U5737 (N_5737,N_4904,N_4515);
or U5738 (N_5738,N_4434,N_4815);
or U5739 (N_5739,N_4163,N_4766);
nor U5740 (N_5740,N_4018,N_4305);
and U5741 (N_5741,N_4714,N_4049);
nor U5742 (N_5742,N_4340,N_4196);
xnor U5743 (N_5743,N_4633,N_4335);
nand U5744 (N_5744,N_4360,N_4620);
nor U5745 (N_5745,N_4343,N_4667);
nor U5746 (N_5746,N_4592,N_4909);
nor U5747 (N_5747,N_4705,N_4038);
nand U5748 (N_5748,N_4758,N_4784);
nand U5749 (N_5749,N_4286,N_4355);
or U5750 (N_5750,N_4768,N_4783);
or U5751 (N_5751,N_4913,N_4696);
and U5752 (N_5752,N_4575,N_4386);
or U5753 (N_5753,N_4985,N_4936);
and U5754 (N_5754,N_4802,N_4741);
or U5755 (N_5755,N_4588,N_4644);
nand U5756 (N_5756,N_4056,N_4821);
or U5757 (N_5757,N_4214,N_4333);
nor U5758 (N_5758,N_4090,N_4174);
nor U5759 (N_5759,N_4549,N_4867);
or U5760 (N_5760,N_4385,N_4399);
or U5761 (N_5761,N_4007,N_4495);
nand U5762 (N_5762,N_4418,N_4157);
and U5763 (N_5763,N_4533,N_4941);
nand U5764 (N_5764,N_4011,N_4638);
nand U5765 (N_5765,N_4593,N_4821);
and U5766 (N_5766,N_4534,N_4550);
and U5767 (N_5767,N_4844,N_4030);
nand U5768 (N_5768,N_4891,N_4587);
nand U5769 (N_5769,N_4148,N_4468);
and U5770 (N_5770,N_4303,N_4998);
nand U5771 (N_5771,N_4790,N_4510);
or U5772 (N_5772,N_4247,N_4692);
nand U5773 (N_5773,N_4008,N_4932);
and U5774 (N_5774,N_4726,N_4456);
nand U5775 (N_5775,N_4120,N_4765);
nor U5776 (N_5776,N_4508,N_4474);
or U5777 (N_5777,N_4239,N_4116);
nand U5778 (N_5778,N_4232,N_4717);
or U5779 (N_5779,N_4308,N_4694);
nor U5780 (N_5780,N_4363,N_4310);
nor U5781 (N_5781,N_4036,N_4473);
and U5782 (N_5782,N_4306,N_4010);
nand U5783 (N_5783,N_4070,N_4844);
or U5784 (N_5784,N_4969,N_4481);
and U5785 (N_5785,N_4667,N_4148);
nand U5786 (N_5786,N_4025,N_4116);
or U5787 (N_5787,N_4791,N_4469);
or U5788 (N_5788,N_4524,N_4529);
xor U5789 (N_5789,N_4854,N_4334);
nand U5790 (N_5790,N_4811,N_4256);
nand U5791 (N_5791,N_4979,N_4735);
nor U5792 (N_5792,N_4147,N_4143);
xor U5793 (N_5793,N_4771,N_4442);
nand U5794 (N_5794,N_4187,N_4156);
nor U5795 (N_5795,N_4813,N_4172);
or U5796 (N_5796,N_4231,N_4695);
and U5797 (N_5797,N_4851,N_4983);
or U5798 (N_5798,N_4558,N_4119);
nor U5799 (N_5799,N_4943,N_4603);
nand U5800 (N_5800,N_4069,N_4802);
or U5801 (N_5801,N_4446,N_4707);
and U5802 (N_5802,N_4621,N_4038);
nor U5803 (N_5803,N_4676,N_4649);
or U5804 (N_5804,N_4787,N_4561);
nand U5805 (N_5805,N_4369,N_4049);
or U5806 (N_5806,N_4394,N_4697);
and U5807 (N_5807,N_4073,N_4509);
or U5808 (N_5808,N_4662,N_4473);
nand U5809 (N_5809,N_4301,N_4244);
or U5810 (N_5810,N_4857,N_4201);
nand U5811 (N_5811,N_4552,N_4314);
or U5812 (N_5812,N_4064,N_4294);
or U5813 (N_5813,N_4062,N_4222);
and U5814 (N_5814,N_4902,N_4419);
nand U5815 (N_5815,N_4723,N_4901);
xnor U5816 (N_5816,N_4488,N_4223);
nand U5817 (N_5817,N_4792,N_4123);
and U5818 (N_5818,N_4951,N_4573);
nand U5819 (N_5819,N_4884,N_4468);
or U5820 (N_5820,N_4683,N_4169);
or U5821 (N_5821,N_4523,N_4500);
xnor U5822 (N_5822,N_4305,N_4837);
nand U5823 (N_5823,N_4807,N_4410);
nor U5824 (N_5824,N_4431,N_4856);
nor U5825 (N_5825,N_4068,N_4650);
nor U5826 (N_5826,N_4646,N_4772);
nand U5827 (N_5827,N_4824,N_4221);
and U5828 (N_5828,N_4522,N_4831);
and U5829 (N_5829,N_4474,N_4930);
and U5830 (N_5830,N_4780,N_4637);
or U5831 (N_5831,N_4371,N_4030);
nand U5832 (N_5832,N_4186,N_4279);
and U5833 (N_5833,N_4541,N_4850);
nor U5834 (N_5834,N_4538,N_4176);
nor U5835 (N_5835,N_4665,N_4308);
nand U5836 (N_5836,N_4364,N_4395);
nand U5837 (N_5837,N_4694,N_4304);
nand U5838 (N_5838,N_4817,N_4652);
and U5839 (N_5839,N_4669,N_4753);
nand U5840 (N_5840,N_4950,N_4785);
nand U5841 (N_5841,N_4518,N_4482);
nor U5842 (N_5842,N_4622,N_4832);
and U5843 (N_5843,N_4643,N_4832);
nor U5844 (N_5844,N_4261,N_4695);
and U5845 (N_5845,N_4431,N_4749);
nor U5846 (N_5846,N_4906,N_4502);
nand U5847 (N_5847,N_4426,N_4584);
nand U5848 (N_5848,N_4481,N_4525);
nand U5849 (N_5849,N_4531,N_4896);
and U5850 (N_5850,N_4354,N_4568);
or U5851 (N_5851,N_4716,N_4828);
or U5852 (N_5852,N_4034,N_4347);
and U5853 (N_5853,N_4973,N_4285);
and U5854 (N_5854,N_4352,N_4157);
nand U5855 (N_5855,N_4876,N_4309);
and U5856 (N_5856,N_4558,N_4435);
and U5857 (N_5857,N_4710,N_4959);
nor U5858 (N_5858,N_4175,N_4852);
nand U5859 (N_5859,N_4640,N_4172);
nor U5860 (N_5860,N_4310,N_4340);
and U5861 (N_5861,N_4758,N_4556);
or U5862 (N_5862,N_4227,N_4308);
nor U5863 (N_5863,N_4577,N_4536);
nand U5864 (N_5864,N_4283,N_4301);
or U5865 (N_5865,N_4094,N_4721);
or U5866 (N_5866,N_4997,N_4214);
nor U5867 (N_5867,N_4687,N_4602);
nand U5868 (N_5868,N_4376,N_4005);
xnor U5869 (N_5869,N_4425,N_4765);
nor U5870 (N_5870,N_4170,N_4415);
and U5871 (N_5871,N_4889,N_4377);
or U5872 (N_5872,N_4879,N_4098);
and U5873 (N_5873,N_4040,N_4348);
and U5874 (N_5874,N_4851,N_4949);
nor U5875 (N_5875,N_4284,N_4117);
nor U5876 (N_5876,N_4677,N_4355);
nor U5877 (N_5877,N_4276,N_4471);
or U5878 (N_5878,N_4337,N_4779);
or U5879 (N_5879,N_4315,N_4502);
or U5880 (N_5880,N_4825,N_4701);
nand U5881 (N_5881,N_4969,N_4344);
and U5882 (N_5882,N_4149,N_4889);
or U5883 (N_5883,N_4470,N_4931);
nand U5884 (N_5884,N_4489,N_4576);
nor U5885 (N_5885,N_4483,N_4460);
or U5886 (N_5886,N_4672,N_4669);
nor U5887 (N_5887,N_4572,N_4782);
nand U5888 (N_5888,N_4290,N_4566);
or U5889 (N_5889,N_4576,N_4376);
or U5890 (N_5890,N_4931,N_4494);
nor U5891 (N_5891,N_4353,N_4708);
or U5892 (N_5892,N_4136,N_4306);
nand U5893 (N_5893,N_4745,N_4856);
nor U5894 (N_5894,N_4527,N_4246);
and U5895 (N_5895,N_4116,N_4104);
or U5896 (N_5896,N_4078,N_4828);
nand U5897 (N_5897,N_4700,N_4025);
and U5898 (N_5898,N_4381,N_4737);
nor U5899 (N_5899,N_4762,N_4993);
or U5900 (N_5900,N_4862,N_4471);
or U5901 (N_5901,N_4224,N_4144);
or U5902 (N_5902,N_4322,N_4618);
and U5903 (N_5903,N_4956,N_4456);
nor U5904 (N_5904,N_4608,N_4538);
nor U5905 (N_5905,N_4667,N_4609);
and U5906 (N_5906,N_4137,N_4334);
or U5907 (N_5907,N_4432,N_4417);
nor U5908 (N_5908,N_4026,N_4950);
and U5909 (N_5909,N_4364,N_4959);
and U5910 (N_5910,N_4171,N_4911);
and U5911 (N_5911,N_4026,N_4429);
nand U5912 (N_5912,N_4459,N_4213);
xnor U5913 (N_5913,N_4020,N_4421);
nand U5914 (N_5914,N_4259,N_4384);
and U5915 (N_5915,N_4558,N_4539);
or U5916 (N_5916,N_4339,N_4318);
nor U5917 (N_5917,N_4832,N_4193);
and U5918 (N_5918,N_4630,N_4873);
or U5919 (N_5919,N_4180,N_4595);
or U5920 (N_5920,N_4233,N_4416);
xor U5921 (N_5921,N_4057,N_4088);
or U5922 (N_5922,N_4367,N_4348);
xnor U5923 (N_5923,N_4860,N_4687);
or U5924 (N_5924,N_4882,N_4626);
nand U5925 (N_5925,N_4010,N_4063);
and U5926 (N_5926,N_4872,N_4049);
or U5927 (N_5927,N_4478,N_4085);
nor U5928 (N_5928,N_4538,N_4190);
xnor U5929 (N_5929,N_4457,N_4256);
or U5930 (N_5930,N_4970,N_4261);
nand U5931 (N_5931,N_4154,N_4253);
nand U5932 (N_5932,N_4585,N_4963);
xnor U5933 (N_5933,N_4570,N_4318);
nand U5934 (N_5934,N_4121,N_4463);
nand U5935 (N_5935,N_4983,N_4861);
nand U5936 (N_5936,N_4022,N_4581);
nand U5937 (N_5937,N_4045,N_4136);
or U5938 (N_5938,N_4856,N_4825);
and U5939 (N_5939,N_4990,N_4714);
and U5940 (N_5940,N_4524,N_4086);
and U5941 (N_5941,N_4404,N_4613);
xnor U5942 (N_5942,N_4236,N_4266);
xnor U5943 (N_5943,N_4735,N_4530);
and U5944 (N_5944,N_4291,N_4112);
nor U5945 (N_5945,N_4601,N_4207);
or U5946 (N_5946,N_4050,N_4783);
nand U5947 (N_5947,N_4092,N_4469);
and U5948 (N_5948,N_4222,N_4934);
nor U5949 (N_5949,N_4790,N_4529);
or U5950 (N_5950,N_4285,N_4289);
or U5951 (N_5951,N_4881,N_4645);
or U5952 (N_5952,N_4371,N_4456);
xnor U5953 (N_5953,N_4449,N_4886);
and U5954 (N_5954,N_4985,N_4212);
nand U5955 (N_5955,N_4047,N_4598);
nor U5956 (N_5956,N_4003,N_4529);
and U5957 (N_5957,N_4319,N_4587);
and U5958 (N_5958,N_4858,N_4256);
and U5959 (N_5959,N_4619,N_4877);
and U5960 (N_5960,N_4240,N_4573);
nand U5961 (N_5961,N_4459,N_4365);
or U5962 (N_5962,N_4790,N_4660);
nor U5963 (N_5963,N_4493,N_4167);
xnor U5964 (N_5964,N_4661,N_4022);
nand U5965 (N_5965,N_4734,N_4286);
and U5966 (N_5966,N_4166,N_4832);
and U5967 (N_5967,N_4098,N_4321);
or U5968 (N_5968,N_4737,N_4877);
and U5969 (N_5969,N_4226,N_4068);
nand U5970 (N_5970,N_4780,N_4460);
nor U5971 (N_5971,N_4739,N_4654);
and U5972 (N_5972,N_4299,N_4699);
or U5973 (N_5973,N_4733,N_4712);
or U5974 (N_5974,N_4009,N_4005);
and U5975 (N_5975,N_4806,N_4371);
nor U5976 (N_5976,N_4214,N_4614);
or U5977 (N_5977,N_4951,N_4983);
or U5978 (N_5978,N_4532,N_4029);
and U5979 (N_5979,N_4270,N_4309);
nor U5980 (N_5980,N_4045,N_4633);
nand U5981 (N_5981,N_4337,N_4875);
nand U5982 (N_5982,N_4469,N_4675);
or U5983 (N_5983,N_4110,N_4738);
nor U5984 (N_5984,N_4363,N_4889);
or U5985 (N_5985,N_4385,N_4537);
and U5986 (N_5986,N_4281,N_4902);
or U5987 (N_5987,N_4792,N_4810);
nand U5988 (N_5988,N_4251,N_4628);
nand U5989 (N_5989,N_4883,N_4271);
or U5990 (N_5990,N_4889,N_4678);
and U5991 (N_5991,N_4826,N_4211);
nor U5992 (N_5992,N_4574,N_4625);
and U5993 (N_5993,N_4350,N_4137);
or U5994 (N_5994,N_4115,N_4484);
or U5995 (N_5995,N_4905,N_4249);
nand U5996 (N_5996,N_4222,N_4890);
or U5997 (N_5997,N_4149,N_4023);
or U5998 (N_5998,N_4592,N_4226);
or U5999 (N_5999,N_4463,N_4748);
or U6000 (N_6000,N_5851,N_5046);
or U6001 (N_6001,N_5711,N_5824);
and U6002 (N_6002,N_5133,N_5609);
and U6003 (N_6003,N_5799,N_5550);
nand U6004 (N_6004,N_5930,N_5559);
or U6005 (N_6005,N_5448,N_5279);
nand U6006 (N_6006,N_5375,N_5118);
nor U6007 (N_6007,N_5592,N_5629);
nor U6008 (N_6008,N_5707,N_5586);
nor U6009 (N_6009,N_5146,N_5812);
or U6010 (N_6010,N_5740,N_5863);
nor U6011 (N_6011,N_5663,N_5410);
or U6012 (N_6012,N_5316,N_5443);
and U6013 (N_6013,N_5092,N_5441);
nand U6014 (N_6014,N_5120,N_5234);
nand U6015 (N_6015,N_5096,N_5540);
nor U6016 (N_6016,N_5357,N_5338);
or U6017 (N_6017,N_5962,N_5767);
nor U6018 (N_6018,N_5001,N_5179);
nor U6019 (N_6019,N_5518,N_5532);
or U6020 (N_6020,N_5560,N_5177);
or U6021 (N_6021,N_5896,N_5318);
and U6022 (N_6022,N_5899,N_5440);
and U6023 (N_6023,N_5045,N_5801);
nor U6024 (N_6024,N_5805,N_5932);
nand U6025 (N_6025,N_5117,N_5906);
nand U6026 (N_6026,N_5429,N_5961);
nand U6027 (N_6027,N_5423,N_5349);
or U6028 (N_6028,N_5821,N_5665);
and U6029 (N_6029,N_5736,N_5753);
nand U6030 (N_6030,N_5090,N_5706);
and U6031 (N_6031,N_5937,N_5446);
and U6032 (N_6032,N_5958,N_5968);
and U6033 (N_6033,N_5342,N_5522);
and U6034 (N_6034,N_5691,N_5565);
and U6035 (N_6035,N_5666,N_5348);
or U6036 (N_6036,N_5798,N_5933);
nor U6037 (N_6037,N_5817,N_5017);
or U6038 (N_6038,N_5310,N_5085);
nor U6039 (N_6039,N_5552,N_5721);
nor U6040 (N_6040,N_5519,N_5359);
or U6041 (N_6041,N_5340,N_5196);
and U6042 (N_6042,N_5876,N_5898);
and U6043 (N_6043,N_5389,N_5329);
and U6044 (N_6044,N_5241,N_5253);
nand U6045 (N_6045,N_5488,N_5744);
nor U6046 (N_6046,N_5047,N_5649);
nand U6047 (N_6047,N_5698,N_5972);
nand U6048 (N_6048,N_5759,N_5861);
nand U6049 (N_6049,N_5315,N_5225);
or U6050 (N_6050,N_5355,N_5347);
or U6051 (N_6051,N_5768,N_5919);
or U6052 (N_6052,N_5844,N_5764);
nor U6053 (N_6053,N_5734,N_5867);
and U6054 (N_6054,N_5800,N_5415);
xor U6055 (N_6055,N_5396,N_5401);
nand U6056 (N_6056,N_5995,N_5549);
nor U6057 (N_6057,N_5266,N_5692);
or U6058 (N_6058,N_5367,N_5135);
nor U6059 (N_6059,N_5322,N_5062);
nand U6060 (N_6060,N_5319,N_5044);
or U6061 (N_6061,N_5198,N_5683);
nor U6062 (N_6062,N_5040,N_5913);
or U6063 (N_6063,N_5137,N_5756);
nor U6064 (N_6064,N_5704,N_5151);
nand U6065 (N_6065,N_5439,N_5110);
nand U6066 (N_6066,N_5466,N_5916);
or U6067 (N_6067,N_5544,N_5645);
and U6068 (N_6068,N_5052,N_5054);
and U6069 (N_6069,N_5395,N_5028);
and U6070 (N_6070,N_5531,N_5255);
nand U6071 (N_6071,N_5681,N_5991);
nand U6072 (N_6072,N_5987,N_5953);
and U6073 (N_6073,N_5712,N_5094);
nor U6074 (N_6074,N_5901,N_5373);
or U6075 (N_6075,N_5067,N_5308);
or U6076 (N_6076,N_5020,N_5783);
nand U6077 (N_6077,N_5637,N_5926);
and U6078 (N_6078,N_5087,N_5945);
or U6079 (N_6079,N_5157,N_5163);
and U6080 (N_6080,N_5569,N_5719);
nand U6081 (N_6081,N_5143,N_5517);
and U6082 (N_6082,N_5320,N_5982);
xor U6083 (N_6083,N_5176,N_5195);
and U6084 (N_6084,N_5004,N_5461);
and U6085 (N_6085,N_5966,N_5976);
nor U6086 (N_6086,N_5141,N_5386);
nand U6087 (N_6087,N_5372,N_5891);
nor U6088 (N_6088,N_5655,N_5224);
nor U6089 (N_6089,N_5601,N_5673);
and U6090 (N_6090,N_5835,N_5999);
nand U6091 (N_6091,N_5282,N_5416);
and U6092 (N_6092,N_5302,N_5741);
nand U6093 (N_6093,N_5538,N_5097);
and U6094 (N_6094,N_5379,N_5873);
nor U6095 (N_6095,N_5589,N_5641);
or U6096 (N_6096,N_5473,N_5728);
nand U6097 (N_6097,N_5848,N_5184);
and U6098 (N_6098,N_5476,N_5152);
nor U6099 (N_6099,N_5625,N_5248);
nand U6100 (N_6100,N_5191,N_5421);
or U6101 (N_6101,N_5868,N_5530);
nand U6102 (N_6102,N_5611,N_5294);
nor U6103 (N_6103,N_5502,N_5875);
nand U6104 (N_6104,N_5053,N_5829);
or U6105 (N_6105,N_5492,N_5727);
and U6106 (N_6106,N_5938,N_5731);
or U6107 (N_6107,N_5670,N_5011);
and U6108 (N_6108,N_5192,N_5145);
and U6109 (N_6109,N_5561,N_5115);
or U6110 (N_6110,N_5831,N_5360);
or U6111 (N_6111,N_5037,N_5748);
nand U6112 (N_6112,N_5624,N_5377);
or U6113 (N_6113,N_5643,N_5159);
nor U6114 (N_6114,N_5134,N_5905);
or U6115 (N_6115,N_5923,N_5908);
nor U6116 (N_6116,N_5607,N_5482);
nand U6117 (N_6117,N_5083,N_5722);
and U6118 (N_6118,N_5022,N_5270);
nor U6119 (N_6119,N_5405,N_5675);
nand U6120 (N_6120,N_5931,N_5714);
and U6121 (N_6121,N_5804,N_5523);
or U6122 (N_6122,N_5434,N_5424);
nor U6123 (N_6123,N_5385,N_5068);
and U6124 (N_6124,N_5445,N_5006);
or U6125 (N_6125,N_5331,N_5076);
or U6126 (N_6126,N_5366,N_5301);
or U6127 (N_6127,N_5242,N_5098);
xnor U6128 (N_6128,N_5285,N_5260);
nand U6129 (N_6129,N_5393,N_5950);
and U6130 (N_6130,N_5686,N_5299);
nand U6131 (N_6131,N_5326,N_5012);
and U6132 (N_6132,N_5880,N_5243);
and U6133 (N_6133,N_5431,N_5506);
nand U6134 (N_6134,N_5892,N_5535);
and U6135 (N_6135,N_5024,N_5776);
or U6136 (N_6136,N_5351,N_5228);
or U6137 (N_6137,N_5303,N_5729);
and U6138 (N_6138,N_5368,N_5409);
or U6139 (N_6139,N_5381,N_5140);
or U6140 (N_6140,N_5955,N_5520);
nand U6141 (N_6141,N_5111,N_5742);
or U6142 (N_6142,N_5109,N_5924);
nand U6143 (N_6143,N_5993,N_5662);
or U6144 (N_6144,N_5713,N_5796);
xnor U6145 (N_6145,N_5739,N_5033);
or U6146 (N_6146,N_5646,N_5306);
nand U6147 (N_6147,N_5826,N_5394);
or U6148 (N_6148,N_5943,N_5103);
and U6149 (N_6149,N_5048,N_5882);
nor U6150 (N_6150,N_5760,N_5579);
xnor U6151 (N_6151,N_5774,N_5834);
nand U6152 (N_6152,N_5153,N_5295);
and U6153 (N_6153,N_5025,N_5564);
nand U6154 (N_6154,N_5185,N_5436);
or U6155 (N_6155,N_5486,N_5696);
nor U6156 (N_6156,N_5269,N_5886);
or U6157 (N_6157,N_5201,N_5703);
or U6158 (N_6158,N_5089,N_5638);
nor U6159 (N_6159,N_5462,N_5494);
nand U6160 (N_6160,N_5989,N_5869);
nor U6161 (N_6161,N_5472,N_5874);
nand U6162 (N_6162,N_5232,N_5178);
nand U6163 (N_6163,N_5330,N_5059);
nand U6164 (N_6164,N_5737,N_5594);
nand U6165 (N_6165,N_5934,N_5509);
nand U6166 (N_6166,N_5658,N_5885);
and U6167 (N_6167,N_5631,N_5644);
nand U6168 (N_6168,N_5197,N_5726);
xor U6169 (N_6169,N_5587,N_5262);
or U6170 (N_6170,N_5407,N_5847);
or U6171 (N_6171,N_5077,N_5674);
nand U6172 (N_6172,N_5558,N_5572);
nand U6173 (N_6173,N_5732,N_5453);
and U6174 (N_6174,N_5165,N_5216);
and U6175 (N_6175,N_5327,N_5361);
and U6176 (N_6176,N_5507,N_5226);
and U6177 (N_6177,N_5581,N_5917);
nand U6178 (N_6178,N_5842,N_5818);
and U6179 (N_6179,N_5596,N_5849);
nor U6180 (N_6180,N_5527,N_5328);
and U6181 (N_6181,N_5632,N_5845);
and U6182 (N_6182,N_5147,N_5480);
and U6183 (N_6183,N_5273,N_5806);
nand U6184 (N_6184,N_5914,N_5451);
and U6185 (N_6185,N_5705,N_5878);
and U6186 (N_6186,N_5156,N_5613);
nand U6187 (N_6187,N_5700,N_5539);
or U6188 (N_6188,N_5129,N_5747);
or U6189 (N_6189,N_5256,N_5803);
or U6190 (N_6190,N_5856,N_5877);
xnor U6191 (N_6191,N_5866,N_5229);
or U6192 (N_6192,N_5682,N_5794);
nand U6193 (N_6193,N_5050,N_5545);
or U6194 (N_6194,N_5939,N_5490);
or U6195 (N_6195,N_5030,N_5775);
and U6196 (N_6196,N_5041,N_5600);
nor U6197 (N_6197,N_5414,N_5819);
or U6198 (N_6198,N_5981,N_5034);
and U6199 (N_6199,N_5701,N_5149);
nor U6200 (N_6200,N_5566,N_5595);
nor U6201 (N_6201,N_5610,N_5404);
and U6202 (N_6202,N_5039,N_5881);
and U6203 (N_6203,N_5093,N_5591);
and U6204 (N_6204,N_5857,N_5464);
nand U6205 (N_6205,N_5419,N_5956);
or U6206 (N_6206,N_5548,N_5664);
or U6207 (N_6207,N_5846,N_5071);
nand U6208 (N_6208,N_5200,N_5936);
or U6209 (N_6209,N_5990,N_5959);
nand U6210 (N_6210,N_5257,N_5314);
and U6211 (N_6211,N_5181,N_5363);
and U6212 (N_6212,N_5227,N_5187);
nand U6213 (N_6213,N_5212,N_5555);
and U6214 (N_6214,N_5108,N_5852);
nor U6215 (N_6215,N_5980,N_5688);
nand U6216 (N_6216,N_5193,N_5026);
nand U6217 (N_6217,N_5390,N_5890);
and U6218 (N_6218,N_5161,N_5679);
and U6219 (N_6219,N_5975,N_5204);
nand U6220 (N_6220,N_5346,N_5321);
or U6221 (N_6221,N_5289,N_5223);
xor U6222 (N_6222,N_5015,N_5828);
and U6223 (N_6223,N_5286,N_5155);
nand U6224 (N_6224,N_5770,N_5944);
nand U6225 (N_6225,N_5717,N_5150);
or U6226 (N_6226,N_5487,N_5927);
and U6227 (N_6227,N_5660,N_5468);
nor U6228 (N_6228,N_5621,N_5101);
or U6229 (N_6229,N_5281,N_5883);
and U6230 (N_6230,N_5013,N_5642);
nor U6231 (N_6231,N_5469,N_5651);
nor U6232 (N_6232,N_5304,N_5554);
or U6233 (N_6233,N_5694,N_5903);
or U6234 (N_6234,N_5463,N_5275);
nor U6235 (N_6235,N_5894,N_5510);
nor U6236 (N_6236,N_5324,N_5007);
and U6237 (N_6237,N_5238,N_5231);
nand U6238 (N_6238,N_5497,N_5005);
and U6239 (N_6239,N_5183,N_5969);
and U6240 (N_6240,N_5733,N_5125);
nor U6241 (N_6241,N_5864,N_5697);
nor U6242 (N_6242,N_5757,N_5912);
or U6243 (N_6243,N_5504,N_5189);
nor U6244 (N_6244,N_5964,N_5049);
nor U6245 (N_6245,N_5259,N_5669);
nand U6246 (N_6246,N_5132,N_5384);
or U6247 (N_6247,N_5702,N_5194);
and U6248 (N_6248,N_5106,N_5751);
nand U6249 (N_6249,N_5210,N_5505);
and U6250 (N_6250,N_5970,N_5684);
nor U6251 (N_6251,N_5808,N_5277);
nor U6252 (N_6252,N_5408,N_5667);
nor U6253 (N_6253,N_5337,N_5537);
and U6254 (N_6254,N_5069,N_5716);
and U6255 (N_6255,N_5648,N_5928);
and U6256 (N_6256,N_5450,N_5075);
and U6257 (N_6257,N_5689,N_5168);
or U6258 (N_6258,N_5618,N_5743);
and U6259 (N_6259,N_5900,N_5814);
nor U6260 (N_6260,N_5317,N_5603);
and U6261 (N_6261,N_5274,N_5166);
and U6262 (N_6262,N_5358,N_5758);
nor U6263 (N_6263,N_5220,N_5810);
or U6264 (N_6264,N_5724,N_5190);
nor U6265 (N_6265,N_5654,N_5465);
and U6266 (N_6266,N_5996,N_5907);
or U6267 (N_6267,N_5915,N_5173);
nor U6268 (N_6268,N_5475,N_5426);
nor U6269 (N_6269,N_5251,N_5400);
nor U6270 (N_6270,N_5174,N_5511);
nand U6271 (N_6271,N_5171,N_5678);
or U6272 (N_6272,N_5795,N_5099);
or U6273 (N_6273,N_5278,N_5622);
and U6274 (N_6274,N_5470,N_5825);
or U6275 (N_6275,N_5895,N_5904);
or U6276 (N_6276,N_5940,N_5433);
or U6277 (N_6277,N_5838,N_5086);
nor U6278 (N_6278,N_5887,N_5571);
nor U6279 (N_6279,N_5219,N_5833);
nor U6280 (N_6280,N_5352,N_5693);
or U6281 (N_6281,N_5977,N_5738);
and U6282 (N_6282,N_5392,N_5154);
nor U6283 (N_6283,N_5640,N_5218);
nand U6284 (N_6284,N_5840,N_5988);
nand U6285 (N_6285,N_5677,N_5122);
and U6286 (N_6286,N_5889,N_5580);
nor U6287 (N_6287,N_5615,N_5634);
nor U6288 (N_6288,N_5657,N_5208);
or U6289 (N_6289,N_5633,N_5457);
nand U6290 (N_6290,N_5449,N_5428);
or U6291 (N_6291,N_5237,N_5855);
or U6292 (N_6292,N_5458,N_5870);
nor U6293 (N_6293,N_5411,N_5583);
and U6294 (N_6294,N_5827,N_5311);
nor U6295 (N_6295,N_5777,N_5807);
nor U6296 (N_6296,N_5762,N_5710);
and U6297 (N_6297,N_5483,N_5008);
or U6298 (N_6298,N_5567,N_5590);
nor U6299 (N_6299,N_5333,N_5965);
or U6300 (N_6300,N_5288,N_5172);
nor U6301 (N_6301,N_5920,N_5547);
and U6302 (N_6302,N_5056,N_5074);
nor U6303 (N_6303,N_5524,N_5388);
nor U6304 (N_6304,N_5602,N_5577);
nand U6305 (N_6305,N_5781,N_5088);
or U6306 (N_6306,N_5832,N_5499);
and U6307 (N_6307,N_5790,N_5112);
nor U6308 (N_6308,N_5459,N_5354);
or U6309 (N_6309,N_5060,N_5138);
or U6310 (N_6310,N_5182,N_5526);
or U6311 (N_6311,N_5661,N_5222);
or U6312 (N_6312,N_5100,N_5746);
and U6313 (N_6313,N_5064,N_5659);
or U6314 (N_6314,N_5160,N_5422);
or U6315 (N_6315,N_5456,N_5513);
and U6316 (N_6316,N_5144,N_5021);
and U6317 (N_6317,N_5551,N_5380);
xnor U6318 (N_6318,N_5859,N_5687);
nand U6319 (N_6319,N_5718,N_5119);
nor U6320 (N_6320,N_5325,N_5780);
or U6321 (N_6321,N_5708,N_5534);
and U6322 (N_6322,N_5065,N_5921);
or U6323 (N_6323,N_5528,N_5496);
or U6324 (N_6324,N_5574,N_5452);
nor U6325 (N_6325,N_5578,N_5576);
nor U6326 (N_6326,N_5843,N_5593);
nor U6327 (N_6327,N_5070,N_5929);
nor U6328 (N_6328,N_5820,N_5647);
and U6329 (N_6329,N_5754,N_5029);
or U6330 (N_6330,N_5822,N_5305);
and U6331 (N_6331,N_5387,N_5170);
and U6332 (N_6332,N_5263,N_5249);
and U6333 (N_6333,N_5623,N_5406);
nor U6334 (N_6334,N_5114,N_5620);
nand U6335 (N_6335,N_5205,N_5720);
or U6336 (N_6336,N_5036,N_5484);
xnor U6337 (N_6337,N_5954,N_5264);
nor U6338 (N_6338,N_5236,N_5809);
nor U6339 (N_6339,N_5180,N_5598);
xnor U6340 (N_6340,N_5376,N_5749);
nand U6341 (N_6341,N_5437,N_5951);
and U6342 (N_6342,N_5214,N_5023);
nor U6343 (N_6343,N_5402,N_5374);
nor U6344 (N_6344,N_5584,N_5058);
and U6345 (N_6345,N_5057,N_5442);
nor U6346 (N_6346,N_5312,N_5323);
and U6347 (N_6347,N_5616,N_5771);
or U6348 (N_6348,N_5252,N_5650);
nor U6349 (N_6349,N_5246,N_5427);
nor U6350 (N_6350,N_5339,N_5430);
and U6351 (N_6351,N_5345,N_5508);
or U6352 (N_6352,N_5211,N_5872);
nand U6353 (N_6353,N_5136,N_5536);
nor U6354 (N_6354,N_5772,N_5897);
nand U6355 (N_6355,N_5879,N_5002);
nor U6356 (N_6356,N_5788,N_5588);
nand U6357 (N_6357,N_5418,N_5568);
nor U6358 (N_6358,N_5126,N_5014);
nor U6359 (N_6359,N_5563,N_5709);
nand U6360 (N_6360,N_5909,N_5515);
nor U6361 (N_6361,N_5032,N_5055);
and U6362 (N_6362,N_5471,N_5091);
nand U6363 (N_6363,N_5862,N_5715);
xor U6364 (N_6364,N_5789,N_5425);
nor U6365 (N_6365,N_5503,N_5000);
and U6366 (N_6366,N_5493,N_5362);
or U6367 (N_6367,N_5910,N_5010);
and U6368 (N_6368,N_5202,N_5617);
or U6369 (N_6369,N_5292,N_5287);
and U6370 (N_6370,N_5350,N_5779);
and U6371 (N_6371,N_5478,N_5334);
xor U6372 (N_6372,N_5925,N_5343);
nor U6373 (N_6373,N_5766,N_5131);
and U6374 (N_6374,N_5290,N_5213);
nor U6375 (N_6375,N_5626,N_5998);
and U6376 (N_6376,N_5356,N_5413);
nor U6377 (N_6377,N_5148,N_5854);
nand U6378 (N_6378,N_5245,N_5474);
nand U6379 (N_6379,N_5562,N_5974);
and U6380 (N_6380,N_5019,N_5209);
and U6381 (N_6381,N_5942,N_5752);
nor U6382 (N_6382,N_5725,N_5495);
or U6383 (N_6383,N_5606,N_5271);
nand U6384 (N_6384,N_5570,N_5250);
and U6385 (N_6385,N_5997,N_5986);
and U6386 (N_6386,N_5630,N_5233);
nor U6387 (N_6387,N_5597,N_5888);
or U6388 (N_6388,N_5438,N_5284);
nor U6389 (N_6389,N_5291,N_5258);
nor U6390 (N_6390,N_5027,N_5336);
and U6391 (N_6391,N_5652,N_5142);
nor U6392 (N_6392,N_5403,N_5239);
nand U6393 (N_6393,N_5038,N_5823);
and U6394 (N_6394,N_5769,N_5957);
nor U6395 (N_6395,N_5382,N_5604);
xor U6396 (N_6396,N_5627,N_5785);
and U6397 (N_6397,N_5063,N_5792);
and U6398 (N_6398,N_5158,N_5787);
and U6399 (N_6399,N_5481,N_5051);
nor U6400 (N_6400,N_5378,N_5841);
or U6401 (N_6401,N_5985,N_5164);
and U6402 (N_6402,N_5297,N_5307);
and U6403 (N_6403,N_5946,N_5546);
or U6404 (N_6404,N_5121,N_5947);
nand U6405 (N_6405,N_5293,N_5763);
or U6406 (N_6406,N_5221,N_5116);
and U6407 (N_6407,N_5745,N_5235);
nor U6408 (N_6408,N_5557,N_5952);
and U6409 (N_6409,N_5949,N_5491);
nand U6410 (N_6410,N_5454,N_5635);
or U6411 (N_6411,N_5072,N_5398);
and U6412 (N_6412,N_5830,N_5653);
nor U6413 (N_6413,N_5203,N_5960);
nand U6414 (N_6414,N_5786,N_5383);
nor U6415 (N_6415,N_5417,N_5501);
and U6416 (N_6416,N_5850,N_5444);
nor U6417 (N_6417,N_5169,N_5217);
or U6418 (N_6418,N_5811,N_5240);
nand U6419 (N_6419,N_5107,N_5902);
or U6420 (N_6420,N_5084,N_5447);
xnor U6421 (N_6421,N_5397,N_5130);
and U6422 (N_6422,N_5298,N_5102);
nand U6423 (N_6423,N_5984,N_5296);
nand U6424 (N_6424,N_5079,N_5994);
and U6425 (N_6425,N_5542,N_5941);
nand U6426 (N_6426,N_5247,N_5477);
or U6427 (N_6427,N_5265,N_5585);
or U6428 (N_6428,N_5128,N_5978);
nor U6429 (N_6429,N_5668,N_5364);
or U6430 (N_6430,N_5365,N_5967);
or U6431 (N_6431,N_5884,N_5516);
and U6432 (N_6432,N_5533,N_5313);
or U6433 (N_6433,N_5272,N_5893);
nor U6434 (N_6434,N_5699,N_5073);
nor U6435 (N_6435,N_5973,N_5676);
and U6436 (N_6436,N_5839,N_5782);
nor U6437 (N_6437,N_5230,N_5188);
nor U6438 (N_6438,N_5061,N_5671);
nand U6439 (N_6439,N_5695,N_5186);
or U6440 (N_6440,N_5628,N_5813);
xnor U6441 (N_6441,N_5935,N_5865);
nor U6442 (N_6442,N_5918,N_5267);
nor U6443 (N_6443,N_5922,N_5018);
nor U6444 (N_6444,N_5003,N_5543);
or U6445 (N_6445,N_5761,N_5573);
nor U6446 (N_6446,N_5344,N_5080);
nor U6447 (N_6447,N_5778,N_5605);
or U6448 (N_6448,N_5199,N_5636);
and U6449 (N_6449,N_5816,N_5514);
nand U6450 (N_6450,N_5371,N_5283);
nor U6451 (N_6451,N_5575,N_5066);
and U6452 (N_6452,N_5016,N_5784);
and U6453 (N_6453,N_5500,N_5723);
nand U6454 (N_6454,N_5685,N_5521);
nor U6455 (N_6455,N_5765,N_5983);
or U6456 (N_6456,N_5948,N_5992);
and U6457 (N_6457,N_5612,N_5105);
and U6458 (N_6458,N_5215,N_5031);
xnor U6459 (N_6459,N_5979,N_5432);
nand U6460 (N_6460,N_5858,N_5435);
nand U6461 (N_6461,N_5582,N_5280);
or U6462 (N_6462,N_5341,N_5391);
or U6463 (N_6463,N_5206,N_5127);
and U6464 (N_6464,N_5479,N_5244);
xor U6465 (N_6465,N_5412,N_5773);
nor U6466 (N_6466,N_5599,N_5735);
or U6467 (N_6467,N_5750,N_5871);
nand U6468 (N_6468,N_5335,N_5971);
nand U6469 (N_6469,N_5860,N_5123);
and U6470 (N_6470,N_5420,N_5078);
or U6471 (N_6471,N_5095,N_5467);
nand U6472 (N_6472,N_5553,N_5489);
or U6473 (N_6473,N_5672,N_5309);
and U6474 (N_6474,N_5167,N_5608);
and U6475 (N_6475,N_5680,N_5369);
nor U6476 (N_6476,N_5113,N_5512);
nor U6477 (N_6477,N_5261,N_5254);
or U6478 (N_6478,N_5963,N_5836);
xor U6479 (N_6479,N_5009,N_5353);
or U6480 (N_6480,N_5104,N_5300);
nor U6481 (N_6481,N_5556,N_5730);
and U6482 (N_6482,N_5639,N_5043);
and U6483 (N_6483,N_5268,N_5656);
nor U6484 (N_6484,N_5541,N_5370);
nor U6485 (N_6485,N_5082,N_5042);
nand U6486 (N_6486,N_5332,N_5455);
nor U6487 (N_6487,N_5525,N_5529);
and U6488 (N_6488,N_5035,N_5276);
xnor U6489 (N_6489,N_5837,N_5797);
or U6490 (N_6490,N_5911,N_5139);
and U6491 (N_6491,N_5755,N_5619);
and U6492 (N_6492,N_5802,N_5175);
nor U6493 (N_6493,N_5498,N_5460);
or U6494 (N_6494,N_5690,N_5124);
nand U6495 (N_6495,N_5815,N_5793);
or U6496 (N_6496,N_5853,N_5207);
or U6497 (N_6497,N_5081,N_5791);
nand U6498 (N_6498,N_5485,N_5614);
xnor U6499 (N_6499,N_5399,N_5162);
and U6500 (N_6500,N_5217,N_5603);
nor U6501 (N_6501,N_5731,N_5560);
nor U6502 (N_6502,N_5861,N_5656);
and U6503 (N_6503,N_5542,N_5897);
or U6504 (N_6504,N_5405,N_5526);
nand U6505 (N_6505,N_5185,N_5132);
xor U6506 (N_6506,N_5550,N_5695);
or U6507 (N_6507,N_5204,N_5625);
and U6508 (N_6508,N_5239,N_5858);
nand U6509 (N_6509,N_5519,N_5972);
and U6510 (N_6510,N_5408,N_5209);
or U6511 (N_6511,N_5736,N_5453);
nand U6512 (N_6512,N_5859,N_5545);
or U6513 (N_6513,N_5950,N_5583);
and U6514 (N_6514,N_5738,N_5540);
nand U6515 (N_6515,N_5059,N_5152);
or U6516 (N_6516,N_5452,N_5381);
nor U6517 (N_6517,N_5292,N_5568);
nor U6518 (N_6518,N_5125,N_5499);
nor U6519 (N_6519,N_5535,N_5480);
and U6520 (N_6520,N_5477,N_5321);
and U6521 (N_6521,N_5057,N_5328);
and U6522 (N_6522,N_5504,N_5718);
or U6523 (N_6523,N_5515,N_5384);
or U6524 (N_6524,N_5251,N_5964);
and U6525 (N_6525,N_5236,N_5774);
and U6526 (N_6526,N_5009,N_5941);
or U6527 (N_6527,N_5099,N_5300);
or U6528 (N_6528,N_5999,N_5990);
or U6529 (N_6529,N_5897,N_5697);
nor U6530 (N_6530,N_5077,N_5683);
or U6531 (N_6531,N_5727,N_5362);
nand U6532 (N_6532,N_5120,N_5563);
nand U6533 (N_6533,N_5633,N_5207);
and U6534 (N_6534,N_5107,N_5942);
or U6535 (N_6535,N_5650,N_5417);
nor U6536 (N_6536,N_5530,N_5069);
nand U6537 (N_6537,N_5705,N_5214);
nand U6538 (N_6538,N_5582,N_5431);
xor U6539 (N_6539,N_5570,N_5869);
and U6540 (N_6540,N_5383,N_5496);
nand U6541 (N_6541,N_5521,N_5086);
nand U6542 (N_6542,N_5472,N_5796);
or U6543 (N_6543,N_5019,N_5531);
nand U6544 (N_6544,N_5928,N_5097);
or U6545 (N_6545,N_5767,N_5116);
and U6546 (N_6546,N_5023,N_5551);
xnor U6547 (N_6547,N_5517,N_5335);
nand U6548 (N_6548,N_5830,N_5053);
nand U6549 (N_6549,N_5410,N_5406);
nand U6550 (N_6550,N_5731,N_5993);
nand U6551 (N_6551,N_5478,N_5555);
nand U6552 (N_6552,N_5679,N_5368);
nor U6553 (N_6553,N_5233,N_5434);
nand U6554 (N_6554,N_5461,N_5003);
nor U6555 (N_6555,N_5611,N_5456);
nand U6556 (N_6556,N_5948,N_5116);
nand U6557 (N_6557,N_5072,N_5181);
xor U6558 (N_6558,N_5640,N_5185);
nand U6559 (N_6559,N_5325,N_5701);
or U6560 (N_6560,N_5447,N_5665);
or U6561 (N_6561,N_5943,N_5071);
or U6562 (N_6562,N_5748,N_5753);
or U6563 (N_6563,N_5336,N_5510);
xnor U6564 (N_6564,N_5041,N_5997);
or U6565 (N_6565,N_5589,N_5335);
nand U6566 (N_6566,N_5892,N_5503);
nor U6567 (N_6567,N_5000,N_5828);
nand U6568 (N_6568,N_5821,N_5998);
or U6569 (N_6569,N_5972,N_5303);
and U6570 (N_6570,N_5342,N_5238);
and U6571 (N_6571,N_5882,N_5968);
nor U6572 (N_6572,N_5934,N_5937);
nor U6573 (N_6573,N_5546,N_5376);
and U6574 (N_6574,N_5618,N_5824);
or U6575 (N_6575,N_5348,N_5512);
nor U6576 (N_6576,N_5387,N_5390);
nand U6577 (N_6577,N_5335,N_5705);
nand U6578 (N_6578,N_5697,N_5729);
nor U6579 (N_6579,N_5107,N_5060);
nor U6580 (N_6580,N_5439,N_5254);
nor U6581 (N_6581,N_5824,N_5507);
or U6582 (N_6582,N_5559,N_5734);
and U6583 (N_6583,N_5236,N_5776);
or U6584 (N_6584,N_5713,N_5596);
and U6585 (N_6585,N_5515,N_5111);
and U6586 (N_6586,N_5280,N_5496);
nand U6587 (N_6587,N_5231,N_5228);
xnor U6588 (N_6588,N_5398,N_5259);
or U6589 (N_6589,N_5810,N_5947);
nor U6590 (N_6590,N_5448,N_5845);
and U6591 (N_6591,N_5468,N_5230);
and U6592 (N_6592,N_5918,N_5189);
or U6593 (N_6593,N_5140,N_5920);
or U6594 (N_6594,N_5241,N_5984);
nand U6595 (N_6595,N_5970,N_5191);
nor U6596 (N_6596,N_5714,N_5295);
nor U6597 (N_6597,N_5914,N_5357);
nor U6598 (N_6598,N_5599,N_5860);
and U6599 (N_6599,N_5241,N_5442);
or U6600 (N_6600,N_5031,N_5353);
nor U6601 (N_6601,N_5060,N_5969);
and U6602 (N_6602,N_5134,N_5887);
and U6603 (N_6603,N_5979,N_5528);
nor U6604 (N_6604,N_5735,N_5109);
or U6605 (N_6605,N_5488,N_5005);
nand U6606 (N_6606,N_5879,N_5544);
nor U6607 (N_6607,N_5697,N_5619);
nand U6608 (N_6608,N_5423,N_5200);
and U6609 (N_6609,N_5743,N_5055);
or U6610 (N_6610,N_5924,N_5200);
and U6611 (N_6611,N_5787,N_5311);
and U6612 (N_6612,N_5177,N_5734);
or U6613 (N_6613,N_5606,N_5679);
nand U6614 (N_6614,N_5710,N_5189);
xor U6615 (N_6615,N_5923,N_5012);
nor U6616 (N_6616,N_5284,N_5942);
nand U6617 (N_6617,N_5728,N_5942);
nor U6618 (N_6618,N_5851,N_5093);
or U6619 (N_6619,N_5800,N_5412);
nand U6620 (N_6620,N_5409,N_5586);
and U6621 (N_6621,N_5175,N_5454);
nand U6622 (N_6622,N_5809,N_5518);
and U6623 (N_6623,N_5498,N_5891);
and U6624 (N_6624,N_5422,N_5196);
nand U6625 (N_6625,N_5936,N_5575);
or U6626 (N_6626,N_5755,N_5070);
nand U6627 (N_6627,N_5169,N_5645);
nand U6628 (N_6628,N_5995,N_5676);
xnor U6629 (N_6629,N_5656,N_5395);
or U6630 (N_6630,N_5757,N_5415);
and U6631 (N_6631,N_5349,N_5236);
and U6632 (N_6632,N_5572,N_5441);
or U6633 (N_6633,N_5186,N_5142);
nor U6634 (N_6634,N_5912,N_5046);
nor U6635 (N_6635,N_5235,N_5664);
nand U6636 (N_6636,N_5532,N_5698);
or U6637 (N_6637,N_5398,N_5793);
and U6638 (N_6638,N_5380,N_5865);
nand U6639 (N_6639,N_5769,N_5722);
nor U6640 (N_6640,N_5172,N_5996);
nand U6641 (N_6641,N_5222,N_5504);
nand U6642 (N_6642,N_5227,N_5132);
or U6643 (N_6643,N_5318,N_5075);
nor U6644 (N_6644,N_5919,N_5191);
and U6645 (N_6645,N_5093,N_5181);
nand U6646 (N_6646,N_5077,N_5794);
and U6647 (N_6647,N_5839,N_5102);
xor U6648 (N_6648,N_5449,N_5593);
nor U6649 (N_6649,N_5852,N_5099);
nor U6650 (N_6650,N_5347,N_5005);
or U6651 (N_6651,N_5990,N_5117);
or U6652 (N_6652,N_5958,N_5592);
and U6653 (N_6653,N_5645,N_5395);
nand U6654 (N_6654,N_5596,N_5743);
nand U6655 (N_6655,N_5087,N_5807);
nor U6656 (N_6656,N_5728,N_5076);
nand U6657 (N_6657,N_5192,N_5960);
and U6658 (N_6658,N_5453,N_5570);
and U6659 (N_6659,N_5877,N_5034);
and U6660 (N_6660,N_5767,N_5098);
or U6661 (N_6661,N_5194,N_5302);
nand U6662 (N_6662,N_5960,N_5860);
and U6663 (N_6663,N_5001,N_5748);
nor U6664 (N_6664,N_5080,N_5410);
or U6665 (N_6665,N_5941,N_5304);
or U6666 (N_6666,N_5098,N_5168);
nor U6667 (N_6667,N_5004,N_5838);
or U6668 (N_6668,N_5143,N_5516);
nand U6669 (N_6669,N_5537,N_5843);
nand U6670 (N_6670,N_5017,N_5053);
and U6671 (N_6671,N_5298,N_5551);
or U6672 (N_6672,N_5040,N_5349);
nor U6673 (N_6673,N_5799,N_5878);
nor U6674 (N_6674,N_5363,N_5340);
nor U6675 (N_6675,N_5922,N_5242);
nand U6676 (N_6676,N_5904,N_5660);
nor U6677 (N_6677,N_5567,N_5065);
nor U6678 (N_6678,N_5670,N_5783);
nand U6679 (N_6679,N_5602,N_5064);
nor U6680 (N_6680,N_5340,N_5741);
nor U6681 (N_6681,N_5675,N_5151);
nand U6682 (N_6682,N_5228,N_5713);
nand U6683 (N_6683,N_5819,N_5654);
nand U6684 (N_6684,N_5585,N_5507);
nor U6685 (N_6685,N_5045,N_5803);
and U6686 (N_6686,N_5085,N_5809);
nand U6687 (N_6687,N_5558,N_5356);
nand U6688 (N_6688,N_5724,N_5526);
nor U6689 (N_6689,N_5296,N_5806);
and U6690 (N_6690,N_5784,N_5650);
nand U6691 (N_6691,N_5616,N_5404);
and U6692 (N_6692,N_5758,N_5812);
nor U6693 (N_6693,N_5395,N_5705);
and U6694 (N_6694,N_5553,N_5344);
and U6695 (N_6695,N_5740,N_5574);
or U6696 (N_6696,N_5751,N_5703);
nand U6697 (N_6697,N_5614,N_5468);
nand U6698 (N_6698,N_5804,N_5227);
and U6699 (N_6699,N_5329,N_5924);
and U6700 (N_6700,N_5517,N_5556);
and U6701 (N_6701,N_5164,N_5716);
or U6702 (N_6702,N_5422,N_5266);
xnor U6703 (N_6703,N_5696,N_5878);
nand U6704 (N_6704,N_5588,N_5301);
and U6705 (N_6705,N_5841,N_5223);
and U6706 (N_6706,N_5365,N_5485);
nand U6707 (N_6707,N_5566,N_5868);
and U6708 (N_6708,N_5411,N_5373);
nor U6709 (N_6709,N_5309,N_5209);
or U6710 (N_6710,N_5243,N_5751);
nand U6711 (N_6711,N_5322,N_5209);
or U6712 (N_6712,N_5067,N_5186);
and U6713 (N_6713,N_5529,N_5112);
nand U6714 (N_6714,N_5314,N_5989);
nor U6715 (N_6715,N_5795,N_5382);
nor U6716 (N_6716,N_5520,N_5245);
nand U6717 (N_6717,N_5794,N_5417);
and U6718 (N_6718,N_5784,N_5677);
and U6719 (N_6719,N_5368,N_5720);
nand U6720 (N_6720,N_5698,N_5909);
nor U6721 (N_6721,N_5253,N_5050);
nor U6722 (N_6722,N_5033,N_5566);
or U6723 (N_6723,N_5535,N_5200);
or U6724 (N_6724,N_5021,N_5193);
or U6725 (N_6725,N_5403,N_5865);
and U6726 (N_6726,N_5695,N_5366);
or U6727 (N_6727,N_5456,N_5190);
nor U6728 (N_6728,N_5717,N_5160);
or U6729 (N_6729,N_5776,N_5913);
nor U6730 (N_6730,N_5385,N_5761);
nor U6731 (N_6731,N_5454,N_5172);
or U6732 (N_6732,N_5251,N_5837);
and U6733 (N_6733,N_5975,N_5507);
nand U6734 (N_6734,N_5841,N_5151);
nor U6735 (N_6735,N_5171,N_5805);
nor U6736 (N_6736,N_5074,N_5239);
nor U6737 (N_6737,N_5817,N_5721);
or U6738 (N_6738,N_5673,N_5066);
or U6739 (N_6739,N_5287,N_5133);
nand U6740 (N_6740,N_5123,N_5850);
or U6741 (N_6741,N_5802,N_5699);
or U6742 (N_6742,N_5480,N_5576);
nor U6743 (N_6743,N_5258,N_5554);
nand U6744 (N_6744,N_5913,N_5392);
and U6745 (N_6745,N_5768,N_5304);
nand U6746 (N_6746,N_5034,N_5748);
nand U6747 (N_6747,N_5041,N_5243);
or U6748 (N_6748,N_5818,N_5579);
nand U6749 (N_6749,N_5360,N_5609);
or U6750 (N_6750,N_5995,N_5200);
xnor U6751 (N_6751,N_5574,N_5287);
or U6752 (N_6752,N_5898,N_5999);
nor U6753 (N_6753,N_5456,N_5018);
or U6754 (N_6754,N_5851,N_5290);
and U6755 (N_6755,N_5844,N_5724);
nor U6756 (N_6756,N_5160,N_5493);
or U6757 (N_6757,N_5691,N_5639);
and U6758 (N_6758,N_5622,N_5993);
nand U6759 (N_6759,N_5604,N_5687);
or U6760 (N_6760,N_5959,N_5319);
and U6761 (N_6761,N_5858,N_5204);
and U6762 (N_6762,N_5932,N_5097);
or U6763 (N_6763,N_5021,N_5410);
and U6764 (N_6764,N_5335,N_5758);
nand U6765 (N_6765,N_5926,N_5477);
nand U6766 (N_6766,N_5475,N_5572);
nand U6767 (N_6767,N_5362,N_5716);
nor U6768 (N_6768,N_5360,N_5260);
nand U6769 (N_6769,N_5309,N_5390);
and U6770 (N_6770,N_5348,N_5220);
nand U6771 (N_6771,N_5757,N_5448);
nor U6772 (N_6772,N_5934,N_5532);
nor U6773 (N_6773,N_5204,N_5706);
or U6774 (N_6774,N_5252,N_5679);
nor U6775 (N_6775,N_5628,N_5593);
nor U6776 (N_6776,N_5751,N_5761);
and U6777 (N_6777,N_5302,N_5845);
or U6778 (N_6778,N_5796,N_5618);
nand U6779 (N_6779,N_5306,N_5629);
or U6780 (N_6780,N_5015,N_5134);
or U6781 (N_6781,N_5649,N_5565);
or U6782 (N_6782,N_5257,N_5716);
and U6783 (N_6783,N_5218,N_5102);
nand U6784 (N_6784,N_5545,N_5635);
nand U6785 (N_6785,N_5461,N_5164);
or U6786 (N_6786,N_5980,N_5396);
nand U6787 (N_6787,N_5777,N_5103);
nand U6788 (N_6788,N_5606,N_5793);
and U6789 (N_6789,N_5808,N_5248);
nor U6790 (N_6790,N_5875,N_5566);
and U6791 (N_6791,N_5160,N_5542);
and U6792 (N_6792,N_5532,N_5606);
or U6793 (N_6793,N_5043,N_5349);
and U6794 (N_6794,N_5924,N_5992);
or U6795 (N_6795,N_5505,N_5442);
or U6796 (N_6796,N_5115,N_5782);
nor U6797 (N_6797,N_5456,N_5302);
or U6798 (N_6798,N_5618,N_5178);
or U6799 (N_6799,N_5099,N_5114);
nor U6800 (N_6800,N_5102,N_5353);
and U6801 (N_6801,N_5678,N_5614);
and U6802 (N_6802,N_5423,N_5131);
and U6803 (N_6803,N_5177,N_5590);
and U6804 (N_6804,N_5944,N_5855);
and U6805 (N_6805,N_5013,N_5103);
nand U6806 (N_6806,N_5725,N_5454);
nor U6807 (N_6807,N_5294,N_5845);
nand U6808 (N_6808,N_5345,N_5846);
or U6809 (N_6809,N_5800,N_5212);
or U6810 (N_6810,N_5300,N_5145);
and U6811 (N_6811,N_5679,N_5480);
nand U6812 (N_6812,N_5226,N_5479);
nor U6813 (N_6813,N_5806,N_5736);
and U6814 (N_6814,N_5871,N_5500);
and U6815 (N_6815,N_5510,N_5135);
nand U6816 (N_6816,N_5993,N_5920);
and U6817 (N_6817,N_5415,N_5165);
nor U6818 (N_6818,N_5599,N_5120);
nor U6819 (N_6819,N_5268,N_5763);
nor U6820 (N_6820,N_5018,N_5308);
or U6821 (N_6821,N_5583,N_5145);
nand U6822 (N_6822,N_5368,N_5738);
nand U6823 (N_6823,N_5725,N_5411);
nand U6824 (N_6824,N_5968,N_5007);
and U6825 (N_6825,N_5982,N_5029);
nor U6826 (N_6826,N_5159,N_5859);
nand U6827 (N_6827,N_5328,N_5711);
nand U6828 (N_6828,N_5677,N_5749);
or U6829 (N_6829,N_5463,N_5545);
and U6830 (N_6830,N_5326,N_5723);
nor U6831 (N_6831,N_5046,N_5868);
and U6832 (N_6832,N_5628,N_5604);
nor U6833 (N_6833,N_5566,N_5732);
nand U6834 (N_6834,N_5062,N_5197);
or U6835 (N_6835,N_5363,N_5667);
or U6836 (N_6836,N_5348,N_5359);
nand U6837 (N_6837,N_5047,N_5485);
or U6838 (N_6838,N_5395,N_5632);
nand U6839 (N_6839,N_5125,N_5504);
nor U6840 (N_6840,N_5977,N_5584);
nand U6841 (N_6841,N_5101,N_5692);
or U6842 (N_6842,N_5890,N_5727);
or U6843 (N_6843,N_5661,N_5718);
nor U6844 (N_6844,N_5665,N_5612);
xor U6845 (N_6845,N_5037,N_5433);
or U6846 (N_6846,N_5130,N_5651);
nor U6847 (N_6847,N_5978,N_5373);
nor U6848 (N_6848,N_5545,N_5454);
nor U6849 (N_6849,N_5920,N_5890);
or U6850 (N_6850,N_5801,N_5332);
nand U6851 (N_6851,N_5573,N_5752);
nand U6852 (N_6852,N_5399,N_5106);
nor U6853 (N_6853,N_5670,N_5398);
nor U6854 (N_6854,N_5607,N_5707);
nor U6855 (N_6855,N_5539,N_5037);
and U6856 (N_6856,N_5030,N_5627);
nand U6857 (N_6857,N_5488,N_5259);
nand U6858 (N_6858,N_5392,N_5281);
nor U6859 (N_6859,N_5294,N_5547);
and U6860 (N_6860,N_5883,N_5208);
or U6861 (N_6861,N_5122,N_5891);
nor U6862 (N_6862,N_5649,N_5786);
nor U6863 (N_6863,N_5432,N_5151);
nor U6864 (N_6864,N_5497,N_5948);
nand U6865 (N_6865,N_5352,N_5708);
and U6866 (N_6866,N_5884,N_5914);
or U6867 (N_6867,N_5913,N_5148);
nor U6868 (N_6868,N_5584,N_5720);
and U6869 (N_6869,N_5582,N_5697);
or U6870 (N_6870,N_5153,N_5195);
xnor U6871 (N_6871,N_5069,N_5467);
nor U6872 (N_6872,N_5897,N_5067);
nor U6873 (N_6873,N_5508,N_5137);
nand U6874 (N_6874,N_5366,N_5120);
nand U6875 (N_6875,N_5034,N_5313);
and U6876 (N_6876,N_5426,N_5458);
or U6877 (N_6877,N_5594,N_5409);
xnor U6878 (N_6878,N_5560,N_5911);
or U6879 (N_6879,N_5164,N_5371);
or U6880 (N_6880,N_5486,N_5213);
or U6881 (N_6881,N_5492,N_5001);
and U6882 (N_6882,N_5052,N_5949);
and U6883 (N_6883,N_5958,N_5768);
nand U6884 (N_6884,N_5616,N_5804);
and U6885 (N_6885,N_5005,N_5255);
xor U6886 (N_6886,N_5699,N_5552);
or U6887 (N_6887,N_5529,N_5279);
nand U6888 (N_6888,N_5916,N_5153);
nor U6889 (N_6889,N_5483,N_5745);
or U6890 (N_6890,N_5240,N_5669);
and U6891 (N_6891,N_5842,N_5664);
nor U6892 (N_6892,N_5523,N_5798);
and U6893 (N_6893,N_5389,N_5412);
or U6894 (N_6894,N_5301,N_5846);
and U6895 (N_6895,N_5219,N_5849);
nor U6896 (N_6896,N_5421,N_5613);
nor U6897 (N_6897,N_5827,N_5449);
or U6898 (N_6898,N_5998,N_5473);
nand U6899 (N_6899,N_5408,N_5524);
or U6900 (N_6900,N_5315,N_5704);
nand U6901 (N_6901,N_5326,N_5199);
or U6902 (N_6902,N_5296,N_5623);
and U6903 (N_6903,N_5769,N_5084);
and U6904 (N_6904,N_5395,N_5129);
or U6905 (N_6905,N_5239,N_5079);
and U6906 (N_6906,N_5210,N_5368);
nand U6907 (N_6907,N_5554,N_5917);
or U6908 (N_6908,N_5663,N_5228);
and U6909 (N_6909,N_5008,N_5865);
or U6910 (N_6910,N_5762,N_5364);
and U6911 (N_6911,N_5348,N_5363);
nand U6912 (N_6912,N_5251,N_5570);
and U6913 (N_6913,N_5452,N_5682);
nor U6914 (N_6914,N_5105,N_5805);
nand U6915 (N_6915,N_5813,N_5378);
and U6916 (N_6916,N_5469,N_5579);
nor U6917 (N_6917,N_5068,N_5115);
nand U6918 (N_6918,N_5004,N_5291);
xnor U6919 (N_6919,N_5282,N_5802);
or U6920 (N_6920,N_5131,N_5039);
and U6921 (N_6921,N_5282,N_5795);
or U6922 (N_6922,N_5327,N_5644);
and U6923 (N_6923,N_5665,N_5560);
or U6924 (N_6924,N_5069,N_5910);
or U6925 (N_6925,N_5866,N_5668);
and U6926 (N_6926,N_5732,N_5009);
nor U6927 (N_6927,N_5433,N_5741);
nand U6928 (N_6928,N_5198,N_5485);
or U6929 (N_6929,N_5012,N_5557);
or U6930 (N_6930,N_5446,N_5861);
and U6931 (N_6931,N_5481,N_5747);
xor U6932 (N_6932,N_5012,N_5434);
and U6933 (N_6933,N_5983,N_5405);
and U6934 (N_6934,N_5106,N_5507);
nor U6935 (N_6935,N_5656,N_5669);
and U6936 (N_6936,N_5155,N_5182);
nand U6937 (N_6937,N_5630,N_5745);
xnor U6938 (N_6938,N_5335,N_5196);
nor U6939 (N_6939,N_5817,N_5540);
and U6940 (N_6940,N_5712,N_5946);
and U6941 (N_6941,N_5003,N_5560);
nand U6942 (N_6942,N_5170,N_5722);
nor U6943 (N_6943,N_5213,N_5137);
and U6944 (N_6944,N_5055,N_5787);
and U6945 (N_6945,N_5023,N_5204);
nor U6946 (N_6946,N_5793,N_5982);
nand U6947 (N_6947,N_5726,N_5251);
nor U6948 (N_6948,N_5325,N_5965);
nand U6949 (N_6949,N_5369,N_5836);
and U6950 (N_6950,N_5345,N_5175);
and U6951 (N_6951,N_5950,N_5759);
or U6952 (N_6952,N_5018,N_5555);
and U6953 (N_6953,N_5670,N_5565);
nor U6954 (N_6954,N_5740,N_5303);
and U6955 (N_6955,N_5180,N_5161);
and U6956 (N_6956,N_5026,N_5797);
nand U6957 (N_6957,N_5294,N_5497);
and U6958 (N_6958,N_5258,N_5422);
nand U6959 (N_6959,N_5926,N_5328);
and U6960 (N_6960,N_5273,N_5532);
nand U6961 (N_6961,N_5250,N_5891);
nand U6962 (N_6962,N_5356,N_5677);
or U6963 (N_6963,N_5551,N_5596);
and U6964 (N_6964,N_5973,N_5951);
or U6965 (N_6965,N_5550,N_5570);
or U6966 (N_6966,N_5883,N_5060);
or U6967 (N_6967,N_5940,N_5388);
or U6968 (N_6968,N_5610,N_5038);
and U6969 (N_6969,N_5024,N_5647);
nand U6970 (N_6970,N_5232,N_5233);
nand U6971 (N_6971,N_5391,N_5316);
and U6972 (N_6972,N_5894,N_5575);
nand U6973 (N_6973,N_5714,N_5475);
nor U6974 (N_6974,N_5232,N_5624);
or U6975 (N_6975,N_5778,N_5391);
nor U6976 (N_6976,N_5641,N_5445);
or U6977 (N_6977,N_5414,N_5161);
and U6978 (N_6978,N_5239,N_5648);
nand U6979 (N_6979,N_5828,N_5430);
or U6980 (N_6980,N_5472,N_5027);
or U6981 (N_6981,N_5130,N_5795);
nor U6982 (N_6982,N_5635,N_5914);
or U6983 (N_6983,N_5363,N_5858);
and U6984 (N_6984,N_5589,N_5034);
nand U6985 (N_6985,N_5147,N_5706);
xor U6986 (N_6986,N_5244,N_5439);
and U6987 (N_6987,N_5735,N_5341);
nor U6988 (N_6988,N_5871,N_5596);
or U6989 (N_6989,N_5824,N_5804);
nand U6990 (N_6990,N_5286,N_5517);
or U6991 (N_6991,N_5651,N_5693);
nor U6992 (N_6992,N_5429,N_5569);
nand U6993 (N_6993,N_5558,N_5671);
nor U6994 (N_6994,N_5254,N_5223);
nand U6995 (N_6995,N_5663,N_5098);
nor U6996 (N_6996,N_5549,N_5747);
and U6997 (N_6997,N_5240,N_5668);
nor U6998 (N_6998,N_5890,N_5646);
nand U6999 (N_6999,N_5894,N_5844);
nand U7000 (N_7000,N_6245,N_6981);
or U7001 (N_7001,N_6272,N_6439);
nor U7002 (N_7002,N_6156,N_6359);
and U7003 (N_7003,N_6696,N_6659);
or U7004 (N_7004,N_6862,N_6276);
or U7005 (N_7005,N_6226,N_6511);
nand U7006 (N_7006,N_6921,N_6767);
or U7007 (N_7007,N_6757,N_6723);
nor U7008 (N_7008,N_6894,N_6325);
nand U7009 (N_7009,N_6642,N_6362);
nand U7010 (N_7010,N_6286,N_6009);
and U7011 (N_7011,N_6728,N_6939);
or U7012 (N_7012,N_6333,N_6338);
and U7013 (N_7013,N_6208,N_6955);
nand U7014 (N_7014,N_6056,N_6024);
nor U7015 (N_7015,N_6320,N_6727);
and U7016 (N_7016,N_6539,N_6097);
and U7017 (N_7017,N_6203,N_6530);
nor U7018 (N_7018,N_6649,N_6755);
and U7019 (N_7019,N_6840,N_6700);
and U7020 (N_7020,N_6904,N_6509);
nand U7021 (N_7021,N_6315,N_6328);
nor U7022 (N_7022,N_6468,N_6706);
and U7023 (N_7023,N_6176,N_6560);
and U7024 (N_7024,N_6020,N_6703);
and U7025 (N_7025,N_6647,N_6332);
nand U7026 (N_7026,N_6622,N_6479);
and U7027 (N_7027,N_6969,N_6403);
or U7028 (N_7028,N_6788,N_6483);
or U7029 (N_7029,N_6271,N_6717);
and U7030 (N_7030,N_6592,N_6873);
or U7031 (N_7031,N_6366,N_6053);
and U7032 (N_7032,N_6316,N_6502);
nor U7033 (N_7033,N_6389,N_6889);
nor U7034 (N_7034,N_6669,N_6925);
nor U7035 (N_7035,N_6327,N_6985);
nand U7036 (N_7036,N_6780,N_6132);
or U7037 (N_7037,N_6111,N_6583);
and U7038 (N_7038,N_6668,N_6336);
or U7039 (N_7039,N_6555,N_6459);
nand U7040 (N_7040,N_6568,N_6593);
and U7041 (N_7041,N_6673,N_6861);
or U7042 (N_7042,N_6446,N_6606);
nand U7043 (N_7043,N_6265,N_6241);
or U7044 (N_7044,N_6756,N_6065);
nor U7045 (N_7045,N_6262,N_6853);
or U7046 (N_7046,N_6972,N_6629);
nor U7047 (N_7047,N_6444,N_6215);
nor U7048 (N_7048,N_6551,N_6712);
nor U7049 (N_7049,N_6405,N_6204);
and U7050 (N_7050,N_6990,N_6297);
and U7051 (N_7051,N_6538,N_6006);
or U7052 (N_7052,N_6372,N_6682);
nor U7053 (N_7053,N_6159,N_6304);
nand U7054 (N_7054,N_6662,N_6736);
and U7055 (N_7055,N_6496,N_6563);
nor U7056 (N_7056,N_6890,N_6870);
and U7057 (N_7057,N_6350,N_6998);
nand U7058 (N_7058,N_6139,N_6956);
or U7059 (N_7059,N_6733,N_6533);
or U7060 (N_7060,N_6070,N_6815);
and U7061 (N_7061,N_6710,N_6602);
nand U7062 (N_7062,N_6101,N_6772);
or U7063 (N_7063,N_6808,N_6819);
nor U7064 (N_7064,N_6516,N_6679);
nor U7065 (N_7065,N_6626,N_6303);
nor U7066 (N_7066,N_6820,N_6000);
or U7067 (N_7067,N_6515,N_6526);
nor U7068 (N_7068,N_6051,N_6517);
or U7069 (N_7069,N_6083,N_6140);
nor U7070 (N_7070,N_6237,N_6388);
or U7071 (N_7071,N_6603,N_6225);
nand U7072 (N_7072,N_6454,N_6043);
and U7073 (N_7073,N_6092,N_6289);
or U7074 (N_7074,N_6027,N_6605);
or U7075 (N_7075,N_6545,N_6506);
or U7076 (N_7076,N_6612,N_6413);
or U7077 (N_7077,N_6234,N_6514);
and U7078 (N_7078,N_6264,N_6246);
and U7079 (N_7079,N_6352,N_6151);
nor U7080 (N_7080,N_6680,N_6950);
nor U7081 (N_7081,N_6034,N_6486);
or U7082 (N_7082,N_6255,N_6404);
and U7083 (N_7083,N_6849,N_6945);
and U7084 (N_7084,N_6007,N_6192);
or U7085 (N_7085,N_6122,N_6050);
nor U7086 (N_7086,N_6635,N_6046);
nor U7087 (N_7087,N_6011,N_6209);
xor U7088 (N_7088,N_6346,N_6628);
nand U7089 (N_7089,N_6038,N_6166);
xor U7090 (N_7090,N_6595,N_6600);
nor U7091 (N_7091,N_6778,N_6010);
and U7092 (N_7092,N_6360,N_6897);
and U7093 (N_7093,N_6982,N_6731);
or U7094 (N_7094,N_6665,N_6368);
or U7095 (N_7095,N_6543,N_6186);
and U7096 (N_7096,N_6369,N_6958);
nand U7097 (N_7097,N_6052,N_6131);
and U7098 (N_7098,N_6268,N_6211);
nor U7099 (N_7099,N_6584,N_6765);
and U7100 (N_7100,N_6689,N_6285);
and U7101 (N_7101,N_6901,N_6223);
or U7102 (N_7102,N_6510,N_6570);
nand U7103 (N_7103,N_6708,N_6860);
and U7104 (N_7104,N_6040,N_6335);
nand U7105 (N_7105,N_6850,N_6764);
nand U7106 (N_7106,N_6451,N_6121);
and U7107 (N_7107,N_6216,N_6334);
nor U7108 (N_7108,N_6929,N_6800);
or U7109 (N_7109,N_6928,N_6054);
or U7110 (N_7110,N_6499,N_6907);
nor U7111 (N_7111,N_6621,N_6423);
nor U7112 (N_7112,N_6442,N_6975);
nand U7113 (N_7113,N_6127,N_6344);
nand U7114 (N_7114,N_6354,N_6089);
and U7115 (N_7115,N_6085,N_6248);
and U7116 (N_7116,N_6966,N_6856);
nand U7117 (N_7117,N_6684,N_6103);
nand U7118 (N_7118,N_6880,N_6697);
nand U7119 (N_7119,N_6394,N_6829);
nor U7120 (N_7120,N_6035,N_6419);
nand U7121 (N_7121,N_6988,N_6742);
and U7122 (N_7122,N_6899,N_6569);
nand U7123 (N_7123,N_6162,N_6702);
nand U7124 (N_7124,N_6576,N_6885);
and U7125 (N_7125,N_6721,N_6913);
and U7126 (N_7126,N_6858,N_6589);
nor U7127 (N_7127,N_6205,N_6771);
or U7128 (N_7128,N_6674,N_6283);
nand U7129 (N_7129,N_6212,N_6571);
and U7130 (N_7130,N_6566,N_6049);
nor U7131 (N_7131,N_6824,N_6746);
nor U7132 (N_7132,N_6760,N_6942);
or U7133 (N_7133,N_6292,N_6959);
nand U7134 (N_7134,N_6910,N_6147);
and U7135 (N_7135,N_6259,N_6866);
or U7136 (N_7136,N_6709,N_6676);
and U7137 (N_7137,N_6409,N_6608);
or U7138 (N_7138,N_6364,N_6830);
nand U7139 (N_7139,N_6003,N_6258);
nand U7140 (N_7140,N_6178,N_6356);
or U7141 (N_7141,N_6920,N_6012);
or U7142 (N_7142,N_6136,N_6524);
nand U7143 (N_7143,N_6585,N_6135);
and U7144 (N_7144,N_6997,N_6180);
nand U7145 (N_7145,N_6022,N_6256);
or U7146 (N_7146,N_6002,N_6298);
or U7147 (N_7147,N_6126,N_6678);
nor U7148 (N_7148,N_6618,N_6343);
nand U7149 (N_7149,N_6342,N_6337);
nor U7150 (N_7150,N_6074,N_6903);
or U7151 (N_7151,N_6695,N_6427);
or U7152 (N_7152,N_6013,N_6953);
nor U7153 (N_7153,N_6658,N_6072);
nor U7154 (N_7154,N_6965,N_6937);
and U7155 (N_7155,N_6112,N_6978);
or U7156 (N_7156,N_6523,N_6616);
nor U7157 (N_7157,N_6711,N_6408);
nand U7158 (N_7158,N_6787,N_6577);
nor U7159 (N_7159,N_6799,N_6993);
and U7160 (N_7160,N_6238,N_6411);
and U7161 (N_7161,N_6844,N_6173);
nand U7162 (N_7162,N_6469,N_6782);
nand U7163 (N_7163,N_6871,N_6923);
nand U7164 (N_7164,N_6852,N_6434);
nand U7165 (N_7165,N_6916,N_6971);
nand U7166 (N_7166,N_6478,N_6317);
or U7167 (N_7167,N_6698,N_6943);
and U7168 (N_7168,N_6888,N_6497);
or U7169 (N_7169,N_6933,N_6094);
xnor U7170 (N_7170,N_6075,N_6339);
nand U7171 (N_7171,N_6387,N_6821);
nand U7172 (N_7172,N_6740,N_6644);
nand U7173 (N_7173,N_6385,N_6763);
and U7174 (N_7174,N_6664,N_6252);
or U7175 (N_7175,N_6290,N_6474);
or U7176 (N_7176,N_6064,N_6081);
or U7177 (N_7177,N_6614,N_6004);
and U7178 (N_7178,N_6500,N_6066);
or U7179 (N_7179,N_6401,N_6519);
nand U7180 (N_7180,N_6219,N_6675);
nor U7181 (N_7181,N_6667,N_6331);
nand U7182 (N_7182,N_6417,N_6938);
and U7183 (N_7183,N_6130,N_6597);
nand U7184 (N_7184,N_6620,N_6416);
and U7185 (N_7185,N_6429,N_6594);
nor U7186 (N_7186,N_6116,N_6504);
nand U7187 (N_7187,N_6715,N_6544);
nor U7188 (N_7188,N_6100,N_6128);
and U7189 (N_7189,N_6155,N_6190);
nor U7190 (N_7190,N_6373,N_6739);
nor U7191 (N_7191,N_6690,N_6704);
xnor U7192 (N_7192,N_6875,N_6572);
nor U7193 (N_7193,N_6441,N_6816);
nand U7194 (N_7194,N_6137,N_6550);
nor U7195 (N_7195,N_6299,N_6177);
or U7196 (N_7196,N_6961,N_6008);
nand U7197 (N_7197,N_6947,N_6613);
nor U7198 (N_7198,N_6383,N_6109);
nand U7199 (N_7199,N_6810,N_6382);
nand U7200 (N_7200,N_6619,N_6438);
nor U7201 (N_7201,N_6279,N_6314);
nand U7202 (N_7202,N_6806,N_6507);
and U7203 (N_7203,N_6029,N_6859);
and U7204 (N_7204,N_6400,N_6805);
nor U7205 (N_7205,N_6573,N_6567);
and U7206 (N_7206,N_6582,N_6774);
nor U7207 (N_7207,N_6206,N_6781);
nor U7208 (N_7208,N_6980,N_6655);
and U7209 (N_7209,N_6308,N_6845);
nor U7210 (N_7210,N_6059,N_6663);
nor U7211 (N_7211,N_6776,N_6017);
xnor U7212 (N_7212,N_6227,N_6912);
or U7213 (N_7213,N_6275,N_6952);
or U7214 (N_7214,N_6872,N_6784);
and U7215 (N_7215,N_6302,N_6591);
nand U7216 (N_7216,N_6836,N_6193);
xor U7217 (N_7217,N_6183,N_6086);
and U7218 (N_7218,N_6087,N_6481);
or U7219 (N_7219,N_6123,N_6609);
nand U7220 (N_7220,N_6951,N_6494);
and U7221 (N_7221,N_6370,N_6380);
or U7222 (N_7222,N_6489,N_6882);
and U7223 (N_7223,N_6777,N_6457);
and U7224 (N_7224,N_6590,N_6179);
and U7225 (N_7225,N_6705,N_6905);
nor U7226 (N_7226,N_6475,N_6798);
nor U7227 (N_7227,N_6537,N_6433);
or U7228 (N_7228,N_6588,N_6039);
and U7229 (N_7229,N_6450,N_6987);
and U7230 (N_7230,N_6743,N_6487);
or U7231 (N_7231,N_6521,N_6527);
nor U7232 (N_7232,N_6542,N_6280);
or U7233 (N_7233,N_6847,N_6979);
nand U7234 (N_7234,N_6745,N_6973);
or U7235 (N_7235,N_6650,N_6701);
or U7236 (N_7236,N_6624,N_6552);
nor U7237 (N_7237,N_6365,N_6804);
and U7238 (N_7238,N_6495,N_6633);
or U7239 (N_7239,N_6832,N_6553);
and U7240 (N_7240,N_6440,N_6358);
nor U7241 (N_7241,N_6549,N_6071);
nor U7242 (N_7242,N_6398,N_6883);
and U7243 (N_7243,N_6986,N_6797);
and U7244 (N_7244,N_6837,N_6863);
and U7245 (N_7245,N_6758,N_6713);
and U7246 (N_7246,N_6738,N_6946);
or U7247 (N_7247,N_6707,N_6102);
nor U7248 (N_7248,N_6976,N_6175);
nor U7249 (N_7249,N_6351,N_6562);
and U7250 (N_7250,N_6324,N_6345);
nand U7251 (N_7251,N_6133,N_6014);
and U7252 (N_7252,N_6599,N_6295);
or U7253 (N_7253,N_6060,N_6250);
or U7254 (N_7254,N_6447,N_6934);
and U7255 (N_7255,N_6381,N_6386);
and U7256 (N_7256,N_6036,N_6498);
nand U7257 (N_7257,N_6586,N_6949);
nor U7258 (N_7258,N_6453,N_6842);
nand U7259 (N_7259,N_6766,N_6093);
or U7260 (N_7260,N_6724,N_6170);
nor U7261 (N_7261,N_6281,N_6813);
and U7262 (N_7262,N_6347,N_6114);
and U7263 (N_7263,N_6376,N_6125);
nand U7264 (N_7264,N_6802,N_6671);
nand U7265 (N_7265,N_6150,N_6561);
and U7266 (N_7266,N_6377,N_6834);
xnor U7267 (N_7267,N_6801,N_6005);
nor U7268 (N_7268,N_6532,N_6522);
and U7269 (N_7269,N_6535,N_6032);
nand U7270 (N_7270,N_6044,N_6967);
and U7271 (N_7271,N_6790,N_6466);
and U7272 (N_7272,N_6160,N_6232);
nand U7273 (N_7273,N_6448,N_6410);
or U7274 (N_7274,N_6931,N_6848);
and U7275 (N_7275,N_6936,N_6452);
nor U7276 (N_7276,N_6026,N_6734);
nor U7277 (N_7277,N_6422,N_6809);
and U7278 (N_7278,N_6045,N_6855);
nor U7279 (N_7279,N_6390,N_6686);
nand U7280 (N_7280,N_6445,N_6421);
nor U7281 (N_7281,N_6751,N_6243);
nand U7282 (N_7282,N_6783,N_6357);
nand U7283 (N_7283,N_6687,N_6182);
and U7284 (N_7284,N_6118,N_6720);
or U7285 (N_7285,N_6536,N_6161);
nand U7286 (N_7286,N_6233,N_6399);
nor U7287 (N_7287,N_6267,N_6718);
and U7288 (N_7288,N_6839,N_6471);
nor U7289 (N_7289,N_6305,N_6415);
and U7290 (N_7290,N_6461,N_6960);
or U7291 (N_7291,N_6754,N_6194);
and U7292 (N_7292,N_6099,N_6753);
xor U7293 (N_7293,N_6531,N_6636);
nand U7294 (N_7294,N_6991,N_6214);
or U7295 (N_7295,N_6240,N_6491);
and U7296 (N_7296,N_6814,N_6493);
nor U7297 (N_7297,N_6348,N_6310);
nor U7298 (N_7298,N_6677,N_6113);
and U7299 (N_7299,N_6048,N_6995);
nand U7300 (N_7300,N_6661,N_6999);
or U7301 (N_7301,N_6187,N_6424);
or U7302 (N_7302,N_6747,N_6490);
nor U7303 (N_7303,N_6854,N_6867);
or U7304 (N_7304,N_6098,N_6581);
nand U7305 (N_7305,N_6231,N_6646);
or U7306 (N_7306,N_6420,N_6908);
nand U7307 (N_7307,N_6886,N_6725);
and U7308 (N_7308,N_6558,N_6055);
and U7309 (N_7309,N_6312,N_6940);
or U7310 (N_7310,N_6235,N_6284);
nand U7311 (N_7311,N_6617,N_6207);
and U7312 (N_7312,N_6470,N_6104);
nand U7313 (N_7313,N_6643,N_6277);
xnor U7314 (N_7314,N_6144,N_6171);
and U7315 (N_7315,N_6230,N_6762);
or U7316 (N_7316,N_6001,N_6068);
nand U7317 (N_7317,N_6088,N_6812);
nor U7318 (N_7318,N_6898,N_6944);
and U7319 (N_7319,N_6775,N_6640);
nand U7320 (N_7320,N_6887,N_6167);
nor U7321 (N_7321,N_6282,N_6748);
and U7322 (N_7322,N_6485,N_6138);
nand U7323 (N_7323,N_6851,N_6120);
and U7324 (N_7324,N_6096,N_6915);
and U7325 (N_7325,N_6737,N_6632);
and U7326 (N_7326,N_6426,N_6463);
or U7327 (N_7327,N_6884,N_6456);
and U7328 (N_7328,N_6031,N_6579);
nand U7329 (N_7329,N_6195,N_6601);
and U7330 (N_7330,N_6393,N_6251);
nor U7331 (N_7331,N_6681,N_6091);
nand U7332 (N_7332,N_6465,N_6141);
nand U7333 (N_7333,N_6146,N_6172);
or U7334 (N_7334,N_6306,N_6768);
and U7335 (N_7335,N_6964,N_6437);
nand U7336 (N_7336,N_6529,N_6513);
and U7337 (N_7337,N_6078,N_6221);
nand U7338 (N_7338,N_6395,N_6458);
nand U7339 (N_7339,N_6648,N_6033);
nor U7340 (N_7340,N_6744,N_6367);
or U7341 (N_7341,N_6165,N_6407);
nor U7342 (N_7342,N_6874,N_6557);
nor U7343 (N_7343,N_6025,N_6021);
nand U7344 (N_7344,N_6770,N_6374);
and U7345 (N_7345,N_6525,N_6828);
or U7346 (N_7346,N_6015,N_6811);
and U7347 (N_7347,N_6287,N_6963);
nor U7348 (N_7348,N_6954,N_6501);
or U7349 (N_7349,N_6917,N_6291);
or U7350 (N_7350,N_6785,N_6418);
and U7351 (N_7351,N_6865,N_6198);
nand U7352 (N_7352,N_6547,N_6909);
or U7353 (N_7353,N_6222,N_6244);
or U7354 (N_7354,N_6154,N_6263);
nand U7355 (N_7355,N_6962,N_6984);
or U7356 (N_7356,N_6028,N_6307);
nand U7357 (N_7357,N_6069,N_6974);
or U7358 (N_7358,N_6833,N_6301);
and U7359 (N_7359,N_6197,N_6108);
and U7360 (N_7360,N_6625,N_6379);
or U7361 (N_7361,N_6846,N_6900);
and U7362 (N_7362,N_6269,N_6106);
nor U7363 (N_7363,N_6266,N_6062);
and U7364 (N_7364,N_6534,N_6587);
nand U7365 (N_7365,N_6341,N_6878);
or U7366 (N_7366,N_6795,N_6164);
and U7367 (N_7367,N_6220,N_6607);
nor U7368 (N_7368,N_6174,N_6670);
or U7369 (N_7369,N_6158,N_6124);
nor U7370 (N_7370,N_6323,N_6425);
and U7371 (N_7371,N_6996,N_6714);
nor U7372 (N_7372,N_6719,N_6631);
nand U7373 (N_7373,N_6691,N_6730);
or U7374 (N_7374,N_6129,N_6941);
nor U7375 (N_7375,N_6864,N_6615);
or U7376 (N_7376,N_6210,N_6397);
nor U7377 (N_7377,N_6548,N_6508);
nand U7378 (N_7378,N_6296,N_6148);
and U7379 (N_7379,N_6278,N_6992);
nor U7380 (N_7380,N_6432,N_6084);
and U7381 (N_7381,N_6293,N_6107);
nand U7382 (N_7382,N_6467,N_6242);
nand U7383 (N_7383,N_6330,N_6835);
nor U7384 (N_7384,N_6692,N_6412);
or U7385 (N_7385,N_6355,N_6492);
xnor U7386 (N_7386,N_6896,N_6321);
nand U7387 (N_7387,N_6857,N_6185);
nor U7388 (N_7388,N_6396,N_6948);
and U7389 (N_7389,N_6922,N_6891);
nor U7390 (N_7390,N_6482,N_6349);
nand U7391 (N_7391,N_6058,N_6391);
and U7392 (N_7392,N_6919,N_6930);
or U7393 (N_7393,N_6528,N_6779);
or U7394 (N_7394,N_6540,N_6329);
nor U7395 (N_7395,N_6803,N_6881);
nor U7396 (N_7396,N_6142,N_6163);
and U7397 (N_7397,N_6911,N_6484);
nand U7398 (N_7398,N_6077,N_6229);
nand U7399 (N_7399,N_6480,N_6565);
or U7400 (N_7400,N_6564,N_6018);
nand U7401 (N_7401,N_6598,N_6503);
or U7402 (N_7402,N_6294,N_6199);
and U7403 (N_7403,N_6634,N_6217);
nor U7404 (N_7404,N_6559,N_6639);
and U7405 (N_7405,N_6924,N_6274);
nand U7406 (N_7406,N_6657,N_6145);
nand U7407 (N_7407,N_6879,N_6823);
nand U7408 (N_7408,N_6057,N_6149);
nand U7409 (N_7409,N_6080,N_6322);
nand U7410 (N_7410,N_6716,N_6042);
nor U7411 (N_7411,N_6115,N_6554);
nor U7412 (N_7412,N_6895,N_6443);
or U7413 (N_7413,N_6968,N_6134);
or U7414 (N_7414,N_6309,N_6876);
nand U7415 (N_7415,N_6773,N_6841);
or U7416 (N_7416,N_6119,N_6652);
xor U7417 (N_7417,N_6970,N_6989);
and U7418 (N_7418,N_6604,N_6638);
and U7419 (N_7419,N_6249,N_6630);
nor U7420 (N_7420,N_6645,N_6627);
and U7421 (N_7421,N_6512,N_6406);
nand U7422 (N_7422,N_6353,N_6318);
or U7423 (N_7423,N_6082,N_6786);
or U7424 (N_7424,N_6476,N_6807);
and U7425 (N_7425,N_6750,N_6694);
nor U7426 (N_7426,N_6030,N_6273);
or U7427 (N_7427,N_6518,N_6428);
nand U7428 (N_7428,N_6983,N_6037);
xor U7429 (N_7429,N_6666,N_6656);
or U7430 (N_7430,N_6654,N_6153);
or U7431 (N_7431,N_6449,N_6201);
or U7432 (N_7432,N_6260,N_6041);
or U7433 (N_7433,N_6651,N_6371);
nand U7434 (N_7434,N_6016,N_6361);
or U7435 (N_7435,N_6090,N_6472);
and U7436 (N_7436,N_6191,N_6300);
or U7437 (N_7437,N_6105,N_6384);
and U7438 (N_7438,N_6574,N_6789);
nand U7439 (N_7439,N_6073,N_6257);
or U7440 (N_7440,N_6505,N_6761);
nor U7441 (N_7441,N_6218,N_6826);
xor U7442 (N_7442,N_6375,N_6977);
or U7443 (N_7443,N_6914,N_6076);
or U7444 (N_7444,N_6236,N_6253);
and U7445 (N_7445,N_6623,N_6430);
nor U7446 (N_7446,N_6796,N_6902);
nor U7447 (N_7447,N_6726,N_6831);
and U7448 (N_7448,N_6462,N_6892);
or U7449 (N_7449,N_6935,N_6455);
and U7450 (N_7450,N_6023,N_6213);
nor U7451 (N_7451,N_6188,N_6752);
nor U7452 (N_7452,N_6994,N_6181);
nor U7453 (N_7453,N_6117,N_6791);
and U7454 (N_7454,N_6906,N_6488);
nor U7455 (N_7455,N_6019,N_6641);
or U7456 (N_7456,N_6464,N_6288);
nor U7457 (N_7457,N_6270,N_6239);
or U7458 (N_7458,N_6957,N_6326);
nand U7459 (N_7459,N_6392,N_6402);
and U7460 (N_7460,N_6378,N_6047);
xnor U7461 (N_7461,N_6683,N_6200);
or U7462 (N_7462,N_6067,N_6869);
xor U7463 (N_7463,N_6825,N_6729);
or U7464 (N_7464,N_6722,N_6063);
nand U7465 (N_7465,N_6261,N_6580);
nor U7466 (N_7466,N_6868,N_6794);
and U7467 (N_7467,N_6313,N_6319);
and U7468 (N_7468,N_6699,N_6224);
nor U7469 (N_7469,N_6822,N_6311);
nand U7470 (N_7470,N_6556,N_6637);
nor U7471 (N_7471,N_6061,N_6672);
or U7472 (N_7472,N_6611,N_6079);
or U7473 (N_7473,N_6732,N_6110);
nor U7474 (N_7474,N_6769,N_6436);
nand U7475 (N_7475,N_6793,N_6660);
or U7476 (N_7476,N_6759,N_6254);
and U7477 (N_7477,N_6157,N_6818);
and U7478 (N_7478,N_6741,N_6228);
or U7479 (N_7479,N_6169,N_6877);
and U7480 (N_7480,N_6749,N_6596);
nand U7481 (N_7481,N_6196,N_6575);
or U7482 (N_7482,N_6578,N_6893);
xnor U7483 (N_7483,N_6610,N_6918);
and U7484 (N_7484,N_6520,N_6152);
or U7485 (N_7485,N_6927,N_6688);
or U7486 (N_7486,N_6817,N_6435);
and U7487 (N_7487,N_6827,N_6541);
nor U7488 (N_7488,N_6168,N_6932);
nand U7489 (N_7489,N_6363,N_6431);
and U7490 (N_7490,N_6693,N_6838);
nor U7491 (N_7491,N_6340,N_6247);
nand U7492 (N_7492,N_6095,N_6546);
nor U7493 (N_7493,N_6685,N_6189);
or U7494 (N_7494,N_6477,N_6473);
nand U7495 (N_7495,N_6414,N_6792);
nor U7496 (N_7496,N_6202,N_6843);
nand U7497 (N_7497,N_6653,N_6926);
nor U7498 (N_7498,N_6460,N_6143);
and U7499 (N_7499,N_6184,N_6735);
and U7500 (N_7500,N_6214,N_6882);
nand U7501 (N_7501,N_6920,N_6529);
or U7502 (N_7502,N_6821,N_6795);
and U7503 (N_7503,N_6817,N_6910);
nand U7504 (N_7504,N_6077,N_6645);
nand U7505 (N_7505,N_6867,N_6754);
nor U7506 (N_7506,N_6818,N_6993);
nand U7507 (N_7507,N_6633,N_6023);
nand U7508 (N_7508,N_6872,N_6463);
nand U7509 (N_7509,N_6103,N_6335);
nand U7510 (N_7510,N_6221,N_6216);
nand U7511 (N_7511,N_6301,N_6073);
nor U7512 (N_7512,N_6032,N_6790);
or U7513 (N_7513,N_6125,N_6998);
or U7514 (N_7514,N_6494,N_6985);
nor U7515 (N_7515,N_6195,N_6630);
nor U7516 (N_7516,N_6440,N_6392);
and U7517 (N_7517,N_6567,N_6270);
nor U7518 (N_7518,N_6095,N_6236);
or U7519 (N_7519,N_6662,N_6472);
nand U7520 (N_7520,N_6829,N_6868);
and U7521 (N_7521,N_6956,N_6428);
or U7522 (N_7522,N_6717,N_6143);
nor U7523 (N_7523,N_6505,N_6569);
or U7524 (N_7524,N_6585,N_6715);
nand U7525 (N_7525,N_6103,N_6992);
nand U7526 (N_7526,N_6574,N_6962);
and U7527 (N_7527,N_6301,N_6451);
nand U7528 (N_7528,N_6527,N_6203);
nand U7529 (N_7529,N_6172,N_6703);
or U7530 (N_7530,N_6066,N_6210);
nand U7531 (N_7531,N_6063,N_6839);
nor U7532 (N_7532,N_6097,N_6749);
nor U7533 (N_7533,N_6745,N_6957);
nor U7534 (N_7534,N_6796,N_6564);
or U7535 (N_7535,N_6622,N_6207);
or U7536 (N_7536,N_6849,N_6003);
or U7537 (N_7537,N_6251,N_6851);
or U7538 (N_7538,N_6651,N_6729);
and U7539 (N_7539,N_6392,N_6788);
nand U7540 (N_7540,N_6890,N_6694);
nand U7541 (N_7541,N_6178,N_6380);
nand U7542 (N_7542,N_6883,N_6213);
nand U7543 (N_7543,N_6961,N_6074);
or U7544 (N_7544,N_6107,N_6096);
or U7545 (N_7545,N_6255,N_6265);
or U7546 (N_7546,N_6327,N_6570);
nand U7547 (N_7547,N_6468,N_6857);
and U7548 (N_7548,N_6001,N_6683);
or U7549 (N_7549,N_6438,N_6377);
nor U7550 (N_7550,N_6838,N_6346);
and U7551 (N_7551,N_6141,N_6875);
xor U7552 (N_7552,N_6678,N_6241);
and U7553 (N_7553,N_6280,N_6290);
or U7554 (N_7554,N_6002,N_6450);
and U7555 (N_7555,N_6839,N_6998);
nand U7556 (N_7556,N_6086,N_6426);
or U7557 (N_7557,N_6348,N_6967);
nor U7558 (N_7558,N_6933,N_6632);
nor U7559 (N_7559,N_6167,N_6247);
or U7560 (N_7560,N_6421,N_6758);
and U7561 (N_7561,N_6424,N_6038);
and U7562 (N_7562,N_6193,N_6371);
and U7563 (N_7563,N_6792,N_6622);
or U7564 (N_7564,N_6349,N_6465);
nand U7565 (N_7565,N_6408,N_6414);
and U7566 (N_7566,N_6854,N_6199);
nor U7567 (N_7567,N_6569,N_6045);
nor U7568 (N_7568,N_6497,N_6180);
nand U7569 (N_7569,N_6844,N_6561);
and U7570 (N_7570,N_6889,N_6239);
or U7571 (N_7571,N_6880,N_6769);
nand U7572 (N_7572,N_6205,N_6267);
nand U7573 (N_7573,N_6708,N_6060);
nand U7574 (N_7574,N_6279,N_6541);
nor U7575 (N_7575,N_6212,N_6768);
and U7576 (N_7576,N_6657,N_6189);
nand U7577 (N_7577,N_6440,N_6255);
nand U7578 (N_7578,N_6325,N_6614);
or U7579 (N_7579,N_6126,N_6606);
nor U7580 (N_7580,N_6531,N_6060);
nand U7581 (N_7581,N_6584,N_6985);
or U7582 (N_7582,N_6276,N_6623);
and U7583 (N_7583,N_6639,N_6950);
nand U7584 (N_7584,N_6659,N_6208);
or U7585 (N_7585,N_6360,N_6676);
nand U7586 (N_7586,N_6804,N_6176);
nand U7587 (N_7587,N_6323,N_6264);
and U7588 (N_7588,N_6286,N_6707);
or U7589 (N_7589,N_6123,N_6836);
or U7590 (N_7590,N_6610,N_6173);
nand U7591 (N_7591,N_6976,N_6493);
nand U7592 (N_7592,N_6351,N_6701);
and U7593 (N_7593,N_6199,N_6515);
and U7594 (N_7594,N_6679,N_6086);
nor U7595 (N_7595,N_6788,N_6127);
and U7596 (N_7596,N_6538,N_6694);
nand U7597 (N_7597,N_6460,N_6952);
nor U7598 (N_7598,N_6296,N_6534);
or U7599 (N_7599,N_6449,N_6707);
or U7600 (N_7600,N_6615,N_6490);
and U7601 (N_7601,N_6861,N_6784);
and U7602 (N_7602,N_6321,N_6144);
or U7603 (N_7603,N_6490,N_6533);
and U7604 (N_7604,N_6372,N_6884);
or U7605 (N_7605,N_6083,N_6756);
nand U7606 (N_7606,N_6636,N_6498);
and U7607 (N_7607,N_6364,N_6057);
nand U7608 (N_7608,N_6080,N_6161);
nor U7609 (N_7609,N_6975,N_6548);
nor U7610 (N_7610,N_6029,N_6986);
and U7611 (N_7611,N_6362,N_6563);
and U7612 (N_7612,N_6222,N_6314);
nand U7613 (N_7613,N_6329,N_6420);
nor U7614 (N_7614,N_6208,N_6685);
or U7615 (N_7615,N_6227,N_6746);
xor U7616 (N_7616,N_6100,N_6394);
and U7617 (N_7617,N_6485,N_6817);
or U7618 (N_7618,N_6469,N_6286);
nor U7619 (N_7619,N_6509,N_6191);
or U7620 (N_7620,N_6546,N_6437);
nand U7621 (N_7621,N_6955,N_6706);
nor U7622 (N_7622,N_6037,N_6675);
nand U7623 (N_7623,N_6403,N_6646);
xnor U7624 (N_7624,N_6029,N_6816);
and U7625 (N_7625,N_6287,N_6939);
xor U7626 (N_7626,N_6008,N_6929);
nor U7627 (N_7627,N_6724,N_6175);
and U7628 (N_7628,N_6669,N_6117);
nor U7629 (N_7629,N_6016,N_6028);
and U7630 (N_7630,N_6216,N_6094);
and U7631 (N_7631,N_6388,N_6208);
xor U7632 (N_7632,N_6178,N_6517);
nor U7633 (N_7633,N_6459,N_6202);
nor U7634 (N_7634,N_6138,N_6109);
and U7635 (N_7635,N_6836,N_6224);
nand U7636 (N_7636,N_6491,N_6369);
nand U7637 (N_7637,N_6271,N_6668);
or U7638 (N_7638,N_6297,N_6047);
and U7639 (N_7639,N_6528,N_6938);
and U7640 (N_7640,N_6118,N_6288);
nor U7641 (N_7641,N_6481,N_6966);
nor U7642 (N_7642,N_6019,N_6732);
and U7643 (N_7643,N_6380,N_6238);
xor U7644 (N_7644,N_6880,N_6864);
nor U7645 (N_7645,N_6839,N_6059);
nor U7646 (N_7646,N_6057,N_6053);
nand U7647 (N_7647,N_6661,N_6275);
or U7648 (N_7648,N_6406,N_6937);
nor U7649 (N_7649,N_6481,N_6712);
and U7650 (N_7650,N_6665,N_6025);
nor U7651 (N_7651,N_6413,N_6146);
or U7652 (N_7652,N_6830,N_6595);
and U7653 (N_7653,N_6018,N_6624);
nand U7654 (N_7654,N_6722,N_6377);
and U7655 (N_7655,N_6862,N_6650);
nand U7656 (N_7656,N_6625,N_6793);
nor U7657 (N_7657,N_6172,N_6975);
nor U7658 (N_7658,N_6168,N_6149);
nand U7659 (N_7659,N_6377,N_6522);
xnor U7660 (N_7660,N_6700,N_6351);
nand U7661 (N_7661,N_6800,N_6089);
or U7662 (N_7662,N_6606,N_6766);
nand U7663 (N_7663,N_6131,N_6294);
or U7664 (N_7664,N_6099,N_6171);
and U7665 (N_7665,N_6006,N_6013);
nor U7666 (N_7666,N_6908,N_6331);
nand U7667 (N_7667,N_6913,N_6116);
nor U7668 (N_7668,N_6194,N_6180);
nor U7669 (N_7669,N_6799,N_6188);
or U7670 (N_7670,N_6379,N_6383);
nor U7671 (N_7671,N_6003,N_6275);
nand U7672 (N_7672,N_6138,N_6871);
nor U7673 (N_7673,N_6979,N_6323);
nor U7674 (N_7674,N_6634,N_6948);
or U7675 (N_7675,N_6117,N_6995);
and U7676 (N_7676,N_6925,N_6606);
and U7677 (N_7677,N_6993,N_6122);
nor U7678 (N_7678,N_6193,N_6204);
and U7679 (N_7679,N_6904,N_6905);
nor U7680 (N_7680,N_6035,N_6409);
or U7681 (N_7681,N_6710,N_6549);
nand U7682 (N_7682,N_6641,N_6658);
nor U7683 (N_7683,N_6192,N_6155);
and U7684 (N_7684,N_6232,N_6236);
nor U7685 (N_7685,N_6733,N_6311);
nand U7686 (N_7686,N_6994,N_6624);
nor U7687 (N_7687,N_6766,N_6719);
nor U7688 (N_7688,N_6478,N_6210);
nor U7689 (N_7689,N_6025,N_6465);
and U7690 (N_7690,N_6193,N_6921);
and U7691 (N_7691,N_6301,N_6949);
nand U7692 (N_7692,N_6712,N_6095);
or U7693 (N_7693,N_6652,N_6247);
nand U7694 (N_7694,N_6274,N_6240);
nor U7695 (N_7695,N_6177,N_6481);
or U7696 (N_7696,N_6939,N_6477);
nor U7697 (N_7697,N_6207,N_6121);
or U7698 (N_7698,N_6080,N_6193);
nor U7699 (N_7699,N_6409,N_6064);
or U7700 (N_7700,N_6380,N_6855);
nor U7701 (N_7701,N_6499,N_6381);
nand U7702 (N_7702,N_6568,N_6525);
nand U7703 (N_7703,N_6005,N_6257);
or U7704 (N_7704,N_6821,N_6519);
and U7705 (N_7705,N_6684,N_6266);
nand U7706 (N_7706,N_6250,N_6095);
nand U7707 (N_7707,N_6743,N_6666);
nand U7708 (N_7708,N_6994,N_6940);
and U7709 (N_7709,N_6273,N_6592);
nand U7710 (N_7710,N_6089,N_6351);
and U7711 (N_7711,N_6874,N_6553);
or U7712 (N_7712,N_6709,N_6139);
and U7713 (N_7713,N_6220,N_6886);
nand U7714 (N_7714,N_6760,N_6815);
xor U7715 (N_7715,N_6730,N_6737);
and U7716 (N_7716,N_6696,N_6390);
nand U7717 (N_7717,N_6702,N_6662);
and U7718 (N_7718,N_6123,N_6875);
nand U7719 (N_7719,N_6043,N_6679);
nor U7720 (N_7720,N_6287,N_6165);
and U7721 (N_7721,N_6860,N_6418);
nand U7722 (N_7722,N_6623,N_6205);
or U7723 (N_7723,N_6153,N_6656);
nand U7724 (N_7724,N_6878,N_6057);
or U7725 (N_7725,N_6719,N_6748);
nand U7726 (N_7726,N_6927,N_6147);
nand U7727 (N_7727,N_6158,N_6714);
nand U7728 (N_7728,N_6691,N_6021);
or U7729 (N_7729,N_6676,N_6342);
nand U7730 (N_7730,N_6109,N_6660);
and U7731 (N_7731,N_6317,N_6887);
nand U7732 (N_7732,N_6993,N_6218);
and U7733 (N_7733,N_6266,N_6094);
and U7734 (N_7734,N_6728,N_6324);
or U7735 (N_7735,N_6565,N_6404);
nand U7736 (N_7736,N_6537,N_6702);
nor U7737 (N_7737,N_6837,N_6042);
nor U7738 (N_7738,N_6738,N_6161);
and U7739 (N_7739,N_6093,N_6704);
nand U7740 (N_7740,N_6054,N_6977);
and U7741 (N_7741,N_6738,N_6275);
nand U7742 (N_7742,N_6168,N_6414);
nor U7743 (N_7743,N_6986,N_6195);
and U7744 (N_7744,N_6537,N_6360);
xor U7745 (N_7745,N_6214,N_6372);
and U7746 (N_7746,N_6181,N_6248);
nor U7747 (N_7747,N_6023,N_6477);
nor U7748 (N_7748,N_6807,N_6921);
nor U7749 (N_7749,N_6216,N_6851);
xnor U7750 (N_7750,N_6137,N_6041);
nand U7751 (N_7751,N_6681,N_6787);
or U7752 (N_7752,N_6074,N_6405);
nand U7753 (N_7753,N_6972,N_6756);
nor U7754 (N_7754,N_6837,N_6500);
nor U7755 (N_7755,N_6855,N_6054);
or U7756 (N_7756,N_6529,N_6951);
nand U7757 (N_7757,N_6736,N_6979);
or U7758 (N_7758,N_6308,N_6372);
nor U7759 (N_7759,N_6781,N_6768);
or U7760 (N_7760,N_6916,N_6052);
nor U7761 (N_7761,N_6255,N_6308);
or U7762 (N_7762,N_6177,N_6609);
nand U7763 (N_7763,N_6509,N_6253);
or U7764 (N_7764,N_6490,N_6655);
nand U7765 (N_7765,N_6311,N_6738);
nand U7766 (N_7766,N_6582,N_6832);
nand U7767 (N_7767,N_6936,N_6480);
nor U7768 (N_7768,N_6504,N_6111);
and U7769 (N_7769,N_6294,N_6740);
nand U7770 (N_7770,N_6517,N_6411);
and U7771 (N_7771,N_6809,N_6975);
nor U7772 (N_7772,N_6250,N_6275);
or U7773 (N_7773,N_6762,N_6998);
xnor U7774 (N_7774,N_6811,N_6500);
xnor U7775 (N_7775,N_6689,N_6241);
nand U7776 (N_7776,N_6065,N_6481);
nor U7777 (N_7777,N_6854,N_6059);
nand U7778 (N_7778,N_6000,N_6861);
nor U7779 (N_7779,N_6986,N_6465);
or U7780 (N_7780,N_6756,N_6355);
or U7781 (N_7781,N_6522,N_6877);
nand U7782 (N_7782,N_6557,N_6134);
or U7783 (N_7783,N_6130,N_6640);
or U7784 (N_7784,N_6020,N_6636);
nand U7785 (N_7785,N_6197,N_6036);
and U7786 (N_7786,N_6245,N_6957);
nor U7787 (N_7787,N_6981,N_6746);
or U7788 (N_7788,N_6058,N_6455);
nor U7789 (N_7789,N_6172,N_6533);
nand U7790 (N_7790,N_6528,N_6376);
and U7791 (N_7791,N_6037,N_6636);
nand U7792 (N_7792,N_6933,N_6580);
nand U7793 (N_7793,N_6416,N_6998);
nor U7794 (N_7794,N_6804,N_6355);
and U7795 (N_7795,N_6270,N_6289);
nand U7796 (N_7796,N_6661,N_6540);
nand U7797 (N_7797,N_6782,N_6638);
nor U7798 (N_7798,N_6963,N_6115);
and U7799 (N_7799,N_6789,N_6039);
xnor U7800 (N_7800,N_6332,N_6730);
xor U7801 (N_7801,N_6805,N_6962);
nand U7802 (N_7802,N_6282,N_6418);
nor U7803 (N_7803,N_6455,N_6712);
and U7804 (N_7804,N_6635,N_6100);
or U7805 (N_7805,N_6688,N_6486);
nand U7806 (N_7806,N_6863,N_6184);
nand U7807 (N_7807,N_6528,N_6937);
or U7808 (N_7808,N_6545,N_6276);
nand U7809 (N_7809,N_6581,N_6019);
nor U7810 (N_7810,N_6249,N_6785);
nor U7811 (N_7811,N_6635,N_6862);
nor U7812 (N_7812,N_6302,N_6028);
or U7813 (N_7813,N_6830,N_6018);
nor U7814 (N_7814,N_6203,N_6334);
and U7815 (N_7815,N_6774,N_6057);
nor U7816 (N_7816,N_6699,N_6394);
and U7817 (N_7817,N_6594,N_6941);
or U7818 (N_7818,N_6569,N_6802);
or U7819 (N_7819,N_6630,N_6567);
xor U7820 (N_7820,N_6477,N_6732);
and U7821 (N_7821,N_6242,N_6081);
nor U7822 (N_7822,N_6606,N_6792);
and U7823 (N_7823,N_6617,N_6609);
xor U7824 (N_7824,N_6868,N_6731);
and U7825 (N_7825,N_6614,N_6038);
nand U7826 (N_7826,N_6386,N_6716);
nor U7827 (N_7827,N_6854,N_6756);
or U7828 (N_7828,N_6857,N_6773);
or U7829 (N_7829,N_6552,N_6611);
nand U7830 (N_7830,N_6736,N_6177);
or U7831 (N_7831,N_6958,N_6629);
or U7832 (N_7832,N_6130,N_6595);
nor U7833 (N_7833,N_6320,N_6703);
xor U7834 (N_7834,N_6861,N_6134);
or U7835 (N_7835,N_6521,N_6157);
nand U7836 (N_7836,N_6396,N_6162);
or U7837 (N_7837,N_6019,N_6179);
nand U7838 (N_7838,N_6045,N_6212);
or U7839 (N_7839,N_6391,N_6813);
nand U7840 (N_7840,N_6284,N_6180);
or U7841 (N_7841,N_6422,N_6330);
nand U7842 (N_7842,N_6146,N_6002);
or U7843 (N_7843,N_6549,N_6572);
nand U7844 (N_7844,N_6496,N_6505);
and U7845 (N_7845,N_6957,N_6877);
or U7846 (N_7846,N_6368,N_6957);
nor U7847 (N_7847,N_6210,N_6209);
nand U7848 (N_7848,N_6244,N_6422);
nor U7849 (N_7849,N_6980,N_6127);
or U7850 (N_7850,N_6750,N_6651);
nand U7851 (N_7851,N_6529,N_6319);
nor U7852 (N_7852,N_6470,N_6578);
nand U7853 (N_7853,N_6205,N_6798);
nor U7854 (N_7854,N_6226,N_6500);
nand U7855 (N_7855,N_6781,N_6983);
nand U7856 (N_7856,N_6334,N_6277);
nor U7857 (N_7857,N_6547,N_6763);
nor U7858 (N_7858,N_6366,N_6869);
or U7859 (N_7859,N_6190,N_6669);
nand U7860 (N_7860,N_6644,N_6225);
and U7861 (N_7861,N_6694,N_6148);
nor U7862 (N_7862,N_6005,N_6748);
and U7863 (N_7863,N_6501,N_6380);
nor U7864 (N_7864,N_6314,N_6711);
nor U7865 (N_7865,N_6590,N_6771);
or U7866 (N_7866,N_6048,N_6780);
nor U7867 (N_7867,N_6608,N_6136);
or U7868 (N_7868,N_6488,N_6273);
and U7869 (N_7869,N_6799,N_6806);
nand U7870 (N_7870,N_6363,N_6100);
and U7871 (N_7871,N_6619,N_6024);
nand U7872 (N_7872,N_6723,N_6924);
nor U7873 (N_7873,N_6005,N_6871);
nand U7874 (N_7874,N_6505,N_6885);
and U7875 (N_7875,N_6982,N_6677);
and U7876 (N_7876,N_6569,N_6133);
and U7877 (N_7877,N_6262,N_6317);
nand U7878 (N_7878,N_6731,N_6322);
or U7879 (N_7879,N_6696,N_6265);
nand U7880 (N_7880,N_6347,N_6950);
or U7881 (N_7881,N_6824,N_6218);
or U7882 (N_7882,N_6608,N_6358);
nor U7883 (N_7883,N_6685,N_6386);
and U7884 (N_7884,N_6658,N_6112);
nor U7885 (N_7885,N_6227,N_6787);
or U7886 (N_7886,N_6844,N_6987);
nor U7887 (N_7887,N_6595,N_6214);
or U7888 (N_7888,N_6656,N_6185);
and U7889 (N_7889,N_6030,N_6952);
nor U7890 (N_7890,N_6327,N_6397);
nand U7891 (N_7891,N_6956,N_6017);
nand U7892 (N_7892,N_6137,N_6975);
or U7893 (N_7893,N_6119,N_6395);
and U7894 (N_7894,N_6187,N_6965);
nand U7895 (N_7895,N_6268,N_6630);
nand U7896 (N_7896,N_6168,N_6916);
and U7897 (N_7897,N_6949,N_6464);
and U7898 (N_7898,N_6220,N_6972);
nand U7899 (N_7899,N_6694,N_6340);
nand U7900 (N_7900,N_6850,N_6070);
nand U7901 (N_7901,N_6736,N_6409);
or U7902 (N_7902,N_6732,N_6442);
or U7903 (N_7903,N_6118,N_6111);
or U7904 (N_7904,N_6137,N_6213);
and U7905 (N_7905,N_6235,N_6766);
nand U7906 (N_7906,N_6068,N_6044);
or U7907 (N_7907,N_6889,N_6612);
nand U7908 (N_7908,N_6529,N_6321);
and U7909 (N_7909,N_6904,N_6352);
nor U7910 (N_7910,N_6451,N_6643);
or U7911 (N_7911,N_6934,N_6469);
or U7912 (N_7912,N_6693,N_6318);
and U7913 (N_7913,N_6046,N_6820);
nor U7914 (N_7914,N_6041,N_6998);
and U7915 (N_7915,N_6297,N_6515);
nor U7916 (N_7916,N_6505,N_6399);
nand U7917 (N_7917,N_6299,N_6132);
or U7918 (N_7918,N_6865,N_6360);
or U7919 (N_7919,N_6367,N_6857);
nor U7920 (N_7920,N_6279,N_6377);
nor U7921 (N_7921,N_6707,N_6358);
nand U7922 (N_7922,N_6773,N_6251);
and U7923 (N_7923,N_6744,N_6872);
nor U7924 (N_7924,N_6071,N_6268);
nor U7925 (N_7925,N_6162,N_6461);
and U7926 (N_7926,N_6861,N_6712);
nor U7927 (N_7927,N_6456,N_6324);
nand U7928 (N_7928,N_6102,N_6279);
nand U7929 (N_7929,N_6700,N_6355);
nor U7930 (N_7930,N_6390,N_6296);
and U7931 (N_7931,N_6217,N_6466);
nand U7932 (N_7932,N_6713,N_6112);
nor U7933 (N_7933,N_6939,N_6357);
and U7934 (N_7934,N_6352,N_6422);
or U7935 (N_7935,N_6382,N_6096);
nor U7936 (N_7936,N_6230,N_6319);
nor U7937 (N_7937,N_6255,N_6387);
nand U7938 (N_7938,N_6916,N_6927);
nor U7939 (N_7939,N_6510,N_6612);
nor U7940 (N_7940,N_6693,N_6367);
or U7941 (N_7941,N_6889,N_6329);
or U7942 (N_7942,N_6217,N_6270);
or U7943 (N_7943,N_6678,N_6725);
nor U7944 (N_7944,N_6617,N_6177);
and U7945 (N_7945,N_6043,N_6056);
or U7946 (N_7946,N_6978,N_6809);
xor U7947 (N_7947,N_6460,N_6692);
nor U7948 (N_7948,N_6700,N_6721);
nor U7949 (N_7949,N_6604,N_6625);
nor U7950 (N_7950,N_6356,N_6993);
and U7951 (N_7951,N_6961,N_6273);
nand U7952 (N_7952,N_6122,N_6558);
and U7953 (N_7953,N_6977,N_6558);
and U7954 (N_7954,N_6530,N_6428);
and U7955 (N_7955,N_6797,N_6047);
or U7956 (N_7956,N_6748,N_6972);
and U7957 (N_7957,N_6984,N_6166);
nand U7958 (N_7958,N_6918,N_6388);
or U7959 (N_7959,N_6827,N_6825);
or U7960 (N_7960,N_6782,N_6669);
nand U7961 (N_7961,N_6762,N_6823);
and U7962 (N_7962,N_6555,N_6976);
nor U7963 (N_7963,N_6737,N_6902);
or U7964 (N_7964,N_6562,N_6920);
and U7965 (N_7965,N_6015,N_6559);
and U7966 (N_7966,N_6332,N_6101);
nor U7967 (N_7967,N_6087,N_6922);
nor U7968 (N_7968,N_6657,N_6861);
or U7969 (N_7969,N_6691,N_6905);
nand U7970 (N_7970,N_6088,N_6223);
nand U7971 (N_7971,N_6098,N_6381);
nor U7972 (N_7972,N_6480,N_6415);
xor U7973 (N_7973,N_6311,N_6264);
nor U7974 (N_7974,N_6448,N_6877);
or U7975 (N_7975,N_6819,N_6504);
and U7976 (N_7976,N_6912,N_6979);
or U7977 (N_7977,N_6665,N_6799);
and U7978 (N_7978,N_6649,N_6268);
nand U7979 (N_7979,N_6710,N_6463);
nor U7980 (N_7980,N_6644,N_6932);
or U7981 (N_7981,N_6296,N_6341);
nand U7982 (N_7982,N_6018,N_6711);
nor U7983 (N_7983,N_6025,N_6269);
nor U7984 (N_7984,N_6892,N_6315);
or U7985 (N_7985,N_6868,N_6496);
and U7986 (N_7986,N_6421,N_6307);
nor U7987 (N_7987,N_6667,N_6918);
nor U7988 (N_7988,N_6467,N_6827);
or U7989 (N_7989,N_6915,N_6331);
or U7990 (N_7990,N_6994,N_6262);
or U7991 (N_7991,N_6900,N_6937);
or U7992 (N_7992,N_6963,N_6943);
or U7993 (N_7993,N_6245,N_6389);
nand U7994 (N_7994,N_6346,N_6101);
nor U7995 (N_7995,N_6868,N_6814);
nand U7996 (N_7996,N_6939,N_6751);
nor U7997 (N_7997,N_6613,N_6070);
or U7998 (N_7998,N_6088,N_6621);
or U7999 (N_7999,N_6520,N_6126);
and U8000 (N_8000,N_7391,N_7676);
and U8001 (N_8001,N_7248,N_7156);
or U8002 (N_8002,N_7850,N_7364);
or U8003 (N_8003,N_7172,N_7401);
nor U8004 (N_8004,N_7501,N_7576);
or U8005 (N_8005,N_7260,N_7509);
or U8006 (N_8006,N_7067,N_7740);
and U8007 (N_8007,N_7794,N_7059);
nand U8008 (N_8008,N_7191,N_7074);
nand U8009 (N_8009,N_7652,N_7249);
or U8010 (N_8010,N_7481,N_7578);
and U8011 (N_8011,N_7962,N_7843);
xor U8012 (N_8012,N_7035,N_7782);
or U8013 (N_8013,N_7650,N_7881);
and U8014 (N_8014,N_7762,N_7193);
nor U8015 (N_8015,N_7678,N_7187);
nand U8016 (N_8016,N_7950,N_7551);
or U8017 (N_8017,N_7824,N_7980);
and U8018 (N_8018,N_7918,N_7791);
nor U8019 (N_8019,N_7241,N_7148);
xnor U8020 (N_8020,N_7434,N_7817);
nor U8021 (N_8021,N_7031,N_7004);
or U8022 (N_8022,N_7381,N_7795);
or U8023 (N_8023,N_7094,N_7251);
nand U8024 (N_8024,N_7126,N_7258);
or U8025 (N_8025,N_7185,N_7211);
or U8026 (N_8026,N_7407,N_7362);
or U8027 (N_8027,N_7750,N_7257);
nand U8028 (N_8028,N_7266,N_7838);
nand U8029 (N_8029,N_7759,N_7468);
nand U8030 (N_8030,N_7237,N_7394);
or U8031 (N_8031,N_7844,N_7463);
nor U8032 (N_8032,N_7124,N_7641);
nand U8033 (N_8033,N_7115,N_7246);
nand U8034 (N_8034,N_7028,N_7596);
nand U8035 (N_8035,N_7776,N_7620);
nor U8036 (N_8036,N_7868,N_7316);
and U8037 (N_8037,N_7546,N_7870);
or U8038 (N_8038,N_7669,N_7693);
and U8039 (N_8039,N_7570,N_7934);
xnor U8040 (N_8040,N_7793,N_7419);
nand U8041 (N_8041,N_7743,N_7819);
nor U8042 (N_8042,N_7517,N_7347);
nand U8043 (N_8043,N_7041,N_7597);
and U8044 (N_8044,N_7385,N_7555);
nor U8045 (N_8045,N_7787,N_7001);
or U8046 (N_8046,N_7536,N_7779);
and U8047 (N_8047,N_7984,N_7305);
and U8048 (N_8048,N_7872,N_7482);
nand U8049 (N_8049,N_7919,N_7282);
or U8050 (N_8050,N_7209,N_7869);
nand U8051 (N_8051,N_7725,N_7814);
or U8052 (N_8052,N_7096,N_7600);
or U8053 (N_8053,N_7013,N_7646);
or U8054 (N_8054,N_7135,N_7447);
or U8055 (N_8055,N_7518,N_7616);
nand U8056 (N_8056,N_7055,N_7681);
nand U8057 (N_8057,N_7890,N_7525);
or U8058 (N_8058,N_7532,N_7489);
and U8059 (N_8059,N_7713,N_7139);
or U8060 (N_8060,N_7704,N_7141);
nand U8061 (N_8061,N_7549,N_7162);
or U8062 (N_8062,N_7125,N_7229);
or U8063 (N_8063,N_7097,N_7803);
nor U8064 (N_8064,N_7076,N_7866);
and U8065 (N_8065,N_7465,N_7886);
nand U8066 (N_8066,N_7163,N_7998);
and U8067 (N_8067,N_7806,N_7816);
nor U8068 (N_8068,N_7330,N_7025);
nor U8069 (N_8069,N_7588,N_7907);
and U8070 (N_8070,N_7580,N_7286);
and U8071 (N_8071,N_7747,N_7414);
nand U8072 (N_8072,N_7514,N_7195);
and U8073 (N_8073,N_7217,N_7686);
or U8074 (N_8074,N_7710,N_7810);
and U8075 (N_8075,N_7512,N_7317);
and U8076 (N_8076,N_7310,N_7508);
nor U8077 (N_8077,N_7994,N_7647);
or U8078 (N_8078,N_7991,N_7622);
and U8079 (N_8079,N_7052,N_7495);
nand U8080 (N_8080,N_7219,N_7377);
or U8081 (N_8081,N_7199,N_7002);
nor U8082 (N_8082,N_7781,N_7638);
and U8083 (N_8083,N_7941,N_7497);
and U8084 (N_8084,N_7812,N_7329);
and U8085 (N_8085,N_7174,N_7021);
nor U8086 (N_8086,N_7978,N_7098);
nor U8087 (N_8087,N_7674,N_7081);
and U8088 (N_8088,N_7830,N_7905);
nor U8089 (N_8089,N_7421,N_7550);
and U8090 (N_8090,N_7823,N_7737);
nand U8091 (N_8091,N_7995,N_7389);
nand U8092 (N_8092,N_7717,N_7348);
nand U8093 (N_8093,N_7661,N_7416);
nor U8094 (N_8094,N_7289,N_7190);
nand U8095 (N_8095,N_7488,N_7937);
nor U8096 (N_8096,N_7399,N_7768);
nand U8097 (N_8097,N_7408,N_7287);
nand U8098 (N_8098,N_7851,N_7105);
nand U8099 (N_8099,N_7775,N_7274);
or U8100 (N_8100,N_7037,N_7335);
nand U8101 (N_8101,N_7227,N_7152);
nand U8102 (N_8102,N_7433,N_7179);
xnor U8103 (N_8103,N_7748,N_7343);
nand U8104 (N_8104,N_7864,N_7757);
or U8105 (N_8105,N_7080,N_7897);
nor U8106 (N_8106,N_7986,N_7077);
nand U8107 (N_8107,N_7023,N_7792);
nor U8108 (N_8108,N_7606,N_7267);
nand U8109 (N_8109,N_7593,N_7261);
xnor U8110 (N_8110,N_7306,N_7507);
nor U8111 (N_8111,N_7671,N_7772);
nor U8112 (N_8112,N_7062,N_7976);
and U8113 (N_8113,N_7208,N_7635);
and U8114 (N_8114,N_7965,N_7624);
or U8115 (N_8115,N_7689,N_7788);
nor U8116 (N_8116,N_7902,N_7605);
or U8117 (N_8117,N_7233,N_7104);
nor U8118 (N_8118,N_7832,N_7958);
and U8119 (N_8119,N_7977,N_7836);
nand U8120 (N_8120,N_7235,N_7140);
nand U8121 (N_8121,N_7167,N_7093);
or U8122 (N_8122,N_7513,N_7018);
or U8123 (N_8123,N_7608,N_7006);
nand U8124 (N_8124,N_7974,N_7559);
or U8125 (N_8125,N_7961,N_7764);
and U8126 (N_8126,N_7545,N_7130);
and U8127 (N_8127,N_7528,N_7665);
nor U8128 (N_8128,N_7276,N_7168);
or U8129 (N_8129,N_7420,N_7904);
nor U8130 (N_8130,N_7415,N_7302);
nand U8131 (N_8131,N_7562,N_7972);
or U8132 (N_8132,N_7291,N_7510);
or U8133 (N_8133,N_7412,N_7715);
nor U8134 (N_8134,N_7034,N_7284);
nor U8135 (N_8135,N_7822,N_7427);
nor U8136 (N_8136,N_7320,N_7595);
and U8137 (N_8137,N_7084,N_7520);
and U8138 (N_8138,N_7075,N_7541);
nand U8139 (N_8139,N_7766,N_7022);
or U8140 (N_8140,N_7802,N_7656);
nor U8141 (N_8141,N_7753,N_7568);
and U8142 (N_8142,N_7090,N_7065);
or U8143 (N_8143,N_7503,N_7631);
nor U8144 (N_8144,N_7540,N_7117);
or U8145 (N_8145,N_7238,N_7042);
nand U8146 (N_8146,N_7599,N_7371);
xnor U8147 (N_8147,N_7672,N_7292);
and U8148 (N_8148,N_7679,N_7591);
and U8149 (N_8149,N_7202,N_7945);
or U8150 (N_8150,N_7829,N_7709);
or U8151 (N_8151,N_7376,N_7259);
and U8152 (N_8152,N_7194,N_7628);
nand U8153 (N_8153,N_7039,N_7040);
nand U8154 (N_8154,N_7275,N_7438);
or U8155 (N_8155,N_7707,N_7192);
nor U8156 (N_8156,N_7048,N_7321);
and U8157 (N_8157,N_7123,N_7724);
or U8158 (N_8158,N_7149,N_7842);
nand U8159 (N_8159,N_7761,N_7845);
nand U8160 (N_8160,N_7653,N_7086);
nor U8161 (N_8161,N_7848,N_7121);
or U8162 (N_8162,N_7887,N_7673);
or U8163 (N_8163,N_7754,N_7563);
nor U8164 (N_8164,N_7623,N_7334);
or U8165 (N_8165,N_7425,N_7240);
nand U8166 (N_8166,N_7129,N_7177);
nor U8167 (N_8167,N_7049,N_7901);
nor U8168 (N_8168,N_7380,N_7144);
xor U8169 (N_8169,N_7437,N_7262);
nand U8170 (N_8170,N_7840,N_7891);
and U8171 (N_8171,N_7307,N_7309);
and U8172 (N_8172,N_7708,N_7223);
and U8173 (N_8173,N_7378,N_7327);
nand U8174 (N_8174,N_7370,N_7756);
nand U8175 (N_8175,N_7279,N_7728);
or U8176 (N_8176,N_7138,N_7429);
or U8177 (N_8177,N_7214,N_7703);
nand U8178 (N_8178,N_7813,N_7346);
or U8179 (N_8179,N_7873,N_7110);
or U8180 (N_8180,N_7175,N_7957);
nand U8181 (N_8181,N_7727,N_7197);
nand U8182 (N_8182,N_7657,N_7083);
and U8183 (N_8183,N_7479,N_7889);
and U8184 (N_8184,N_7831,N_7734);
nand U8185 (N_8185,N_7614,N_7119);
and U8186 (N_8186,N_7044,N_7353);
or U8187 (N_8187,N_7594,N_7150);
or U8188 (N_8188,N_7752,N_7230);
or U8189 (N_8189,N_7894,N_7494);
nor U8190 (N_8190,N_7103,N_7397);
and U8191 (N_8191,N_7472,N_7553);
or U8192 (N_8192,N_7629,N_7654);
and U8193 (N_8193,N_7834,N_7592);
and U8194 (N_8194,N_7527,N_7383);
or U8195 (N_8195,N_7366,N_7454);
xor U8196 (N_8196,N_7966,N_7224);
nand U8197 (N_8197,N_7645,N_7981);
and U8198 (N_8198,N_7572,N_7443);
nand U8199 (N_8199,N_7263,N_7712);
nor U8200 (N_8200,N_7231,N_7091);
and U8201 (N_8201,N_7045,N_7333);
and U8202 (N_8202,N_7642,N_7909);
nand U8203 (N_8203,N_7272,N_7535);
nand U8204 (N_8204,N_7145,N_7344);
and U8205 (N_8205,N_7804,N_7243);
nor U8206 (N_8206,N_7604,N_7173);
or U8207 (N_8207,N_7992,N_7906);
nor U8208 (N_8208,N_7456,N_7565);
nor U8209 (N_8209,N_7921,N_7644);
nand U8210 (N_8210,N_7648,N_7867);
nand U8211 (N_8211,N_7032,N_7857);
nor U8212 (N_8212,N_7127,N_7484);
nand U8213 (N_8213,N_7863,N_7351);
nor U8214 (N_8214,N_7726,N_7388);
and U8215 (N_8215,N_7200,N_7337);
or U8216 (N_8216,N_7999,N_7422);
xnor U8217 (N_8217,N_7714,N_7155);
and U8218 (N_8218,N_7960,N_7982);
nand U8219 (N_8219,N_7809,N_7464);
or U8220 (N_8220,N_7142,N_7521);
or U8221 (N_8221,N_7692,N_7931);
and U8222 (N_8222,N_7170,N_7970);
nor U8223 (N_8223,N_7896,N_7137);
nor U8224 (N_8224,N_7690,N_7299);
and U8225 (N_8225,N_7837,N_7893);
or U8226 (N_8226,N_7213,N_7718);
nor U8227 (N_8227,N_7311,N_7232);
nor U8228 (N_8228,N_7607,N_7016);
or U8229 (N_8229,N_7496,N_7092);
and U8230 (N_8230,N_7571,N_7448);
nor U8231 (N_8231,N_7908,N_7892);
or U8232 (N_8232,N_7057,N_7051);
or U8233 (N_8233,N_7858,N_7393);
nor U8234 (N_8234,N_7273,N_7332);
nand U8235 (N_8235,N_7755,N_7552);
nor U8236 (N_8236,N_7988,N_7786);
and U8237 (N_8237,N_7739,N_7574);
or U8238 (N_8238,N_7298,N_7108);
nor U8239 (N_8239,N_7369,N_7916);
nand U8240 (N_8240,N_7296,N_7205);
nand U8241 (N_8241,N_7968,N_7914);
or U8242 (N_8242,N_7539,N_7688);
and U8243 (N_8243,N_7349,N_7630);
nand U8244 (N_8244,N_7668,N_7418);
and U8245 (N_8245,N_7354,N_7825);
nand U8246 (N_8246,N_7491,N_7312);
or U8247 (N_8247,N_7745,N_7112);
or U8248 (N_8248,N_7967,N_7729);
nor U8249 (N_8249,N_7885,N_7963);
and U8250 (N_8250,N_7506,N_7923);
nor U8251 (N_8251,N_7461,N_7722);
and U8252 (N_8252,N_7721,N_7070);
or U8253 (N_8253,N_7660,N_7345);
nor U8254 (N_8254,N_7990,N_7053);
nand U8255 (N_8255,N_7038,N_7453);
and U8256 (N_8256,N_7993,N_7392);
and U8257 (N_8257,N_7949,N_7452);
or U8258 (N_8258,N_7969,N_7424);
and U8259 (N_8259,N_7365,N_7435);
xor U8260 (N_8260,N_7774,N_7212);
or U8261 (N_8261,N_7181,N_7439);
nand U8262 (N_8262,N_7485,N_7655);
and U8263 (N_8263,N_7701,N_7581);
nor U8264 (N_8264,N_7475,N_7387);
or U8265 (N_8265,N_7215,N_7490);
and U8266 (N_8266,N_7136,N_7043);
nand U8267 (N_8267,N_7164,N_7723);
and U8268 (N_8268,N_7944,N_7663);
nor U8269 (N_8269,N_7883,N_7114);
and U8270 (N_8270,N_7856,N_7554);
and U8271 (N_8271,N_7132,N_7171);
and U8272 (N_8272,N_7471,N_7297);
or U8273 (N_8273,N_7796,N_7303);
or U8274 (N_8274,N_7113,N_7880);
and U8275 (N_8275,N_7178,N_7293);
nor U8276 (N_8276,N_7165,N_7011);
and U8277 (N_8277,N_7158,N_7854);
and U8278 (N_8278,N_7504,N_7799);
or U8279 (N_8279,N_7499,N_7470);
and U8280 (N_8280,N_7946,N_7698);
nor U8281 (N_8281,N_7106,N_7515);
nor U8282 (N_8282,N_7151,N_7010);
or U8283 (N_8283,N_7069,N_7033);
nand U8284 (N_8284,N_7860,N_7947);
or U8285 (N_8285,N_7898,N_7085);
or U8286 (N_8286,N_7102,N_7847);
nor U8287 (N_8287,N_7956,N_7820);
nor U8288 (N_8288,N_7411,N_7537);
and U8289 (N_8289,N_7720,N_7524);
nand U8290 (N_8290,N_7483,N_7939);
nand U8291 (N_8291,N_7543,N_7256);
nand U8292 (N_8292,N_7073,N_7015);
or U8293 (N_8293,N_7811,N_7331);
nand U8294 (N_8294,N_7458,N_7245);
and U8295 (N_8295,N_7099,N_7875);
or U8296 (N_8296,N_7615,N_7128);
nand U8297 (N_8297,N_7818,N_7925);
nand U8298 (N_8298,N_7575,N_7500);
and U8299 (N_8299,N_7932,N_7254);
and U8300 (N_8300,N_7912,N_7432);
nor U8301 (N_8301,N_7498,N_7785);
or U8302 (N_8302,N_7882,N_7473);
and U8303 (N_8303,N_7560,N_7783);
nand U8304 (N_8304,N_7955,N_7928);
and U8305 (N_8305,N_7402,N_7198);
or U8306 (N_8306,N_7731,N_7460);
nand U8307 (N_8307,N_7161,N_7627);
or U8308 (N_8308,N_7180,N_7643);
nand U8309 (N_8309,N_7711,N_7079);
or U8310 (N_8310,N_7670,N_7544);
nor U8311 (N_8311,N_7603,N_7699);
nand U8312 (N_8312,N_7884,N_7801);
or U8313 (N_8313,N_7784,N_7072);
or U8314 (N_8314,N_7933,N_7036);
nand U8315 (N_8315,N_7579,N_7954);
or U8316 (N_8316,N_7691,N_7428);
nand U8317 (N_8317,N_7805,N_7056);
or U8318 (N_8318,N_7935,N_7511);
and U8319 (N_8319,N_7147,N_7095);
nand U8320 (N_8320,N_7294,N_7538);
nor U8321 (N_8321,N_7278,N_7859);
nor U8322 (N_8322,N_7462,N_7236);
nand U8323 (N_8323,N_7012,N_7295);
xnor U8324 (N_8324,N_7697,N_7000);
nor U8325 (N_8325,N_7478,N_7951);
nand U8326 (N_8326,N_7913,N_7154);
nor U8327 (N_8327,N_7852,N_7242);
nor U8328 (N_8328,N_7009,N_7066);
nand U8329 (N_8329,N_7373,N_7474);
nor U8330 (N_8330,N_7457,N_7153);
nand U8331 (N_8331,N_7952,N_7610);
nor U8332 (N_8332,N_7247,N_7706);
or U8333 (N_8333,N_7220,N_7780);
and U8334 (N_8334,N_7542,N_7502);
and U8335 (N_8335,N_7221,N_7157);
or U8336 (N_8336,N_7319,N_7064);
nor U8337 (N_8337,N_7953,N_7100);
nor U8338 (N_8338,N_7336,N_7915);
or U8339 (N_8339,N_7027,N_7751);
nand U8340 (N_8340,N_7736,N_7683);
nand U8341 (N_8341,N_7210,N_7798);
or U8342 (N_8342,N_7547,N_7760);
or U8343 (N_8343,N_7398,N_7356);
and U8344 (N_8344,N_7228,N_7900);
and U8345 (N_8345,N_7390,N_7612);
nor U8346 (N_8346,N_7815,N_7446);
and U8347 (N_8347,N_7451,N_7973);
nor U8348 (N_8348,N_7531,N_7586);
nor U8349 (N_8349,N_7030,N_7269);
or U8350 (N_8350,N_7871,N_7618);
nor U8351 (N_8351,N_7146,N_7120);
or U8352 (N_8352,N_7265,N_7361);
nor U8353 (N_8353,N_7455,N_7003);
and U8354 (N_8354,N_7417,N_7878);
or U8355 (N_8355,N_7664,N_7920);
and U8356 (N_8356,N_7216,N_7324);
nand U8357 (N_8357,N_7938,N_7116);
nor U8358 (N_8358,N_7322,N_7403);
or U8359 (N_8359,N_7964,N_7617);
nor U8360 (N_8360,N_7800,N_7008);
nor U8361 (N_8361,N_7839,N_7476);
and U8362 (N_8362,N_7060,N_7078);
and U8363 (N_8363,N_7328,N_7583);
nand U8364 (N_8364,N_7063,N_7379);
nand U8365 (N_8365,N_7625,N_7769);
nand U8366 (N_8366,N_7087,N_7619);
nor U8367 (N_8367,N_7742,N_7926);
nor U8368 (N_8368,N_7410,N_7109);
and U8369 (N_8369,N_7395,N_7314);
or U8370 (N_8370,N_7971,N_7406);
or U8371 (N_8371,N_7133,N_7758);
and U8372 (N_8372,N_7024,N_7469);
nand U8373 (N_8373,N_7684,N_7253);
nand U8374 (N_8374,N_7268,N_7225);
or U8375 (N_8375,N_7396,N_7855);
and U8376 (N_8376,N_7738,N_7640);
or U8377 (N_8377,N_7061,N_7649);
nand U8378 (N_8378,N_7598,N_7888);
nor U8379 (N_8379,N_7368,N_7765);
nor U8380 (N_8380,N_7413,N_7360);
nor U8381 (N_8381,N_7749,N_7930);
nor U8382 (N_8382,N_7486,N_7404);
or U8383 (N_8383,N_7522,N_7300);
or U8384 (N_8384,N_7985,N_7493);
nand U8385 (N_8385,N_7621,N_7874);
and U8386 (N_8386,N_7357,N_7771);
nor U8387 (N_8387,N_7735,N_7534);
or U8388 (N_8388,N_7666,N_7853);
nor U8389 (N_8389,N_7088,N_7778);
and U8390 (N_8390,N_7677,N_7160);
or U8391 (N_8391,N_7741,N_7876);
nand U8392 (N_8392,N_7903,N_7341);
and U8393 (N_8393,N_7505,N_7071);
nand U8394 (N_8394,N_7255,N_7548);
or U8395 (N_8395,N_7558,N_7271);
nand U8396 (N_8396,N_7444,N_7226);
or U8397 (N_8397,N_7182,N_7050);
nor U8398 (N_8398,N_7359,N_7441);
and U8399 (N_8399,N_7917,N_7252);
nand U8400 (N_8400,N_7662,N_7516);
and U8401 (N_8401,N_7440,N_7431);
or U8402 (N_8402,N_7323,N_7667);
nor U8403 (N_8403,N_7639,N_7459);
nor U8404 (N_8404,N_7201,N_7636);
and U8405 (N_8405,N_7005,N_7702);
xor U8406 (N_8406,N_7159,N_7131);
or U8407 (N_8407,N_7582,N_7340);
nor U8408 (N_8408,N_7445,N_7046);
or U8409 (N_8409,N_7218,N_7899);
or U8410 (N_8410,N_7204,N_7118);
nor U8411 (N_8411,N_7358,N_7590);
and U8412 (N_8412,N_7849,N_7339);
nor U8413 (N_8413,N_7487,N_7313);
nand U8414 (N_8414,N_7658,N_7659);
nor U8415 (N_8415,N_7283,N_7557);
or U8416 (N_8416,N_7700,N_7315);
and U8417 (N_8417,N_7694,N_7533);
or U8418 (N_8418,N_7601,N_7430);
and U8419 (N_8419,N_7355,N_7405);
or U8420 (N_8420,N_7186,N_7007);
nand U8421 (N_8421,N_7277,N_7996);
xor U8422 (N_8422,N_7566,N_7111);
nor U8423 (N_8423,N_7573,N_7338);
and U8424 (N_8424,N_7014,N_7523);
nand U8425 (N_8425,N_7746,N_7234);
nand U8426 (N_8426,N_7047,N_7196);
and U8427 (N_8427,N_7569,N_7342);
or U8428 (N_8428,N_7927,N_7203);
nor U8429 (N_8429,N_7773,N_7763);
nand U8430 (N_8430,N_7288,N_7979);
or U8431 (N_8431,N_7632,N_7790);
and U8432 (N_8432,N_7068,N_7910);
nor U8433 (N_8433,N_7318,N_7519);
or U8434 (N_8434,N_7375,N_7634);
nand U8435 (N_8435,N_7280,N_7695);
or U8436 (N_8436,N_7019,N_7244);
or U8437 (N_8437,N_7384,N_7101);
or U8438 (N_8438,N_7166,N_7530);
nor U8439 (N_8439,N_7367,N_7833);
nor U8440 (N_8440,N_7222,N_7026);
nor U8441 (N_8441,N_7685,N_7556);
or U8442 (N_8442,N_7449,N_7959);
and U8443 (N_8443,N_7564,N_7911);
and U8444 (N_8444,N_7730,N_7719);
and U8445 (N_8445,N_7054,N_7997);
and U8446 (N_8446,N_7651,N_7613);
nor U8447 (N_8447,N_7602,N_7058);
or U8448 (N_8448,N_7584,N_7477);
nand U8449 (N_8449,N_7480,N_7561);
or U8450 (N_8450,N_7442,N_7983);
or U8451 (N_8451,N_7020,N_7895);
nand U8452 (N_8452,N_7675,N_7176);
and U8453 (N_8453,N_7924,N_7936);
and U8454 (N_8454,N_7865,N_7325);
nand U8455 (N_8455,N_7363,N_7987);
or U8456 (N_8456,N_7821,N_7436);
or U8457 (N_8457,N_7029,N_7922);
nor U8458 (N_8458,N_7777,N_7835);
nor U8459 (N_8459,N_7732,N_7169);
or U8460 (N_8460,N_7352,N_7637);
or U8461 (N_8461,N_7250,N_7687);
and U8462 (N_8462,N_7807,N_7290);
or U8463 (N_8463,N_7877,N_7089);
nand U8464 (N_8464,N_7285,N_7948);
nor U8465 (N_8465,N_7633,N_7301);
nand U8466 (N_8466,N_7861,N_7716);
and U8467 (N_8467,N_7270,N_7989);
or U8468 (N_8468,N_7770,N_7450);
nor U8469 (N_8469,N_7400,N_7183);
nor U8470 (N_8470,N_7841,N_7589);
and U8471 (N_8471,N_7281,N_7350);
nor U8472 (N_8472,N_7386,N_7696);
and U8473 (N_8473,N_7188,N_7107);
and U8474 (N_8474,N_7239,N_7567);
xor U8475 (N_8475,N_7082,N_7308);
and U8476 (N_8476,N_7492,N_7372);
nor U8477 (N_8477,N_7467,N_7304);
and U8478 (N_8478,N_7767,N_7326);
or U8479 (N_8479,N_7846,N_7943);
or U8480 (N_8480,N_7942,N_7797);
nor U8481 (N_8481,N_7587,N_7206);
and U8482 (N_8482,N_7577,N_7017);
nand U8483 (N_8483,N_7134,N_7466);
nand U8484 (N_8484,N_7808,N_7862);
nor U8485 (N_8485,N_7609,N_7207);
or U8486 (N_8486,N_7382,N_7426);
nor U8487 (N_8487,N_7122,N_7682);
or U8488 (N_8488,N_7940,N_7184);
nand U8489 (N_8489,N_7423,N_7733);
nand U8490 (N_8490,N_7264,N_7585);
nand U8491 (N_8491,N_7526,N_7374);
and U8492 (N_8492,N_7929,N_7789);
nor U8493 (N_8493,N_7879,N_7744);
xnor U8494 (N_8494,N_7680,N_7143);
nand U8495 (N_8495,N_7705,N_7827);
and U8496 (N_8496,N_7828,N_7626);
or U8497 (N_8497,N_7409,N_7826);
or U8498 (N_8498,N_7975,N_7529);
nand U8499 (N_8499,N_7611,N_7189);
or U8500 (N_8500,N_7203,N_7056);
or U8501 (N_8501,N_7315,N_7580);
nand U8502 (N_8502,N_7122,N_7698);
nand U8503 (N_8503,N_7071,N_7364);
and U8504 (N_8504,N_7441,N_7620);
nand U8505 (N_8505,N_7097,N_7376);
and U8506 (N_8506,N_7682,N_7226);
and U8507 (N_8507,N_7757,N_7772);
or U8508 (N_8508,N_7761,N_7841);
nand U8509 (N_8509,N_7306,N_7763);
or U8510 (N_8510,N_7389,N_7319);
and U8511 (N_8511,N_7445,N_7323);
or U8512 (N_8512,N_7631,N_7778);
nand U8513 (N_8513,N_7384,N_7978);
nor U8514 (N_8514,N_7697,N_7797);
nor U8515 (N_8515,N_7821,N_7205);
nor U8516 (N_8516,N_7282,N_7622);
and U8517 (N_8517,N_7247,N_7501);
and U8518 (N_8518,N_7590,N_7938);
nand U8519 (N_8519,N_7305,N_7827);
or U8520 (N_8520,N_7772,N_7204);
nand U8521 (N_8521,N_7245,N_7675);
nand U8522 (N_8522,N_7687,N_7913);
and U8523 (N_8523,N_7732,N_7595);
or U8524 (N_8524,N_7074,N_7775);
xor U8525 (N_8525,N_7597,N_7281);
xor U8526 (N_8526,N_7790,N_7135);
nand U8527 (N_8527,N_7037,N_7887);
or U8528 (N_8528,N_7425,N_7721);
nand U8529 (N_8529,N_7594,N_7219);
or U8530 (N_8530,N_7639,N_7380);
or U8531 (N_8531,N_7283,N_7510);
and U8532 (N_8532,N_7786,N_7037);
nor U8533 (N_8533,N_7926,N_7804);
and U8534 (N_8534,N_7545,N_7723);
xor U8535 (N_8535,N_7797,N_7936);
or U8536 (N_8536,N_7980,N_7438);
and U8537 (N_8537,N_7478,N_7810);
or U8538 (N_8538,N_7552,N_7390);
or U8539 (N_8539,N_7768,N_7995);
nand U8540 (N_8540,N_7046,N_7426);
or U8541 (N_8541,N_7051,N_7411);
and U8542 (N_8542,N_7401,N_7100);
and U8543 (N_8543,N_7245,N_7429);
nand U8544 (N_8544,N_7931,N_7613);
nand U8545 (N_8545,N_7917,N_7007);
and U8546 (N_8546,N_7150,N_7628);
nor U8547 (N_8547,N_7601,N_7983);
nor U8548 (N_8548,N_7677,N_7629);
and U8549 (N_8549,N_7766,N_7784);
nand U8550 (N_8550,N_7814,N_7238);
and U8551 (N_8551,N_7376,N_7326);
and U8552 (N_8552,N_7185,N_7318);
or U8553 (N_8553,N_7821,N_7859);
nand U8554 (N_8554,N_7827,N_7140);
or U8555 (N_8555,N_7279,N_7830);
and U8556 (N_8556,N_7198,N_7965);
and U8557 (N_8557,N_7326,N_7365);
or U8558 (N_8558,N_7493,N_7355);
and U8559 (N_8559,N_7954,N_7040);
xor U8560 (N_8560,N_7732,N_7138);
and U8561 (N_8561,N_7938,N_7783);
and U8562 (N_8562,N_7191,N_7940);
and U8563 (N_8563,N_7563,N_7268);
nand U8564 (N_8564,N_7813,N_7581);
nor U8565 (N_8565,N_7316,N_7344);
nand U8566 (N_8566,N_7132,N_7018);
and U8567 (N_8567,N_7797,N_7103);
nor U8568 (N_8568,N_7714,N_7231);
and U8569 (N_8569,N_7310,N_7083);
or U8570 (N_8570,N_7022,N_7216);
or U8571 (N_8571,N_7552,N_7530);
nand U8572 (N_8572,N_7376,N_7123);
and U8573 (N_8573,N_7092,N_7333);
and U8574 (N_8574,N_7343,N_7231);
and U8575 (N_8575,N_7653,N_7626);
nor U8576 (N_8576,N_7992,N_7058);
nand U8577 (N_8577,N_7962,N_7139);
and U8578 (N_8578,N_7313,N_7782);
nand U8579 (N_8579,N_7872,N_7064);
or U8580 (N_8580,N_7947,N_7065);
xor U8581 (N_8581,N_7226,N_7653);
nand U8582 (N_8582,N_7291,N_7840);
and U8583 (N_8583,N_7874,N_7484);
or U8584 (N_8584,N_7720,N_7773);
xor U8585 (N_8585,N_7149,N_7490);
nand U8586 (N_8586,N_7388,N_7745);
and U8587 (N_8587,N_7301,N_7367);
or U8588 (N_8588,N_7575,N_7290);
or U8589 (N_8589,N_7484,N_7518);
or U8590 (N_8590,N_7468,N_7778);
or U8591 (N_8591,N_7693,N_7757);
nor U8592 (N_8592,N_7491,N_7371);
and U8593 (N_8593,N_7291,N_7480);
or U8594 (N_8594,N_7766,N_7867);
nor U8595 (N_8595,N_7272,N_7961);
nor U8596 (N_8596,N_7146,N_7160);
or U8597 (N_8597,N_7878,N_7107);
nor U8598 (N_8598,N_7014,N_7004);
nor U8599 (N_8599,N_7801,N_7714);
nand U8600 (N_8600,N_7060,N_7197);
and U8601 (N_8601,N_7941,N_7676);
nor U8602 (N_8602,N_7180,N_7874);
xnor U8603 (N_8603,N_7237,N_7590);
nor U8604 (N_8604,N_7628,N_7328);
nand U8605 (N_8605,N_7715,N_7588);
or U8606 (N_8606,N_7375,N_7810);
or U8607 (N_8607,N_7410,N_7975);
nand U8608 (N_8608,N_7084,N_7872);
and U8609 (N_8609,N_7171,N_7493);
nor U8610 (N_8610,N_7434,N_7509);
xor U8611 (N_8611,N_7796,N_7069);
nor U8612 (N_8612,N_7666,N_7516);
and U8613 (N_8613,N_7507,N_7403);
or U8614 (N_8614,N_7823,N_7643);
nor U8615 (N_8615,N_7158,N_7762);
nand U8616 (N_8616,N_7764,N_7553);
or U8617 (N_8617,N_7572,N_7157);
nor U8618 (N_8618,N_7586,N_7699);
nand U8619 (N_8619,N_7276,N_7164);
xor U8620 (N_8620,N_7321,N_7528);
xnor U8621 (N_8621,N_7069,N_7344);
nand U8622 (N_8622,N_7944,N_7046);
nor U8623 (N_8623,N_7879,N_7966);
nand U8624 (N_8624,N_7860,N_7695);
and U8625 (N_8625,N_7379,N_7879);
nor U8626 (N_8626,N_7260,N_7621);
and U8627 (N_8627,N_7797,N_7826);
nand U8628 (N_8628,N_7346,N_7143);
or U8629 (N_8629,N_7321,N_7044);
nand U8630 (N_8630,N_7709,N_7022);
nand U8631 (N_8631,N_7472,N_7463);
or U8632 (N_8632,N_7383,N_7205);
and U8633 (N_8633,N_7850,N_7601);
and U8634 (N_8634,N_7005,N_7462);
nor U8635 (N_8635,N_7449,N_7072);
or U8636 (N_8636,N_7794,N_7855);
nor U8637 (N_8637,N_7576,N_7723);
and U8638 (N_8638,N_7640,N_7879);
nand U8639 (N_8639,N_7968,N_7420);
nand U8640 (N_8640,N_7207,N_7645);
or U8641 (N_8641,N_7473,N_7965);
nor U8642 (N_8642,N_7158,N_7029);
nand U8643 (N_8643,N_7975,N_7392);
or U8644 (N_8644,N_7754,N_7562);
or U8645 (N_8645,N_7460,N_7705);
nand U8646 (N_8646,N_7357,N_7092);
nand U8647 (N_8647,N_7123,N_7922);
nand U8648 (N_8648,N_7296,N_7793);
nand U8649 (N_8649,N_7361,N_7432);
or U8650 (N_8650,N_7776,N_7427);
nor U8651 (N_8651,N_7707,N_7560);
nand U8652 (N_8652,N_7082,N_7800);
xor U8653 (N_8653,N_7347,N_7328);
and U8654 (N_8654,N_7423,N_7863);
or U8655 (N_8655,N_7090,N_7561);
and U8656 (N_8656,N_7234,N_7549);
or U8657 (N_8657,N_7282,N_7051);
or U8658 (N_8658,N_7277,N_7305);
nor U8659 (N_8659,N_7767,N_7583);
or U8660 (N_8660,N_7017,N_7040);
or U8661 (N_8661,N_7201,N_7573);
nand U8662 (N_8662,N_7473,N_7219);
nor U8663 (N_8663,N_7941,N_7158);
and U8664 (N_8664,N_7742,N_7706);
nor U8665 (N_8665,N_7781,N_7386);
and U8666 (N_8666,N_7719,N_7482);
and U8667 (N_8667,N_7574,N_7421);
nor U8668 (N_8668,N_7709,N_7854);
nor U8669 (N_8669,N_7108,N_7746);
nor U8670 (N_8670,N_7555,N_7086);
nand U8671 (N_8671,N_7291,N_7500);
nand U8672 (N_8672,N_7708,N_7011);
nor U8673 (N_8673,N_7194,N_7432);
nor U8674 (N_8674,N_7179,N_7874);
or U8675 (N_8675,N_7205,N_7464);
nor U8676 (N_8676,N_7551,N_7261);
nand U8677 (N_8677,N_7536,N_7127);
or U8678 (N_8678,N_7577,N_7357);
and U8679 (N_8679,N_7884,N_7316);
or U8680 (N_8680,N_7592,N_7128);
nor U8681 (N_8681,N_7468,N_7400);
nor U8682 (N_8682,N_7027,N_7877);
xor U8683 (N_8683,N_7329,N_7078);
nor U8684 (N_8684,N_7001,N_7492);
or U8685 (N_8685,N_7493,N_7695);
or U8686 (N_8686,N_7543,N_7552);
and U8687 (N_8687,N_7386,N_7788);
and U8688 (N_8688,N_7729,N_7338);
or U8689 (N_8689,N_7270,N_7633);
and U8690 (N_8690,N_7503,N_7723);
or U8691 (N_8691,N_7428,N_7900);
and U8692 (N_8692,N_7119,N_7583);
nor U8693 (N_8693,N_7750,N_7788);
nor U8694 (N_8694,N_7686,N_7023);
or U8695 (N_8695,N_7875,N_7323);
and U8696 (N_8696,N_7269,N_7683);
and U8697 (N_8697,N_7592,N_7032);
nor U8698 (N_8698,N_7337,N_7995);
nand U8699 (N_8699,N_7681,N_7608);
or U8700 (N_8700,N_7462,N_7782);
and U8701 (N_8701,N_7862,N_7782);
or U8702 (N_8702,N_7306,N_7180);
nor U8703 (N_8703,N_7949,N_7226);
nor U8704 (N_8704,N_7179,N_7249);
nor U8705 (N_8705,N_7624,N_7605);
or U8706 (N_8706,N_7036,N_7717);
nor U8707 (N_8707,N_7576,N_7165);
nor U8708 (N_8708,N_7289,N_7284);
or U8709 (N_8709,N_7307,N_7734);
nor U8710 (N_8710,N_7193,N_7212);
nor U8711 (N_8711,N_7233,N_7389);
and U8712 (N_8712,N_7543,N_7492);
and U8713 (N_8713,N_7226,N_7194);
xor U8714 (N_8714,N_7642,N_7030);
nor U8715 (N_8715,N_7743,N_7592);
nor U8716 (N_8716,N_7346,N_7960);
nor U8717 (N_8717,N_7792,N_7213);
and U8718 (N_8718,N_7773,N_7525);
nand U8719 (N_8719,N_7026,N_7639);
xor U8720 (N_8720,N_7194,N_7451);
and U8721 (N_8721,N_7063,N_7993);
or U8722 (N_8722,N_7529,N_7310);
nor U8723 (N_8723,N_7347,N_7553);
nor U8724 (N_8724,N_7955,N_7305);
nor U8725 (N_8725,N_7054,N_7942);
nand U8726 (N_8726,N_7261,N_7397);
nand U8727 (N_8727,N_7131,N_7267);
and U8728 (N_8728,N_7579,N_7565);
nor U8729 (N_8729,N_7673,N_7630);
or U8730 (N_8730,N_7617,N_7774);
nand U8731 (N_8731,N_7131,N_7165);
or U8732 (N_8732,N_7574,N_7625);
nand U8733 (N_8733,N_7597,N_7851);
nand U8734 (N_8734,N_7030,N_7638);
nand U8735 (N_8735,N_7698,N_7714);
nor U8736 (N_8736,N_7281,N_7321);
and U8737 (N_8737,N_7256,N_7188);
nor U8738 (N_8738,N_7858,N_7130);
and U8739 (N_8739,N_7244,N_7329);
nand U8740 (N_8740,N_7685,N_7150);
and U8741 (N_8741,N_7853,N_7351);
or U8742 (N_8742,N_7185,N_7594);
and U8743 (N_8743,N_7307,N_7851);
and U8744 (N_8744,N_7792,N_7616);
nand U8745 (N_8745,N_7907,N_7182);
or U8746 (N_8746,N_7158,N_7234);
and U8747 (N_8747,N_7056,N_7312);
nor U8748 (N_8748,N_7614,N_7701);
or U8749 (N_8749,N_7050,N_7766);
nand U8750 (N_8750,N_7942,N_7636);
and U8751 (N_8751,N_7311,N_7258);
nor U8752 (N_8752,N_7125,N_7773);
nor U8753 (N_8753,N_7227,N_7390);
and U8754 (N_8754,N_7274,N_7457);
nor U8755 (N_8755,N_7435,N_7893);
nand U8756 (N_8756,N_7184,N_7125);
or U8757 (N_8757,N_7618,N_7036);
xor U8758 (N_8758,N_7556,N_7115);
or U8759 (N_8759,N_7822,N_7861);
and U8760 (N_8760,N_7642,N_7702);
nor U8761 (N_8761,N_7133,N_7610);
nand U8762 (N_8762,N_7240,N_7813);
nand U8763 (N_8763,N_7883,N_7488);
and U8764 (N_8764,N_7266,N_7228);
or U8765 (N_8765,N_7907,N_7005);
xnor U8766 (N_8766,N_7523,N_7953);
and U8767 (N_8767,N_7501,N_7407);
and U8768 (N_8768,N_7406,N_7589);
or U8769 (N_8769,N_7444,N_7627);
or U8770 (N_8770,N_7534,N_7985);
and U8771 (N_8771,N_7004,N_7305);
and U8772 (N_8772,N_7581,N_7492);
nor U8773 (N_8773,N_7935,N_7589);
and U8774 (N_8774,N_7238,N_7524);
or U8775 (N_8775,N_7869,N_7264);
nor U8776 (N_8776,N_7061,N_7790);
and U8777 (N_8777,N_7551,N_7058);
nor U8778 (N_8778,N_7633,N_7494);
and U8779 (N_8779,N_7295,N_7165);
nor U8780 (N_8780,N_7772,N_7537);
nand U8781 (N_8781,N_7524,N_7984);
or U8782 (N_8782,N_7726,N_7917);
and U8783 (N_8783,N_7633,N_7074);
and U8784 (N_8784,N_7106,N_7267);
nand U8785 (N_8785,N_7045,N_7266);
or U8786 (N_8786,N_7363,N_7914);
or U8787 (N_8787,N_7868,N_7874);
or U8788 (N_8788,N_7193,N_7651);
nor U8789 (N_8789,N_7755,N_7624);
nor U8790 (N_8790,N_7473,N_7316);
nand U8791 (N_8791,N_7429,N_7903);
or U8792 (N_8792,N_7172,N_7523);
and U8793 (N_8793,N_7854,N_7607);
or U8794 (N_8794,N_7602,N_7104);
nor U8795 (N_8795,N_7254,N_7033);
and U8796 (N_8796,N_7838,N_7307);
or U8797 (N_8797,N_7227,N_7774);
nand U8798 (N_8798,N_7712,N_7558);
nor U8799 (N_8799,N_7179,N_7370);
nor U8800 (N_8800,N_7606,N_7251);
or U8801 (N_8801,N_7118,N_7561);
and U8802 (N_8802,N_7073,N_7395);
nand U8803 (N_8803,N_7463,N_7071);
and U8804 (N_8804,N_7045,N_7940);
nand U8805 (N_8805,N_7307,N_7310);
nand U8806 (N_8806,N_7542,N_7584);
nor U8807 (N_8807,N_7483,N_7024);
nand U8808 (N_8808,N_7609,N_7581);
and U8809 (N_8809,N_7456,N_7244);
or U8810 (N_8810,N_7131,N_7971);
xnor U8811 (N_8811,N_7651,N_7882);
or U8812 (N_8812,N_7911,N_7678);
nor U8813 (N_8813,N_7652,N_7596);
or U8814 (N_8814,N_7704,N_7964);
or U8815 (N_8815,N_7206,N_7571);
or U8816 (N_8816,N_7660,N_7515);
nand U8817 (N_8817,N_7956,N_7794);
and U8818 (N_8818,N_7454,N_7339);
nand U8819 (N_8819,N_7291,N_7509);
and U8820 (N_8820,N_7473,N_7955);
nand U8821 (N_8821,N_7102,N_7022);
nand U8822 (N_8822,N_7727,N_7667);
and U8823 (N_8823,N_7251,N_7539);
or U8824 (N_8824,N_7192,N_7235);
nor U8825 (N_8825,N_7763,N_7898);
xor U8826 (N_8826,N_7135,N_7563);
nor U8827 (N_8827,N_7892,N_7442);
and U8828 (N_8828,N_7209,N_7219);
nand U8829 (N_8829,N_7261,N_7505);
or U8830 (N_8830,N_7542,N_7708);
nand U8831 (N_8831,N_7252,N_7608);
or U8832 (N_8832,N_7884,N_7666);
or U8833 (N_8833,N_7687,N_7389);
or U8834 (N_8834,N_7567,N_7967);
nand U8835 (N_8835,N_7871,N_7951);
or U8836 (N_8836,N_7201,N_7048);
or U8837 (N_8837,N_7186,N_7572);
and U8838 (N_8838,N_7935,N_7455);
or U8839 (N_8839,N_7630,N_7236);
nor U8840 (N_8840,N_7652,N_7210);
or U8841 (N_8841,N_7089,N_7976);
or U8842 (N_8842,N_7783,N_7522);
nand U8843 (N_8843,N_7122,N_7243);
and U8844 (N_8844,N_7032,N_7974);
or U8845 (N_8845,N_7708,N_7044);
or U8846 (N_8846,N_7232,N_7649);
or U8847 (N_8847,N_7508,N_7479);
nand U8848 (N_8848,N_7546,N_7217);
or U8849 (N_8849,N_7381,N_7141);
nor U8850 (N_8850,N_7191,N_7994);
nor U8851 (N_8851,N_7701,N_7593);
nand U8852 (N_8852,N_7514,N_7094);
nand U8853 (N_8853,N_7556,N_7431);
nor U8854 (N_8854,N_7810,N_7942);
and U8855 (N_8855,N_7670,N_7229);
nor U8856 (N_8856,N_7768,N_7843);
or U8857 (N_8857,N_7279,N_7933);
or U8858 (N_8858,N_7031,N_7736);
and U8859 (N_8859,N_7964,N_7432);
and U8860 (N_8860,N_7455,N_7964);
nor U8861 (N_8861,N_7658,N_7889);
nor U8862 (N_8862,N_7729,N_7127);
and U8863 (N_8863,N_7736,N_7910);
nor U8864 (N_8864,N_7150,N_7545);
nor U8865 (N_8865,N_7344,N_7867);
and U8866 (N_8866,N_7741,N_7972);
nand U8867 (N_8867,N_7424,N_7940);
nand U8868 (N_8868,N_7233,N_7522);
nand U8869 (N_8869,N_7614,N_7374);
and U8870 (N_8870,N_7216,N_7263);
and U8871 (N_8871,N_7380,N_7660);
and U8872 (N_8872,N_7531,N_7707);
nand U8873 (N_8873,N_7662,N_7981);
and U8874 (N_8874,N_7686,N_7338);
or U8875 (N_8875,N_7067,N_7364);
nor U8876 (N_8876,N_7096,N_7393);
or U8877 (N_8877,N_7476,N_7997);
or U8878 (N_8878,N_7065,N_7685);
and U8879 (N_8879,N_7924,N_7215);
nand U8880 (N_8880,N_7810,N_7861);
nor U8881 (N_8881,N_7889,N_7820);
nor U8882 (N_8882,N_7345,N_7811);
or U8883 (N_8883,N_7923,N_7431);
or U8884 (N_8884,N_7102,N_7489);
and U8885 (N_8885,N_7113,N_7199);
or U8886 (N_8886,N_7849,N_7218);
nor U8887 (N_8887,N_7997,N_7361);
nand U8888 (N_8888,N_7340,N_7376);
and U8889 (N_8889,N_7129,N_7304);
or U8890 (N_8890,N_7134,N_7902);
and U8891 (N_8891,N_7317,N_7231);
and U8892 (N_8892,N_7012,N_7120);
and U8893 (N_8893,N_7049,N_7197);
or U8894 (N_8894,N_7009,N_7783);
or U8895 (N_8895,N_7020,N_7007);
and U8896 (N_8896,N_7401,N_7262);
and U8897 (N_8897,N_7292,N_7498);
and U8898 (N_8898,N_7242,N_7094);
nand U8899 (N_8899,N_7752,N_7042);
nand U8900 (N_8900,N_7259,N_7417);
nor U8901 (N_8901,N_7962,N_7038);
or U8902 (N_8902,N_7024,N_7699);
or U8903 (N_8903,N_7286,N_7622);
or U8904 (N_8904,N_7829,N_7813);
nor U8905 (N_8905,N_7687,N_7404);
or U8906 (N_8906,N_7118,N_7901);
nand U8907 (N_8907,N_7615,N_7946);
nand U8908 (N_8908,N_7065,N_7568);
nor U8909 (N_8909,N_7622,N_7911);
nor U8910 (N_8910,N_7482,N_7530);
or U8911 (N_8911,N_7906,N_7451);
nor U8912 (N_8912,N_7284,N_7330);
nor U8913 (N_8913,N_7677,N_7892);
xnor U8914 (N_8914,N_7878,N_7354);
nand U8915 (N_8915,N_7761,N_7681);
nor U8916 (N_8916,N_7763,N_7794);
nand U8917 (N_8917,N_7425,N_7202);
and U8918 (N_8918,N_7652,N_7283);
nor U8919 (N_8919,N_7711,N_7342);
and U8920 (N_8920,N_7364,N_7665);
and U8921 (N_8921,N_7201,N_7355);
nor U8922 (N_8922,N_7129,N_7496);
nand U8923 (N_8923,N_7221,N_7360);
nor U8924 (N_8924,N_7874,N_7447);
xnor U8925 (N_8925,N_7712,N_7907);
or U8926 (N_8926,N_7403,N_7007);
or U8927 (N_8927,N_7938,N_7690);
and U8928 (N_8928,N_7555,N_7432);
nand U8929 (N_8929,N_7476,N_7764);
nor U8930 (N_8930,N_7172,N_7882);
nand U8931 (N_8931,N_7640,N_7716);
nand U8932 (N_8932,N_7999,N_7519);
nand U8933 (N_8933,N_7498,N_7269);
nand U8934 (N_8934,N_7130,N_7398);
xnor U8935 (N_8935,N_7381,N_7662);
or U8936 (N_8936,N_7944,N_7383);
or U8937 (N_8937,N_7961,N_7557);
nand U8938 (N_8938,N_7790,N_7164);
nor U8939 (N_8939,N_7084,N_7394);
nand U8940 (N_8940,N_7749,N_7785);
and U8941 (N_8941,N_7136,N_7516);
or U8942 (N_8942,N_7598,N_7575);
and U8943 (N_8943,N_7820,N_7139);
or U8944 (N_8944,N_7968,N_7767);
nor U8945 (N_8945,N_7927,N_7043);
xor U8946 (N_8946,N_7269,N_7697);
or U8947 (N_8947,N_7418,N_7883);
nand U8948 (N_8948,N_7279,N_7242);
nor U8949 (N_8949,N_7943,N_7049);
nand U8950 (N_8950,N_7318,N_7495);
nand U8951 (N_8951,N_7776,N_7510);
or U8952 (N_8952,N_7959,N_7181);
nor U8953 (N_8953,N_7347,N_7709);
nand U8954 (N_8954,N_7039,N_7866);
and U8955 (N_8955,N_7233,N_7703);
or U8956 (N_8956,N_7719,N_7656);
nor U8957 (N_8957,N_7873,N_7179);
and U8958 (N_8958,N_7750,N_7426);
and U8959 (N_8959,N_7969,N_7594);
xnor U8960 (N_8960,N_7583,N_7800);
or U8961 (N_8961,N_7449,N_7195);
and U8962 (N_8962,N_7779,N_7321);
and U8963 (N_8963,N_7147,N_7198);
and U8964 (N_8964,N_7836,N_7154);
or U8965 (N_8965,N_7550,N_7317);
nand U8966 (N_8966,N_7342,N_7709);
or U8967 (N_8967,N_7991,N_7646);
or U8968 (N_8968,N_7098,N_7651);
or U8969 (N_8969,N_7919,N_7219);
nor U8970 (N_8970,N_7108,N_7851);
and U8971 (N_8971,N_7175,N_7602);
nor U8972 (N_8972,N_7711,N_7883);
xor U8973 (N_8973,N_7328,N_7870);
and U8974 (N_8974,N_7283,N_7981);
or U8975 (N_8975,N_7556,N_7101);
nand U8976 (N_8976,N_7991,N_7319);
and U8977 (N_8977,N_7002,N_7610);
and U8978 (N_8978,N_7101,N_7403);
nand U8979 (N_8979,N_7838,N_7160);
or U8980 (N_8980,N_7339,N_7784);
and U8981 (N_8981,N_7055,N_7400);
nor U8982 (N_8982,N_7962,N_7421);
nand U8983 (N_8983,N_7403,N_7662);
or U8984 (N_8984,N_7177,N_7347);
nand U8985 (N_8985,N_7640,N_7625);
or U8986 (N_8986,N_7512,N_7363);
and U8987 (N_8987,N_7260,N_7011);
nor U8988 (N_8988,N_7286,N_7306);
or U8989 (N_8989,N_7904,N_7640);
nand U8990 (N_8990,N_7863,N_7271);
nand U8991 (N_8991,N_7863,N_7035);
and U8992 (N_8992,N_7303,N_7612);
or U8993 (N_8993,N_7893,N_7367);
and U8994 (N_8994,N_7447,N_7743);
xnor U8995 (N_8995,N_7285,N_7951);
nand U8996 (N_8996,N_7547,N_7266);
and U8997 (N_8997,N_7331,N_7762);
and U8998 (N_8998,N_7790,N_7170);
and U8999 (N_8999,N_7628,N_7871);
and U9000 (N_9000,N_8496,N_8899);
and U9001 (N_9001,N_8345,N_8070);
nor U9002 (N_9002,N_8926,N_8501);
or U9003 (N_9003,N_8124,N_8554);
nor U9004 (N_9004,N_8118,N_8651);
and U9005 (N_9005,N_8234,N_8869);
nand U9006 (N_9006,N_8789,N_8941);
and U9007 (N_9007,N_8109,N_8062);
nor U9008 (N_9008,N_8037,N_8671);
and U9009 (N_9009,N_8590,N_8003);
or U9010 (N_9010,N_8721,N_8014);
xor U9011 (N_9011,N_8279,N_8361);
or U9012 (N_9012,N_8558,N_8967);
nor U9013 (N_9013,N_8173,N_8143);
or U9014 (N_9014,N_8659,N_8834);
and U9015 (N_9015,N_8809,N_8565);
nor U9016 (N_9016,N_8597,N_8186);
or U9017 (N_9017,N_8050,N_8807);
or U9018 (N_9018,N_8678,N_8910);
nor U9019 (N_9019,N_8581,N_8564);
and U9020 (N_9020,N_8650,N_8931);
nor U9021 (N_9021,N_8170,N_8171);
nor U9022 (N_9022,N_8935,N_8540);
or U9023 (N_9023,N_8606,N_8850);
nand U9024 (N_9024,N_8624,N_8356);
nor U9025 (N_9025,N_8432,N_8242);
and U9026 (N_9026,N_8491,N_8623);
and U9027 (N_9027,N_8755,N_8669);
nor U9028 (N_9028,N_8603,N_8896);
or U9029 (N_9029,N_8589,N_8131);
nand U9030 (N_9030,N_8828,N_8878);
nand U9031 (N_9031,N_8113,N_8660);
nand U9032 (N_9032,N_8007,N_8567);
nor U9033 (N_9033,N_8505,N_8368);
nor U9034 (N_9034,N_8796,N_8295);
or U9035 (N_9035,N_8736,N_8183);
or U9036 (N_9036,N_8788,N_8398);
and U9037 (N_9037,N_8212,N_8914);
nand U9038 (N_9038,N_8031,N_8381);
nor U9039 (N_9039,N_8853,N_8805);
nor U9040 (N_9040,N_8304,N_8799);
and U9041 (N_9041,N_8535,N_8060);
nand U9042 (N_9042,N_8400,N_8619);
nand U9043 (N_9043,N_8702,N_8605);
xnor U9044 (N_9044,N_8919,N_8323);
nand U9045 (N_9045,N_8785,N_8239);
nor U9046 (N_9046,N_8454,N_8577);
nor U9047 (N_9047,N_8962,N_8808);
nor U9048 (N_9048,N_8810,N_8065);
or U9049 (N_9049,N_8579,N_8228);
or U9050 (N_9050,N_8775,N_8359);
or U9051 (N_9051,N_8078,N_8887);
and U9052 (N_9052,N_8610,N_8169);
nand U9053 (N_9053,N_8717,N_8649);
nand U9054 (N_9054,N_8916,N_8331);
and U9055 (N_9055,N_8327,N_8397);
and U9056 (N_9056,N_8248,N_8987);
or U9057 (N_9057,N_8001,N_8319);
nor U9058 (N_9058,N_8519,N_8394);
and U9059 (N_9059,N_8376,N_8436);
nor U9060 (N_9060,N_8572,N_8348);
nand U9061 (N_9061,N_8665,N_8042);
nor U9062 (N_9062,N_8451,N_8291);
and U9063 (N_9063,N_8192,N_8645);
nand U9064 (N_9064,N_8800,N_8691);
and U9065 (N_9065,N_8907,N_8393);
and U9066 (N_9066,N_8993,N_8561);
and U9067 (N_9067,N_8823,N_8602);
nand U9068 (N_9068,N_8929,N_8444);
xnor U9069 (N_9069,N_8750,N_8608);
nand U9070 (N_9070,N_8832,N_8421);
nand U9071 (N_9071,N_8483,N_8695);
nor U9072 (N_9072,N_8149,N_8842);
nor U9073 (N_9073,N_8117,N_8628);
nor U9074 (N_9074,N_8103,N_8133);
and U9075 (N_9075,N_8971,N_8321);
or U9076 (N_9076,N_8395,N_8879);
nand U9077 (N_9077,N_8954,N_8445);
and U9078 (N_9078,N_8865,N_8229);
or U9079 (N_9079,N_8245,N_8043);
nand U9080 (N_9080,N_8293,N_8284);
and U9081 (N_9081,N_8989,N_8417);
nor U9082 (N_9082,N_8674,N_8246);
nor U9083 (N_9083,N_8144,N_8515);
xnor U9084 (N_9084,N_8071,N_8763);
or U9085 (N_9085,N_8240,N_8197);
and U9086 (N_9086,N_8227,N_8613);
nand U9087 (N_9087,N_8487,N_8803);
nor U9088 (N_9088,N_8885,N_8034);
nor U9089 (N_9089,N_8604,N_8438);
or U9090 (N_9090,N_8254,N_8326);
or U9091 (N_9091,N_8902,N_8922);
and U9092 (N_9092,N_8854,N_8531);
and U9093 (N_9093,N_8302,N_8666);
nand U9094 (N_9094,N_8614,N_8375);
nor U9095 (N_9095,N_8708,N_8662);
nor U9096 (N_9096,N_8325,N_8524);
nand U9097 (N_9097,N_8725,N_8758);
nor U9098 (N_9098,N_8706,N_8575);
nand U9099 (N_9099,N_8867,N_8046);
xor U9100 (N_9100,N_8313,N_8092);
or U9101 (N_9101,N_8968,N_8029);
and U9102 (N_9102,N_8748,N_8988);
nor U9103 (N_9103,N_8960,N_8557);
nand U9104 (N_9104,N_8292,N_8693);
nor U9105 (N_9105,N_8928,N_8396);
nand U9106 (N_9106,N_8670,N_8985);
and U9107 (N_9107,N_8038,N_8735);
and U9108 (N_9108,N_8679,N_8108);
nand U9109 (N_9109,N_8552,N_8656);
or U9110 (N_9110,N_8517,N_8159);
nor U9111 (N_9111,N_8544,N_8860);
nand U9112 (N_9112,N_8664,N_8714);
nor U9113 (N_9113,N_8508,N_8819);
nand U9114 (N_9114,N_8719,N_8209);
or U9115 (N_9115,N_8891,N_8536);
nor U9116 (N_9116,N_8430,N_8844);
or U9117 (N_9117,N_8354,N_8503);
or U9118 (N_9118,N_8526,N_8045);
nand U9119 (N_9119,N_8482,N_8843);
or U9120 (N_9120,N_8626,N_8768);
nor U9121 (N_9121,N_8587,N_8801);
nor U9122 (N_9122,N_8551,N_8663);
nand U9123 (N_9123,N_8120,N_8868);
or U9124 (N_9124,N_8855,N_8465);
and U9125 (N_9125,N_8792,N_8163);
or U9126 (N_9126,N_8213,N_8897);
nor U9127 (N_9127,N_8274,N_8371);
nand U9128 (N_9128,N_8407,N_8739);
nor U9129 (N_9129,N_8779,N_8439);
and U9130 (N_9130,N_8514,N_8222);
and U9131 (N_9131,N_8179,N_8731);
xnor U9132 (N_9132,N_8235,N_8635);
nand U9133 (N_9133,N_8250,N_8214);
nand U9134 (N_9134,N_8265,N_8399);
nand U9135 (N_9135,N_8106,N_8220);
nand U9136 (N_9136,N_8329,N_8181);
nor U9137 (N_9137,N_8692,N_8475);
nand U9138 (N_9138,N_8629,N_8986);
nor U9139 (N_9139,N_8294,N_8688);
nor U9140 (N_9140,N_8324,N_8090);
and U9141 (N_9141,N_8104,N_8364);
or U9142 (N_9142,N_8949,N_8538);
nor U9143 (N_9143,N_8009,N_8727);
or U9144 (N_9144,N_8711,N_8480);
nand U9145 (N_9145,N_8370,N_8571);
or U9146 (N_9146,N_8894,N_8028);
or U9147 (N_9147,N_8848,N_8252);
xnor U9148 (N_9148,N_8724,N_8172);
nand U9149 (N_9149,N_8094,N_8040);
nor U9150 (N_9150,N_8115,N_8264);
and U9151 (N_9151,N_8908,N_8784);
and U9152 (N_9152,N_8906,N_8917);
xnor U9153 (N_9153,N_8733,N_8580);
nand U9154 (N_9154,N_8699,N_8957);
and U9155 (N_9155,N_8460,N_8548);
nand U9156 (N_9156,N_8521,N_8940);
nor U9157 (N_9157,N_8138,N_8905);
nor U9158 (N_9158,N_8627,N_8648);
or U9159 (N_9159,N_8886,N_8365);
and U9160 (N_9160,N_8208,N_8328);
or U9161 (N_9161,N_8225,N_8497);
nor U9162 (N_9162,N_8995,N_8041);
nand U9163 (N_9163,N_8336,N_8523);
or U9164 (N_9164,N_8632,N_8201);
and U9165 (N_9165,N_8574,N_8925);
or U9166 (N_9166,N_8273,N_8435);
nor U9167 (N_9167,N_8509,N_8493);
or U9168 (N_9168,N_8573,N_8039);
nand U9169 (N_9169,N_8205,N_8990);
nand U9170 (N_9170,N_8114,N_8713);
nand U9171 (N_9171,N_8697,N_8424);
and U9172 (N_9172,N_8760,N_8369);
nand U9173 (N_9173,N_8765,N_8271);
nand U9174 (N_9174,N_8742,N_8654);
nor U9175 (N_9175,N_8099,N_8857);
and U9176 (N_9176,N_8952,N_8403);
nor U9177 (N_9177,N_8450,N_8944);
nor U9178 (N_9178,N_8927,N_8513);
and U9179 (N_9179,N_8686,N_8522);
nand U9180 (N_9180,N_8948,N_8311);
nor U9181 (N_9181,N_8024,N_8193);
and U9182 (N_9182,N_8787,N_8640);
nor U9183 (N_9183,N_8226,N_8932);
or U9184 (N_9184,N_8056,N_8478);
nand U9185 (N_9185,N_8261,N_8794);
nand U9186 (N_9186,N_8730,N_8119);
nand U9187 (N_9187,N_8915,N_8741);
and U9188 (N_9188,N_8020,N_8342);
nand U9189 (N_9189,N_8266,N_8840);
and U9190 (N_9190,N_8655,N_8738);
and U9191 (N_9191,N_8017,N_8647);
xnor U9192 (N_9192,N_8428,N_8077);
or U9193 (N_9193,N_8946,N_8959);
or U9194 (N_9194,N_8998,N_8105);
nor U9195 (N_9195,N_8055,N_8392);
nand U9196 (N_9196,N_8155,N_8303);
nand U9197 (N_9197,N_8539,N_8140);
and U9198 (N_9198,N_8937,N_8633);
xnor U9199 (N_9199,N_8534,N_8873);
and U9200 (N_9200,N_8773,N_8463);
and U9201 (N_9201,N_8086,N_8797);
nand U9202 (N_9202,N_8530,N_8468);
and U9203 (N_9203,N_8756,N_8901);
nor U9204 (N_9204,N_8723,N_8909);
nor U9205 (N_9205,N_8722,N_8685);
nor U9206 (N_9206,N_8469,N_8344);
nor U9207 (N_9207,N_8533,N_8849);
nand U9208 (N_9208,N_8484,N_8970);
and U9209 (N_9209,N_8732,N_8506);
or U9210 (N_9210,N_8746,N_8818);
nand U9211 (N_9211,N_8537,N_8161);
and U9212 (N_9212,N_8025,N_8578);
nand U9213 (N_9213,N_8776,N_8427);
or U9214 (N_9214,N_8022,N_8263);
nand U9215 (N_9215,N_8139,N_8676);
nand U9216 (N_9216,N_8459,N_8032);
nor U9217 (N_9217,N_8806,N_8991);
or U9218 (N_9218,N_8956,N_8786);
and U9219 (N_9219,N_8030,N_8821);
nand U9220 (N_9220,N_8550,N_8419);
or U9221 (N_9221,N_8426,N_8997);
nand U9222 (N_9222,N_8983,N_8595);
and U9223 (N_9223,N_8249,N_8277);
and U9224 (N_9224,N_8474,N_8203);
nand U9225 (N_9225,N_8858,N_8236);
or U9226 (N_9226,N_8027,N_8198);
or U9227 (N_9227,N_8673,N_8672);
nand U9228 (N_9228,N_8458,N_8141);
nand U9229 (N_9229,N_8500,N_8618);
and U9230 (N_9230,N_8880,N_8363);
nand U9231 (N_9231,N_8272,N_8101);
nor U9232 (N_9232,N_8076,N_8740);
or U9233 (N_9233,N_8044,N_8745);
nor U9234 (N_9234,N_8123,N_8638);
nand U9235 (N_9235,N_8390,N_8631);
nor U9236 (N_9236,N_8116,N_8188);
or U9237 (N_9237,N_8013,N_8795);
nor U9238 (N_9238,N_8620,N_8762);
and U9239 (N_9239,N_8333,N_8726);
and U9240 (N_9240,N_8838,N_8884);
nor U9241 (N_9241,N_8945,N_8667);
and U9242 (N_9242,N_8831,N_8243);
or U9243 (N_9243,N_8851,N_8529);
or U9244 (N_9244,N_8682,N_8247);
nor U9245 (N_9245,N_8033,N_8830);
and U9246 (N_9246,N_8337,N_8175);
nand U9247 (N_9247,N_8625,N_8296);
or U9248 (N_9248,N_8063,N_8021);
and U9249 (N_9249,N_8979,N_8471);
or U9250 (N_9250,N_8977,N_8507);
and U9251 (N_9251,N_8241,N_8377);
nand U9252 (N_9252,N_8846,N_8955);
and U9253 (N_9253,N_8969,N_8898);
or U9254 (N_9254,N_8476,N_8267);
nor U9255 (N_9255,N_8754,N_8704);
nor U9256 (N_9256,N_8980,N_8617);
and U9257 (N_9257,N_8637,N_8005);
or U9258 (N_9258,N_8452,N_8683);
nand U9259 (N_9259,N_8446,N_8877);
and U9260 (N_9260,N_8408,N_8048);
nor U9261 (N_9261,N_8467,N_8084);
nor U9262 (N_9262,N_8232,N_8689);
nand U9263 (N_9263,N_8130,N_8165);
or U9264 (N_9264,N_8418,N_8479);
and U9265 (N_9265,N_8639,N_8824);
and U9266 (N_9266,N_8871,N_8545);
nand U9267 (N_9267,N_8047,N_8317);
nand U9268 (N_9268,N_8135,N_8059);
nor U9269 (N_9269,N_8999,N_8449);
or U9270 (N_9270,N_8943,N_8006);
nand U9271 (N_9271,N_8401,N_8772);
nor U9272 (N_9272,N_8072,N_8315);
or U9273 (N_9273,N_8258,N_8180);
and U9274 (N_9274,N_8994,N_8134);
nor U9275 (N_9275,N_8307,N_8111);
nor U9276 (N_9276,N_8287,N_8253);
nor U9277 (N_9277,N_8751,N_8757);
nor U9278 (N_9278,N_8996,N_8498);
or U9279 (N_9279,N_8298,N_8387);
and U9280 (N_9280,N_8875,N_8528);
nand U9281 (N_9281,N_8904,N_8816);
nor U9282 (N_9282,N_8184,N_8568);
nand U9283 (N_9283,N_8716,N_8541);
nand U9284 (N_9284,N_8516,N_8251);
or U9285 (N_9285,N_8802,N_8332);
or U9286 (N_9286,N_8859,N_8856);
nor U9287 (N_9287,N_8185,N_8053);
and U9288 (N_9288,N_8622,N_8644);
and U9289 (N_9289,N_8817,N_8338);
or U9290 (N_9290,N_8367,N_8309);
or U9291 (N_9291,N_8168,N_8036);
nand U9292 (N_9292,N_8592,N_8079);
and U9293 (N_9293,N_8687,N_8352);
nand U9294 (N_9294,N_8391,N_8833);
xor U9295 (N_9295,N_8152,N_8488);
nor U9296 (N_9296,N_8729,N_8583);
and U9297 (N_9297,N_8889,N_8314);
and U9298 (N_9298,N_8698,N_8194);
nand U9299 (N_9299,N_8643,N_8494);
or U9300 (N_9300,N_8893,N_8646);
nand U9301 (N_9301,N_8798,N_8972);
nor U9302 (N_9302,N_8316,N_8431);
nor U9303 (N_9303,N_8462,N_8260);
nor U9304 (N_9304,N_8609,N_8412);
and U9305 (N_9305,N_8542,N_8189);
or U9306 (N_9306,N_8191,N_8137);
nor U9307 (N_9307,N_8978,N_8826);
nor U9308 (N_9308,N_8000,N_8362);
or U9309 (N_9309,N_8965,N_8058);
nand U9310 (N_9310,N_8154,N_8930);
and U9311 (N_9311,N_8696,N_8812);
nand U9312 (N_9312,N_8196,N_8839);
nor U9313 (N_9313,N_8011,N_8947);
nand U9314 (N_9314,N_8598,N_8268);
nor U9315 (N_9315,N_8002,N_8835);
or U9316 (N_9316,N_8023,N_8012);
nor U9317 (N_9317,N_8582,N_8527);
nand U9318 (N_9318,N_8749,N_8158);
or U9319 (N_9319,N_8499,N_8127);
nor U9320 (N_9320,N_8095,N_8811);
and U9321 (N_9321,N_8933,N_8767);
and U9322 (N_9322,N_8016,N_8384);
nor U9323 (N_9323,N_8569,N_8900);
or U9324 (N_9324,N_8984,N_8008);
nor U9325 (N_9325,N_8286,N_8167);
nor U9326 (N_9326,N_8512,N_8976);
and U9327 (N_9327,N_8146,N_8347);
nor U9328 (N_9328,N_8774,N_8349);
nand U9329 (N_9329,N_8425,N_8255);
nand U9330 (N_9330,N_8010,N_8636);
xnor U9331 (N_9331,N_8963,N_8281);
nand U9332 (N_9332,N_8136,N_8477);
and U9333 (N_9333,N_8718,N_8299);
nand U9334 (N_9334,N_8199,N_8122);
nor U9335 (N_9335,N_8936,N_8318);
and U9336 (N_9336,N_8766,N_8206);
nand U9337 (N_9337,N_8335,N_8360);
xor U9338 (N_9338,N_8211,N_8437);
nor U9339 (N_9339,N_8098,N_8770);
nand U9340 (N_9340,N_8288,N_8543);
and U9341 (N_9341,N_8492,N_8156);
or U9342 (N_9342,N_8820,N_8642);
and U9343 (N_9343,N_8472,N_8150);
and U9344 (N_9344,N_8903,N_8276);
nor U9345 (N_9345,N_8950,N_8334);
or U9346 (N_9346,N_8383,N_8982);
or U9347 (N_9347,N_8566,N_8883);
and U9348 (N_9348,N_8067,N_8675);
nand U9349 (N_9349,N_8709,N_8087);
nand U9350 (N_9350,N_8223,N_8862);
nor U9351 (N_9351,N_8411,N_8594);
nand U9352 (N_9352,N_8737,N_8473);
or U9353 (N_9353,N_8330,N_8420);
xor U9354 (N_9354,N_8813,N_8864);
nor U9355 (N_9355,N_8380,N_8780);
nand U9356 (N_9356,N_8791,N_8202);
nor U9357 (N_9357,N_8074,N_8981);
nand U9358 (N_9358,N_8876,N_8781);
and U9359 (N_9359,N_8657,N_8921);
or U9360 (N_9360,N_8340,N_8555);
nor U9361 (N_9361,N_8720,N_8461);
or U9362 (N_9362,N_8847,N_8630);
nand U9363 (N_9363,N_8747,N_8546);
or U9364 (N_9364,N_8607,N_8586);
and U9365 (N_9365,N_8100,N_8129);
nor U9366 (N_9366,N_8061,N_8374);
or U9367 (N_9367,N_8953,N_8320);
nand U9368 (N_9368,N_8049,N_8951);
or U9369 (N_9369,N_8453,N_8224);
nand U9370 (N_9370,N_8157,N_8083);
nand U9371 (N_9371,N_8081,N_8404);
and U9372 (N_9372,N_8378,N_8771);
and U9373 (N_9373,N_8782,N_8210);
nand U9374 (N_9374,N_8525,N_8052);
or U9375 (N_9375,N_8178,N_8621);
nand U9376 (N_9376,N_8703,N_8690);
nand U9377 (N_9377,N_8744,N_8018);
and U9378 (N_9378,N_8406,N_8218);
nand U9379 (N_9379,N_8836,N_8485);
or U9380 (N_9380,N_8684,N_8448);
nor U9381 (N_9381,N_8600,N_8339);
nand U9382 (N_9382,N_8372,N_8861);
nand U9383 (N_9383,N_8761,N_8547);
nand U9384 (N_9384,N_8312,N_8486);
nand U9385 (N_9385,N_8423,N_8641);
or U9386 (N_9386,N_8285,N_8096);
nor U9387 (N_9387,N_8694,N_8357);
or U9388 (N_9388,N_8290,N_8837);
nor U9389 (N_9389,N_8490,N_8221);
and U9390 (N_9390,N_8593,N_8257);
and U9391 (N_9391,N_8164,N_8102);
or U9392 (N_9392,N_8511,N_8142);
nand U9393 (N_9393,N_8872,N_8707);
nor U9394 (N_9394,N_8217,N_8825);
or U9395 (N_9395,N_8238,N_8961);
nor U9396 (N_9396,N_8700,N_8470);
and U9397 (N_9397,N_8599,N_8097);
nand U9398 (N_9398,N_8495,N_8126);
nor U9399 (N_9399,N_8911,N_8019);
and U9400 (N_9400,N_8195,N_8615);
and U9401 (N_9401,N_8308,N_8416);
nor U9402 (N_9402,N_8804,N_8405);
nand U9403 (N_9403,N_8346,N_8305);
nand U9404 (N_9404,N_8814,N_8358);
and U9405 (N_9405,N_8681,N_8563);
or U9406 (N_9406,N_8068,N_8066);
and U9407 (N_9407,N_8591,N_8456);
or U9408 (N_9408,N_8237,N_8004);
or U9409 (N_9409,N_8093,N_8964);
nand U9410 (N_9410,N_8777,N_8743);
or U9411 (N_9411,N_8585,N_8764);
nor U9412 (N_9412,N_8588,N_8215);
or U9413 (N_9413,N_8570,N_8341);
and U9414 (N_9414,N_8256,N_8379);
and U9415 (N_9415,N_8481,N_8166);
nand U9416 (N_9416,N_8442,N_8553);
nand U9417 (N_9417,N_8110,N_8413);
and U9418 (N_9418,N_8701,N_8918);
or U9419 (N_9419,N_8920,N_8231);
or U9420 (N_9420,N_8504,N_8057);
or U9421 (N_9421,N_8388,N_8556);
nand U9422 (N_9422,N_8200,N_8728);
and U9423 (N_9423,N_8852,N_8913);
nor U9424 (N_9424,N_8715,N_8790);
and U9425 (N_9425,N_8863,N_8306);
nor U9426 (N_9426,N_8447,N_8652);
or U9427 (N_9427,N_8280,N_8680);
and U9428 (N_9428,N_8270,N_8355);
nand U9429 (N_9429,N_8148,N_8187);
nor U9430 (N_9430,N_8874,N_8658);
or U9431 (N_9431,N_8054,N_8174);
or U9432 (N_9432,N_8560,N_8892);
and U9433 (N_9433,N_8350,N_8866);
nand U9434 (N_9434,N_8441,N_8300);
xnor U9435 (N_9435,N_8244,N_8783);
or U9436 (N_9436,N_8502,N_8415);
nand U9437 (N_9437,N_8386,N_8125);
or U9438 (N_9438,N_8882,N_8705);
and U9439 (N_9439,N_8440,N_8233);
nor U9440 (N_9440,N_8841,N_8938);
nor U9441 (N_9441,N_8677,N_8443);
nor U9442 (N_9442,N_8177,N_8230);
or U9443 (N_9443,N_8353,N_8601);
nor U9444 (N_9444,N_8026,N_8282);
and U9445 (N_9445,N_8822,N_8297);
nor U9446 (N_9446,N_8035,N_8219);
and U9447 (N_9447,N_8373,N_8351);
nor U9448 (N_9448,N_8069,N_8015);
nor U9449 (N_9449,N_8710,N_8259);
xnor U9450 (N_9450,N_8753,N_8389);
nand U9451 (N_9451,N_8845,N_8612);
nor U9452 (N_9452,N_8429,N_8283);
and U9453 (N_9453,N_8385,N_8661);
or U9454 (N_9454,N_8275,N_8769);
xor U9455 (N_9455,N_8827,N_8402);
nor U9456 (N_9456,N_8966,N_8075);
and U9457 (N_9457,N_8973,N_8410);
xnor U9458 (N_9458,N_8322,N_8422);
or U9459 (N_9459,N_8455,N_8559);
or U9460 (N_9460,N_8778,N_8112);
nand U9461 (N_9461,N_8457,N_8939);
nor U9462 (N_9462,N_8182,N_8958);
nand U9463 (N_9463,N_8634,N_8734);
or U9464 (N_9464,N_8190,N_8888);
or U9465 (N_9465,N_8759,N_8890);
or U9466 (N_9466,N_8549,N_8162);
nor U9467 (N_9467,N_8091,N_8414);
nand U9468 (N_9468,N_8912,N_8923);
nand U9469 (N_9469,N_8520,N_8596);
and U9470 (N_9470,N_8085,N_8216);
nor U9471 (N_9471,N_8176,N_8942);
nand U9472 (N_9472,N_8653,N_8160);
or U9473 (N_9473,N_8584,N_8532);
and U9474 (N_9474,N_8204,N_8975);
nand U9475 (N_9475,N_8089,N_8466);
nor U9476 (N_9476,N_8668,N_8562);
nand U9477 (N_9477,N_8433,N_8051);
and U9478 (N_9478,N_8616,N_8829);
nand U9479 (N_9479,N_8934,N_8262);
nand U9480 (N_9480,N_8924,N_8489);
nor U9481 (N_9481,N_8343,N_8107);
and U9482 (N_9482,N_8464,N_8366);
and U9483 (N_9483,N_8992,N_8576);
nand U9484 (N_9484,N_8382,N_8712);
nor U9485 (N_9485,N_8870,N_8278);
nand U9486 (N_9486,N_8132,N_8145);
nand U9487 (N_9487,N_8434,N_8088);
and U9488 (N_9488,N_8974,N_8409);
or U9489 (N_9489,N_8082,N_8269);
or U9490 (N_9490,N_8301,N_8153);
nand U9491 (N_9491,N_8289,N_8881);
and U9492 (N_9492,N_8793,N_8128);
and U9493 (N_9493,N_8073,N_8518);
or U9494 (N_9494,N_8310,N_8151);
and U9495 (N_9495,N_8510,N_8895);
nor U9496 (N_9496,N_8815,N_8064);
and U9497 (N_9497,N_8611,N_8080);
and U9498 (N_9498,N_8147,N_8121);
or U9499 (N_9499,N_8752,N_8207);
nor U9500 (N_9500,N_8263,N_8670);
or U9501 (N_9501,N_8879,N_8898);
and U9502 (N_9502,N_8069,N_8280);
nor U9503 (N_9503,N_8505,N_8163);
nor U9504 (N_9504,N_8631,N_8560);
nor U9505 (N_9505,N_8041,N_8560);
nand U9506 (N_9506,N_8909,N_8309);
nor U9507 (N_9507,N_8475,N_8942);
and U9508 (N_9508,N_8626,N_8069);
and U9509 (N_9509,N_8710,N_8315);
nand U9510 (N_9510,N_8122,N_8966);
nand U9511 (N_9511,N_8638,N_8811);
nand U9512 (N_9512,N_8464,N_8122);
xor U9513 (N_9513,N_8477,N_8334);
nor U9514 (N_9514,N_8003,N_8985);
nor U9515 (N_9515,N_8512,N_8638);
nor U9516 (N_9516,N_8182,N_8129);
or U9517 (N_9517,N_8328,N_8985);
xnor U9518 (N_9518,N_8795,N_8373);
or U9519 (N_9519,N_8678,N_8061);
nor U9520 (N_9520,N_8261,N_8260);
or U9521 (N_9521,N_8199,N_8908);
or U9522 (N_9522,N_8582,N_8993);
nor U9523 (N_9523,N_8325,N_8377);
or U9524 (N_9524,N_8997,N_8662);
and U9525 (N_9525,N_8494,N_8295);
xor U9526 (N_9526,N_8755,N_8269);
and U9527 (N_9527,N_8126,N_8163);
nor U9528 (N_9528,N_8126,N_8187);
xnor U9529 (N_9529,N_8601,N_8187);
nor U9530 (N_9530,N_8585,N_8314);
nor U9531 (N_9531,N_8617,N_8539);
nor U9532 (N_9532,N_8130,N_8092);
or U9533 (N_9533,N_8685,N_8665);
or U9534 (N_9534,N_8806,N_8165);
or U9535 (N_9535,N_8824,N_8759);
and U9536 (N_9536,N_8967,N_8060);
and U9537 (N_9537,N_8615,N_8069);
nor U9538 (N_9538,N_8166,N_8229);
nand U9539 (N_9539,N_8449,N_8968);
and U9540 (N_9540,N_8173,N_8481);
nand U9541 (N_9541,N_8380,N_8243);
or U9542 (N_9542,N_8814,N_8912);
and U9543 (N_9543,N_8819,N_8746);
nand U9544 (N_9544,N_8202,N_8941);
or U9545 (N_9545,N_8760,N_8703);
nor U9546 (N_9546,N_8024,N_8207);
nand U9547 (N_9547,N_8167,N_8442);
nand U9548 (N_9548,N_8720,N_8669);
and U9549 (N_9549,N_8776,N_8392);
or U9550 (N_9550,N_8661,N_8499);
and U9551 (N_9551,N_8599,N_8608);
nand U9552 (N_9552,N_8252,N_8602);
nor U9553 (N_9553,N_8523,N_8040);
nand U9554 (N_9554,N_8828,N_8291);
and U9555 (N_9555,N_8052,N_8907);
nand U9556 (N_9556,N_8031,N_8386);
or U9557 (N_9557,N_8109,N_8830);
or U9558 (N_9558,N_8779,N_8465);
nor U9559 (N_9559,N_8020,N_8264);
nand U9560 (N_9560,N_8840,N_8716);
or U9561 (N_9561,N_8736,N_8455);
nand U9562 (N_9562,N_8313,N_8402);
nor U9563 (N_9563,N_8231,N_8884);
and U9564 (N_9564,N_8360,N_8305);
nor U9565 (N_9565,N_8439,N_8515);
and U9566 (N_9566,N_8530,N_8197);
nand U9567 (N_9567,N_8680,N_8397);
nor U9568 (N_9568,N_8599,N_8383);
and U9569 (N_9569,N_8011,N_8432);
nor U9570 (N_9570,N_8252,N_8907);
nor U9571 (N_9571,N_8394,N_8090);
and U9572 (N_9572,N_8365,N_8761);
nor U9573 (N_9573,N_8125,N_8720);
or U9574 (N_9574,N_8039,N_8588);
nor U9575 (N_9575,N_8204,N_8383);
and U9576 (N_9576,N_8473,N_8112);
nand U9577 (N_9577,N_8045,N_8474);
nand U9578 (N_9578,N_8647,N_8053);
nand U9579 (N_9579,N_8845,N_8819);
and U9580 (N_9580,N_8729,N_8315);
nor U9581 (N_9581,N_8209,N_8517);
or U9582 (N_9582,N_8056,N_8624);
nand U9583 (N_9583,N_8491,N_8773);
and U9584 (N_9584,N_8746,N_8933);
nor U9585 (N_9585,N_8118,N_8627);
and U9586 (N_9586,N_8418,N_8143);
nand U9587 (N_9587,N_8339,N_8765);
nor U9588 (N_9588,N_8625,N_8710);
nand U9589 (N_9589,N_8328,N_8842);
and U9590 (N_9590,N_8954,N_8862);
and U9591 (N_9591,N_8514,N_8632);
or U9592 (N_9592,N_8292,N_8863);
and U9593 (N_9593,N_8861,N_8696);
and U9594 (N_9594,N_8060,N_8229);
nor U9595 (N_9595,N_8469,N_8476);
nor U9596 (N_9596,N_8385,N_8061);
or U9597 (N_9597,N_8654,N_8320);
or U9598 (N_9598,N_8436,N_8283);
and U9599 (N_9599,N_8730,N_8418);
xnor U9600 (N_9600,N_8653,N_8193);
and U9601 (N_9601,N_8441,N_8336);
or U9602 (N_9602,N_8370,N_8368);
nand U9603 (N_9603,N_8512,N_8740);
or U9604 (N_9604,N_8366,N_8154);
or U9605 (N_9605,N_8878,N_8792);
nand U9606 (N_9606,N_8705,N_8040);
or U9607 (N_9607,N_8775,N_8117);
and U9608 (N_9608,N_8581,N_8017);
or U9609 (N_9609,N_8190,N_8969);
nor U9610 (N_9610,N_8664,N_8470);
nor U9611 (N_9611,N_8147,N_8764);
nand U9612 (N_9612,N_8203,N_8995);
nand U9613 (N_9613,N_8875,N_8759);
and U9614 (N_9614,N_8554,N_8347);
or U9615 (N_9615,N_8769,N_8095);
and U9616 (N_9616,N_8183,N_8744);
nor U9617 (N_9617,N_8558,N_8107);
and U9618 (N_9618,N_8400,N_8346);
or U9619 (N_9619,N_8257,N_8583);
nand U9620 (N_9620,N_8267,N_8724);
nor U9621 (N_9621,N_8097,N_8738);
or U9622 (N_9622,N_8214,N_8560);
nor U9623 (N_9623,N_8883,N_8878);
xor U9624 (N_9624,N_8557,N_8985);
or U9625 (N_9625,N_8852,N_8930);
and U9626 (N_9626,N_8264,N_8512);
nand U9627 (N_9627,N_8864,N_8409);
and U9628 (N_9628,N_8937,N_8866);
nand U9629 (N_9629,N_8743,N_8493);
nand U9630 (N_9630,N_8140,N_8857);
nor U9631 (N_9631,N_8752,N_8043);
nor U9632 (N_9632,N_8695,N_8296);
nor U9633 (N_9633,N_8792,N_8448);
nor U9634 (N_9634,N_8047,N_8790);
or U9635 (N_9635,N_8032,N_8408);
and U9636 (N_9636,N_8210,N_8184);
and U9637 (N_9637,N_8904,N_8808);
nor U9638 (N_9638,N_8667,N_8106);
xnor U9639 (N_9639,N_8543,N_8935);
and U9640 (N_9640,N_8550,N_8485);
or U9641 (N_9641,N_8780,N_8297);
nand U9642 (N_9642,N_8744,N_8230);
and U9643 (N_9643,N_8539,N_8294);
nor U9644 (N_9644,N_8382,N_8561);
and U9645 (N_9645,N_8903,N_8842);
nand U9646 (N_9646,N_8479,N_8826);
and U9647 (N_9647,N_8969,N_8883);
and U9648 (N_9648,N_8807,N_8107);
nor U9649 (N_9649,N_8681,N_8943);
or U9650 (N_9650,N_8088,N_8697);
xnor U9651 (N_9651,N_8974,N_8178);
nand U9652 (N_9652,N_8326,N_8754);
or U9653 (N_9653,N_8873,N_8658);
nand U9654 (N_9654,N_8558,N_8625);
nor U9655 (N_9655,N_8146,N_8024);
or U9656 (N_9656,N_8914,N_8050);
and U9657 (N_9657,N_8609,N_8544);
nor U9658 (N_9658,N_8232,N_8852);
nor U9659 (N_9659,N_8304,N_8284);
and U9660 (N_9660,N_8939,N_8398);
or U9661 (N_9661,N_8423,N_8960);
and U9662 (N_9662,N_8576,N_8146);
and U9663 (N_9663,N_8887,N_8690);
and U9664 (N_9664,N_8098,N_8970);
xor U9665 (N_9665,N_8515,N_8901);
and U9666 (N_9666,N_8374,N_8665);
nor U9667 (N_9667,N_8407,N_8059);
nand U9668 (N_9668,N_8261,N_8738);
and U9669 (N_9669,N_8847,N_8039);
and U9670 (N_9670,N_8155,N_8128);
xor U9671 (N_9671,N_8578,N_8985);
nand U9672 (N_9672,N_8446,N_8709);
nor U9673 (N_9673,N_8183,N_8933);
nand U9674 (N_9674,N_8407,N_8903);
nand U9675 (N_9675,N_8774,N_8438);
nor U9676 (N_9676,N_8210,N_8924);
nand U9677 (N_9677,N_8846,N_8619);
or U9678 (N_9678,N_8441,N_8284);
and U9679 (N_9679,N_8888,N_8136);
nor U9680 (N_9680,N_8151,N_8921);
nor U9681 (N_9681,N_8472,N_8996);
nand U9682 (N_9682,N_8315,N_8984);
nor U9683 (N_9683,N_8707,N_8083);
nor U9684 (N_9684,N_8128,N_8298);
nand U9685 (N_9685,N_8790,N_8512);
nor U9686 (N_9686,N_8008,N_8818);
and U9687 (N_9687,N_8808,N_8590);
xnor U9688 (N_9688,N_8547,N_8012);
nand U9689 (N_9689,N_8659,N_8272);
and U9690 (N_9690,N_8522,N_8125);
or U9691 (N_9691,N_8515,N_8460);
xnor U9692 (N_9692,N_8728,N_8445);
nand U9693 (N_9693,N_8333,N_8679);
nor U9694 (N_9694,N_8875,N_8411);
nor U9695 (N_9695,N_8172,N_8628);
or U9696 (N_9696,N_8102,N_8939);
nor U9697 (N_9697,N_8593,N_8081);
or U9698 (N_9698,N_8287,N_8135);
and U9699 (N_9699,N_8312,N_8188);
or U9700 (N_9700,N_8246,N_8358);
and U9701 (N_9701,N_8482,N_8633);
or U9702 (N_9702,N_8163,N_8546);
nand U9703 (N_9703,N_8802,N_8504);
nor U9704 (N_9704,N_8574,N_8051);
or U9705 (N_9705,N_8297,N_8806);
or U9706 (N_9706,N_8403,N_8110);
nor U9707 (N_9707,N_8380,N_8460);
nor U9708 (N_9708,N_8591,N_8125);
and U9709 (N_9709,N_8907,N_8326);
nor U9710 (N_9710,N_8249,N_8274);
nand U9711 (N_9711,N_8569,N_8602);
nor U9712 (N_9712,N_8555,N_8354);
xor U9713 (N_9713,N_8520,N_8794);
nor U9714 (N_9714,N_8653,N_8281);
nor U9715 (N_9715,N_8969,N_8506);
nand U9716 (N_9716,N_8665,N_8593);
nand U9717 (N_9717,N_8449,N_8906);
nor U9718 (N_9718,N_8194,N_8289);
or U9719 (N_9719,N_8905,N_8026);
nor U9720 (N_9720,N_8390,N_8203);
nor U9721 (N_9721,N_8965,N_8076);
and U9722 (N_9722,N_8833,N_8318);
or U9723 (N_9723,N_8397,N_8418);
nor U9724 (N_9724,N_8959,N_8301);
or U9725 (N_9725,N_8453,N_8467);
nor U9726 (N_9726,N_8311,N_8093);
nand U9727 (N_9727,N_8882,N_8933);
or U9728 (N_9728,N_8711,N_8349);
nor U9729 (N_9729,N_8593,N_8771);
and U9730 (N_9730,N_8850,N_8201);
or U9731 (N_9731,N_8876,N_8322);
and U9732 (N_9732,N_8254,N_8190);
or U9733 (N_9733,N_8554,N_8548);
xnor U9734 (N_9734,N_8695,N_8395);
and U9735 (N_9735,N_8265,N_8500);
nor U9736 (N_9736,N_8191,N_8386);
nor U9737 (N_9737,N_8676,N_8952);
nand U9738 (N_9738,N_8326,N_8849);
and U9739 (N_9739,N_8279,N_8674);
nor U9740 (N_9740,N_8857,N_8239);
nand U9741 (N_9741,N_8001,N_8241);
nor U9742 (N_9742,N_8415,N_8757);
nor U9743 (N_9743,N_8460,N_8480);
xnor U9744 (N_9744,N_8721,N_8032);
nor U9745 (N_9745,N_8077,N_8039);
nor U9746 (N_9746,N_8277,N_8288);
nor U9747 (N_9747,N_8452,N_8190);
nor U9748 (N_9748,N_8836,N_8607);
nor U9749 (N_9749,N_8097,N_8270);
and U9750 (N_9750,N_8714,N_8948);
nor U9751 (N_9751,N_8101,N_8680);
nor U9752 (N_9752,N_8728,N_8417);
nand U9753 (N_9753,N_8501,N_8184);
nor U9754 (N_9754,N_8614,N_8984);
nand U9755 (N_9755,N_8407,N_8642);
nand U9756 (N_9756,N_8473,N_8216);
nor U9757 (N_9757,N_8669,N_8844);
and U9758 (N_9758,N_8420,N_8537);
and U9759 (N_9759,N_8631,N_8817);
nor U9760 (N_9760,N_8970,N_8629);
or U9761 (N_9761,N_8187,N_8750);
and U9762 (N_9762,N_8118,N_8556);
and U9763 (N_9763,N_8842,N_8006);
and U9764 (N_9764,N_8824,N_8410);
xnor U9765 (N_9765,N_8076,N_8195);
or U9766 (N_9766,N_8809,N_8668);
nand U9767 (N_9767,N_8326,N_8474);
or U9768 (N_9768,N_8722,N_8243);
nand U9769 (N_9769,N_8470,N_8980);
nand U9770 (N_9770,N_8364,N_8855);
nor U9771 (N_9771,N_8777,N_8601);
or U9772 (N_9772,N_8796,N_8000);
nand U9773 (N_9773,N_8420,N_8052);
nor U9774 (N_9774,N_8559,N_8764);
and U9775 (N_9775,N_8229,N_8913);
and U9776 (N_9776,N_8486,N_8488);
xor U9777 (N_9777,N_8041,N_8877);
nand U9778 (N_9778,N_8955,N_8044);
or U9779 (N_9779,N_8783,N_8682);
nor U9780 (N_9780,N_8783,N_8296);
nor U9781 (N_9781,N_8536,N_8717);
and U9782 (N_9782,N_8018,N_8025);
nor U9783 (N_9783,N_8212,N_8218);
nand U9784 (N_9784,N_8198,N_8658);
nor U9785 (N_9785,N_8977,N_8518);
nand U9786 (N_9786,N_8145,N_8478);
nand U9787 (N_9787,N_8293,N_8039);
nor U9788 (N_9788,N_8800,N_8382);
or U9789 (N_9789,N_8701,N_8392);
nor U9790 (N_9790,N_8799,N_8709);
and U9791 (N_9791,N_8180,N_8467);
and U9792 (N_9792,N_8997,N_8896);
nor U9793 (N_9793,N_8692,N_8527);
nand U9794 (N_9794,N_8973,N_8279);
nor U9795 (N_9795,N_8036,N_8678);
and U9796 (N_9796,N_8148,N_8792);
nand U9797 (N_9797,N_8559,N_8041);
nor U9798 (N_9798,N_8969,N_8740);
or U9799 (N_9799,N_8153,N_8762);
nor U9800 (N_9800,N_8297,N_8207);
and U9801 (N_9801,N_8656,N_8864);
nand U9802 (N_9802,N_8088,N_8429);
and U9803 (N_9803,N_8159,N_8451);
or U9804 (N_9804,N_8591,N_8063);
nand U9805 (N_9805,N_8280,N_8972);
nand U9806 (N_9806,N_8945,N_8742);
nor U9807 (N_9807,N_8012,N_8686);
xor U9808 (N_9808,N_8903,N_8392);
and U9809 (N_9809,N_8414,N_8030);
or U9810 (N_9810,N_8555,N_8421);
nand U9811 (N_9811,N_8044,N_8441);
or U9812 (N_9812,N_8412,N_8768);
nor U9813 (N_9813,N_8298,N_8700);
or U9814 (N_9814,N_8130,N_8084);
nand U9815 (N_9815,N_8818,N_8497);
nor U9816 (N_9816,N_8115,N_8624);
or U9817 (N_9817,N_8194,N_8768);
nor U9818 (N_9818,N_8710,N_8833);
and U9819 (N_9819,N_8168,N_8020);
and U9820 (N_9820,N_8483,N_8396);
or U9821 (N_9821,N_8199,N_8468);
and U9822 (N_9822,N_8698,N_8598);
nand U9823 (N_9823,N_8214,N_8151);
nor U9824 (N_9824,N_8955,N_8705);
or U9825 (N_9825,N_8946,N_8267);
and U9826 (N_9826,N_8699,N_8672);
and U9827 (N_9827,N_8162,N_8894);
nand U9828 (N_9828,N_8741,N_8100);
nor U9829 (N_9829,N_8944,N_8272);
nand U9830 (N_9830,N_8410,N_8929);
and U9831 (N_9831,N_8822,N_8399);
nand U9832 (N_9832,N_8637,N_8355);
or U9833 (N_9833,N_8202,N_8370);
nand U9834 (N_9834,N_8493,N_8611);
or U9835 (N_9835,N_8143,N_8337);
and U9836 (N_9836,N_8536,N_8187);
or U9837 (N_9837,N_8642,N_8177);
nand U9838 (N_9838,N_8131,N_8914);
nand U9839 (N_9839,N_8419,N_8500);
and U9840 (N_9840,N_8104,N_8717);
xnor U9841 (N_9841,N_8321,N_8446);
and U9842 (N_9842,N_8142,N_8176);
nor U9843 (N_9843,N_8073,N_8469);
nand U9844 (N_9844,N_8318,N_8238);
and U9845 (N_9845,N_8985,N_8008);
nand U9846 (N_9846,N_8358,N_8296);
nor U9847 (N_9847,N_8478,N_8225);
or U9848 (N_9848,N_8495,N_8365);
or U9849 (N_9849,N_8459,N_8969);
and U9850 (N_9850,N_8140,N_8204);
nor U9851 (N_9851,N_8781,N_8837);
nand U9852 (N_9852,N_8305,N_8386);
nand U9853 (N_9853,N_8274,N_8132);
nor U9854 (N_9854,N_8866,N_8064);
nor U9855 (N_9855,N_8326,N_8552);
nand U9856 (N_9856,N_8010,N_8776);
nand U9857 (N_9857,N_8983,N_8236);
and U9858 (N_9858,N_8362,N_8902);
or U9859 (N_9859,N_8739,N_8745);
nand U9860 (N_9860,N_8277,N_8593);
or U9861 (N_9861,N_8239,N_8195);
nand U9862 (N_9862,N_8949,N_8317);
or U9863 (N_9863,N_8358,N_8542);
and U9864 (N_9864,N_8062,N_8374);
or U9865 (N_9865,N_8260,N_8464);
or U9866 (N_9866,N_8598,N_8697);
nand U9867 (N_9867,N_8365,N_8297);
xor U9868 (N_9868,N_8290,N_8766);
nand U9869 (N_9869,N_8161,N_8924);
nor U9870 (N_9870,N_8696,N_8859);
or U9871 (N_9871,N_8250,N_8697);
nor U9872 (N_9872,N_8088,N_8567);
or U9873 (N_9873,N_8589,N_8135);
or U9874 (N_9874,N_8978,N_8956);
or U9875 (N_9875,N_8806,N_8527);
nor U9876 (N_9876,N_8375,N_8073);
or U9877 (N_9877,N_8318,N_8577);
nand U9878 (N_9878,N_8823,N_8957);
and U9879 (N_9879,N_8928,N_8862);
and U9880 (N_9880,N_8832,N_8112);
nor U9881 (N_9881,N_8659,N_8586);
and U9882 (N_9882,N_8800,N_8328);
or U9883 (N_9883,N_8422,N_8012);
or U9884 (N_9884,N_8985,N_8937);
nor U9885 (N_9885,N_8503,N_8658);
nor U9886 (N_9886,N_8004,N_8771);
nor U9887 (N_9887,N_8462,N_8010);
and U9888 (N_9888,N_8784,N_8216);
nand U9889 (N_9889,N_8196,N_8088);
nor U9890 (N_9890,N_8749,N_8078);
and U9891 (N_9891,N_8366,N_8167);
and U9892 (N_9892,N_8661,N_8141);
nor U9893 (N_9893,N_8668,N_8367);
nor U9894 (N_9894,N_8804,N_8863);
nor U9895 (N_9895,N_8685,N_8986);
nand U9896 (N_9896,N_8250,N_8807);
or U9897 (N_9897,N_8393,N_8568);
and U9898 (N_9898,N_8369,N_8045);
nand U9899 (N_9899,N_8517,N_8752);
and U9900 (N_9900,N_8755,N_8425);
nand U9901 (N_9901,N_8397,N_8827);
nand U9902 (N_9902,N_8084,N_8816);
or U9903 (N_9903,N_8913,N_8921);
xor U9904 (N_9904,N_8663,N_8714);
or U9905 (N_9905,N_8892,N_8652);
nand U9906 (N_9906,N_8975,N_8631);
or U9907 (N_9907,N_8899,N_8203);
nand U9908 (N_9908,N_8507,N_8131);
or U9909 (N_9909,N_8276,N_8771);
nand U9910 (N_9910,N_8907,N_8064);
nand U9911 (N_9911,N_8375,N_8844);
nand U9912 (N_9912,N_8662,N_8828);
and U9913 (N_9913,N_8168,N_8196);
and U9914 (N_9914,N_8659,N_8747);
and U9915 (N_9915,N_8375,N_8231);
nor U9916 (N_9916,N_8172,N_8217);
nor U9917 (N_9917,N_8219,N_8142);
nand U9918 (N_9918,N_8381,N_8879);
nor U9919 (N_9919,N_8161,N_8417);
and U9920 (N_9920,N_8799,N_8392);
nand U9921 (N_9921,N_8529,N_8432);
xor U9922 (N_9922,N_8029,N_8113);
and U9923 (N_9923,N_8070,N_8463);
or U9924 (N_9924,N_8737,N_8070);
nand U9925 (N_9925,N_8607,N_8463);
xor U9926 (N_9926,N_8657,N_8770);
and U9927 (N_9927,N_8148,N_8785);
or U9928 (N_9928,N_8988,N_8132);
xor U9929 (N_9929,N_8806,N_8208);
or U9930 (N_9930,N_8582,N_8906);
nor U9931 (N_9931,N_8811,N_8463);
or U9932 (N_9932,N_8490,N_8270);
nor U9933 (N_9933,N_8405,N_8221);
or U9934 (N_9934,N_8729,N_8340);
nand U9935 (N_9935,N_8574,N_8189);
nor U9936 (N_9936,N_8652,N_8107);
nor U9937 (N_9937,N_8146,N_8752);
or U9938 (N_9938,N_8490,N_8585);
or U9939 (N_9939,N_8715,N_8992);
nor U9940 (N_9940,N_8159,N_8576);
or U9941 (N_9941,N_8717,N_8439);
nor U9942 (N_9942,N_8809,N_8209);
or U9943 (N_9943,N_8954,N_8802);
or U9944 (N_9944,N_8884,N_8428);
or U9945 (N_9945,N_8845,N_8869);
xnor U9946 (N_9946,N_8295,N_8835);
and U9947 (N_9947,N_8578,N_8747);
nand U9948 (N_9948,N_8554,N_8187);
nand U9949 (N_9949,N_8600,N_8667);
nor U9950 (N_9950,N_8151,N_8168);
nand U9951 (N_9951,N_8864,N_8550);
and U9952 (N_9952,N_8850,N_8794);
and U9953 (N_9953,N_8093,N_8662);
and U9954 (N_9954,N_8262,N_8417);
and U9955 (N_9955,N_8542,N_8057);
or U9956 (N_9956,N_8467,N_8861);
or U9957 (N_9957,N_8173,N_8431);
or U9958 (N_9958,N_8662,N_8777);
nor U9959 (N_9959,N_8132,N_8229);
and U9960 (N_9960,N_8245,N_8427);
nor U9961 (N_9961,N_8354,N_8413);
nand U9962 (N_9962,N_8090,N_8685);
or U9963 (N_9963,N_8274,N_8911);
or U9964 (N_9964,N_8454,N_8787);
xor U9965 (N_9965,N_8236,N_8894);
nor U9966 (N_9966,N_8614,N_8734);
and U9967 (N_9967,N_8115,N_8495);
and U9968 (N_9968,N_8142,N_8931);
nor U9969 (N_9969,N_8274,N_8358);
nor U9970 (N_9970,N_8333,N_8520);
nor U9971 (N_9971,N_8101,N_8520);
xor U9972 (N_9972,N_8935,N_8544);
or U9973 (N_9973,N_8642,N_8238);
and U9974 (N_9974,N_8333,N_8904);
xor U9975 (N_9975,N_8819,N_8040);
and U9976 (N_9976,N_8984,N_8692);
and U9977 (N_9977,N_8220,N_8330);
nand U9978 (N_9978,N_8835,N_8870);
nor U9979 (N_9979,N_8889,N_8391);
and U9980 (N_9980,N_8167,N_8850);
nor U9981 (N_9981,N_8552,N_8462);
and U9982 (N_9982,N_8520,N_8291);
and U9983 (N_9983,N_8338,N_8180);
or U9984 (N_9984,N_8479,N_8892);
nor U9985 (N_9985,N_8302,N_8534);
nor U9986 (N_9986,N_8914,N_8730);
nand U9987 (N_9987,N_8364,N_8188);
or U9988 (N_9988,N_8197,N_8363);
nand U9989 (N_9989,N_8346,N_8638);
and U9990 (N_9990,N_8805,N_8747);
nor U9991 (N_9991,N_8220,N_8721);
nand U9992 (N_9992,N_8683,N_8588);
nand U9993 (N_9993,N_8438,N_8437);
nor U9994 (N_9994,N_8416,N_8598);
nor U9995 (N_9995,N_8586,N_8412);
nand U9996 (N_9996,N_8044,N_8666);
nor U9997 (N_9997,N_8841,N_8849);
nand U9998 (N_9998,N_8529,N_8256);
nor U9999 (N_9999,N_8101,N_8583);
nand UO_0 (O_0,N_9420,N_9365);
nand UO_1 (O_1,N_9873,N_9599);
and UO_2 (O_2,N_9082,N_9581);
and UO_3 (O_3,N_9959,N_9839);
or UO_4 (O_4,N_9096,N_9467);
and UO_5 (O_5,N_9616,N_9194);
xnor UO_6 (O_6,N_9484,N_9674);
and UO_7 (O_7,N_9097,N_9042);
or UO_8 (O_8,N_9753,N_9047);
or UO_9 (O_9,N_9626,N_9689);
and UO_10 (O_10,N_9911,N_9174);
nor UO_11 (O_11,N_9267,N_9727);
or UO_12 (O_12,N_9854,N_9140);
nand UO_13 (O_13,N_9395,N_9255);
nor UO_14 (O_14,N_9747,N_9981);
and UO_15 (O_15,N_9299,N_9790);
and UO_16 (O_16,N_9912,N_9593);
nor UO_17 (O_17,N_9410,N_9202);
nand UO_18 (O_18,N_9906,N_9373);
or UO_19 (O_19,N_9745,N_9837);
nand UO_20 (O_20,N_9519,N_9513);
and UO_21 (O_21,N_9640,N_9526);
or UO_22 (O_22,N_9243,N_9936);
nor UO_23 (O_23,N_9233,N_9273);
nor UO_24 (O_24,N_9230,N_9771);
nor UO_25 (O_25,N_9154,N_9320);
nand UO_26 (O_26,N_9792,N_9662);
or UO_27 (O_27,N_9426,N_9547);
and UO_28 (O_28,N_9372,N_9666);
xnor UO_29 (O_29,N_9432,N_9163);
or UO_30 (O_30,N_9677,N_9569);
or UO_31 (O_31,N_9788,N_9014);
and UO_32 (O_32,N_9356,N_9653);
nor UO_33 (O_33,N_9607,N_9774);
nor UO_34 (O_34,N_9120,N_9483);
and UO_35 (O_35,N_9425,N_9785);
xnor UO_36 (O_36,N_9571,N_9590);
nand UO_37 (O_37,N_9602,N_9656);
nor UO_38 (O_38,N_9704,N_9846);
nor UO_39 (O_39,N_9076,N_9214);
and UO_40 (O_40,N_9634,N_9831);
nand UO_41 (O_41,N_9364,N_9709);
or UO_42 (O_42,N_9326,N_9274);
and UO_43 (O_43,N_9242,N_9754);
nand UO_44 (O_44,N_9670,N_9206);
nand UO_45 (O_45,N_9861,N_9324);
nand UO_46 (O_46,N_9800,N_9770);
or UO_47 (O_47,N_9405,N_9300);
and UO_48 (O_48,N_9226,N_9333);
nand UO_49 (O_49,N_9366,N_9717);
or UO_50 (O_50,N_9996,N_9284);
or UO_51 (O_51,N_9892,N_9382);
nand UO_52 (O_52,N_9714,N_9841);
nand UO_53 (O_53,N_9811,N_9787);
and UO_54 (O_54,N_9789,N_9624);
or UO_55 (O_55,N_9357,N_9767);
nor UO_56 (O_56,N_9481,N_9972);
or UO_57 (O_57,N_9227,N_9309);
and UO_58 (O_58,N_9168,N_9428);
and UO_59 (O_59,N_9715,N_9583);
or UO_60 (O_60,N_9259,N_9612);
or UO_61 (O_61,N_9575,N_9535);
xnor UO_62 (O_62,N_9148,N_9024);
and UO_63 (O_63,N_9947,N_9396);
and UO_64 (O_64,N_9292,N_9471);
nor UO_65 (O_65,N_9825,N_9904);
and UO_66 (O_66,N_9118,N_9129);
nand UO_67 (O_67,N_9700,N_9948);
nor UO_68 (O_68,N_9500,N_9701);
or UO_69 (O_69,N_9399,N_9564);
and UO_70 (O_70,N_9751,N_9992);
nand UO_71 (O_71,N_9113,N_9030);
nor UO_72 (O_72,N_9252,N_9253);
nand UO_73 (O_73,N_9625,N_9492);
or UO_74 (O_74,N_9728,N_9560);
or UO_75 (O_75,N_9541,N_9695);
or UO_76 (O_76,N_9524,N_9977);
or UO_77 (O_77,N_9147,N_9777);
or UO_78 (O_78,N_9065,N_9195);
and UO_79 (O_79,N_9579,N_9203);
nor UO_80 (O_80,N_9759,N_9720);
or UO_81 (O_81,N_9217,N_9848);
and UO_82 (O_82,N_9190,N_9394);
nand UO_83 (O_83,N_9974,N_9013);
or UO_84 (O_84,N_9312,N_9922);
nor UO_85 (O_85,N_9913,N_9982);
and UO_86 (O_86,N_9235,N_9946);
or UO_87 (O_87,N_9875,N_9802);
and UO_88 (O_88,N_9872,N_9028);
or UO_89 (O_89,N_9288,N_9139);
and UO_90 (O_90,N_9534,N_9725);
and UO_91 (O_91,N_9138,N_9707);
nor UO_92 (O_92,N_9657,N_9597);
nand UO_93 (O_93,N_9303,N_9499);
nand UO_94 (O_94,N_9810,N_9176);
nor UO_95 (O_95,N_9169,N_9931);
xnor UO_96 (O_96,N_9383,N_9941);
nor UO_97 (O_97,N_9359,N_9536);
xnor UO_98 (O_98,N_9368,N_9048);
nand UO_99 (O_99,N_9291,N_9183);
nand UO_100 (O_100,N_9676,N_9406);
and UO_101 (O_101,N_9488,N_9098);
and UO_102 (O_102,N_9191,N_9845);
or UO_103 (O_103,N_9505,N_9313);
nand UO_104 (O_104,N_9944,N_9463);
and UO_105 (O_105,N_9156,N_9131);
nor UO_106 (O_106,N_9887,N_9630);
nor UO_107 (O_107,N_9344,N_9457);
or UO_108 (O_108,N_9239,N_9315);
or UO_109 (O_109,N_9693,N_9122);
nand UO_110 (O_110,N_9102,N_9298);
nand UO_111 (O_111,N_9671,N_9940);
or UO_112 (O_112,N_9920,N_9991);
or UO_113 (O_113,N_9899,N_9317);
nand UO_114 (O_114,N_9673,N_9658);
and UO_115 (O_115,N_9355,N_9398);
nor UO_116 (O_116,N_9543,N_9108);
nand UO_117 (O_117,N_9435,N_9557);
or UO_118 (O_118,N_9548,N_9863);
nand UO_119 (O_119,N_9971,N_9290);
nand UO_120 (O_120,N_9180,N_9000);
or UO_121 (O_121,N_9185,N_9275);
nor UO_122 (O_122,N_9092,N_9508);
nor UO_123 (O_123,N_9649,N_9330);
nor UO_124 (O_124,N_9442,N_9815);
and UO_125 (O_125,N_9123,N_9026);
nand UO_126 (O_126,N_9043,N_9506);
nor UO_127 (O_127,N_9251,N_9135);
nor UO_128 (O_128,N_9970,N_9393);
xor UO_129 (O_129,N_9350,N_9244);
nand UO_130 (O_130,N_9308,N_9939);
and UO_131 (O_131,N_9145,N_9258);
nor UO_132 (O_132,N_9604,N_9456);
nand UO_133 (O_133,N_9523,N_9278);
or UO_134 (O_134,N_9053,N_9719);
and UO_135 (O_135,N_9149,N_9094);
nand UO_136 (O_136,N_9891,N_9807);
xor UO_137 (O_137,N_9103,N_9472);
nor UO_138 (O_138,N_9723,N_9694);
and UO_139 (O_139,N_9329,N_9306);
nand UO_140 (O_140,N_9438,N_9726);
nor UO_141 (O_141,N_9414,N_9295);
nor UO_142 (O_142,N_9402,N_9808);
nand UO_143 (O_143,N_9384,N_9004);
nand UO_144 (O_144,N_9084,N_9852);
xor UO_145 (O_145,N_9204,N_9124);
nand UO_146 (O_146,N_9431,N_9159);
or UO_147 (O_147,N_9254,N_9083);
or UO_148 (O_148,N_9167,N_9160);
and UO_149 (O_149,N_9611,N_9780);
and UO_150 (O_150,N_9712,N_9552);
nor UO_151 (O_151,N_9462,N_9562);
nor UO_152 (O_152,N_9224,N_9544);
and UO_153 (O_153,N_9563,N_9844);
nand UO_154 (O_154,N_9377,N_9691);
nand UO_155 (O_155,N_9491,N_9933);
or UO_156 (O_156,N_9010,N_9229);
nand UO_157 (O_157,N_9783,N_9647);
and UO_158 (O_158,N_9403,N_9369);
or UO_159 (O_159,N_9280,N_9623);
and UO_160 (O_160,N_9494,N_9928);
nand UO_161 (O_161,N_9137,N_9960);
nand UO_162 (O_162,N_9990,N_9998);
or UO_163 (O_163,N_9056,N_9858);
or UO_164 (O_164,N_9830,N_9643);
nand UO_165 (O_165,N_9521,N_9698);
nor UO_166 (O_166,N_9404,N_9276);
and UO_167 (O_167,N_9018,N_9376);
xnor UO_168 (O_168,N_9595,N_9874);
nand UO_169 (O_169,N_9126,N_9201);
or UO_170 (O_170,N_9798,N_9570);
nand UO_171 (O_171,N_9188,N_9965);
or UO_172 (O_172,N_9900,N_9086);
nor UO_173 (O_173,N_9311,N_9703);
nand UO_174 (O_174,N_9119,N_9460);
nor UO_175 (O_175,N_9989,N_9450);
and UO_176 (O_176,N_9054,N_9121);
nand UO_177 (O_177,N_9757,N_9601);
or UO_178 (O_178,N_9436,N_9710);
nand UO_179 (O_179,N_9608,N_9870);
nand UO_180 (O_180,N_9454,N_9078);
nand UO_181 (O_181,N_9134,N_9824);
or UO_182 (O_182,N_9144,N_9755);
or UO_183 (O_183,N_9015,N_9157);
and UO_184 (O_184,N_9718,N_9504);
or UO_185 (O_185,N_9681,N_9555);
nand UO_186 (O_186,N_9101,N_9627);
or UO_187 (O_187,N_9150,N_9937);
nor UO_188 (O_188,N_9988,N_9877);
or UO_189 (O_189,N_9002,N_9272);
nor UO_190 (O_190,N_9642,N_9051);
nand UO_191 (O_191,N_9896,N_9328);
and UO_192 (O_192,N_9956,N_9071);
nand UO_193 (O_193,N_9060,N_9136);
nand UO_194 (O_194,N_9553,N_9061);
and UO_195 (O_195,N_9832,N_9884);
nor UO_196 (O_196,N_9917,N_9475);
nor UO_197 (O_197,N_9902,N_9362);
and UO_198 (O_198,N_9213,N_9302);
nor UO_199 (O_199,N_9529,N_9908);
or UO_200 (O_200,N_9349,N_9835);
xnor UO_201 (O_201,N_9088,N_9200);
or UO_202 (O_202,N_9155,N_9385);
or UO_203 (O_203,N_9517,N_9577);
nor UO_204 (O_204,N_9423,N_9301);
and UO_205 (O_205,N_9059,N_9542);
and UO_206 (O_206,N_9198,N_9029);
or UO_207 (O_207,N_9584,N_9269);
or UO_208 (O_208,N_9829,N_9044);
and UO_209 (O_209,N_9261,N_9045);
and UO_210 (O_210,N_9158,N_9905);
or UO_211 (O_211,N_9737,N_9687);
and UO_212 (O_212,N_9976,N_9245);
and UO_213 (O_213,N_9983,N_9722);
nor UO_214 (O_214,N_9617,N_9778);
nand UO_215 (O_215,N_9942,N_9416);
or UO_216 (O_216,N_9818,N_9744);
nor UO_217 (O_217,N_9323,N_9938);
nor UO_218 (O_218,N_9378,N_9692);
nand UO_219 (O_219,N_9321,N_9035);
nor UO_220 (O_220,N_9153,N_9146);
or UO_221 (O_221,N_9784,N_9193);
or UO_222 (O_222,N_9424,N_9401);
or UO_223 (O_223,N_9994,N_9479);
or UO_224 (O_224,N_9646,N_9619);
nand UO_225 (O_225,N_9304,N_9192);
nor UO_226 (O_226,N_9008,N_9429);
nand UO_227 (O_227,N_9683,N_9448);
nor UO_228 (O_228,N_9885,N_9455);
nor UO_229 (O_229,N_9133,N_9143);
nor UO_230 (O_230,N_9012,N_9099);
nand UO_231 (O_231,N_9205,N_9470);
xor UO_232 (O_232,N_9182,N_9958);
and UO_233 (O_233,N_9752,N_9980);
nand UO_234 (O_234,N_9476,N_9843);
nor UO_235 (O_235,N_9090,N_9897);
and UO_236 (O_236,N_9164,N_9162);
or UO_237 (O_237,N_9005,N_9016);
nor UO_238 (O_238,N_9019,N_9361);
and UO_239 (O_239,N_9215,N_9865);
and UO_240 (O_240,N_9461,N_9923);
or UO_241 (O_241,N_9170,N_9518);
nand UO_242 (O_242,N_9225,N_9466);
nand UO_243 (O_243,N_9813,N_9417);
nor UO_244 (O_244,N_9914,N_9104);
nand UO_245 (O_245,N_9540,N_9596);
nor UO_246 (O_246,N_9050,N_9111);
or UO_247 (O_247,N_9085,N_9287);
nand UO_248 (O_248,N_9776,N_9352);
nand UO_249 (O_249,N_9172,N_9591);
nand UO_250 (O_250,N_9733,N_9660);
nand UO_251 (O_251,N_9890,N_9341);
xnor UO_252 (O_252,N_9866,N_9696);
or UO_253 (O_253,N_9211,N_9445);
or UO_254 (O_254,N_9270,N_9268);
or UO_255 (O_255,N_9973,N_9685);
nand UO_256 (O_256,N_9550,N_9761);
and UO_257 (O_257,N_9549,N_9916);
nor UO_258 (O_258,N_9978,N_9629);
or UO_259 (O_259,N_9075,N_9794);
nor UO_260 (O_260,N_9801,N_9661);
and UO_261 (O_261,N_9860,N_9963);
nand UO_262 (O_262,N_9294,N_9222);
or UO_263 (O_263,N_9069,N_9052);
nand UO_264 (O_264,N_9574,N_9343);
nand UO_265 (O_265,N_9605,N_9115);
or UO_266 (O_266,N_9446,N_9370);
nand UO_267 (O_267,N_9915,N_9165);
and UO_268 (O_268,N_9512,N_9951);
nand UO_269 (O_269,N_9256,N_9573);
nand UO_270 (O_270,N_9434,N_9567);
or UO_271 (O_271,N_9007,N_9995);
nor UO_272 (O_272,N_9580,N_9477);
xnor UO_273 (O_273,N_9522,N_9207);
or UO_274 (O_274,N_9568,N_9077);
nor UO_275 (O_275,N_9246,N_9561);
nand UO_276 (O_276,N_9351,N_9918);
nand UO_277 (O_277,N_9212,N_9731);
and UO_278 (O_278,N_9682,N_9447);
and UO_279 (O_279,N_9871,N_9708);
and UO_280 (O_280,N_9586,N_9598);
nand UO_281 (O_281,N_9614,N_9651);
nand UO_282 (O_282,N_9697,N_9117);
nor UO_283 (O_283,N_9793,N_9025);
nor UO_284 (O_284,N_9487,N_9836);
or UO_285 (O_285,N_9468,N_9786);
nor UO_286 (O_286,N_9705,N_9441);
or UO_287 (O_287,N_9949,N_9622);
nor UO_288 (O_288,N_9022,N_9859);
and UO_289 (O_289,N_9228,N_9927);
nor UO_290 (O_290,N_9006,N_9699);
or UO_291 (O_291,N_9888,N_9680);
or UO_292 (O_292,N_9023,N_9421);
nand UO_293 (O_293,N_9781,N_9823);
nand UO_294 (O_294,N_9842,N_9663);
or UO_295 (O_295,N_9849,N_9381);
nand UO_296 (O_296,N_9107,N_9391);
nand UO_297 (O_297,N_9110,N_9509);
and UO_298 (O_298,N_9764,N_9934);
or UO_299 (O_299,N_9285,N_9750);
nor UO_300 (O_300,N_9411,N_9910);
or UO_301 (O_301,N_9566,N_9729);
nor UO_302 (O_302,N_9511,N_9962);
nor UO_303 (O_303,N_9089,N_9443);
nor UO_304 (O_304,N_9296,N_9514);
nor UO_305 (O_305,N_9452,N_9017);
and UO_306 (O_306,N_9223,N_9820);
nor UO_307 (O_307,N_9473,N_9062);
and UO_308 (O_308,N_9880,N_9812);
nand UO_309 (O_309,N_9358,N_9072);
nand UO_310 (O_310,N_9894,N_9070);
and UO_311 (O_311,N_9664,N_9773);
and UO_312 (O_312,N_9882,N_9620);
and UO_313 (O_313,N_9641,N_9074);
nor UO_314 (O_314,N_9063,N_9589);
and UO_315 (O_315,N_9679,N_9178);
nor UO_316 (O_316,N_9756,N_9209);
nand UO_317 (O_317,N_9093,N_9392);
and UO_318 (O_318,N_9730,N_9482);
and UO_319 (O_319,N_9895,N_9128);
and UO_320 (O_320,N_9850,N_9307);
or UO_321 (O_321,N_9969,N_9189);
nor UO_322 (O_322,N_9688,N_9503);
nand UO_323 (O_323,N_9868,N_9578);
or UO_324 (O_324,N_9289,N_9961);
nor UO_325 (O_325,N_9112,N_9498);
and UO_326 (O_326,N_9142,N_9458);
and UO_327 (O_327,N_9855,N_9247);
nand UO_328 (O_328,N_9655,N_9449);
or UO_329 (O_329,N_9046,N_9331);
nor UO_330 (O_330,N_9546,N_9415);
nor UO_331 (O_331,N_9100,N_9758);
nor UO_332 (O_332,N_9817,N_9967);
or UO_333 (O_333,N_9430,N_9867);
nor UO_334 (O_334,N_9525,N_9250);
nor UO_335 (O_335,N_9279,N_9265);
xnor UO_336 (O_336,N_9263,N_9496);
and UO_337 (O_337,N_9537,N_9763);
or UO_338 (O_338,N_9125,N_9600);
nor UO_339 (O_339,N_9073,N_9009);
nor UO_340 (O_340,N_9397,N_9637);
or UO_341 (O_341,N_9721,N_9338);
and UO_342 (O_342,N_9132,N_9531);
nand UO_343 (O_343,N_9856,N_9635);
nand UO_344 (O_344,N_9116,N_9196);
and UO_345 (O_345,N_9638,N_9530);
nor UO_346 (O_346,N_9407,N_9277);
nor UO_347 (O_347,N_9502,N_9804);
nor UO_348 (O_348,N_9208,N_9650);
nand UO_349 (O_349,N_9654,N_9197);
xor UO_350 (O_350,N_9186,N_9768);
or UO_351 (O_351,N_9011,N_9316);
and UO_352 (O_352,N_9345,N_9743);
nand UO_353 (O_353,N_9055,N_9171);
or UO_354 (O_354,N_9851,N_9184);
nand UO_355 (O_355,N_9437,N_9440);
or UO_356 (O_356,N_9659,N_9738);
nor UO_357 (O_357,N_9953,N_9878);
nand UO_358 (O_358,N_9489,N_9081);
and UO_359 (O_359,N_9556,N_9732);
nor UO_360 (O_360,N_9652,N_9572);
or UO_361 (O_361,N_9999,N_9027);
and UO_362 (O_362,N_9293,N_9621);
or UO_363 (O_363,N_9827,N_9893);
nand UO_364 (O_364,N_9886,N_9809);
nand UO_365 (O_365,N_9826,N_9672);
and UO_366 (O_366,N_9576,N_9067);
nand UO_367 (O_367,N_9805,N_9422);
nand UO_368 (O_368,N_9327,N_9702);
or UO_369 (O_369,N_9353,N_9985);
or UO_370 (O_370,N_9987,N_9610);
nor UO_371 (O_371,N_9644,N_9390);
and UO_372 (O_372,N_9001,N_9114);
or UO_373 (O_373,N_9332,N_9924);
nor UO_374 (O_374,N_9314,N_9930);
or UO_375 (O_375,N_9706,N_9975);
xnor UO_376 (O_376,N_9806,N_9881);
nor UO_377 (O_377,N_9979,N_9618);
or UO_378 (O_378,N_9955,N_9795);
or UO_379 (O_379,N_9510,N_9734);
nor UO_380 (O_380,N_9935,N_9427);
xor UO_381 (O_381,N_9986,N_9864);
and UO_382 (O_382,N_9889,N_9371);
nand UO_383 (O_383,N_9444,N_9716);
nor UO_384 (O_384,N_9822,N_9876);
nand UO_385 (O_385,N_9954,N_9486);
nor UO_386 (O_386,N_9003,N_9310);
or UO_387 (O_387,N_9565,N_9926);
and UO_388 (O_388,N_9495,N_9907);
and UO_389 (O_389,N_9675,N_9814);
nor UO_390 (O_390,N_9419,N_9337);
nor UO_391 (O_391,N_9857,N_9628);
nor UO_392 (O_392,N_9412,N_9713);
nand UO_393 (O_393,N_9527,N_9236);
or UO_394 (O_394,N_9480,N_9901);
nor UO_395 (O_395,N_9187,N_9558);
nand UO_396 (O_396,N_9742,N_9796);
nor UO_397 (O_397,N_9588,N_9141);
and UO_398 (O_398,N_9746,N_9161);
and UO_399 (O_399,N_9439,N_9058);
nor UO_400 (O_400,N_9997,N_9769);
nor UO_401 (O_401,N_9847,N_9354);
and UO_402 (O_402,N_9219,N_9038);
and UO_403 (O_403,N_9367,N_9966);
nor UO_404 (O_404,N_9049,N_9037);
and UO_405 (O_405,N_9834,N_9179);
or UO_406 (O_406,N_9238,N_9501);
and UO_407 (O_407,N_9903,N_9216);
nor UO_408 (O_408,N_9633,N_9379);
or UO_409 (O_409,N_9057,N_9921);
nand UO_410 (O_410,N_9177,N_9603);
nor UO_411 (O_411,N_9340,N_9465);
or UO_412 (O_412,N_9739,N_9765);
nor UO_413 (O_413,N_9957,N_9816);
nand UO_414 (O_414,N_9068,N_9039);
and UO_415 (O_415,N_9690,N_9181);
nand UO_416 (O_416,N_9741,N_9021);
or UO_417 (O_417,N_9319,N_9532);
or UO_418 (O_418,N_9606,N_9582);
nand UO_419 (O_419,N_9400,N_9380);
or UO_420 (O_420,N_9669,N_9632);
nand UO_421 (O_421,N_9684,N_9388);
or UO_422 (O_422,N_9418,N_9952);
xnor UO_423 (O_423,N_9231,N_9968);
or UO_424 (O_424,N_9232,N_9533);
nand UO_425 (O_425,N_9066,N_9262);
and UO_426 (O_426,N_9749,N_9087);
nand UO_427 (O_427,N_9587,N_9221);
and UO_428 (O_428,N_9993,N_9109);
or UO_429 (O_429,N_9363,N_9929);
nand UO_430 (O_430,N_9469,N_9516);
nand UO_431 (O_431,N_9668,N_9199);
nand UO_432 (O_432,N_9984,N_9240);
and UO_433 (O_433,N_9735,N_9032);
nand UO_434 (O_434,N_9678,N_9945);
and UO_435 (O_435,N_9964,N_9932);
and UO_436 (O_436,N_9853,N_9648);
and UO_437 (O_437,N_9545,N_9515);
nor UO_438 (O_438,N_9031,N_9507);
and UO_439 (O_439,N_9838,N_9775);
and UO_440 (O_440,N_9130,N_9318);
nor UO_441 (O_441,N_9950,N_9869);
nand UO_442 (O_442,N_9478,N_9305);
and UO_443 (O_443,N_9724,N_9551);
nand UO_444 (O_444,N_9336,N_9520);
nand UO_445 (O_445,N_9879,N_9493);
or UO_446 (O_446,N_9408,N_9762);
and UO_447 (O_447,N_9539,N_9271);
nand UO_448 (O_448,N_9791,N_9594);
nand UO_449 (O_449,N_9374,N_9106);
and UO_450 (O_450,N_9898,N_9220);
and UO_451 (O_451,N_9631,N_9218);
nand UO_452 (O_452,N_9281,N_9464);
nor UO_453 (O_453,N_9615,N_9386);
and UO_454 (O_454,N_9833,N_9840);
nor UO_455 (O_455,N_9766,N_9033);
nand UO_456 (O_456,N_9782,N_9339);
nand UO_457 (O_457,N_9645,N_9409);
nand UO_458 (O_458,N_9283,N_9248);
and UO_459 (O_459,N_9485,N_9925);
or UO_460 (O_460,N_9528,N_9282);
and UO_461 (O_461,N_9451,N_9779);
nor UO_462 (O_462,N_9609,N_9020);
nand UO_463 (O_463,N_9210,N_9335);
nand UO_464 (O_464,N_9883,N_9554);
or UO_465 (O_465,N_9387,N_9667);
nor UO_466 (O_466,N_9828,N_9080);
or UO_467 (O_467,N_9413,N_9748);
nor UO_468 (O_468,N_9538,N_9257);
or UO_469 (O_469,N_9234,N_9862);
nand UO_470 (O_470,N_9490,N_9166);
nor UO_471 (O_471,N_9613,N_9799);
nor UO_472 (O_472,N_9105,N_9091);
nand UO_473 (O_473,N_9041,N_9760);
and UO_474 (O_474,N_9433,N_9497);
or UO_475 (O_475,N_9453,N_9036);
nand UO_476 (O_476,N_9297,N_9249);
nand UO_477 (O_477,N_9375,N_9175);
and UO_478 (O_478,N_9346,N_9360);
or UO_479 (O_479,N_9459,N_9322);
or UO_480 (O_480,N_9127,N_9639);
nor UO_481 (O_481,N_9559,N_9909);
nor UO_482 (O_482,N_9665,N_9152);
nand UO_483 (O_483,N_9474,N_9325);
and UO_484 (O_484,N_9347,N_9286);
and UO_485 (O_485,N_9740,N_9237);
or UO_486 (O_486,N_9686,N_9241);
nand UO_487 (O_487,N_9821,N_9173);
and UO_488 (O_488,N_9592,N_9797);
xor UO_489 (O_489,N_9034,N_9943);
or UO_490 (O_490,N_9348,N_9040);
and UO_491 (O_491,N_9919,N_9585);
or UO_492 (O_492,N_9819,N_9342);
and UO_493 (O_493,N_9389,N_9260);
nand UO_494 (O_494,N_9064,N_9266);
and UO_495 (O_495,N_9334,N_9772);
nor UO_496 (O_496,N_9803,N_9736);
and UO_497 (O_497,N_9079,N_9711);
nor UO_498 (O_498,N_9636,N_9264);
and UO_499 (O_499,N_9151,N_9095);
nor UO_500 (O_500,N_9952,N_9597);
and UO_501 (O_501,N_9796,N_9684);
and UO_502 (O_502,N_9932,N_9094);
xnor UO_503 (O_503,N_9159,N_9269);
nand UO_504 (O_504,N_9992,N_9312);
or UO_505 (O_505,N_9524,N_9095);
and UO_506 (O_506,N_9698,N_9309);
and UO_507 (O_507,N_9186,N_9243);
or UO_508 (O_508,N_9333,N_9821);
and UO_509 (O_509,N_9835,N_9473);
or UO_510 (O_510,N_9594,N_9390);
nand UO_511 (O_511,N_9924,N_9667);
nor UO_512 (O_512,N_9038,N_9279);
and UO_513 (O_513,N_9909,N_9711);
and UO_514 (O_514,N_9770,N_9242);
or UO_515 (O_515,N_9362,N_9030);
nor UO_516 (O_516,N_9246,N_9116);
or UO_517 (O_517,N_9921,N_9927);
nor UO_518 (O_518,N_9429,N_9825);
and UO_519 (O_519,N_9437,N_9846);
nand UO_520 (O_520,N_9559,N_9163);
or UO_521 (O_521,N_9052,N_9959);
nand UO_522 (O_522,N_9585,N_9914);
nand UO_523 (O_523,N_9413,N_9737);
nor UO_524 (O_524,N_9378,N_9243);
or UO_525 (O_525,N_9719,N_9701);
or UO_526 (O_526,N_9738,N_9157);
or UO_527 (O_527,N_9941,N_9765);
nor UO_528 (O_528,N_9188,N_9244);
nor UO_529 (O_529,N_9875,N_9264);
nand UO_530 (O_530,N_9761,N_9557);
nand UO_531 (O_531,N_9271,N_9048);
nor UO_532 (O_532,N_9287,N_9985);
or UO_533 (O_533,N_9524,N_9376);
nand UO_534 (O_534,N_9628,N_9960);
nand UO_535 (O_535,N_9316,N_9047);
or UO_536 (O_536,N_9267,N_9795);
and UO_537 (O_537,N_9280,N_9696);
nor UO_538 (O_538,N_9095,N_9871);
nor UO_539 (O_539,N_9673,N_9746);
or UO_540 (O_540,N_9720,N_9784);
or UO_541 (O_541,N_9109,N_9571);
or UO_542 (O_542,N_9441,N_9361);
nand UO_543 (O_543,N_9806,N_9769);
and UO_544 (O_544,N_9457,N_9945);
or UO_545 (O_545,N_9118,N_9568);
and UO_546 (O_546,N_9131,N_9161);
nand UO_547 (O_547,N_9541,N_9534);
nand UO_548 (O_548,N_9712,N_9063);
nand UO_549 (O_549,N_9931,N_9922);
nand UO_550 (O_550,N_9282,N_9502);
nand UO_551 (O_551,N_9683,N_9650);
or UO_552 (O_552,N_9351,N_9922);
nand UO_553 (O_553,N_9582,N_9494);
and UO_554 (O_554,N_9274,N_9410);
or UO_555 (O_555,N_9782,N_9271);
nor UO_556 (O_556,N_9230,N_9697);
or UO_557 (O_557,N_9602,N_9900);
and UO_558 (O_558,N_9358,N_9391);
nor UO_559 (O_559,N_9435,N_9291);
nand UO_560 (O_560,N_9491,N_9247);
nand UO_561 (O_561,N_9857,N_9503);
nand UO_562 (O_562,N_9492,N_9089);
nand UO_563 (O_563,N_9216,N_9576);
or UO_564 (O_564,N_9096,N_9956);
and UO_565 (O_565,N_9511,N_9988);
or UO_566 (O_566,N_9373,N_9244);
and UO_567 (O_567,N_9217,N_9305);
and UO_568 (O_568,N_9895,N_9817);
or UO_569 (O_569,N_9609,N_9408);
or UO_570 (O_570,N_9024,N_9929);
and UO_571 (O_571,N_9372,N_9942);
and UO_572 (O_572,N_9012,N_9726);
nor UO_573 (O_573,N_9520,N_9287);
or UO_574 (O_574,N_9749,N_9083);
or UO_575 (O_575,N_9175,N_9038);
or UO_576 (O_576,N_9172,N_9611);
nand UO_577 (O_577,N_9150,N_9517);
or UO_578 (O_578,N_9271,N_9609);
nor UO_579 (O_579,N_9514,N_9168);
nor UO_580 (O_580,N_9251,N_9194);
and UO_581 (O_581,N_9058,N_9920);
and UO_582 (O_582,N_9528,N_9559);
or UO_583 (O_583,N_9304,N_9700);
or UO_584 (O_584,N_9167,N_9930);
and UO_585 (O_585,N_9153,N_9802);
and UO_586 (O_586,N_9750,N_9211);
nand UO_587 (O_587,N_9507,N_9711);
and UO_588 (O_588,N_9507,N_9120);
nand UO_589 (O_589,N_9006,N_9277);
and UO_590 (O_590,N_9860,N_9533);
nand UO_591 (O_591,N_9027,N_9419);
and UO_592 (O_592,N_9639,N_9229);
and UO_593 (O_593,N_9544,N_9232);
nor UO_594 (O_594,N_9123,N_9324);
or UO_595 (O_595,N_9738,N_9371);
nor UO_596 (O_596,N_9268,N_9155);
and UO_597 (O_597,N_9404,N_9436);
and UO_598 (O_598,N_9106,N_9428);
and UO_599 (O_599,N_9417,N_9548);
nand UO_600 (O_600,N_9314,N_9682);
nor UO_601 (O_601,N_9422,N_9892);
nor UO_602 (O_602,N_9515,N_9585);
nor UO_603 (O_603,N_9869,N_9817);
or UO_604 (O_604,N_9198,N_9390);
and UO_605 (O_605,N_9912,N_9972);
or UO_606 (O_606,N_9025,N_9372);
nor UO_607 (O_607,N_9779,N_9065);
and UO_608 (O_608,N_9457,N_9188);
nand UO_609 (O_609,N_9241,N_9404);
nand UO_610 (O_610,N_9316,N_9936);
and UO_611 (O_611,N_9516,N_9193);
xor UO_612 (O_612,N_9149,N_9560);
nor UO_613 (O_613,N_9904,N_9976);
or UO_614 (O_614,N_9686,N_9584);
or UO_615 (O_615,N_9615,N_9586);
nor UO_616 (O_616,N_9123,N_9831);
nor UO_617 (O_617,N_9587,N_9013);
nor UO_618 (O_618,N_9724,N_9648);
and UO_619 (O_619,N_9682,N_9528);
or UO_620 (O_620,N_9869,N_9043);
nand UO_621 (O_621,N_9065,N_9497);
nand UO_622 (O_622,N_9785,N_9376);
nor UO_623 (O_623,N_9677,N_9666);
nor UO_624 (O_624,N_9455,N_9659);
and UO_625 (O_625,N_9352,N_9118);
nand UO_626 (O_626,N_9214,N_9613);
or UO_627 (O_627,N_9099,N_9754);
nor UO_628 (O_628,N_9482,N_9958);
and UO_629 (O_629,N_9615,N_9735);
or UO_630 (O_630,N_9436,N_9149);
or UO_631 (O_631,N_9904,N_9486);
nor UO_632 (O_632,N_9878,N_9234);
or UO_633 (O_633,N_9813,N_9810);
nor UO_634 (O_634,N_9261,N_9132);
or UO_635 (O_635,N_9902,N_9150);
nand UO_636 (O_636,N_9022,N_9372);
or UO_637 (O_637,N_9074,N_9104);
and UO_638 (O_638,N_9598,N_9508);
and UO_639 (O_639,N_9904,N_9468);
or UO_640 (O_640,N_9985,N_9836);
or UO_641 (O_641,N_9773,N_9734);
or UO_642 (O_642,N_9345,N_9390);
nand UO_643 (O_643,N_9437,N_9767);
and UO_644 (O_644,N_9766,N_9291);
and UO_645 (O_645,N_9136,N_9837);
nand UO_646 (O_646,N_9808,N_9580);
nor UO_647 (O_647,N_9457,N_9900);
nand UO_648 (O_648,N_9800,N_9223);
or UO_649 (O_649,N_9309,N_9073);
nor UO_650 (O_650,N_9197,N_9081);
nand UO_651 (O_651,N_9313,N_9972);
and UO_652 (O_652,N_9409,N_9674);
and UO_653 (O_653,N_9543,N_9492);
or UO_654 (O_654,N_9710,N_9392);
nor UO_655 (O_655,N_9012,N_9413);
and UO_656 (O_656,N_9886,N_9642);
and UO_657 (O_657,N_9971,N_9796);
nor UO_658 (O_658,N_9378,N_9531);
and UO_659 (O_659,N_9003,N_9470);
nand UO_660 (O_660,N_9268,N_9699);
nor UO_661 (O_661,N_9024,N_9346);
or UO_662 (O_662,N_9921,N_9846);
nand UO_663 (O_663,N_9983,N_9045);
nor UO_664 (O_664,N_9564,N_9126);
or UO_665 (O_665,N_9817,N_9709);
xor UO_666 (O_666,N_9541,N_9976);
nor UO_667 (O_667,N_9591,N_9366);
and UO_668 (O_668,N_9293,N_9915);
or UO_669 (O_669,N_9020,N_9373);
or UO_670 (O_670,N_9221,N_9358);
nor UO_671 (O_671,N_9910,N_9366);
or UO_672 (O_672,N_9543,N_9471);
and UO_673 (O_673,N_9477,N_9937);
and UO_674 (O_674,N_9214,N_9229);
and UO_675 (O_675,N_9148,N_9829);
and UO_676 (O_676,N_9527,N_9970);
nor UO_677 (O_677,N_9879,N_9133);
or UO_678 (O_678,N_9044,N_9013);
nand UO_679 (O_679,N_9190,N_9246);
nand UO_680 (O_680,N_9552,N_9884);
nor UO_681 (O_681,N_9226,N_9117);
nor UO_682 (O_682,N_9865,N_9473);
nand UO_683 (O_683,N_9181,N_9763);
or UO_684 (O_684,N_9057,N_9337);
or UO_685 (O_685,N_9319,N_9081);
nor UO_686 (O_686,N_9147,N_9650);
nor UO_687 (O_687,N_9451,N_9260);
or UO_688 (O_688,N_9449,N_9320);
and UO_689 (O_689,N_9692,N_9644);
nor UO_690 (O_690,N_9633,N_9304);
nand UO_691 (O_691,N_9223,N_9592);
nor UO_692 (O_692,N_9234,N_9392);
nand UO_693 (O_693,N_9934,N_9207);
and UO_694 (O_694,N_9710,N_9329);
xnor UO_695 (O_695,N_9512,N_9948);
nor UO_696 (O_696,N_9766,N_9991);
xor UO_697 (O_697,N_9365,N_9051);
and UO_698 (O_698,N_9110,N_9692);
and UO_699 (O_699,N_9146,N_9819);
nor UO_700 (O_700,N_9852,N_9748);
and UO_701 (O_701,N_9818,N_9056);
or UO_702 (O_702,N_9524,N_9071);
nand UO_703 (O_703,N_9039,N_9121);
nand UO_704 (O_704,N_9170,N_9885);
and UO_705 (O_705,N_9190,N_9626);
nor UO_706 (O_706,N_9493,N_9119);
or UO_707 (O_707,N_9576,N_9812);
nor UO_708 (O_708,N_9922,N_9361);
and UO_709 (O_709,N_9581,N_9034);
and UO_710 (O_710,N_9091,N_9894);
or UO_711 (O_711,N_9429,N_9786);
nor UO_712 (O_712,N_9074,N_9057);
nor UO_713 (O_713,N_9245,N_9611);
or UO_714 (O_714,N_9222,N_9395);
or UO_715 (O_715,N_9481,N_9663);
or UO_716 (O_716,N_9871,N_9965);
nor UO_717 (O_717,N_9353,N_9817);
nand UO_718 (O_718,N_9933,N_9552);
nand UO_719 (O_719,N_9876,N_9035);
or UO_720 (O_720,N_9097,N_9489);
nand UO_721 (O_721,N_9675,N_9683);
nor UO_722 (O_722,N_9277,N_9387);
nand UO_723 (O_723,N_9695,N_9427);
or UO_724 (O_724,N_9805,N_9864);
nand UO_725 (O_725,N_9651,N_9421);
nor UO_726 (O_726,N_9046,N_9986);
nand UO_727 (O_727,N_9033,N_9135);
nor UO_728 (O_728,N_9829,N_9143);
or UO_729 (O_729,N_9294,N_9531);
nand UO_730 (O_730,N_9698,N_9891);
and UO_731 (O_731,N_9498,N_9896);
nor UO_732 (O_732,N_9262,N_9330);
and UO_733 (O_733,N_9408,N_9009);
or UO_734 (O_734,N_9436,N_9727);
nand UO_735 (O_735,N_9601,N_9094);
nor UO_736 (O_736,N_9035,N_9936);
or UO_737 (O_737,N_9317,N_9489);
and UO_738 (O_738,N_9802,N_9065);
and UO_739 (O_739,N_9199,N_9055);
or UO_740 (O_740,N_9363,N_9037);
and UO_741 (O_741,N_9676,N_9397);
nor UO_742 (O_742,N_9293,N_9077);
nand UO_743 (O_743,N_9838,N_9691);
and UO_744 (O_744,N_9814,N_9844);
nand UO_745 (O_745,N_9835,N_9952);
nand UO_746 (O_746,N_9650,N_9536);
nor UO_747 (O_747,N_9675,N_9046);
or UO_748 (O_748,N_9377,N_9363);
nor UO_749 (O_749,N_9027,N_9895);
nor UO_750 (O_750,N_9173,N_9934);
and UO_751 (O_751,N_9040,N_9556);
nand UO_752 (O_752,N_9315,N_9746);
or UO_753 (O_753,N_9657,N_9610);
nand UO_754 (O_754,N_9955,N_9894);
nor UO_755 (O_755,N_9031,N_9522);
nand UO_756 (O_756,N_9461,N_9995);
and UO_757 (O_757,N_9669,N_9347);
nor UO_758 (O_758,N_9160,N_9144);
or UO_759 (O_759,N_9023,N_9941);
nand UO_760 (O_760,N_9855,N_9542);
nor UO_761 (O_761,N_9504,N_9827);
nand UO_762 (O_762,N_9128,N_9025);
and UO_763 (O_763,N_9889,N_9245);
or UO_764 (O_764,N_9264,N_9253);
and UO_765 (O_765,N_9323,N_9664);
and UO_766 (O_766,N_9608,N_9702);
nor UO_767 (O_767,N_9792,N_9489);
nor UO_768 (O_768,N_9235,N_9277);
or UO_769 (O_769,N_9396,N_9770);
nand UO_770 (O_770,N_9543,N_9358);
nor UO_771 (O_771,N_9008,N_9708);
and UO_772 (O_772,N_9850,N_9711);
and UO_773 (O_773,N_9640,N_9445);
and UO_774 (O_774,N_9071,N_9965);
and UO_775 (O_775,N_9733,N_9116);
and UO_776 (O_776,N_9652,N_9515);
nand UO_777 (O_777,N_9615,N_9555);
nor UO_778 (O_778,N_9996,N_9568);
or UO_779 (O_779,N_9512,N_9720);
nor UO_780 (O_780,N_9643,N_9142);
nand UO_781 (O_781,N_9975,N_9663);
and UO_782 (O_782,N_9635,N_9143);
or UO_783 (O_783,N_9251,N_9613);
and UO_784 (O_784,N_9824,N_9639);
nand UO_785 (O_785,N_9465,N_9143);
or UO_786 (O_786,N_9655,N_9417);
nor UO_787 (O_787,N_9104,N_9035);
or UO_788 (O_788,N_9945,N_9047);
nand UO_789 (O_789,N_9726,N_9823);
nand UO_790 (O_790,N_9609,N_9040);
nand UO_791 (O_791,N_9431,N_9162);
or UO_792 (O_792,N_9926,N_9200);
or UO_793 (O_793,N_9299,N_9610);
nor UO_794 (O_794,N_9421,N_9545);
or UO_795 (O_795,N_9698,N_9530);
nand UO_796 (O_796,N_9627,N_9605);
nand UO_797 (O_797,N_9962,N_9226);
and UO_798 (O_798,N_9560,N_9240);
nand UO_799 (O_799,N_9855,N_9835);
or UO_800 (O_800,N_9066,N_9475);
nor UO_801 (O_801,N_9143,N_9921);
nor UO_802 (O_802,N_9106,N_9104);
nor UO_803 (O_803,N_9619,N_9805);
nor UO_804 (O_804,N_9183,N_9219);
and UO_805 (O_805,N_9790,N_9161);
or UO_806 (O_806,N_9587,N_9970);
or UO_807 (O_807,N_9871,N_9250);
and UO_808 (O_808,N_9432,N_9681);
xnor UO_809 (O_809,N_9367,N_9526);
nor UO_810 (O_810,N_9967,N_9212);
and UO_811 (O_811,N_9897,N_9088);
or UO_812 (O_812,N_9188,N_9736);
nand UO_813 (O_813,N_9866,N_9045);
nand UO_814 (O_814,N_9345,N_9289);
nand UO_815 (O_815,N_9466,N_9677);
and UO_816 (O_816,N_9759,N_9883);
or UO_817 (O_817,N_9047,N_9386);
and UO_818 (O_818,N_9094,N_9762);
or UO_819 (O_819,N_9584,N_9504);
nand UO_820 (O_820,N_9563,N_9556);
or UO_821 (O_821,N_9202,N_9829);
or UO_822 (O_822,N_9612,N_9192);
and UO_823 (O_823,N_9478,N_9725);
and UO_824 (O_824,N_9945,N_9249);
nand UO_825 (O_825,N_9388,N_9662);
or UO_826 (O_826,N_9666,N_9082);
nor UO_827 (O_827,N_9067,N_9704);
nand UO_828 (O_828,N_9646,N_9523);
or UO_829 (O_829,N_9785,N_9965);
and UO_830 (O_830,N_9861,N_9417);
nand UO_831 (O_831,N_9456,N_9347);
nand UO_832 (O_832,N_9026,N_9771);
or UO_833 (O_833,N_9440,N_9835);
or UO_834 (O_834,N_9249,N_9566);
and UO_835 (O_835,N_9219,N_9737);
and UO_836 (O_836,N_9041,N_9878);
and UO_837 (O_837,N_9796,N_9818);
nand UO_838 (O_838,N_9005,N_9041);
nor UO_839 (O_839,N_9036,N_9422);
nand UO_840 (O_840,N_9205,N_9258);
and UO_841 (O_841,N_9979,N_9427);
nor UO_842 (O_842,N_9357,N_9102);
nand UO_843 (O_843,N_9258,N_9609);
xnor UO_844 (O_844,N_9878,N_9290);
or UO_845 (O_845,N_9738,N_9519);
and UO_846 (O_846,N_9321,N_9264);
nor UO_847 (O_847,N_9183,N_9675);
and UO_848 (O_848,N_9933,N_9715);
and UO_849 (O_849,N_9797,N_9514);
nand UO_850 (O_850,N_9335,N_9347);
and UO_851 (O_851,N_9038,N_9330);
nor UO_852 (O_852,N_9607,N_9405);
and UO_853 (O_853,N_9683,N_9325);
nand UO_854 (O_854,N_9380,N_9433);
and UO_855 (O_855,N_9872,N_9975);
or UO_856 (O_856,N_9597,N_9250);
or UO_857 (O_857,N_9705,N_9744);
or UO_858 (O_858,N_9909,N_9137);
or UO_859 (O_859,N_9823,N_9007);
nand UO_860 (O_860,N_9830,N_9453);
nand UO_861 (O_861,N_9604,N_9419);
or UO_862 (O_862,N_9966,N_9872);
nor UO_863 (O_863,N_9541,N_9249);
and UO_864 (O_864,N_9413,N_9802);
or UO_865 (O_865,N_9876,N_9111);
and UO_866 (O_866,N_9138,N_9325);
nand UO_867 (O_867,N_9465,N_9079);
and UO_868 (O_868,N_9726,N_9683);
and UO_869 (O_869,N_9564,N_9059);
nand UO_870 (O_870,N_9699,N_9226);
and UO_871 (O_871,N_9308,N_9212);
and UO_872 (O_872,N_9270,N_9092);
and UO_873 (O_873,N_9781,N_9892);
or UO_874 (O_874,N_9850,N_9804);
and UO_875 (O_875,N_9452,N_9403);
or UO_876 (O_876,N_9231,N_9948);
or UO_877 (O_877,N_9458,N_9789);
and UO_878 (O_878,N_9516,N_9610);
and UO_879 (O_879,N_9508,N_9736);
or UO_880 (O_880,N_9081,N_9823);
and UO_881 (O_881,N_9216,N_9391);
and UO_882 (O_882,N_9621,N_9816);
and UO_883 (O_883,N_9843,N_9830);
nand UO_884 (O_884,N_9730,N_9020);
or UO_885 (O_885,N_9782,N_9958);
nand UO_886 (O_886,N_9893,N_9193);
nand UO_887 (O_887,N_9025,N_9804);
and UO_888 (O_888,N_9051,N_9154);
or UO_889 (O_889,N_9436,N_9539);
nor UO_890 (O_890,N_9012,N_9004);
nor UO_891 (O_891,N_9063,N_9428);
nor UO_892 (O_892,N_9377,N_9972);
and UO_893 (O_893,N_9351,N_9793);
and UO_894 (O_894,N_9061,N_9368);
and UO_895 (O_895,N_9053,N_9026);
nor UO_896 (O_896,N_9642,N_9937);
nand UO_897 (O_897,N_9336,N_9139);
nand UO_898 (O_898,N_9105,N_9005);
and UO_899 (O_899,N_9470,N_9127);
and UO_900 (O_900,N_9971,N_9062);
nor UO_901 (O_901,N_9709,N_9706);
nor UO_902 (O_902,N_9392,N_9509);
nor UO_903 (O_903,N_9808,N_9335);
and UO_904 (O_904,N_9262,N_9780);
nor UO_905 (O_905,N_9323,N_9455);
and UO_906 (O_906,N_9858,N_9069);
nand UO_907 (O_907,N_9334,N_9462);
and UO_908 (O_908,N_9773,N_9927);
nor UO_909 (O_909,N_9196,N_9159);
nor UO_910 (O_910,N_9077,N_9597);
nor UO_911 (O_911,N_9104,N_9642);
and UO_912 (O_912,N_9828,N_9873);
and UO_913 (O_913,N_9322,N_9885);
or UO_914 (O_914,N_9432,N_9566);
nor UO_915 (O_915,N_9204,N_9412);
nor UO_916 (O_916,N_9441,N_9261);
or UO_917 (O_917,N_9759,N_9982);
nor UO_918 (O_918,N_9486,N_9656);
or UO_919 (O_919,N_9747,N_9133);
or UO_920 (O_920,N_9280,N_9439);
xnor UO_921 (O_921,N_9286,N_9793);
and UO_922 (O_922,N_9677,N_9210);
and UO_923 (O_923,N_9044,N_9149);
or UO_924 (O_924,N_9740,N_9415);
nand UO_925 (O_925,N_9353,N_9674);
nor UO_926 (O_926,N_9999,N_9030);
xnor UO_927 (O_927,N_9740,N_9580);
or UO_928 (O_928,N_9608,N_9121);
and UO_929 (O_929,N_9600,N_9189);
nand UO_930 (O_930,N_9581,N_9316);
or UO_931 (O_931,N_9024,N_9882);
or UO_932 (O_932,N_9311,N_9138);
nor UO_933 (O_933,N_9219,N_9927);
or UO_934 (O_934,N_9847,N_9983);
nor UO_935 (O_935,N_9707,N_9540);
xnor UO_936 (O_936,N_9683,N_9472);
nand UO_937 (O_937,N_9809,N_9953);
or UO_938 (O_938,N_9390,N_9292);
nor UO_939 (O_939,N_9862,N_9385);
and UO_940 (O_940,N_9421,N_9707);
nand UO_941 (O_941,N_9103,N_9316);
nor UO_942 (O_942,N_9676,N_9420);
nand UO_943 (O_943,N_9311,N_9275);
nand UO_944 (O_944,N_9321,N_9512);
or UO_945 (O_945,N_9611,N_9334);
nand UO_946 (O_946,N_9536,N_9970);
nand UO_947 (O_947,N_9520,N_9066);
or UO_948 (O_948,N_9522,N_9419);
nor UO_949 (O_949,N_9757,N_9382);
nand UO_950 (O_950,N_9761,N_9043);
and UO_951 (O_951,N_9905,N_9715);
nor UO_952 (O_952,N_9275,N_9721);
nand UO_953 (O_953,N_9222,N_9788);
and UO_954 (O_954,N_9222,N_9343);
nand UO_955 (O_955,N_9725,N_9297);
nand UO_956 (O_956,N_9617,N_9439);
nand UO_957 (O_957,N_9364,N_9091);
and UO_958 (O_958,N_9073,N_9166);
nand UO_959 (O_959,N_9032,N_9262);
and UO_960 (O_960,N_9265,N_9756);
nand UO_961 (O_961,N_9024,N_9235);
nand UO_962 (O_962,N_9006,N_9730);
nand UO_963 (O_963,N_9688,N_9496);
and UO_964 (O_964,N_9629,N_9565);
nor UO_965 (O_965,N_9035,N_9620);
nor UO_966 (O_966,N_9961,N_9363);
and UO_967 (O_967,N_9663,N_9459);
and UO_968 (O_968,N_9479,N_9767);
and UO_969 (O_969,N_9090,N_9314);
or UO_970 (O_970,N_9221,N_9688);
xor UO_971 (O_971,N_9751,N_9489);
nand UO_972 (O_972,N_9563,N_9776);
and UO_973 (O_973,N_9352,N_9185);
or UO_974 (O_974,N_9103,N_9489);
and UO_975 (O_975,N_9295,N_9252);
xnor UO_976 (O_976,N_9757,N_9738);
and UO_977 (O_977,N_9473,N_9739);
or UO_978 (O_978,N_9751,N_9019);
xor UO_979 (O_979,N_9576,N_9910);
nor UO_980 (O_980,N_9387,N_9099);
nor UO_981 (O_981,N_9141,N_9707);
and UO_982 (O_982,N_9204,N_9926);
and UO_983 (O_983,N_9926,N_9478);
and UO_984 (O_984,N_9840,N_9808);
nor UO_985 (O_985,N_9303,N_9249);
nor UO_986 (O_986,N_9576,N_9818);
nor UO_987 (O_987,N_9721,N_9994);
nor UO_988 (O_988,N_9459,N_9782);
and UO_989 (O_989,N_9771,N_9179);
or UO_990 (O_990,N_9861,N_9995);
or UO_991 (O_991,N_9487,N_9605);
or UO_992 (O_992,N_9311,N_9935);
or UO_993 (O_993,N_9686,N_9277);
nand UO_994 (O_994,N_9163,N_9214);
nand UO_995 (O_995,N_9324,N_9491);
or UO_996 (O_996,N_9505,N_9003);
and UO_997 (O_997,N_9553,N_9514);
or UO_998 (O_998,N_9819,N_9984);
nor UO_999 (O_999,N_9648,N_9992);
or UO_1000 (O_1000,N_9304,N_9951);
or UO_1001 (O_1001,N_9011,N_9022);
nor UO_1002 (O_1002,N_9822,N_9054);
or UO_1003 (O_1003,N_9797,N_9121);
and UO_1004 (O_1004,N_9444,N_9481);
nor UO_1005 (O_1005,N_9744,N_9460);
nor UO_1006 (O_1006,N_9011,N_9080);
nand UO_1007 (O_1007,N_9752,N_9774);
nand UO_1008 (O_1008,N_9294,N_9126);
nand UO_1009 (O_1009,N_9137,N_9260);
nand UO_1010 (O_1010,N_9876,N_9759);
or UO_1011 (O_1011,N_9760,N_9681);
nor UO_1012 (O_1012,N_9727,N_9692);
xnor UO_1013 (O_1013,N_9931,N_9849);
nand UO_1014 (O_1014,N_9054,N_9191);
and UO_1015 (O_1015,N_9117,N_9399);
and UO_1016 (O_1016,N_9070,N_9241);
nand UO_1017 (O_1017,N_9855,N_9000);
nand UO_1018 (O_1018,N_9256,N_9675);
or UO_1019 (O_1019,N_9932,N_9488);
and UO_1020 (O_1020,N_9963,N_9409);
nor UO_1021 (O_1021,N_9769,N_9962);
or UO_1022 (O_1022,N_9777,N_9752);
xnor UO_1023 (O_1023,N_9784,N_9944);
or UO_1024 (O_1024,N_9308,N_9808);
nor UO_1025 (O_1025,N_9796,N_9998);
or UO_1026 (O_1026,N_9514,N_9681);
nor UO_1027 (O_1027,N_9843,N_9026);
and UO_1028 (O_1028,N_9540,N_9081);
or UO_1029 (O_1029,N_9216,N_9302);
and UO_1030 (O_1030,N_9828,N_9491);
nand UO_1031 (O_1031,N_9437,N_9611);
nand UO_1032 (O_1032,N_9694,N_9595);
nand UO_1033 (O_1033,N_9591,N_9921);
and UO_1034 (O_1034,N_9708,N_9439);
or UO_1035 (O_1035,N_9343,N_9931);
and UO_1036 (O_1036,N_9355,N_9386);
or UO_1037 (O_1037,N_9993,N_9265);
or UO_1038 (O_1038,N_9221,N_9637);
nor UO_1039 (O_1039,N_9014,N_9994);
and UO_1040 (O_1040,N_9059,N_9686);
nor UO_1041 (O_1041,N_9015,N_9694);
nor UO_1042 (O_1042,N_9141,N_9933);
nor UO_1043 (O_1043,N_9866,N_9177);
or UO_1044 (O_1044,N_9096,N_9734);
or UO_1045 (O_1045,N_9966,N_9571);
or UO_1046 (O_1046,N_9711,N_9642);
and UO_1047 (O_1047,N_9600,N_9440);
or UO_1048 (O_1048,N_9998,N_9342);
nand UO_1049 (O_1049,N_9077,N_9671);
nand UO_1050 (O_1050,N_9537,N_9698);
nand UO_1051 (O_1051,N_9253,N_9090);
nor UO_1052 (O_1052,N_9741,N_9676);
and UO_1053 (O_1053,N_9717,N_9774);
nor UO_1054 (O_1054,N_9562,N_9989);
nand UO_1055 (O_1055,N_9696,N_9716);
nand UO_1056 (O_1056,N_9036,N_9273);
nand UO_1057 (O_1057,N_9738,N_9366);
or UO_1058 (O_1058,N_9118,N_9521);
nor UO_1059 (O_1059,N_9653,N_9013);
or UO_1060 (O_1060,N_9697,N_9426);
nor UO_1061 (O_1061,N_9367,N_9490);
nand UO_1062 (O_1062,N_9865,N_9053);
and UO_1063 (O_1063,N_9631,N_9871);
and UO_1064 (O_1064,N_9579,N_9835);
nor UO_1065 (O_1065,N_9913,N_9902);
and UO_1066 (O_1066,N_9819,N_9530);
nand UO_1067 (O_1067,N_9457,N_9498);
and UO_1068 (O_1068,N_9328,N_9545);
nand UO_1069 (O_1069,N_9573,N_9401);
and UO_1070 (O_1070,N_9183,N_9970);
nor UO_1071 (O_1071,N_9854,N_9625);
nand UO_1072 (O_1072,N_9984,N_9677);
nor UO_1073 (O_1073,N_9078,N_9913);
or UO_1074 (O_1074,N_9415,N_9187);
nor UO_1075 (O_1075,N_9186,N_9622);
or UO_1076 (O_1076,N_9055,N_9761);
and UO_1077 (O_1077,N_9628,N_9615);
nand UO_1078 (O_1078,N_9428,N_9389);
and UO_1079 (O_1079,N_9810,N_9297);
nor UO_1080 (O_1080,N_9237,N_9466);
and UO_1081 (O_1081,N_9949,N_9145);
or UO_1082 (O_1082,N_9222,N_9096);
nor UO_1083 (O_1083,N_9715,N_9030);
nand UO_1084 (O_1084,N_9679,N_9176);
or UO_1085 (O_1085,N_9275,N_9625);
nor UO_1086 (O_1086,N_9250,N_9780);
and UO_1087 (O_1087,N_9970,N_9197);
or UO_1088 (O_1088,N_9906,N_9097);
nand UO_1089 (O_1089,N_9244,N_9393);
or UO_1090 (O_1090,N_9460,N_9555);
nor UO_1091 (O_1091,N_9648,N_9219);
nand UO_1092 (O_1092,N_9759,N_9964);
or UO_1093 (O_1093,N_9703,N_9601);
and UO_1094 (O_1094,N_9095,N_9941);
nand UO_1095 (O_1095,N_9869,N_9515);
and UO_1096 (O_1096,N_9555,N_9126);
and UO_1097 (O_1097,N_9789,N_9411);
and UO_1098 (O_1098,N_9377,N_9638);
nand UO_1099 (O_1099,N_9597,N_9755);
nand UO_1100 (O_1100,N_9569,N_9555);
nand UO_1101 (O_1101,N_9005,N_9841);
or UO_1102 (O_1102,N_9927,N_9098);
nor UO_1103 (O_1103,N_9705,N_9666);
or UO_1104 (O_1104,N_9881,N_9610);
nor UO_1105 (O_1105,N_9254,N_9582);
nor UO_1106 (O_1106,N_9987,N_9051);
nor UO_1107 (O_1107,N_9795,N_9299);
nand UO_1108 (O_1108,N_9300,N_9629);
nor UO_1109 (O_1109,N_9277,N_9096);
or UO_1110 (O_1110,N_9641,N_9089);
nor UO_1111 (O_1111,N_9820,N_9375);
nand UO_1112 (O_1112,N_9659,N_9560);
and UO_1113 (O_1113,N_9213,N_9607);
nand UO_1114 (O_1114,N_9097,N_9685);
xnor UO_1115 (O_1115,N_9337,N_9392);
nor UO_1116 (O_1116,N_9239,N_9937);
or UO_1117 (O_1117,N_9731,N_9626);
and UO_1118 (O_1118,N_9327,N_9066);
or UO_1119 (O_1119,N_9206,N_9690);
xnor UO_1120 (O_1120,N_9949,N_9500);
nor UO_1121 (O_1121,N_9746,N_9743);
nand UO_1122 (O_1122,N_9542,N_9671);
or UO_1123 (O_1123,N_9034,N_9545);
and UO_1124 (O_1124,N_9239,N_9764);
and UO_1125 (O_1125,N_9024,N_9059);
nor UO_1126 (O_1126,N_9573,N_9077);
or UO_1127 (O_1127,N_9503,N_9556);
nor UO_1128 (O_1128,N_9498,N_9156);
and UO_1129 (O_1129,N_9667,N_9193);
nand UO_1130 (O_1130,N_9284,N_9973);
nor UO_1131 (O_1131,N_9592,N_9212);
or UO_1132 (O_1132,N_9260,N_9029);
or UO_1133 (O_1133,N_9344,N_9275);
or UO_1134 (O_1134,N_9225,N_9344);
and UO_1135 (O_1135,N_9948,N_9091);
or UO_1136 (O_1136,N_9870,N_9767);
and UO_1137 (O_1137,N_9354,N_9363);
nand UO_1138 (O_1138,N_9128,N_9567);
and UO_1139 (O_1139,N_9962,N_9828);
or UO_1140 (O_1140,N_9000,N_9111);
nand UO_1141 (O_1141,N_9318,N_9164);
nand UO_1142 (O_1142,N_9758,N_9866);
nand UO_1143 (O_1143,N_9669,N_9865);
nand UO_1144 (O_1144,N_9026,N_9700);
nor UO_1145 (O_1145,N_9888,N_9840);
or UO_1146 (O_1146,N_9232,N_9435);
nand UO_1147 (O_1147,N_9977,N_9065);
or UO_1148 (O_1148,N_9423,N_9277);
and UO_1149 (O_1149,N_9704,N_9110);
nand UO_1150 (O_1150,N_9124,N_9256);
nand UO_1151 (O_1151,N_9834,N_9449);
nor UO_1152 (O_1152,N_9063,N_9385);
or UO_1153 (O_1153,N_9320,N_9745);
nand UO_1154 (O_1154,N_9349,N_9854);
and UO_1155 (O_1155,N_9284,N_9213);
or UO_1156 (O_1156,N_9121,N_9038);
or UO_1157 (O_1157,N_9302,N_9990);
and UO_1158 (O_1158,N_9339,N_9832);
and UO_1159 (O_1159,N_9643,N_9088);
and UO_1160 (O_1160,N_9548,N_9561);
or UO_1161 (O_1161,N_9346,N_9858);
nor UO_1162 (O_1162,N_9339,N_9134);
or UO_1163 (O_1163,N_9623,N_9762);
and UO_1164 (O_1164,N_9752,N_9265);
or UO_1165 (O_1165,N_9351,N_9045);
nand UO_1166 (O_1166,N_9145,N_9979);
nor UO_1167 (O_1167,N_9345,N_9445);
nand UO_1168 (O_1168,N_9662,N_9414);
nor UO_1169 (O_1169,N_9592,N_9977);
xnor UO_1170 (O_1170,N_9840,N_9425);
nand UO_1171 (O_1171,N_9648,N_9772);
or UO_1172 (O_1172,N_9957,N_9080);
nor UO_1173 (O_1173,N_9786,N_9718);
nand UO_1174 (O_1174,N_9765,N_9867);
and UO_1175 (O_1175,N_9077,N_9303);
and UO_1176 (O_1176,N_9449,N_9289);
and UO_1177 (O_1177,N_9993,N_9719);
nand UO_1178 (O_1178,N_9464,N_9330);
or UO_1179 (O_1179,N_9093,N_9203);
xor UO_1180 (O_1180,N_9271,N_9702);
nand UO_1181 (O_1181,N_9327,N_9887);
or UO_1182 (O_1182,N_9161,N_9459);
nor UO_1183 (O_1183,N_9040,N_9504);
and UO_1184 (O_1184,N_9091,N_9945);
nand UO_1185 (O_1185,N_9663,N_9124);
and UO_1186 (O_1186,N_9955,N_9683);
nor UO_1187 (O_1187,N_9975,N_9931);
nand UO_1188 (O_1188,N_9519,N_9459);
nand UO_1189 (O_1189,N_9089,N_9820);
nand UO_1190 (O_1190,N_9476,N_9870);
nand UO_1191 (O_1191,N_9634,N_9057);
or UO_1192 (O_1192,N_9582,N_9554);
and UO_1193 (O_1193,N_9502,N_9012);
or UO_1194 (O_1194,N_9568,N_9375);
or UO_1195 (O_1195,N_9630,N_9767);
or UO_1196 (O_1196,N_9650,N_9295);
or UO_1197 (O_1197,N_9029,N_9882);
or UO_1198 (O_1198,N_9051,N_9765);
nor UO_1199 (O_1199,N_9918,N_9021);
nor UO_1200 (O_1200,N_9079,N_9945);
nor UO_1201 (O_1201,N_9436,N_9431);
nand UO_1202 (O_1202,N_9971,N_9665);
and UO_1203 (O_1203,N_9652,N_9777);
or UO_1204 (O_1204,N_9615,N_9823);
and UO_1205 (O_1205,N_9821,N_9597);
nand UO_1206 (O_1206,N_9204,N_9915);
and UO_1207 (O_1207,N_9567,N_9683);
nor UO_1208 (O_1208,N_9222,N_9540);
xor UO_1209 (O_1209,N_9249,N_9512);
nor UO_1210 (O_1210,N_9697,N_9761);
and UO_1211 (O_1211,N_9483,N_9899);
nand UO_1212 (O_1212,N_9976,N_9744);
or UO_1213 (O_1213,N_9323,N_9317);
and UO_1214 (O_1214,N_9483,N_9684);
or UO_1215 (O_1215,N_9868,N_9720);
and UO_1216 (O_1216,N_9995,N_9773);
nand UO_1217 (O_1217,N_9449,N_9266);
nand UO_1218 (O_1218,N_9272,N_9069);
nor UO_1219 (O_1219,N_9492,N_9676);
or UO_1220 (O_1220,N_9490,N_9720);
or UO_1221 (O_1221,N_9313,N_9487);
and UO_1222 (O_1222,N_9476,N_9009);
or UO_1223 (O_1223,N_9097,N_9393);
nor UO_1224 (O_1224,N_9663,N_9520);
nand UO_1225 (O_1225,N_9058,N_9803);
nor UO_1226 (O_1226,N_9121,N_9094);
or UO_1227 (O_1227,N_9580,N_9825);
nor UO_1228 (O_1228,N_9965,N_9686);
nand UO_1229 (O_1229,N_9297,N_9873);
nor UO_1230 (O_1230,N_9678,N_9684);
nand UO_1231 (O_1231,N_9054,N_9074);
or UO_1232 (O_1232,N_9513,N_9542);
or UO_1233 (O_1233,N_9861,N_9352);
nand UO_1234 (O_1234,N_9854,N_9476);
xnor UO_1235 (O_1235,N_9573,N_9052);
nand UO_1236 (O_1236,N_9623,N_9485);
nand UO_1237 (O_1237,N_9370,N_9101);
xor UO_1238 (O_1238,N_9696,N_9339);
or UO_1239 (O_1239,N_9292,N_9250);
or UO_1240 (O_1240,N_9267,N_9801);
nand UO_1241 (O_1241,N_9888,N_9259);
and UO_1242 (O_1242,N_9616,N_9127);
or UO_1243 (O_1243,N_9394,N_9203);
or UO_1244 (O_1244,N_9506,N_9155);
xnor UO_1245 (O_1245,N_9162,N_9789);
nor UO_1246 (O_1246,N_9199,N_9482);
and UO_1247 (O_1247,N_9956,N_9421);
nor UO_1248 (O_1248,N_9202,N_9366);
or UO_1249 (O_1249,N_9030,N_9250);
or UO_1250 (O_1250,N_9943,N_9254);
or UO_1251 (O_1251,N_9045,N_9915);
and UO_1252 (O_1252,N_9347,N_9608);
and UO_1253 (O_1253,N_9762,N_9078);
nor UO_1254 (O_1254,N_9447,N_9067);
nand UO_1255 (O_1255,N_9533,N_9118);
or UO_1256 (O_1256,N_9215,N_9763);
nand UO_1257 (O_1257,N_9630,N_9785);
nor UO_1258 (O_1258,N_9057,N_9311);
nor UO_1259 (O_1259,N_9466,N_9099);
and UO_1260 (O_1260,N_9809,N_9411);
and UO_1261 (O_1261,N_9579,N_9853);
and UO_1262 (O_1262,N_9820,N_9497);
nor UO_1263 (O_1263,N_9967,N_9431);
nor UO_1264 (O_1264,N_9410,N_9002);
nor UO_1265 (O_1265,N_9890,N_9440);
or UO_1266 (O_1266,N_9709,N_9363);
nand UO_1267 (O_1267,N_9994,N_9178);
or UO_1268 (O_1268,N_9771,N_9004);
and UO_1269 (O_1269,N_9043,N_9029);
nor UO_1270 (O_1270,N_9815,N_9102);
and UO_1271 (O_1271,N_9315,N_9409);
nand UO_1272 (O_1272,N_9096,N_9097);
nor UO_1273 (O_1273,N_9642,N_9452);
nor UO_1274 (O_1274,N_9095,N_9131);
or UO_1275 (O_1275,N_9687,N_9361);
nor UO_1276 (O_1276,N_9812,N_9452);
nor UO_1277 (O_1277,N_9018,N_9389);
nor UO_1278 (O_1278,N_9645,N_9106);
nor UO_1279 (O_1279,N_9526,N_9274);
or UO_1280 (O_1280,N_9939,N_9562);
nand UO_1281 (O_1281,N_9244,N_9115);
nor UO_1282 (O_1282,N_9941,N_9371);
nor UO_1283 (O_1283,N_9450,N_9409);
nor UO_1284 (O_1284,N_9249,N_9649);
and UO_1285 (O_1285,N_9344,N_9006);
nand UO_1286 (O_1286,N_9326,N_9882);
or UO_1287 (O_1287,N_9557,N_9617);
or UO_1288 (O_1288,N_9094,N_9471);
nand UO_1289 (O_1289,N_9247,N_9648);
nor UO_1290 (O_1290,N_9357,N_9310);
nor UO_1291 (O_1291,N_9467,N_9402);
nand UO_1292 (O_1292,N_9427,N_9112);
xor UO_1293 (O_1293,N_9300,N_9697);
or UO_1294 (O_1294,N_9713,N_9022);
and UO_1295 (O_1295,N_9795,N_9859);
nand UO_1296 (O_1296,N_9958,N_9197);
and UO_1297 (O_1297,N_9725,N_9635);
and UO_1298 (O_1298,N_9047,N_9730);
or UO_1299 (O_1299,N_9610,N_9022);
nor UO_1300 (O_1300,N_9026,N_9614);
or UO_1301 (O_1301,N_9801,N_9750);
nand UO_1302 (O_1302,N_9459,N_9188);
nor UO_1303 (O_1303,N_9263,N_9661);
nor UO_1304 (O_1304,N_9771,N_9977);
nand UO_1305 (O_1305,N_9045,N_9324);
nand UO_1306 (O_1306,N_9668,N_9210);
and UO_1307 (O_1307,N_9489,N_9398);
nand UO_1308 (O_1308,N_9616,N_9722);
and UO_1309 (O_1309,N_9926,N_9979);
or UO_1310 (O_1310,N_9031,N_9007);
and UO_1311 (O_1311,N_9465,N_9700);
nand UO_1312 (O_1312,N_9772,N_9120);
or UO_1313 (O_1313,N_9919,N_9781);
and UO_1314 (O_1314,N_9946,N_9737);
and UO_1315 (O_1315,N_9543,N_9159);
and UO_1316 (O_1316,N_9290,N_9378);
or UO_1317 (O_1317,N_9557,N_9216);
and UO_1318 (O_1318,N_9092,N_9015);
or UO_1319 (O_1319,N_9495,N_9938);
and UO_1320 (O_1320,N_9384,N_9395);
or UO_1321 (O_1321,N_9340,N_9830);
or UO_1322 (O_1322,N_9042,N_9572);
and UO_1323 (O_1323,N_9713,N_9621);
xor UO_1324 (O_1324,N_9063,N_9220);
and UO_1325 (O_1325,N_9884,N_9969);
nand UO_1326 (O_1326,N_9880,N_9609);
nand UO_1327 (O_1327,N_9920,N_9098);
nor UO_1328 (O_1328,N_9767,N_9309);
and UO_1329 (O_1329,N_9846,N_9054);
nand UO_1330 (O_1330,N_9111,N_9796);
nand UO_1331 (O_1331,N_9985,N_9315);
nand UO_1332 (O_1332,N_9540,N_9729);
or UO_1333 (O_1333,N_9504,N_9671);
and UO_1334 (O_1334,N_9809,N_9163);
and UO_1335 (O_1335,N_9537,N_9668);
nand UO_1336 (O_1336,N_9273,N_9055);
nand UO_1337 (O_1337,N_9918,N_9023);
nand UO_1338 (O_1338,N_9506,N_9975);
nand UO_1339 (O_1339,N_9428,N_9314);
nand UO_1340 (O_1340,N_9899,N_9366);
and UO_1341 (O_1341,N_9918,N_9803);
and UO_1342 (O_1342,N_9654,N_9258);
and UO_1343 (O_1343,N_9387,N_9347);
or UO_1344 (O_1344,N_9043,N_9372);
or UO_1345 (O_1345,N_9075,N_9502);
and UO_1346 (O_1346,N_9084,N_9133);
nand UO_1347 (O_1347,N_9384,N_9409);
or UO_1348 (O_1348,N_9490,N_9514);
nand UO_1349 (O_1349,N_9718,N_9208);
nand UO_1350 (O_1350,N_9548,N_9097);
xnor UO_1351 (O_1351,N_9165,N_9056);
or UO_1352 (O_1352,N_9201,N_9421);
nand UO_1353 (O_1353,N_9263,N_9534);
and UO_1354 (O_1354,N_9655,N_9359);
or UO_1355 (O_1355,N_9804,N_9028);
and UO_1356 (O_1356,N_9332,N_9557);
and UO_1357 (O_1357,N_9251,N_9018);
nand UO_1358 (O_1358,N_9319,N_9380);
nand UO_1359 (O_1359,N_9141,N_9468);
and UO_1360 (O_1360,N_9498,N_9996);
xnor UO_1361 (O_1361,N_9634,N_9037);
nor UO_1362 (O_1362,N_9366,N_9413);
or UO_1363 (O_1363,N_9317,N_9032);
nor UO_1364 (O_1364,N_9920,N_9994);
or UO_1365 (O_1365,N_9558,N_9854);
and UO_1366 (O_1366,N_9878,N_9264);
and UO_1367 (O_1367,N_9018,N_9237);
or UO_1368 (O_1368,N_9269,N_9533);
and UO_1369 (O_1369,N_9604,N_9006);
and UO_1370 (O_1370,N_9067,N_9436);
or UO_1371 (O_1371,N_9974,N_9307);
and UO_1372 (O_1372,N_9329,N_9140);
or UO_1373 (O_1373,N_9861,N_9985);
nand UO_1374 (O_1374,N_9255,N_9262);
nor UO_1375 (O_1375,N_9793,N_9709);
xnor UO_1376 (O_1376,N_9791,N_9200);
and UO_1377 (O_1377,N_9756,N_9784);
or UO_1378 (O_1378,N_9384,N_9439);
or UO_1379 (O_1379,N_9996,N_9201);
xnor UO_1380 (O_1380,N_9033,N_9424);
nor UO_1381 (O_1381,N_9121,N_9600);
or UO_1382 (O_1382,N_9864,N_9629);
nand UO_1383 (O_1383,N_9407,N_9046);
or UO_1384 (O_1384,N_9037,N_9658);
xor UO_1385 (O_1385,N_9897,N_9009);
and UO_1386 (O_1386,N_9598,N_9262);
and UO_1387 (O_1387,N_9104,N_9672);
nor UO_1388 (O_1388,N_9435,N_9622);
or UO_1389 (O_1389,N_9560,N_9122);
nand UO_1390 (O_1390,N_9706,N_9881);
or UO_1391 (O_1391,N_9985,N_9537);
nor UO_1392 (O_1392,N_9913,N_9388);
nand UO_1393 (O_1393,N_9117,N_9906);
or UO_1394 (O_1394,N_9450,N_9439);
or UO_1395 (O_1395,N_9351,N_9949);
nand UO_1396 (O_1396,N_9212,N_9998);
nand UO_1397 (O_1397,N_9427,N_9938);
and UO_1398 (O_1398,N_9034,N_9446);
nor UO_1399 (O_1399,N_9806,N_9709);
nand UO_1400 (O_1400,N_9548,N_9377);
nand UO_1401 (O_1401,N_9356,N_9281);
and UO_1402 (O_1402,N_9958,N_9313);
and UO_1403 (O_1403,N_9928,N_9443);
or UO_1404 (O_1404,N_9849,N_9221);
and UO_1405 (O_1405,N_9916,N_9570);
and UO_1406 (O_1406,N_9719,N_9033);
nor UO_1407 (O_1407,N_9733,N_9476);
nand UO_1408 (O_1408,N_9271,N_9504);
nand UO_1409 (O_1409,N_9238,N_9397);
nor UO_1410 (O_1410,N_9584,N_9371);
nand UO_1411 (O_1411,N_9086,N_9775);
nand UO_1412 (O_1412,N_9637,N_9600);
and UO_1413 (O_1413,N_9750,N_9475);
and UO_1414 (O_1414,N_9072,N_9600);
or UO_1415 (O_1415,N_9998,N_9860);
or UO_1416 (O_1416,N_9502,N_9908);
nor UO_1417 (O_1417,N_9141,N_9873);
and UO_1418 (O_1418,N_9092,N_9177);
or UO_1419 (O_1419,N_9135,N_9786);
and UO_1420 (O_1420,N_9202,N_9197);
nor UO_1421 (O_1421,N_9766,N_9817);
nand UO_1422 (O_1422,N_9228,N_9639);
nand UO_1423 (O_1423,N_9132,N_9226);
nor UO_1424 (O_1424,N_9281,N_9463);
xor UO_1425 (O_1425,N_9082,N_9338);
and UO_1426 (O_1426,N_9687,N_9790);
nand UO_1427 (O_1427,N_9984,N_9469);
and UO_1428 (O_1428,N_9065,N_9333);
xnor UO_1429 (O_1429,N_9892,N_9250);
or UO_1430 (O_1430,N_9080,N_9614);
nand UO_1431 (O_1431,N_9064,N_9271);
nor UO_1432 (O_1432,N_9363,N_9055);
nor UO_1433 (O_1433,N_9097,N_9141);
or UO_1434 (O_1434,N_9162,N_9844);
and UO_1435 (O_1435,N_9908,N_9175);
or UO_1436 (O_1436,N_9483,N_9395);
or UO_1437 (O_1437,N_9751,N_9726);
or UO_1438 (O_1438,N_9275,N_9941);
or UO_1439 (O_1439,N_9797,N_9854);
nand UO_1440 (O_1440,N_9691,N_9524);
nor UO_1441 (O_1441,N_9478,N_9951);
and UO_1442 (O_1442,N_9810,N_9531);
nor UO_1443 (O_1443,N_9277,N_9230);
nor UO_1444 (O_1444,N_9870,N_9795);
nand UO_1445 (O_1445,N_9168,N_9475);
or UO_1446 (O_1446,N_9496,N_9680);
or UO_1447 (O_1447,N_9648,N_9282);
or UO_1448 (O_1448,N_9261,N_9733);
nand UO_1449 (O_1449,N_9034,N_9931);
or UO_1450 (O_1450,N_9933,N_9670);
nand UO_1451 (O_1451,N_9169,N_9666);
or UO_1452 (O_1452,N_9465,N_9309);
and UO_1453 (O_1453,N_9208,N_9318);
nand UO_1454 (O_1454,N_9896,N_9491);
and UO_1455 (O_1455,N_9348,N_9030);
and UO_1456 (O_1456,N_9999,N_9671);
or UO_1457 (O_1457,N_9131,N_9838);
nand UO_1458 (O_1458,N_9743,N_9800);
and UO_1459 (O_1459,N_9017,N_9288);
nor UO_1460 (O_1460,N_9240,N_9500);
nor UO_1461 (O_1461,N_9813,N_9783);
nand UO_1462 (O_1462,N_9976,N_9971);
nor UO_1463 (O_1463,N_9147,N_9607);
xnor UO_1464 (O_1464,N_9972,N_9475);
nand UO_1465 (O_1465,N_9232,N_9255);
nor UO_1466 (O_1466,N_9700,N_9503);
or UO_1467 (O_1467,N_9679,N_9441);
or UO_1468 (O_1468,N_9109,N_9580);
or UO_1469 (O_1469,N_9844,N_9680);
nand UO_1470 (O_1470,N_9125,N_9860);
and UO_1471 (O_1471,N_9570,N_9513);
nor UO_1472 (O_1472,N_9597,N_9223);
nand UO_1473 (O_1473,N_9888,N_9625);
nand UO_1474 (O_1474,N_9130,N_9823);
or UO_1475 (O_1475,N_9798,N_9766);
nor UO_1476 (O_1476,N_9996,N_9473);
and UO_1477 (O_1477,N_9172,N_9929);
nor UO_1478 (O_1478,N_9730,N_9376);
nor UO_1479 (O_1479,N_9035,N_9530);
nand UO_1480 (O_1480,N_9975,N_9375);
xor UO_1481 (O_1481,N_9153,N_9140);
or UO_1482 (O_1482,N_9510,N_9519);
nand UO_1483 (O_1483,N_9319,N_9589);
nor UO_1484 (O_1484,N_9994,N_9886);
or UO_1485 (O_1485,N_9372,N_9819);
or UO_1486 (O_1486,N_9488,N_9012);
and UO_1487 (O_1487,N_9425,N_9506);
or UO_1488 (O_1488,N_9517,N_9266);
or UO_1489 (O_1489,N_9196,N_9390);
nor UO_1490 (O_1490,N_9915,N_9134);
nand UO_1491 (O_1491,N_9359,N_9919);
and UO_1492 (O_1492,N_9460,N_9541);
or UO_1493 (O_1493,N_9710,N_9188);
nand UO_1494 (O_1494,N_9793,N_9336);
nor UO_1495 (O_1495,N_9030,N_9643);
nor UO_1496 (O_1496,N_9020,N_9583);
nand UO_1497 (O_1497,N_9519,N_9066);
nor UO_1498 (O_1498,N_9306,N_9330);
nor UO_1499 (O_1499,N_9140,N_9829);
endmodule