module basic_500_3000_500_30_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_307,In_359);
or U1 (N_1,In_50,In_324);
and U2 (N_2,In_62,In_314);
or U3 (N_3,In_187,In_145);
or U4 (N_4,In_199,In_432);
nand U5 (N_5,In_107,In_373);
xor U6 (N_6,In_451,In_56);
or U7 (N_7,In_477,In_177);
and U8 (N_8,In_156,In_424);
or U9 (N_9,In_97,In_89);
nor U10 (N_10,In_384,In_208);
xnor U11 (N_11,In_102,In_498);
nor U12 (N_12,In_281,In_457);
or U13 (N_13,In_261,In_288);
or U14 (N_14,In_455,In_146);
or U15 (N_15,In_106,In_226);
xnor U16 (N_16,In_240,In_2);
and U17 (N_17,In_257,In_118);
nand U18 (N_18,In_55,In_139);
xnor U19 (N_19,In_313,In_248);
nand U20 (N_20,In_27,In_178);
nor U21 (N_21,In_181,In_399);
nor U22 (N_22,In_166,In_251);
nor U23 (N_23,In_31,In_459);
or U24 (N_24,In_273,In_265);
or U25 (N_25,In_300,In_380);
xnor U26 (N_26,In_236,In_35);
and U27 (N_27,In_354,In_452);
nand U28 (N_28,In_174,In_425);
xor U29 (N_29,In_168,In_374);
nand U30 (N_30,In_47,In_271);
and U31 (N_31,In_329,In_194);
xnor U32 (N_32,In_103,In_396);
nand U33 (N_33,In_496,In_165);
xnor U34 (N_34,In_244,In_392);
nand U35 (N_35,In_88,In_376);
nand U36 (N_36,In_317,In_95);
and U37 (N_37,In_119,In_91);
xnor U38 (N_38,In_293,In_440);
nand U39 (N_39,In_339,In_475);
xnor U40 (N_40,In_90,In_442);
xnor U41 (N_41,In_254,In_70);
nor U42 (N_42,In_344,In_435);
nand U43 (N_43,In_110,In_80);
xnor U44 (N_44,In_382,In_332);
or U45 (N_45,In_113,In_25);
or U46 (N_46,In_169,In_355);
nor U47 (N_47,In_338,In_22);
and U48 (N_48,In_356,In_108);
nor U49 (N_49,In_426,In_397);
or U50 (N_50,In_465,In_391);
nor U51 (N_51,In_492,In_176);
nor U52 (N_52,In_137,In_231);
xor U53 (N_53,In_65,In_147);
or U54 (N_54,In_164,In_403);
nor U55 (N_55,In_441,In_390);
and U56 (N_56,In_245,In_429);
or U57 (N_57,In_476,In_252);
or U58 (N_58,In_310,In_109);
or U59 (N_59,In_283,In_234);
or U60 (N_60,In_469,In_458);
nor U61 (N_61,In_93,In_184);
xor U62 (N_62,In_454,In_152);
xor U63 (N_63,In_61,In_287);
nor U64 (N_64,In_79,In_453);
xnor U65 (N_65,In_331,In_82);
and U66 (N_66,In_418,In_279);
xor U67 (N_67,In_294,In_23);
xnor U68 (N_68,In_328,In_112);
nor U69 (N_69,In_73,In_34);
nor U70 (N_70,In_346,In_488);
nand U71 (N_71,In_48,In_189);
and U72 (N_72,In_437,In_198);
xor U73 (N_73,In_436,In_431);
nor U74 (N_74,In_158,In_408);
xor U75 (N_75,In_214,In_282);
and U76 (N_76,In_49,In_303);
xnor U77 (N_77,In_446,In_207);
and U78 (N_78,In_370,In_149);
nand U79 (N_79,In_443,In_215);
xnor U80 (N_80,In_341,In_201);
or U81 (N_81,In_378,In_77);
nand U82 (N_82,In_179,In_100);
nor U83 (N_83,In_369,In_220);
and U84 (N_84,In_362,In_241);
or U85 (N_85,In_84,In_322);
and U86 (N_86,In_232,In_98);
or U87 (N_87,In_182,In_306);
nor U88 (N_88,In_301,In_81);
xor U89 (N_89,In_143,In_447);
nor U90 (N_90,In_71,In_327);
nand U91 (N_91,In_1,In_272);
and U92 (N_92,In_197,In_295);
or U93 (N_93,In_337,In_478);
xor U94 (N_94,In_123,In_490);
nor U95 (N_95,In_404,In_167);
nor U96 (N_96,In_37,In_414);
nor U97 (N_97,In_0,In_218);
nand U98 (N_98,In_239,In_308);
nand U99 (N_99,In_290,In_489);
nand U100 (N_100,In_473,N_23);
xor U101 (N_101,In_188,N_1);
xor U102 (N_102,In_333,In_52);
xor U103 (N_103,N_9,In_63);
or U104 (N_104,In_230,In_227);
and U105 (N_105,In_450,In_135);
xor U106 (N_106,In_468,In_334);
xnor U107 (N_107,In_367,N_11);
nand U108 (N_108,In_266,In_379);
and U109 (N_109,In_321,N_81);
nor U110 (N_110,In_32,In_402);
nand U111 (N_111,N_18,In_40);
and U112 (N_112,N_6,In_438);
and U113 (N_113,In_330,In_368);
xor U114 (N_114,In_345,In_246);
or U115 (N_115,In_289,N_32);
xnor U116 (N_116,N_83,In_250);
nand U117 (N_117,In_161,In_15);
and U118 (N_118,In_284,In_213);
and U119 (N_119,In_260,In_92);
nand U120 (N_120,In_38,N_51);
or U121 (N_121,In_115,In_54);
and U122 (N_122,In_43,In_130);
xnor U123 (N_123,In_150,In_393);
nand U124 (N_124,In_493,In_361);
and U125 (N_125,N_56,N_28);
nand U126 (N_126,In_39,In_263);
nand U127 (N_127,In_316,N_24);
or U128 (N_128,In_280,N_59);
nor U129 (N_129,In_340,In_401);
xnor U130 (N_130,N_61,In_170);
or U131 (N_131,N_96,N_25);
xnor U132 (N_132,In_5,In_302);
xor U133 (N_133,N_63,In_444);
nand U134 (N_134,In_256,In_409);
and U135 (N_135,In_372,In_315);
or U136 (N_136,N_8,In_242);
nand U137 (N_137,In_190,In_153);
nor U138 (N_138,In_486,N_3);
xnor U139 (N_139,In_375,In_292);
nor U140 (N_140,In_462,In_223);
and U141 (N_141,In_349,N_19);
or U142 (N_142,In_212,In_456);
or U143 (N_143,In_229,In_318);
xor U144 (N_144,In_472,In_268);
or U145 (N_145,N_88,In_175);
nand U146 (N_146,In_484,In_383);
nand U147 (N_147,In_258,N_84);
xor U148 (N_148,N_50,In_445);
and U149 (N_149,In_66,In_204);
or U150 (N_150,In_124,In_78);
nand U151 (N_151,In_36,N_16);
xor U152 (N_152,In_466,In_304);
or U153 (N_153,In_16,In_99);
or U154 (N_154,In_427,In_497);
nand U155 (N_155,In_159,In_148);
nand U156 (N_156,N_20,N_2);
or U157 (N_157,N_94,In_395);
xnor U158 (N_158,N_82,N_33);
xnor U159 (N_159,In_157,In_224);
and U160 (N_160,N_67,N_38);
nor U161 (N_161,N_34,In_68);
or U162 (N_162,N_41,In_243);
xnor U163 (N_163,In_342,N_60);
nand U164 (N_164,In_144,In_28);
nor U165 (N_165,In_96,In_311);
nand U166 (N_166,N_86,In_494);
nand U167 (N_167,In_365,In_267);
nor U168 (N_168,In_186,In_298);
nor U169 (N_169,N_48,In_377);
or U170 (N_170,In_479,In_196);
and U171 (N_171,In_86,In_64);
nand U172 (N_172,In_275,In_128);
nand U173 (N_173,In_210,N_7);
nor U174 (N_174,In_195,In_485);
nor U175 (N_175,In_480,In_471);
or U176 (N_176,In_151,N_47);
xnor U177 (N_177,N_57,In_495);
xnor U178 (N_178,In_417,In_117);
nand U179 (N_179,In_12,In_274);
or U180 (N_180,In_323,In_398);
nor U181 (N_181,N_80,In_219);
and U182 (N_182,In_421,N_40);
or U183 (N_183,N_89,N_26);
or U184 (N_184,In_228,N_71);
nor U185 (N_185,In_30,In_413);
or U186 (N_186,N_99,In_101);
xor U187 (N_187,In_141,In_385);
nand U188 (N_188,In_448,In_138);
nor U189 (N_189,In_114,N_12);
nand U190 (N_190,In_60,In_222);
and U191 (N_191,In_21,In_312);
nor U192 (N_192,In_449,In_430);
xor U193 (N_193,In_7,N_66);
and U194 (N_194,In_129,In_203);
or U195 (N_195,N_70,N_39);
xor U196 (N_196,In_26,In_132);
xor U197 (N_197,In_405,In_121);
and U198 (N_198,In_45,N_17);
xnor U199 (N_199,In_255,In_76);
nand U200 (N_200,In_131,N_105);
nand U201 (N_201,In_59,In_155);
or U202 (N_202,In_343,N_168);
or U203 (N_203,N_58,N_134);
nand U204 (N_204,N_77,N_150);
nand U205 (N_205,In_238,N_175);
or U206 (N_206,N_187,In_416);
and U207 (N_207,In_154,In_217);
or U208 (N_208,N_198,In_42);
nor U209 (N_209,N_189,In_360);
nor U210 (N_210,In_353,In_185);
and U211 (N_211,In_8,In_269);
and U212 (N_212,In_352,In_400);
and U213 (N_213,In_24,N_75);
nand U214 (N_214,In_20,N_164);
nand U215 (N_215,In_72,N_0);
xnor U216 (N_216,In_183,N_186);
and U217 (N_217,N_120,In_193);
nor U218 (N_218,In_134,N_153);
and U219 (N_219,N_142,N_76);
nand U220 (N_220,In_297,N_95);
nor U221 (N_221,In_122,In_309);
nor U222 (N_222,In_57,In_180);
nor U223 (N_223,In_299,In_433);
or U224 (N_224,N_114,N_46);
or U225 (N_225,In_14,N_112);
nand U226 (N_226,N_167,In_51);
or U227 (N_227,In_83,In_461);
and U228 (N_228,In_348,N_193);
nor U229 (N_229,In_74,N_144);
nor U230 (N_230,In_120,In_225);
nand U231 (N_231,In_411,In_336);
nand U232 (N_232,N_136,N_45);
nand U233 (N_233,N_68,In_85);
nor U234 (N_234,N_10,N_30);
nand U235 (N_235,In_171,N_54);
nand U236 (N_236,N_5,N_107);
nor U237 (N_237,In_216,N_180);
and U238 (N_238,N_103,N_163);
or U239 (N_239,In_163,In_285);
nand U240 (N_240,In_10,N_73);
nor U241 (N_241,In_202,In_192);
xnor U242 (N_242,In_286,In_162);
xnor U243 (N_243,In_364,N_139);
nor U244 (N_244,N_104,N_129);
xor U245 (N_245,In_277,N_156);
and U246 (N_246,In_44,N_171);
xor U247 (N_247,N_159,In_491);
or U248 (N_248,N_151,In_464);
xnor U249 (N_249,In_319,In_233);
xor U250 (N_250,In_264,N_141);
nor U251 (N_251,In_278,In_420);
or U252 (N_252,N_170,In_116);
nor U253 (N_253,In_406,N_35);
or U254 (N_254,In_487,N_160);
nand U255 (N_255,N_62,In_335);
nand U256 (N_256,N_121,N_143);
or U257 (N_257,In_18,In_387);
xnor U258 (N_258,In_13,In_6);
nand U259 (N_259,N_145,N_190);
nor U260 (N_260,In_415,In_276);
nor U261 (N_261,In_67,In_235);
nand U262 (N_262,In_211,N_53);
nand U263 (N_263,N_192,N_102);
or U264 (N_264,N_55,N_147);
nor U265 (N_265,In_17,N_87);
or U266 (N_266,In_41,N_52);
nand U267 (N_267,In_419,N_98);
and U268 (N_268,N_65,In_291);
or U269 (N_269,N_146,In_75);
or U270 (N_270,N_124,In_388);
xnor U271 (N_271,In_136,In_237);
xnor U272 (N_272,N_122,In_160);
xor U273 (N_273,N_15,N_78);
nand U274 (N_274,In_463,N_131);
nor U275 (N_275,N_108,In_29);
and U276 (N_276,N_194,In_69);
nand U277 (N_277,In_46,N_79);
or U278 (N_278,N_93,N_161);
nor U279 (N_279,N_140,N_85);
nor U280 (N_280,In_140,N_174);
nand U281 (N_281,N_64,N_123);
and U282 (N_282,N_29,N_135);
nor U283 (N_283,N_22,N_4);
xnor U284 (N_284,In_407,In_259);
nor U285 (N_285,N_74,In_386);
nand U286 (N_286,N_176,N_92);
and U287 (N_287,In_53,N_155);
nor U288 (N_288,N_36,In_19);
or U289 (N_289,N_127,N_169);
nor U290 (N_290,N_181,In_423);
nor U291 (N_291,In_125,N_115);
and U292 (N_292,N_13,In_200);
nand U293 (N_293,In_262,N_109);
nor U294 (N_294,In_363,In_173);
nand U295 (N_295,In_470,In_127);
nor U296 (N_296,In_9,In_206);
xnor U297 (N_297,N_157,In_247);
or U298 (N_298,N_138,N_43);
nand U299 (N_299,N_111,In_94);
or U300 (N_300,N_196,N_148);
and U301 (N_301,N_154,N_228);
xor U302 (N_302,N_249,N_128);
xnor U303 (N_303,In_460,N_297);
nor U304 (N_304,N_231,N_276);
and U305 (N_305,In_358,N_256);
xor U306 (N_306,N_183,N_27);
xnor U307 (N_307,N_226,In_371);
or U308 (N_308,In_347,N_217);
and U309 (N_309,N_91,N_191);
or U310 (N_310,N_130,In_351);
nand U311 (N_311,N_218,N_233);
or U312 (N_312,N_90,In_357);
nor U313 (N_313,N_230,N_125);
or U314 (N_314,N_287,N_229);
nand U315 (N_315,N_210,In_270);
xor U316 (N_316,In_474,In_104);
nand U317 (N_317,N_296,In_249);
xor U318 (N_318,In_320,N_201);
or U319 (N_319,In_428,N_290);
and U320 (N_320,N_243,N_227);
nand U321 (N_321,N_44,N_298);
nor U322 (N_322,N_208,N_279);
or U323 (N_323,N_283,In_394);
nand U324 (N_324,N_236,N_247);
xnor U325 (N_325,N_110,N_21);
xor U326 (N_326,N_289,N_267);
and U327 (N_327,N_252,In_296);
nand U328 (N_328,N_200,In_381);
nor U329 (N_329,N_237,N_266);
and U330 (N_330,N_224,In_350);
or U331 (N_331,N_240,N_254);
and U332 (N_332,In_412,In_172);
xnor U333 (N_333,In_11,N_37);
and U334 (N_334,N_261,N_158);
or U335 (N_335,N_101,N_250);
and U336 (N_336,N_100,N_179);
nor U337 (N_337,N_215,N_216);
xor U338 (N_338,In_3,N_262);
or U339 (N_339,N_207,In_434);
and U340 (N_340,N_49,N_264);
nor U341 (N_341,In_422,N_205);
nor U342 (N_342,In_482,N_282);
nor U343 (N_343,N_195,In_467);
nand U344 (N_344,N_212,N_185);
xnor U345 (N_345,In_483,In_191);
xor U346 (N_346,In_410,In_221);
xnor U347 (N_347,N_223,N_72);
and U348 (N_348,N_241,N_31);
and U349 (N_349,In_253,N_271);
and U350 (N_350,N_268,In_439);
and U351 (N_351,N_270,N_278);
nand U352 (N_352,N_178,N_221);
and U353 (N_353,N_204,N_106);
nor U354 (N_354,In_305,N_199);
nor U355 (N_355,N_291,N_172);
nor U356 (N_356,N_166,N_272);
or U357 (N_357,N_238,N_42);
or U358 (N_358,N_248,N_292);
nand U359 (N_359,N_234,N_284);
nand U360 (N_360,N_14,N_286);
xor U361 (N_361,N_225,In_58);
nand U362 (N_362,N_119,N_177);
xnor U363 (N_363,N_184,N_258);
and U364 (N_364,In_205,In_209);
xor U365 (N_365,N_232,N_244);
and U366 (N_366,N_213,N_235);
nand U367 (N_367,N_188,N_295);
and U368 (N_368,N_118,N_220);
xnor U369 (N_369,N_152,N_257);
and U370 (N_370,In_87,N_280);
and U371 (N_371,N_285,N_260);
xor U372 (N_372,N_165,N_133);
xor U373 (N_373,N_273,N_242);
nor U374 (N_374,N_294,N_222);
xor U375 (N_375,N_203,In_326);
nor U376 (N_376,N_126,N_251);
nand U377 (N_377,N_209,N_214);
xnor U378 (N_378,N_275,In_481);
nand U379 (N_379,In_126,In_33);
xnor U380 (N_380,N_206,In_133);
nand U381 (N_381,N_299,N_137);
nand U382 (N_382,N_69,In_499);
or U383 (N_383,In_4,N_246);
and U384 (N_384,N_277,In_142);
and U385 (N_385,N_182,N_149);
xor U386 (N_386,N_259,N_255);
nor U387 (N_387,N_263,In_325);
nand U388 (N_388,N_281,N_265);
and U389 (N_389,N_211,N_269);
nor U390 (N_390,N_245,N_239);
nand U391 (N_391,In_366,In_111);
xor U392 (N_392,N_293,In_389);
nor U393 (N_393,N_173,In_105);
nor U394 (N_394,N_219,N_288);
or U395 (N_395,N_132,N_117);
xnor U396 (N_396,N_253,N_97);
or U397 (N_397,N_202,N_162);
or U398 (N_398,N_197,N_116);
xnor U399 (N_399,N_113,N_274);
or U400 (N_400,N_384,N_306);
nor U401 (N_401,N_334,N_330);
nor U402 (N_402,N_344,N_343);
and U403 (N_403,N_388,N_386);
or U404 (N_404,N_316,N_369);
xnor U405 (N_405,N_320,N_350);
nand U406 (N_406,N_321,N_362);
xnor U407 (N_407,N_300,N_385);
nand U408 (N_408,N_302,N_315);
nor U409 (N_409,N_374,N_383);
nor U410 (N_410,N_340,N_305);
or U411 (N_411,N_389,N_336);
and U412 (N_412,N_394,N_317);
and U413 (N_413,N_393,N_318);
xor U414 (N_414,N_373,N_301);
nor U415 (N_415,N_328,N_363);
or U416 (N_416,N_391,N_333);
nor U417 (N_417,N_365,N_364);
nand U418 (N_418,N_370,N_390);
xor U419 (N_419,N_339,N_352);
nand U420 (N_420,N_322,N_338);
nor U421 (N_421,N_307,N_380);
nand U422 (N_422,N_329,N_375);
nor U423 (N_423,N_371,N_304);
and U424 (N_424,N_327,N_331);
and U425 (N_425,N_381,N_367);
xnor U426 (N_426,N_382,N_353);
or U427 (N_427,N_358,N_324);
and U428 (N_428,N_347,N_356);
or U429 (N_429,N_359,N_313);
or U430 (N_430,N_355,N_372);
xor U431 (N_431,N_314,N_308);
or U432 (N_432,N_341,N_346);
nor U433 (N_433,N_379,N_395);
nor U434 (N_434,N_377,N_351);
or U435 (N_435,N_323,N_319);
and U436 (N_436,N_349,N_312);
and U437 (N_437,N_396,N_392);
nor U438 (N_438,N_397,N_378);
nand U439 (N_439,N_310,N_335);
nor U440 (N_440,N_325,N_360);
xor U441 (N_441,N_398,N_303);
or U442 (N_442,N_399,N_332);
xnor U443 (N_443,N_368,N_311);
nand U444 (N_444,N_354,N_387);
and U445 (N_445,N_366,N_342);
nor U446 (N_446,N_376,N_348);
nor U447 (N_447,N_326,N_357);
and U448 (N_448,N_309,N_345);
or U449 (N_449,N_337,N_361);
and U450 (N_450,N_398,N_363);
and U451 (N_451,N_328,N_331);
xnor U452 (N_452,N_388,N_336);
xor U453 (N_453,N_383,N_303);
or U454 (N_454,N_397,N_360);
xnor U455 (N_455,N_351,N_392);
or U456 (N_456,N_387,N_353);
and U457 (N_457,N_395,N_317);
nor U458 (N_458,N_346,N_316);
xor U459 (N_459,N_306,N_354);
or U460 (N_460,N_363,N_305);
and U461 (N_461,N_361,N_388);
or U462 (N_462,N_305,N_362);
nor U463 (N_463,N_351,N_321);
and U464 (N_464,N_344,N_368);
or U465 (N_465,N_312,N_351);
nand U466 (N_466,N_393,N_330);
xor U467 (N_467,N_375,N_387);
nand U468 (N_468,N_387,N_302);
and U469 (N_469,N_333,N_375);
and U470 (N_470,N_356,N_377);
xnor U471 (N_471,N_341,N_310);
or U472 (N_472,N_386,N_362);
xor U473 (N_473,N_303,N_333);
nand U474 (N_474,N_395,N_311);
xor U475 (N_475,N_379,N_383);
nand U476 (N_476,N_330,N_327);
and U477 (N_477,N_395,N_390);
or U478 (N_478,N_321,N_355);
xnor U479 (N_479,N_350,N_367);
or U480 (N_480,N_308,N_341);
nand U481 (N_481,N_344,N_358);
nor U482 (N_482,N_363,N_324);
nor U483 (N_483,N_336,N_366);
and U484 (N_484,N_313,N_378);
or U485 (N_485,N_397,N_358);
and U486 (N_486,N_345,N_383);
nand U487 (N_487,N_373,N_306);
nor U488 (N_488,N_306,N_377);
or U489 (N_489,N_324,N_302);
xnor U490 (N_490,N_338,N_325);
or U491 (N_491,N_311,N_393);
or U492 (N_492,N_390,N_376);
and U493 (N_493,N_356,N_333);
nand U494 (N_494,N_379,N_385);
nor U495 (N_495,N_321,N_343);
xor U496 (N_496,N_399,N_306);
nor U497 (N_497,N_346,N_375);
nand U498 (N_498,N_324,N_366);
and U499 (N_499,N_379,N_328);
xnor U500 (N_500,N_402,N_460);
and U501 (N_501,N_473,N_405);
xnor U502 (N_502,N_406,N_463);
nand U503 (N_503,N_490,N_469);
or U504 (N_504,N_457,N_413);
or U505 (N_505,N_474,N_441);
and U506 (N_506,N_414,N_481);
nand U507 (N_507,N_432,N_475);
or U508 (N_508,N_487,N_415);
or U509 (N_509,N_466,N_494);
xor U510 (N_510,N_429,N_461);
or U511 (N_511,N_440,N_489);
xor U512 (N_512,N_496,N_418);
and U513 (N_513,N_446,N_499);
or U514 (N_514,N_433,N_424);
xor U515 (N_515,N_409,N_465);
xor U516 (N_516,N_456,N_448);
xor U517 (N_517,N_412,N_479);
or U518 (N_518,N_485,N_428);
and U519 (N_519,N_491,N_482);
xnor U520 (N_520,N_449,N_403);
and U521 (N_521,N_458,N_472);
nor U522 (N_522,N_421,N_427);
and U523 (N_523,N_453,N_455);
nor U524 (N_524,N_425,N_417);
nand U525 (N_525,N_451,N_419);
xor U526 (N_526,N_437,N_401);
nand U527 (N_527,N_436,N_400);
or U528 (N_528,N_430,N_493);
nor U529 (N_529,N_464,N_488);
and U530 (N_530,N_444,N_404);
nor U531 (N_531,N_439,N_434);
nand U532 (N_532,N_470,N_438);
nand U533 (N_533,N_483,N_486);
nor U534 (N_534,N_423,N_416);
or U535 (N_535,N_478,N_471);
nand U536 (N_536,N_452,N_420);
nand U537 (N_537,N_498,N_495);
xor U538 (N_538,N_480,N_484);
nand U539 (N_539,N_426,N_450);
or U540 (N_540,N_468,N_410);
xor U541 (N_541,N_422,N_431);
xor U542 (N_542,N_435,N_408);
and U543 (N_543,N_492,N_445);
nand U544 (N_544,N_477,N_443);
xor U545 (N_545,N_454,N_476);
nor U546 (N_546,N_407,N_447);
nand U547 (N_547,N_497,N_467);
nor U548 (N_548,N_411,N_462);
xnor U549 (N_549,N_442,N_459);
xnor U550 (N_550,N_413,N_414);
or U551 (N_551,N_484,N_498);
and U552 (N_552,N_499,N_419);
and U553 (N_553,N_481,N_498);
and U554 (N_554,N_422,N_494);
nand U555 (N_555,N_479,N_488);
xnor U556 (N_556,N_405,N_419);
or U557 (N_557,N_428,N_421);
nor U558 (N_558,N_498,N_406);
nand U559 (N_559,N_486,N_423);
xor U560 (N_560,N_458,N_424);
nand U561 (N_561,N_483,N_415);
nand U562 (N_562,N_459,N_402);
nor U563 (N_563,N_422,N_419);
or U564 (N_564,N_490,N_472);
xnor U565 (N_565,N_488,N_497);
xnor U566 (N_566,N_424,N_417);
xnor U567 (N_567,N_424,N_476);
xnor U568 (N_568,N_479,N_426);
or U569 (N_569,N_425,N_482);
or U570 (N_570,N_458,N_457);
nand U571 (N_571,N_441,N_463);
xor U572 (N_572,N_449,N_408);
or U573 (N_573,N_400,N_492);
nor U574 (N_574,N_446,N_413);
nand U575 (N_575,N_439,N_436);
and U576 (N_576,N_471,N_433);
nand U577 (N_577,N_409,N_472);
and U578 (N_578,N_489,N_442);
nand U579 (N_579,N_454,N_468);
and U580 (N_580,N_491,N_480);
nand U581 (N_581,N_402,N_416);
or U582 (N_582,N_460,N_414);
nand U583 (N_583,N_461,N_424);
xnor U584 (N_584,N_413,N_439);
and U585 (N_585,N_467,N_432);
nand U586 (N_586,N_440,N_499);
nor U587 (N_587,N_404,N_428);
nor U588 (N_588,N_415,N_457);
and U589 (N_589,N_466,N_449);
nand U590 (N_590,N_417,N_444);
and U591 (N_591,N_446,N_427);
or U592 (N_592,N_483,N_402);
or U593 (N_593,N_438,N_487);
nand U594 (N_594,N_491,N_497);
nor U595 (N_595,N_442,N_491);
or U596 (N_596,N_498,N_493);
xnor U597 (N_597,N_452,N_478);
or U598 (N_598,N_459,N_486);
and U599 (N_599,N_454,N_447);
and U600 (N_600,N_583,N_539);
nand U601 (N_601,N_507,N_518);
nand U602 (N_602,N_515,N_533);
nand U603 (N_603,N_520,N_597);
and U604 (N_604,N_558,N_564);
nor U605 (N_605,N_501,N_567);
nand U606 (N_606,N_530,N_570);
nand U607 (N_607,N_512,N_553);
xnor U608 (N_608,N_529,N_527);
and U609 (N_609,N_513,N_588);
and U610 (N_610,N_587,N_582);
xnor U611 (N_611,N_516,N_580);
nor U612 (N_612,N_522,N_584);
xnor U613 (N_613,N_525,N_545);
xor U614 (N_614,N_538,N_537);
or U615 (N_615,N_581,N_571);
xnor U616 (N_616,N_562,N_504);
nor U617 (N_617,N_535,N_521);
xor U618 (N_618,N_547,N_566);
nand U619 (N_619,N_551,N_573);
nor U620 (N_620,N_544,N_598);
and U621 (N_621,N_565,N_578);
xnor U622 (N_622,N_503,N_593);
xor U623 (N_623,N_579,N_526);
nand U624 (N_624,N_549,N_532);
nor U625 (N_625,N_595,N_508);
and U626 (N_626,N_586,N_591);
or U627 (N_627,N_523,N_531);
nor U628 (N_628,N_576,N_528);
nor U629 (N_629,N_563,N_509);
xnor U630 (N_630,N_514,N_534);
nor U631 (N_631,N_575,N_524);
nor U632 (N_632,N_517,N_519);
xor U633 (N_633,N_568,N_552);
xor U634 (N_634,N_502,N_594);
nand U635 (N_635,N_557,N_590);
and U636 (N_636,N_536,N_511);
nor U637 (N_637,N_550,N_596);
or U638 (N_638,N_546,N_574);
nor U639 (N_639,N_561,N_555);
nand U640 (N_640,N_592,N_599);
xor U641 (N_641,N_548,N_554);
and U642 (N_642,N_559,N_560);
and U643 (N_643,N_543,N_572);
xor U644 (N_644,N_500,N_556);
and U645 (N_645,N_506,N_540);
nand U646 (N_646,N_569,N_589);
nor U647 (N_647,N_510,N_585);
xor U648 (N_648,N_541,N_542);
or U649 (N_649,N_505,N_577);
nor U650 (N_650,N_509,N_546);
xnor U651 (N_651,N_558,N_524);
xnor U652 (N_652,N_551,N_542);
nor U653 (N_653,N_504,N_531);
xor U654 (N_654,N_500,N_536);
nor U655 (N_655,N_565,N_545);
nor U656 (N_656,N_586,N_505);
or U657 (N_657,N_575,N_512);
or U658 (N_658,N_555,N_577);
or U659 (N_659,N_588,N_566);
or U660 (N_660,N_530,N_520);
nor U661 (N_661,N_576,N_547);
nor U662 (N_662,N_519,N_512);
nor U663 (N_663,N_574,N_534);
or U664 (N_664,N_588,N_505);
xnor U665 (N_665,N_526,N_549);
or U666 (N_666,N_507,N_552);
nand U667 (N_667,N_518,N_558);
xnor U668 (N_668,N_574,N_515);
or U669 (N_669,N_592,N_581);
nand U670 (N_670,N_589,N_543);
and U671 (N_671,N_582,N_596);
and U672 (N_672,N_560,N_557);
or U673 (N_673,N_541,N_579);
and U674 (N_674,N_582,N_565);
nand U675 (N_675,N_503,N_573);
and U676 (N_676,N_581,N_552);
nor U677 (N_677,N_584,N_565);
xnor U678 (N_678,N_525,N_574);
xor U679 (N_679,N_577,N_573);
nor U680 (N_680,N_513,N_547);
or U681 (N_681,N_525,N_513);
xor U682 (N_682,N_594,N_579);
xnor U683 (N_683,N_547,N_594);
nand U684 (N_684,N_511,N_525);
xor U685 (N_685,N_505,N_511);
and U686 (N_686,N_594,N_556);
xor U687 (N_687,N_562,N_501);
nand U688 (N_688,N_574,N_591);
nor U689 (N_689,N_558,N_554);
and U690 (N_690,N_555,N_512);
and U691 (N_691,N_546,N_503);
nor U692 (N_692,N_567,N_583);
or U693 (N_693,N_585,N_582);
or U694 (N_694,N_512,N_586);
xor U695 (N_695,N_529,N_582);
and U696 (N_696,N_554,N_580);
nor U697 (N_697,N_505,N_551);
or U698 (N_698,N_528,N_541);
and U699 (N_699,N_565,N_541);
or U700 (N_700,N_646,N_629);
and U701 (N_701,N_619,N_624);
nand U702 (N_702,N_618,N_610);
and U703 (N_703,N_684,N_695);
nor U704 (N_704,N_689,N_601);
or U705 (N_705,N_690,N_686);
or U706 (N_706,N_635,N_678);
nand U707 (N_707,N_651,N_634);
xnor U708 (N_708,N_687,N_631);
nand U709 (N_709,N_667,N_632);
and U710 (N_710,N_677,N_665);
and U711 (N_711,N_611,N_602);
or U712 (N_712,N_633,N_604);
and U713 (N_713,N_616,N_676);
nand U714 (N_714,N_636,N_642);
xor U715 (N_715,N_692,N_620);
nand U716 (N_716,N_666,N_614);
and U717 (N_717,N_679,N_648);
and U718 (N_718,N_658,N_696);
nor U719 (N_719,N_672,N_623);
xor U720 (N_720,N_673,N_699);
nor U721 (N_721,N_664,N_693);
nand U722 (N_722,N_650,N_606);
nor U723 (N_723,N_652,N_697);
and U724 (N_724,N_649,N_671);
or U725 (N_725,N_637,N_644);
and U726 (N_726,N_622,N_613);
nor U727 (N_727,N_661,N_612);
nand U728 (N_728,N_656,N_608);
and U729 (N_729,N_605,N_660);
or U730 (N_730,N_691,N_640);
nand U731 (N_731,N_615,N_680);
and U732 (N_732,N_674,N_688);
or U733 (N_733,N_645,N_681);
and U734 (N_734,N_625,N_630);
nand U735 (N_735,N_653,N_685);
nand U736 (N_736,N_603,N_647);
nand U737 (N_737,N_617,N_654);
xor U738 (N_738,N_668,N_682);
xor U739 (N_739,N_628,N_627);
nand U740 (N_740,N_639,N_621);
or U741 (N_741,N_609,N_626);
nand U742 (N_742,N_669,N_600);
or U743 (N_743,N_607,N_698);
and U744 (N_744,N_659,N_675);
nand U745 (N_745,N_670,N_657);
and U746 (N_746,N_655,N_641);
nor U747 (N_747,N_694,N_638);
xor U748 (N_748,N_662,N_643);
nor U749 (N_749,N_663,N_683);
xor U750 (N_750,N_653,N_641);
and U751 (N_751,N_657,N_644);
and U752 (N_752,N_633,N_670);
or U753 (N_753,N_668,N_612);
and U754 (N_754,N_687,N_612);
nor U755 (N_755,N_660,N_636);
and U756 (N_756,N_644,N_614);
nor U757 (N_757,N_632,N_633);
and U758 (N_758,N_682,N_621);
xnor U759 (N_759,N_639,N_655);
xnor U760 (N_760,N_673,N_619);
nor U761 (N_761,N_637,N_694);
and U762 (N_762,N_613,N_603);
nor U763 (N_763,N_638,N_606);
and U764 (N_764,N_619,N_669);
or U765 (N_765,N_601,N_648);
xor U766 (N_766,N_632,N_610);
xor U767 (N_767,N_655,N_665);
nand U768 (N_768,N_604,N_626);
and U769 (N_769,N_679,N_632);
nor U770 (N_770,N_603,N_691);
xor U771 (N_771,N_619,N_683);
nand U772 (N_772,N_624,N_697);
nor U773 (N_773,N_691,N_696);
nand U774 (N_774,N_619,N_696);
nand U775 (N_775,N_601,N_630);
or U776 (N_776,N_600,N_603);
and U777 (N_777,N_683,N_637);
nand U778 (N_778,N_631,N_695);
or U779 (N_779,N_655,N_635);
xnor U780 (N_780,N_646,N_663);
or U781 (N_781,N_696,N_655);
xnor U782 (N_782,N_697,N_681);
or U783 (N_783,N_639,N_686);
or U784 (N_784,N_632,N_639);
nand U785 (N_785,N_661,N_688);
nand U786 (N_786,N_629,N_674);
nor U787 (N_787,N_667,N_661);
xnor U788 (N_788,N_634,N_645);
nand U789 (N_789,N_610,N_625);
and U790 (N_790,N_649,N_626);
xnor U791 (N_791,N_666,N_619);
and U792 (N_792,N_602,N_639);
nand U793 (N_793,N_694,N_607);
xnor U794 (N_794,N_651,N_652);
and U795 (N_795,N_658,N_670);
or U796 (N_796,N_631,N_640);
nor U797 (N_797,N_686,N_695);
and U798 (N_798,N_665,N_633);
xnor U799 (N_799,N_609,N_641);
and U800 (N_800,N_792,N_709);
and U801 (N_801,N_791,N_705);
nand U802 (N_802,N_793,N_708);
xor U803 (N_803,N_706,N_751);
xnor U804 (N_804,N_720,N_760);
and U805 (N_805,N_780,N_772);
and U806 (N_806,N_788,N_797);
or U807 (N_807,N_714,N_785);
nor U808 (N_808,N_761,N_722);
or U809 (N_809,N_731,N_732);
or U810 (N_810,N_752,N_764);
or U811 (N_811,N_784,N_717);
nor U812 (N_812,N_723,N_715);
nor U813 (N_813,N_739,N_744);
xnor U814 (N_814,N_724,N_700);
nor U815 (N_815,N_740,N_721);
and U816 (N_816,N_726,N_738);
xnor U817 (N_817,N_755,N_707);
or U818 (N_818,N_786,N_796);
and U819 (N_819,N_753,N_771);
or U820 (N_820,N_735,N_776);
or U821 (N_821,N_711,N_748);
nand U822 (N_822,N_778,N_773);
or U823 (N_823,N_750,N_728);
xor U824 (N_824,N_762,N_733);
xnor U825 (N_825,N_747,N_736);
and U826 (N_826,N_765,N_741);
and U827 (N_827,N_756,N_787);
and U828 (N_828,N_768,N_712);
nor U829 (N_829,N_781,N_704);
xnor U830 (N_830,N_775,N_798);
xor U831 (N_831,N_716,N_737);
or U832 (N_832,N_719,N_782);
nand U833 (N_833,N_769,N_734);
nor U834 (N_834,N_727,N_794);
nor U835 (N_835,N_749,N_757);
or U836 (N_836,N_758,N_779);
or U837 (N_837,N_743,N_725);
or U838 (N_838,N_710,N_701);
or U839 (N_839,N_763,N_789);
xor U840 (N_840,N_783,N_770);
or U841 (N_841,N_729,N_799);
nor U842 (N_842,N_742,N_767);
xnor U843 (N_843,N_754,N_766);
nor U844 (N_844,N_777,N_702);
and U845 (N_845,N_718,N_730);
or U846 (N_846,N_713,N_703);
nor U847 (N_847,N_774,N_759);
and U848 (N_848,N_790,N_795);
nor U849 (N_849,N_745,N_746);
xnor U850 (N_850,N_772,N_721);
nor U851 (N_851,N_785,N_752);
nor U852 (N_852,N_784,N_773);
or U853 (N_853,N_782,N_740);
or U854 (N_854,N_758,N_705);
nor U855 (N_855,N_712,N_749);
xor U856 (N_856,N_773,N_763);
and U857 (N_857,N_775,N_760);
and U858 (N_858,N_766,N_749);
nor U859 (N_859,N_795,N_777);
nor U860 (N_860,N_711,N_790);
nor U861 (N_861,N_703,N_760);
nand U862 (N_862,N_788,N_742);
and U863 (N_863,N_751,N_705);
nor U864 (N_864,N_725,N_716);
and U865 (N_865,N_703,N_766);
nand U866 (N_866,N_715,N_789);
and U867 (N_867,N_774,N_788);
nor U868 (N_868,N_741,N_747);
nor U869 (N_869,N_756,N_776);
and U870 (N_870,N_715,N_708);
and U871 (N_871,N_779,N_725);
nor U872 (N_872,N_714,N_744);
and U873 (N_873,N_796,N_748);
xor U874 (N_874,N_743,N_798);
xor U875 (N_875,N_756,N_793);
or U876 (N_876,N_762,N_756);
nand U877 (N_877,N_737,N_730);
and U878 (N_878,N_785,N_737);
nand U879 (N_879,N_783,N_718);
or U880 (N_880,N_747,N_703);
or U881 (N_881,N_749,N_741);
and U882 (N_882,N_723,N_781);
and U883 (N_883,N_760,N_704);
or U884 (N_884,N_740,N_778);
and U885 (N_885,N_747,N_758);
and U886 (N_886,N_771,N_744);
nor U887 (N_887,N_769,N_766);
nand U888 (N_888,N_749,N_739);
nor U889 (N_889,N_707,N_794);
and U890 (N_890,N_774,N_701);
or U891 (N_891,N_707,N_746);
xor U892 (N_892,N_740,N_748);
and U893 (N_893,N_712,N_705);
or U894 (N_894,N_746,N_791);
nand U895 (N_895,N_745,N_748);
or U896 (N_896,N_759,N_709);
xnor U897 (N_897,N_786,N_722);
nand U898 (N_898,N_767,N_798);
and U899 (N_899,N_714,N_745);
and U900 (N_900,N_888,N_809);
nor U901 (N_901,N_870,N_863);
nand U902 (N_902,N_866,N_882);
nand U903 (N_903,N_874,N_875);
or U904 (N_904,N_878,N_831);
nor U905 (N_905,N_816,N_849);
or U906 (N_906,N_810,N_872);
and U907 (N_907,N_841,N_879);
nand U908 (N_908,N_853,N_820);
xnor U909 (N_909,N_830,N_898);
and U910 (N_910,N_836,N_806);
nand U911 (N_911,N_821,N_807);
nor U912 (N_912,N_834,N_881);
or U913 (N_913,N_860,N_823);
nand U914 (N_914,N_889,N_801);
xnor U915 (N_915,N_838,N_873);
or U916 (N_916,N_802,N_822);
nor U917 (N_917,N_800,N_887);
or U918 (N_918,N_843,N_867);
xnor U919 (N_919,N_859,N_855);
nand U920 (N_920,N_829,N_892);
and U921 (N_921,N_824,N_869);
or U922 (N_922,N_813,N_847);
nor U923 (N_923,N_856,N_818);
xnor U924 (N_924,N_840,N_845);
and U925 (N_925,N_884,N_844);
or U926 (N_926,N_891,N_803);
nor U927 (N_927,N_832,N_893);
or U928 (N_928,N_857,N_871);
and U929 (N_929,N_811,N_826);
nand U930 (N_930,N_833,N_850);
or U931 (N_931,N_864,N_899);
nand U932 (N_932,N_885,N_897);
nand U933 (N_933,N_854,N_880);
or U934 (N_934,N_890,N_846);
and U935 (N_935,N_865,N_848);
and U936 (N_936,N_896,N_815);
and U937 (N_937,N_851,N_876);
nand U938 (N_938,N_812,N_886);
and U939 (N_939,N_808,N_842);
nor U940 (N_940,N_805,N_862);
or U941 (N_941,N_895,N_828);
nor U942 (N_942,N_814,N_837);
or U943 (N_943,N_883,N_819);
xor U944 (N_944,N_861,N_858);
nor U945 (N_945,N_825,N_835);
nor U946 (N_946,N_852,N_877);
or U947 (N_947,N_839,N_894);
xor U948 (N_948,N_804,N_817);
nand U949 (N_949,N_827,N_868);
or U950 (N_950,N_819,N_878);
nor U951 (N_951,N_826,N_822);
or U952 (N_952,N_891,N_892);
and U953 (N_953,N_858,N_840);
xnor U954 (N_954,N_862,N_882);
nor U955 (N_955,N_864,N_810);
or U956 (N_956,N_866,N_877);
or U957 (N_957,N_813,N_832);
xor U958 (N_958,N_873,N_880);
nor U959 (N_959,N_818,N_866);
xnor U960 (N_960,N_857,N_838);
xnor U961 (N_961,N_842,N_843);
or U962 (N_962,N_888,N_835);
nor U963 (N_963,N_853,N_826);
or U964 (N_964,N_819,N_816);
nand U965 (N_965,N_845,N_817);
xor U966 (N_966,N_853,N_862);
nor U967 (N_967,N_887,N_811);
and U968 (N_968,N_879,N_882);
nand U969 (N_969,N_872,N_809);
and U970 (N_970,N_882,N_823);
xnor U971 (N_971,N_833,N_818);
xnor U972 (N_972,N_892,N_830);
nand U973 (N_973,N_861,N_897);
nor U974 (N_974,N_888,N_832);
and U975 (N_975,N_838,N_821);
and U976 (N_976,N_884,N_855);
and U977 (N_977,N_808,N_838);
xor U978 (N_978,N_800,N_898);
and U979 (N_979,N_861,N_878);
nand U980 (N_980,N_875,N_899);
nand U981 (N_981,N_822,N_891);
and U982 (N_982,N_861,N_837);
nand U983 (N_983,N_842,N_846);
and U984 (N_984,N_891,N_874);
xor U985 (N_985,N_809,N_880);
or U986 (N_986,N_861,N_894);
nor U987 (N_987,N_856,N_859);
or U988 (N_988,N_802,N_827);
xor U989 (N_989,N_815,N_850);
and U990 (N_990,N_818,N_834);
or U991 (N_991,N_842,N_864);
xor U992 (N_992,N_832,N_815);
xor U993 (N_993,N_819,N_830);
nor U994 (N_994,N_818,N_889);
nor U995 (N_995,N_889,N_873);
or U996 (N_996,N_898,N_835);
nand U997 (N_997,N_875,N_844);
and U998 (N_998,N_832,N_807);
xnor U999 (N_999,N_858,N_849);
or U1000 (N_1000,N_952,N_972);
xnor U1001 (N_1001,N_970,N_955);
nor U1002 (N_1002,N_935,N_966);
xor U1003 (N_1003,N_987,N_901);
and U1004 (N_1004,N_976,N_912);
and U1005 (N_1005,N_974,N_928);
or U1006 (N_1006,N_961,N_965);
or U1007 (N_1007,N_998,N_945);
xnor U1008 (N_1008,N_948,N_931);
or U1009 (N_1009,N_913,N_943);
nand U1010 (N_1010,N_908,N_944);
or U1011 (N_1011,N_906,N_997);
nand U1012 (N_1012,N_907,N_969);
nor U1013 (N_1013,N_940,N_927);
nand U1014 (N_1014,N_990,N_973);
or U1015 (N_1015,N_900,N_959);
xnor U1016 (N_1016,N_993,N_904);
nand U1017 (N_1017,N_934,N_916);
or U1018 (N_1018,N_930,N_938);
or U1019 (N_1019,N_921,N_957);
nand U1020 (N_1020,N_920,N_992);
and U1021 (N_1021,N_963,N_975);
nor U1022 (N_1022,N_956,N_979);
nor U1023 (N_1023,N_926,N_985);
nand U1024 (N_1024,N_994,N_910);
and U1025 (N_1025,N_933,N_937);
or U1026 (N_1026,N_942,N_960);
or U1027 (N_1027,N_917,N_936);
or U1028 (N_1028,N_903,N_950);
or U1029 (N_1029,N_962,N_999);
xor U1030 (N_1030,N_922,N_914);
xor U1031 (N_1031,N_919,N_971);
or U1032 (N_1032,N_947,N_978);
nor U1033 (N_1033,N_939,N_988);
and U1034 (N_1034,N_932,N_958);
nand U1035 (N_1035,N_929,N_982);
and U1036 (N_1036,N_905,N_924);
and U1037 (N_1037,N_902,N_951);
nor U1038 (N_1038,N_980,N_911);
nor U1039 (N_1039,N_953,N_995);
nand U1040 (N_1040,N_968,N_989);
nor U1041 (N_1041,N_946,N_949);
xnor U1042 (N_1042,N_986,N_983);
xnor U1043 (N_1043,N_991,N_967);
nor U1044 (N_1044,N_964,N_909);
nor U1045 (N_1045,N_941,N_954);
or U1046 (N_1046,N_915,N_977);
or U1047 (N_1047,N_984,N_923);
nor U1048 (N_1048,N_918,N_981);
or U1049 (N_1049,N_996,N_925);
and U1050 (N_1050,N_901,N_952);
nand U1051 (N_1051,N_951,N_948);
or U1052 (N_1052,N_907,N_909);
and U1053 (N_1053,N_952,N_924);
xor U1054 (N_1054,N_998,N_914);
or U1055 (N_1055,N_996,N_916);
nand U1056 (N_1056,N_900,N_979);
nand U1057 (N_1057,N_965,N_934);
nor U1058 (N_1058,N_923,N_959);
nor U1059 (N_1059,N_956,N_911);
and U1060 (N_1060,N_924,N_999);
nand U1061 (N_1061,N_990,N_904);
nor U1062 (N_1062,N_930,N_948);
or U1063 (N_1063,N_992,N_908);
nor U1064 (N_1064,N_910,N_940);
and U1065 (N_1065,N_980,N_906);
nor U1066 (N_1066,N_926,N_953);
or U1067 (N_1067,N_937,N_965);
or U1068 (N_1068,N_984,N_945);
nor U1069 (N_1069,N_990,N_994);
and U1070 (N_1070,N_998,N_954);
nand U1071 (N_1071,N_994,N_931);
or U1072 (N_1072,N_995,N_917);
nand U1073 (N_1073,N_913,N_938);
or U1074 (N_1074,N_973,N_941);
and U1075 (N_1075,N_940,N_926);
nor U1076 (N_1076,N_956,N_903);
nor U1077 (N_1077,N_992,N_914);
xor U1078 (N_1078,N_943,N_979);
nor U1079 (N_1079,N_941,N_938);
nand U1080 (N_1080,N_904,N_991);
xnor U1081 (N_1081,N_917,N_946);
nor U1082 (N_1082,N_928,N_933);
or U1083 (N_1083,N_947,N_934);
nor U1084 (N_1084,N_994,N_975);
xnor U1085 (N_1085,N_919,N_901);
and U1086 (N_1086,N_937,N_926);
and U1087 (N_1087,N_947,N_913);
or U1088 (N_1088,N_988,N_953);
nand U1089 (N_1089,N_967,N_988);
nor U1090 (N_1090,N_913,N_914);
nand U1091 (N_1091,N_918,N_941);
and U1092 (N_1092,N_979,N_974);
and U1093 (N_1093,N_951,N_963);
nor U1094 (N_1094,N_936,N_940);
xor U1095 (N_1095,N_977,N_944);
nand U1096 (N_1096,N_992,N_964);
nand U1097 (N_1097,N_976,N_910);
xor U1098 (N_1098,N_949,N_950);
xnor U1099 (N_1099,N_916,N_959);
nor U1100 (N_1100,N_1098,N_1016);
nand U1101 (N_1101,N_1087,N_1031);
and U1102 (N_1102,N_1083,N_1091);
nand U1103 (N_1103,N_1063,N_1064);
xnor U1104 (N_1104,N_1092,N_1096);
nand U1105 (N_1105,N_1055,N_1034);
and U1106 (N_1106,N_1088,N_1057);
or U1107 (N_1107,N_1067,N_1068);
or U1108 (N_1108,N_1081,N_1053);
nand U1109 (N_1109,N_1089,N_1086);
or U1110 (N_1110,N_1022,N_1026);
and U1111 (N_1111,N_1090,N_1014);
and U1112 (N_1112,N_1069,N_1006);
xnor U1113 (N_1113,N_1077,N_1038);
and U1114 (N_1114,N_1076,N_1079);
nand U1115 (N_1115,N_1017,N_1033);
nand U1116 (N_1116,N_1070,N_1048);
and U1117 (N_1117,N_1060,N_1001);
xor U1118 (N_1118,N_1036,N_1042);
nand U1119 (N_1119,N_1099,N_1093);
nand U1120 (N_1120,N_1084,N_1052);
and U1121 (N_1121,N_1015,N_1012);
nor U1122 (N_1122,N_1002,N_1085);
nor U1123 (N_1123,N_1075,N_1065);
nand U1124 (N_1124,N_1024,N_1020);
xor U1125 (N_1125,N_1018,N_1032);
xor U1126 (N_1126,N_1061,N_1005);
xor U1127 (N_1127,N_1045,N_1013);
nor U1128 (N_1128,N_1027,N_1043);
xnor U1129 (N_1129,N_1000,N_1044);
and U1130 (N_1130,N_1058,N_1025);
or U1131 (N_1131,N_1008,N_1011);
and U1132 (N_1132,N_1019,N_1059);
and U1133 (N_1133,N_1073,N_1041);
or U1134 (N_1134,N_1050,N_1078);
xor U1135 (N_1135,N_1097,N_1094);
xor U1136 (N_1136,N_1074,N_1054);
nand U1137 (N_1137,N_1004,N_1066);
and U1138 (N_1138,N_1049,N_1072);
xor U1139 (N_1139,N_1095,N_1003);
nand U1140 (N_1140,N_1035,N_1007);
xor U1141 (N_1141,N_1051,N_1062);
nand U1142 (N_1142,N_1046,N_1030);
and U1143 (N_1143,N_1028,N_1071);
nor U1144 (N_1144,N_1009,N_1021);
and U1145 (N_1145,N_1023,N_1056);
nor U1146 (N_1146,N_1010,N_1040);
nor U1147 (N_1147,N_1082,N_1039);
nand U1148 (N_1148,N_1080,N_1037);
or U1149 (N_1149,N_1029,N_1047);
nor U1150 (N_1150,N_1081,N_1093);
xnor U1151 (N_1151,N_1029,N_1017);
or U1152 (N_1152,N_1021,N_1064);
nor U1153 (N_1153,N_1048,N_1011);
nand U1154 (N_1154,N_1008,N_1069);
xor U1155 (N_1155,N_1084,N_1021);
xnor U1156 (N_1156,N_1042,N_1086);
nand U1157 (N_1157,N_1089,N_1085);
nand U1158 (N_1158,N_1014,N_1087);
xnor U1159 (N_1159,N_1089,N_1064);
nand U1160 (N_1160,N_1084,N_1079);
and U1161 (N_1161,N_1093,N_1071);
or U1162 (N_1162,N_1010,N_1075);
nand U1163 (N_1163,N_1042,N_1018);
or U1164 (N_1164,N_1075,N_1033);
nor U1165 (N_1165,N_1016,N_1068);
nand U1166 (N_1166,N_1054,N_1066);
or U1167 (N_1167,N_1018,N_1087);
nand U1168 (N_1168,N_1054,N_1069);
or U1169 (N_1169,N_1064,N_1094);
and U1170 (N_1170,N_1061,N_1002);
nor U1171 (N_1171,N_1042,N_1010);
or U1172 (N_1172,N_1001,N_1061);
and U1173 (N_1173,N_1097,N_1000);
nor U1174 (N_1174,N_1023,N_1067);
or U1175 (N_1175,N_1071,N_1034);
nand U1176 (N_1176,N_1036,N_1015);
and U1177 (N_1177,N_1069,N_1041);
and U1178 (N_1178,N_1003,N_1097);
and U1179 (N_1179,N_1070,N_1082);
xnor U1180 (N_1180,N_1073,N_1070);
xnor U1181 (N_1181,N_1044,N_1054);
nor U1182 (N_1182,N_1076,N_1071);
nand U1183 (N_1183,N_1045,N_1014);
or U1184 (N_1184,N_1043,N_1010);
and U1185 (N_1185,N_1060,N_1045);
or U1186 (N_1186,N_1034,N_1050);
xor U1187 (N_1187,N_1042,N_1015);
and U1188 (N_1188,N_1060,N_1019);
xor U1189 (N_1189,N_1015,N_1091);
xnor U1190 (N_1190,N_1082,N_1026);
or U1191 (N_1191,N_1050,N_1066);
nand U1192 (N_1192,N_1046,N_1084);
nor U1193 (N_1193,N_1072,N_1023);
xnor U1194 (N_1194,N_1014,N_1039);
and U1195 (N_1195,N_1056,N_1048);
nand U1196 (N_1196,N_1034,N_1023);
and U1197 (N_1197,N_1004,N_1015);
xor U1198 (N_1198,N_1017,N_1052);
and U1199 (N_1199,N_1059,N_1080);
nand U1200 (N_1200,N_1101,N_1115);
xor U1201 (N_1201,N_1112,N_1151);
nor U1202 (N_1202,N_1150,N_1111);
and U1203 (N_1203,N_1109,N_1195);
or U1204 (N_1204,N_1144,N_1135);
xnor U1205 (N_1205,N_1106,N_1149);
nand U1206 (N_1206,N_1124,N_1136);
xnor U1207 (N_1207,N_1129,N_1110);
nor U1208 (N_1208,N_1103,N_1185);
nand U1209 (N_1209,N_1160,N_1145);
xor U1210 (N_1210,N_1148,N_1137);
nor U1211 (N_1211,N_1133,N_1159);
and U1212 (N_1212,N_1190,N_1198);
nor U1213 (N_1213,N_1139,N_1174);
xor U1214 (N_1214,N_1178,N_1141);
nand U1215 (N_1215,N_1187,N_1119);
nand U1216 (N_1216,N_1177,N_1114);
or U1217 (N_1217,N_1113,N_1171);
or U1218 (N_1218,N_1147,N_1193);
nor U1219 (N_1219,N_1197,N_1140);
and U1220 (N_1220,N_1118,N_1126);
and U1221 (N_1221,N_1123,N_1165);
nor U1222 (N_1222,N_1125,N_1134);
nor U1223 (N_1223,N_1192,N_1131);
or U1224 (N_1224,N_1130,N_1156);
and U1225 (N_1225,N_1180,N_1173);
xnor U1226 (N_1226,N_1116,N_1127);
nand U1227 (N_1227,N_1183,N_1132);
or U1228 (N_1228,N_1152,N_1166);
nand U1229 (N_1229,N_1162,N_1108);
xnor U1230 (N_1230,N_1191,N_1196);
nor U1231 (N_1231,N_1142,N_1102);
and U1232 (N_1232,N_1107,N_1163);
xor U1233 (N_1233,N_1164,N_1188);
nor U1234 (N_1234,N_1167,N_1117);
nand U1235 (N_1235,N_1176,N_1100);
or U1236 (N_1236,N_1128,N_1105);
nor U1237 (N_1237,N_1121,N_1172);
nand U1238 (N_1238,N_1157,N_1186);
and U1239 (N_1239,N_1182,N_1122);
nand U1240 (N_1240,N_1194,N_1169);
nand U1241 (N_1241,N_1168,N_1184);
or U1242 (N_1242,N_1146,N_1158);
and U1243 (N_1243,N_1161,N_1104);
nand U1244 (N_1244,N_1154,N_1170);
and U1245 (N_1245,N_1199,N_1120);
and U1246 (N_1246,N_1155,N_1189);
and U1247 (N_1247,N_1153,N_1143);
nand U1248 (N_1248,N_1175,N_1179);
nand U1249 (N_1249,N_1138,N_1181);
nand U1250 (N_1250,N_1159,N_1122);
nor U1251 (N_1251,N_1154,N_1125);
xnor U1252 (N_1252,N_1102,N_1173);
or U1253 (N_1253,N_1125,N_1111);
xor U1254 (N_1254,N_1135,N_1101);
nor U1255 (N_1255,N_1199,N_1118);
or U1256 (N_1256,N_1176,N_1195);
nor U1257 (N_1257,N_1103,N_1154);
nor U1258 (N_1258,N_1123,N_1103);
nor U1259 (N_1259,N_1116,N_1170);
nor U1260 (N_1260,N_1104,N_1120);
and U1261 (N_1261,N_1111,N_1192);
nor U1262 (N_1262,N_1193,N_1166);
or U1263 (N_1263,N_1177,N_1185);
and U1264 (N_1264,N_1142,N_1144);
xnor U1265 (N_1265,N_1116,N_1131);
nand U1266 (N_1266,N_1149,N_1150);
and U1267 (N_1267,N_1111,N_1155);
nor U1268 (N_1268,N_1137,N_1116);
nor U1269 (N_1269,N_1176,N_1179);
xnor U1270 (N_1270,N_1153,N_1117);
nand U1271 (N_1271,N_1146,N_1105);
nor U1272 (N_1272,N_1179,N_1131);
xor U1273 (N_1273,N_1114,N_1191);
or U1274 (N_1274,N_1100,N_1153);
nor U1275 (N_1275,N_1144,N_1123);
nor U1276 (N_1276,N_1199,N_1102);
xor U1277 (N_1277,N_1147,N_1159);
nor U1278 (N_1278,N_1183,N_1169);
nand U1279 (N_1279,N_1190,N_1168);
nand U1280 (N_1280,N_1158,N_1122);
nand U1281 (N_1281,N_1116,N_1196);
nor U1282 (N_1282,N_1194,N_1198);
and U1283 (N_1283,N_1177,N_1151);
nand U1284 (N_1284,N_1178,N_1172);
and U1285 (N_1285,N_1136,N_1143);
nor U1286 (N_1286,N_1177,N_1127);
and U1287 (N_1287,N_1170,N_1134);
and U1288 (N_1288,N_1176,N_1182);
nand U1289 (N_1289,N_1155,N_1195);
xnor U1290 (N_1290,N_1191,N_1193);
or U1291 (N_1291,N_1115,N_1163);
xor U1292 (N_1292,N_1108,N_1160);
nand U1293 (N_1293,N_1131,N_1173);
or U1294 (N_1294,N_1135,N_1173);
xor U1295 (N_1295,N_1124,N_1171);
nor U1296 (N_1296,N_1158,N_1154);
xnor U1297 (N_1297,N_1129,N_1130);
or U1298 (N_1298,N_1133,N_1137);
or U1299 (N_1299,N_1114,N_1181);
nor U1300 (N_1300,N_1243,N_1242);
and U1301 (N_1301,N_1231,N_1250);
nor U1302 (N_1302,N_1227,N_1294);
xor U1303 (N_1303,N_1272,N_1274);
or U1304 (N_1304,N_1234,N_1251);
or U1305 (N_1305,N_1265,N_1273);
xnor U1306 (N_1306,N_1254,N_1286);
and U1307 (N_1307,N_1223,N_1293);
or U1308 (N_1308,N_1210,N_1233);
and U1309 (N_1309,N_1263,N_1288);
xnor U1310 (N_1310,N_1200,N_1236);
nand U1311 (N_1311,N_1270,N_1228);
nand U1312 (N_1312,N_1252,N_1203);
nor U1313 (N_1313,N_1204,N_1207);
or U1314 (N_1314,N_1298,N_1259);
nor U1315 (N_1315,N_1230,N_1229);
and U1316 (N_1316,N_1261,N_1245);
nor U1317 (N_1317,N_1267,N_1280);
and U1318 (N_1318,N_1283,N_1269);
nand U1319 (N_1319,N_1296,N_1249);
and U1320 (N_1320,N_1277,N_1235);
xor U1321 (N_1321,N_1262,N_1211);
xnor U1322 (N_1322,N_1206,N_1276);
and U1323 (N_1323,N_1297,N_1208);
nor U1324 (N_1324,N_1248,N_1291);
nor U1325 (N_1325,N_1221,N_1258);
and U1326 (N_1326,N_1278,N_1226);
xnor U1327 (N_1327,N_1219,N_1205);
xnor U1328 (N_1328,N_1284,N_1290);
and U1329 (N_1329,N_1253,N_1232);
or U1330 (N_1330,N_1217,N_1260);
or U1331 (N_1331,N_1224,N_1237);
xor U1332 (N_1332,N_1222,N_1268);
and U1333 (N_1333,N_1209,N_1247);
nor U1334 (N_1334,N_1266,N_1295);
and U1335 (N_1335,N_1282,N_1281);
nor U1336 (N_1336,N_1241,N_1289);
xor U1337 (N_1337,N_1271,N_1216);
nand U1338 (N_1338,N_1285,N_1275);
or U1339 (N_1339,N_1218,N_1292);
nor U1340 (N_1340,N_1212,N_1244);
xnor U1341 (N_1341,N_1213,N_1279);
and U1342 (N_1342,N_1255,N_1246);
or U1343 (N_1343,N_1257,N_1220);
nand U1344 (N_1344,N_1239,N_1214);
xor U1345 (N_1345,N_1264,N_1215);
or U1346 (N_1346,N_1201,N_1238);
nor U1347 (N_1347,N_1202,N_1225);
or U1348 (N_1348,N_1287,N_1299);
xnor U1349 (N_1349,N_1256,N_1240);
or U1350 (N_1350,N_1235,N_1268);
nor U1351 (N_1351,N_1270,N_1273);
or U1352 (N_1352,N_1253,N_1251);
and U1353 (N_1353,N_1289,N_1290);
and U1354 (N_1354,N_1210,N_1292);
nor U1355 (N_1355,N_1279,N_1234);
xor U1356 (N_1356,N_1249,N_1265);
nand U1357 (N_1357,N_1279,N_1265);
xnor U1358 (N_1358,N_1294,N_1257);
nor U1359 (N_1359,N_1219,N_1264);
or U1360 (N_1360,N_1224,N_1235);
xor U1361 (N_1361,N_1264,N_1298);
xor U1362 (N_1362,N_1200,N_1219);
xor U1363 (N_1363,N_1247,N_1295);
nor U1364 (N_1364,N_1262,N_1233);
and U1365 (N_1365,N_1234,N_1254);
and U1366 (N_1366,N_1200,N_1204);
or U1367 (N_1367,N_1219,N_1240);
nor U1368 (N_1368,N_1233,N_1279);
or U1369 (N_1369,N_1284,N_1239);
xnor U1370 (N_1370,N_1262,N_1257);
or U1371 (N_1371,N_1256,N_1273);
xnor U1372 (N_1372,N_1275,N_1219);
nor U1373 (N_1373,N_1216,N_1277);
and U1374 (N_1374,N_1232,N_1219);
nand U1375 (N_1375,N_1227,N_1263);
or U1376 (N_1376,N_1274,N_1221);
nand U1377 (N_1377,N_1286,N_1214);
nand U1378 (N_1378,N_1219,N_1222);
xnor U1379 (N_1379,N_1298,N_1268);
or U1380 (N_1380,N_1273,N_1235);
and U1381 (N_1381,N_1258,N_1236);
and U1382 (N_1382,N_1297,N_1249);
and U1383 (N_1383,N_1285,N_1237);
nor U1384 (N_1384,N_1235,N_1209);
or U1385 (N_1385,N_1249,N_1277);
nand U1386 (N_1386,N_1205,N_1268);
or U1387 (N_1387,N_1290,N_1272);
nor U1388 (N_1388,N_1293,N_1235);
and U1389 (N_1389,N_1292,N_1219);
or U1390 (N_1390,N_1265,N_1200);
xnor U1391 (N_1391,N_1243,N_1287);
and U1392 (N_1392,N_1262,N_1272);
nor U1393 (N_1393,N_1207,N_1248);
and U1394 (N_1394,N_1243,N_1294);
xnor U1395 (N_1395,N_1231,N_1235);
or U1396 (N_1396,N_1241,N_1218);
and U1397 (N_1397,N_1218,N_1244);
or U1398 (N_1398,N_1287,N_1271);
nor U1399 (N_1399,N_1229,N_1267);
nor U1400 (N_1400,N_1396,N_1346);
nor U1401 (N_1401,N_1370,N_1390);
nor U1402 (N_1402,N_1395,N_1382);
nand U1403 (N_1403,N_1369,N_1366);
xnor U1404 (N_1404,N_1340,N_1356);
nor U1405 (N_1405,N_1355,N_1373);
xor U1406 (N_1406,N_1361,N_1306);
nor U1407 (N_1407,N_1334,N_1351);
and U1408 (N_1408,N_1399,N_1378);
xnor U1409 (N_1409,N_1342,N_1393);
nor U1410 (N_1410,N_1341,N_1332);
xor U1411 (N_1411,N_1321,N_1364);
and U1412 (N_1412,N_1352,N_1335);
or U1413 (N_1413,N_1329,N_1380);
and U1414 (N_1414,N_1363,N_1338);
nand U1415 (N_1415,N_1319,N_1372);
and U1416 (N_1416,N_1349,N_1314);
nand U1417 (N_1417,N_1337,N_1345);
nor U1418 (N_1418,N_1307,N_1384);
nand U1419 (N_1419,N_1360,N_1339);
xor U1420 (N_1420,N_1347,N_1315);
nand U1421 (N_1421,N_1310,N_1331);
and U1422 (N_1422,N_1381,N_1376);
or U1423 (N_1423,N_1397,N_1377);
nand U1424 (N_1424,N_1316,N_1388);
nand U1425 (N_1425,N_1385,N_1354);
nand U1426 (N_1426,N_1365,N_1322);
xor U1427 (N_1427,N_1398,N_1375);
and U1428 (N_1428,N_1301,N_1300);
and U1429 (N_1429,N_1350,N_1312);
and U1430 (N_1430,N_1368,N_1323);
or U1431 (N_1431,N_1383,N_1386);
xnor U1432 (N_1432,N_1302,N_1327);
xor U1433 (N_1433,N_1320,N_1379);
or U1434 (N_1434,N_1367,N_1371);
xor U1435 (N_1435,N_1305,N_1325);
and U1436 (N_1436,N_1326,N_1308);
nor U1437 (N_1437,N_1311,N_1389);
nand U1438 (N_1438,N_1313,N_1303);
and U1439 (N_1439,N_1391,N_1304);
or U1440 (N_1440,N_1394,N_1362);
nand U1441 (N_1441,N_1348,N_1359);
or U1442 (N_1442,N_1357,N_1330);
xor U1443 (N_1443,N_1324,N_1353);
nor U1444 (N_1444,N_1392,N_1317);
nand U1445 (N_1445,N_1328,N_1387);
nor U1446 (N_1446,N_1358,N_1333);
and U1447 (N_1447,N_1309,N_1318);
nor U1448 (N_1448,N_1374,N_1343);
nor U1449 (N_1449,N_1336,N_1344);
or U1450 (N_1450,N_1303,N_1329);
nand U1451 (N_1451,N_1334,N_1390);
nor U1452 (N_1452,N_1312,N_1377);
or U1453 (N_1453,N_1332,N_1377);
or U1454 (N_1454,N_1318,N_1394);
or U1455 (N_1455,N_1385,N_1346);
and U1456 (N_1456,N_1334,N_1342);
nand U1457 (N_1457,N_1370,N_1355);
and U1458 (N_1458,N_1392,N_1371);
xor U1459 (N_1459,N_1322,N_1328);
and U1460 (N_1460,N_1361,N_1346);
or U1461 (N_1461,N_1353,N_1307);
or U1462 (N_1462,N_1371,N_1348);
xor U1463 (N_1463,N_1319,N_1335);
nor U1464 (N_1464,N_1344,N_1310);
nand U1465 (N_1465,N_1389,N_1398);
or U1466 (N_1466,N_1394,N_1390);
or U1467 (N_1467,N_1301,N_1398);
nand U1468 (N_1468,N_1350,N_1384);
or U1469 (N_1469,N_1332,N_1350);
xor U1470 (N_1470,N_1397,N_1312);
nor U1471 (N_1471,N_1351,N_1324);
nand U1472 (N_1472,N_1383,N_1393);
and U1473 (N_1473,N_1343,N_1303);
or U1474 (N_1474,N_1323,N_1374);
nor U1475 (N_1475,N_1304,N_1378);
or U1476 (N_1476,N_1393,N_1395);
xnor U1477 (N_1477,N_1394,N_1342);
nor U1478 (N_1478,N_1382,N_1310);
nor U1479 (N_1479,N_1355,N_1318);
xor U1480 (N_1480,N_1380,N_1392);
xnor U1481 (N_1481,N_1355,N_1360);
xnor U1482 (N_1482,N_1350,N_1378);
nand U1483 (N_1483,N_1352,N_1316);
xor U1484 (N_1484,N_1393,N_1340);
nand U1485 (N_1485,N_1377,N_1393);
and U1486 (N_1486,N_1366,N_1355);
or U1487 (N_1487,N_1376,N_1355);
nand U1488 (N_1488,N_1376,N_1313);
and U1489 (N_1489,N_1374,N_1386);
xor U1490 (N_1490,N_1341,N_1363);
or U1491 (N_1491,N_1304,N_1366);
nor U1492 (N_1492,N_1326,N_1374);
xnor U1493 (N_1493,N_1318,N_1399);
and U1494 (N_1494,N_1356,N_1305);
and U1495 (N_1495,N_1378,N_1331);
nand U1496 (N_1496,N_1301,N_1333);
or U1497 (N_1497,N_1349,N_1357);
nand U1498 (N_1498,N_1310,N_1343);
nor U1499 (N_1499,N_1346,N_1310);
or U1500 (N_1500,N_1497,N_1480);
nor U1501 (N_1501,N_1447,N_1440);
nor U1502 (N_1502,N_1420,N_1448);
nor U1503 (N_1503,N_1479,N_1494);
xor U1504 (N_1504,N_1462,N_1449);
or U1505 (N_1505,N_1476,N_1438);
or U1506 (N_1506,N_1419,N_1423);
nand U1507 (N_1507,N_1490,N_1445);
or U1508 (N_1508,N_1468,N_1492);
nand U1509 (N_1509,N_1401,N_1416);
or U1510 (N_1510,N_1463,N_1426);
or U1511 (N_1511,N_1433,N_1483);
xnor U1512 (N_1512,N_1487,N_1422);
xnor U1513 (N_1513,N_1495,N_1457);
and U1514 (N_1514,N_1417,N_1439);
or U1515 (N_1515,N_1436,N_1407);
xnor U1516 (N_1516,N_1486,N_1460);
nand U1517 (N_1517,N_1435,N_1405);
nor U1518 (N_1518,N_1499,N_1446);
nor U1519 (N_1519,N_1465,N_1461);
or U1520 (N_1520,N_1451,N_1458);
nor U1521 (N_1521,N_1471,N_1418);
nand U1522 (N_1522,N_1474,N_1482);
nor U1523 (N_1523,N_1441,N_1469);
nand U1524 (N_1524,N_1489,N_1477);
or U1525 (N_1525,N_1466,N_1475);
nor U1526 (N_1526,N_1430,N_1484);
and U1527 (N_1527,N_1481,N_1455);
and U1528 (N_1528,N_1444,N_1425);
xnor U1529 (N_1529,N_1453,N_1403);
or U1530 (N_1530,N_1456,N_1434);
nor U1531 (N_1531,N_1424,N_1415);
or U1532 (N_1532,N_1450,N_1409);
or U1533 (N_1533,N_1454,N_1431);
or U1534 (N_1534,N_1443,N_1437);
or U1535 (N_1535,N_1411,N_1421);
nand U1536 (N_1536,N_1464,N_1413);
and U1537 (N_1537,N_1442,N_1412);
or U1538 (N_1538,N_1491,N_1428);
xnor U1539 (N_1539,N_1485,N_1452);
or U1540 (N_1540,N_1470,N_1427);
and U1541 (N_1541,N_1472,N_1402);
and U1542 (N_1542,N_1488,N_1406);
nor U1543 (N_1543,N_1459,N_1414);
xor U1544 (N_1544,N_1408,N_1410);
or U1545 (N_1545,N_1498,N_1478);
nor U1546 (N_1546,N_1432,N_1473);
xor U1547 (N_1547,N_1467,N_1496);
nor U1548 (N_1548,N_1493,N_1400);
or U1549 (N_1549,N_1429,N_1404);
xor U1550 (N_1550,N_1427,N_1486);
and U1551 (N_1551,N_1462,N_1407);
nand U1552 (N_1552,N_1435,N_1495);
xnor U1553 (N_1553,N_1448,N_1426);
and U1554 (N_1554,N_1494,N_1445);
or U1555 (N_1555,N_1440,N_1490);
xor U1556 (N_1556,N_1451,N_1461);
and U1557 (N_1557,N_1480,N_1459);
xnor U1558 (N_1558,N_1467,N_1474);
nor U1559 (N_1559,N_1471,N_1462);
and U1560 (N_1560,N_1476,N_1457);
xor U1561 (N_1561,N_1486,N_1498);
xor U1562 (N_1562,N_1426,N_1418);
nor U1563 (N_1563,N_1429,N_1415);
or U1564 (N_1564,N_1421,N_1462);
nand U1565 (N_1565,N_1433,N_1451);
and U1566 (N_1566,N_1455,N_1454);
xnor U1567 (N_1567,N_1438,N_1478);
and U1568 (N_1568,N_1400,N_1489);
and U1569 (N_1569,N_1427,N_1465);
or U1570 (N_1570,N_1434,N_1477);
xnor U1571 (N_1571,N_1484,N_1413);
or U1572 (N_1572,N_1413,N_1451);
or U1573 (N_1573,N_1432,N_1493);
or U1574 (N_1574,N_1412,N_1438);
nor U1575 (N_1575,N_1420,N_1404);
xor U1576 (N_1576,N_1410,N_1411);
or U1577 (N_1577,N_1411,N_1445);
xnor U1578 (N_1578,N_1438,N_1475);
xor U1579 (N_1579,N_1424,N_1439);
or U1580 (N_1580,N_1471,N_1465);
xnor U1581 (N_1581,N_1491,N_1417);
and U1582 (N_1582,N_1440,N_1477);
nand U1583 (N_1583,N_1416,N_1417);
and U1584 (N_1584,N_1487,N_1474);
xor U1585 (N_1585,N_1469,N_1495);
or U1586 (N_1586,N_1444,N_1450);
nor U1587 (N_1587,N_1455,N_1476);
nand U1588 (N_1588,N_1426,N_1415);
or U1589 (N_1589,N_1486,N_1418);
nand U1590 (N_1590,N_1452,N_1469);
xnor U1591 (N_1591,N_1400,N_1440);
nand U1592 (N_1592,N_1474,N_1419);
nor U1593 (N_1593,N_1489,N_1452);
xor U1594 (N_1594,N_1477,N_1454);
and U1595 (N_1595,N_1485,N_1470);
xnor U1596 (N_1596,N_1464,N_1438);
or U1597 (N_1597,N_1490,N_1408);
nand U1598 (N_1598,N_1487,N_1460);
nor U1599 (N_1599,N_1473,N_1450);
nor U1600 (N_1600,N_1588,N_1553);
and U1601 (N_1601,N_1591,N_1572);
or U1602 (N_1602,N_1534,N_1501);
nand U1603 (N_1603,N_1571,N_1516);
or U1604 (N_1604,N_1586,N_1511);
and U1605 (N_1605,N_1543,N_1545);
nor U1606 (N_1606,N_1554,N_1584);
xor U1607 (N_1607,N_1559,N_1592);
nor U1608 (N_1608,N_1564,N_1565);
and U1609 (N_1609,N_1529,N_1527);
nand U1610 (N_1610,N_1575,N_1558);
nand U1611 (N_1611,N_1519,N_1552);
nor U1612 (N_1612,N_1585,N_1589);
nor U1613 (N_1613,N_1518,N_1582);
or U1614 (N_1614,N_1581,N_1544);
xor U1615 (N_1615,N_1583,N_1557);
or U1616 (N_1616,N_1576,N_1577);
and U1617 (N_1617,N_1566,N_1508);
xnor U1618 (N_1618,N_1512,N_1547);
and U1619 (N_1619,N_1533,N_1517);
nand U1620 (N_1620,N_1541,N_1530);
and U1621 (N_1621,N_1567,N_1574);
nand U1622 (N_1622,N_1509,N_1590);
nor U1623 (N_1623,N_1546,N_1521);
nor U1624 (N_1624,N_1536,N_1526);
nand U1625 (N_1625,N_1555,N_1548);
xnor U1626 (N_1626,N_1515,N_1513);
nor U1627 (N_1627,N_1596,N_1579);
nor U1628 (N_1628,N_1549,N_1510);
or U1629 (N_1629,N_1525,N_1522);
nand U1630 (N_1630,N_1550,N_1524);
and U1631 (N_1631,N_1540,N_1504);
nor U1632 (N_1632,N_1560,N_1563);
or U1633 (N_1633,N_1505,N_1503);
nor U1634 (N_1634,N_1556,N_1531);
or U1635 (N_1635,N_1593,N_1562);
nor U1636 (N_1636,N_1580,N_1595);
or U1637 (N_1637,N_1535,N_1500);
nand U1638 (N_1638,N_1597,N_1507);
and U1639 (N_1639,N_1528,N_1538);
xor U1640 (N_1640,N_1570,N_1514);
nand U1641 (N_1641,N_1506,N_1532);
or U1642 (N_1642,N_1523,N_1520);
and U1643 (N_1643,N_1594,N_1587);
nor U1644 (N_1644,N_1568,N_1578);
nand U1645 (N_1645,N_1569,N_1551);
nor U1646 (N_1646,N_1573,N_1561);
and U1647 (N_1647,N_1542,N_1599);
and U1648 (N_1648,N_1537,N_1502);
nor U1649 (N_1649,N_1598,N_1539);
xnor U1650 (N_1650,N_1590,N_1521);
xor U1651 (N_1651,N_1523,N_1579);
xor U1652 (N_1652,N_1567,N_1503);
nor U1653 (N_1653,N_1598,N_1555);
xnor U1654 (N_1654,N_1509,N_1529);
or U1655 (N_1655,N_1517,N_1514);
nand U1656 (N_1656,N_1506,N_1545);
nor U1657 (N_1657,N_1506,N_1527);
nor U1658 (N_1658,N_1593,N_1594);
nor U1659 (N_1659,N_1550,N_1583);
nand U1660 (N_1660,N_1567,N_1512);
and U1661 (N_1661,N_1500,N_1528);
and U1662 (N_1662,N_1526,N_1540);
and U1663 (N_1663,N_1554,N_1590);
and U1664 (N_1664,N_1556,N_1530);
nor U1665 (N_1665,N_1547,N_1532);
nand U1666 (N_1666,N_1591,N_1598);
nor U1667 (N_1667,N_1574,N_1553);
nor U1668 (N_1668,N_1595,N_1582);
xor U1669 (N_1669,N_1552,N_1516);
nor U1670 (N_1670,N_1537,N_1531);
and U1671 (N_1671,N_1596,N_1534);
or U1672 (N_1672,N_1593,N_1571);
nand U1673 (N_1673,N_1540,N_1512);
and U1674 (N_1674,N_1523,N_1502);
or U1675 (N_1675,N_1555,N_1576);
nand U1676 (N_1676,N_1593,N_1504);
nor U1677 (N_1677,N_1549,N_1563);
xnor U1678 (N_1678,N_1524,N_1549);
and U1679 (N_1679,N_1562,N_1590);
xor U1680 (N_1680,N_1561,N_1517);
nand U1681 (N_1681,N_1552,N_1513);
and U1682 (N_1682,N_1528,N_1540);
nand U1683 (N_1683,N_1548,N_1568);
nand U1684 (N_1684,N_1577,N_1514);
nand U1685 (N_1685,N_1558,N_1576);
and U1686 (N_1686,N_1517,N_1593);
nand U1687 (N_1687,N_1572,N_1574);
nor U1688 (N_1688,N_1510,N_1572);
nor U1689 (N_1689,N_1548,N_1537);
nand U1690 (N_1690,N_1508,N_1546);
or U1691 (N_1691,N_1547,N_1587);
or U1692 (N_1692,N_1501,N_1567);
nand U1693 (N_1693,N_1543,N_1566);
or U1694 (N_1694,N_1517,N_1503);
xor U1695 (N_1695,N_1594,N_1551);
and U1696 (N_1696,N_1523,N_1545);
nand U1697 (N_1697,N_1512,N_1554);
nand U1698 (N_1698,N_1591,N_1502);
and U1699 (N_1699,N_1506,N_1566);
xnor U1700 (N_1700,N_1665,N_1630);
and U1701 (N_1701,N_1603,N_1681);
nand U1702 (N_1702,N_1628,N_1656);
or U1703 (N_1703,N_1644,N_1674);
xor U1704 (N_1704,N_1649,N_1671);
nor U1705 (N_1705,N_1648,N_1608);
or U1706 (N_1706,N_1660,N_1658);
and U1707 (N_1707,N_1634,N_1633);
xor U1708 (N_1708,N_1646,N_1676);
xnor U1709 (N_1709,N_1638,N_1667);
nand U1710 (N_1710,N_1695,N_1659);
nand U1711 (N_1711,N_1618,N_1636);
nand U1712 (N_1712,N_1631,N_1621);
or U1713 (N_1713,N_1668,N_1664);
and U1714 (N_1714,N_1647,N_1645);
and U1715 (N_1715,N_1690,N_1696);
nand U1716 (N_1716,N_1652,N_1611);
nor U1717 (N_1717,N_1672,N_1657);
and U1718 (N_1718,N_1691,N_1605);
or U1719 (N_1719,N_1686,N_1625);
nand U1720 (N_1720,N_1688,N_1643);
or U1721 (N_1721,N_1602,N_1600);
and U1722 (N_1722,N_1612,N_1616);
nor U1723 (N_1723,N_1609,N_1615);
xor U1724 (N_1724,N_1626,N_1639);
nor U1725 (N_1725,N_1607,N_1683);
nor U1726 (N_1726,N_1629,N_1679);
nand U1727 (N_1727,N_1669,N_1617);
nor U1728 (N_1728,N_1640,N_1651);
nor U1729 (N_1729,N_1613,N_1662);
or U1730 (N_1730,N_1689,N_1624);
and U1731 (N_1731,N_1601,N_1675);
or U1732 (N_1732,N_1632,N_1677);
and U1733 (N_1733,N_1698,N_1673);
xnor U1734 (N_1734,N_1614,N_1682);
nand U1735 (N_1735,N_1692,N_1661);
and U1736 (N_1736,N_1687,N_1642);
xor U1737 (N_1737,N_1685,N_1655);
and U1738 (N_1738,N_1637,N_1606);
and U1739 (N_1739,N_1678,N_1684);
nor U1740 (N_1740,N_1627,N_1663);
or U1741 (N_1741,N_1654,N_1635);
nor U1742 (N_1742,N_1604,N_1697);
xor U1743 (N_1743,N_1670,N_1620);
and U1744 (N_1744,N_1610,N_1666);
nor U1745 (N_1745,N_1623,N_1680);
nor U1746 (N_1746,N_1641,N_1653);
or U1747 (N_1747,N_1699,N_1619);
xnor U1748 (N_1748,N_1694,N_1693);
and U1749 (N_1749,N_1622,N_1650);
nor U1750 (N_1750,N_1661,N_1697);
nor U1751 (N_1751,N_1668,N_1673);
nor U1752 (N_1752,N_1698,N_1662);
and U1753 (N_1753,N_1616,N_1646);
or U1754 (N_1754,N_1686,N_1665);
xnor U1755 (N_1755,N_1666,N_1678);
nor U1756 (N_1756,N_1698,N_1692);
or U1757 (N_1757,N_1655,N_1687);
nand U1758 (N_1758,N_1603,N_1660);
nand U1759 (N_1759,N_1638,N_1622);
nand U1760 (N_1760,N_1666,N_1620);
nor U1761 (N_1761,N_1692,N_1626);
xnor U1762 (N_1762,N_1664,N_1602);
nand U1763 (N_1763,N_1693,N_1644);
nor U1764 (N_1764,N_1667,N_1665);
or U1765 (N_1765,N_1647,N_1698);
xnor U1766 (N_1766,N_1610,N_1637);
xnor U1767 (N_1767,N_1695,N_1696);
nand U1768 (N_1768,N_1601,N_1688);
or U1769 (N_1769,N_1680,N_1666);
and U1770 (N_1770,N_1651,N_1606);
nand U1771 (N_1771,N_1662,N_1690);
or U1772 (N_1772,N_1626,N_1699);
and U1773 (N_1773,N_1619,N_1634);
nor U1774 (N_1774,N_1617,N_1689);
and U1775 (N_1775,N_1627,N_1618);
nand U1776 (N_1776,N_1619,N_1665);
or U1777 (N_1777,N_1664,N_1646);
nor U1778 (N_1778,N_1608,N_1680);
xor U1779 (N_1779,N_1653,N_1628);
nor U1780 (N_1780,N_1678,N_1617);
and U1781 (N_1781,N_1627,N_1694);
xor U1782 (N_1782,N_1609,N_1623);
or U1783 (N_1783,N_1644,N_1688);
nor U1784 (N_1784,N_1694,N_1626);
xnor U1785 (N_1785,N_1624,N_1664);
and U1786 (N_1786,N_1675,N_1644);
or U1787 (N_1787,N_1602,N_1663);
xnor U1788 (N_1788,N_1697,N_1626);
and U1789 (N_1789,N_1657,N_1677);
nor U1790 (N_1790,N_1631,N_1672);
or U1791 (N_1791,N_1644,N_1686);
and U1792 (N_1792,N_1674,N_1655);
or U1793 (N_1793,N_1657,N_1642);
nand U1794 (N_1794,N_1693,N_1683);
xnor U1795 (N_1795,N_1683,N_1652);
and U1796 (N_1796,N_1644,N_1634);
xor U1797 (N_1797,N_1611,N_1622);
nand U1798 (N_1798,N_1615,N_1629);
nand U1799 (N_1799,N_1608,N_1687);
or U1800 (N_1800,N_1773,N_1766);
nand U1801 (N_1801,N_1748,N_1732);
xor U1802 (N_1802,N_1775,N_1763);
xnor U1803 (N_1803,N_1781,N_1795);
nor U1804 (N_1804,N_1799,N_1724);
and U1805 (N_1805,N_1790,N_1741);
nand U1806 (N_1806,N_1780,N_1735);
xnor U1807 (N_1807,N_1788,N_1752);
and U1808 (N_1808,N_1722,N_1747);
nand U1809 (N_1809,N_1708,N_1789);
nand U1810 (N_1810,N_1716,N_1756);
nor U1811 (N_1811,N_1729,N_1743);
xor U1812 (N_1812,N_1737,N_1719);
or U1813 (N_1813,N_1726,N_1755);
or U1814 (N_1814,N_1721,N_1717);
nand U1815 (N_1815,N_1706,N_1768);
xor U1816 (N_1816,N_1749,N_1778);
nor U1817 (N_1817,N_1711,N_1727);
nand U1818 (N_1818,N_1715,N_1776);
nor U1819 (N_1819,N_1734,N_1760);
nand U1820 (N_1820,N_1725,N_1736);
nand U1821 (N_1821,N_1797,N_1786);
and U1822 (N_1822,N_1731,N_1718);
and U1823 (N_1823,N_1779,N_1701);
xnor U1824 (N_1824,N_1770,N_1787);
and U1825 (N_1825,N_1753,N_1709);
nand U1826 (N_1826,N_1771,N_1772);
xnor U1827 (N_1827,N_1744,N_1769);
nor U1828 (N_1828,N_1762,N_1767);
or U1829 (N_1829,N_1746,N_1782);
and U1830 (N_1830,N_1728,N_1792);
nor U1831 (N_1831,N_1798,N_1785);
nand U1832 (N_1832,N_1751,N_1740);
xor U1833 (N_1833,N_1713,N_1704);
xor U1834 (N_1834,N_1700,N_1730);
nor U1835 (N_1835,N_1742,N_1777);
and U1836 (N_1836,N_1765,N_1796);
xor U1837 (N_1837,N_1703,N_1793);
xor U1838 (N_1838,N_1794,N_1738);
nand U1839 (N_1839,N_1710,N_1745);
and U1840 (N_1840,N_1739,N_1733);
and U1841 (N_1841,N_1714,N_1783);
xnor U1842 (N_1842,N_1720,N_1712);
nor U1843 (N_1843,N_1761,N_1784);
xor U1844 (N_1844,N_1723,N_1758);
nor U1845 (N_1845,N_1774,N_1750);
nor U1846 (N_1846,N_1707,N_1757);
xnor U1847 (N_1847,N_1764,N_1759);
nand U1848 (N_1848,N_1705,N_1791);
nand U1849 (N_1849,N_1702,N_1754);
and U1850 (N_1850,N_1743,N_1742);
nand U1851 (N_1851,N_1702,N_1792);
xor U1852 (N_1852,N_1711,N_1728);
and U1853 (N_1853,N_1778,N_1709);
and U1854 (N_1854,N_1781,N_1717);
and U1855 (N_1855,N_1739,N_1757);
and U1856 (N_1856,N_1771,N_1784);
or U1857 (N_1857,N_1780,N_1706);
xnor U1858 (N_1858,N_1716,N_1753);
nor U1859 (N_1859,N_1727,N_1756);
and U1860 (N_1860,N_1714,N_1756);
or U1861 (N_1861,N_1778,N_1751);
or U1862 (N_1862,N_1781,N_1734);
or U1863 (N_1863,N_1749,N_1713);
nand U1864 (N_1864,N_1740,N_1728);
nand U1865 (N_1865,N_1712,N_1793);
nor U1866 (N_1866,N_1720,N_1791);
nor U1867 (N_1867,N_1782,N_1715);
nor U1868 (N_1868,N_1710,N_1790);
or U1869 (N_1869,N_1771,N_1726);
and U1870 (N_1870,N_1741,N_1774);
nand U1871 (N_1871,N_1721,N_1742);
and U1872 (N_1872,N_1717,N_1736);
or U1873 (N_1873,N_1758,N_1743);
nand U1874 (N_1874,N_1774,N_1752);
nor U1875 (N_1875,N_1770,N_1749);
xor U1876 (N_1876,N_1700,N_1701);
or U1877 (N_1877,N_1795,N_1789);
nand U1878 (N_1878,N_1702,N_1773);
xnor U1879 (N_1879,N_1792,N_1753);
and U1880 (N_1880,N_1742,N_1700);
nand U1881 (N_1881,N_1720,N_1721);
or U1882 (N_1882,N_1745,N_1727);
xor U1883 (N_1883,N_1702,N_1727);
nand U1884 (N_1884,N_1758,N_1764);
and U1885 (N_1885,N_1724,N_1747);
nor U1886 (N_1886,N_1729,N_1754);
and U1887 (N_1887,N_1789,N_1703);
xor U1888 (N_1888,N_1764,N_1726);
nor U1889 (N_1889,N_1773,N_1768);
xnor U1890 (N_1890,N_1777,N_1770);
nor U1891 (N_1891,N_1737,N_1708);
and U1892 (N_1892,N_1789,N_1713);
or U1893 (N_1893,N_1700,N_1798);
nor U1894 (N_1894,N_1751,N_1729);
xnor U1895 (N_1895,N_1725,N_1778);
or U1896 (N_1896,N_1726,N_1700);
or U1897 (N_1897,N_1787,N_1723);
nor U1898 (N_1898,N_1720,N_1705);
xor U1899 (N_1899,N_1713,N_1745);
nand U1900 (N_1900,N_1804,N_1824);
nand U1901 (N_1901,N_1807,N_1815);
xor U1902 (N_1902,N_1868,N_1858);
xor U1903 (N_1903,N_1846,N_1895);
or U1904 (N_1904,N_1898,N_1866);
nand U1905 (N_1905,N_1844,N_1826);
xor U1906 (N_1906,N_1878,N_1876);
or U1907 (N_1907,N_1862,N_1819);
nand U1908 (N_1908,N_1861,N_1872);
and U1909 (N_1909,N_1889,N_1892);
nor U1910 (N_1910,N_1829,N_1883);
nor U1911 (N_1911,N_1870,N_1837);
or U1912 (N_1912,N_1896,N_1809);
or U1913 (N_1913,N_1875,N_1882);
nor U1914 (N_1914,N_1843,N_1893);
or U1915 (N_1915,N_1820,N_1802);
or U1916 (N_1916,N_1888,N_1849);
and U1917 (N_1917,N_1836,N_1814);
or U1918 (N_1918,N_1884,N_1856);
nand U1919 (N_1919,N_1874,N_1854);
and U1920 (N_1920,N_1812,N_1801);
and U1921 (N_1921,N_1833,N_1886);
and U1922 (N_1922,N_1879,N_1852);
nor U1923 (N_1923,N_1851,N_1871);
and U1924 (N_1924,N_1873,N_1890);
nand U1925 (N_1925,N_1841,N_1877);
or U1926 (N_1926,N_1897,N_1865);
nand U1927 (N_1927,N_1828,N_1887);
nor U1928 (N_1928,N_1821,N_1853);
and U1929 (N_1929,N_1832,N_1827);
nor U1930 (N_1930,N_1811,N_1848);
or U1931 (N_1931,N_1803,N_1806);
nand U1932 (N_1932,N_1891,N_1805);
and U1933 (N_1933,N_1830,N_1899);
and U1934 (N_1934,N_1818,N_1855);
xnor U1935 (N_1935,N_1880,N_1869);
nand U1936 (N_1936,N_1822,N_1838);
xnor U1937 (N_1937,N_1867,N_1885);
nand U1938 (N_1938,N_1810,N_1860);
and U1939 (N_1939,N_1842,N_1859);
nand U1940 (N_1940,N_1857,N_1808);
or U1941 (N_1941,N_1839,N_1840);
xor U1942 (N_1942,N_1834,N_1831);
nand U1943 (N_1943,N_1825,N_1817);
nand U1944 (N_1944,N_1813,N_1847);
and U1945 (N_1945,N_1850,N_1845);
and U1946 (N_1946,N_1894,N_1835);
nand U1947 (N_1947,N_1800,N_1823);
nand U1948 (N_1948,N_1816,N_1863);
nor U1949 (N_1949,N_1864,N_1881);
xnor U1950 (N_1950,N_1876,N_1872);
and U1951 (N_1951,N_1823,N_1850);
nand U1952 (N_1952,N_1834,N_1849);
nor U1953 (N_1953,N_1827,N_1802);
and U1954 (N_1954,N_1885,N_1854);
or U1955 (N_1955,N_1806,N_1814);
nor U1956 (N_1956,N_1885,N_1801);
nand U1957 (N_1957,N_1899,N_1829);
nand U1958 (N_1958,N_1848,N_1832);
xnor U1959 (N_1959,N_1899,N_1890);
nor U1960 (N_1960,N_1890,N_1836);
and U1961 (N_1961,N_1859,N_1885);
and U1962 (N_1962,N_1841,N_1892);
and U1963 (N_1963,N_1819,N_1877);
and U1964 (N_1964,N_1801,N_1841);
and U1965 (N_1965,N_1808,N_1869);
nand U1966 (N_1966,N_1817,N_1898);
xor U1967 (N_1967,N_1859,N_1873);
nor U1968 (N_1968,N_1883,N_1825);
nand U1969 (N_1969,N_1830,N_1859);
nor U1970 (N_1970,N_1874,N_1872);
nand U1971 (N_1971,N_1827,N_1846);
or U1972 (N_1972,N_1855,N_1830);
or U1973 (N_1973,N_1803,N_1841);
xor U1974 (N_1974,N_1851,N_1897);
and U1975 (N_1975,N_1831,N_1808);
xnor U1976 (N_1976,N_1857,N_1813);
nor U1977 (N_1977,N_1841,N_1872);
or U1978 (N_1978,N_1817,N_1869);
nand U1979 (N_1979,N_1857,N_1872);
and U1980 (N_1980,N_1895,N_1823);
nor U1981 (N_1981,N_1823,N_1813);
nor U1982 (N_1982,N_1849,N_1889);
nor U1983 (N_1983,N_1833,N_1820);
or U1984 (N_1984,N_1818,N_1850);
and U1985 (N_1985,N_1848,N_1867);
and U1986 (N_1986,N_1896,N_1842);
nor U1987 (N_1987,N_1882,N_1888);
and U1988 (N_1988,N_1846,N_1836);
and U1989 (N_1989,N_1816,N_1874);
nand U1990 (N_1990,N_1894,N_1828);
or U1991 (N_1991,N_1878,N_1832);
xor U1992 (N_1992,N_1811,N_1818);
nand U1993 (N_1993,N_1804,N_1831);
nand U1994 (N_1994,N_1850,N_1827);
or U1995 (N_1995,N_1860,N_1802);
nor U1996 (N_1996,N_1895,N_1892);
nand U1997 (N_1997,N_1854,N_1898);
or U1998 (N_1998,N_1857,N_1890);
nand U1999 (N_1999,N_1844,N_1810);
and U2000 (N_2000,N_1909,N_1922);
and U2001 (N_2001,N_1932,N_1993);
xor U2002 (N_2002,N_1940,N_1926);
or U2003 (N_2003,N_1924,N_1937);
xor U2004 (N_2004,N_1930,N_1989);
and U2005 (N_2005,N_1929,N_1950);
xnor U2006 (N_2006,N_1910,N_1935);
nand U2007 (N_2007,N_1980,N_1971);
nand U2008 (N_2008,N_1943,N_1942);
and U2009 (N_2009,N_1988,N_1976);
or U2010 (N_2010,N_1961,N_1965);
nor U2011 (N_2011,N_1949,N_1933);
nor U2012 (N_2012,N_1995,N_1906);
xnor U2013 (N_2013,N_1948,N_1954);
xnor U2014 (N_2014,N_1928,N_1915);
nand U2015 (N_2015,N_1964,N_1962);
or U2016 (N_2016,N_1939,N_1905);
xnor U2017 (N_2017,N_1904,N_1934);
xnor U2018 (N_2018,N_1912,N_1984);
nand U2019 (N_2019,N_1990,N_1955);
or U2020 (N_2020,N_1913,N_1973);
nor U2021 (N_2021,N_1936,N_1956);
xor U2022 (N_2022,N_1947,N_1959);
nor U2023 (N_2023,N_1979,N_1917);
nand U2024 (N_2024,N_1946,N_1966);
or U2025 (N_2025,N_1914,N_1941);
nand U2026 (N_2026,N_1970,N_1911);
or U2027 (N_2027,N_1997,N_1921);
or U2028 (N_2028,N_1983,N_1919);
nand U2029 (N_2029,N_1944,N_1953);
xor U2030 (N_2030,N_1952,N_1972);
nand U2031 (N_2031,N_1969,N_1938);
xor U2032 (N_2032,N_1927,N_1902);
nor U2033 (N_2033,N_1974,N_1987);
nand U2034 (N_2034,N_1978,N_1907);
nand U2035 (N_2035,N_1931,N_1901);
nand U2036 (N_2036,N_1908,N_1918);
nor U2037 (N_2037,N_1996,N_1903);
or U2038 (N_2038,N_1991,N_1900);
or U2039 (N_2039,N_1998,N_1985);
nor U2040 (N_2040,N_1982,N_1923);
or U2041 (N_2041,N_1975,N_1958);
or U2042 (N_2042,N_1968,N_1981);
nor U2043 (N_2043,N_1925,N_1986);
nand U2044 (N_2044,N_1977,N_1967);
nand U2045 (N_2045,N_1951,N_1945);
nand U2046 (N_2046,N_1916,N_1999);
nor U2047 (N_2047,N_1994,N_1960);
xnor U2048 (N_2048,N_1992,N_1920);
and U2049 (N_2049,N_1957,N_1963);
or U2050 (N_2050,N_1909,N_1963);
nor U2051 (N_2051,N_1943,N_1979);
nand U2052 (N_2052,N_1980,N_1990);
nand U2053 (N_2053,N_1901,N_1959);
and U2054 (N_2054,N_1995,N_1991);
nor U2055 (N_2055,N_1939,N_1977);
nor U2056 (N_2056,N_1959,N_1939);
nand U2057 (N_2057,N_1943,N_1973);
xor U2058 (N_2058,N_1956,N_1909);
or U2059 (N_2059,N_1989,N_1935);
and U2060 (N_2060,N_1902,N_1936);
and U2061 (N_2061,N_1955,N_1917);
or U2062 (N_2062,N_1934,N_1986);
or U2063 (N_2063,N_1989,N_1927);
or U2064 (N_2064,N_1961,N_1997);
nand U2065 (N_2065,N_1920,N_1903);
and U2066 (N_2066,N_1967,N_1987);
or U2067 (N_2067,N_1958,N_1957);
or U2068 (N_2068,N_1971,N_1905);
nor U2069 (N_2069,N_1906,N_1932);
nand U2070 (N_2070,N_1931,N_1919);
nand U2071 (N_2071,N_1962,N_1988);
nor U2072 (N_2072,N_1924,N_1950);
or U2073 (N_2073,N_1992,N_1994);
nor U2074 (N_2074,N_1974,N_1937);
nand U2075 (N_2075,N_1969,N_1927);
nor U2076 (N_2076,N_1916,N_1946);
or U2077 (N_2077,N_1960,N_1918);
nand U2078 (N_2078,N_1950,N_1987);
or U2079 (N_2079,N_1922,N_1978);
xnor U2080 (N_2080,N_1963,N_1983);
nor U2081 (N_2081,N_1995,N_1929);
or U2082 (N_2082,N_1989,N_1971);
and U2083 (N_2083,N_1919,N_1918);
or U2084 (N_2084,N_1964,N_1994);
or U2085 (N_2085,N_1978,N_1904);
xnor U2086 (N_2086,N_1987,N_1979);
xor U2087 (N_2087,N_1970,N_1920);
nand U2088 (N_2088,N_1989,N_1918);
and U2089 (N_2089,N_1972,N_1959);
nand U2090 (N_2090,N_1948,N_1981);
and U2091 (N_2091,N_1902,N_1906);
xnor U2092 (N_2092,N_1943,N_1938);
nand U2093 (N_2093,N_1982,N_1916);
or U2094 (N_2094,N_1934,N_1944);
xnor U2095 (N_2095,N_1964,N_1904);
nor U2096 (N_2096,N_1969,N_1901);
and U2097 (N_2097,N_1980,N_1979);
nand U2098 (N_2098,N_1988,N_1934);
or U2099 (N_2099,N_1953,N_1963);
nor U2100 (N_2100,N_2056,N_2028);
nor U2101 (N_2101,N_2070,N_2096);
xor U2102 (N_2102,N_2054,N_2006);
or U2103 (N_2103,N_2052,N_2073);
xnor U2104 (N_2104,N_2010,N_2090);
xor U2105 (N_2105,N_2024,N_2067);
nor U2106 (N_2106,N_2057,N_2032);
or U2107 (N_2107,N_2017,N_2012);
or U2108 (N_2108,N_2077,N_2045);
nor U2109 (N_2109,N_2088,N_2040);
nand U2110 (N_2110,N_2036,N_2043);
and U2111 (N_2111,N_2029,N_2086);
or U2112 (N_2112,N_2015,N_2019);
xnor U2113 (N_2113,N_2031,N_2072);
or U2114 (N_2114,N_2030,N_2009);
nand U2115 (N_2115,N_2047,N_2074);
nand U2116 (N_2116,N_2081,N_2049);
nand U2117 (N_2117,N_2008,N_2071);
or U2118 (N_2118,N_2061,N_2039);
or U2119 (N_2119,N_2060,N_2000);
or U2120 (N_2120,N_2002,N_2014);
nor U2121 (N_2121,N_2016,N_2011);
xnor U2122 (N_2122,N_2064,N_2003);
and U2123 (N_2123,N_2093,N_2075);
nor U2124 (N_2124,N_2050,N_2041);
or U2125 (N_2125,N_2053,N_2058);
and U2126 (N_2126,N_2084,N_2094);
nand U2127 (N_2127,N_2042,N_2001);
nor U2128 (N_2128,N_2020,N_2007);
nor U2129 (N_2129,N_2092,N_2097);
xor U2130 (N_2130,N_2098,N_2062);
nor U2131 (N_2131,N_2091,N_2026);
and U2132 (N_2132,N_2055,N_2018);
nor U2133 (N_2133,N_2025,N_2004);
nand U2134 (N_2134,N_2051,N_2065);
xor U2135 (N_2135,N_2037,N_2044);
nand U2136 (N_2136,N_2059,N_2087);
xnor U2137 (N_2137,N_2013,N_2080);
xor U2138 (N_2138,N_2022,N_2089);
and U2139 (N_2139,N_2033,N_2034);
nor U2140 (N_2140,N_2035,N_2076);
nand U2141 (N_2141,N_2046,N_2063);
xnor U2142 (N_2142,N_2068,N_2066);
xnor U2143 (N_2143,N_2099,N_2082);
nor U2144 (N_2144,N_2023,N_2048);
or U2145 (N_2145,N_2095,N_2021);
nand U2146 (N_2146,N_2079,N_2027);
nand U2147 (N_2147,N_2069,N_2005);
nand U2148 (N_2148,N_2078,N_2038);
nor U2149 (N_2149,N_2083,N_2085);
or U2150 (N_2150,N_2001,N_2084);
or U2151 (N_2151,N_2079,N_2041);
nor U2152 (N_2152,N_2051,N_2054);
nor U2153 (N_2153,N_2031,N_2073);
nand U2154 (N_2154,N_2007,N_2055);
xor U2155 (N_2155,N_2011,N_2084);
or U2156 (N_2156,N_2037,N_2059);
nand U2157 (N_2157,N_2008,N_2056);
nand U2158 (N_2158,N_2007,N_2004);
xor U2159 (N_2159,N_2026,N_2020);
or U2160 (N_2160,N_2064,N_2052);
and U2161 (N_2161,N_2028,N_2062);
xor U2162 (N_2162,N_2075,N_2053);
nand U2163 (N_2163,N_2010,N_2007);
nand U2164 (N_2164,N_2025,N_2046);
and U2165 (N_2165,N_2089,N_2078);
nand U2166 (N_2166,N_2061,N_2013);
or U2167 (N_2167,N_2057,N_2016);
or U2168 (N_2168,N_2055,N_2056);
nor U2169 (N_2169,N_2061,N_2089);
nor U2170 (N_2170,N_2090,N_2064);
nand U2171 (N_2171,N_2085,N_2025);
or U2172 (N_2172,N_2002,N_2088);
and U2173 (N_2173,N_2036,N_2011);
nand U2174 (N_2174,N_2071,N_2095);
nor U2175 (N_2175,N_2079,N_2047);
or U2176 (N_2176,N_2085,N_2016);
nor U2177 (N_2177,N_2078,N_2075);
nor U2178 (N_2178,N_2027,N_2018);
nor U2179 (N_2179,N_2087,N_2019);
or U2180 (N_2180,N_2067,N_2009);
or U2181 (N_2181,N_2002,N_2048);
and U2182 (N_2182,N_2008,N_2064);
or U2183 (N_2183,N_2078,N_2027);
xor U2184 (N_2184,N_2060,N_2073);
nor U2185 (N_2185,N_2064,N_2077);
nor U2186 (N_2186,N_2027,N_2082);
nor U2187 (N_2187,N_2058,N_2080);
or U2188 (N_2188,N_2083,N_2084);
xnor U2189 (N_2189,N_2021,N_2084);
nand U2190 (N_2190,N_2011,N_2037);
and U2191 (N_2191,N_2072,N_2087);
and U2192 (N_2192,N_2007,N_2075);
and U2193 (N_2193,N_2026,N_2068);
and U2194 (N_2194,N_2024,N_2088);
nor U2195 (N_2195,N_2006,N_2012);
xnor U2196 (N_2196,N_2028,N_2047);
nor U2197 (N_2197,N_2029,N_2087);
nand U2198 (N_2198,N_2051,N_2090);
nor U2199 (N_2199,N_2041,N_2004);
and U2200 (N_2200,N_2175,N_2117);
or U2201 (N_2201,N_2186,N_2101);
nor U2202 (N_2202,N_2141,N_2157);
or U2203 (N_2203,N_2178,N_2124);
or U2204 (N_2204,N_2112,N_2159);
or U2205 (N_2205,N_2174,N_2160);
and U2206 (N_2206,N_2187,N_2193);
nor U2207 (N_2207,N_2171,N_2122);
or U2208 (N_2208,N_2153,N_2177);
xnor U2209 (N_2209,N_2138,N_2179);
nand U2210 (N_2210,N_2111,N_2142);
and U2211 (N_2211,N_2170,N_2162);
nor U2212 (N_2212,N_2182,N_2125);
nand U2213 (N_2213,N_2189,N_2133);
nand U2214 (N_2214,N_2150,N_2169);
nor U2215 (N_2215,N_2176,N_2144);
and U2216 (N_2216,N_2195,N_2132);
nand U2217 (N_2217,N_2184,N_2198);
nor U2218 (N_2218,N_2135,N_2103);
nand U2219 (N_2219,N_2143,N_2163);
xnor U2220 (N_2220,N_2105,N_2197);
xor U2221 (N_2221,N_2155,N_2167);
xnor U2222 (N_2222,N_2131,N_2139);
nand U2223 (N_2223,N_2100,N_2108);
nor U2224 (N_2224,N_2196,N_2119);
and U2225 (N_2225,N_2129,N_2154);
and U2226 (N_2226,N_2115,N_2116);
nand U2227 (N_2227,N_2147,N_2158);
and U2228 (N_2228,N_2165,N_2191);
and U2229 (N_2229,N_2128,N_2130);
xnor U2230 (N_2230,N_2152,N_2109);
nor U2231 (N_2231,N_2145,N_2199);
nand U2232 (N_2232,N_2149,N_2118);
and U2233 (N_2233,N_2123,N_2161);
nor U2234 (N_2234,N_2120,N_2194);
nor U2235 (N_2235,N_2136,N_2121);
and U2236 (N_2236,N_2140,N_2173);
nand U2237 (N_2237,N_2192,N_2134);
nor U2238 (N_2238,N_2172,N_2168);
and U2239 (N_2239,N_2126,N_2183);
and U2240 (N_2240,N_2190,N_2146);
or U2241 (N_2241,N_2137,N_2127);
or U2242 (N_2242,N_2180,N_2188);
nand U2243 (N_2243,N_2181,N_2151);
nor U2244 (N_2244,N_2102,N_2106);
nor U2245 (N_2245,N_2148,N_2164);
and U2246 (N_2246,N_2104,N_2166);
nand U2247 (N_2247,N_2107,N_2110);
nand U2248 (N_2248,N_2114,N_2185);
and U2249 (N_2249,N_2156,N_2113);
nand U2250 (N_2250,N_2175,N_2116);
nand U2251 (N_2251,N_2103,N_2138);
nor U2252 (N_2252,N_2127,N_2117);
nor U2253 (N_2253,N_2191,N_2147);
nor U2254 (N_2254,N_2138,N_2176);
xor U2255 (N_2255,N_2165,N_2104);
or U2256 (N_2256,N_2123,N_2178);
nor U2257 (N_2257,N_2104,N_2105);
or U2258 (N_2258,N_2114,N_2110);
nor U2259 (N_2259,N_2139,N_2192);
and U2260 (N_2260,N_2140,N_2141);
or U2261 (N_2261,N_2124,N_2188);
or U2262 (N_2262,N_2115,N_2179);
xnor U2263 (N_2263,N_2151,N_2142);
xor U2264 (N_2264,N_2123,N_2141);
or U2265 (N_2265,N_2177,N_2172);
or U2266 (N_2266,N_2151,N_2165);
or U2267 (N_2267,N_2186,N_2181);
nor U2268 (N_2268,N_2188,N_2161);
and U2269 (N_2269,N_2108,N_2143);
nand U2270 (N_2270,N_2101,N_2174);
nor U2271 (N_2271,N_2150,N_2102);
nor U2272 (N_2272,N_2105,N_2152);
nand U2273 (N_2273,N_2114,N_2121);
nand U2274 (N_2274,N_2136,N_2124);
xor U2275 (N_2275,N_2155,N_2182);
and U2276 (N_2276,N_2128,N_2185);
or U2277 (N_2277,N_2104,N_2187);
or U2278 (N_2278,N_2128,N_2192);
nand U2279 (N_2279,N_2141,N_2180);
nor U2280 (N_2280,N_2125,N_2146);
or U2281 (N_2281,N_2181,N_2146);
nor U2282 (N_2282,N_2163,N_2190);
and U2283 (N_2283,N_2158,N_2134);
xor U2284 (N_2284,N_2197,N_2186);
nand U2285 (N_2285,N_2124,N_2153);
nand U2286 (N_2286,N_2129,N_2100);
nor U2287 (N_2287,N_2157,N_2111);
or U2288 (N_2288,N_2161,N_2139);
or U2289 (N_2289,N_2130,N_2196);
and U2290 (N_2290,N_2155,N_2188);
nand U2291 (N_2291,N_2116,N_2169);
and U2292 (N_2292,N_2135,N_2131);
xor U2293 (N_2293,N_2187,N_2182);
or U2294 (N_2294,N_2168,N_2117);
nand U2295 (N_2295,N_2128,N_2166);
or U2296 (N_2296,N_2101,N_2128);
nand U2297 (N_2297,N_2121,N_2115);
or U2298 (N_2298,N_2117,N_2149);
nand U2299 (N_2299,N_2142,N_2101);
xor U2300 (N_2300,N_2280,N_2226);
or U2301 (N_2301,N_2261,N_2231);
nand U2302 (N_2302,N_2225,N_2237);
nand U2303 (N_2303,N_2282,N_2294);
nand U2304 (N_2304,N_2287,N_2299);
and U2305 (N_2305,N_2286,N_2218);
xor U2306 (N_2306,N_2281,N_2283);
and U2307 (N_2307,N_2242,N_2267);
or U2308 (N_2308,N_2247,N_2271);
and U2309 (N_2309,N_2222,N_2268);
nor U2310 (N_2310,N_2213,N_2252);
xor U2311 (N_2311,N_2227,N_2262);
and U2312 (N_2312,N_2243,N_2290);
nand U2313 (N_2313,N_2248,N_2206);
or U2314 (N_2314,N_2263,N_2256);
or U2315 (N_2315,N_2273,N_2291);
nor U2316 (N_2316,N_2288,N_2224);
nor U2317 (N_2317,N_2204,N_2238);
xor U2318 (N_2318,N_2296,N_2279);
nor U2319 (N_2319,N_2239,N_2245);
and U2320 (N_2320,N_2285,N_2244);
nand U2321 (N_2321,N_2295,N_2232);
or U2322 (N_2322,N_2275,N_2253);
nor U2323 (N_2323,N_2235,N_2258);
or U2324 (N_2324,N_2223,N_2249);
nor U2325 (N_2325,N_2208,N_2212);
xnor U2326 (N_2326,N_2229,N_2298);
xnor U2327 (N_2327,N_2221,N_2257);
or U2328 (N_2328,N_2254,N_2210);
nand U2329 (N_2329,N_2207,N_2217);
and U2330 (N_2330,N_2277,N_2250);
nor U2331 (N_2331,N_2284,N_2293);
nor U2332 (N_2332,N_2297,N_2203);
or U2333 (N_2333,N_2202,N_2240);
nand U2334 (N_2334,N_2266,N_2236);
and U2335 (N_2335,N_2289,N_2234);
or U2336 (N_2336,N_2201,N_2205);
nor U2337 (N_2337,N_2264,N_2260);
and U2338 (N_2338,N_2219,N_2270);
xnor U2339 (N_2339,N_2209,N_2276);
nor U2340 (N_2340,N_2216,N_2214);
and U2341 (N_2341,N_2233,N_2292);
and U2342 (N_2342,N_2228,N_2278);
or U2343 (N_2343,N_2265,N_2215);
xnor U2344 (N_2344,N_2230,N_2259);
nor U2345 (N_2345,N_2246,N_2211);
xor U2346 (N_2346,N_2220,N_2272);
and U2347 (N_2347,N_2255,N_2200);
nand U2348 (N_2348,N_2251,N_2274);
and U2349 (N_2349,N_2269,N_2241);
or U2350 (N_2350,N_2286,N_2209);
nor U2351 (N_2351,N_2273,N_2246);
xnor U2352 (N_2352,N_2280,N_2218);
or U2353 (N_2353,N_2209,N_2293);
or U2354 (N_2354,N_2235,N_2275);
xor U2355 (N_2355,N_2256,N_2241);
nand U2356 (N_2356,N_2211,N_2251);
and U2357 (N_2357,N_2231,N_2292);
and U2358 (N_2358,N_2212,N_2283);
and U2359 (N_2359,N_2210,N_2237);
xnor U2360 (N_2360,N_2221,N_2237);
and U2361 (N_2361,N_2259,N_2279);
and U2362 (N_2362,N_2209,N_2239);
nand U2363 (N_2363,N_2226,N_2272);
nor U2364 (N_2364,N_2258,N_2234);
or U2365 (N_2365,N_2262,N_2282);
and U2366 (N_2366,N_2225,N_2299);
xor U2367 (N_2367,N_2274,N_2237);
or U2368 (N_2368,N_2290,N_2257);
xor U2369 (N_2369,N_2252,N_2242);
nor U2370 (N_2370,N_2226,N_2227);
nand U2371 (N_2371,N_2220,N_2285);
xor U2372 (N_2372,N_2239,N_2284);
xor U2373 (N_2373,N_2294,N_2298);
xor U2374 (N_2374,N_2259,N_2241);
or U2375 (N_2375,N_2245,N_2297);
or U2376 (N_2376,N_2264,N_2212);
or U2377 (N_2377,N_2291,N_2245);
and U2378 (N_2378,N_2217,N_2296);
nor U2379 (N_2379,N_2264,N_2219);
and U2380 (N_2380,N_2259,N_2211);
or U2381 (N_2381,N_2248,N_2241);
xnor U2382 (N_2382,N_2212,N_2265);
nand U2383 (N_2383,N_2221,N_2290);
nor U2384 (N_2384,N_2244,N_2251);
and U2385 (N_2385,N_2283,N_2221);
or U2386 (N_2386,N_2220,N_2293);
or U2387 (N_2387,N_2267,N_2227);
xnor U2388 (N_2388,N_2244,N_2238);
xor U2389 (N_2389,N_2291,N_2265);
nor U2390 (N_2390,N_2280,N_2291);
nor U2391 (N_2391,N_2249,N_2207);
or U2392 (N_2392,N_2217,N_2288);
nand U2393 (N_2393,N_2290,N_2200);
nor U2394 (N_2394,N_2246,N_2279);
and U2395 (N_2395,N_2211,N_2236);
xnor U2396 (N_2396,N_2200,N_2249);
xor U2397 (N_2397,N_2229,N_2240);
nor U2398 (N_2398,N_2269,N_2282);
nor U2399 (N_2399,N_2266,N_2220);
nor U2400 (N_2400,N_2324,N_2304);
nand U2401 (N_2401,N_2322,N_2364);
nor U2402 (N_2402,N_2384,N_2332);
nor U2403 (N_2403,N_2378,N_2360);
xor U2404 (N_2404,N_2350,N_2312);
nand U2405 (N_2405,N_2338,N_2363);
nor U2406 (N_2406,N_2357,N_2301);
or U2407 (N_2407,N_2300,N_2348);
or U2408 (N_2408,N_2305,N_2316);
and U2409 (N_2409,N_2377,N_2394);
or U2410 (N_2410,N_2358,N_2388);
and U2411 (N_2411,N_2331,N_2379);
nor U2412 (N_2412,N_2370,N_2335);
nor U2413 (N_2413,N_2376,N_2337);
or U2414 (N_2414,N_2302,N_2343);
nand U2415 (N_2415,N_2375,N_2395);
nand U2416 (N_2416,N_2303,N_2380);
nand U2417 (N_2417,N_2385,N_2361);
or U2418 (N_2418,N_2330,N_2310);
nand U2419 (N_2419,N_2342,N_2349);
or U2420 (N_2420,N_2355,N_2398);
nor U2421 (N_2421,N_2315,N_2387);
nand U2422 (N_2422,N_2340,N_2399);
xor U2423 (N_2423,N_2346,N_2323);
xor U2424 (N_2424,N_2329,N_2369);
or U2425 (N_2425,N_2389,N_2366);
nor U2426 (N_2426,N_2371,N_2333);
xnor U2427 (N_2427,N_2372,N_2374);
xor U2428 (N_2428,N_2311,N_2344);
nand U2429 (N_2429,N_2336,N_2327);
nand U2430 (N_2430,N_2353,N_2318);
or U2431 (N_2431,N_2391,N_2306);
nor U2432 (N_2432,N_2362,N_2314);
nand U2433 (N_2433,N_2339,N_2368);
or U2434 (N_2434,N_2397,N_2334);
nand U2435 (N_2435,N_2341,N_2390);
nand U2436 (N_2436,N_2309,N_2392);
or U2437 (N_2437,N_2328,N_2354);
nand U2438 (N_2438,N_2308,N_2383);
or U2439 (N_2439,N_2365,N_2381);
nor U2440 (N_2440,N_2313,N_2382);
or U2441 (N_2441,N_2345,N_2356);
or U2442 (N_2442,N_2326,N_2319);
xor U2443 (N_2443,N_2317,N_2359);
xnor U2444 (N_2444,N_2325,N_2396);
xor U2445 (N_2445,N_2393,N_2351);
and U2446 (N_2446,N_2386,N_2347);
and U2447 (N_2447,N_2352,N_2320);
xor U2448 (N_2448,N_2321,N_2373);
xor U2449 (N_2449,N_2307,N_2367);
nand U2450 (N_2450,N_2377,N_2348);
nand U2451 (N_2451,N_2309,N_2390);
nand U2452 (N_2452,N_2349,N_2352);
xor U2453 (N_2453,N_2378,N_2325);
nor U2454 (N_2454,N_2378,N_2328);
and U2455 (N_2455,N_2312,N_2399);
or U2456 (N_2456,N_2357,N_2327);
nand U2457 (N_2457,N_2386,N_2394);
or U2458 (N_2458,N_2399,N_2308);
nand U2459 (N_2459,N_2303,N_2383);
xnor U2460 (N_2460,N_2362,N_2391);
xnor U2461 (N_2461,N_2329,N_2324);
xnor U2462 (N_2462,N_2314,N_2395);
xnor U2463 (N_2463,N_2375,N_2310);
or U2464 (N_2464,N_2337,N_2300);
xor U2465 (N_2465,N_2322,N_2382);
or U2466 (N_2466,N_2360,N_2372);
or U2467 (N_2467,N_2394,N_2390);
nand U2468 (N_2468,N_2350,N_2363);
xnor U2469 (N_2469,N_2347,N_2321);
or U2470 (N_2470,N_2379,N_2358);
and U2471 (N_2471,N_2306,N_2355);
xor U2472 (N_2472,N_2388,N_2342);
nor U2473 (N_2473,N_2325,N_2398);
xnor U2474 (N_2474,N_2311,N_2369);
nor U2475 (N_2475,N_2306,N_2329);
nand U2476 (N_2476,N_2361,N_2380);
nand U2477 (N_2477,N_2392,N_2383);
nor U2478 (N_2478,N_2374,N_2389);
and U2479 (N_2479,N_2343,N_2397);
xnor U2480 (N_2480,N_2385,N_2306);
nand U2481 (N_2481,N_2346,N_2397);
xnor U2482 (N_2482,N_2388,N_2337);
xnor U2483 (N_2483,N_2315,N_2391);
or U2484 (N_2484,N_2320,N_2312);
xor U2485 (N_2485,N_2380,N_2345);
and U2486 (N_2486,N_2377,N_2374);
and U2487 (N_2487,N_2348,N_2302);
xnor U2488 (N_2488,N_2380,N_2326);
and U2489 (N_2489,N_2365,N_2331);
nand U2490 (N_2490,N_2334,N_2381);
nand U2491 (N_2491,N_2303,N_2353);
nor U2492 (N_2492,N_2397,N_2395);
xnor U2493 (N_2493,N_2367,N_2383);
or U2494 (N_2494,N_2320,N_2341);
xnor U2495 (N_2495,N_2369,N_2387);
and U2496 (N_2496,N_2392,N_2385);
nand U2497 (N_2497,N_2321,N_2306);
nand U2498 (N_2498,N_2313,N_2358);
nor U2499 (N_2499,N_2307,N_2315);
nand U2500 (N_2500,N_2446,N_2456);
nor U2501 (N_2501,N_2408,N_2473);
nor U2502 (N_2502,N_2487,N_2438);
nand U2503 (N_2503,N_2450,N_2442);
nand U2504 (N_2504,N_2451,N_2428);
xnor U2505 (N_2505,N_2415,N_2478);
nor U2506 (N_2506,N_2469,N_2427);
nor U2507 (N_2507,N_2494,N_2412);
and U2508 (N_2508,N_2437,N_2470);
and U2509 (N_2509,N_2432,N_2493);
nand U2510 (N_2510,N_2477,N_2460);
nand U2511 (N_2511,N_2439,N_2454);
xor U2512 (N_2512,N_2490,N_2472);
or U2513 (N_2513,N_2453,N_2463);
and U2514 (N_2514,N_2422,N_2409);
xnor U2515 (N_2515,N_2475,N_2496);
and U2516 (N_2516,N_2457,N_2418);
nand U2517 (N_2517,N_2402,N_2459);
and U2518 (N_2518,N_2420,N_2462);
and U2519 (N_2519,N_2474,N_2497);
nand U2520 (N_2520,N_2486,N_2476);
and U2521 (N_2521,N_2464,N_2467);
or U2522 (N_2522,N_2492,N_2421);
and U2523 (N_2523,N_2488,N_2465);
nand U2524 (N_2524,N_2424,N_2405);
and U2525 (N_2525,N_2491,N_2483);
nor U2526 (N_2526,N_2434,N_2406);
nor U2527 (N_2527,N_2435,N_2426);
nor U2528 (N_2528,N_2468,N_2461);
or U2529 (N_2529,N_2404,N_2480);
or U2530 (N_2530,N_2449,N_2433);
nor U2531 (N_2531,N_2429,N_2455);
nand U2532 (N_2532,N_2400,N_2413);
nand U2533 (N_2533,N_2410,N_2458);
or U2534 (N_2534,N_2414,N_2443);
and U2535 (N_2535,N_2445,N_2489);
or U2536 (N_2536,N_2481,N_2452);
or U2537 (N_2537,N_2495,N_2407);
nand U2538 (N_2538,N_2485,N_2417);
xor U2539 (N_2539,N_2440,N_2479);
xor U2540 (N_2540,N_2482,N_2447);
nor U2541 (N_2541,N_2441,N_2444);
xor U2542 (N_2542,N_2448,N_2471);
and U2543 (N_2543,N_2430,N_2416);
and U2544 (N_2544,N_2425,N_2419);
nand U2545 (N_2545,N_2499,N_2403);
and U2546 (N_2546,N_2401,N_2436);
and U2547 (N_2547,N_2498,N_2466);
and U2548 (N_2548,N_2423,N_2484);
or U2549 (N_2549,N_2431,N_2411);
nand U2550 (N_2550,N_2435,N_2449);
nand U2551 (N_2551,N_2419,N_2421);
nor U2552 (N_2552,N_2480,N_2407);
xnor U2553 (N_2553,N_2468,N_2479);
nor U2554 (N_2554,N_2484,N_2480);
nor U2555 (N_2555,N_2435,N_2488);
nand U2556 (N_2556,N_2485,N_2406);
or U2557 (N_2557,N_2402,N_2479);
nor U2558 (N_2558,N_2478,N_2419);
nor U2559 (N_2559,N_2413,N_2476);
xnor U2560 (N_2560,N_2445,N_2433);
nor U2561 (N_2561,N_2499,N_2476);
or U2562 (N_2562,N_2448,N_2460);
or U2563 (N_2563,N_2479,N_2458);
or U2564 (N_2564,N_2437,N_2469);
and U2565 (N_2565,N_2408,N_2490);
nand U2566 (N_2566,N_2409,N_2485);
xnor U2567 (N_2567,N_2416,N_2424);
xnor U2568 (N_2568,N_2463,N_2494);
and U2569 (N_2569,N_2478,N_2494);
or U2570 (N_2570,N_2450,N_2406);
or U2571 (N_2571,N_2426,N_2458);
xnor U2572 (N_2572,N_2478,N_2433);
or U2573 (N_2573,N_2415,N_2472);
xor U2574 (N_2574,N_2400,N_2489);
xor U2575 (N_2575,N_2474,N_2410);
xnor U2576 (N_2576,N_2432,N_2472);
nor U2577 (N_2577,N_2483,N_2456);
nor U2578 (N_2578,N_2474,N_2496);
and U2579 (N_2579,N_2485,N_2418);
nand U2580 (N_2580,N_2482,N_2498);
or U2581 (N_2581,N_2493,N_2408);
xor U2582 (N_2582,N_2436,N_2461);
and U2583 (N_2583,N_2414,N_2485);
xnor U2584 (N_2584,N_2441,N_2438);
and U2585 (N_2585,N_2467,N_2496);
nand U2586 (N_2586,N_2485,N_2486);
xor U2587 (N_2587,N_2461,N_2470);
nand U2588 (N_2588,N_2423,N_2415);
nor U2589 (N_2589,N_2439,N_2465);
and U2590 (N_2590,N_2464,N_2413);
xnor U2591 (N_2591,N_2451,N_2456);
or U2592 (N_2592,N_2424,N_2488);
nor U2593 (N_2593,N_2490,N_2420);
or U2594 (N_2594,N_2472,N_2494);
or U2595 (N_2595,N_2467,N_2420);
nand U2596 (N_2596,N_2450,N_2433);
and U2597 (N_2597,N_2490,N_2471);
or U2598 (N_2598,N_2414,N_2452);
or U2599 (N_2599,N_2435,N_2487);
and U2600 (N_2600,N_2573,N_2543);
or U2601 (N_2601,N_2545,N_2597);
and U2602 (N_2602,N_2539,N_2508);
or U2603 (N_2603,N_2533,N_2546);
nor U2604 (N_2604,N_2564,N_2561);
nand U2605 (N_2605,N_2535,N_2563);
nand U2606 (N_2606,N_2532,N_2522);
and U2607 (N_2607,N_2588,N_2550);
and U2608 (N_2608,N_2523,N_2529);
nand U2609 (N_2609,N_2575,N_2500);
xnor U2610 (N_2610,N_2507,N_2574);
and U2611 (N_2611,N_2526,N_2520);
nor U2612 (N_2612,N_2599,N_2540);
nand U2613 (N_2613,N_2547,N_2583);
xnor U2614 (N_2614,N_2586,N_2571);
or U2615 (N_2615,N_2514,N_2534);
nand U2616 (N_2616,N_2506,N_2578);
nor U2617 (N_2617,N_2565,N_2556);
nor U2618 (N_2618,N_2515,N_2509);
nand U2619 (N_2619,N_2552,N_2592);
or U2620 (N_2620,N_2555,N_2585);
nand U2621 (N_2621,N_2551,N_2582);
and U2622 (N_2622,N_2549,N_2570);
xor U2623 (N_2623,N_2544,N_2593);
nand U2624 (N_2624,N_2572,N_2530);
nor U2625 (N_2625,N_2519,N_2568);
xor U2626 (N_2626,N_2538,N_2516);
or U2627 (N_2627,N_2581,N_2521);
nand U2628 (N_2628,N_2566,N_2542);
nand U2629 (N_2629,N_2580,N_2576);
or U2630 (N_2630,N_2503,N_2584);
xor U2631 (N_2631,N_2595,N_2502);
or U2632 (N_2632,N_2510,N_2587);
xnor U2633 (N_2633,N_2589,N_2569);
nand U2634 (N_2634,N_2505,N_2537);
nor U2635 (N_2635,N_2591,N_2531);
and U2636 (N_2636,N_2596,N_2559);
xor U2637 (N_2637,N_2554,N_2536);
nand U2638 (N_2638,N_2553,N_2598);
xor U2639 (N_2639,N_2513,N_2558);
or U2640 (N_2640,N_2557,N_2562);
and U2641 (N_2641,N_2560,N_2504);
and U2642 (N_2642,N_2528,N_2524);
and U2643 (N_2643,N_2541,N_2512);
nand U2644 (N_2644,N_2518,N_2567);
nand U2645 (N_2645,N_2511,N_2579);
nor U2646 (N_2646,N_2577,N_2590);
nor U2647 (N_2647,N_2548,N_2517);
nand U2648 (N_2648,N_2594,N_2527);
nor U2649 (N_2649,N_2501,N_2525);
nor U2650 (N_2650,N_2582,N_2562);
nand U2651 (N_2651,N_2576,N_2589);
xor U2652 (N_2652,N_2521,N_2533);
and U2653 (N_2653,N_2555,N_2570);
xnor U2654 (N_2654,N_2528,N_2521);
xor U2655 (N_2655,N_2517,N_2554);
nand U2656 (N_2656,N_2501,N_2510);
and U2657 (N_2657,N_2555,N_2518);
or U2658 (N_2658,N_2599,N_2516);
and U2659 (N_2659,N_2512,N_2588);
nor U2660 (N_2660,N_2562,N_2515);
nor U2661 (N_2661,N_2528,N_2511);
nor U2662 (N_2662,N_2512,N_2536);
and U2663 (N_2663,N_2550,N_2555);
and U2664 (N_2664,N_2504,N_2501);
nand U2665 (N_2665,N_2561,N_2529);
xor U2666 (N_2666,N_2530,N_2594);
xor U2667 (N_2667,N_2590,N_2566);
xor U2668 (N_2668,N_2561,N_2587);
or U2669 (N_2669,N_2568,N_2509);
and U2670 (N_2670,N_2508,N_2530);
nand U2671 (N_2671,N_2554,N_2588);
or U2672 (N_2672,N_2546,N_2578);
nor U2673 (N_2673,N_2540,N_2500);
and U2674 (N_2674,N_2527,N_2511);
nand U2675 (N_2675,N_2502,N_2561);
or U2676 (N_2676,N_2554,N_2506);
or U2677 (N_2677,N_2509,N_2532);
and U2678 (N_2678,N_2505,N_2583);
and U2679 (N_2679,N_2528,N_2512);
or U2680 (N_2680,N_2508,N_2549);
nor U2681 (N_2681,N_2590,N_2521);
or U2682 (N_2682,N_2510,N_2583);
nor U2683 (N_2683,N_2546,N_2540);
and U2684 (N_2684,N_2566,N_2558);
or U2685 (N_2685,N_2521,N_2540);
nand U2686 (N_2686,N_2524,N_2569);
nand U2687 (N_2687,N_2530,N_2548);
and U2688 (N_2688,N_2584,N_2556);
xnor U2689 (N_2689,N_2545,N_2522);
and U2690 (N_2690,N_2527,N_2588);
xnor U2691 (N_2691,N_2523,N_2557);
nand U2692 (N_2692,N_2552,N_2511);
xor U2693 (N_2693,N_2552,N_2564);
nand U2694 (N_2694,N_2565,N_2594);
and U2695 (N_2695,N_2518,N_2549);
or U2696 (N_2696,N_2573,N_2539);
and U2697 (N_2697,N_2593,N_2585);
nand U2698 (N_2698,N_2563,N_2571);
or U2699 (N_2699,N_2563,N_2577);
or U2700 (N_2700,N_2630,N_2610);
and U2701 (N_2701,N_2628,N_2688);
nor U2702 (N_2702,N_2643,N_2662);
xnor U2703 (N_2703,N_2616,N_2670);
xor U2704 (N_2704,N_2698,N_2673);
nand U2705 (N_2705,N_2693,N_2666);
nor U2706 (N_2706,N_2667,N_2695);
and U2707 (N_2707,N_2655,N_2625);
xor U2708 (N_2708,N_2638,N_2682);
and U2709 (N_2709,N_2674,N_2653);
and U2710 (N_2710,N_2680,N_2632);
nand U2711 (N_2711,N_2622,N_2637);
nand U2712 (N_2712,N_2664,N_2627);
nand U2713 (N_2713,N_2671,N_2651);
nor U2714 (N_2714,N_2629,N_2665);
nand U2715 (N_2715,N_2634,N_2642);
xnor U2716 (N_2716,N_2648,N_2645);
or U2717 (N_2717,N_2601,N_2613);
xnor U2718 (N_2718,N_2657,N_2621);
nand U2719 (N_2719,N_2668,N_2681);
xor U2720 (N_2720,N_2606,N_2672);
or U2721 (N_2721,N_2635,N_2611);
nand U2722 (N_2722,N_2663,N_2615);
or U2723 (N_2723,N_2603,N_2640);
and U2724 (N_2724,N_2609,N_2683);
xnor U2725 (N_2725,N_2626,N_2639);
nor U2726 (N_2726,N_2600,N_2676);
and U2727 (N_2727,N_2602,N_2661);
nor U2728 (N_2728,N_2654,N_2608);
nor U2729 (N_2729,N_2677,N_2612);
nand U2730 (N_2730,N_2624,N_2694);
and U2731 (N_2731,N_2660,N_2650);
nand U2732 (N_2732,N_2618,N_2689);
nand U2733 (N_2733,N_2614,N_2690);
nand U2734 (N_2734,N_2652,N_2696);
or U2735 (N_2735,N_2649,N_2636);
or U2736 (N_2736,N_2678,N_2669);
nand U2737 (N_2737,N_2684,N_2675);
nor U2738 (N_2738,N_2631,N_2697);
xor U2739 (N_2739,N_2686,N_2658);
xor U2740 (N_2740,N_2641,N_2607);
and U2741 (N_2741,N_2692,N_2604);
nor U2742 (N_2742,N_2679,N_2620);
nand U2743 (N_2743,N_2691,N_2699);
or U2744 (N_2744,N_2647,N_2656);
xor U2745 (N_2745,N_2617,N_2619);
and U2746 (N_2746,N_2659,N_2687);
nand U2747 (N_2747,N_2633,N_2644);
or U2748 (N_2748,N_2646,N_2623);
nand U2749 (N_2749,N_2605,N_2685);
xor U2750 (N_2750,N_2635,N_2644);
or U2751 (N_2751,N_2689,N_2697);
xor U2752 (N_2752,N_2671,N_2656);
and U2753 (N_2753,N_2629,N_2617);
or U2754 (N_2754,N_2697,N_2668);
or U2755 (N_2755,N_2600,N_2665);
nor U2756 (N_2756,N_2697,N_2628);
or U2757 (N_2757,N_2608,N_2638);
nand U2758 (N_2758,N_2685,N_2600);
and U2759 (N_2759,N_2600,N_2666);
nand U2760 (N_2760,N_2692,N_2631);
nand U2761 (N_2761,N_2691,N_2667);
xnor U2762 (N_2762,N_2605,N_2696);
and U2763 (N_2763,N_2691,N_2638);
or U2764 (N_2764,N_2657,N_2671);
nand U2765 (N_2765,N_2642,N_2606);
nor U2766 (N_2766,N_2681,N_2652);
nor U2767 (N_2767,N_2600,N_2684);
nand U2768 (N_2768,N_2623,N_2687);
nor U2769 (N_2769,N_2646,N_2689);
and U2770 (N_2770,N_2686,N_2691);
and U2771 (N_2771,N_2604,N_2615);
xnor U2772 (N_2772,N_2625,N_2672);
or U2773 (N_2773,N_2607,N_2600);
and U2774 (N_2774,N_2697,N_2600);
or U2775 (N_2775,N_2619,N_2624);
nand U2776 (N_2776,N_2667,N_2644);
and U2777 (N_2777,N_2673,N_2649);
and U2778 (N_2778,N_2647,N_2603);
and U2779 (N_2779,N_2633,N_2638);
or U2780 (N_2780,N_2615,N_2648);
nor U2781 (N_2781,N_2624,N_2631);
xnor U2782 (N_2782,N_2666,N_2673);
xnor U2783 (N_2783,N_2600,N_2627);
nand U2784 (N_2784,N_2690,N_2627);
xnor U2785 (N_2785,N_2656,N_2691);
nor U2786 (N_2786,N_2650,N_2661);
nor U2787 (N_2787,N_2627,N_2652);
xnor U2788 (N_2788,N_2647,N_2642);
xor U2789 (N_2789,N_2697,N_2614);
or U2790 (N_2790,N_2606,N_2614);
nor U2791 (N_2791,N_2697,N_2635);
xnor U2792 (N_2792,N_2693,N_2687);
xnor U2793 (N_2793,N_2629,N_2649);
or U2794 (N_2794,N_2638,N_2672);
and U2795 (N_2795,N_2630,N_2619);
xor U2796 (N_2796,N_2654,N_2694);
and U2797 (N_2797,N_2634,N_2668);
nor U2798 (N_2798,N_2686,N_2699);
and U2799 (N_2799,N_2600,N_2624);
nand U2800 (N_2800,N_2778,N_2701);
xor U2801 (N_2801,N_2709,N_2759);
or U2802 (N_2802,N_2768,N_2782);
and U2803 (N_2803,N_2748,N_2738);
nand U2804 (N_2804,N_2716,N_2733);
or U2805 (N_2805,N_2773,N_2711);
or U2806 (N_2806,N_2740,N_2749);
or U2807 (N_2807,N_2770,N_2702);
nor U2808 (N_2808,N_2783,N_2751);
or U2809 (N_2809,N_2721,N_2758);
or U2810 (N_2810,N_2752,N_2750);
and U2811 (N_2811,N_2786,N_2784);
nor U2812 (N_2812,N_2706,N_2717);
or U2813 (N_2813,N_2710,N_2776);
nand U2814 (N_2814,N_2728,N_2700);
or U2815 (N_2815,N_2798,N_2777);
xnor U2816 (N_2816,N_2739,N_2722);
nand U2817 (N_2817,N_2703,N_2771);
nand U2818 (N_2818,N_2742,N_2719);
nor U2819 (N_2819,N_2767,N_2724);
or U2820 (N_2820,N_2705,N_2743);
or U2821 (N_2821,N_2720,N_2741);
and U2822 (N_2822,N_2761,N_2760);
xor U2823 (N_2823,N_2779,N_2789);
nand U2824 (N_2824,N_2745,N_2723);
nand U2825 (N_2825,N_2726,N_2796);
or U2826 (N_2826,N_2762,N_2736);
xor U2827 (N_2827,N_2785,N_2708);
and U2828 (N_2828,N_2769,N_2788);
and U2829 (N_2829,N_2764,N_2714);
xnor U2830 (N_2830,N_2732,N_2730);
nor U2831 (N_2831,N_2731,N_2757);
or U2832 (N_2832,N_2765,N_2780);
and U2833 (N_2833,N_2737,N_2755);
nand U2834 (N_2834,N_2766,N_2747);
nor U2835 (N_2835,N_2754,N_2787);
xnor U2836 (N_2836,N_2797,N_2763);
nor U2837 (N_2837,N_2746,N_2729);
and U2838 (N_2838,N_2713,N_2735);
nor U2839 (N_2839,N_2727,N_2715);
nor U2840 (N_2840,N_2781,N_2753);
xor U2841 (N_2841,N_2718,N_2794);
or U2842 (N_2842,N_2799,N_2744);
xor U2843 (N_2843,N_2791,N_2775);
xor U2844 (N_2844,N_2734,N_2792);
and U2845 (N_2845,N_2793,N_2725);
nand U2846 (N_2846,N_2772,N_2774);
nand U2847 (N_2847,N_2790,N_2712);
nor U2848 (N_2848,N_2795,N_2756);
nor U2849 (N_2849,N_2704,N_2707);
nor U2850 (N_2850,N_2706,N_2781);
or U2851 (N_2851,N_2766,N_2774);
or U2852 (N_2852,N_2749,N_2788);
xnor U2853 (N_2853,N_2731,N_2711);
or U2854 (N_2854,N_2769,N_2756);
nor U2855 (N_2855,N_2742,N_2764);
or U2856 (N_2856,N_2763,N_2760);
nor U2857 (N_2857,N_2702,N_2747);
or U2858 (N_2858,N_2701,N_2716);
and U2859 (N_2859,N_2731,N_2726);
or U2860 (N_2860,N_2786,N_2773);
or U2861 (N_2861,N_2754,N_2755);
nand U2862 (N_2862,N_2720,N_2737);
and U2863 (N_2863,N_2713,N_2784);
nand U2864 (N_2864,N_2734,N_2710);
xor U2865 (N_2865,N_2712,N_2773);
nor U2866 (N_2866,N_2706,N_2734);
and U2867 (N_2867,N_2799,N_2775);
or U2868 (N_2868,N_2797,N_2781);
or U2869 (N_2869,N_2788,N_2716);
and U2870 (N_2870,N_2733,N_2721);
or U2871 (N_2871,N_2719,N_2792);
and U2872 (N_2872,N_2711,N_2782);
and U2873 (N_2873,N_2777,N_2734);
nor U2874 (N_2874,N_2786,N_2779);
xor U2875 (N_2875,N_2761,N_2794);
nand U2876 (N_2876,N_2797,N_2725);
nor U2877 (N_2877,N_2749,N_2704);
and U2878 (N_2878,N_2790,N_2768);
and U2879 (N_2879,N_2795,N_2753);
or U2880 (N_2880,N_2748,N_2783);
nor U2881 (N_2881,N_2724,N_2733);
xnor U2882 (N_2882,N_2749,N_2790);
nand U2883 (N_2883,N_2759,N_2732);
xor U2884 (N_2884,N_2724,N_2714);
nor U2885 (N_2885,N_2790,N_2727);
and U2886 (N_2886,N_2742,N_2753);
xnor U2887 (N_2887,N_2735,N_2721);
or U2888 (N_2888,N_2748,N_2751);
xor U2889 (N_2889,N_2701,N_2702);
and U2890 (N_2890,N_2756,N_2787);
xor U2891 (N_2891,N_2737,N_2733);
and U2892 (N_2892,N_2725,N_2775);
nor U2893 (N_2893,N_2746,N_2753);
nand U2894 (N_2894,N_2781,N_2769);
and U2895 (N_2895,N_2728,N_2720);
and U2896 (N_2896,N_2797,N_2743);
or U2897 (N_2897,N_2746,N_2719);
nand U2898 (N_2898,N_2786,N_2723);
nor U2899 (N_2899,N_2773,N_2716);
nand U2900 (N_2900,N_2861,N_2844);
and U2901 (N_2901,N_2865,N_2873);
nor U2902 (N_2902,N_2819,N_2802);
and U2903 (N_2903,N_2858,N_2875);
nor U2904 (N_2904,N_2808,N_2816);
nor U2905 (N_2905,N_2830,N_2837);
xor U2906 (N_2906,N_2892,N_2843);
xor U2907 (N_2907,N_2870,N_2871);
and U2908 (N_2908,N_2853,N_2867);
nor U2909 (N_2909,N_2863,N_2860);
xor U2910 (N_2910,N_2852,N_2874);
nand U2911 (N_2911,N_2803,N_2869);
nor U2912 (N_2912,N_2888,N_2818);
nor U2913 (N_2913,N_2847,N_2801);
nor U2914 (N_2914,N_2890,N_2856);
and U2915 (N_2915,N_2879,N_2887);
nand U2916 (N_2916,N_2895,N_2809);
xnor U2917 (N_2917,N_2850,N_2824);
xnor U2918 (N_2918,N_2845,N_2827);
and U2919 (N_2919,N_2831,N_2834);
and U2920 (N_2920,N_2848,N_2817);
nor U2921 (N_2921,N_2810,N_2804);
or U2922 (N_2922,N_2898,N_2807);
nand U2923 (N_2923,N_2812,N_2899);
nand U2924 (N_2924,N_2882,N_2893);
and U2925 (N_2925,N_2805,N_2823);
nor U2926 (N_2926,N_2866,N_2857);
nor U2927 (N_2927,N_2897,N_2881);
nand U2928 (N_2928,N_2806,N_2862);
and U2929 (N_2929,N_2822,N_2864);
nor U2930 (N_2930,N_2855,N_2883);
nand U2931 (N_2931,N_2885,N_2886);
and U2932 (N_2932,N_2896,N_2813);
and U2933 (N_2933,N_2841,N_2815);
and U2934 (N_2934,N_2839,N_2811);
nor U2935 (N_2935,N_2836,N_2854);
nor U2936 (N_2936,N_2820,N_2825);
nand U2937 (N_2937,N_2833,N_2878);
xor U2938 (N_2938,N_2868,N_2880);
and U2939 (N_2939,N_2849,N_2884);
nand U2940 (N_2940,N_2800,N_2877);
nor U2941 (N_2941,N_2832,N_2828);
or U2942 (N_2942,N_2876,N_2851);
and U2943 (N_2943,N_2814,N_2859);
and U2944 (N_2944,N_2835,N_2840);
or U2945 (N_2945,N_2891,N_2846);
and U2946 (N_2946,N_2838,N_2889);
xor U2947 (N_2947,N_2842,N_2821);
nor U2948 (N_2948,N_2826,N_2894);
nor U2949 (N_2949,N_2829,N_2872);
nor U2950 (N_2950,N_2835,N_2862);
xnor U2951 (N_2951,N_2873,N_2800);
or U2952 (N_2952,N_2822,N_2874);
nand U2953 (N_2953,N_2811,N_2825);
and U2954 (N_2954,N_2830,N_2823);
nand U2955 (N_2955,N_2894,N_2802);
nand U2956 (N_2956,N_2813,N_2830);
and U2957 (N_2957,N_2812,N_2874);
nor U2958 (N_2958,N_2832,N_2859);
and U2959 (N_2959,N_2816,N_2857);
nor U2960 (N_2960,N_2806,N_2809);
xor U2961 (N_2961,N_2876,N_2808);
nor U2962 (N_2962,N_2805,N_2827);
nor U2963 (N_2963,N_2831,N_2830);
nor U2964 (N_2964,N_2856,N_2875);
and U2965 (N_2965,N_2849,N_2885);
or U2966 (N_2966,N_2876,N_2826);
nand U2967 (N_2967,N_2816,N_2817);
nor U2968 (N_2968,N_2881,N_2888);
and U2969 (N_2969,N_2865,N_2826);
or U2970 (N_2970,N_2847,N_2877);
or U2971 (N_2971,N_2833,N_2844);
nor U2972 (N_2972,N_2833,N_2874);
nor U2973 (N_2973,N_2827,N_2823);
or U2974 (N_2974,N_2828,N_2801);
or U2975 (N_2975,N_2832,N_2827);
and U2976 (N_2976,N_2873,N_2841);
nor U2977 (N_2977,N_2814,N_2889);
or U2978 (N_2978,N_2811,N_2888);
and U2979 (N_2979,N_2864,N_2824);
or U2980 (N_2980,N_2887,N_2801);
nand U2981 (N_2981,N_2884,N_2848);
and U2982 (N_2982,N_2853,N_2874);
xor U2983 (N_2983,N_2842,N_2818);
nand U2984 (N_2984,N_2890,N_2835);
nor U2985 (N_2985,N_2897,N_2882);
nand U2986 (N_2986,N_2843,N_2870);
and U2987 (N_2987,N_2818,N_2889);
and U2988 (N_2988,N_2884,N_2837);
nand U2989 (N_2989,N_2807,N_2852);
xor U2990 (N_2990,N_2836,N_2887);
or U2991 (N_2991,N_2848,N_2815);
nor U2992 (N_2992,N_2824,N_2884);
and U2993 (N_2993,N_2866,N_2891);
and U2994 (N_2994,N_2807,N_2833);
and U2995 (N_2995,N_2812,N_2890);
and U2996 (N_2996,N_2834,N_2889);
nand U2997 (N_2997,N_2824,N_2866);
or U2998 (N_2998,N_2893,N_2878);
and U2999 (N_2999,N_2826,N_2820);
xor UO_0 (O_0,N_2982,N_2973);
nand UO_1 (O_1,N_2944,N_2913);
or UO_2 (O_2,N_2922,N_2917);
and UO_3 (O_3,N_2919,N_2906);
and UO_4 (O_4,N_2992,N_2926);
or UO_5 (O_5,N_2950,N_2966);
xor UO_6 (O_6,N_2946,N_2957);
xor UO_7 (O_7,N_2972,N_2938);
xnor UO_8 (O_8,N_2930,N_2940);
or UO_9 (O_9,N_2912,N_2942);
and UO_10 (O_10,N_2995,N_2905);
nor UO_11 (O_11,N_2978,N_2969);
nor UO_12 (O_12,N_2910,N_2999);
or UO_13 (O_13,N_2907,N_2923);
or UO_14 (O_14,N_2920,N_2932);
nand UO_15 (O_15,N_2997,N_2963);
and UO_16 (O_16,N_2918,N_2996);
xnor UO_17 (O_17,N_2953,N_2904);
nor UO_18 (O_18,N_2927,N_2988);
nor UO_19 (O_19,N_2962,N_2947);
nor UO_20 (O_20,N_2970,N_2901);
nor UO_21 (O_21,N_2937,N_2935);
xnor UO_22 (O_22,N_2921,N_2961);
or UO_23 (O_23,N_2949,N_2960);
nand UO_24 (O_24,N_2986,N_2959);
nor UO_25 (O_25,N_2990,N_2916);
and UO_26 (O_26,N_2928,N_2925);
and UO_27 (O_27,N_2943,N_2964);
or UO_28 (O_28,N_2931,N_2985);
and UO_29 (O_29,N_2902,N_2976);
and UO_30 (O_30,N_2915,N_2975);
nand UO_31 (O_31,N_2909,N_2974);
nand UO_32 (O_32,N_2936,N_2929);
or UO_33 (O_33,N_2941,N_2945);
and UO_34 (O_34,N_2993,N_2987);
nand UO_35 (O_35,N_2951,N_2952);
or UO_36 (O_36,N_2983,N_2956);
or UO_37 (O_37,N_2939,N_2971);
xor UO_38 (O_38,N_2965,N_2981);
nor UO_39 (O_39,N_2934,N_2955);
nand UO_40 (O_40,N_2911,N_2989);
xnor UO_41 (O_41,N_2977,N_2948);
xor UO_42 (O_42,N_2924,N_2979);
xnor UO_43 (O_43,N_2914,N_2933);
xnor UO_44 (O_44,N_2991,N_2903);
and UO_45 (O_45,N_2994,N_2954);
or UO_46 (O_46,N_2967,N_2958);
nand UO_47 (O_47,N_2998,N_2968);
nand UO_48 (O_48,N_2984,N_2908);
or UO_49 (O_49,N_2900,N_2980);
nor UO_50 (O_50,N_2935,N_2970);
or UO_51 (O_51,N_2900,N_2940);
xor UO_52 (O_52,N_2990,N_2998);
xnor UO_53 (O_53,N_2972,N_2946);
xnor UO_54 (O_54,N_2912,N_2995);
nand UO_55 (O_55,N_2943,N_2952);
xor UO_56 (O_56,N_2952,N_2929);
or UO_57 (O_57,N_2960,N_2971);
or UO_58 (O_58,N_2954,N_2975);
or UO_59 (O_59,N_2908,N_2987);
nand UO_60 (O_60,N_2900,N_2901);
xor UO_61 (O_61,N_2917,N_2976);
nand UO_62 (O_62,N_2995,N_2970);
nand UO_63 (O_63,N_2905,N_2909);
xor UO_64 (O_64,N_2981,N_2978);
and UO_65 (O_65,N_2924,N_2947);
or UO_66 (O_66,N_2981,N_2963);
nor UO_67 (O_67,N_2974,N_2962);
nor UO_68 (O_68,N_2927,N_2951);
nand UO_69 (O_69,N_2962,N_2970);
xor UO_70 (O_70,N_2933,N_2907);
or UO_71 (O_71,N_2974,N_2920);
or UO_72 (O_72,N_2943,N_2940);
or UO_73 (O_73,N_2999,N_2908);
xor UO_74 (O_74,N_2943,N_2983);
nor UO_75 (O_75,N_2936,N_2909);
nand UO_76 (O_76,N_2952,N_2930);
nand UO_77 (O_77,N_2970,N_2930);
nor UO_78 (O_78,N_2959,N_2932);
xor UO_79 (O_79,N_2982,N_2934);
or UO_80 (O_80,N_2975,N_2916);
nand UO_81 (O_81,N_2962,N_2918);
or UO_82 (O_82,N_2916,N_2995);
or UO_83 (O_83,N_2947,N_2970);
xor UO_84 (O_84,N_2942,N_2964);
nand UO_85 (O_85,N_2960,N_2933);
nand UO_86 (O_86,N_2921,N_2939);
nand UO_87 (O_87,N_2984,N_2927);
and UO_88 (O_88,N_2974,N_2934);
or UO_89 (O_89,N_2920,N_2955);
xnor UO_90 (O_90,N_2920,N_2996);
nand UO_91 (O_91,N_2985,N_2994);
xnor UO_92 (O_92,N_2984,N_2904);
xnor UO_93 (O_93,N_2903,N_2978);
nand UO_94 (O_94,N_2987,N_2926);
or UO_95 (O_95,N_2953,N_2982);
xnor UO_96 (O_96,N_2928,N_2927);
or UO_97 (O_97,N_2966,N_2921);
nand UO_98 (O_98,N_2935,N_2915);
or UO_99 (O_99,N_2996,N_2988);
or UO_100 (O_100,N_2971,N_2933);
nand UO_101 (O_101,N_2957,N_2942);
xnor UO_102 (O_102,N_2901,N_2953);
nor UO_103 (O_103,N_2920,N_2977);
nor UO_104 (O_104,N_2906,N_2902);
nor UO_105 (O_105,N_2958,N_2924);
nand UO_106 (O_106,N_2965,N_2950);
and UO_107 (O_107,N_2926,N_2939);
nor UO_108 (O_108,N_2991,N_2906);
or UO_109 (O_109,N_2928,N_2909);
or UO_110 (O_110,N_2925,N_2940);
and UO_111 (O_111,N_2981,N_2977);
nor UO_112 (O_112,N_2961,N_2976);
and UO_113 (O_113,N_2933,N_2936);
xnor UO_114 (O_114,N_2919,N_2930);
xor UO_115 (O_115,N_2978,N_2999);
nor UO_116 (O_116,N_2955,N_2902);
xnor UO_117 (O_117,N_2956,N_2948);
nor UO_118 (O_118,N_2973,N_2935);
xnor UO_119 (O_119,N_2989,N_2956);
or UO_120 (O_120,N_2948,N_2986);
xor UO_121 (O_121,N_2998,N_2901);
or UO_122 (O_122,N_2910,N_2959);
or UO_123 (O_123,N_2902,N_2963);
or UO_124 (O_124,N_2957,N_2984);
nand UO_125 (O_125,N_2949,N_2957);
nor UO_126 (O_126,N_2965,N_2975);
xnor UO_127 (O_127,N_2919,N_2925);
nor UO_128 (O_128,N_2986,N_2903);
and UO_129 (O_129,N_2975,N_2946);
nand UO_130 (O_130,N_2965,N_2930);
nand UO_131 (O_131,N_2956,N_2974);
nor UO_132 (O_132,N_2982,N_2998);
xnor UO_133 (O_133,N_2954,N_2916);
nand UO_134 (O_134,N_2913,N_2905);
nor UO_135 (O_135,N_2908,N_2926);
nor UO_136 (O_136,N_2912,N_2919);
nand UO_137 (O_137,N_2963,N_2925);
or UO_138 (O_138,N_2949,N_2971);
nor UO_139 (O_139,N_2937,N_2992);
or UO_140 (O_140,N_2946,N_2910);
and UO_141 (O_141,N_2968,N_2978);
or UO_142 (O_142,N_2984,N_2968);
or UO_143 (O_143,N_2991,N_2993);
xnor UO_144 (O_144,N_2986,N_2973);
or UO_145 (O_145,N_2978,N_2982);
and UO_146 (O_146,N_2923,N_2952);
and UO_147 (O_147,N_2962,N_2984);
or UO_148 (O_148,N_2916,N_2969);
or UO_149 (O_149,N_2921,N_2933);
nor UO_150 (O_150,N_2924,N_2955);
nor UO_151 (O_151,N_2914,N_2901);
xor UO_152 (O_152,N_2946,N_2920);
or UO_153 (O_153,N_2990,N_2910);
or UO_154 (O_154,N_2973,N_2944);
and UO_155 (O_155,N_2915,N_2917);
nor UO_156 (O_156,N_2926,N_2998);
nor UO_157 (O_157,N_2900,N_2906);
xnor UO_158 (O_158,N_2941,N_2909);
or UO_159 (O_159,N_2910,N_2964);
nand UO_160 (O_160,N_2986,N_2931);
or UO_161 (O_161,N_2990,N_2941);
nor UO_162 (O_162,N_2977,N_2914);
nor UO_163 (O_163,N_2987,N_2997);
nor UO_164 (O_164,N_2959,N_2907);
nor UO_165 (O_165,N_2954,N_2987);
and UO_166 (O_166,N_2915,N_2969);
and UO_167 (O_167,N_2949,N_2959);
and UO_168 (O_168,N_2983,N_2955);
or UO_169 (O_169,N_2916,N_2922);
nand UO_170 (O_170,N_2993,N_2947);
and UO_171 (O_171,N_2958,N_2954);
or UO_172 (O_172,N_2904,N_2992);
or UO_173 (O_173,N_2979,N_2945);
and UO_174 (O_174,N_2955,N_2944);
nand UO_175 (O_175,N_2968,N_2907);
nor UO_176 (O_176,N_2913,N_2941);
or UO_177 (O_177,N_2968,N_2952);
nor UO_178 (O_178,N_2916,N_2911);
or UO_179 (O_179,N_2976,N_2930);
xnor UO_180 (O_180,N_2950,N_2946);
or UO_181 (O_181,N_2906,N_2934);
xor UO_182 (O_182,N_2971,N_2921);
or UO_183 (O_183,N_2950,N_2960);
nor UO_184 (O_184,N_2929,N_2972);
nor UO_185 (O_185,N_2912,N_2946);
and UO_186 (O_186,N_2966,N_2953);
xnor UO_187 (O_187,N_2953,N_2992);
or UO_188 (O_188,N_2974,N_2953);
xnor UO_189 (O_189,N_2978,N_2917);
nand UO_190 (O_190,N_2976,N_2970);
and UO_191 (O_191,N_2936,N_2920);
xor UO_192 (O_192,N_2905,N_2924);
and UO_193 (O_193,N_2964,N_2936);
or UO_194 (O_194,N_2909,N_2978);
xor UO_195 (O_195,N_2977,N_2928);
nand UO_196 (O_196,N_2914,N_2907);
nand UO_197 (O_197,N_2970,N_2960);
or UO_198 (O_198,N_2922,N_2996);
xor UO_199 (O_199,N_2980,N_2999);
nand UO_200 (O_200,N_2988,N_2936);
and UO_201 (O_201,N_2991,N_2946);
nor UO_202 (O_202,N_2999,N_2934);
nand UO_203 (O_203,N_2986,N_2981);
or UO_204 (O_204,N_2991,N_2947);
or UO_205 (O_205,N_2978,N_2992);
xor UO_206 (O_206,N_2910,N_2916);
nand UO_207 (O_207,N_2977,N_2990);
nand UO_208 (O_208,N_2918,N_2930);
or UO_209 (O_209,N_2933,N_2978);
and UO_210 (O_210,N_2969,N_2935);
nor UO_211 (O_211,N_2915,N_2971);
nor UO_212 (O_212,N_2995,N_2971);
xnor UO_213 (O_213,N_2981,N_2983);
and UO_214 (O_214,N_2930,N_2961);
nand UO_215 (O_215,N_2901,N_2925);
xnor UO_216 (O_216,N_2991,N_2958);
or UO_217 (O_217,N_2993,N_2956);
nor UO_218 (O_218,N_2959,N_2983);
nand UO_219 (O_219,N_2931,N_2926);
nor UO_220 (O_220,N_2932,N_2935);
nand UO_221 (O_221,N_2912,N_2992);
and UO_222 (O_222,N_2998,N_2949);
nand UO_223 (O_223,N_2940,N_2986);
or UO_224 (O_224,N_2979,N_2930);
and UO_225 (O_225,N_2983,N_2919);
and UO_226 (O_226,N_2960,N_2906);
and UO_227 (O_227,N_2914,N_2994);
nand UO_228 (O_228,N_2991,N_2992);
nand UO_229 (O_229,N_2931,N_2900);
and UO_230 (O_230,N_2972,N_2981);
xnor UO_231 (O_231,N_2994,N_2905);
or UO_232 (O_232,N_2958,N_2956);
nand UO_233 (O_233,N_2957,N_2910);
or UO_234 (O_234,N_2914,N_2997);
and UO_235 (O_235,N_2908,N_2932);
or UO_236 (O_236,N_2927,N_2979);
nand UO_237 (O_237,N_2987,N_2967);
nor UO_238 (O_238,N_2987,N_2988);
nor UO_239 (O_239,N_2974,N_2937);
and UO_240 (O_240,N_2909,N_2995);
nor UO_241 (O_241,N_2970,N_2977);
and UO_242 (O_242,N_2994,N_2968);
nand UO_243 (O_243,N_2978,N_2950);
or UO_244 (O_244,N_2971,N_2917);
xnor UO_245 (O_245,N_2966,N_2968);
or UO_246 (O_246,N_2919,N_2980);
nand UO_247 (O_247,N_2913,N_2914);
nand UO_248 (O_248,N_2980,N_2940);
nand UO_249 (O_249,N_2955,N_2961);
nor UO_250 (O_250,N_2924,N_2988);
and UO_251 (O_251,N_2950,N_2939);
nor UO_252 (O_252,N_2987,N_2930);
or UO_253 (O_253,N_2906,N_2995);
and UO_254 (O_254,N_2981,N_2951);
and UO_255 (O_255,N_2957,N_2906);
nor UO_256 (O_256,N_2998,N_2985);
xnor UO_257 (O_257,N_2970,N_2940);
xnor UO_258 (O_258,N_2936,N_2944);
nor UO_259 (O_259,N_2922,N_2968);
nand UO_260 (O_260,N_2950,N_2986);
nor UO_261 (O_261,N_2996,N_2928);
nand UO_262 (O_262,N_2999,N_2989);
or UO_263 (O_263,N_2938,N_2921);
xnor UO_264 (O_264,N_2932,N_2902);
and UO_265 (O_265,N_2903,N_2988);
nand UO_266 (O_266,N_2988,N_2968);
nand UO_267 (O_267,N_2929,N_2949);
nand UO_268 (O_268,N_2985,N_2977);
nor UO_269 (O_269,N_2933,N_2928);
and UO_270 (O_270,N_2954,N_2900);
xnor UO_271 (O_271,N_2916,N_2907);
and UO_272 (O_272,N_2923,N_2973);
and UO_273 (O_273,N_2967,N_2981);
and UO_274 (O_274,N_2935,N_2992);
and UO_275 (O_275,N_2985,N_2921);
and UO_276 (O_276,N_2996,N_2933);
or UO_277 (O_277,N_2988,N_2998);
nand UO_278 (O_278,N_2933,N_2959);
and UO_279 (O_279,N_2906,N_2992);
xnor UO_280 (O_280,N_2975,N_2956);
or UO_281 (O_281,N_2990,N_2964);
nand UO_282 (O_282,N_2910,N_2920);
and UO_283 (O_283,N_2969,N_2920);
and UO_284 (O_284,N_2901,N_2911);
nor UO_285 (O_285,N_2935,N_2994);
nor UO_286 (O_286,N_2924,N_2972);
or UO_287 (O_287,N_2956,N_2980);
and UO_288 (O_288,N_2925,N_2976);
nor UO_289 (O_289,N_2902,N_2912);
and UO_290 (O_290,N_2997,N_2957);
nor UO_291 (O_291,N_2942,N_2913);
nand UO_292 (O_292,N_2997,N_2990);
nor UO_293 (O_293,N_2917,N_2935);
and UO_294 (O_294,N_2913,N_2933);
nor UO_295 (O_295,N_2913,N_2934);
or UO_296 (O_296,N_2998,N_2932);
or UO_297 (O_297,N_2966,N_2911);
or UO_298 (O_298,N_2962,N_2995);
nor UO_299 (O_299,N_2982,N_2933);
and UO_300 (O_300,N_2905,N_2923);
nor UO_301 (O_301,N_2934,N_2985);
and UO_302 (O_302,N_2967,N_2995);
and UO_303 (O_303,N_2940,N_2969);
xnor UO_304 (O_304,N_2993,N_2900);
nand UO_305 (O_305,N_2983,N_2949);
nand UO_306 (O_306,N_2948,N_2910);
nor UO_307 (O_307,N_2904,N_2954);
nand UO_308 (O_308,N_2902,N_2939);
nor UO_309 (O_309,N_2969,N_2942);
xnor UO_310 (O_310,N_2946,N_2960);
and UO_311 (O_311,N_2942,N_2996);
nand UO_312 (O_312,N_2920,N_2970);
and UO_313 (O_313,N_2949,N_2936);
nand UO_314 (O_314,N_2942,N_2951);
and UO_315 (O_315,N_2970,N_2932);
xnor UO_316 (O_316,N_2946,N_2941);
nand UO_317 (O_317,N_2929,N_2917);
and UO_318 (O_318,N_2919,N_2926);
nor UO_319 (O_319,N_2917,N_2924);
nand UO_320 (O_320,N_2934,N_2901);
nand UO_321 (O_321,N_2953,N_2925);
or UO_322 (O_322,N_2920,N_2966);
or UO_323 (O_323,N_2933,N_2969);
nand UO_324 (O_324,N_2964,N_2978);
and UO_325 (O_325,N_2951,N_2988);
nand UO_326 (O_326,N_2983,N_2929);
and UO_327 (O_327,N_2999,N_2947);
nor UO_328 (O_328,N_2968,N_2955);
nor UO_329 (O_329,N_2905,N_2982);
and UO_330 (O_330,N_2918,N_2964);
nand UO_331 (O_331,N_2922,N_2934);
and UO_332 (O_332,N_2962,N_2986);
or UO_333 (O_333,N_2967,N_2916);
nor UO_334 (O_334,N_2965,N_2996);
nor UO_335 (O_335,N_2906,N_2921);
and UO_336 (O_336,N_2907,N_2990);
and UO_337 (O_337,N_2994,N_2996);
or UO_338 (O_338,N_2948,N_2940);
nand UO_339 (O_339,N_2975,N_2987);
nor UO_340 (O_340,N_2963,N_2960);
and UO_341 (O_341,N_2979,N_2929);
xnor UO_342 (O_342,N_2981,N_2953);
nor UO_343 (O_343,N_2973,N_2967);
and UO_344 (O_344,N_2940,N_2913);
or UO_345 (O_345,N_2916,N_2937);
or UO_346 (O_346,N_2915,N_2902);
nor UO_347 (O_347,N_2969,N_2988);
xnor UO_348 (O_348,N_2980,N_2944);
nand UO_349 (O_349,N_2941,N_2938);
xnor UO_350 (O_350,N_2947,N_2954);
nand UO_351 (O_351,N_2931,N_2955);
xnor UO_352 (O_352,N_2929,N_2925);
or UO_353 (O_353,N_2908,N_2920);
xor UO_354 (O_354,N_2962,N_2988);
or UO_355 (O_355,N_2919,N_2981);
nor UO_356 (O_356,N_2999,N_2956);
or UO_357 (O_357,N_2995,N_2921);
nand UO_358 (O_358,N_2954,N_2921);
and UO_359 (O_359,N_2927,N_2914);
xor UO_360 (O_360,N_2912,N_2962);
nor UO_361 (O_361,N_2975,N_2993);
nor UO_362 (O_362,N_2986,N_2902);
and UO_363 (O_363,N_2967,N_2955);
nand UO_364 (O_364,N_2967,N_2956);
and UO_365 (O_365,N_2989,N_2967);
and UO_366 (O_366,N_2945,N_2959);
xnor UO_367 (O_367,N_2921,N_2988);
nor UO_368 (O_368,N_2959,N_2901);
nor UO_369 (O_369,N_2933,N_2965);
and UO_370 (O_370,N_2934,N_2953);
or UO_371 (O_371,N_2906,N_2956);
xnor UO_372 (O_372,N_2951,N_2928);
nand UO_373 (O_373,N_2930,N_2955);
and UO_374 (O_374,N_2924,N_2956);
nand UO_375 (O_375,N_2992,N_2990);
or UO_376 (O_376,N_2963,N_2928);
or UO_377 (O_377,N_2910,N_2938);
nand UO_378 (O_378,N_2928,N_2912);
nor UO_379 (O_379,N_2983,N_2921);
xor UO_380 (O_380,N_2986,N_2991);
nor UO_381 (O_381,N_2938,N_2948);
or UO_382 (O_382,N_2933,N_2966);
xnor UO_383 (O_383,N_2994,N_2943);
nand UO_384 (O_384,N_2906,N_2909);
xor UO_385 (O_385,N_2964,N_2915);
or UO_386 (O_386,N_2960,N_2905);
xnor UO_387 (O_387,N_2986,N_2995);
and UO_388 (O_388,N_2902,N_2997);
or UO_389 (O_389,N_2930,N_2931);
nor UO_390 (O_390,N_2924,N_2935);
xor UO_391 (O_391,N_2940,N_2956);
nor UO_392 (O_392,N_2958,N_2909);
and UO_393 (O_393,N_2954,N_2966);
nand UO_394 (O_394,N_2925,N_2930);
and UO_395 (O_395,N_2991,N_2931);
nor UO_396 (O_396,N_2999,N_2909);
nor UO_397 (O_397,N_2920,N_2978);
nand UO_398 (O_398,N_2917,N_2972);
or UO_399 (O_399,N_2960,N_2993);
xor UO_400 (O_400,N_2981,N_2979);
xor UO_401 (O_401,N_2951,N_2992);
nor UO_402 (O_402,N_2936,N_2916);
or UO_403 (O_403,N_2952,N_2946);
or UO_404 (O_404,N_2991,N_2943);
or UO_405 (O_405,N_2968,N_2967);
and UO_406 (O_406,N_2980,N_2913);
xnor UO_407 (O_407,N_2987,N_2961);
xnor UO_408 (O_408,N_2972,N_2999);
or UO_409 (O_409,N_2906,N_2981);
nor UO_410 (O_410,N_2906,N_2987);
xnor UO_411 (O_411,N_2957,N_2944);
nand UO_412 (O_412,N_2988,N_2970);
nor UO_413 (O_413,N_2975,N_2979);
xnor UO_414 (O_414,N_2921,N_2973);
nand UO_415 (O_415,N_2964,N_2940);
or UO_416 (O_416,N_2982,N_2922);
nand UO_417 (O_417,N_2910,N_2905);
nor UO_418 (O_418,N_2968,N_2956);
nor UO_419 (O_419,N_2940,N_2991);
nor UO_420 (O_420,N_2940,N_2963);
nor UO_421 (O_421,N_2925,N_2911);
and UO_422 (O_422,N_2935,N_2978);
or UO_423 (O_423,N_2972,N_2978);
xnor UO_424 (O_424,N_2975,N_2928);
xnor UO_425 (O_425,N_2966,N_2994);
and UO_426 (O_426,N_2998,N_2963);
or UO_427 (O_427,N_2917,N_2989);
xor UO_428 (O_428,N_2907,N_2991);
and UO_429 (O_429,N_2963,N_2976);
nor UO_430 (O_430,N_2919,N_2967);
nand UO_431 (O_431,N_2984,N_2910);
nand UO_432 (O_432,N_2960,N_2959);
and UO_433 (O_433,N_2909,N_2973);
or UO_434 (O_434,N_2982,N_2950);
nand UO_435 (O_435,N_2948,N_2947);
xnor UO_436 (O_436,N_2991,N_2956);
nand UO_437 (O_437,N_2939,N_2984);
nand UO_438 (O_438,N_2969,N_2908);
xor UO_439 (O_439,N_2917,N_2943);
nor UO_440 (O_440,N_2916,N_2970);
nor UO_441 (O_441,N_2905,N_2967);
or UO_442 (O_442,N_2930,N_2959);
xnor UO_443 (O_443,N_2976,N_2957);
and UO_444 (O_444,N_2974,N_2961);
nor UO_445 (O_445,N_2939,N_2912);
and UO_446 (O_446,N_2961,N_2964);
xor UO_447 (O_447,N_2984,N_2979);
nand UO_448 (O_448,N_2961,N_2932);
nor UO_449 (O_449,N_2977,N_2967);
and UO_450 (O_450,N_2976,N_2975);
nand UO_451 (O_451,N_2927,N_2926);
or UO_452 (O_452,N_2944,N_2935);
nand UO_453 (O_453,N_2948,N_2915);
nand UO_454 (O_454,N_2967,N_2949);
xor UO_455 (O_455,N_2937,N_2989);
and UO_456 (O_456,N_2934,N_2928);
and UO_457 (O_457,N_2919,N_2979);
nor UO_458 (O_458,N_2930,N_2914);
nand UO_459 (O_459,N_2921,N_2901);
nand UO_460 (O_460,N_2998,N_2903);
or UO_461 (O_461,N_2900,N_2950);
or UO_462 (O_462,N_2985,N_2912);
nand UO_463 (O_463,N_2995,N_2919);
nand UO_464 (O_464,N_2945,N_2978);
or UO_465 (O_465,N_2916,N_2962);
nand UO_466 (O_466,N_2909,N_2940);
xor UO_467 (O_467,N_2988,N_2925);
and UO_468 (O_468,N_2936,N_2992);
and UO_469 (O_469,N_2949,N_2916);
or UO_470 (O_470,N_2974,N_2970);
and UO_471 (O_471,N_2901,N_2938);
and UO_472 (O_472,N_2991,N_2953);
or UO_473 (O_473,N_2913,N_2938);
nor UO_474 (O_474,N_2986,N_2980);
nor UO_475 (O_475,N_2945,N_2942);
xor UO_476 (O_476,N_2928,N_2959);
nor UO_477 (O_477,N_2987,N_2958);
xor UO_478 (O_478,N_2961,N_2928);
xor UO_479 (O_479,N_2994,N_2902);
or UO_480 (O_480,N_2935,N_2990);
or UO_481 (O_481,N_2998,N_2987);
and UO_482 (O_482,N_2910,N_2904);
nand UO_483 (O_483,N_2928,N_2920);
nand UO_484 (O_484,N_2925,N_2958);
nor UO_485 (O_485,N_2996,N_2959);
nand UO_486 (O_486,N_2963,N_2935);
xor UO_487 (O_487,N_2980,N_2933);
and UO_488 (O_488,N_2954,N_2932);
and UO_489 (O_489,N_2951,N_2954);
nor UO_490 (O_490,N_2933,N_2994);
nor UO_491 (O_491,N_2974,N_2921);
or UO_492 (O_492,N_2937,N_2909);
nand UO_493 (O_493,N_2983,N_2977);
nand UO_494 (O_494,N_2927,N_2949);
and UO_495 (O_495,N_2918,N_2900);
or UO_496 (O_496,N_2955,N_2949);
or UO_497 (O_497,N_2979,N_2937);
nor UO_498 (O_498,N_2958,N_2971);
nor UO_499 (O_499,N_2955,N_2911);
endmodule