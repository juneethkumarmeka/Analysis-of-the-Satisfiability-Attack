module basic_1000_10000_1500_50_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_522,In_892);
nor U1 (N_1,In_786,In_176);
or U2 (N_2,In_262,In_371);
xor U3 (N_3,In_875,In_234);
nor U4 (N_4,In_747,In_886);
or U5 (N_5,In_225,In_963);
and U6 (N_6,In_964,In_622);
xor U7 (N_7,In_128,In_563);
or U8 (N_8,In_19,In_75);
and U9 (N_9,In_383,In_69);
xnor U10 (N_10,In_707,In_310);
and U11 (N_11,In_161,In_788);
or U12 (N_12,In_903,In_385);
xor U13 (N_13,In_384,In_490);
and U14 (N_14,In_609,In_560);
and U15 (N_15,In_743,In_917);
nand U16 (N_16,In_977,In_315);
nand U17 (N_17,In_338,In_257);
or U18 (N_18,In_523,In_95);
nor U19 (N_19,In_779,In_773);
nor U20 (N_20,In_712,In_35);
and U21 (N_21,In_246,In_623);
and U22 (N_22,In_555,In_568);
and U23 (N_23,In_227,In_954);
xor U24 (N_24,In_153,In_601);
or U25 (N_25,In_143,In_898);
nand U26 (N_26,In_349,In_0);
xnor U27 (N_27,In_540,In_855);
and U28 (N_28,In_108,In_758);
xnor U29 (N_29,In_214,In_993);
or U30 (N_30,In_27,In_318);
nand U31 (N_31,In_33,In_613);
or U32 (N_32,In_413,In_579);
nand U33 (N_33,In_115,In_183);
and U34 (N_34,In_147,In_746);
nor U35 (N_35,In_137,In_829);
nor U36 (N_36,In_464,In_37);
or U37 (N_37,In_317,In_967);
nand U38 (N_38,In_651,In_703);
and U39 (N_39,In_530,In_485);
or U40 (N_40,In_419,In_333);
xnor U41 (N_41,In_269,In_483);
nand U42 (N_42,In_918,In_253);
and U43 (N_43,In_52,In_996);
and U44 (N_44,In_70,In_665);
nor U45 (N_45,In_328,In_500);
nor U46 (N_46,In_724,In_201);
and U47 (N_47,In_495,In_940);
nand U48 (N_48,In_685,In_438);
and U49 (N_49,In_840,In_787);
xnor U50 (N_50,In_29,In_66);
nand U51 (N_51,In_529,In_185);
and U52 (N_52,In_586,In_812);
xor U53 (N_53,In_451,In_138);
nand U54 (N_54,In_297,In_804);
nand U55 (N_55,In_611,In_193);
nand U56 (N_56,In_430,In_99);
nand U57 (N_57,In_345,In_591);
and U58 (N_58,In_380,In_843);
xnor U59 (N_59,In_807,In_484);
nor U60 (N_60,In_157,In_325);
nor U61 (N_61,In_550,In_7);
or U62 (N_62,In_145,In_155);
and U63 (N_63,In_352,In_23);
nand U64 (N_64,In_179,In_369);
or U65 (N_65,In_319,In_684);
and U66 (N_66,In_302,In_267);
nand U67 (N_67,In_806,In_111);
xor U68 (N_68,In_882,In_344);
xnor U69 (N_69,In_753,In_931);
and U70 (N_70,In_661,In_113);
nor U71 (N_71,In_312,In_721);
nor U72 (N_72,In_229,In_629);
nand U73 (N_73,In_190,In_49);
nand U74 (N_74,In_194,In_182);
xnor U75 (N_75,In_224,In_118);
nor U76 (N_76,In_838,In_507);
xor U77 (N_77,In_503,In_238);
or U78 (N_78,In_402,In_744);
or U79 (N_79,In_720,In_250);
or U80 (N_80,In_915,In_696);
nor U81 (N_81,In_578,In_283);
and U82 (N_82,In_692,In_22);
xnor U83 (N_83,In_277,In_204);
xor U84 (N_84,In_78,In_471);
or U85 (N_85,In_114,In_274);
nand U86 (N_86,In_705,In_637);
and U87 (N_87,In_472,In_48);
nor U88 (N_88,In_899,In_988);
nor U89 (N_89,In_557,In_859);
nor U90 (N_90,In_442,In_947);
and U91 (N_91,In_361,In_456);
nand U92 (N_92,In_872,In_924);
nor U93 (N_93,In_458,In_534);
and U94 (N_94,In_434,In_187);
nor U95 (N_95,In_945,In_978);
xnor U96 (N_96,In_748,In_429);
nor U97 (N_97,In_482,In_687);
or U98 (N_98,In_156,In_62);
xnor U99 (N_99,In_63,In_260);
or U100 (N_100,In_842,In_248);
nand U101 (N_101,In_850,In_223);
and U102 (N_102,In_97,In_528);
nor U103 (N_103,In_314,In_981);
nand U104 (N_104,In_533,In_195);
nand U105 (N_105,In_904,In_643);
or U106 (N_106,In_307,In_331);
xor U107 (N_107,In_5,In_837);
nand U108 (N_108,In_551,In_582);
and U109 (N_109,In_891,In_572);
xnor U110 (N_110,In_895,In_293);
xor U111 (N_111,In_83,In_202);
or U112 (N_112,In_117,In_87);
xnor U113 (N_113,In_868,In_184);
xnor U114 (N_114,In_491,In_818);
and U115 (N_115,In_514,In_797);
nor U116 (N_116,In_865,In_864);
nand U117 (N_117,In_85,In_570);
nor U118 (N_118,In_771,In_760);
xor U119 (N_119,In_2,In_695);
or U120 (N_120,In_16,In_792);
xnor U121 (N_121,In_324,In_520);
or U122 (N_122,In_10,In_391);
nor U123 (N_123,In_50,In_706);
and U124 (N_124,In_857,In_228);
or U125 (N_125,In_765,In_326);
xnor U126 (N_126,In_983,In_997);
nor U127 (N_127,In_546,In_732);
nand U128 (N_128,In_263,In_406);
xor U129 (N_129,In_477,In_962);
or U130 (N_130,In_286,In_112);
nor U131 (N_131,In_603,In_496);
xnor U132 (N_132,In_284,In_498);
or U133 (N_133,In_306,In_989);
or U134 (N_134,In_770,In_71);
and U135 (N_135,In_34,In_614);
or U136 (N_136,In_766,In_567);
xnor U137 (N_137,In_655,In_359);
nor U138 (N_138,In_251,In_921);
xnor U139 (N_139,In_254,In_60);
nor U140 (N_140,In_606,In_679);
nor U141 (N_141,In_144,In_207);
and U142 (N_142,In_473,In_203);
and U143 (N_143,In_59,In_965);
nor U144 (N_144,In_311,In_971);
or U145 (N_145,In_320,In_119);
and U146 (N_146,In_421,In_11);
or U147 (N_147,In_803,In_437);
nand U148 (N_148,In_608,In_780);
or U149 (N_149,In_387,In_15);
xor U150 (N_150,In_124,In_913);
xor U151 (N_151,In_681,In_98);
or U152 (N_152,In_39,In_762);
and U153 (N_153,In_823,In_867);
and U154 (N_154,In_175,In_920);
nand U155 (N_155,In_313,In_463);
and U156 (N_156,In_493,In_726);
xor U157 (N_157,In_628,In_951);
nand U158 (N_158,In_937,In_12);
nand U159 (N_159,In_43,In_862);
and U160 (N_160,In_191,In_552);
nor U161 (N_161,In_105,In_616);
or U162 (N_162,In_300,In_32);
or U163 (N_163,In_587,In_44);
nor U164 (N_164,In_497,In_755);
or U165 (N_165,In_648,In_357);
nor U166 (N_166,In_537,In_288);
nor U167 (N_167,In_475,In_833);
nand U168 (N_168,In_217,In_323);
or U169 (N_169,In_30,In_411);
nor U170 (N_170,In_824,In_372);
and U171 (N_171,In_970,In_708);
xor U172 (N_172,In_26,In_410);
nand U173 (N_173,In_960,In_910);
xor U174 (N_174,In_795,In_258);
nand U175 (N_175,In_660,In_730);
and U176 (N_176,In_856,In_925);
or U177 (N_177,In_547,In_757);
and U178 (N_178,In_675,In_177);
xnor U179 (N_179,In_256,In_88);
nor U180 (N_180,In_104,In_991);
nand U181 (N_181,In_447,In_426);
nand U182 (N_182,In_948,In_337);
or U183 (N_183,In_285,In_908);
nand U184 (N_184,In_887,In_249);
xor U185 (N_185,In_198,In_569);
nand U186 (N_186,In_649,In_662);
nor U187 (N_187,In_336,In_735);
nand U188 (N_188,In_96,In_602);
and U189 (N_189,In_393,In_992);
and U190 (N_190,In_102,In_47);
nand U191 (N_191,In_808,In_553);
and U192 (N_192,In_536,In_308);
nand U193 (N_193,In_222,In_682);
xor U194 (N_194,In_358,In_980);
nor U195 (N_195,In_819,In_860);
xnor U196 (N_196,In_723,In_683);
and U197 (N_197,In_929,In_905);
xnor U198 (N_198,In_135,In_890);
or U199 (N_199,In_132,In_666);
or U200 (N_200,In_470,N_36);
and U201 (N_201,In_226,In_825);
nand U202 (N_202,In_186,In_301);
xor U203 (N_203,In_424,N_7);
xnor U204 (N_204,In_509,In_631);
xor U205 (N_205,In_621,In_901);
xnor U206 (N_206,In_531,In_791);
xnor U207 (N_207,In_973,In_211);
xnor U208 (N_208,N_97,N_62);
xnor U209 (N_209,N_124,In_669);
nand U210 (N_210,In_617,In_640);
and U211 (N_211,N_106,In_14);
xor U212 (N_212,In_366,N_59);
and U213 (N_213,In_577,In_386);
xor U214 (N_214,In_756,In_524);
or U215 (N_215,In_869,In_879);
or U216 (N_216,In_441,N_127);
nor U217 (N_217,In_595,N_185);
nand U218 (N_218,In_738,N_177);
nor U219 (N_219,In_150,In_428);
nand U220 (N_220,N_0,In_405);
or U221 (N_221,In_374,In_581);
nand U222 (N_222,In_893,In_133);
and U223 (N_223,In_987,In_761);
nand U224 (N_224,In_65,N_33);
xnor U225 (N_225,In_403,In_585);
xor U226 (N_226,In_916,N_32);
nand U227 (N_227,In_782,N_152);
and U228 (N_228,N_56,In_880);
or U229 (N_229,N_120,In_299);
nor U230 (N_230,In_169,In_445);
nand U231 (N_231,In_180,In_774);
and U232 (N_232,In_691,In_487);
and U233 (N_233,In_734,In_953);
xnor U234 (N_234,In_397,In_433);
nand U235 (N_235,In_443,In_517);
xor U236 (N_236,In_516,In_21);
nor U237 (N_237,N_2,In_817);
nor U238 (N_238,In_273,In_478);
or U239 (N_239,N_49,In_363);
nor U240 (N_240,In_479,In_172);
nor U241 (N_241,In_474,In_876);
and U242 (N_242,N_176,In_995);
nor U243 (N_243,In_664,N_61);
or U244 (N_244,In_233,N_137);
xor U245 (N_245,N_25,In_573);
xnor U246 (N_246,In_844,N_20);
xnor U247 (N_247,N_28,In_106);
and U248 (N_248,In_330,In_676);
nand U249 (N_249,N_156,N_86);
and U250 (N_250,In_266,N_47);
xnor U251 (N_251,In_545,In_519);
or U252 (N_252,In_165,In_515);
nor U253 (N_253,In_728,N_46);
nor U254 (N_254,In_392,In_670);
nor U255 (N_255,N_128,N_15);
or U256 (N_256,In_206,In_576);
or U257 (N_257,In_943,In_784);
and U258 (N_258,In_835,In_541);
or U259 (N_259,In_974,N_38);
or U260 (N_260,In_466,In_914);
and U261 (N_261,In_923,In_151);
and U262 (N_262,In_526,In_972);
and U263 (N_263,N_173,In_42);
xnor U264 (N_264,N_72,In_134);
or U265 (N_265,In_295,In_814);
xnor U266 (N_266,N_68,In_84);
or U267 (N_267,In_455,In_239);
nand U268 (N_268,In_598,In_863);
nand U269 (N_269,In_334,In_713);
xor U270 (N_270,In_122,In_347);
nor U271 (N_271,In_240,In_874);
or U272 (N_272,N_90,N_44);
and U273 (N_273,N_50,In_715);
nand U274 (N_274,In_241,In_298);
nor U275 (N_275,In_3,In_28);
and U276 (N_276,In_316,N_163);
nor U277 (N_277,In_982,In_457);
or U278 (N_278,In_909,N_27);
and U279 (N_279,In_750,In_73);
and U280 (N_280,In_271,In_830);
nor U281 (N_281,In_678,N_131);
and U282 (N_282,In_689,In_367);
xnor U283 (N_283,In_976,In_373);
and U284 (N_284,In_646,N_85);
and U285 (N_285,In_31,In_499);
nand U286 (N_286,In_813,In_647);
nor U287 (N_287,N_89,N_79);
and U288 (N_288,In_645,In_189);
nor U289 (N_289,N_111,In_290);
xor U290 (N_290,In_884,In_615);
nor U291 (N_291,In_638,In_61);
nor U292 (N_292,In_408,In_17);
xnor U293 (N_293,In_170,N_114);
nor U294 (N_294,In_888,N_199);
xnor U295 (N_295,In_955,In_751);
or U296 (N_296,N_103,N_21);
xor U297 (N_297,N_112,In_130);
and U298 (N_298,N_149,In_8);
xnor U299 (N_299,In_894,In_624);
or U300 (N_300,N_168,N_166);
xor U301 (N_301,In_208,In_821);
and U302 (N_302,N_117,In_140);
xor U303 (N_303,N_3,In_449);
nor U304 (N_304,N_40,In_935);
nand U305 (N_305,In_321,In_816);
nand U306 (N_306,N_133,In_627);
nand U307 (N_307,In_532,In_435);
and U308 (N_308,In_854,N_75);
nand U309 (N_309,In_396,In_303);
and U310 (N_310,N_6,In_858);
xor U311 (N_311,In_348,In_527);
and U312 (N_312,In_4,In_938);
xor U313 (N_313,In_282,In_467);
nor U314 (N_314,In_412,In_196);
nor U315 (N_315,In_716,In_346);
and U316 (N_316,In_439,In_985);
xor U317 (N_317,In_242,N_78);
nor U318 (N_318,In_680,In_535);
nand U319 (N_319,In_969,N_150);
and U320 (N_320,In_959,In_852);
nand U321 (N_321,In_593,In_107);
and U322 (N_322,In_356,In_469);
nand U323 (N_323,In_53,In_45);
nor U324 (N_324,In_436,In_604);
nand U325 (N_325,N_9,In_897);
xor U326 (N_326,In_230,In_278);
or U327 (N_327,In_280,N_188);
nor U328 (N_328,In_861,N_161);
and U329 (N_329,In_141,In_763);
and U330 (N_330,In_889,In_885);
or U331 (N_331,In_600,In_740);
nand U332 (N_332,In_801,In_453);
xnor U333 (N_333,In_832,In_178);
xor U334 (N_334,N_109,In_998);
or U335 (N_335,In_166,In_667);
xnor U336 (N_336,N_57,In_544);
nor U337 (N_337,N_34,In_116);
xnor U338 (N_338,In_902,In_272);
and U339 (N_339,In_494,In_120);
nand U340 (N_340,In_422,In_364);
nor U341 (N_341,N_157,In_936);
and U342 (N_342,In_163,In_827);
xnor U343 (N_343,In_244,In_919);
xor U344 (N_344,N_64,In_934);
nor U345 (N_345,In_454,In_719);
nand U346 (N_346,In_745,In_231);
nor U347 (N_347,In_409,N_105);
xnor U348 (N_348,N_71,In_376);
nand U349 (N_349,In_633,In_332);
nor U350 (N_350,In_561,In_710);
nand U351 (N_351,In_656,N_180);
xor U352 (N_352,In_944,In_404);
and U353 (N_353,N_193,In_518);
or U354 (N_354,In_462,In_381);
nor U355 (N_355,In_619,In_820);
nor U356 (N_356,In_146,In_18);
nor U357 (N_357,In_459,N_186);
nor U358 (N_358,In_542,In_778);
nor U359 (N_359,In_79,In_41);
xnor U360 (N_360,In_711,In_802);
or U361 (N_361,In_956,In_181);
and U362 (N_362,In_737,In_704);
or U363 (N_363,In_164,In_407);
nor U364 (N_364,In_583,N_4);
or U365 (N_365,N_122,In_123);
nor U366 (N_366,N_43,N_140);
xnor U367 (N_367,N_91,In_939);
nor U368 (N_368,In_883,In_360);
and U369 (N_369,N_100,In_370);
and U370 (N_370,In_694,In_121);
or U371 (N_371,In_510,N_23);
nand U372 (N_372,N_102,In_235);
or U373 (N_373,In_160,In_663);
and U374 (N_374,In_129,In_793);
xor U375 (N_375,In_390,In_975);
nand U376 (N_376,N_74,In_846);
and U377 (N_377,In_539,In_736);
and U378 (N_378,In_605,In_174);
nand U379 (N_379,In_722,In_871);
nand U380 (N_380,In_218,In_91);
nand U381 (N_381,N_169,In_72);
nor U382 (N_382,In_109,In_565);
nand U383 (N_383,In_610,In_866);
or U384 (N_384,In_543,In_36);
xor U385 (N_385,In_221,N_42);
nand U386 (N_386,In_574,In_1);
or U387 (N_387,N_70,In_968);
or U388 (N_388,In_461,N_179);
nor U389 (N_389,In_775,N_10);
nor U390 (N_390,In_417,In_949);
nor U391 (N_391,In_725,In_168);
and U392 (N_392,In_54,In_425);
xnor U393 (N_393,N_51,In_329);
or U394 (N_394,N_13,In_268);
or U395 (N_395,In_768,In_596);
and U396 (N_396,N_58,In_13);
xnor U397 (N_397,N_191,In_566);
xnor U398 (N_398,In_922,N_184);
or U399 (N_399,In_486,In_379);
and U400 (N_400,In_783,In_252);
nand U401 (N_401,N_12,N_383);
or U402 (N_402,N_96,N_260);
nor U403 (N_403,In_100,N_339);
and U404 (N_404,In_154,N_116);
or U405 (N_405,In_94,In_158);
xnor U406 (N_406,In_382,N_393);
nor U407 (N_407,In_580,N_235);
nor U408 (N_408,In_831,N_282);
nor U409 (N_409,In_632,N_175);
xnor U410 (N_410,In_673,N_160);
nor U411 (N_411,N_305,In_847);
xnor U412 (N_412,N_347,In_492);
xor U413 (N_413,N_399,N_215);
nand U414 (N_414,In_64,N_349);
xnor U415 (N_415,In_279,In_353);
xor U416 (N_416,N_338,N_333);
and U417 (N_417,In_148,In_607);
or U418 (N_418,In_489,N_182);
nand U419 (N_419,In_237,In_834);
nand U420 (N_420,In_247,N_181);
nand U421 (N_421,N_95,In_618);
nand U422 (N_422,N_279,N_172);
xor U423 (N_423,In_167,In_504);
xor U424 (N_424,In_139,N_225);
xor U425 (N_425,In_769,N_315);
nand U426 (N_426,In_400,In_809);
xnor U427 (N_427,N_271,In_521);
and U428 (N_428,In_912,In_414);
or U429 (N_429,In_811,N_217);
and U430 (N_430,N_190,N_17);
and U431 (N_431,N_368,In_709);
and U432 (N_432,N_321,N_268);
nand U433 (N_433,N_344,N_266);
xnor U434 (N_434,N_272,In_418);
and U435 (N_435,In_597,N_8);
nor U436 (N_436,In_839,In_990);
nand U437 (N_437,In_508,In_209);
or U438 (N_438,In_512,N_234);
xor U439 (N_439,In_92,N_285);
nor U440 (N_440,N_247,In_881);
or U441 (N_441,N_357,N_249);
or U442 (N_442,N_206,N_54);
nand U443 (N_443,In_432,N_269);
or U444 (N_444,N_147,N_389);
and U445 (N_445,N_262,In_501);
xor U446 (N_446,N_76,In_671);
or U447 (N_447,N_297,In_717);
nand U448 (N_448,N_370,N_108);
xor U449 (N_449,N_259,N_65);
nor U450 (N_450,N_245,In_986);
nor U451 (N_451,N_254,N_376);
or U452 (N_452,N_45,In_688);
or U453 (N_453,In_625,In_245);
or U454 (N_454,In_25,In_575);
nand U455 (N_455,N_1,N_159);
xor U456 (N_456,In_700,In_80);
nor U457 (N_457,N_380,N_350);
or U458 (N_458,N_126,In_742);
nor U459 (N_459,N_165,In_415);
nor U460 (N_460,N_301,N_219);
and U461 (N_461,In_327,N_312);
or U462 (N_462,In_427,In_767);
xor U463 (N_463,In_562,In_296);
nand U464 (N_464,In_828,N_281);
and U465 (N_465,In_335,N_31);
or U466 (N_466,N_200,N_293);
and U467 (N_467,N_369,N_80);
xor U468 (N_468,In_354,N_53);
nor U469 (N_469,N_241,N_29);
nand U470 (N_470,In_729,In_588);
nand U471 (N_471,N_385,In_878);
or U472 (N_472,In_136,N_387);
xnor U473 (N_473,In_220,In_261);
or U474 (N_474,In_900,N_208);
nand U475 (N_475,In_255,N_189);
or U476 (N_476,N_130,N_290);
nand U477 (N_477,In_961,N_198);
nand U478 (N_478,N_238,In_873);
nand U479 (N_479,N_224,In_906);
or U480 (N_480,N_278,N_244);
and U481 (N_481,N_318,In_110);
nand U482 (N_482,N_360,N_107);
and U483 (N_483,In_86,N_231);
nor U484 (N_484,N_221,N_248);
nor U485 (N_485,In_171,In_126);
xnor U486 (N_486,N_220,In_309);
nor U487 (N_487,In_232,In_644);
xnor U488 (N_488,In_173,N_382);
and U489 (N_489,In_481,In_636);
nor U490 (N_490,N_311,N_288);
and U491 (N_491,In_423,In_375);
nand U492 (N_492,In_594,N_30);
nand U493 (N_493,N_125,In_103);
nor U494 (N_494,In_957,N_313);
or U495 (N_495,N_243,In_243);
xnor U496 (N_496,In_394,In_657);
xnor U497 (N_497,N_320,In_210);
xor U498 (N_498,N_236,N_202);
or U499 (N_499,In_641,N_162);
nor U500 (N_500,N_246,N_229);
or U501 (N_501,N_194,N_303);
and U502 (N_502,In_450,N_239);
xor U503 (N_503,In_149,In_815);
or U504 (N_504,In_294,In_589);
nand U505 (N_505,N_227,N_232);
or U506 (N_506,N_222,N_60);
nand U507 (N_507,In_548,In_810);
nand U508 (N_508,N_135,In_749);
and U509 (N_509,In_790,In_89);
or U510 (N_510,N_300,N_286);
nand U511 (N_511,N_309,N_237);
and U512 (N_512,In_907,In_505);
nor U513 (N_513,N_324,In_448);
xnor U514 (N_514,In_219,In_200);
nor U515 (N_515,In_468,In_668);
nand U516 (N_516,In_74,In_764);
nor U517 (N_517,N_374,In_592);
and U518 (N_518,N_69,N_251);
nand U519 (N_519,In_630,N_230);
xor U520 (N_520,N_277,N_330);
and U521 (N_521,N_136,In_51);
nor U522 (N_522,In_538,In_197);
nor U523 (N_523,N_81,In_942);
nand U524 (N_524,N_336,N_343);
xnor U525 (N_525,N_35,N_270);
xnor U526 (N_526,N_348,In_870);
and U527 (N_527,In_800,N_294);
and U528 (N_528,N_213,N_77);
and U529 (N_529,In_702,In_845);
or U530 (N_530,N_123,N_328);
and U531 (N_531,In_727,N_228);
nor U532 (N_532,N_63,In_556);
nand U533 (N_533,In_984,In_93);
xnor U534 (N_534,N_207,In_564);
nand U535 (N_535,N_332,N_195);
and U536 (N_536,N_284,In_67);
nor U537 (N_537,N_205,In_731);
xor U538 (N_538,N_84,N_296);
or U539 (N_539,In_446,In_420);
or U540 (N_540,In_952,N_214);
xor U541 (N_541,N_18,In_506);
nor U542 (N_542,N_154,In_999);
or U543 (N_543,N_151,In_927);
nor U544 (N_544,N_319,N_275);
and U545 (N_545,In_896,In_77);
nand U546 (N_546,In_159,N_365);
nor U547 (N_547,N_298,N_337);
or U548 (N_548,In_926,N_92);
xor U549 (N_549,N_52,In_38);
or U550 (N_550,In_822,N_158);
nand U551 (N_551,N_386,In_188);
nor U552 (N_552,N_295,In_24);
and U553 (N_553,In_794,N_171);
and U554 (N_554,In_264,In_851);
nor U555 (N_555,In_933,N_327);
nor U556 (N_556,In_292,In_698);
nand U557 (N_557,In_958,N_142);
or U558 (N_558,In_752,In_56);
nand U559 (N_559,In_826,N_395);
nor U560 (N_560,N_375,N_233);
nor U561 (N_561,N_196,In_612);
and U562 (N_562,In_378,In_20);
xnor U563 (N_563,In_398,N_132);
or U564 (N_564,N_121,N_384);
and U565 (N_565,In_853,N_99);
xnor U566 (N_566,N_19,In_776);
nor U567 (N_567,N_351,In_125);
and U568 (N_568,In_287,In_304);
nand U569 (N_569,N_345,N_326);
nand U570 (N_570,N_302,In_152);
nor U571 (N_571,N_253,N_267);
and U572 (N_572,In_452,In_690);
nor U573 (N_573,N_240,In_772);
nor U574 (N_574,N_14,In_58);
nand U575 (N_575,In_342,In_620);
or U576 (N_576,In_480,N_371);
or U577 (N_577,N_322,N_210);
xor U578 (N_578,N_183,In_559);
or U579 (N_579,N_352,N_104);
nand U580 (N_580,N_129,N_264);
nand U581 (N_581,In_259,N_310);
nor U582 (N_582,N_364,N_226);
xor U583 (N_583,N_201,N_361);
nor U584 (N_584,In_697,N_379);
and U585 (N_585,In_584,N_362);
nand U586 (N_586,In_395,N_354);
or U587 (N_587,N_48,N_274);
nand U588 (N_588,N_367,In_276);
and U589 (N_589,In_511,In_741);
nand U590 (N_590,In_142,In_343);
nor U591 (N_591,N_26,In_476);
nand U592 (N_592,In_754,In_440);
and U593 (N_593,N_396,N_212);
and U594 (N_594,N_388,In_799);
nor U595 (N_595,N_263,N_211);
or U596 (N_596,In_805,N_22);
nand U597 (N_597,In_677,In_659);
xor U598 (N_598,In_639,In_362);
or U599 (N_599,N_359,In_849);
or U600 (N_600,N_353,N_408);
and U601 (N_601,N_554,N_287);
nor U602 (N_602,N_439,N_590);
nor U603 (N_603,N_443,N_555);
nor U604 (N_604,In_281,N_533);
xor U605 (N_605,N_547,N_358);
and U606 (N_606,In_652,N_257);
nor U607 (N_607,In_55,N_561);
and U608 (N_608,N_280,N_209);
xnor U609 (N_609,In_877,N_447);
and U610 (N_610,N_417,N_544);
and U611 (N_611,In_950,N_534);
nor U612 (N_612,N_517,In_127);
xnor U613 (N_613,N_575,N_425);
xnor U614 (N_614,N_145,In_635);
or U615 (N_615,N_289,N_402);
nor U616 (N_616,N_82,N_373);
nand U617 (N_617,In_9,N_557);
nand U618 (N_618,N_475,In_131);
nand U619 (N_619,N_355,N_470);
xor U620 (N_620,N_520,N_469);
nand U621 (N_621,N_398,In_341);
and U622 (N_622,N_492,N_482);
or U623 (N_623,N_483,N_452);
and U624 (N_624,N_255,In_693);
xor U625 (N_625,N_487,In_911);
nor U626 (N_626,In_339,N_428);
and U627 (N_627,N_465,N_499);
nor U628 (N_628,In_6,In_401);
nor U629 (N_629,N_537,N_460);
or U630 (N_630,N_392,N_559);
nand U631 (N_631,N_574,N_558);
nand U632 (N_632,N_66,In_599);
or U633 (N_633,N_377,In_265);
or U634 (N_634,N_496,N_510);
nor U635 (N_635,In_571,N_479);
nor U636 (N_636,N_426,In_465);
and U637 (N_637,N_540,N_329);
xnor U638 (N_638,N_518,N_440);
or U639 (N_639,In_930,N_504);
xor U640 (N_640,N_144,N_187);
nand U641 (N_641,N_317,N_568);
xor U642 (N_642,In_634,N_174);
nor U643 (N_643,N_515,In_979);
nor U644 (N_644,In_275,N_258);
or U645 (N_645,N_578,N_404);
and U646 (N_646,N_170,N_491);
or U647 (N_647,N_88,In_460);
xnor U648 (N_648,N_306,N_261);
nand U649 (N_649,N_197,N_391);
or U650 (N_650,N_340,N_273);
nor U651 (N_651,In_714,N_591);
nand U652 (N_652,N_532,In_781);
and U653 (N_653,N_37,In_733);
xnor U654 (N_654,N_250,In_90);
nand U655 (N_655,N_586,N_594);
nand U656 (N_656,In_40,N_543);
or U657 (N_657,N_509,In_699);
and U658 (N_658,N_418,N_441);
and U659 (N_659,N_138,N_98);
xnor U660 (N_660,N_87,N_334);
nor U661 (N_661,N_454,N_477);
xnor U662 (N_662,N_372,In_76);
and U663 (N_663,N_463,N_299);
or U664 (N_664,N_83,N_456);
and U665 (N_665,N_505,N_437);
and U666 (N_666,In_377,In_289);
nand U667 (N_667,N_525,N_503);
nor U668 (N_668,N_67,N_589);
nor U669 (N_669,In_739,N_451);
or U670 (N_670,N_256,N_581);
or U671 (N_671,N_73,N_432);
or U672 (N_672,N_522,N_421);
xnor U673 (N_673,N_342,N_216);
and U674 (N_674,N_412,N_523);
nor U675 (N_675,In_68,N_41);
and U676 (N_676,N_401,In_355);
xnor U677 (N_677,N_560,N_419);
nand U678 (N_678,N_573,N_153);
nor U679 (N_679,N_597,N_405);
nor U680 (N_680,N_242,N_599);
and U681 (N_681,N_536,N_363);
or U682 (N_682,N_55,N_450);
or U683 (N_683,N_203,N_24);
nand U684 (N_684,N_580,In_431);
nor U685 (N_685,N_307,N_472);
xnor U686 (N_686,N_276,N_549);
xnor U687 (N_687,N_218,N_118);
nand U688 (N_688,In_46,In_759);
nor U689 (N_689,N_446,In_199);
xor U690 (N_690,N_508,N_435);
nand U691 (N_691,N_423,In_81);
nor U692 (N_692,In_270,N_464);
nand U693 (N_693,N_445,N_223);
and U694 (N_694,In_399,In_654);
and U695 (N_695,In_525,N_436);
nand U696 (N_696,N_596,N_473);
xnor U697 (N_697,N_94,In_836);
xnor U698 (N_698,N_119,N_502);
and U699 (N_699,N_314,N_164);
nor U700 (N_700,N_511,N_556);
nand U701 (N_701,In_365,In_928);
nor U702 (N_702,N_498,N_414);
nor U703 (N_703,N_572,In_212);
xor U704 (N_704,N_427,N_304);
xnor U705 (N_705,N_565,N_521);
nand U706 (N_706,N_474,N_430);
nor U707 (N_707,N_507,N_481);
and U708 (N_708,In_626,N_252);
nor U709 (N_709,In_213,In_701);
nand U710 (N_710,N_512,N_527);
nor U711 (N_711,In_674,N_113);
or U712 (N_712,N_553,In_444);
nor U713 (N_713,N_291,N_468);
nand U714 (N_714,N_5,N_308);
and U715 (N_715,N_514,In_590);
or U716 (N_716,N_494,N_366);
or U717 (N_717,N_429,N_587);
or U718 (N_718,N_434,In_513);
and U719 (N_719,N_459,N_592);
nand U720 (N_720,In_162,In_488);
xor U721 (N_721,In_215,N_476);
or U722 (N_722,N_415,In_192);
or U723 (N_723,In_351,N_431);
nor U724 (N_724,N_397,N_115);
and U725 (N_725,N_466,N_449);
or U726 (N_726,In_658,N_551);
or U727 (N_727,In_672,N_531);
nand U728 (N_728,N_562,N_569);
xor U729 (N_729,In_236,In_291);
nand U730 (N_730,In_932,N_486);
nor U731 (N_731,In_368,N_155);
nor U732 (N_732,N_566,N_576);
or U733 (N_733,In_686,N_192);
nand U734 (N_734,N_598,N_538);
xnor U735 (N_735,N_16,In_322);
nand U736 (N_736,N_528,N_563);
xor U737 (N_737,N_485,In_558);
nand U738 (N_738,N_410,N_541);
nand U739 (N_739,N_148,N_501);
and U740 (N_740,N_101,N_325);
xnor U741 (N_741,N_539,N_265);
nor U742 (N_742,N_519,In_848);
and U743 (N_743,N_457,In_554);
nand U744 (N_744,N_283,N_341);
nand U745 (N_745,N_292,N_461);
xnor U746 (N_746,In_994,N_546);
and U747 (N_747,N_110,N_467);
xnor U748 (N_748,In_650,N_584);
nor U749 (N_749,N_407,N_455);
or U750 (N_750,N_356,N_593);
or U751 (N_751,N_550,N_478);
xnor U752 (N_752,N_500,In_841);
nor U753 (N_753,In_789,In_642);
nand U754 (N_754,N_583,N_570);
and U755 (N_755,N_582,N_390);
xor U756 (N_756,N_378,N_524);
or U757 (N_757,N_346,N_585);
nand U758 (N_758,N_39,N_204);
nand U759 (N_759,In_941,In_653);
nand U760 (N_760,N_413,N_381);
nand U761 (N_761,N_493,N_433);
nor U762 (N_762,N_416,In_82);
nand U763 (N_763,N_424,In_101);
nor U764 (N_764,In_305,N_488);
nand U765 (N_765,N_529,N_93);
and U766 (N_766,N_403,In_340);
nor U767 (N_767,N_134,In_796);
or U768 (N_768,N_178,In_798);
and U769 (N_769,N_462,N_438);
xor U770 (N_770,N_571,In_718);
nand U771 (N_771,N_420,N_484);
nand U772 (N_772,N_167,N_448);
and U773 (N_773,N_490,N_143);
and U774 (N_774,In_205,N_453);
nor U775 (N_775,N_411,N_506);
or U776 (N_776,N_444,In_549);
xor U777 (N_777,N_564,In_57);
xor U778 (N_778,N_516,In_502);
or U779 (N_779,N_480,N_545);
and U780 (N_780,In_350,N_535);
xnor U781 (N_781,N_331,N_394);
and U782 (N_782,N_11,N_595);
and U783 (N_783,In_416,N_139);
or U784 (N_784,In_389,N_409);
nor U785 (N_785,In_388,N_335);
or U786 (N_786,N_489,N_567);
nor U787 (N_787,In_216,N_579);
or U788 (N_788,N_552,N_588);
and U789 (N_789,N_422,N_316);
nand U790 (N_790,In_777,N_141);
xnor U791 (N_791,N_400,N_513);
or U792 (N_792,In_785,N_323);
nand U793 (N_793,N_406,N_497);
or U794 (N_794,N_458,N_542);
or U795 (N_795,N_530,N_471);
and U796 (N_796,In_946,N_442);
xnor U797 (N_797,N_577,N_495);
and U798 (N_798,N_548,In_966);
and U799 (N_799,N_146,N_526);
nor U800 (N_800,N_684,N_689);
nand U801 (N_801,N_773,N_612);
or U802 (N_802,N_710,N_696);
nand U803 (N_803,N_775,N_691);
or U804 (N_804,N_789,N_704);
or U805 (N_805,N_651,N_607);
or U806 (N_806,N_660,N_767);
and U807 (N_807,N_796,N_698);
nand U808 (N_808,N_749,N_680);
and U809 (N_809,N_735,N_601);
nor U810 (N_810,N_793,N_643);
nand U811 (N_811,N_711,N_746);
nand U812 (N_812,N_731,N_743);
nand U813 (N_813,N_633,N_645);
nand U814 (N_814,N_752,N_699);
and U815 (N_815,N_730,N_750);
nand U816 (N_816,N_609,N_715);
nor U817 (N_817,N_656,N_611);
nand U818 (N_818,N_799,N_785);
xnor U819 (N_819,N_650,N_676);
xnor U820 (N_820,N_622,N_700);
and U821 (N_821,N_687,N_638);
nor U822 (N_822,N_641,N_602);
or U823 (N_823,N_690,N_647);
xor U824 (N_824,N_794,N_774);
nand U825 (N_825,N_778,N_702);
and U826 (N_826,N_649,N_631);
and U827 (N_827,N_624,N_619);
and U828 (N_828,N_783,N_616);
nand U829 (N_829,N_717,N_606);
and U830 (N_830,N_629,N_714);
or U831 (N_831,N_781,N_639);
nand U832 (N_832,N_666,N_719);
nor U833 (N_833,N_608,N_720);
xor U834 (N_834,N_748,N_603);
and U835 (N_835,N_644,N_692);
and U836 (N_836,N_669,N_784);
or U837 (N_837,N_621,N_701);
xnor U838 (N_838,N_740,N_628);
xor U839 (N_839,N_635,N_663);
nor U840 (N_840,N_648,N_758);
and U841 (N_841,N_797,N_705);
xnor U842 (N_842,N_664,N_665);
or U843 (N_843,N_770,N_654);
nand U844 (N_844,N_625,N_737);
xor U845 (N_845,N_792,N_718);
xnor U846 (N_846,N_615,N_780);
or U847 (N_847,N_769,N_693);
and U848 (N_848,N_766,N_779);
and U849 (N_849,N_655,N_677);
or U850 (N_850,N_726,N_617);
nand U851 (N_851,N_642,N_653);
xor U852 (N_852,N_682,N_678);
nand U853 (N_853,N_672,N_632);
or U854 (N_854,N_753,N_754);
and U855 (N_855,N_600,N_728);
and U856 (N_856,N_636,N_686);
xor U857 (N_857,N_736,N_791);
xnor U858 (N_858,N_661,N_685);
nor U859 (N_859,N_733,N_721);
or U860 (N_860,N_659,N_763);
nor U861 (N_861,N_623,N_755);
nand U862 (N_862,N_634,N_742);
or U863 (N_863,N_673,N_662);
nor U864 (N_864,N_637,N_681);
or U865 (N_865,N_729,N_688);
nor U866 (N_866,N_786,N_762);
nor U867 (N_867,N_798,N_725);
xor U868 (N_868,N_670,N_658);
nor U869 (N_869,N_695,N_765);
or U870 (N_870,N_795,N_747);
or U871 (N_871,N_759,N_723);
or U872 (N_872,N_613,N_761);
nor U873 (N_873,N_620,N_652);
xor U874 (N_874,N_777,N_734);
or U875 (N_875,N_716,N_614);
nand U876 (N_876,N_744,N_604);
or U877 (N_877,N_757,N_703);
nand U878 (N_878,N_668,N_712);
or U879 (N_879,N_630,N_709);
xor U880 (N_880,N_768,N_671);
xnor U881 (N_881,N_707,N_787);
and U882 (N_882,N_618,N_745);
nand U883 (N_883,N_640,N_605);
and U884 (N_884,N_741,N_708);
or U885 (N_885,N_756,N_732);
xor U886 (N_886,N_739,N_724);
xnor U887 (N_887,N_760,N_610);
and U888 (N_888,N_706,N_738);
or U889 (N_889,N_771,N_679);
and U890 (N_890,N_790,N_722);
nand U891 (N_891,N_788,N_646);
xnor U892 (N_892,N_776,N_697);
nor U893 (N_893,N_627,N_667);
and U894 (N_894,N_727,N_683);
nor U895 (N_895,N_713,N_764);
and U896 (N_896,N_626,N_657);
nand U897 (N_897,N_694,N_772);
nand U898 (N_898,N_675,N_751);
and U899 (N_899,N_782,N_674);
xor U900 (N_900,N_762,N_601);
nor U901 (N_901,N_676,N_748);
nand U902 (N_902,N_778,N_631);
xnor U903 (N_903,N_638,N_798);
and U904 (N_904,N_708,N_798);
or U905 (N_905,N_692,N_618);
and U906 (N_906,N_676,N_651);
and U907 (N_907,N_705,N_642);
xnor U908 (N_908,N_609,N_683);
or U909 (N_909,N_739,N_781);
or U910 (N_910,N_699,N_764);
and U911 (N_911,N_701,N_772);
nor U912 (N_912,N_799,N_724);
and U913 (N_913,N_620,N_637);
and U914 (N_914,N_786,N_770);
xor U915 (N_915,N_622,N_767);
nor U916 (N_916,N_619,N_780);
and U917 (N_917,N_672,N_757);
xor U918 (N_918,N_754,N_711);
nand U919 (N_919,N_723,N_664);
or U920 (N_920,N_700,N_621);
or U921 (N_921,N_770,N_695);
xor U922 (N_922,N_683,N_687);
and U923 (N_923,N_779,N_616);
xor U924 (N_924,N_630,N_615);
or U925 (N_925,N_717,N_673);
nor U926 (N_926,N_788,N_737);
nor U927 (N_927,N_734,N_623);
nor U928 (N_928,N_772,N_605);
nand U929 (N_929,N_631,N_766);
or U930 (N_930,N_637,N_645);
nand U931 (N_931,N_664,N_623);
and U932 (N_932,N_735,N_771);
nor U933 (N_933,N_704,N_781);
nand U934 (N_934,N_682,N_677);
and U935 (N_935,N_694,N_689);
or U936 (N_936,N_736,N_604);
or U937 (N_937,N_673,N_609);
nand U938 (N_938,N_605,N_793);
nor U939 (N_939,N_750,N_741);
nor U940 (N_940,N_634,N_790);
and U941 (N_941,N_605,N_737);
xnor U942 (N_942,N_634,N_757);
nor U943 (N_943,N_623,N_768);
xor U944 (N_944,N_735,N_738);
and U945 (N_945,N_641,N_646);
nand U946 (N_946,N_652,N_794);
or U947 (N_947,N_771,N_745);
xor U948 (N_948,N_788,N_630);
nand U949 (N_949,N_747,N_760);
or U950 (N_950,N_645,N_666);
nand U951 (N_951,N_687,N_787);
and U952 (N_952,N_663,N_690);
and U953 (N_953,N_627,N_689);
nand U954 (N_954,N_755,N_626);
and U955 (N_955,N_611,N_771);
nor U956 (N_956,N_663,N_795);
nor U957 (N_957,N_718,N_747);
nand U958 (N_958,N_709,N_673);
or U959 (N_959,N_749,N_662);
nand U960 (N_960,N_742,N_694);
and U961 (N_961,N_796,N_787);
xor U962 (N_962,N_689,N_695);
xor U963 (N_963,N_605,N_773);
or U964 (N_964,N_743,N_753);
and U965 (N_965,N_794,N_666);
nor U966 (N_966,N_779,N_621);
and U967 (N_967,N_760,N_797);
or U968 (N_968,N_723,N_666);
nand U969 (N_969,N_624,N_693);
xor U970 (N_970,N_717,N_707);
xnor U971 (N_971,N_718,N_737);
nor U972 (N_972,N_645,N_733);
and U973 (N_973,N_658,N_728);
nand U974 (N_974,N_675,N_636);
xnor U975 (N_975,N_661,N_626);
or U976 (N_976,N_684,N_711);
nor U977 (N_977,N_678,N_763);
nor U978 (N_978,N_653,N_639);
or U979 (N_979,N_683,N_647);
xor U980 (N_980,N_744,N_703);
xor U981 (N_981,N_711,N_610);
xor U982 (N_982,N_706,N_715);
nor U983 (N_983,N_722,N_712);
xor U984 (N_984,N_735,N_741);
or U985 (N_985,N_720,N_684);
or U986 (N_986,N_630,N_731);
xnor U987 (N_987,N_789,N_769);
or U988 (N_988,N_794,N_676);
and U989 (N_989,N_767,N_699);
or U990 (N_990,N_698,N_677);
or U991 (N_991,N_714,N_672);
and U992 (N_992,N_756,N_679);
and U993 (N_993,N_720,N_671);
nor U994 (N_994,N_610,N_665);
and U995 (N_995,N_693,N_755);
or U996 (N_996,N_732,N_641);
or U997 (N_997,N_604,N_773);
nand U998 (N_998,N_662,N_702);
nor U999 (N_999,N_736,N_793);
or U1000 (N_1000,N_952,N_930);
and U1001 (N_1001,N_812,N_977);
nor U1002 (N_1002,N_859,N_971);
or U1003 (N_1003,N_996,N_988);
nor U1004 (N_1004,N_913,N_808);
or U1005 (N_1005,N_824,N_850);
nor U1006 (N_1006,N_845,N_816);
and U1007 (N_1007,N_833,N_828);
xnor U1008 (N_1008,N_964,N_814);
nand U1009 (N_1009,N_836,N_928);
nor U1010 (N_1010,N_938,N_980);
xnor U1011 (N_1011,N_869,N_831);
xor U1012 (N_1012,N_901,N_925);
and U1013 (N_1013,N_851,N_888);
and U1014 (N_1014,N_872,N_982);
nor U1015 (N_1015,N_835,N_852);
or U1016 (N_1016,N_960,N_847);
nand U1017 (N_1017,N_923,N_909);
nand U1018 (N_1018,N_896,N_922);
and U1019 (N_1019,N_946,N_939);
or U1020 (N_1020,N_951,N_958);
and U1021 (N_1021,N_968,N_804);
or U1022 (N_1022,N_815,N_955);
nor U1023 (N_1023,N_947,N_953);
or U1024 (N_1024,N_825,N_881);
and U1025 (N_1025,N_983,N_967);
or U1026 (N_1026,N_999,N_877);
nand U1027 (N_1027,N_826,N_878);
xnor U1028 (N_1028,N_853,N_935);
and U1029 (N_1029,N_990,N_843);
xnor U1030 (N_1030,N_823,N_950);
xor U1031 (N_1031,N_864,N_854);
and U1032 (N_1032,N_921,N_918);
nand U1033 (N_1033,N_856,N_803);
and U1034 (N_1034,N_897,N_956);
nand U1035 (N_1035,N_801,N_885);
or U1036 (N_1036,N_855,N_972);
and U1037 (N_1037,N_842,N_933);
nand U1038 (N_1038,N_929,N_916);
or U1039 (N_1039,N_893,N_883);
nand U1040 (N_1040,N_811,N_873);
and U1041 (N_1041,N_817,N_906);
and U1042 (N_1042,N_800,N_900);
nand U1043 (N_1043,N_832,N_805);
or U1044 (N_1044,N_992,N_862);
or U1045 (N_1045,N_818,N_895);
nand U1046 (N_1046,N_807,N_834);
and U1047 (N_1047,N_910,N_932);
and U1048 (N_1048,N_827,N_905);
or U1049 (N_1049,N_974,N_844);
nand U1050 (N_1050,N_802,N_995);
nand U1051 (N_1051,N_865,N_927);
or U1052 (N_1052,N_970,N_886);
nor U1053 (N_1053,N_991,N_945);
nor U1054 (N_1054,N_941,N_839);
and U1055 (N_1055,N_959,N_907);
and U1056 (N_1056,N_966,N_963);
or U1057 (N_1057,N_860,N_838);
or U1058 (N_1058,N_940,N_849);
nor U1059 (N_1059,N_870,N_961);
xnor U1060 (N_1060,N_846,N_949);
nor U1061 (N_1061,N_908,N_861);
nor U1062 (N_1062,N_943,N_965);
xnor U1063 (N_1063,N_858,N_934);
and U1064 (N_1064,N_978,N_898);
or U1065 (N_1065,N_942,N_868);
nand U1066 (N_1066,N_890,N_819);
nand U1067 (N_1067,N_954,N_924);
xor U1068 (N_1068,N_903,N_882);
nand U1069 (N_1069,N_830,N_911);
nand U1070 (N_1070,N_944,N_936);
or U1071 (N_1071,N_998,N_919);
nor U1072 (N_1072,N_857,N_871);
nand U1073 (N_1073,N_985,N_987);
or U1074 (N_1074,N_889,N_874);
nand U1075 (N_1075,N_829,N_904);
and U1076 (N_1076,N_979,N_867);
nor U1077 (N_1077,N_822,N_891);
nor U1078 (N_1078,N_813,N_899);
nand U1079 (N_1079,N_969,N_820);
nand U1080 (N_1080,N_806,N_986);
or U1081 (N_1081,N_984,N_841);
xnor U1082 (N_1082,N_894,N_976);
or U1083 (N_1083,N_848,N_821);
or U1084 (N_1084,N_957,N_997);
and U1085 (N_1085,N_937,N_837);
nor U1086 (N_1086,N_914,N_880);
xor U1087 (N_1087,N_926,N_981);
or U1088 (N_1088,N_875,N_879);
and U1089 (N_1089,N_915,N_912);
and U1090 (N_1090,N_810,N_863);
nand U1091 (N_1091,N_917,N_884);
xnor U1092 (N_1092,N_948,N_887);
and U1093 (N_1093,N_994,N_809);
and U1094 (N_1094,N_892,N_973);
and U1095 (N_1095,N_962,N_975);
or U1096 (N_1096,N_989,N_902);
nor U1097 (N_1097,N_931,N_920);
nand U1098 (N_1098,N_876,N_993);
and U1099 (N_1099,N_840,N_866);
nand U1100 (N_1100,N_808,N_833);
or U1101 (N_1101,N_962,N_898);
nand U1102 (N_1102,N_861,N_827);
nand U1103 (N_1103,N_983,N_856);
nor U1104 (N_1104,N_954,N_875);
and U1105 (N_1105,N_879,N_898);
nand U1106 (N_1106,N_918,N_986);
nand U1107 (N_1107,N_887,N_822);
nor U1108 (N_1108,N_827,N_838);
nor U1109 (N_1109,N_813,N_917);
nand U1110 (N_1110,N_995,N_968);
nor U1111 (N_1111,N_899,N_860);
nand U1112 (N_1112,N_811,N_819);
and U1113 (N_1113,N_933,N_937);
or U1114 (N_1114,N_858,N_810);
and U1115 (N_1115,N_857,N_854);
or U1116 (N_1116,N_920,N_944);
nand U1117 (N_1117,N_869,N_903);
and U1118 (N_1118,N_912,N_980);
nor U1119 (N_1119,N_910,N_865);
and U1120 (N_1120,N_858,N_930);
nand U1121 (N_1121,N_918,N_893);
nand U1122 (N_1122,N_925,N_883);
and U1123 (N_1123,N_865,N_997);
xnor U1124 (N_1124,N_817,N_909);
xnor U1125 (N_1125,N_904,N_834);
and U1126 (N_1126,N_884,N_895);
or U1127 (N_1127,N_830,N_886);
xnor U1128 (N_1128,N_840,N_996);
nor U1129 (N_1129,N_832,N_851);
xnor U1130 (N_1130,N_991,N_960);
or U1131 (N_1131,N_801,N_977);
nand U1132 (N_1132,N_897,N_953);
or U1133 (N_1133,N_922,N_910);
or U1134 (N_1134,N_984,N_825);
or U1135 (N_1135,N_990,N_888);
and U1136 (N_1136,N_969,N_998);
nand U1137 (N_1137,N_832,N_906);
or U1138 (N_1138,N_976,N_828);
nand U1139 (N_1139,N_827,N_959);
and U1140 (N_1140,N_852,N_904);
or U1141 (N_1141,N_919,N_904);
or U1142 (N_1142,N_810,N_883);
and U1143 (N_1143,N_850,N_902);
nand U1144 (N_1144,N_912,N_923);
and U1145 (N_1145,N_869,N_853);
nor U1146 (N_1146,N_958,N_991);
or U1147 (N_1147,N_877,N_894);
nor U1148 (N_1148,N_905,N_967);
nor U1149 (N_1149,N_890,N_853);
and U1150 (N_1150,N_974,N_878);
or U1151 (N_1151,N_934,N_925);
or U1152 (N_1152,N_990,N_864);
xor U1153 (N_1153,N_880,N_984);
xnor U1154 (N_1154,N_902,N_974);
or U1155 (N_1155,N_908,N_961);
nor U1156 (N_1156,N_835,N_830);
nand U1157 (N_1157,N_906,N_931);
and U1158 (N_1158,N_992,N_964);
nand U1159 (N_1159,N_831,N_922);
xnor U1160 (N_1160,N_843,N_945);
and U1161 (N_1161,N_925,N_958);
nor U1162 (N_1162,N_921,N_947);
nand U1163 (N_1163,N_965,N_893);
and U1164 (N_1164,N_818,N_998);
xor U1165 (N_1165,N_886,N_993);
xor U1166 (N_1166,N_958,N_843);
nor U1167 (N_1167,N_976,N_844);
xnor U1168 (N_1168,N_968,N_908);
nor U1169 (N_1169,N_918,N_929);
xnor U1170 (N_1170,N_861,N_921);
or U1171 (N_1171,N_800,N_954);
nand U1172 (N_1172,N_897,N_890);
and U1173 (N_1173,N_837,N_968);
nor U1174 (N_1174,N_840,N_991);
and U1175 (N_1175,N_902,N_837);
or U1176 (N_1176,N_839,N_824);
xor U1177 (N_1177,N_933,N_847);
nand U1178 (N_1178,N_995,N_874);
xor U1179 (N_1179,N_907,N_958);
nor U1180 (N_1180,N_855,N_964);
nand U1181 (N_1181,N_951,N_803);
or U1182 (N_1182,N_838,N_813);
nand U1183 (N_1183,N_956,N_996);
xnor U1184 (N_1184,N_976,N_888);
nand U1185 (N_1185,N_997,N_871);
or U1186 (N_1186,N_868,N_979);
xor U1187 (N_1187,N_983,N_990);
xnor U1188 (N_1188,N_974,N_912);
nor U1189 (N_1189,N_973,N_825);
or U1190 (N_1190,N_970,N_867);
nor U1191 (N_1191,N_928,N_857);
xnor U1192 (N_1192,N_886,N_831);
and U1193 (N_1193,N_893,N_845);
nor U1194 (N_1194,N_880,N_876);
or U1195 (N_1195,N_938,N_880);
nand U1196 (N_1196,N_879,N_844);
nor U1197 (N_1197,N_965,N_835);
nor U1198 (N_1198,N_919,N_808);
or U1199 (N_1199,N_903,N_846);
or U1200 (N_1200,N_1195,N_1160);
nand U1201 (N_1201,N_1024,N_1083);
xor U1202 (N_1202,N_1091,N_1162);
and U1203 (N_1203,N_1165,N_1025);
nor U1204 (N_1204,N_1168,N_1075);
and U1205 (N_1205,N_1046,N_1177);
or U1206 (N_1206,N_1108,N_1153);
and U1207 (N_1207,N_1131,N_1064);
nor U1208 (N_1208,N_1088,N_1019);
and U1209 (N_1209,N_1065,N_1134);
xnor U1210 (N_1210,N_1185,N_1102);
nand U1211 (N_1211,N_1032,N_1147);
and U1212 (N_1212,N_1186,N_1066);
nand U1213 (N_1213,N_1192,N_1179);
and U1214 (N_1214,N_1116,N_1123);
xor U1215 (N_1215,N_1174,N_1144);
nand U1216 (N_1216,N_1048,N_1181);
xnor U1217 (N_1217,N_1073,N_1127);
and U1218 (N_1218,N_1107,N_1000);
or U1219 (N_1219,N_1189,N_1047);
or U1220 (N_1220,N_1051,N_1169);
xnor U1221 (N_1221,N_1035,N_1054);
and U1222 (N_1222,N_1038,N_1062);
nor U1223 (N_1223,N_1059,N_1037);
nand U1224 (N_1224,N_1045,N_1060);
nor U1225 (N_1225,N_1175,N_1128);
and U1226 (N_1226,N_1005,N_1004);
xnor U1227 (N_1227,N_1133,N_1136);
and U1228 (N_1228,N_1158,N_1104);
or U1229 (N_1229,N_1125,N_1145);
and U1230 (N_1230,N_1183,N_1089);
nor U1231 (N_1231,N_1092,N_1018);
and U1232 (N_1232,N_1101,N_1085);
and U1233 (N_1233,N_1132,N_1188);
xor U1234 (N_1234,N_1042,N_1034);
xor U1235 (N_1235,N_1002,N_1022);
xor U1236 (N_1236,N_1167,N_1187);
nand U1237 (N_1237,N_1033,N_1198);
and U1238 (N_1238,N_1040,N_1070);
nor U1239 (N_1239,N_1090,N_1171);
xnor U1240 (N_1240,N_1163,N_1084);
or U1241 (N_1241,N_1079,N_1093);
nand U1242 (N_1242,N_1098,N_1067);
and U1243 (N_1243,N_1043,N_1159);
or U1244 (N_1244,N_1056,N_1013);
nand U1245 (N_1245,N_1191,N_1021);
nor U1246 (N_1246,N_1112,N_1126);
or U1247 (N_1247,N_1055,N_1197);
nor U1248 (N_1248,N_1053,N_1016);
and U1249 (N_1249,N_1069,N_1026);
xor U1250 (N_1250,N_1003,N_1182);
or U1251 (N_1251,N_1148,N_1029);
nor U1252 (N_1252,N_1041,N_1078);
and U1253 (N_1253,N_1050,N_1155);
xor U1254 (N_1254,N_1120,N_1149);
nand U1255 (N_1255,N_1130,N_1086);
nand U1256 (N_1256,N_1012,N_1142);
nand U1257 (N_1257,N_1199,N_1170);
nand U1258 (N_1258,N_1010,N_1173);
nand U1259 (N_1259,N_1063,N_1166);
or U1260 (N_1260,N_1014,N_1193);
nand U1261 (N_1261,N_1015,N_1156);
nand U1262 (N_1262,N_1190,N_1039);
and U1263 (N_1263,N_1007,N_1082);
nor U1264 (N_1264,N_1184,N_1139);
nor U1265 (N_1265,N_1140,N_1194);
nand U1266 (N_1266,N_1076,N_1049);
and U1267 (N_1267,N_1157,N_1097);
nand U1268 (N_1268,N_1110,N_1103);
nand U1269 (N_1269,N_1137,N_1017);
and U1270 (N_1270,N_1172,N_1146);
xnor U1271 (N_1271,N_1057,N_1109);
or U1272 (N_1272,N_1122,N_1028);
nand U1273 (N_1273,N_1121,N_1052);
xor U1274 (N_1274,N_1113,N_1176);
xor U1275 (N_1275,N_1058,N_1099);
nor U1276 (N_1276,N_1068,N_1023);
nand U1277 (N_1277,N_1020,N_1080);
nand U1278 (N_1278,N_1071,N_1027);
nand U1279 (N_1279,N_1154,N_1164);
and U1280 (N_1280,N_1129,N_1150);
nand U1281 (N_1281,N_1115,N_1178);
nor U1282 (N_1282,N_1106,N_1036);
and U1283 (N_1283,N_1124,N_1119);
or U1284 (N_1284,N_1105,N_1096);
nand U1285 (N_1285,N_1143,N_1152);
nand U1286 (N_1286,N_1072,N_1094);
and U1287 (N_1287,N_1151,N_1117);
and U1288 (N_1288,N_1031,N_1138);
xnor U1289 (N_1289,N_1074,N_1081);
nand U1290 (N_1290,N_1111,N_1077);
nand U1291 (N_1291,N_1135,N_1196);
xnor U1292 (N_1292,N_1100,N_1006);
and U1293 (N_1293,N_1011,N_1061);
and U1294 (N_1294,N_1008,N_1009);
or U1295 (N_1295,N_1141,N_1095);
or U1296 (N_1296,N_1114,N_1087);
xnor U1297 (N_1297,N_1118,N_1044);
nor U1298 (N_1298,N_1001,N_1180);
nor U1299 (N_1299,N_1161,N_1030);
xor U1300 (N_1300,N_1112,N_1019);
nand U1301 (N_1301,N_1111,N_1106);
and U1302 (N_1302,N_1053,N_1022);
or U1303 (N_1303,N_1191,N_1135);
nor U1304 (N_1304,N_1196,N_1088);
and U1305 (N_1305,N_1164,N_1121);
nor U1306 (N_1306,N_1057,N_1084);
nor U1307 (N_1307,N_1126,N_1132);
nor U1308 (N_1308,N_1127,N_1062);
xnor U1309 (N_1309,N_1090,N_1168);
xor U1310 (N_1310,N_1012,N_1147);
nor U1311 (N_1311,N_1134,N_1151);
and U1312 (N_1312,N_1120,N_1099);
or U1313 (N_1313,N_1014,N_1015);
or U1314 (N_1314,N_1177,N_1112);
nand U1315 (N_1315,N_1163,N_1177);
nand U1316 (N_1316,N_1103,N_1115);
xor U1317 (N_1317,N_1093,N_1090);
xnor U1318 (N_1318,N_1091,N_1098);
xor U1319 (N_1319,N_1145,N_1191);
or U1320 (N_1320,N_1008,N_1021);
nor U1321 (N_1321,N_1144,N_1044);
xor U1322 (N_1322,N_1197,N_1139);
or U1323 (N_1323,N_1036,N_1152);
and U1324 (N_1324,N_1006,N_1013);
nor U1325 (N_1325,N_1143,N_1066);
and U1326 (N_1326,N_1070,N_1186);
xor U1327 (N_1327,N_1100,N_1008);
xnor U1328 (N_1328,N_1076,N_1124);
xnor U1329 (N_1329,N_1019,N_1169);
and U1330 (N_1330,N_1161,N_1141);
and U1331 (N_1331,N_1037,N_1024);
nor U1332 (N_1332,N_1009,N_1059);
or U1333 (N_1333,N_1141,N_1187);
and U1334 (N_1334,N_1108,N_1095);
or U1335 (N_1335,N_1020,N_1003);
nand U1336 (N_1336,N_1051,N_1080);
and U1337 (N_1337,N_1096,N_1198);
nor U1338 (N_1338,N_1161,N_1018);
or U1339 (N_1339,N_1093,N_1034);
and U1340 (N_1340,N_1188,N_1073);
or U1341 (N_1341,N_1003,N_1067);
or U1342 (N_1342,N_1004,N_1144);
nand U1343 (N_1343,N_1024,N_1196);
nand U1344 (N_1344,N_1055,N_1127);
or U1345 (N_1345,N_1006,N_1102);
and U1346 (N_1346,N_1065,N_1157);
xnor U1347 (N_1347,N_1117,N_1068);
xnor U1348 (N_1348,N_1159,N_1081);
xor U1349 (N_1349,N_1094,N_1018);
and U1350 (N_1350,N_1178,N_1159);
nand U1351 (N_1351,N_1026,N_1164);
nor U1352 (N_1352,N_1107,N_1055);
and U1353 (N_1353,N_1082,N_1140);
nor U1354 (N_1354,N_1168,N_1063);
or U1355 (N_1355,N_1061,N_1114);
nor U1356 (N_1356,N_1000,N_1118);
or U1357 (N_1357,N_1106,N_1147);
nor U1358 (N_1358,N_1056,N_1097);
or U1359 (N_1359,N_1177,N_1043);
xnor U1360 (N_1360,N_1057,N_1153);
nand U1361 (N_1361,N_1041,N_1062);
nor U1362 (N_1362,N_1079,N_1142);
nand U1363 (N_1363,N_1066,N_1125);
nor U1364 (N_1364,N_1067,N_1134);
xor U1365 (N_1365,N_1079,N_1060);
nor U1366 (N_1366,N_1177,N_1128);
xnor U1367 (N_1367,N_1111,N_1104);
nand U1368 (N_1368,N_1084,N_1186);
nor U1369 (N_1369,N_1195,N_1097);
or U1370 (N_1370,N_1119,N_1090);
or U1371 (N_1371,N_1087,N_1028);
xor U1372 (N_1372,N_1142,N_1162);
or U1373 (N_1373,N_1026,N_1046);
and U1374 (N_1374,N_1015,N_1049);
or U1375 (N_1375,N_1106,N_1034);
or U1376 (N_1376,N_1186,N_1133);
nand U1377 (N_1377,N_1173,N_1195);
nand U1378 (N_1378,N_1198,N_1041);
nand U1379 (N_1379,N_1116,N_1096);
xor U1380 (N_1380,N_1094,N_1125);
xor U1381 (N_1381,N_1196,N_1169);
nand U1382 (N_1382,N_1012,N_1016);
nand U1383 (N_1383,N_1009,N_1011);
and U1384 (N_1384,N_1019,N_1043);
nand U1385 (N_1385,N_1079,N_1062);
or U1386 (N_1386,N_1016,N_1014);
or U1387 (N_1387,N_1085,N_1120);
nor U1388 (N_1388,N_1127,N_1082);
and U1389 (N_1389,N_1050,N_1194);
nand U1390 (N_1390,N_1197,N_1093);
or U1391 (N_1391,N_1137,N_1058);
xnor U1392 (N_1392,N_1083,N_1047);
nand U1393 (N_1393,N_1040,N_1166);
xnor U1394 (N_1394,N_1154,N_1034);
xor U1395 (N_1395,N_1142,N_1092);
nor U1396 (N_1396,N_1071,N_1090);
nor U1397 (N_1397,N_1096,N_1082);
and U1398 (N_1398,N_1127,N_1050);
nand U1399 (N_1399,N_1178,N_1010);
xor U1400 (N_1400,N_1243,N_1213);
xnor U1401 (N_1401,N_1311,N_1253);
xnor U1402 (N_1402,N_1260,N_1273);
or U1403 (N_1403,N_1383,N_1327);
or U1404 (N_1404,N_1219,N_1355);
xnor U1405 (N_1405,N_1325,N_1397);
or U1406 (N_1406,N_1282,N_1294);
xnor U1407 (N_1407,N_1255,N_1240);
nand U1408 (N_1408,N_1399,N_1258);
nor U1409 (N_1409,N_1335,N_1344);
xnor U1410 (N_1410,N_1370,N_1387);
nor U1411 (N_1411,N_1205,N_1295);
nand U1412 (N_1412,N_1338,N_1236);
nand U1413 (N_1413,N_1284,N_1220);
nand U1414 (N_1414,N_1334,N_1352);
xor U1415 (N_1415,N_1283,N_1376);
xor U1416 (N_1416,N_1365,N_1238);
and U1417 (N_1417,N_1249,N_1268);
or U1418 (N_1418,N_1230,N_1209);
nand U1419 (N_1419,N_1218,N_1277);
xor U1420 (N_1420,N_1200,N_1212);
or U1421 (N_1421,N_1287,N_1224);
or U1422 (N_1422,N_1392,N_1321);
nand U1423 (N_1423,N_1271,N_1278);
nand U1424 (N_1424,N_1329,N_1353);
and U1425 (N_1425,N_1225,N_1281);
and U1426 (N_1426,N_1201,N_1292);
and U1427 (N_1427,N_1246,N_1342);
nand U1428 (N_1428,N_1316,N_1384);
xnor U1429 (N_1429,N_1211,N_1233);
or U1430 (N_1430,N_1214,N_1361);
xnor U1431 (N_1431,N_1366,N_1373);
nor U1432 (N_1432,N_1296,N_1336);
or U1433 (N_1433,N_1259,N_1324);
or U1434 (N_1434,N_1377,N_1279);
nor U1435 (N_1435,N_1348,N_1252);
nand U1436 (N_1436,N_1322,N_1363);
or U1437 (N_1437,N_1326,N_1372);
and U1438 (N_1438,N_1378,N_1358);
nor U1439 (N_1439,N_1379,N_1398);
xor U1440 (N_1440,N_1306,N_1232);
and U1441 (N_1441,N_1202,N_1264);
and U1442 (N_1442,N_1333,N_1357);
nor U1443 (N_1443,N_1257,N_1339);
xor U1444 (N_1444,N_1234,N_1263);
nor U1445 (N_1445,N_1269,N_1347);
xor U1446 (N_1446,N_1204,N_1251);
nor U1447 (N_1447,N_1275,N_1228);
or U1448 (N_1448,N_1297,N_1315);
or U1449 (N_1449,N_1276,N_1368);
and U1450 (N_1450,N_1262,N_1291);
or U1451 (N_1451,N_1305,N_1394);
and U1452 (N_1452,N_1288,N_1300);
nand U1453 (N_1453,N_1241,N_1235);
xnor U1454 (N_1454,N_1239,N_1345);
nor U1455 (N_1455,N_1303,N_1266);
and U1456 (N_1456,N_1364,N_1286);
and U1457 (N_1457,N_1261,N_1391);
xor U1458 (N_1458,N_1285,N_1307);
xor U1459 (N_1459,N_1270,N_1374);
nor U1460 (N_1460,N_1362,N_1237);
xnor U1461 (N_1461,N_1346,N_1280);
nor U1462 (N_1462,N_1308,N_1371);
or U1463 (N_1463,N_1317,N_1393);
and U1464 (N_1464,N_1227,N_1385);
nor U1465 (N_1465,N_1206,N_1369);
nand U1466 (N_1466,N_1323,N_1267);
nor U1467 (N_1467,N_1331,N_1217);
nor U1468 (N_1468,N_1229,N_1254);
or U1469 (N_1469,N_1312,N_1203);
xor U1470 (N_1470,N_1247,N_1386);
nor U1471 (N_1471,N_1256,N_1349);
xnor U1472 (N_1472,N_1341,N_1210);
or U1473 (N_1473,N_1265,N_1223);
or U1474 (N_1474,N_1304,N_1375);
or U1475 (N_1475,N_1222,N_1299);
and U1476 (N_1476,N_1290,N_1302);
or U1477 (N_1477,N_1388,N_1359);
nor U1478 (N_1478,N_1343,N_1293);
or U1479 (N_1479,N_1298,N_1367);
or U1480 (N_1480,N_1313,N_1340);
nor U1481 (N_1481,N_1314,N_1250);
nand U1482 (N_1482,N_1382,N_1389);
or U1483 (N_1483,N_1350,N_1318);
and U1484 (N_1484,N_1330,N_1272);
xor U1485 (N_1485,N_1289,N_1309);
nor U1486 (N_1486,N_1390,N_1301);
and U1487 (N_1487,N_1221,N_1310);
nor U1488 (N_1488,N_1351,N_1274);
nor U1489 (N_1489,N_1231,N_1207);
and U1490 (N_1490,N_1337,N_1208);
xnor U1491 (N_1491,N_1396,N_1395);
xnor U1492 (N_1492,N_1319,N_1332);
and U1493 (N_1493,N_1380,N_1245);
or U1494 (N_1494,N_1360,N_1215);
nand U1495 (N_1495,N_1248,N_1216);
xor U1496 (N_1496,N_1226,N_1356);
or U1497 (N_1497,N_1242,N_1381);
xor U1498 (N_1498,N_1354,N_1320);
or U1499 (N_1499,N_1244,N_1328);
nand U1500 (N_1500,N_1322,N_1328);
xor U1501 (N_1501,N_1226,N_1365);
nand U1502 (N_1502,N_1207,N_1318);
or U1503 (N_1503,N_1218,N_1281);
nor U1504 (N_1504,N_1360,N_1307);
nor U1505 (N_1505,N_1262,N_1267);
xor U1506 (N_1506,N_1347,N_1237);
and U1507 (N_1507,N_1239,N_1309);
xnor U1508 (N_1508,N_1394,N_1221);
xnor U1509 (N_1509,N_1339,N_1309);
xnor U1510 (N_1510,N_1363,N_1224);
and U1511 (N_1511,N_1325,N_1351);
nand U1512 (N_1512,N_1204,N_1202);
nand U1513 (N_1513,N_1366,N_1328);
and U1514 (N_1514,N_1263,N_1250);
nand U1515 (N_1515,N_1358,N_1329);
xor U1516 (N_1516,N_1326,N_1283);
nand U1517 (N_1517,N_1236,N_1322);
or U1518 (N_1518,N_1389,N_1279);
nor U1519 (N_1519,N_1390,N_1335);
xnor U1520 (N_1520,N_1388,N_1363);
or U1521 (N_1521,N_1258,N_1338);
and U1522 (N_1522,N_1270,N_1361);
and U1523 (N_1523,N_1254,N_1396);
xor U1524 (N_1524,N_1272,N_1232);
or U1525 (N_1525,N_1237,N_1357);
or U1526 (N_1526,N_1290,N_1372);
nor U1527 (N_1527,N_1244,N_1308);
nand U1528 (N_1528,N_1384,N_1329);
nor U1529 (N_1529,N_1379,N_1272);
and U1530 (N_1530,N_1240,N_1344);
or U1531 (N_1531,N_1232,N_1376);
nor U1532 (N_1532,N_1323,N_1266);
nand U1533 (N_1533,N_1212,N_1306);
or U1534 (N_1534,N_1228,N_1288);
or U1535 (N_1535,N_1369,N_1216);
and U1536 (N_1536,N_1375,N_1289);
and U1537 (N_1537,N_1237,N_1234);
and U1538 (N_1538,N_1327,N_1268);
nor U1539 (N_1539,N_1223,N_1369);
nand U1540 (N_1540,N_1294,N_1249);
and U1541 (N_1541,N_1335,N_1363);
nor U1542 (N_1542,N_1287,N_1337);
nand U1543 (N_1543,N_1325,N_1213);
nor U1544 (N_1544,N_1323,N_1369);
or U1545 (N_1545,N_1357,N_1242);
nor U1546 (N_1546,N_1390,N_1253);
or U1547 (N_1547,N_1315,N_1221);
and U1548 (N_1548,N_1203,N_1345);
nand U1549 (N_1549,N_1296,N_1241);
nor U1550 (N_1550,N_1304,N_1204);
nand U1551 (N_1551,N_1318,N_1292);
nor U1552 (N_1552,N_1283,N_1319);
nand U1553 (N_1553,N_1275,N_1236);
nand U1554 (N_1554,N_1225,N_1221);
and U1555 (N_1555,N_1256,N_1253);
nor U1556 (N_1556,N_1352,N_1360);
nand U1557 (N_1557,N_1300,N_1274);
xnor U1558 (N_1558,N_1236,N_1309);
nor U1559 (N_1559,N_1322,N_1375);
and U1560 (N_1560,N_1206,N_1229);
nor U1561 (N_1561,N_1319,N_1292);
or U1562 (N_1562,N_1281,N_1203);
and U1563 (N_1563,N_1383,N_1212);
nand U1564 (N_1564,N_1279,N_1280);
xnor U1565 (N_1565,N_1235,N_1322);
nand U1566 (N_1566,N_1208,N_1344);
nor U1567 (N_1567,N_1271,N_1248);
and U1568 (N_1568,N_1322,N_1387);
or U1569 (N_1569,N_1382,N_1319);
or U1570 (N_1570,N_1294,N_1338);
or U1571 (N_1571,N_1398,N_1233);
nor U1572 (N_1572,N_1365,N_1237);
and U1573 (N_1573,N_1306,N_1251);
or U1574 (N_1574,N_1371,N_1337);
and U1575 (N_1575,N_1386,N_1283);
nor U1576 (N_1576,N_1238,N_1331);
nor U1577 (N_1577,N_1305,N_1328);
and U1578 (N_1578,N_1214,N_1251);
nand U1579 (N_1579,N_1364,N_1317);
and U1580 (N_1580,N_1353,N_1350);
nor U1581 (N_1581,N_1385,N_1392);
and U1582 (N_1582,N_1386,N_1378);
and U1583 (N_1583,N_1389,N_1398);
nand U1584 (N_1584,N_1246,N_1215);
nand U1585 (N_1585,N_1312,N_1383);
nor U1586 (N_1586,N_1227,N_1318);
or U1587 (N_1587,N_1324,N_1216);
or U1588 (N_1588,N_1326,N_1282);
nor U1589 (N_1589,N_1321,N_1209);
and U1590 (N_1590,N_1287,N_1353);
and U1591 (N_1591,N_1329,N_1307);
or U1592 (N_1592,N_1284,N_1295);
nand U1593 (N_1593,N_1312,N_1238);
nor U1594 (N_1594,N_1396,N_1238);
xor U1595 (N_1595,N_1260,N_1367);
and U1596 (N_1596,N_1340,N_1240);
xnor U1597 (N_1597,N_1225,N_1368);
or U1598 (N_1598,N_1312,N_1391);
nand U1599 (N_1599,N_1223,N_1356);
and U1600 (N_1600,N_1514,N_1564);
xor U1601 (N_1601,N_1455,N_1597);
or U1602 (N_1602,N_1596,N_1434);
nor U1603 (N_1603,N_1568,N_1582);
xnor U1604 (N_1604,N_1433,N_1479);
nor U1605 (N_1605,N_1586,N_1456);
nand U1606 (N_1606,N_1452,N_1449);
nand U1607 (N_1607,N_1497,N_1553);
nor U1608 (N_1608,N_1448,N_1579);
or U1609 (N_1609,N_1400,N_1439);
nand U1610 (N_1610,N_1559,N_1469);
or U1611 (N_1611,N_1570,N_1598);
xnor U1612 (N_1612,N_1577,N_1499);
and U1613 (N_1613,N_1571,N_1556);
nor U1614 (N_1614,N_1583,N_1515);
nand U1615 (N_1615,N_1493,N_1401);
nor U1616 (N_1616,N_1555,N_1405);
nor U1617 (N_1617,N_1422,N_1413);
and U1618 (N_1618,N_1410,N_1591);
nand U1619 (N_1619,N_1446,N_1522);
nand U1620 (N_1620,N_1545,N_1462);
nor U1621 (N_1621,N_1560,N_1421);
xnor U1622 (N_1622,N_1593,N_1411);
nor U1623 (N_1623,N_1454,N_1489);
or U1624 (N_1624,N_1572,N_1477);
nand U1625 (N_1625,N_1415,N_1471);
xor U1626 (N_1626,N_1594,N_1419);
nand U1627 (N_1627,N_1547,N_1408);
nor U1628 (N_1628,N_1500,N_1566);
and U1629 (N_1629,N_1428,N_1531);
nand U1630 (N_1630,N_1552,N_1460);
nor U1631 (N_1631,N_1447,N_1534);
or U1632 (N_1632,N_1521,N_1474);
nor U1633 (N_1633,N_1498,N_1403);
nand U1634 (N_1634,N_1592,N_1540);
or U1635 (N_1635,N_1542,N_1561);
nor U1636 (N_1636,N_1416,N_1520);
and U1637 (N_1637,N_1495,N_1588);
nor U1638 (N_1638,N_1412,N_1490);
or U1639 (N_1639,N_1453,N_1457);
xnor U1640 (N_1640,N_1506,N_1575);
nor U1641 (N_1641,N_1461,N_1476);
nor U1642 (N_1642,N_1468,N_1539);
nand U1643 (N_1643,N_1451,N_1525);
or U1644 (N_1644,N_1440,N_1536);
xor U1645 (N_1645,N_1424,N_1507);
and U1646 (N_1646,N_1427,N_1423);
xnor U1647 (N_1647,N_1426,N_1523);
xnor U1648 (N_1648,N_1467,N_1546);
and U1649 (N_1649,N_1470,N_1535);
nand U1650 (N_1650,N_1492,N_1578);
or U1651 (N_1651,N_1431,N_1524);
and U1652 (N_1652,N_1502,N_1409);
and U1653 (N_1653,N_1541,N_1558);
xnor U1654 (N_1654,N_1458,N_1473);
and U1655 (N_1655,N_1406,N_1543);
and U1656 (N_1656,N_1436,N_1425);
and U1657 (N_1657,N_1587,N_1528);
or U1658 (N_1658,N_1450,N_1465);
xor U1659 (N_1659,N_1483,N_1438);
or U1660 (N_1660,N_1418,N_1485);
nor U1661 (N_1661,N_1513,N_1445);
nor U1662 (N_1662,N_1501,N_1517);
nor U1663 (N_1663,N_1565,N_1420);
and U1664 (N_1664,N_1519,N_1494);
and U1665 (N_1665,N_1437,N_1576);
and U1666 (N_1666,N_1590,N_1538);
and U1667 (N_1667,N_1599,N_1487);
xor U1668 (N_1668,N_1488,N_1585);
or U1669 (N_1669,N_1484,N_1402);
nand U1670 (N_1670,N_1509,N_1532);
or U1671 (N_1671,N_1518,N_1404);
nand U1672 (N_1672,N_1595,N_1512);
or U1673 (N_1673,N_1526,N_1580);
nor U1674 (N_1674,N_1527,N_1510);
and U1675 (N_1675,N_1491,N_1511);
and U1676 (N_1676,N_1463,N_1549);
nand U1677 (N_1677,N_1464,N_1504);
nand U1678 (N_1678,N_1472,N_1430);
nor U1679 (N_1679,N_1466,N_1533);
or U1680 (N_1680,N_1569,N_1567);
nand U1681 (N_1681,N_1589,N_1486);
xnor U1682 (N_1682,N_1435,N_1459);
xor U1683 (N_1683,N_1505,N_1562);
nand U1684 (N_1684,N_1478,N_1530);
or U1685 (N_1685,N_1496,N_1481);
nand U1686 (N_1686,N_1508,N_1444);
nand U1687 (N_1687,N_1557,N_1550);
nor U1688 (N_1688,N_1407,N_1581);
xor U1689 (N_1689,N_1551,N_1516);
and U1690 (N_1690,N_1443,N_1573);
nor U1691 (N_1691,N_1414,N_1563);
xor U1692 (N_1692,N_1503,N_1544);
and U1693 (N_1693,N_1417,N_1529);
and U1694 (N_1694,N_1584,N_1548);
xnor U1695 (N_1695,N_1480,N_1482);
nand U1696 (N_1696,N_1475,N_1441);
or U1697 (N_1697,N_1574,N_1554);
nor U1698 (N_1698,N_1432,N_1442);
nor U1699 (N_1699,N_1429,N_1537);
nor U1700 (N_1700,N_1525,N_1498);
nand U1701 (N_1701,N_1560,N_1475);
xor U1702 (N_1702,N_1490,N_1543);
xor U1703 (N_1703,N_1432,N_1556);
nand U1704 (N_1704,N_1454,N_1467);
xor U1705 (N_1705,N_1401,N_1578);
and U1706 (N_1706,N_1551,N_1462);
nor U1707 (N_1707,N_1548,N_1449);
nand U1708 (N_1708,N_1533,N_1525);
and U1709 (N_1709,N_1490,N_1526);
xnor U1710 (N_1710,N_1578,N_1534);
or U1711 (N_1711,N_1524,N_1440);
nand U1712 (N_1712,N_1440,N_1427);
nor U1713 (N_1713,N_1536,N_1579);
nand U1714 (N_1714,N_1415,N_1427);
nor U1715 (N_1715,N_1427,N_1490);
xor U1716 (N_1716,N_1588,N_1443);
nor U1717 (N_1717,N_1571,N_1551);
and U1718 (N_1718,N_1531,N_1403);
or U1719 (N_1719,N_1450,N_1570);
and U1720 (N_1720,N_1568,N_1579);
or U1721 (N_1721,N_1583,N_1565);
nand U1722 (N_1722,N_1560,N_1423);
nand U1723 (N_1723,N_1432,N_1423);
nand U1724 (N_1724,N_1531,N_1409);
xor U1725 (N_1725,N_1446,N_1448);
nor U1726 (N_1726,N_1448,N_1586);
nor U1727 (N_1727,N_1498,N_1406);
nor U1728 (N_1728,N_1440,N_1528);
nand U1729 (N_1729,N_1584,N_1591);
or U1730 (N_1730,N_1554,N_1466);
nand U1731 (N_1731,N_1540,N_1446);
and U1732 (N_1732,N_1454,N_1518);
xor U1733 (N_1733,N_1579,N_1584);
nand U1734 (N_1734,N_1427,N_1417);
nand U1735 (N_1735,N_1502,N_1453);
and U1736 (N_1736,N_1571,N_1568);
nor U1737 (N_1737,N_1465,N_1569);
nor U1738 (N_1738,N_1572,N_1415);
xor U1739 (N_1739,N_1536,N_1589);
xnor U1740 (N_1740,N_1408,N_1543);
xnor U1741 (N_1741,N_1520,N_1466);
or U1742 (N_1742,N_1588,N_1520);
xor U1743 (N_1743,N_1525,N_1551);
or U1744 (N_1744,N_1439,N_1544);
and U1745 (N_1745,N_1473,N_1571);
nor U1746 (N_1746,N_1448,N_1533);
xnor U1747 (N_1747,N_1550,N_1437);
nor U1748 (N_1748,N_1427,N_1550);
and U1749 (N_1749,N_1414,N_1519);
xor U1750 (N_1750,N_1400,N_1517);
or U1751 (N_1751,N_1405,N_1433);
or U1752 (N_1752,N_1519,N_1416);
and U1753 (N_1753,N_1531,N_1463);
and U1754 (N_1754,N_1547,N_1579);
xor U1755 (N_1755,N_1556,N_1481);
nor U1756 (N_1756,N_1504,N_1454);
xor U1757 (N_1757,N_1470,N_1421);
nand U1758 (N_1758,N_1535,N_1539);
and U1759 (N_1759,N_1551,N_1543);
nor U1760 (N_1760,N_1435,N_1495);
and U1761 (N_1761,N_1532,N_1597);
or U1762 (N_1762,N_1505,N_1448);
or U1763 (N_1763,N_1476,N_1480);
and U1764 (N_1764,N_1459,N_1546);
nor U1765 (N_1765,N_1568,N_1532);
xor U1766 (N_1766,N_1549,N_1565);
and U1767 (N_1767,N_1562,N_1408);
nor U1768 (N_1768,N_1535,N_1543);
xor U1769 (N_1769,N_1594,N_1554);
xor U1770 (N_1770,N_1408,N_1585);
xnor U1771 (N_1771,N_1538,N_1474);
and U1772 (N_1772,N_1421,N_1484);
xnor U1773 (N_1773,N_1486,N_1536);
or U1774 (N_1774,N_1516,N_1500);
nand U1775 (N_1775,N_1489,N_1421);
xor U1776 (N_1776,N_1437,N_1416);
nor U1777 (N_1777,N_1469,N_1582);
or U1778 (N_1778,N_1527,N_1514);
or U1779 (N_1779,N_1561,N_1587);
nor U1780 (N_1780,N_1472,N_1576);
nand U1781 (N_1781,N_1491,N_1449);
nor U1782 (N_1782,N_1471,N_1458);
xnor U1783 (N_1783,N_1482,N_1559);
nand U1784 (N_1784,N_1514,N_1404);
nor U1785 (N_1785,N_1425,N_1582);
or U1786 (N_1786,N_1487,N_1458);
and U1787 (N_1787,N_1545,N_1575);
or U1788 (N_1788,N_1581,N_1483);
nand U1789 (N_1789,N_1518,N_1554);
xor U1790 (N_1790,N_1440,N_1489);
and U1791 (N_1791,N_1478,N_1571);
xor U1792 (N_1792,N_1548,N_1560);
xnor U1793 (N_1793,N_1484,N_1442);
xor U1794 (N_1794,N_1556,N_1539);
and U1795 (N_1795,N_1475,N_1574);
xnor U1796 (N_1796,N_1501,N_1450);
nor U1797 (N_1797,N_1491,N_1413);
and U1798 (N_1798,N_1420,N_1541);
and U1799 (N_1799,N_1521,N_1498);
and U1800 (N_1800,N_1677,N_1741);
xnor U1801 (N_1801,N_1634,N_1715);
xor U1802 (N_1802,N_1629,N_1797);
and U1803 (N_1803,N_1753,N_1725);
nor U1804 (N_1804,N_1652,N_1746);
nor U1805 (N_1805,N_1603,N_1720);
xnor U1806 (N_1806,N_1617,N_1755);
and U1807 (N_1807,N_1718,N_1689);
nor U1808 (N_1808,N_1742,N_1692);
nand U1809 (N_1809,N_1666,N_1782);
xnor U1810 (N_1810,N_1748,N_1616);
xor U1811 (N_1811,N_1785,N_1735);
and U1812 (N_1812,N_1710,N_1767);
nand U1813 (N_1813,N_1757,N_1758);
nand U1814 (N_1814,N_1698,N_1705);
or U1815 (N_1815,N_1685,N_1632);
nand U1816 (N_1816,N_1633,N_1795);
or U1817 (N_1817,N_1619,N_1605);
nand U1818 (N_1818,N_1607,N_1769);
nor U1819 (N_1819,N_1671,N_1760);
nand U1820 (N_1820,N_1655,N_1793);
xnor U1821 (N_1821,N_1790,N_1747);
or U1822 (N_1822,N_1602,N_1611);
nand U1823 (N_1823,N_1764,N_1623);
xnor U1824 (N_1824,N_1660,N_1700);
and U1825 (N_1825,N_1686,N_1657);
and U1826 (N_1826,N_1658,N_1749);
nand U1827 (N_1827,N_1775,N_1676);
and U1828 (N_1828,N_1640,N_1631);
or U1829 (N_1829,N_1745,N_1601);
or U1830 (N_1830,N_1636,N_1643);
or U1831 (N_1831,N_1694,N_1739);
nand U1832 (N_1832,N_1699,N_1743);
or U1833 (N_1833,N_1615,N_1695);
xor U1834 (N_1834,N_1754,N_1794);
nor U1835 (N_1835,N_1609,N_1621);
and U1836 (N_1836,N_1774,N_1721);
and U1837 (N_1837,N_1722,N_1751);
nand U1838 (N_1838,N_1687,N_1723);
xnor U1839 (N_1839,N_1620,N_1724);
and U1840 (N_1840,N_1780,N_1702);
and U1841 (N_1841,N_1708,N_1712);
xnor U1842 (N_1842,N_1777,N_1784);
or U1843 (N_1843,N_1740,N_1681);
nor U1844 (N_1844,N_1679,N_1642);
nor U1845 (N_1845,N_1759,N_1690);
nand U1846 (N_1846,N_1618,N_1726);
or U1847 (N_1847,N_1661,N_1651);
and U1848 (N_1848,N_1761,N_1783);
nor U1849 (N_1849,N_1637,N_1647);
nor U1850 (N_1850,N_1664,N_1706);
xor U1851 (N_1851,N_1614,N_1675);
xnor U1852 (N_1852,N_1798,N_1772);
nor U1853 (N_1853,N_1729,N_1737);
nand U1854 (N_1854,N_1734,N_1613);
xnor U1855 (N_1855,N_1799,N_1779);
nand U1856 (N_1856,N_1683,N_1771);
or U1857 (N_1857,N_1778,N_1731);
xnor U1858 (N_1858,N_1670,N_1752);
and U1859 (N_1859,N_1641,N_1688);
nand U1860 (N_1860,N_1668,N_1682);
or U1861 (N_1861,N_1606,N_1669);
nand U1862 (N_1862,N_1768,N_1628);
nor U1863 (N_1863,N_1717,N_1714);
or U1864 (N_1864,N_1604,N_1646);
or U1865 (N_1865,N_1719,N_1659);
xor U1866 (N_1866,N_1787,N_1770);
xor U1867 (N_1867,N_1704,N_1762);
nor U1868 (N_1868,N_1750,N_1736);
nand U1869 (N_1869,N_1674,N_1709);
xnor U1870 (N_1870,N_1766,N_1733);
and U1871 (N_1871,N_1678,N_1638);
or U1872 (N_1872,N_1622,N_1791);
or U1873 (N_1873,N_1716,N_1744);
nand U1874 (N_1874,N_1789,N_1612);
and U1875 (N_1875,N_1765,N_1663);
and U1876 (N_1876,N_1653,N_1667);
nand U1877 (N_1877,N_1707,N_1672);
and U1878 (N_1878,N_1630,N_1773);
and U1879 (N_1879,N_1673,N_1713);
nor U1880 (N_1880,N_1639,N_1732);
nor U1881 (N_1881,N_1786,N_1796);
or U1882 (N_1882,N_1756,N_1624);
and U1883 (N_1883,N_1691,N_1697);
nor U1884 (N_1884,N_1781,N_1645);
nand U1885 (N_1885,N_1792,N_1656);
nand U1886 (N_1886,N_1680,N_1684);
nor U1887 (N_1887,N_1788,N_1711);
xnor U1888 (N_1888,N_1693,N_1650);
nor U1889 (N_1889,N_1610,N_1625);
nand U1890 (N_1890,N_1703,N_1654);
or U1891 (N_1891,N_1763,N_1648);
and U1892 (N_1892,N_1627,N_1665);
and U1893 (N_1893,N_1696,N_1626);
xor U1894 (N_1894,N_1644,N_1730);
nand U1895 (N_1895,N_1776,N_1727);
and U1896 (N_1896,N_1600,N_1701);
xor U1897 (N_1897,N_1662,N_1738);
and U1898 (N_1898,N_1635,N_1728);
xor U1899 (N_1899,N_1608,N_1649);
and U1900 (N_1900,N_1670,N_1740);
xor U1901 (N_1901,N_1717,N_1683);
and U1902 (N_1902,N_1740,N_1754);
and U1903 (N_1903,N_1781,N_1793);
nand U1904 (N_1904,N_1779,N_1705);
and U1905 (N_1905,N_1653,N_1794);
nand U1906 (N_1906,N_1719,N_1740);
xnor U1907 (N_1907,N_1719,N_1785);
nand U1908 (N_1908,N_1667,N_1610);
nand U1909 (N_1909,N_1756,N_1646);
nand U1910 (N_1910,N_1776,N_1614);
and U1911 (N_1911,N_1613,N_1663);
xnor U1912 (N_1912,N_1743,N_1790);
xor U1913 (N_1913,N_1740,N_1690);
xnor U1914 (N_1914,N_1727,N_1716);
xnor U1915 (N_1915,N_1730,N_1726);
and U1916 (N_1916,N_1625,N_1679);
or U1917 (N_1917,N_1658,N_1656);
nand U1918 (N_1918,N_1767,N_1761);
nand U1919 (N_1919,N_1732,N_1638);
and U1920 (N_1920,N_1741,N_1615);
or U1921 (N_1921,N_1672,N_1683);
nor U1922 (N_1922,N_1606,N_1698);
xor U1923 (N_1923,N_1644,N_1628);
nand U1924 (N_1924,N_1681,N_1704);
and U1925 (N_1925,N_1791,N_1630);
and U1926 (N_1926,N_1729,N_1750);
nand U1927 (N_1927,N_1685,N_1704);
or U1928 (N_1928,N_1744,N_1691);
nor U1929 (N_1929,N_1655,N_1727);
and U1930 (N_1930,N_1708,N_1677);
nor U1931 (N_1931,N_1704,N_1651);
xor U1932 (N_1932,N_1774,N_1613);
or U1933 (N_1933,N_1654,N_1659);
nand U1934 (N_1934,N_1619,N_1712);
xor U1935 (N_1935,N_1798,N_1633);
xnor U1936 (N_1936,N_1702,N_1662);
nor U1937 (N_1937,N_1739,N_1657);
nor U1938 (N_1938,N_1656,N_1744);
nand U1939 (N_1939,N_1702,N_1756);
nor U1940 (N_1940,N_1639,N_1765);
nand U1941 (N_1941,N_1658,N_1733);
nand U1942 (N_1942,N_1706,N_1613);
nor U1943 (N_1943,N_1742,N_1641);
nand U1944 (N_1944,N_1796,N_1731);
nand U1945 (N_1945,N_1790,N_1780);
nor U1946 (N_1946,N_1692,N_1740);
xnor U1947 (N_1947,N_1796,N_1724);
nor U1948 (N_1948,N_1627,N_1694);
or U1949 (N_1949,N_1634,N_1747);
nand U1950 (N_1950,N_1705,N_1706);
and U1951 (N_1951,N_1721,N_1737);
and U1952 (N_1952,N_1774,N_1719);
nor U1953 (N_1953,N_1637,N_1639);
and U1954 (N_1954,N_1772,N_1729);
nand U1955 (N_1955,N_1757,N_1676);
and U1956 (N_1956,N_1767,N_1666);
nor U1957 (N_1957,N_1680,N_1724);
nand U1958 (N_1958,N_1653,N_1744);
or U1959 (N_1959,N_1639,N_1610);
or U1960 (N_1960,N_1684,N_1782);
and U1961 (N_1961,N_1738,N_1751);
nand U1962 (N_1962,N_1739,N_1781);
or U1963 (N_1963,N_1615,N_1606);
or U1964 (N_1964,N_1641,N_1690);
and U1965 (N_1965,N_1708,N_1605);
nand U1966 (N_1966,N_1746,N_1717);
and U1967 (N_1967,N_1758,N_1621);
xnor U1968 (N_1968,N_1789,N_1781);
and U1969 (N_1969,N_1771,N_1613);
nand U1970 (N_1970,N_1730,N_1676);
and U1971 (N_1971,N_1683,N_1668);
nand U1972 (N_1972,N_1758,N_1730);
nor U1973 (N_1973,N_1641,N_1653);
or U1974 (N_1974,N_1722,N_1768);
and U1975 (N_1975,N_1742,N_1728);
and U1976 (N_1976,N_1773,N_1724);
xor U1977 (N_1977,N_1603,N_1799);
nand U1978 (N_1978,N_1706,N_1615);
xnor U1979 (N_1979,N_1663,N_1614);
or U1980 (N_1980,N_1672,N_1682);
nor U1981 (N_1981,N_1787,N_1624);
nand U1982 (N_1982,N_1788,N_1621);
xor U1983 (N_1983,N_1656,N_1643);
or U1984 (N_1984,N_1723,N_1647);
nand U1985 (N_1985,N_1680,N_1721);
nand U1986 (N_1986,N_1697,N_1645);
nand U1987 (N_1987,N_1637,N_1785);
or U1988 (N_1988,N_1794,N_1650);
xor U1989 (N_1989,N_1641,N_1708);
xnor U1990 (N_1990,N_1647,N_1628);
xnor U1991 (N_1991,N_1795,N_1731);
or U1992 (N_1992,N_1600,N_1647);
xor U1993 (N_1993,N_1765,N_1621);
or U1994 (N_1994,N_1665,N_1734);
nand U1995 (N_1995,N_1634,N_1617);
nor U1996 (N_1996,N_1650,N_1610);
and U1997 (N_1997,N_1671,N_1673);
nand U1998 (N_1998,N_1744,N_1642);
xor U1999 (N_1999,N_1748,N_1761);
or U2000 (N_2000,N_1982,N_1822);
or U2001 (N_2001,N_1827,N_1862);
or U2002 (N_2002,N_1857,N_1931);
and U2003 (N_2003,N_1996,N_1881);
nand U2004 (N_2004,N_1979,N_1856);
nor U2005 (N_2005,N_1945,N_1898);
and U2006 (N_2006,N_1937,N_1904);
and U2007 (N_2007,N_1861,N_1914);
nor U2008 (N_2008,N_1884,N_1954);
or U2009 (N_2009,N_1850,N_1915);
or U2010 (N_2010,N_1895,N_1909);
or U2011 (N_2011,N_1829,N_1941);
xnor U2012 (N_2012,N_1831,N_1913);
xor U2013 (N_2013,N_1835,N_1845);
nand U2014 (N_2014,N_1837,N_1801);
xnor U2015 (N_2015,N_1876,N_1974);
xnor U2016 (N_2016,N_1947,N_1965);
nor U2017 (N_2017,N_1961,N_1820);
nand U2018 (N_2018,N_1810,N_1806);
xnor U2019 (N_2019,N_1886,N_1929);
nor U2020 (N_2020,N_1936,N_1940);
and U2021 (N_2021,N_1891,N_1815);
nor U2022 (N_2022,N_1847,N_1848);
or U2023 (N_2023,N_1997,N_1869);
xor U2024 (N_2024,N_1853,N_1993);
xor U2025 (N_2025,N_1867,N_1935);
nor U2026 (N_2026,N_1973,N_1819);
and U2027 (N_2027,N_1870,N_1933);
and U2028 (N_2028,N_1934,N_1999);
or U2029 (N_2029,N_1920,N_1894);
xnor U2030 (N_2030,N_1800,N_1926);
nand U2031 (N_2031,N_1901,N_1987);
xnor U2032 (N_2032,N_1854,N_1988);
nor U2033 (N_2033,N_1942,N_1900);
and U2034 (N_2034,N_1991,N_1946);
nand U2035 (N_2035,N_1813,N_1808);
nor U2036 (N_2036,N_1834,N_1842);
and U2037 (N_2037,N_1989,N_1975);
nand U2038 (N_2038,N_1978,N_1922);
or U2039 (N_2039,N_1980,N_1944);
or U2040 (N_2040,N_1889,N_1849);
or U2041 (N_2041,N_1832,N_1807);
or U2042 (N_2042,N_1907,N_1938);
nor U2043 (N_2043,N_1874,N_1956);
and U2044 (N_2044,N_1983,N_1963);
xor U2045 (N_2045,N_1841,N_1921);
or U2046 (N_2046,N_1851,N_1888);
and U2047 (N_2047,N_1966,N_1868);
and U2048 (N_2048,N_1802,N_1823);
or U2049 (N_2049,N_1959,N_1899);
nand U2050 (N_2050,N_1878,N_1871);
nand U2051 (N_2051,N_1866,N_1836);
or U2052 (N_2052,N_1817,N_1830);
nand U2053 (N_2053,N_1890,N_1846);
nor U2054 (N_2054,N_1928,N_1984);
and U2055 (N_2055,N_1838,N_1863);
nand U2056 (N_2056,N_1818,N_1814);
xor U2057 (N_2057,N_1964,N_1967);
nor U2058 (N_2058,N_1816,N_1803);
nor U2059 (N_2059,N_1908,N_1952);
and U2060 (N_2060,N_1981,N_1809);
nand U2061 (N_2061,N_1804,N_1924);
xnor U2062 (N_2062,N_1925,N_1821);
and U2063 (N_2063,N_1958,N_1902);
nand U2064 (N_2064,N_1855,N_1805);
or U2065 (N_2065,N_1887,N_1918);
or U2066 (N_2066,N_1885,N_1950);
nor U2067 (N_2067,N_1949,N_1919);
and U2068 (N_2068,N_1923,N_1824);
xnor U2069 (N_2069,N_1916,N_1977);
xnor U2070 (N_2070,N_1873,N_1872);
and U2071 (N_2071,N_1828,N_1839);
nor U2072 (N_2072,N_1840,N_1972);
nor U2073 (N_2073,N_1833,N_1976);
nand U2074 (N_2074,N_1826,N_1843);
xnor U2075 (N_2075,N_1943,N_1852);
or U2076 (N_2076,N_1906,N_1892);
xor U2077 (N_2077,N_1932,N_1948);
or U2078 (N_2078,N_1992,N_1953);
and U2079 (N_2079,N_1875,N_1994);
xnor U2080 (N_2080,N_1910,N_1968);
nand U2081 (N_2081,N_1812,N_1939);
xor U2082 (N_2082,N_1917,N_1825);
and U2083 (N_2083,N_1877,N_1995);
and U2084 (N_2084,N_1990,N_1970);
nand U2085 (N_2085,N_1860,N_1883);
and U2086 (N_2086,N_1811,N_1912);
xor U2087 (N_2087,N_1962,N_1865);
and U2088 (N_2088,N_1858,N_1927);
nor U2089 (N_2089,N_1882,N_1960);
xor U2090 (N_2090,N_1985,N_1897);
and U2091 (N_2091,N_1864,N_1969);
and U2092 (N_2092,N_1844,N_1951);
and U2093 (N_2093,N_1911,N_1971);
nor U2094 (N_2094,N_1905,N_1957);
nand U2095 (N_2095,N_1896,N_1930);
nor U2096 (N_2096,N_1903,N_1893);
nor U2097 (N_2097,N_1859,N_1879);
nand U2098 (N_2098,N_1998,N_1880);
nor U2099 (N_2099,N_1955,N_1986);
and U2100 (N_2100,N_1945,N_1960);
nor U2101 (N_2101,N_1855,N_1884);
xor U2102 (N_2102,N_1800,N_1973);
or U2103 (N_2103,N_1910,N_1848);
nor U2104 (N_2104,N_1873,N_1851);
xor U2105 (N_2105,N_1973,N_1806);
nand U2106 (N_2106,N_1962,N_1889);
and U2107 (N_2107,N_1928,N_1831);
xor U2108 (N_2108,N_1973,N_1933);
and U2109 (N_2109,N_1960,N_1888);
nor U2110 (N_2110,N_1865,N_1973);
and U2111 (N_2111,N_1981,N_1986);
or U2112 (N_2112,N_1938,N_1849);
nand U2113 (N_2113,N_1802,N_1868);
and U2114 (N_2114,N_1998,N_1868);
xor U2115 (N_2115,N_1993,N_1893);
nor U2116 (N_2116,N_1989,N_1943);
or U2117 (N_2117,N_1996,N_1878);
nand U2118 (N_2118,N_1966,N_1825);
and U2119 (N_2119,N_1879,N_1823);
xor U2120 (N_2120,N_1910,N_1842);
nand U2121 (N_2121,N_1998,N_1838);
nand U2122 (N_2122,N_1876,N_1975);
or U2123 (N_2123,N_1822,N_1942);
nand U2124 (N_2124,N_1996,N_1981);
nor U2125 (N_2125,N_1912,N_1843);
nor U2126 (N_2126,N_1821,N_1806);
or U2127 (N_2127,N_1917,N_1961);
and U2128 (N_2128,N_1917,N_1953);
xnor U2129 (N_2129,N_1996,N_1833);
and U2130 (N_2130,N_1974,N_1911);
xor U2131 (N_2131,N_1904,N_1885);
and U2132 (N_2132,N_1875,N_1938);
or U2133 (N_2133,N_1847,N_1805);
nor U2134 (N_2134,N_1977,N_1950);
xor U2135 (N_2135,N_1978,N_1970);
and U2136 (N_2136,N_1813,N_1822);
xnor U2137 (N_2137,N_1923,N_1926);
nor U2138 (N_2138,N_1841,N_1948);
nor U2139 (N_2139,N_1847,N_1829);
nand U2140 (N_2140,N_1814,N_1906);
and U2141 (N_2141,N_1806,N_1873);
nand U2142 (N_2142,N_1938,N_1964);
and U2143 (N_2143,N_1815,N_1927);
nand U2144 (N_2144,N_1882,N_1878);
nand U2145 (N_2145,N_1914,N_1976);
nor U2146 (N_2146,N_1938,N_1806);
or U2147 (N_2147,N_1940,N_1889);
nor U2148 (N_2148,N_1935,N_1820);
xor U2149 (N_2149,N_1957,N_1831);
or U2150 (N_2150,N_1960,N_1845);
and U2151 (N_2151,N_1978,N_1891);
nor U2152 (N_2152,N_1813,N_1918);
or U2153 (N_2153,N_1975,N_1936);
xnor U2154 (N_2154,N_1816,N_1883);
nand U2155 (N_2155,N_1997,N_1820);
or U2156 (N_2156,N_1868,N_1936);
and U2157 (N_2157,N_1878,N_1832);
xor U2158 (N_2158,N_1976,N_1814);
nor U2159 (N_2159,N_1800,N_1809);
nor U2160 (N_2160,N_1899,N_1927);
or U2161 (N_2161,N_1933,N_1878);
and U2162 (N_2162,N_1858,N_1847);
or U2163 (N_2163,N_1973,N_1957);
and U2164 (N_2164,N_1863,N_1866);
or U2165 (N_2165,N_1924,N_1859);
nor U2166 (N_2166,N_1903,N_1833);
nand U2167 (N_2167,N_1973,N_1919);
xnor U2168 (N_2168,N_1882,N_1818);
nor U2169 (N_2169,N_1981,N_1849);
nor U2170 (N_2170,N_1856,N_1833);
or U2171 (N_2171,N_1996,N_1942);
nand U2172 (N_2172,N_1893,N_1886);
and U2173 (N_2173,N_1869,N_1991);
or U2174 (N_2174,N_1953,N_1804);
xor U2175 (N_2175,N_1933,N_1950);
and U2176 (N_2176,N_1905,N_1886);
nor U2177 (N_2177,N_1884,N_1835);
or U2178 (N_2178,N_1975,N_1966);
nand U2179 (N_2179,N_1885,N_1859);
nor U2180 (N_2180,N_1973,N_1949);
and U2181 (N_2181,N_1917,N_1983);
nand U2182 (N_2182,N_1822,N_1880);
and U2183 (N_2183,N_1846,N_1833);
nor U2184 (N_2184,N_1845,N_1881);
or U2185 (N_2185,N_1868,N_1880);
nand U2186 (N_2186,N_1859,N_1992);
and U2187 (N_2187,N_1828,N_1832);
or U2188 (N_2188,N_1882,N_1812);
xor U2189 (N_2189,N_1874,N_1801);
xnor U2190 (N_2190,N_1888,N_1903);
nor U2191 (N_2191,N_1803,N_1870);
and U2192 (N_2192,N_1899,N_1978);
xor U2193 (N_2193,N_1857,N_1809);
nor U2194 (N_2194,N_1880,N_1944);
and U2195 (N_2195,N_1885,N_1883);
xor U2196 (N_2196,N_1916,N_1844);
xnor U2197 (N_2197,N_1850,N_1855);
and U2198 (N_2198,N_1863,N_1814);
and U2199 (N_2199,N_1905,N_1962);
nand U2200 (N_2200,N_2088,N_2058);
nand U2201 (N_2201,N_2076,N_2027);
or U2202 (N_2202,N_2004,N_2104);
and U2203 (N_2203,N_2108,N_2073);
xnor U2204 (N_2204,N_2018,N_2143);
or U2205 (N_2205,N_2109,N_2006);
xnor U2206 (N_2206,N_2194,N_2033);
nor U2207 (N_2207,N_2131,N_2068);
nor U2208 (N_2208,N_2130,N_2064);
nand U2209 (N_2209,N_2127,N_2193);
and U2210 (N_2210,N_2145,N_2043);
nand U2211 (N_2211,N_2197,N_2053);
xor U2212 (N_2212,N_2045,N_2129);
nor U2213 (N_2213,N_2037,N_2132);
nand U2214 (N_2214,N_2093,N_2080);
and U2215 (N_2215,N_2026,N_2159);
nand U2216 (N_2216,N_2092,N_2103);
nor U2217 (N_2217,N_2141,N_2106);
and U2218 (N_2218,N_2154,N_2151);
nor U2219 (N_2219,N_2056,N_2126);
or U2220 (N_2220,N_2136,N_2015);
xor U2221 (N_2221,N_2157,N_2177);
and U2222 (N_2222,N_2101,N_2060);
xor U2223 (N_2223,N_2081,N_2147);
or U2224 (N_2224,N_2048,N_2174);
and U2225 (N_2225,N_2083,N_2155);
nor U2226 (N_2226,N_2114,N_2191);
nand U2227 (N_2227,N_2122,N_2019);
nor U2228 (N_2228,N_2119,N_2057);
nor U2229 (N_2229,N_2050,N_2062);
xnor U2230 (N_2230,N_2040,N_2002);
and U2231 (N_2231,N_2036,N_2035);
or U2232 (N_2232,N_2032,N_2166);
xor U2233 (N_2233,N_2051,N_2100);
and U2234 (N_2234,N_2180,N_2042);
and U2235 (N_2235,N_2156,N_2188);
and U2236 (N_2236,N_2117,N_2000);
and U2237 (N_2237,N_2094,N_2077);
and U2238 (N_2238,N_2190,N_2074);
xnor U2239 (N_2239,N_2063,N_2195);
xnor U2240 (N_2240,N_2181,N_2137);
nand U2241 (N_2241,N_2183,N_2008);
or U2242 (N_2242,N_2124,N_2087);
nor U2243 (N_2243,N_2164,N_2167);
nor U2244 (N_2244,N_2049,N_2084);
nand U2245 (N_2245,N_2070,N_2176);
or U2246 (N_2246,N_2171,N_2116);
nor U2247 (N_2247,N_2086,N_2115);
nand U2248 (N_2248,N_2091,N_2158);
nor U2249 (N_2249,N_2182,N_2142);
xnor U2250 (N_2250,N_2111,N_2067);
and U2251 (N_2251,N_2110,N_2134);
xnor U2252 (N_2252,N_2061,N_2007);
nor U2253 (N_2253,N_2003,N_2118);
nor U2254 (N_2254,N_2102,N_2113);
or U2255 (N_2255,N_2029,N_2161);
and U2256 (N_2256,N_2112,N_2028);
nand U2257 (N_2257,N_2082,N_2178);
and U2258 (N_2258,N_2135,N_2017);
nand U2259 (N_2259,N_2160,N_2005);
or U2260 (N_2260,N_2069,N_2123);
and U2261 (N_2261,N_2098,N_2184);
nand U2262 (N_2262,N_2031,N_2046);
nor U2263 (N_2263,N_2090,N_2079);
xnor U2264 (N_2264,N_2153,N_2140);
and U2265 (N_2265,N_2023,N_2096);
and U2266 (N_2266,N_2089,N_2075);
nand U2267 (N_2267,N_2199,N_2030);
and U2268 (N_2268,N_2144,N_2022);
or U2269 (N_2269,N_2078,N_2055);
nand U2270 (N_2270,N_2149,N_2010);
xor U2271 (N_2271,N_2001,N_2189);
nor U2272 (N_2272,N_2150,N_2196);
nor U2273 (N_2273,N_2009,N_2163);
and U2274 (N_2274,N_2138,N_2175);
xor U2275 (N_2275,N_2016,N_2165);
and U2276 (N_2276,N_2121,N_2024);
and U2277 (N_2277,N_2085,N_2128);
nor U2278 (N_2278,N_2152,N_2170);
nand U2279 (N_2279,N_2039,N_2162);
nand U2280 (N_2280,N_2059,N_2172);
xor U2281 (N_2281,N_2169,N_2139);
nand U2282 (N_2282,N_2125,N_2192);
or U2283 (N_2283,N_2052,N_2107);
xnor U2284 (N_2284,N_2025,N_2097);
or U2285 (N_2285,N_2148,N_2173);
or U2286 (N_2286,N_2099,N_2120);
or U2287 (N_2287,N_2198,N_2071);
and U2288 (N_2288,N_2187,N_2179);
or U2289 (N_2289,N_2105,N_2021);
xnor U2290 (N_2290,N_2012,N_2041);
nand U2291 (N_2291,N_2054,N_2186);
and U2292 (N_2292,N_2095,N_2034);
and U2293 (N_2293,N_2185,N_2168);
nand U2294 (N_2294,N_2020,N_2065);
or U2295 (N_2295,N_2047,N_2038);
and U2296 (N_2296,N_2072,N_2066);
or U2297 (N_2297,N_2044,N_2146);
xnor U2298 (N_2298,N_2011,N_2133);
or U2299 (N_2299,N_2013,N_2014);
or U2300 (N_2300,N_2156,N_2034);
nand U2301 (N_2301,N_2074,N_2182);
nor U2302 (N_2302,N_2072,N_2170);
and U2303 (N_2303,N_2132,N_2189);
or U2304 (N_2304,N_2025,N_2129);
and U2305 (N_2305,N_2038,N_2163);
or U2306 (N_2306,N_2174,N_2071);
or U2307 (N_2307,N_2145,N_2166);
or U2308 (N_2308,N_2113,N_2131);
or U2309 (N_2309,N_2040,N_2124);
and U2310 (N_2310,N_2100,N_2138);
or U2311 (N_2311,N_2119,N_2022);
nor U2312 (N_2312,N_2062,N_2110);
xnor U2313 (N_2313,N_2011,N_2028);
and U2314 (N_2314,N_2151,N_2063);
nand U2315 (N_2315,N_2023,N_2006);
xor U2316 (N_2316,N_2117,N_2136);
nor U2317 (N_2317,N_2108,N_2051);
xnor U2318 (N_2318,N_2178,N_2065);
or U2319 (N_2319,N_2066,N_2087);
or U2320 (N_2320,N_2098,N_2002);
or U2321 (N_2321,N_2166,N_2082);
and U2322 (N_2322,N_2020,N_2120);
or U2323 (N_2323,N_2073,N_2180);
nor U2324 (N_2324,N_2195,N_2072);
xor U2325 (N_2325,N_2156,N_2059);
nand U2326 (N_2326,N_2131,N_2159);
and U2327 (N_2327,N_2108,N_2034);
and U2328 (N_2328,N_2002,N_2028);
and U2329 (N_2329,N_2008,N_2049);
nor U2330 (N_2330,N_2061,N_2017);
or U2331 (N_2331,N_2077,N_2085);
or U2332 (N_2332,N_2181,N_2191);
nor U2333 (N_2333,N_2002,N_2092);
or U2334 (N_2334,N_2049,N_2035);
nor U2335 (N_2335,N_2159,N_2112);
and U2336 (N_2336,N_2023,N_2174);
xor U2337 (N_2337,N_2184,N_2188);
nor U2338 (N_2338,N_2049,N_2151);
xor U2339 (N_2339,N_2123,N_2004);
or U2340 (N_2340,N_2038,N_2152);
nor U2341 (N_2341,N_2127,N_2092);
and U2342 (N_2342,N_2043,N_2137);
or U2343 (N_2343,N_2095,N_2017);
nand U2344 (N_2344,N_2125,N_2185);
xnor U2345 (N_2345,N_2009,N_2119);
nand U2346 (N_2346,N_2092,N_2021);
nand U2347 (N_2347,N_2047,N_2009);
nor U2348 (N_2348,N_2126,N_2057);
or U2349 (N_2349,N_2133,N_2148);
nor U2350 (N_2350,N_2187,N_2027);
nor U2351 (N_2351,N_2007,N_2075);
nand U2352 (N_2352,N_2051,N_2192);
nand U2353 (N_2353,N_2069,N_2148);
nand U2354 (N_2354,N_2175,N_2098);
nand U2355 (N_2355,N_2153,N_2030);
or U2356 (N_2356,N_2109,N_2156);
or U2357 (N_2357,N_2184,N_2136);
xnor U2358 (N_2358,N_2013,N_2164);
and U2359 (N_2359,N_2137,N_2023);
xor U2360 (N_2360,N_2146,N_2064);
or U2361 (N_2361,N_2126,N_2166);
nand U2362 (N_2362,N_2091,N_2022);
nand U2363 (N_2363,N_2177,N_2185);
and U2364 (N_2364,N_2142,N_2050);
nor U2365 (N_2365,N_2064,N_2103);
or U2366 (N_2366,N_2077,N_2192);
xor U2367 (N_2367,N_2195,N_2146);
xor U2368 (N_2368,N_2027,N_2042);
nor U2369 (N_2369,N_2133,N_2010);
or U2370 (N_2370,N_2143,N_2154);
or U2371 (N_2371,N_2126,N_2161);
nor U2372 (N_2372,N_2106,N_2024);
nand U2373 (N_2373,N_2190,N_2016);
xor U2374 (N_2374,N_2033,N_2007);
nor U2375 (N_2375,N_2131,N_2144);
nor U2376 (N_2376,N_2006,N_2097);
or U2377 (N_2377,N_2165,N_2062);
xnor U2378 (N_2378,N_2043,N_2076);
xor U2379 (N_2379,N_2112,N_2111);
nor U2380 (N_2380,N_2097,N_2112);
and U2381 (N_2381,N_2104,N_2020);
or U2382 (N_2382,N_2023,N_2102);
nor U2383 (N_2383,N_2098,N_2139);
or U2384 (N_2384,N_2018,N_2149);
or U2385 (N_2385,N_2019,N_2149);
or U2386 (N_2386,N_2089,N_2103);
and U2387 (N_2387,N_2132,N_2150);
and U2388 (N_2388,N_2158,N_2105);
nor U2389 (N_2389,N_2024,N_2178);
or U2390 (N_2390,N_2120,N_2197);
xnor U2391 (N_2391,N_2137,N_2036);
xnor U2392 (N_2392,N_2167,N_2014);
nor U2393 (N_2393,N_2001,N_2157);
or U2394 (N_2394,N_2195,N_2022);
nand U2395 (N_2395,N_2164,N_2062);
nor U2396 (N_2396,N_2113,N_2044);
xnor U2397 (N_2397,N_2109,N_2159);
nand U2398 (N_2398,N_2113,N_2127);
xnor U2399 (N_2399,N_2081,N_2051);
xor U2400 (N_2400,N_2331,N_2260);
and U2401 (N_2401,N_2355,N_2387);
or U2402 (N_2402,N_2334,N_2245);
nand U2403 (N_2403,N_2290,N_2292);
and U2404 (N_2404,N_2218,N_2354);
and U2405 (N_2405,N_2214,N_2391);
nand U2406 (N_2406,N_2254,N_2266);
nor U2407 (N_2407,N_2208,N_2212);
and U2408 (N_2408,N_2207,N_2365);
and U2409 (N_2409,N_2313,N_2399);
or U2410 (N_2410,N_2251,N_2328);
or U2411 (N_2411,N_2318,N_2302);
or U2412 (N_2412,N_2264,N_2224);
nor U2413 (N_2413,N_2258,N_2368);
and U2414 (N_2414,N_2321,N_2378);
nor U2415 (N_2415,N_2351,N_2303);
nand U2416 (N_2416,N_2268,N_2291);
nand U2417 (N_2417,N_2263,N_2294);
and U2418 (N_2418,N_2228,N_2307);
nand U2419 (N_2419,N_2398,N_2246);
or U2420 (N_2420,N_2359,N_2211);
or U2421 (N_2421,N_2225,N_2297);
nand U2422 (N_2422,N_2308,N_2248);
nand U2423 (N_2423,N_2327,N_2395);
or U2424 (N_2424,N_2240,N_2227);
xor U2425 (N_2425,N_2366,N_2338);
and U2426 (N_2426,N_2386,N_2316);
nor U2427 (N_2427,N_2319,N_2220);
xnor U2428 (N_2428,N_2323,N_2341);
and U2429 (N_2429,N_2340,N_2262);
or U2430 (N_2430,N_2377,N_2234);
xor U2431 (N_2431,N_2279,N_2272);
or U2432 (N_2432,N_2216,N_2210);
nand U2433 (N_2433,N_2285,N_2371);
nor U2434 (N_2434,N_2283,N_2310);
or U2435 (N_2435,N_2353,N_2286);
nor U2436 (N_2436,N_2202,N_2201);
xnor U2437 (N_2437,N_2244,N_2293);
or U2438 (N_2438,N_2345,N_2332);
or U2439 (N_2439,N_2253,N_2325);
or U2440 (N_2440,N_2363,N_2273);
nor U2441 (N_2441,N_2288,N_2339);
xnor U2442 (N_2442,N_2396,N_2370);
and U2443 (N_2443,N_2255,N_2280);
or U2444 (N_2444,N_2229,N_2367);
and U2445 (N_2445,N_2320,N_2343);
and U2446 (N_2446,N_2349,N_2333);
nand U2447 (N_2447,N_2375,N_2311);
or U2448 (N_2448,N_2267,N_2394);
and U2449 (N_2449,N_2239,N_2296);
xnor U2450 (N_2450,N_2206,N_2250);
or U2451 (N_2451,N_2204,N_2300);
nor U2452 (N_2452,N_2236,N_2282);
nor U2453 (N_2453,N_2237,N_2223);
nand U2454 (N_2454,N_2221,N_2231);
or U2455 (N_2455,N_2298,N_2241);
or U2456 (N_2456,N_2350,N_2352);
nor U2457 (N_2457,N_2299,N_2215);
or U2458 (N_2458,N_2360,N_2392);
or U2459 (N_2459,N_2379,N_2329);
nand U2460 (N_2460,N_2274,N_2362);
or U2461 (N_2461,N_2304,N_2346);
and U2462 (N_2462,N_2257,N_2380);
and U2463 (N_2463,N_2301,N_2306);
xor U2464 (N_2464,N_2393,N_2390);
nand U2465 (N_2465,N_2374,N_2347);
and U2466 (N_2466,N_2256,N_2200);
or U2467 (N_2467,N_2335,N_2383);
xor U2468 (N_2468,N_2322,N_2259);
nand U2469 (N_2469,N_2348,N_2287);
xnor U2470 (N_2470,N_2203,N_2249);
nor U2471 (N_2471,N_2269,N_2226);
or U2472 (N_2472,N_2385,N_2252);
or U2473 (N_2473,N_2372,N_2364);
nor U2474 (N_2474,N_2369,N_2361);
xor U2475 (N_2475,N_2337,N_2315);
nor U2476 (N_2476,N_2376,N_2270);
xor U2477 (N_2477,N_2342,N_2289);
and U2478 (N_2478,N_2242,N_2358);
nand U2479 (N_2479,N_2275,N_2357);
nand U2480 (N_2480,N_2381,N_2235);
xnor U2481 (N_2481,N_2312,N_2336);
or U2482 (N_2482,N_2261,N_2233);
or U2483 (N_2483,N_2397,N_2205);
nand U2484 (N_2484,N_2324,N_2247);
or U2485 (N_2485,N_2238,N_2281);
or U2486 (N_2486,N_2356,N_2384);
or U2487 (N_2487,N_2277,N_2388);
or U2488 (N_2488,N_2271,N_2230);
nand U2489 (N_2489,N_2389,N_2219);
nor U2490 (N_2490,N_2344,N_2217);
xnor U2491 (N_2491,N_2243,N_2284);
or U2492 (N_2492,N_2232,N_2382);
and U2493 (N_2493,N_2309,N_2222);
and U2494 (N_2494,N_2330,N_2295);
or U2495 (N_2495,N_2209,N_2326);
xnor U2496 (N_2496,N_2265,N_2213);
or U2497 (N_2497,N_2317,N_2278);
and U2498 (N_2498,N_2314,N_2373);
and U2499 (N_2499,N_2276,N_2305);
or U2500 (N_2500,N_2383,N_2312);
xor U2501 (N_2501,N_2251,N_2243);
nor U2502 (N_2502,N_2385,N_2319);
nor U2503 (N_2503,N_2358,N_2338);
xnor U2504 (N_2504,N_2354,N_2246);
nand U2505 (N_2505,N_2357,N_2203);
nor U2506 (N_2506,N_2263,N_2239);
or U2507 (N_2507,N_2201,N_2367);
nor U2508 (N_2508,N_2332,N_2352);
nor U2509 (N_2509,N_2298,N_2348);
nand U2510 (N_2510,N_2372,N_2227);
or U2511 (N_2511,N_2294,N_2320);
and U2512 (N_2512,N_2327,N_2398);
or U2513 (N_2513,N_2350,N_2376);
and U2514 (N_2514,N_2240,N_2318);
nand U2515 (N_2515,N_2241,N_2356);
or U2516 (N_2516,N_2316,N_2269);
and U2517 (N_2517,N_2262,N_2344);
or U2518 (N_2518,N_2319,N_2350);
or U2519 (N_2519,N_2251,N_2228);
or U2520 (N_2520,N_2307,N_2292);
xnor U2521 (N_2521,N_2248,N_2296);
xor U2522 (N_2522,N_2220,N_2390);
nor U2523 (N_2523,N_2366,N_2247);
nand U2524 (N_2524,N_2393,N_2259);
nand U2525 (N_2525,N_2279,N_2268);
and U2526 (N_2526,N_2365,N_2369);
or U2527 (N_2527,N_2358,N_2306);
xor U2528 (N_2528,N_2322,N_2275);
xor U2529 (N_2529,N_2268,N_2344);
nor U2530 (N_2530,N_2289,N_2236);
nor U2531 (N_2531,N_2334,N_2305);
nor U2532 (N_2532,N_2394,N_2295);
nor U2533 (N_2533,N_2213,N_2349);
nand U2534 (N_2534,N_2201,N_2374);
nor U2535 (N_2535,N_2304,N_2305);
and U2536 (N_2536,N_2318,N_2207);
nor U2537 (N_2537,N_2362,N_2319);
or U2538 (N_2538,N_2329,N_2215);
and U2539 (N_2539,N_2258,N_2309);
nor U2540 (N_2540,N_2210,N_2272);
nand U2541 (N_2541,N_2366,N_2226);
nand U2542 (N_2542,N_2359,N_2310);
xnor U2543 (N_2543,N_2219,N_2354);
nor U2544 (N_2544,N_2225,N_2303);
nor U2545 (N_2545,N_2360,N_2372);
xor U2546 (N_2546,N_2356,N_2281);
or U2547 (N_2547,N_2218,N_2353);
xnor U2548 (N_2548,N_2301,N_2292);
and U2549 (N_2549,N_2381,N_2221);
nand U2550 (N_2550,N_2250,N_2249);
and U2551 (N_2551,N_2237,N_2391);
xor U2552 (N_2552,N_2277,N_2317);
xnor U2553 (N_2553,N_2322,N_2226);
xnor U2554 (N_2554,N_2292,N_2263);
and U2555 (N_2555,N_2279,N_2358);
nor U2556 (N_2556,N_2286,N_2327);
nand U2557 (N_2557,N_2271,N_2258);
and U2558 (N_2558,N_2357,N_2322);
xor U2559 (N_2559,N_2299,N_2303);
nand U2560 (N_2560,N_2325,N_2294);
nand U2561 (N_2561,N_2293,N_2394);
or U2562 (N_2562,N_2355,N_2390);
xor U2563 (N_2563,N_2348,N_2296);
or U2564 (N_2564,N_2242,N_2350);
nand U2565 (N_2565,N_2300,N_2344);
nor U2566 (N_2566,N_2314,N_2246);
nand U2567 (N_2567,N_2267,N_2232);
nor U2568 (N_2568,N_2260,N_2275);
and U2569 (N_2569,N_2227,N_2327);
or U2570 (N_2570,N_2266,N_2334);
xor U2571 (N_2571,N_2367,N_2381);
or U2572 (N_2572,N_2329,N_2299);
xnor U2573 (N_2573,N_2299,N_2346);
or U2574 (N_2574,N_2276,N_2336);
or U2575 (N_2575,N_2261,N_2313);
nand U2576 (N_2576,N_2262,N_2252);
nand U2577 (N_2577,N_2213,N_2252);
nand U2578 (N_2578,N_2262,N_2236);
xnor U2579 (N_2579,N_2331,N_2283);
or U2580 (N_2580,N_2369,N_2313);
xor U2581 (N_2581,N_2270,N_2285);
nor U2582 (N_2582,N_2298,N_2364);
and U2583 (N_2583,N_2333,N_2256);
and U2584 (N_2584,N_2287,N_2321);
or U2585 (N_2585,N_2386,N_2339);
or U2586 (N_2586,N_2237,N_2215);
xnor U2587 (N_2587,N_2288,N_2340);
nand U2588 (N_2588,N_2213,N_2390);
nor U2589 (N_2589,N_2238,N_2253);
nand U2590 (N_2590,N_2321,N_2296);
or U2591 (N_2591,N_2201,N_2350);
nand U2592 (N_2592,N_2334,N_2273);
or U2593 (N_2593,N_2338,N_2319);
xnor U2594 (N_2594,N_2381,N_2270);
or U2595 (N_2595,N_2389,N_2322);
nand U2596 (N_2596,N_2339,N_2307);
nand U2597 (N_2597,N_2255,N_2251);
and U2598 (N_2598,N_2205,N_2231);
xor U2599 (N_2599,N_2299,N_2240);
nand U2600 (N_2600,N_2563,N_2427);
xnor U2601 (N_2601,N_2430,N_2418);
nor U2602 (N_2602,N_2540,N_2595);
nand U2603 (N_2603,N_2508,N_2484);
nor U2604 (N_2604,N_2501,N_2436);
and U2605 (N_2605,N_2528,N_2476);
nor U2606 (N_2606,N_2471,N_2575);
nand U2607 (N_2607,N_2470,N_2521);
nor U2608 (N_2608,N_2593,N_2530);
nor U2609 (N_2609,N_2583,N_2455);
or U2610 (N_2610,N_2475,N_2569);
or U2611 (N_2611,N_2532,N_2465);
and U2612 (N_2612,N_2485,N_2535);
xor U2613 (N_2613,N_2545,N_2403);
nand U2614 (N_2614,N_2558,N_2454);
xnor U2615 (N_2615,N_2510,N_2522);
nand U2616 (N_2616,N_2462,N_2426);
and U2617 (N_2617,N_2445,N_2442);
nor U2618 (N_2618,N_2498,N_2513);
and U2619 (N_2619,N_2585,N_2481);
nand U2620 (N_2620,N_2538,N_2495);
nor U2621 (N_2621,N_2568,N_2435);
or U2622 (N_2622,N_2460,N_2416);
or U2623 (N_2623,N_2429,N_2443);
xor U2624 (N_2624,N_2556,N_2401);
xor U2625 (N_2625,N_2587,N_2577);
nand U2626 (N_2626,N_2467,N_2597);
and U2627 (N_2627,N_2449,N_2591);
nor U2628 (N_2628,N_2448,N_2490);
or U2629 (N_2629,N_2567,N_2534);
xnor U2630 (N_2630,N_2419,N_2548);
xor U2631 (N_2631,N_2566,N_2497);
and U2632 (N_2632,N_2555,N_2482);
nand U2633 (N_2633,N_2573,N_2584);
nand U2634 (N_2634,N_2493,N_2526);
xor U2635 (N_2635,N_2542,N_2564);
nor U2636 (N_2636,N_2589,N_2486);
nor U2637 (N_2637,N_2405,N_2433);
nand U2638 (N_2638,N_2415,N_2507);
nand U2639 (N_2639,N_2483,N_2414);
or U2640 (N_2640,N_2421,N_2447);
nor U2641 (N_2641,N_2547,N_2459);
nand U2642 (N_2642,N_2588,N_2565);
nor U2643 (N_2643,N_2599,N_2582);
or U2644 (N_2644,N_2503,N_2516);
nor U2645 (N_2645,N_2524,N_2514);
nand U2646 (N_2646,N_2425,N_2472);
nor U2647 (N_2647,N_2550,N_2559);
or U2648 (N_2648,N_2438,N_2519);
or U2649 (N_2649,N_2408,N_2473);
or U2650 (N_2650,N_2413,N_2463);
or U2651 (N_2651,N_2404,N_2432);
xnor U2652 (N_2652,N_2543,N_2505);
and U2653 (N_2653,N_2400,N_2451);
xnor U2654 (N_2654,N_2499,N_2504);
and U2655 (N_2655,N_2491,N_2596);
or U2656 (N_2656,N_2598,N_2488);
xor U2657 (N_2657,N_2494,N_2478);
and U2658 (N_2658,N_2456,N_2512);
nand U2659 (N_2659,N_2431,N_2544);
or U2660 (N_2660,N_2411,N_2571);
nor U2661 (N_2661,N_2517,N_2511);
xnor U2662 (N_2662,N_2402,N_2580);
nand U2663 (N_2663,N_2492,N_2434);
nor U2664 (N_2664,N_2529,N_2424);
and U2665 (N_2665,N_2592,N_2464);
xnor U2666 (N_2666,N_2572,N_2553);
and U2667 (N_2667,N_2506,N_2515);
nor U2668 (N_2668,N_2446,N_2537);
xnor U2669 (N_2669,N_2581,N_2458);
or U2670 (N_2670,N_2509,N_2574);
nor U2671 (N_2671,N_2496,N_2439);
xnor U2672 (N_2672,N_2461,N_2502);
nor U2673 (N_2673,N_2546,N_2477);
or U2674 (N_2674,N_2560,N_2487);
and U2675 (N_2675,N_2578,N_2410);
or U2676 (N_2676,N_2406,N_2479);
nand U2677 (N_2677,N_2576,N_2453);
nand U2678 (N_2678,N_2452,N_2541);
nand U2679 (N_2679,N_2590,N_2579);
xnor U2680 (N_2680,N_2570,N_2586);
nand U2681 (N_2681,N_2480,N_2417);
and U2682 (N_2682,N_2466,N_2468);
and U2683 (N_2683,N_2551,N_2428);
xor U2684 (N_2684,N_2420,N_2554);
nor U2685 (N_2685,N_2423,N_2562);
xnor U2686 (N_2686,N_2552,N_2422);
and U2687 (N_2687,N_2489,N_2539);
nor U2688 (N_2688,N_2444,N_2500);
nor U2689 (N_2689,N_2474,N_2594);
or U2690 (N_2690,N_2412,N_2525);
nor U2691 (N_2691,N_2437,N_2533);
and U2692 (N_2692,N_2536,N_2531);
nor U2693 (N_2693,N_2469,N_2409);
nand U2694 (N_2694,N_2450,N_2441);
or U2695 (N_2695,N_2520,N_2440);
or U2696 (N_2696,N_2549,N_2518);
and U2697 (N_2697,N_2523,N_2557);
nand U2698 (N_2698,N_2527,N_2407);
or U2699 (N_2699,N_2561,N_2457);
or U2700 (N_2700,N_2408,N_2598);
and U2701 (N_2701,N_2526,N_2566);
nand U2702 (N_2702,N_2515,N_2421);
xnor U2703 (N_2703,N_2504,N_2533);
xnor U2704 (N_2704,N_2479,N_2495);
nand U2705 (N_2705,N_2557,N_2471);
nor U2706 (N_2706,N_2491,N_2487);
nand U2707 (N_2707,N_2568,N_2473);
and U2708 (N_2708,N_2511,N_2569);
or U2709 (N_2709,N_2581,N_2536);
or U2710 (N_2710,N_2507,N_2538);
and U2711 (N_2711,N_2404,N_2532);
nand U2712 (N_2712,N_2581,N_2582);
nor U2713 (N_2713,N_2545,N_2406);
or U2714 (N_2714,N_2542,N_2532);
nand U2715 (N_2715,N_2531,N_2573);
nor U2716 (N_2716,N_2527,N_2532);
and U2717 (N_2717,N_2517,N_2451);
nor U2718 (N_2718,N_2524,N_2523);
and U2719 (N_2719,N_2538,N_2450);
xnor U2720 (N_2720,N_2556,N_2515);
and U2721 (N_2721,N_2522,N_2491);
xor U2722 (N_2722,N_2514,N_2489);
xnor U2723 (N_2723,N_2509,N_2422);
or U2724 (N_2724,N_2440,N_2582);
xnor U2725 (N_2725,N_2539,N_2583);
nor U2726 (N_2726,N_2454,N_2409);
nor U2727 (N_2727,N_2594,N_2498);
xor U2728 (N_2728,N_2592,N_2537);
or U2729 (N_2729,N_2472,N_2481);
xor U2730 (N_2730,N_2587,N_2417);
xnor U2731 (N_2731,N_2487,N_2430);
or U2732 (N_2732,N_2532,N_2515);
xnor U2733 (N_2733,N_2596,N_2472);
nor U2734 (N_2734,N_2518,N_2559);
xor U2735 (N_2735,N_2553,N_2462);
nand U2736 (N_2736,N_2422,N_2429);
nor U2737 (N_2737,N_2487,N_2591);
nand U2738 (N_2738,N_2586,N_2535);
or U2739 (N_2739,N_2445,N_2428);
nand U2740 (N_2740,N_2579,N_2403);
nand U2741 (N_2741,N_2597,N_2526);
nand U2742 (N_2742,N_2404,N_2579);
nand U2743 (N_2743,N_2558,N_2570);
and U2744 (N_2744,N_2529,N_2557);
and U2745 (N_2745,N_2513,N_2545);
xnor U2746 (N_2746,N_2518,N_2453);
xnor U2747 (N_2747,N_2595,N_2567);
nand U2748 (N_2748,N_2563,N_2453);
xor U2749 (N_2749,N_2452,N_2489);
nand U2750 (N_2750,N_2516,N_2403);
nand U2751 (N_2751,N_2440,N_2491);
and U2752 (N_2752,N_2550,N_2599);
xor U2753 (N_2753,N_2517,N_2558);
nor U2754 (N_2754,N_2537,N_2522);
nor U2755 (N_2755,N_2553,N_2559);
and U2756 (N_2756,N_2497,N_2531);
nor U2757 (N_2757,N_2416,N_2433);
nor U2758 (N_2758,N_2530,N_2406);
or U2759 (N_2759,N_2419,N_2555);
and U2760 (N_2760,N_2545,N_2445);
or U2761 (N_2761,N_2403,N_2497);
or U2762 (N_2762,N_2427,N_2576);
and U2763 (N_2763,N_2403,N_2520);
and U2764 (N_2764,N_2447,N_2581);
or U2765 (N_2765,N_2402,N_2424);
nand U2766 (N_2766,N_2422,N_2570);
and U2767 (N_2767,N_2572,N_2449);
and U2768 (N_2768,N_2513,N_2456);
or U2769 (N_2769,N_2485,N_2548);
and U2770 (N_2770,N_2491,N_2526);
and U2771 (N_2771,N_2401,N_2420);
xnor U2772 (N_2772,N_2500,N_2475);
xor U2773 (N_2773,N_2464,N_2578);
nand U2774 (N_2774,N_2432,N_2591);
nor U2775 (N_2775,N_2438,N_2472);
and U2776 (N_2776,N_2523,N_2491);
and U2777 (N_2777,N_2549,N_2516);
xor U2778 (N_2778,N_2568,N_2475);
nor U2779 (N_2779,N_2485,N_2539);
nor U2780 (N_2780,N_2444,N_2498);
or U2781 (N_2781,N_2436,N_2467);
nor U2782 (N_2782,N_2483,N_2423);
or U2783 (N_2783,N_2559,N_2513);
nor U2784 (N_2784,N_2594,N_2491);
xor U2785 (N_2785,N_2443,N_2565);
nor U2786 (N_2786,N_2539,N_2441);
xnor U2787 (N_2787,N_2531,N_2455);
xor U2788 (N_2788,N_2528,N_2416);
xnor U2789 (N_2789,N_2425,N_2585);
nand U2790 (N_2790,N_2435,N_2580);
nor U2791 (N_2791,N_2477,N_2557);
nand U2792 (N_2792,N_2454,N_2435);
or U2793 (N_2793,N_2536,N_2543);
xor U2794 (N_2794,N_2553,N_2451);
nor U2795 (N_2795,N_2546,N_2443);
or U2796 (N_2796,N_2503,N_2402);
nor U2797 (N_2797,N_2483,N_2502);
or U2798 (N_2798,N_2563,N_2401);
nand U2799 (N_2799,N_2547,N_2534);
xor U2800 (N_2800,N_2786,N_2657);
and U2801 (N_2801,N_2754,N_2621);
or U2802 (N_2802,N_2662,N_2681);
nand U2803 (N_2803,N_2654,N_2640);
and U2804 (N_2804,N_2726,N_2706);
xnor U2805 (N_2805,N_2620,N_2610);
nand U2806 (N_2806,N_2724,N_2729);
nand U2807 (N_2807,N_2650,N_2787);
nor U2808 (N_2808,N_2735,N_2617);
nor U2809 (N_2809,N_2635,N_2698);
or U2810 (N_2810,N_2741,N_2601);
xor U2811 (N_2811,N_2661,N_2694);
xnor U2812 (N_2812,N_2765,N_2695);
and U2813 (N_2813,N_2634,N_2710);
or U2814 (N_2814,N_2779,N_2714);
nor U2815 (N_2815,N_2728,N_2700);
nand U2816 (N_2816,N_2623,N_2675);
or U2817 (N_2817,N_2774,N_2701);
or U2818 (N_2818,N_2684,N_2709);
or U2819 (N_2819,N_2749,N_2782);
nand U2820 (N_2820,N_2707,N_2771);
and U2821 (N_2821,N_2730,N_2781);
xnor U2822 (N_2822,N_2615,N_2719);
or U2823 (N_2823,N_2685,N_2751);
xnor U2824 (N_2824,N_2680,N_2705);
and U2825 (N_2825,N_2792,N_2677);
or U2826 (N_2826,N_2733,N_2718);
xnor U2827 (N_2827,N_2666,N_2644);
and U2828 (N_2828,N_2760,N_2699);
or U2829 (N_2829,N_2756,N_2772);
and U2830 (N_2830,N_2607,N_2626);
nand U2831 (N_2831,N_2778,N_2748);
and U2832 (N_2832,N_2618,N_2664);
and U2833 (N_2833,N_2750,N_2791);
xor U2834 (N_2834,N_2630,N_2723);
or U2835 (N_2835,N_2627,N_2720);
nand U2836 (N_2836,N_2788,N_2638);
nand U2837 (N_2837,N_2777,N_2672);
nand U2838 (N_2838,N_2674,N_2797);
and U2839 (N_2839,N_2757,N_2682);
nand U2840 (N_2840,N_2648,N_2688);
and U2841 (N_2841,N_2746,N_2667);
and U2842 (N_2842,N_2651,N_2708);
nor U2843 (N_2843,N_2670,N_2646);
xnor U2844 (N_2844,N_2637,N_2609);
or U2845 (N_2845,N_2669,N_2704);
and U2846 (N_2846,N_2776,N_2734);
xnor U2847 (N_2847,N_2612,N_2783);
and U2848 (N_2848,N_2668,N_2613);
and U2849 (N_2849,N_2737,N_2702);
and U2850 (N_2850,N_2636,N_2736);
nand U2851 (N_2851,N_2649,N_2799);
nand U2852 (N_2852,N_2652,N_2602);
nand U2853 (N_2853,N_2686,N_2608);
and U2854 (N_2854,N_2656,N_2606);
and U2855 (N_2855,N_2732,N_2773);
nand U2856 (N_2856,N_2611,N_2780);
nand U2857 (N_2857,N_2691,N_2796);
nor U2858 (N_2858,N_2696,N_2747);
or U2859 (N_2859,N_2614,N_2716);
nor U2860 (N_2860,N_2671,N_2655);
nand U2861 (N_2861,N_2717,N_2761);
nor U2862 (N_2862,N_2790,N_2763);
nor U2863 (N_2863,N_2766,N_2703);
xor U2864 (N_2864,N_2647,N_2762);
xor U2865 (N_2865,N_2693,N_2769);
and U2866 (N_2866,N_2738,N_2753);
or U2867 (N_2867,N_2755,N_2663);
and U2868 (N_2868,N_2628,N_2785);
nand U2869 (N_2869,N_2624,N_2795);
xnor U2870 (N_2870,N_2744,N_2764);
nor U2871 (N_2871,N_2740,N_2616);
or U2872 (N_2872,N_2659,N_2793);
or U2873 (N_2873,N_2784,N_2633);
nor U2874 (N_2874,N_2619,N_2689);
xor U2875 (N_2875,N_2711,N_2742);
xnor U2876 (N_2876,N_2789,N_2745);
nor U2877 (N_2877,N_2722,N_2758);
and U2878 (N_2878,N_2660,N_2631);
or U2879 (N_2879,N_2770,N_2697);
and U2880 (N_2880,N_2605,N_2687);
nand U2881 (N_2881,N_2676,N_2645);
or U2882 (N_2882,N_2768,N_2798);
xnor U2883 (N_2883,N_2658,N_2604);
or U2884 (N_2884,N_2673,N_2622);
and U2885 (N_2885,N_2679,N_2632);
or U2886 (N_2886,N_2683,N_2712);
nor U2887 (N_2887,N_2759,N_2642);
nor U2888 (N_2888,N_2625,N_2678);
and U2889 (N_2889,N_2725,N_2692);
and U2890 (N_2890,N_2629,N_2690);
xor U2891 (N_2891,N_2739,N_2775);
or U2892 (N_2892,N_2665,N_2767);
and U2893 (N_2893,N_2653,N_2752);
nor U2894 (N_2894,N_2639,N_2643);
nand U2895 (N_2895,N_2727,N_2743);
and U2896 (N_2896,N_2715,N_2603);
and U2897 (N_2897,N_2794,N_2600);
nor U2898 (N_2898,N_2713,N_2641);
xnor U2899 (N_2899,N_2721,N_2731);
nand U2900 (N_2900,N_2798,N_2647);
or U2901 (N_2901,N_2776,N_2675);
nand U2902 (N_2902,N_2606,N_2675);
xnor U2903 (N_2903,N_2665,N_2685);
xor U2904 (N_2904,N_2605,N_2773);
nor U2905 (N_2905,N_2649,N_2783);
nor U2906 (N_2906,N_2690,N_2754);
xnor U2907 (N_2907,N_2735,N_2776);
nor U2908 (N_2908,N_2776,N_2778);
or U2909 (N_2909,N_2744,N_2628);
xnor U2910 (N_2910,N_2760,N_2784);
xnor U2911 (N_2911,N_2749,N_2769);
and U2912 (N_2912,N_2691,N_2683);
nor U2913 (N_2913,N_2675,N_2750);
nor U2914 (N_2914,N_2725,N_2697);
nor U2915 (N_2915,N_2758,N_2669);
xor U2916 (N_2916,N_2755,N_2677);
or U2917 (N_2917,N_2775,N_2793);
and U2918 (N_2918,N_2675,N_2759);
and U2919 (N_2919,N_2619,N_2620);
or U2920 (N_2920,N_2703,N_2742);
nand U2921 (N_2921,N_2616,N_2693);
or U2922 (N_2922,N_2729,N_2681);
xor U2923 (N_2923,N_2612,N_2698);
or U2924 (N_2924,N_2662,N_2790);
or U2925 (N_2925,N_2714,N_2621);
nor U2926 (N_2926,N_2725,N_2780);
or U2927 (N_2927,N_2701,N_2779);
nand U2928 (N_2928,N_2684,N_2788);
xor U2929 (N_2929,N_2659,N_2615);
and U2930 (N_2930,N_2762,N_2756);
or U2931 (N_2931,N_2724,N_2703);
nand U2932 (N_2932,N_2603,N_2725);
nor U2933 (N_2933,N_2761,N_2766);
and U2934 (N_2934,N_2749,N_2750);
nand U2935 (N_2935,N_2659,N_2640);
and U2936 (N_2936,N_2624,N_2788);
nand U2937 (N_2937,N_2677,N_2669);
nor U2938 (N_2938,N_2711,N_2745);
nor U2939 (N_2939,N_2633,N_2751);
and U2940 (N_2940,N_2691,N_2752);
and U2941 (N_2941,N_2686,N_2657);
nand U2942 (N_2942,N_2755,N_2701);
nand U2943 (N_2943,N_2661,N_2793);
and U2944 (N_2944,N_2760,N_2609);
nor U2945 (N_2945,N_2720,N_2668);
or U2946 (N_2946,N_2659,N_2671);
nand U2947 (N_2947,N_2643,N_2733);
or U2948 (N_2948,N_2734,N_2729);
xnor U2949 (N_2949,N_2636,N_2713);
and U2950 (N_2950,N_2658,N_2673);
xnor U2951 (N_2951,N_2759,N_2653);
nor U2952 (N_2952,N_2782,N_2605);
xnor U2953 (N_2953,N_2685,N_2730);
and U2954 (N_2954,N_2748,N_2615);
xor U2955 (N_2955,N_2712,N_2772);
nand U2956 (N_2956,N_2637,N_2658);
and U2957 (N_2957,N_2635,N_2715);
nand U2958 (N_2958,N_2721,N_2660);
and U2959 (N_2959,N_2757,N_2705);
xor U2960 (N_2960,N_2771,N_2723);
nor U2961 (N_2961,N_2728,N_2701);
xor U2962 (N_2962,N_2611,N_2685);
or U2963 (N_2963,N_2601,N_2734);
nand U2964 (N_2964,N_2745,N_2782);
nand U2965 (N_2965,N_2601,N_2698);
or U2966 (N_2966,N_2630,N_2604);
xnor U2967 (N_2967,N_2708,N_2611);
and U2968 (N_2968,N_2709,N_2678);
or U2969 (N_2969,N_2676,N_2762);
or U2970 (N_2970,N_2771,N_2746);
and U2971 (N_2971,N_2651,N_2672);
nand U2972 (N_2972,N_2673,N_2706);
and U2973 (N_2973,N_2660,N_2768);
or U2974 (N_2974,N_2682,N_2787);
and U2975 (N_2975,N_2779,N_2742);
and U2976 (N_2976,N_2665,N_2622);
nor U2977 (N_2977,N_2694,N_2602);
nor U2978 (N_2978,N_2744,N_2784);
nor U2979 (N_2979,N_2761,N_2728);
nor U2980 (N_2980,N_2685,N_2612);
or U2981 (N_2981,N_2767,N_2752);
nor U2982 (N_2982,N_2761,N_2656);
nand U2983 (N_2983,N_2728,N_2683);
nand U2984 (N_2984,N_2709,N_2794);
xnor U2985 (N_2985,N_2631,N_2718);
or U2986 (N_2986,N_2737,N_2731);
nor U2987 (N_2987,N_2672,N_2683);
xor U2988 (N_2988,N_2662,N_2718);
xor U2989 (N_2989,N_2685,N_2723);
or U2990 (N_2990,N_2659,N_2644);
or U2991 (N_2991,N_2660,N_2640);
nor U2992 (N_2992,N_2699,N_2626);
or U2993 (N_2993,N_2660,N_2678);
and U2994 (N_2994,N_2746,N_2679);
xnor U2995 (N_2995,N_2706,N_2779);
and U2996 (N_2996,N_2778,N_2688);
and U2997 (N_2997,N_2659,N_2601);
or U2998 (N_2998,N_2737,N_2793);
nor U2999 (N_2999,N_2781,N_2634);
nand U3000 (N_3000,N_2821,N_2875);
nand U3001 (N_3001,N_2996,N_2911);
xnor U3002 (N_3002,N_2814,N_2833);
or U3003 (N_3003,N_2829,N_2981);
or U3004 (N_3004,N_2809,N_2824);
nand U3005 (N_3005,N_2820,N_2985);
xnor U3006 (N_3006,N_2927,N_2853);
nor U3007 (N_3007,N_2825,N_2885);
or U3008 (N_3008,N_2858,N_2913);
xnor U3009 (N_3009,N_2977,N_2940);
or U3010 (N_3010,N_2964,N_2871);
and U3011 (N_3011,N_2992,N_2854);
xor U3012 (N_3012,N_2950,N_2863);
nor U3013 (N_3013,N_2961,N_2883);
nand U3014 (N_3014,N_2906,N_2966);
and U3015 (N_3015,N_2801,N_2956);
or U3016 (N_3016,N_2969,N_2962);
and U3017 (N_3017,N_2840,N_2959);
and U3018 (N_3018,N_2953,N_2932);
xnor U3019 (N_3019,N_2846,N_2915);
or U3020 (N_3020,N_2997,N_2931);
and U3021 (N_3021,N_2974,N_2888);
or U3022 (N_3022,N_2910,N_2847);
nand U3023 (N_3023,N_2816,N_2984);
or U3024 (N_3024,N_2803,N_2946);
nand U3025 (N_3025,N_2819,N_2861);
or U3026 (N_3026,N_2860,N_2952);
xnor U3027 (N_3027,N_2926,N_2935);
nor U3028 (N_3028,N_2949,N_2893);
and U3029 (N_3029,N_2999,N_2866);
and U3030 (N_3030,N_2934,N_2830);
or U3031 (N_3031,N_2806,N_2876);
xor U3032 (N_3032,N_2900,N_2813);
and U3033 (N_3033,N_2912,N_2972);
and U3034 (N_3034,N_2933,N_2901);
nand U3035 (N_3035,N_2898,N_2874);
nand U3036 (N_3036,N_2957,N_2832);
and U3037 (N_3037,N_2988,N_2823);
nor U3038 (N_3038,N_2839,N_2842);
and U3039 (N_3039,N_2802,N_2945);
or U3040 (N_3040,N_2845,N_2978);
xnor U3041 (N_3041,N_2947,N_2890);
xnor U3042 (N_3042,N_2834,N_2908);
nand U3043 (N_3043,N_2921,N_2818);
and U3044 (N_3044,N_2887,N_2835);
or U3045 (N_3045,N_2980,N_2852);
and U3046 (N_3046,N_2810,N_2919);
xor U3047 (N_3047,N_2936,N_2800);
nand U3048 (N_3048,N_2951,N_2944);
xor U3049 (N_3049,N_2862,N_2827);
xnor U3050 (N_3050,N_2897,N_2937);
xnor U3051 (N_3051,N_2889,N_2841);
nand U3052 (N_3052,N_2989,N_2994);
or U3053 (N_3053,N_2867,N_2916);
nand U3054 (N_3054,N_2987,N_2879);
nand U3055 (N_3055,N_2877,N_2983);
nor U3056 (N_3056,N_2836,N_2998);
or U3057 (N_3057,N_2902,N_2857);
or U3058 (N_3058,N_2865,N_2975);
nand U3059 (N_3059,N_2955,N_2870);
or U3060 (N_3060,N_2849,N_2923);
xor U3061 (N_3061,N_2864,N_2873);
or U3062 (N_3062,N_2943,N_2848);
nand U3063 (N_3063,N_2914,N_2963);
nand U3064 (N_3064,N_2850,N_2986);
nand U3065 (N_3065,N_2941,N_2807);
or U3066 (N_3066,N_2884,N_2811);
xor U3067 (N_3067,N_2880,N_2970);
and U3068 (N_3068,N_2979,N_2881);
nor U3069 (N_3069,N_2817,N_2907);
or U3070 (N_3070,N_2918,N_2922);
and U3071 (N_3071,N_2899,N_2868);
nand U3072 (N_3072,N_2929,N_2822);
nor U3073 (N_3073,N_2928,N_2990);
nand U3074 (N_3074,N_2973,N_2804);
nand U3075 (N_3075,N_2925,N_2882);
nor U3076 (N_3076,N_2917,N_2942);
nor U3077 (N_3077,N_2831,N_2924);
and U3078 (N_3078,N_2920,N_2948);
nand U3079 (N_3079,N_2903,N_2844);
and U3080 (N_3080,N_2826,N_2968);
and U3081 (N_3081,N_2895,N_2894);
nor U3082 (N_3082,N_2958,N_2967);
nor U3083 (N_3083,N_2991,N_2859);
nand U3084 (N_3084,N_2938,N_2869);
or U3085 (N_3085,N_2904,N_2965);
and U3086 (N_3086,N_2878,N_2843);
xor U3087 (N_3087,N_2930,N_2851);
and U3088 (N_3088,N_2954,N_2856);
nand U3089 (N_3089,N_2808,N_2828);
nor U3090 (N_3090,N_2939,N_2892);
nand U3091 (N_3091,N_2812,N_2855);
and U3092 (N_3092,N_2995,N_2976);
or U3093 (N_3093,N_2837,N_2886);
xnor U3094 (N_3094,N_2909,N_2896);
or U3095 (N_3095,N_2905,N_2815);
or U3096 (N_3096,N_2960,N_2872);
nand U3097 (N_3097,N_2993,N_2971);
xnor U3098 (N_3098,N_2805,N_2891);
nor U3099 (N_3099,N_2982,N_2838);
nor U3100 (N_3100,N_2907,N_2923);
xnor U3101 (N_3101,N_2845,N_2826);
or U3102 (N_3102,N_2917,N_2947);
nor U3103 (N_3103,N_2880,N_2949);
nor U3104 (N_3104,N_2807,N_2902);
and U3105 (N_3105,N_2996,N_2973);
and U3106 (N_3106,N_2836,N_2913);
xor U3107 (N_3107,N_2881,N_2996);
and U3108 (N_3108,N_2986,N_2834);
or U3109 (N_3109,N_2984,N_2939);
and U3110 (N_3110,N_2837,N_2895);
nor U3111 (N_3111,N_2919,N_2966);
xnor U3112 (N_3112,N_2964,N_2905);
and U3113 (N_3113,N_2852,N_2960);
and U3114 (N_3114,N_2950,N_2888);
nor U3115 (N_3115,N_2830,N_2981);
or U3116 (N_3116,N_2917,N_2858);
nor U3117 (N_3117,N_2957,N_2803);
xor U3118 (N_3118,N_2861,N_2853);
nor U3119 (N_3119,N_2885,N_2935);
xnor U3120 (N_3120,N_2989,N_2930);
and U3121 (N_3121,N_2929,N_2827);
xor U3122 (N_3122,N_2832,N_2963);
or U3123 (N_3123,N_2868,N_2845);
xnor U3124 (N_3124,N_2975,N_2931);
nor U3125 (N_3125,N_2924,N_2817);
nand U3126 (N_3126,N_2824,N_2939);
or U3127 (N_3127,N_2871,N_2848);
and U3128 (N_3128,N_2961,N_2825);
nand U3129 (N_3129,N_2916,N_2850);
nand U3130 (N_3130,N_2965,N_2839);
or U3131 (N_3131,N_2830,N_2828);
nand U3132 (N_3132,N_2878,N_2906);
or U3133 (N_3133,N_2855,N_2892);
nand U3134 (N_3134,N_2918,N_2875);
or U3135 (N_3135,N_2836,N_2983);
xnor U3136 (N_3136,N_2869,N_2949);
and U3137 (N_3137,N_2805,N_2842);
and U3138 (N_3138,N_2948,N_2988);
nand U3139 (N_3139,N_2961,N_2840);
nand U3140 (N_3140,N_2962,N_2851);
nand U3141 (N_3141,N_2919,N_2816);
xnor U3142 (N_3142,N_2889,N_2947);
nor U3143 (N_3143,N_2807,N_2804);
and U3144 (N_3144,N_2889,N_2936);
or U3145 (N_3145,N_2872,N_2893);
and U3146 (N_3146,N_2874,N_2812);
and U3147 (N_3147,N_2945,N_2903);
nand U3148 (N_3148,N_2827,N_2945);
and U3149 (N_3149,N_2824,N_2811);
and U3150 (N_3150,N_2875,N_2925);
xnor U3151 (N_3151,N_2874,N_2978);
nand U3152 (N_3152,N_2947,N_2869);
or U3153 (N_3153,N_2841,N_2881);
nor U3154 (N_3154,N_2812,N_2809);
or U3155 (N_3155,N_2832,N_2916);
or U3156 (N_3156,N_2844,N_2976);
xor U3157 (N_3157,N_2933,N_2875);
or U3158 (N_3158,N_2894,N_2805);
xnor U3159 (N_3159,N_2917,N_2807);
and U3160 (N_3160,N_2987,N_2800);
nor U3161 (N_3161,N_2947,N_2831);
nor U3162 (N_3162,N_2847,N_2815);
xor U3163 (N_3163,N_2830,N_2876);
or U3164 (N_3164,N_2909,N_2834);
nand U3165 (N_3165,N_2919,N_2941);
nand U3166 (N_3166,N_2840,N_2882);
xnor U3167 (N_3167,N_2995,N_2890);
and U3168 (N_3168,N_2957,N_2901);
xnor U3169 (N_3169,N_2888,N_2832);
nor U3170 (N_3170,N_2905,N_2933);
nor U3171 (N_3171,N_2830,N_2945);
nand U3172 (N_3172,N_2922,N_2901);
and U3173 (N_3173,N_2847,N_2923);
nand U3174 (N_3174,N_2922,N_2844);
xnor U3175 (N_3175,N_2902,N_2912);
xor U3176 (N_3176,N_2875,N_2987);
or U3177 (N_3177,N_2984,N_2898);
and U3178 (N_3178,N_2842,N_2919);
xnor U3179 (N_3179,N_2827,N_2944);
and U3180 (N_3180,N_2968,N_2807);
xor U3181 (N_3181,N_2950,N_2919);
and U3182 (N_3182,N_2829,N_2928);
or U3183 (N_3183,N_2912,N_2830);
or U3184 (N_3184,N_2858,N_2947);
xnor U3185 (N_3185,N_2895,N_2964);
xnor U3186 (N_3186,N_2840,N_2973);
or U3187 (N_3187,N_2951,N_2803);
or U3188 (N_3188,N_2811,N_2932);
xnor U3189 (N_3189,N_2960,N_2966);
nand U3190 (N_3190,N_2998,N_2936);
xor U3191 (N_3191,N_2867,N_2902);
or U3192 (N_3192,N_2810,N_2860);
or U3193 (N_3193,N_2835,N_2864);
xnor U3194 (N_3194,N_2857,N_2937);
or U3195 (N_3195,N_2867,N_2963);
xor U3196 (N_3196,N_2975,N_2807);
or U3197 (N_3197,N_2836,N_2838);
nor U3198 (N_3198,N_2914,N_2999);
nand U3199 (N_3199,N_2863,N_2851);
nand U3200 (N_3200,N_3090,N_3020);
or U3201 (N_3201,N_3069,N_3171);
xnor U3202 (N_3202,N_3098,N_3093);
nor U3203 (N_3203,N_3148,N_3100);
nand U3204 (N_3204,N_3134,N_3008);
xnor U3205 (N_3205,N_3136,N_3092);
xor U3206 (N_3206,N_3183,N_3048);
nand U3207 (N_3207,N_3055,N_3094);
xor U3208 (N_3208,N_3182,N_3140);
nand U3209 (N_3209,N_3033,N_3066);
or U3210 (N_3210,N_3103,N_3119);
or U3211 (N_3211,N_3000,N_3147);
or U3212 (N_3212,N_3052,N_3190);
and U3213 (N_3213,N_3196,N_3101);
and U3214 (N_3214,N_3152,N_3081);
and U3215 (N_3215,N_3121,N_3029);
xnor U3216 (N_3216,N_3115,N_3145);
xnor U3217 (N_3217,N_3111,N_3001);
nand U3218 (N_3218,N_3120,N_3137);
or U3219 (N_3219,N_3022,N_3075);
and U3220 (N_3220,N_3072,N_3181);
nand U3221 (N_3221,N_3155,N_3021);
nor U3222 (N_3222,N_3080,N_3151);
nand U3223 (N_3223,N_3028,N_3025);
xnor U3224 (N_3224,N_3146,N_3161);
xnor U3225 (N_3225,N_3054,N_3178);
xor U3226 (N_3226,N_3009,N_3040);
nand U3227 (N_3227,N_3049,N_3032);
or U3228 (N_3228,N_3050,N_3014);
nor U3229 (N_3229,N_3010,N_3011);
and U3230 (N_3230,N_3106,N_3159);
nor U3231 (N_3231,N_3051,N_3174);
or U3232 (N_3232,N_3193,N_3061);
nor U3233 (N_3233,N_3097,N_3114);
nand U3234 (N_3234,N_3089,N_3086);
nor U3235 (N_3235,N_3124,N_3004);
and U3236 (N_3236,N_3150,N_3012);
or U3237 (N_3237,N_3199,N_3160);
and U3238 (N_3238,N_3179,N_3099);
or U3239 (N_3239,N_3044,N_3060);
xnor U3240 (N_3240,N_3068,N_3073);
and U3241 (N_3241,N_3059,N_3195);
nand U3242 (N_3242,N_3180,N_3118);
and U3243 (N_3243,N_3107,N_3041);
nor U3244 (N_3244,N_3085,N_3185);
nand U3245 (N_3245,N_3153,N_3053);
xor U3246 (N_3246,N_3168,N_3003);
nand U3247 (N_3247,N_3078,N_3194);
or U3248 (N_3248,N_3016,N_3113);
nor U3249 (N_3249,N_3125,N_3005);
or U3250 (N_3250,N_3177,N_3058);
xnor U3251 (N_3251,N_3074,N_3128);
or U3252 (N_3252,N_3141,N_3095);
or U3253 (N_3253,N_3042,N_3126);
or U3254 (N_3254,N_3176,N_3198);
nor U3255 (N_3255,N_3186,N_3175);
and U3256 (N_3256,N_3169,N_3036);
nor U3257 (N_3257,N_3139,N_3189);
and U3258 (N_3258,N_3144,N_3067);
and U3259 (N_3259,N_3065,N_3132);
xnor U3260 (N_3260,N_3027,N_3026);
or U3261 (N_3261,N_3019,N_3034);
nand U3262 (N_3262,N_3046,N_3015);
and U3263 (N_3263,N_3043,N_3082);
nand U3264 (N_3264,N_3064,N_3197);
nand U3265 (N_3265,N_3131,N_3117);
xnor U3266 (N_3266,N_3133,N_3087);
xor U3267 (N_3267,N_3123,N_3079);
and U3268 (N_3268,N_3023,N_3167);
nand U3269 (N_3269,N_3149,N_3156);
or U3270 (N_3270,N_3083,N_3035);
nor U3271 (N_3271,N_3007,N_3170);
xnor U3272 (N_3272,N_3091,N_3077);
xnor U3273 (N_3273,N_3138,N_3047);
xor U3274 (N_3274,N_3164,N_3102);
nand U3275 (N_3275,N_3030,N_3063);
nand U3276 (N_3276,N_3127,N_3129);
xor U3277 (N_3277,N_3096,N_3037);
nor U3278 (N_3278,N_3142,N_3112);
nand U3279 (N_3279,N_3122,N_3184);
nand U3280 (N_3280,N_3024,N_3088);
nor U3281 (N_3281,N_3110,N_3165);
xnor U3282 (N_3282,N_3173,N_3031);
xnor U3283 (N_3283,N_3172,N_3045);
or U3284 (N_3284,N_3070,N_3162);
nor U3285 (N_3285,N_3038,N_3191);
xor U3286 (N_3286,N_3071,N_3084);
nand U3287 (N_3287,N_3039,N_3109);
xnor U3288 (N_3288,N_3062,N_3018);
and U3289 (N_3289,N_3108,N_3163);
nand U3290 (N_3290,N_3166,N_3017);
nand U3291 (N_3291,N_3076,N_3143);
nand U3292 (N_3292,N_3135,N_3116);
xor U3293 (N_3293,N_3192,N_3157);
or U3294 (N_3294,N_3056,N_3188);
and U3295 (N_3295,N_3002,N_3006);
nand U3296 (N_3296,N_3154,N_3187);
xnor U3297 (N_3297,N_3105,N_3104);
and U3298 (N_3298,N_3057,N_3158);
nor U3299 (N_3299,N_3013,N_3130);
or U3300 (N_3300,N_3047,N_3166);
xor U3301 (N_3301,N_3144,N_3116);
and U3302 (N_3302,N_3154,N_3161);
or U3303 (N_3303,N_3145,N_3196);
or U3304 (N_3304,N_3108,N_3121);
or U3305 (N_3305,N_3179,N_3001);
or U3306 (N_3306,N_3052,N_3059);
or U3307 (N_3307,N_3031,N_3007);
xor U3308 (N_3308,N_3140,N_3193);
nand U3309 (N_3309,N_3168,N_3135);
or U3310 (N_3310,N_3041,N_3104);
nor U3311 (N_3311,N_3058,N_3147);
and U3312 (N_3312,N_3198,N_3105);
and U3313 (N_3313,N_3088,N_3072);
nand U3314 (N_3314,N_3108,N_3025);
xnor U3315 (N_3315,N_3174,N_3001);
and U3316 (N_3316,N_3024,N_3139);
nor U3317 (N_3317,N_3167,N_3147);
nand U3318 (N_3318,N_3180,N_3130);
nor U3319 (N_3319,N_3133,N_3128);
nor U3320 (N_3320,N_3102,N_3152);
nor U3321 (N_3321,N_3114,N_3065);
and U3322 (N_3322,N_3106,N_3022);
nand U3323 (N_3323,N_3079,N_3124);
nand U3324 (N_3324,N_3021,N_3167);
or U3325 (N_3325,N_3163,N_3066);
xnor U3326 (N_3326,N_3060,N_3105);
and U3327 (N_3327,N_3040,N_3042);
xnor U3328 (N_3328,N_3042,N_3028);
nand U3329 (N_3329,N_3109,N_3086);
or U3330 (N_3330,N_3018,N_3013);
or U3331 (N_3331,N_3033,N_3031);
or U3332 (N_3332,N_3053,N_3072);
xor U3333 (N_3333,N_3025,N_3068);
xor U3334 (N_3334,N_3112,N_3024);
and U3335 (N_3335,N_3149,N_3010);
and U3336 (N_3336,N_3076,N_3084);
nand U3337 (N_3337,N_3077,N_3134);
xor U3338 (N_3338,N_3004,N_3111);
nor U3339 (N_3339,N_3143,N_3079);
and U3340 (N_3340,N_3158,N_3088);
xor U3341 (N_3341,N_3113,N_3127);
and U3342 (N_3342,N_3145,N_3156);
xor U3343 (N_3343,N_3187,N_3144);
and U3344 (N_3344,N_3195,N_3188);
or U3345 (N_3345,N_3065,N_3067);
nand U3346 (N_3346,N_3191,N_3052);
xor U3347 (N_3347,N_3054,N_3140);
and U3348 (N_3348,N_3141,N_3059);
xor U3349 (N_3349,N_3102,N_3072);
or U3350 (N_3350,N_3068,N_3143);
or U3351 (N_3351,N_3110,N_3014);
nand U3352 (N_3352,N_3175,N_3040);
and U3353 (N_3353,N_3060,N_3147);
or U3354 (N_3354,N_3029,N_3183);
xor U3355 (N_3355,N_3150,N_3094);
or U3356 (N_3356,N_3103,N_3016);
or U3357 (N_3357,N_3018,N_3067);
xor U3358 (N_3358,N_3070,N_3080);
nor U3359 (N_3359,N_3102,N_3129);
or U3360 (N_3360,N_3184,N_3087);
nand U3361 (N_3361,N_3110,N_3108);
xnor U3362 (N_3362,N_3047,N_3172);
or U3363 (N_3363,N_3116,N_3183);
nor U3364 (N_3364,N_3100,N_3142);
nor U3365 (N_3365,N_3139,N_3122);
and U3366 (N_3366,N_3156,N_3194);
and U3367 (N_3367,N_3161,N_3115);
nand U3368 (N_3368,N_3122,N_3141);
xnor U3369 (N_3369,N_3129,N_3016);
or U3370 (N_3370,N_3102,N_3134);
and U3371 (N_3371,N_3151,N_3083);
nand U3372 (N_3372,N_3041,N_3191);
nand U3373 (N_3373,N_3164,N_3109);
nor U3374 (N_3374,N_3092,N_3095);
nand U3375 (N_3375,N_3078,N_3185);
and U3376 (N_3376,N_3029,N_3098);
nor U3377 (N_3377,N_3092,N_3169);
nand U3378 (N_3378,N_3097,N_3157);
nand U3379 (N_3379,N_3079,N_3092);
nor U3380 (N_3380,N_3020,N_3152);
xor U3381 (N_3381,N_3060,N_3182);
nor U3382 (N_3382,N_3076,N_3010);
and U3383 (N_3383,N_3085,N_3181);
nand U3384 (N_3384,N_3134,N_3053);
nor U3385 (N_3385,N_3108,N_3148);
nor U3386 (N_3386,N_3183,N_3147);
or U3387 (N_3387,N_3197,N_3075);
xnor U3388 (N_3388,N_3059,N_3130);
or U3389 (N_3389,N_3054,N_3182);
or U3390 (N_3390,N_3112,N_3114);
or U3391 (N_3391,N_3098,N_3038);
or U3392 (N_3392,N_3195,N_3158);
nor U3393 (N_3393,N_3156,N_3189);
nand U3394 (N_3394,N_3125,N_3142);
xor U3395 (N_3395,N_3079,N_3051);
or U3396 (N_3396,N_3114,N_3109);
nand U3397 (N_3397,N_3076,N_3081);
nand U3398 (N_3398,N_3166,N_3100);
nand U3399 (N_3399,N_3068,N_3199);
or U3400 (N_3400,N_3335,N_3267);
and U3401 (N_3401,N_3206,N_3346);
nand U3402 (N_3402,N_3311,N_3255);
xnor U3403 (N_3403,N_3247,N_3373);
or U3404 (N_3404,N_3351,N_3269);
nand U3405 (N_3405,N_3222,N_3388);
or U3406 (N_3406,N_3333,N_3298);
or U3407 (N_3407,N_3262,N_3245);
or U3408 (N_3408,N_3358,N_3397);
xor U3409 (N_3409,N_3341,N_3290);
nand U3410 (N_3410,N_3279,N_3238);
nand U3411 (N_3411,N_3256,N_3359);
or U3412 (N_3412,N_3220,N_3379);
or U3413 (N_3413,N_3211,N_3216);
nor U3414 (N_3414,N_3319,N_3234);
xor U3415 (N_3415,N_3337,N_3203);
nand U3416 (N_3416,N_3309,N_3350);
nand U3417 (N_3417,N_3249,N_3324);
nand U3418 (N_3418,N_3280,N_3328);
and U3419 (N_3419,N_3225,N_3297);
xor U3420 (N_3420,N_3229,N_3292);
and U3421 (N_3421,N_3381,N_3382);
nor U3422 (N_3422,N_3268,N_3361);
xor U3423 (N_3423,N_3342,N_3261);
nor U3424 (N_3424,N_3248,N_3364);
nand U3425 (N_3425,N_3375,N_3369);
and U3426 (N_3426,N_3398,N_3305);
nand U3427 (N_3427,N_3274,N_3212);
nor U3428 (N_3428,N_3224,N_3242);
nor U3429 (N_3429,N_3231,N_3352);
or U3430 (N_3430,N_3362,N_3227);
nor U3431 (N_3431,N_3370,N_3380);
xnor U3432 (N_3432,N_3217,N_3260);
nor U3433 (N_3433,N_3284,N_3276);
or U3434 (N_3434,N_3377,N_3330);
nand U3435 (N_3435,N_3254,N_3295);
and U3436 (N_3436,N_3208,N_3259);
nand U3437 (N_3437,N_3326,N_3201);
nand U3438 (N_3438,N_3243,N_3293);
or U3439 (N_3439,N_3288,N_3313);
and U3440 (N_3440,N_3396,N_3307);
and U3441 (N_3441,N_3393,N_3365);
nor U3442 (N_3442,N_3289,N_3334);
or U3443 (N_3443,N_3285,N_3232);
and U3444 (N_3444,N_3310,N_3300);
nor U3445 (N_3445,N_3219,N_3320);
nand U3446 (N_3446,N_3383,N_3270);
or U3447 (N_3447,N_3278,N_3221);
nor U3448 (N_3448,N_3282,N_3391);
or U3449 (N_3449,N_3389,N_3258);
or U3450 (N_3450,N_3317,N_3318);
and U3451 (N_3451,N_3360,N_3392);
nand U3452 (N_3452,N_3348,N_3271);
nand U3453 (N_3453,N_3343,N_3336);
nand U3454 (N_3454,N_3240,N_3325);
or U3455 (N_3455,N_3299,N_3399);
nor U3456 (N_3456,N_3390,N_3226);
or U3457 (N_3457,N_3252,N_3344);
and U3458 (N_3458,N_3304,N_3287);
or U3459 (N_3459,N_3296,N_3327);
or U3460 (N_3460,N_3306,N_3347);
nand U3461 (N_3461,N_3257,N_3209);
or U3462 (N_3462,N_3236,N_3387);
nand U3463 (N_3463,N_3230,N_3338);
and U3464 (N_3464,N_3356,N_3349);
nand U3465 (N_3465,N_3291,N_3384);
and U3466 (N_3466,N_3214,N_3367);
or U3467 (N_3467,N_3237,N_3283);
and U3468 (N_3468,N_3277,N_3395);
xor U3469 (N_3469,N_3385,N_3345);
nand U3470 (N_3470,N_3264,N_3376);
nor U3471 (N_3471,N_3202,N_3331);
nand U3472 (N_3472,N_3272,N_3235);
xor U3473 (N_3473,N_3215,N_3339);
and U3474 (N_3474,N_3213,N_3250);
or U3475 (N_3475,N_3303,N_3354);
or U3476 (N_3476,N_3378,N_3312);
nor U3477 (N_3477,N_3241,N_3265);
nand U3478 (N_3478,N_3314,N_3322);
and U3479 (N_3479,N_3205,N_3368);
and U3480 (N_3480,N_3273,N_3372);
and U3481 (N_3481,N_3357,N_3218);
nor U3482 (N_3482,N_3315,N_3210);
or U3483 (N_3483,N_3316,N_3394);
and U3484 (N_3484,N_3332,N_3275);
xor U3485 (N_3485,N_3266,N_3207);
or U3486 (N_3486,N_3233,N_3244);
nand U3487 (N_3487,N_3386,N_3200);
or U3488 (N_3488,N_3374,N_3355);
and U3489 (N_3489,N_3366,N_3340);
nand U3490 (N_3490,N_3251,N_3239);
nand U3491 (N_3491,N_3294,N_3281);
nand U3492 (N_3492,N_3353,N_3253);
xor U3493 (N_3493,N_3321,N_3286);
or U3494 (N_3494,N_3204,N_3371);
xor U3495 (N_3495,N_3246,N_3223);
or U3496 (N_3496,N_3329,N_3323);
nand U3497 (N_3497,N_3308,N_3302);
or U3498 (N_3498,N_3363,N_3228);
nor U3499 (N_3499,N_3301,N_3263);
nand U3500 (N_3500,N_3372,N_3367);
or U3501 (N_3501,N_3221,N_3259);
xor U3502 (N_3502,N_3385,N_3339);
xnor U3503 (N_3503,N_3309,N_3360);
nor U3504 (N_3504,N_3211,N_3321);
xnor U3505 (N_3505,N_3396,N_3302);
nand U3506 (N_3506,N_3362,N_3264);
and U3507 (N_3507,N_3373,N_3378);
nor U3508 (N_3508,N_3269,N_3369);
and U3509 (N_3509,N_3254,N_3322);
nand U3510 (N_3510,N_3356,N_3301);
and U3511 (N_3511,N_3238,N_3356);
and U3512 (N_3512,N_3239,N_3244);
xor U3513 (N_3513,N_3296,N_3324);
and U3514 (N_3514,N_3370,N_3275);
nand U3515 (N_3515,N_3337,N_3397);
nand U3516 (N_3516,N_3285,N_3226);
xor U3517 (N_3517,N_3306,N_3323);
or U3518 (N_3518,N_3395,N_3219);
xor U3519 (N_3519,N_3302,N_3274);
nor U3520 (N_3520,N_3398,N_3378);
nand U3521 (N_3521,N_3357,N_3257);
or U3522 (N_3522,N_3368,N_3234);
xnor U3523 (N_3523,N_3390,N_3256);
nand U3524 (N_3524,N_3364,N_3300);
nand U3525 (N_3525,N_3221,N_3372);
nor U3526 (N_3526,N_3241,N_3349);
nor U3527 (N_3527,N_3377,N_3370);
and U3528 (N_3528,N_3351,N_3307);
and U3529 (N_3529,N_3351,N_3335);
xor U3530 (N_3530,N_3203,N_3310);
and U3531 (N_3531,N_3219,N_3313);
nand U3532 (N_3532,N_3357,N_3228);
xor U3533 (N_3533,N_3274,N_3252);
or U3534 (N_3534,N_3231,N_3291);
xor U3535 (N_3535,N_3202,N_3325);
nand U3536 (N_3536,N_3397,N_3294);
xor U3537 (N_3537,N_3241,N_3225);
xnor U3538 (N_3538,N_3345,N_3354);
and U3539 (N_3539,N_3373,N_3323);
nor U3540 (N_3540,N_3205,N_3310);
xnor U3541 (N_3541,N_3226,N_3361);
nand U3542 (N_3542,N_3306,N_3248);
and U3543 (N_3543,N_3269,N_3290);
and U3544 (N_3544,N_3371,N_3346);
nand U3545 (N_3545,N_3375,N_3305);
or U3546 (N_3546,N_3326,N_3332);
nand U3547 (N_3547,N_3208,N_3316);
nand U3548 (N_3548,N_3390,N_3388);
and U3549 (N_3549,N_3200,N_3354);
or U3550 (N_3550,N_3254,N_3351);
and U3551 (N_3551,N_3273,N_3281);
and U3552 (N_3552,N_3243,N_3338);
or U3553 (N_3553,N_3393,N_3262);
nand U3554 (N_3554,N_3309,N_3392);
or U3555 (N_3555,N_3263,N_3280);
and U3556 (N_3556,N_3305,N_3372);
and U3557 (N_3557,N_3221,N_3338);
xor U3558 (N_3558,N_3390,N_3237);
nor U3559 (N_3559,N_3242,N_3262);
and U3560 (N_3560,N_3321,N_3274);
or U3561 (N_3561,N_3346,N_3327);
xnor U3562 (N_3562,N_3360,N_3244);
and U3563 (N_3563,N_3378,N_3389);
or U3564 (N_3564,N_3213,N_3358);
or U3565 (N_3565,N_3379,N_3393);
or U3566 (N_3566,N_3354,N_3277);
and U3567 (N_3567,N_3398,N_3220);
and U3568 (N_3568,N_3301,N_3248);
nor U3569 (N_3569,N_3282,N_3352);
nand U3570 (N_3570,N_3210,N_3336);
and U3571 (N_3571,N_3261,N_3357);
and U3572 (N_3572,N_3319,N_3250);
and U3573 (N_3573,N_3254,N_3266);
and U3574 (N_3574,N_3257,N_3388);
or U3575 (N_3575,N_3235,N_3281);
nor U3576 (N_3576,N_3226,N_3268);
and U3577 (N_3577,N_3236,N_3301);
nand U3578 (N_3578,N_3358,N_3243);
nor U3579 (N_3579,N_3336,N_3250);
nand U3580 (N_3580,N_3370,N_3358);
xor U3581 (N_3581,N_3335,N_3324);
xor U3582 (N_3582,N_3321,N_3351);
and U3583 (N_3583,N_3306,N_3387);
nor U3584 (N_3584,N_3260,N_3222);
or U3585 (N_3585,N_3384,N_3239);
and U3586 (N_3586,N_3264,N_3299);
nor U3587 (N_3587,N_3203,N_3204);
or U3588 (N_3588,N_3233,N_3210);
nor U3589 (N_3589,N_3290,N_3249);
xor U3590 (N_3590,N_3369,N_3286);
and U3591 (N_3591,N_3281,N_3329);
nor U3592 (N_3592,N_3389,N_3228);
nand U3593 (N_3593,N_3269,N_3324);
nor U3594 (N_3594,N_3276,N_3378);
and U3595 (N_3595,N_3344,N_3353);
xnor U3596 (N_3596,N_3226,N_3385);
and U3597 (N_3597,N_3384,N_3315);
and U3598 (N_3598,N_3262,N_3363);
nand U3599 (N_3599,N_3331,N_3258);
xnor U3600 (N_3600,N_3458,N_3471);
xnor U3601 (N_3601,N_3537,N_3414);
nand U3602 (N_3602,N_3542,N_3520);
nor U3603 (N_3603,N_3490,N_3565);
nor U3604 (N_3604,N_3541,N_3512);
and U3605 (N_3605,N_3494,N_3474);
and U3606 (N_3606,N_3462,N_3488);
and U3607 (N_3607,N_3440,N_3487);
or U3608 (N_3608,N_3500,N_3405);
xnor U3609 (N_3609,N_3485,N_3588);
xnor U3610 (N_3610,N_3453,N_3548);
nor U3611 (N_3611,N_3577,N_3468);
or U3612 (N_3612,N_3590,N_3563);
nand U3613 (N_3613,N_3492,N_3409);
xnor U3614 (N_3614,N_3460,N_3429);
nand U3615 (N_3615,N_3401,N_3427);
nor U3616 (N_3616,N_3554,N_3599);
xnor U3617 (N_3617,N_3421,N_3523);
and U3618 (N_3618,N_3435,N_3406);
and U3619 (N_3619,N_3549,N_3477);
xor U3620 (N_3620,N_3529,N_3594);
and U3621 (N_3621,N_3498,N_3502);
nor U3622 (N_3622,N_3459,N_3596);
and U3623 (N_3623,N_3457,N_3410);
or U3624 (N_3624,N_3572,N_3568);
nor U3625 (N_3625,N_3546,N_3522);
xnor U3626 (N_3626,N_3438,N_3569);
and U3627 (N_3627,N_3455,N_3432);
nor U3628 (N_3628,N_3595,N_3499);
and U3629 (N_3629,N_3493,N_3430);
or U3630 (N_3630,N_3422,N_3579);
and U3631 (N_3631,N_3570,N_3456);
xnor U3632 (N_3632,N_3504,N_3558);
nor U3633 (N_3633,N_3425,N_3575);
and U3634 (N_3634,N_3479,N_3519);
or U3635 (N_3635,N_3553,N_3413);
xnor U3636 (N_3636,N_3449,N_3545);
or U3637 (N_3637,N_3517,N_3495);
and U3638 (N_3638,N_3564,N_3528);
and U3639 (N_3639,N_3431,N_3551);
or U3640 (N_3640,N_3521,N_3497);
and U3641 (N_3641,N_3589,N_3445);
nand U3642 (N_3642,N_3581,N_3547);
nand U3643 (N_3643,N_3481,N_3583);
nand U3644 (N_3644,N_3446,N_3559);
and U3645 (N_3645,N_3505,N_3424);
or U3646 (N_3646,N_3411,N_3403);
nor U3647 (N_3647,N_3514,N_3451);
xor U3648 (N_3648,N_3530,N_3496);
or U3649 (N_3649,N_3472,N_3557);
nor U3650 (N_3650,N_3400,N_3540);
nor U3651 (N_3651,N_3544,N_3543);
or U3652 (N_3652,N_3452,N_3586);
nand U3653 (N_3653,N_3417,N_3437);
or U3654 (N_3654,N_3503,N_3527);
xnor U3655 (N_3655,N_3473,N_3464);
xor U3656 (N_3656,N_3584,N_3415);
xnor U3657 (N_3657,N_3566,N_3571);
and U3658 (N_3658,N_3592,N_3513);
or U3659 (N_3659,N_3478,N_3442);
nand U3660 (N_3660,N_3454,N_3484);
and U3661 (N_3661,N_3573,N_3536);
nor U3662 (N_3662,N_3448,N_3436);
and U3663 (N_3663,N_3418,N_3524);
nor U3664 (N_3664,N_3469,N_3574);
or U3665 (N_3665,N_3526,N_3516);
xor U3666 (N_3666,N_3518,N_3561);
nand U3667 (N_3667,N_3423,N_3463);
or U3668 (N_3668,N_3531,N_3585);
nand U3669 (N_3669,N_3408,N_3426);
xor U3670 (N_3670,N_3447,N_3465);
or U3671 (N_3671,N_3501,N_3412);
or U3672 (N_3672,N_3482,N_3587);
and U3673 (N_3673,N_3476,N_3552);
nor U3674 (N_3674,N_3538,N_3535);
nand U3675 (N_3675,N_3489,N_3402);
nand U3676 (N_3676,N_3508,N_3576);
nor U3677 (N_3677,N_3555,N_3539);
or U3678 (N_3678,N_3506,N_3560);
nor U3679 (N_3679,N_3598,N_3593);
nand U3680 (N_3680,N_3443,N_3515);
nand U3681 (N_3681,N_3509,N_3556);
nor U3682 (N_3682,N_3461,N_3470);
nand U3683 (N_3683,N_3533,N_3407);
and U3684 (N_3684,N_3511,N_3420);
xnor U3685 (N_3685,N_3404,N_3507);
nor U3686 (N_3686,N_3419,N_3466);
and U3687 (N_3687,N_3591,N_3525);
nand U3688 (N_3688,N_3550,N_3428);
xor U3689 (N_3689,N_3534,N_3567);
or U3690 (N_3690,N_3510,N_3450);
nand U3691 (N_3691,N_3416,N_3562);
or U3692 (N_3692,N_3480,N_3467);
nand U3693 (N_3693,N_3491,N_3582);
or U3694 (N_3694,N_3483,N_3444);
xnor U3695 (N_3695,N_3578,N_3475);
nand U3696 (N_3696,N_3532,N_3433);
nor U3697 (N_3697,N_3441,N_3486);
xnor U3698 (N_3698,N_3439,N_3434);
nor U3699 (N_3699,N_3580,N_3597);
and U3700 (N_3700,N_3413,N_3483);
xor U3701 (N_3701,N_3408,N_3556);
or U3702 (N_3702,N_3440,N_3578);
xor U3703 (N_3703,N_3488,N_3510);
and U3704 (N_3704,N_3550,N_3481);
nand U3705 (N_3705,N_3555,N_3502);
and U3706 (N_3706,N_3478,N_3485);
nand U3707 (N_3707,N_3421,N_3453);
and U3708 (N_3708,N_3492,N_3534);
xnor U3709 (N_3709,N_3449,N_3452);
xnor U3710 (N_3710,N_3504,N_3464);
nor U3711 (N_3711,N_3525,N_3519);
nand U3712 (N_3712,N_3436,N_3431);
and U3713 (N_3713,N_3578,N_3552);
nor U3714 (N_3714,N_3506,N_3536);
xor U3715 (N_3715,N_3585,N_3489);
and U3716 (N_3716,N_3576,N_3582);
nand U3717 (N_3717,N_3500,N_3474);
or U3718 (N_3718,N_3437,N_3595);
nor U3719 (N_3719,N_3491,N_3561);
nor U3720 (N_3720,N_3452,N_3562);
or U3721 (N_3721,N_3551,N_3506);
nor U3722 (N_3722,N_3415,N_3520);
or U3723 (N_3723,N_3570,N_3436);
nand U3724 (N_3724,N_3443,N_3590);
and U3725 (N_3725,N_3478,N_3534);
nor U3726 (N_3726,N_3442,N_3409);
xnor U3727 (N_3727,N_3490,N_3497);
and U3728 (N_3728,N_3561,N_3454);
nor U3729 (N_3729,N_3502,N_3595);
nor U3730 (N_3730,N_3575,N_3522);
xor U3731 (N_3731,N_3483,N_3469);
nand U3732 (N_3732,N_3494,N_3506);
nor U3733 (N_3733,N_3445,N_3577);
xor U3734 (N_3734,N_3476,N_3490);
nor U3735 (N_3735,N_3574,N_3584);
nor U3736 (N_3736,N_3539,N_3404);
xor U3737 (N_3737,N_3470,N_3434);
or U3738 (N_3738,N_3475,N_3497);
and U3739 (N_3739,N_3561,N_3504);
xnor U3740 (N_3740,N_3531,N_3435);
nor U3741 (N_3741,N_3532,N_3430);
and U3742 (N_3742,N_3444,N_3409);
and U3743 (N_3743,N_3425,N_3529);
nand U3744 (N_3744,N_3406,N_3517);
and U3745 (N_3745,N_3529,N_3454);
and U3746 (N_3746,N_3446,N_3412);
xnor U3747 (N_3747,N_3474,N_3580);
nor U3748 (N_3748,N_3434,N_3563);
nor U3749 (N_3749,N_3446,N_3439);
or U3750 (N_3750,N_3491,N_3573);
or U3751 (N_3751,N_3424,N_3499);
xor U3752 (N_3752,N_3479,N_3545);
or U3753 (N_3753,N_3457,N_3597);
nand U3754 (N_3754,N_3529,N_3429);
nand U3755 (N_3755,N_3409,N_3407);
xnor U3756 (N_3756,N_3573,N_3578);
xnor U3757 (N_3757,N_3553,N_3422);
or U3758 (N_3758,N_3556,N_3447);
nor U3759 (N_3759,N_3496,N_3429);
or U3760 (N_3760,N_3433,N_3491);
nor U3761 (N_3761,N_3469,N_3464);
and U3762 (N_3762,N_3447,N_3494);
and U3763 (N_3763,N_3512,N_3569);
nand U3764 (N_3764,N_3497,N_3482);
and U3765 (N_3765,N_3458,N_3548);
and U3766 (N_3766,N_3495,N_3591);
nand U3767 (N_3767,N_3435,N_3570);
nand U3768 (N_3768,N_3413,N_3590);
or U3769 (N_3769,N_3485,N_3567);
and U3770 (N_3770,N_3461,N_3592);
and U3771 (N_3771,N_3449,N_3567);
nand U3772 (N_3772,N_3507,N_3577);
nand U3773 (N_3773,N_3549,N_3453);
nand U3774 (N_3774,N_3544,N_3467);
nand U3775 (N_3775,N_3436,N_3492);
nor U3776 (N_3776,N_3548,N_3499);
and U3777 (N_3777,N_3528,N_3485);
or U3778 (N_3778,N_3404,N_3403);
and U3779 (N_3779,N_3582,N_3483);
xor U3780 (N_3780,N_3503,N_3417);
xor U3781 (N_3781,N_3428,N_3519);
or U3782 (N_3782,N_3445,N_3567);
xnor U3783 (N_3783,N_3425,N_3475);
or U3784 (N_3784,N_3593,N_3515);
and U3785 (N_3785,N_3551,N_3461);
nor U3786 (N_3786,N_3537,N_3559);
or U3787 (N_3787,N_3423,N_3471);
xnor U3788 (N_3788,N_3553,N_3557);
and U3789 (N_3789,N_3405,N_3465);
and U3790 (N_3790,N_3581,N_3582);
or U3791 (N_3791,N_3489,N_3512);
xor U3792 (N_3792,N_3478,N_3465);
nand U3793 (N_3793,N_3550,N_3557);
nor U3794 (N_3794,N_3501,N_3558);
xnor U3795 (N_3795,N_3527,N_3485);
xnor U3796 (N_3796,N_3456,N_3443);
nor U3797 (N_3797,N_3461,N_3595);
and U3798 (N_3798,N_3446,N_3576);
and U3799 (N_3799,N_3412,N_3513);
nor U3800 (N_3800,N_3662,N_3765);
or U3801 (N_3801,N_3664,N_3611);
nand U3802 (N_3802,N_3630,N_3787);
nor U3803 (N_3803,N_3767,N_3704);
and U3804 (N_3804,N_3797,N_3741);
nand U3805 (N_3805,N_3724,N_3676);
nor U3806 (N_3806,N_3792,N_3673);
and U3807 (N_3807,N_3694,N_3693);
xnor U3808 (N_3808,N_3682,N_3723);
and U3809 (N_3809,N_3698,N_3614);
or U3810 (N_3810,N_3701,N_3622);
or U3811 (N_3811,N_3768,N_3715);
and U3812 (N_3812,N_3669,N_3601);
or U3813 (N_3813,N_3660,N_3631);
nor U3814 (N_3814,N_3779,N_3729);
nand U3815 (N_3815,N_3613,N_3790);
xor U3816 (N_3816,N_3685,N_3720);
xor U3817 (N_3817,N_3702,N_3726);
nand U3818 (N_3818,N_3670,N_3760);
nor U3819 (N_3819,N_3788,N_3713);
or U3820 (N_3820,N_3684,N_3647);
and U3821 (N_3821,N_3616,N_3759);
and U3822 (N_3822,N_3652,N_3712);
xor U3823 (N_3823,N_3785,N_3755);
and U3824 (N_3824,N_3776,N_3757);
nor U3825 (N_3825,N_3608,N_3615);
xor U3826 (N_3826,N_3653,N_3744);
xnor U3827 (N_3827,N_3783,N_3777);
nor U3828 (N_3828,N_3665,N_3738);
xor U3829 (N_3829,N_3707,N_3706);
nor U3830 (N_3830,N_3648,N_3633);
or U3831 (N_3831,N_3716,N_3742);
and U3832 (N_3832,N_3600,N_3617);
nand U3833 (N_3833,N_3714,N_3740);
xnor U3834 (N_3834,N_3644,N_3634);
or U3835 (N_3835,N_3639,N_3773);
nor U3836 (N_3836,N_3780,N_3678);
xnor U3837 (N_3837,N_3679,N_3717);
or U3838 (N_3838,N_3672,N_3656);
nand U3839 (N_3839,N_3705,N_3733);
nor U3840 (N_3840,N_3753,N_3642);
nand U3841 (N_3841,N_3756,N_3754);
nand U3842 (N_3842,N_3654,N_3624);
nand U3843 (N_3843,N_3671,N_3677);
and U3844 (N_3844,N_3771,N_3609);
nand U3845 (N_3845,N_3650,N_3782);
nor U3846 (N_3846,N_3764,N_3668);
nand U3847 (N_3847,N_3623,N_3766);
and U3848 (N_3848,N_3703,N_3657);
nand U3849 (N_3849,N_3745,N_3789);
nor U3850 (N_3850,N_3725,N_3603);
or U3851 (N_3851,N_3637,N_3735);
nand U3852 (N_3852,N_3667,N_3618);
xor U3853 (N_3853,N_3646,N_3620);
xnor U3854 (N_3854,N_3688,N_3711);
nor U3855 (N_3855,N_3697,N_3649);
nor U3856 (N_3856,N_3791,N_3629);
and U3857 (N_3857,N_3749,N_3619);
nand U3858 (N_3858,N_3718,N_3674);
or U3859 (N_3859,N_3612,N_3610);
nor U3860 (N_3860,N_3778,N_3748);
or U3861 (N_3861,N_3643,N_3736);
or U3862 (N_3862,N_3728,N_3763);
nand U3863 (N_3863,N_3722,N_3770);
nand U3864 (N_3864,N_3627,N_3795);
nand U3865 (N_3865,N_3746,N_3604);
nor U3866 (N_3866,N_3680,N_3645);
nand U3867 (N_3867,N_3659,N_3625);
and U3868 (N_3868,N_3750,N_3699);
or U3869 (N_3869,N_3663,N_3621);
or U3870 (N_3870,N_3793,N_3727);
nand U3871 (N_3871,N_3607,N_3761);
nand U3872 (N_3872,N_3758,N_3762);
or U3873 (N_3873,N_3686,N_3794);
nor U3874 (N_3874,N_3632,N_3798);
nand U3875 (N_3875,N_3730,N_3721);
and U3876 (N_3876,N_3638,N_3695);
nor U3877 (N_3877,N_3690,N_3655);
nand U3878 (N_3878,N_3658,N_3799);
and U3879 (N_3879,N_3692,N_3786);
xor U3880 (N_3880,N_3635,N_3719);
and U3881 (N_3881,N_3606,N_3769);
xor U3882 (N_3882,N_3666,N_3640);
or U3883 (N_3883,N_3734,N_3774);
and U3884 (N_3884,N_3775,N_3641);
xor U3885 (N_3885,N_3709,N_3696);
nor U3886 (N_3886,N_3732,N_3626);
nor U3887 (N_3887,N_3784,N_3751);
nor U3888 (N_3888,N_3772,N_3710);
nand U3889 (N_3889,N_3636,N_3747);
nor U3890 (N_3890,N_3661,N_3781);
or U3891 (N_3891,N_3737,N_3651);
or U3892 (N_3892,N_3700,N_3691);
nand U3893 (N_3893,N_3675,N_3628);
and U3894 (N_3894,N_3681,N_3743);
nand U3895 (N_3895,N_3683,N_3731);
nor U3896 (N_3896,N_3708,N_3752);
nor U3897 (N_3897,N_3689,N_3605);
and U3898 (N_3898,N_3687,N_3739);
nand U3899 (N_3899,N_3796,N_3602);
xor U3900 (N_3900,N_3654,N_3730);
nand U3901 (N_3901,N_3760,N_3645);
and U3902 (N_3902,N_3768,N_3642);
xor U3903 (N_3903,N_3646,N_3734);
or U3904 (N_3904,N_3785,N_3688);
xor U3905 (N_3905,N_3767,N_3605);
nand U3906 (N_3906,N_3741,N_3652);
xnor U3907 (N_3907,N_3682,N_3745);
nand U3908 (N_3908,N_3675,N_3715);
xor U3909 (N_3909,N_3703,N_3789);
and U3910 (N_3910,N_3763,N_3778);
nor U3911 (N_3911,N_3622,N_3736);
xor U3912 (N_3912,N_3732,N_3756);
and U3913 (N_3913,N_3720,N_3735);
or U3914 (N_3914,N_3642,N_3712);
xor U3915 (N_3915,N_3770,N_3698);
xnor U3916 (N_3916,N_3628,N_3619);
nor U3917 (N_3917,N_3611,N_3660);
nand U3918 (N_3918,N_3620,N_3633);
or U3919 (N_3919,N_3694,N_3653);
nand U3920 (N_3920,N_3787,N_3782);
and U3921 (N_3921,N_3667,N_3616);
and U3922 (N_3922,N_3785,N_3660);
nand U3923 (N_3923,N_3721,N_3690);
and U3924 (N_3924,N_3634,N_3698);
and U3925 (N_3925,N_3780,N_3766);
and U3926 (N_3926,N_3713,N_3641);
nor U3927 (N_3927,N_3741,N_3710);
or U3928 (N_3928,N_3766,N_3608);
and U3929 (N_3929,N_3795,N_3702);
and U3930 (N_3930,N_3713,N_3733);
or U3931 (N_3931,N_3760,N_3762);
nor U3932 (N_3932,N_3612,N_3673);
nor U3933 (N_3933,N_3738,N_3678);
nor U3934 (N_3934,N_3728,N_3616);
and U3935 (N_3935,N_3635,N_3744);
or U3936 (N_3936,N_3747,N_3683);
xor U3937 (N_3937,N_3747,N_3797);
xor U3938 (N_3938,N_3744,N_3738);
or U3939 (N_3939,N_3679,N_3703);
and U3940 (N_3940,N_3736,N_3723);
nor U3941 (N_3941,N_3623,N_3661);
xor U3942 (N_3942,N_3684,N_3715);
xnor U3943 (N_3943,N_3610,N_3754);
nand U3944 (N_3944,N_3738,N_3633);
and U3945 (N_3945,N_3607,N_3685);
and U3946 (N_3946,N_3683,N_3703);
nand U3947 (N_3947,N_3613,N_3791);
nand U3948 (N_3948,N_3741,N_3762);
and U3949 (N_3949,N_3743,N_3749);
and U3950 (N_3950,N_3629,N_3706);
nor U3951 (N_3951,N_3758,N_3626);
or U3952 (N_3952,N_3736,N_3658);
nand U3953 (N_3953,N_3703,N_3614);
or U3954 (N_3954,N_3622,N_3716);
xor U3955 (N_3955,N_3624,N_3726);
xor U3956 (N_3956,N_3786,N_3784);
xor U3957 (N_3957,N_3749,N_3797);
xor U3958 (N_3958,N_3703,N_3782);
xnor U3959 (N_3959,N_3675,N_3648);
nand U3960 (N_3960,N_3604,N_3699);
xnor U3961 (N_3961,N_3693,N_3797);
nor U3962 (N_3962,N_3644,N_3756);
nand U3963 (N_3963,N_3656,N_3605);
or U3964 (N_3964,N_3765,N_3671);
xor U3965 (N_3965,N_3741,N_3753);
xor U3966 (N_3966,N_3707,N_3641);
and U3967 (N_3967,N_3767,N_3783);
or U3968 (N_3968,N_3790,N_3797);
nand U3969 (N_3969,N_3726,N_3711);
nand U3970 (N_3970,N_3797,N_3799);
xnor U3971 (N_3971,N_3615,N_3613);
nor U3972 (N_3972,N_3637,N_3685);
and U3973 (N_3973,N_3607,N_3705);
or U3974 (N_3974,N_3661,N_3644);
and U3975 (N_3975,N_3722,N_3619);
and U3976 (N_3976,N_3623,N_3761);
nor U3977 (N_3977,N_3622,N_3733);
and U3978 (N_3978,N_3773,N_3781);
nand U3979 (N_3979,N_3687,N_3776);
nand U3980 (N_3980,N_3794,N_3753);
or U3981 (N_3981,N_3673,N_3635);
or U3982 (N_3982,N_3634,N_3649);
or U3983 (N_3983,N_3699,N_3757);
nor U3984 (N_3984,N_3799,N_3721);
or U3985 (N_3985,N_3789,N_3767);
nand U3986 (N_3986,N_3776,N_3611);
and U3987 (N_3987,N_3609,N_3765);
nand U3988 (N_3988,N_3677,N_3689);
or U3989 (N_3989,N_3654,N_3749);
and U3990 (N_3990,N_3713,N_3741);
or U3991 (N_3991,N_3638,N_3622);
xor U3992 (N_3992,N_3712,N_3783);
and U3993 (N_3993,N_3673,N_3659);
and U3994 (N_3994,N_3705,N_3672);
nor U3995 (N_3995,N_3764,N_3609);
nor U3996 (N_3996,N_3701,N_3729);
and U3997 (N_3997,N_3678,N_3795);
and U3998 (N_3998,N_3760,N_3612);
nor U3999 (N_3999,N_3781,N_3637);
nand U4000 (N_4000,N_3966,N_3889);
nand U4001 (N_4001,N_3880,N_3943);
nand U4002 (N_4002,N_3802,N_3863);
nand U4003 (N_4003,N_3940,N_3814);
nor U4004 (N_4004,N_3952,N_3977);
xor U4005 (N_4005,N_3998,N_3894);
xnor U4006 (N_4006,N_3861,N_3807);
or U4007 (N_4007,N_3905,N_3804);
nor U4008 (N_4008,N_3835,N_3926);
and U4009 (N_4009,N_3860,N_3806);
nand U4010 (N_4010,N_3873,N_3929);
or U4011 (N_4011,N_3920,N_3946);
nand U4012 (N_4012,N_3812,N_3906);
and U4013 (N_4013,N_3840,N_3949);
nor U4014 (N_4014,N_3980,N_3999);
xor U4015 (N_4015,N_3988,N_3992);
and U4016 (N_4016,N_3884,N_3984);
nand U4017 (N_4017,N_3847,N_3936);
nor U4018 (N_4018,N_3848,N_3883);
xnor U4019 (N_4019,N_3886,N_3978);
and U4020 (N_4020,N_3831,N_3991);
xnor U4021 (N_4021,N_3826,N_3827);
and U4022 (N_4022,N_3972,N_3959);
xor U4023 (N_4023,N_3960,N_3918);
and U4024 (N_4024,N_3934,N_3979);
nor U4025 (N_4025,N_3830,N_3904);
xor U4026 (N_4026,N_3842,N_3938);
and U4027 (N_4027,N_3907,N_3866);
xnor U4028 (N_4028,N_3834,N_3951);
nand U4029 (N_4029,N_3963,N_3933);
and U4030 (N_4030,N_3879,N_3947);
and U4031 (N_4031,N_3898,N_3981);
or U4032 (N_4032,N_3955,N_3822);
and U4033 (N_4033,N_3912,N_3810);
nor U4034 (N_4034,N_3893,N_3817);
or U4035 (N_4035,N_3876,N_3865);
or U4036 (N_4036,N_3924,N_3870);
xnor U4037 (N_4037,N_3950,N_3954);
and U4038 (N_4038,N_3890,N_3844);
nor U4039 (N_4039,N_3996,N_3922);
or U4040 (N_4040,N_3909,N_3815);
xor U4041 (N_4041,N_3864,N_3994);
and U4042 (N_4042,N_3986,N_3975);
and U4043 (N_4043,N_3900,N_3921);
or U4044 (N_4044,N_3902,N_3816);
nand U4045 (N_4045,N_3857,N_3813);
xor U4046 (N_4046,N_3843,N_3897);
or U4047 (N_4047,N_3976,N_3925);
and U4048 (N_4048,N_3995,N_3881);
or U4049 (N_4049,N_3962,N_3961);
nor U4050 (N_4050,N_3927,N_3916);
nand U4051 (N_4051,N_3837,N_3930);
and U4052 (N_4052,N_3803,N_3868);
nand U4053 (N_4053,N_3821,N_3948);
and U4054 (N_4054,N_3973,N_3850);
and U4055 (N_4055,N_3832,N_3913);
nor U4056 (N_4056,N_3958,N_3856);
nor U4057 (N_4057,N_3862,N_3932);
and U4058 (N_4058,N_3941,N_3945);
or U4059 (N_4059,N_3872,N_3852);
or U4060 (N_4060,N_3935,N_3923);
and U4061 (N_4061,N_3841,N_3855);
xor U4062 (N_4062,N_3937,N_3811);
nor U4063 (N_4063,N_3944,N_3805);
xor U4064 (N_4064,N_3895,N_3915);
or U4065 (N_4065,N_3888,N_3956);
nor U4066 (N_4066,N_3983,N_3899);
xnor U4067 (N_4067,N_3896,N_3989);
xor U4068 (N_4068,N_3820,N_3970);
nor U4069 (N_4069,N_3942,N_3953);
nand U4070 (N_4070,N_3971,N_3969);
and U4071 (N_4071,N_3823,N_3982);
and U4072 (N_4072,N_3964,N_3800);
or U4073 (N_4073,N_3851,N_3987);
nor U4074 (N_4074,N_3859,N_3839);
nor U4075 (N_4075,N_3974,N_3845);
xor U4076 (N_4076,N_3997,N_3993);
and U4077 (N_4077,N_3846,N_3928);
nor U4078 (N_4078,N_3828,N_3869);
xor U4079 (N_4079,N_3874,N_3858);
nor U4080 (N_4080,N_3849,N_3824);
xnor U4081 (N_4081,N_3808,N_3809);
nor U4082 (N_4082,N_3908,N_3911);
and U4083 (N_4083,N_3965,N_3917);
and U4084 (N_4084,N_3967,N_3878);
or U4085 (N_4085,N_3957,N_3903);
xnor U4086 (N_4086,N_3833,N_3985);
or U4087 (N_4087,N_3871,N_3853);
or U4088 (N_4088,N_3854,N_3829);
xnor U4089 (N_4089,N_3885,N_3818);
xnor U4090 (N_4090,N_3877,N_3801);
nand U4091 (N_4091,N_3914,N_3990);
and U4092 (N_4092,N_3892,N_3919);
nor U4093 (N_4093,N_3891,N_3819);
and U4094 (N_4094,N_3875,N_3910);
nor U4095 (N_4095,N_3838,N_3836);
nor U4096 (N_4096,N_3825,N_3939);
or U4097 (N_4097,N_3882,N_3901);
nand U4098 (N_4098,N_3968,N_3887);
xor U4099 (N_4099,N_3867,N_3931);
nor U4100 (N_4100,N_3882,N_3978);
nand U4101 (N_4101,N_3907,N_3975);
and U4102 (N_4102,N_3992,N_3813);
nand U4103 (N_4103,N_3860,N_3906);
nor U4104 (N_4104,N_3877,N_3986);
nand U4105 (N_4105,N_3852,N_3922);
and U4106 (N_4106,N_3924,N_3988);
xnor U4107 (N_4107,N_3891,N_3867);
and U4108 (N_4108,N_3831,N_3892);
nand U4109 (N_4109,N_3910,N_3905);
nand U4110 (N_4110,N_3913,N_3997);
nor U4111 (N_4111,N_3874,N_3893);
and U4112 (N_4112,N_3976,N_3935);
xnor U4113 (N_4113,N_3824,N_3997);
xor U4114 (N_4114,N_3935,N_3815);
and U4115 (N_4115,N_3912,N_3827);
and U4116 (N_4116,N_3895,N_3802);
nand U4117 (N_4117,N_3906,N_3851);
nor U4118 (N_4118,N_3941,N_3900);
xor U4119 (N_4119,N_3806,N_3941);
nand U4120 (N_4120,N_3949,N_3847);
xnor U4121 (N_4121,N_3891,N_3991);
nand U4122 (N_4122,N_3837,N_3905);
and U4123 (N_4123,N_3843,N_3876);
nand U4124 (N_4124,N_3895,N_3862);
nand U4125 (N_4125,N_3993,N_3851);
nand U4126 (N_4126,N_3814,N_3949);
nor U4127 (N_4127,N_3911,N_3950);
and U4128 (N_4128,N_3863,N_3822);
nor U4129 (N_4129,N_3814,N_3876);
nor U4130 (N_4130,N_3823,N_3951);
and U4131 (N_4131,N_3963,N_3961);
nand U4132 (N_4132,N_3804,N_3960);
or U4133 (N_4133,N_3809,N_3816);
and U4134 (N_4134,N_3922,N_3898);
nand U4135 (N_4135,N_3853,N_3900);
xor U4136 (N_4136,N_3806,N_3988);
and U4137 (N_4137,N_3919,N_3984);
xnor U4138 (N_4138,N_3971,N_3886);
or U4139 (N_4139,N_3924,N_3807);
nor U4140 (N_4140,N_3988,N_3913);
nor U4141 (N_4141,N_3899,N_3877);
xor U4142 (N_4142,N_3927,N_3969);
or U4143 (N_4143,N_3909,N_3883);
nand U4144 (N_4144,N_3891,N_3933);
nor U4145 (N_4145,N_3958,N_3852);
xor U4146 (N_4146,N_3929,N_3974);
and U4147 (N_4147,N_3872,N_3998);
nand U4148 (N_4148,N_3800,N_3812);
nor U4149 (N_4149,N_3865,N_3835);
and U4150 (N_4150,N_3992,N_3867);
nand U4151 (N_4151,N_3942,N_3828);
nor U4152 (N_4152,N_3842,N_3881);
nand U4153 (N_4153,N_3982,N_3904);
nand U4154 (N_4154,N_3816,N_3874);
or U4155 (N_4155,N_3891,N_3818);
nand U4156 (N_4156,N_3894,N_3990);
nand U4157 (N_4157,N_3985,N_3836);
nand U4158 (N_4158,N_3807,N_3850);
nand U4159 (N_4159,N_3878,N_3838);
nor U4160 (N_4160,N_3877,N_3902);
or U4161 (N_4161,N_3843,N_3983);
xnor U4162 (N_4162,N_3811,N_3867);
nand U4163 (N_4163,N_3958,N_3948);
or U4164 (N_4164,N_3961,N_3812);
and U4165 (N_4165,N_3975,N_3946);
or U4166 (N_4166,N_3912,N_3856);
xor U4167 (N_4167,N_3886,N_3938);
and U4168 (N_4168,N_3997,N_3860);
and U4169 (N_4169,N_3843,N_3996);
nand U4170 (N_4170,N_3818,N_3850);
nand U4171 (N_4171,N_3924,N_3932);
or U4172 (N_4172,N_3837,N_3916);
or U4173 (N_4173,N_3982,N_3818);
nand U4174 (N_4174,N_3817,N_3883);
nand U4175 (N_4175,N_3888,N_3963);
xnor U4176 (N_4176,N_3927,N_3899);
xor U4177 (N_4177,N_3843,N_3884);
and U4178 (N_4178,N_3844,N_3943);
nand U4179 (N_4179,N_3984,N_3848);
nand U4180 (N_4180,N_3804,N_3903);
or U4181 (N_4181,N_3819,N_3934);
nor U4182 (N_4182,N_3946,N_3999);
and U4183 (N_4183,N_3821,N_3958);
or U4184 (N_4184,N_3953,N_3897);
nor U4185 (N_4185,N_3976,N_3828);
or U4186 (N_4186,N_3939,N_3966);
or U4187 (N_4187,N_3936,N_3816);
or U4188 (N_4188,N_3838,N_3955);
or U4189 (N_4189,N_3917,N_3992);
or U4190 (N_4190,N_3866,N_3945);
xor U4191 (N_4191,N_3803,N_3990);
nand U4192 (N_4192,N_3964,N_3882);
and U4193 (N_4193,N_3885,N_3957);
nor U4194 (N_4194,N_3912,N_3942);
or U4195 (N_4195,N_3998,N_3965);
nor U4196 (N_4196,N_3949,N_3816);
or U4197 (N_4197,N_3849,N_3877);
and U4198 (N_4198,N_3971,N_3827);
or U4199 (N_4199,N_3961,N_3871);
nor U4200 (N_4200,N_4136,N_4013);
and U4201 (N_4201,N_4021,N_4102);
xnor U4202 (N_4202,N_4054,N_4169);
or U4203 (N_4203,N_4189,N_4104);
and U4204 (N_4204,N_4178,N_4108);
nor U4205 (N_4205,N_4044,N_4122);
nor U4206 (N_4206,N_4014,N_4167);
and U4207 (N_4207,N_4026,N_4056);
and U4208 (N_4208,N_4139,N_4164);
nand U4209 (N_4209,N_4138,N_4153);
and U4210 (N_4210,N_4035,N_4128);
and U4211 (N_4211,N_4076,N_4019);
xor U4212 (N_4212,N_4006,N_4043);
xnor U4213 (N_4213,N_4093,N_4143);
and U4214 (N_4214,N_4158,N_4074);
nand U4215 (N_4215,N_4116,N_4110);
or U4216 (N_4216,N_4194,N_4015);
and U4217 (N_4217,N_4050,N_4011);
xor U4218 (N_4218,N_4047,N_4068);
or U4219 (N_4219,N_4003,N_4127);
or U4220 (N_4220,N_4062,N_4132);
nand U4221 (N_4221,N_4072,N_4126);
and U4222 (N_4222,N_4082,N_4195);
nor U4223 (N_4223,N_4109,N_4106);
nor U4224 (N_4224,N_4005,N_4030);
xnor U4225 (N_4225,N_4075,N_4087);
xor U4226 (N_4226,N_4103,N_4029);
and U4227 (N_4227,N_4060,N_4041);
and U4228 (N_4228,N_4010,N_4089);
or U4229 (N_4229,N_4079,N_4114);
nand U4230 (N_4230,N_4168,N_4183);
nand U4231 (N_4231,N_4152,N_4192);
and U4232 (N_4232,N_4187,N_4184);
nor U4233 (N_4233,N_4023,N_4179);
and U4234 (N_4234,N_4193,N_4070);
and U4235 (N_4235,N_4053,N_4022);
and U4236 (N_4236,N_4000,N_4049);
and U4237 (N_4237,N_4171,N_4159);
or U4238 (N_4238,N_4197,N_4190);
xnor U4239 (N_4239,N_4131,N_4095);
nor U4240 (N_4240,N_4088,N_4124);
xnor U4241 (N_4241,N_4042,N_4092);
or U4242 (N_4242,N_4162,N_4154);
and U4243 (N_4243,N_4174,N_4170);
or U4244 (N_4244,N_4129,N_4039);
nand U4245 (N_4245,N_4028,N_4155);
nand U4246 (N_4246,N_4017,N_4172);
or U4247 (N_4247,N_4134,N_4161);
nand U4248 (N_4248,N_4094,N_4181);
or U4249 (N_4249,N_4165,N_4099);
xnor U4250 (N_4250,N_4101,N_4166);
and U4251 (N_4251,N_4051,N_4133);
nand U4252 (N_4252,N_4185,N_4113);
and U4253 (N_4253,N_4065,N_4182);
or U4254 (N_4254,N_4078,N_4037);
and U4255 (N_4255,N_4057,N_4148);
and U4256 (N_4256,N_4020,N_4173);
and U4257 (N_4257,N_4111,N_4100);
nor U4258 (N_4258,N_4118,N_4191);
nor U4259 (N_4259,N_4081,N_4024);
and U4260 (N_4260,N_4177,N_4142);
nand U4261 (N_4261,N_4098,N_4069);
nor U4262 (N_4262,N_4115,N_4071);
xnor U4263 (N_4263,N_4033,N_4137);
and U4264 (N_4264,N_4058,N_4150);
xnor U4265 (N_4265,N_4196,N_4135);
xor U4266 (N_4266,N_4107,N_4151);
and U4267 (N_4267,N_4186,N_4198);
or U4268 (N_4268,N_4121,N_4097);
nand U4269 (N_4269,N_4160,N_4105);
and U4270 (N_4270,N_4077,N_4018);
nor U4271 (N_4271,N_4016,N_4149);
nand U4272 (N_4272,N_4085,N_4038);
nand U4273 (N_4273,N_4001,N_4141);
and U4274 (N_4274,N_4004,N_4008);
xnor U4275 (N_4275,N_4055,N_4145);
nor U4276 (N_4276,N_4032,N_4123);
nand U4277 (N_4277,N_4009,N_4091);
or U4278 (N_4278,N_4048,N_4176);
and U4279 (N_4279,N_4188,N_4090);
nand U4280 (N_4280,N_4163,N_4059);
and U4281 (N_4281,N_4064,N_4061);
nor U4282 (N_4282,N_4086,N_4036);
xor U4283 (N_4283,N_4119,N_4147);
xor U4284 (N_4284,N_4063,N_4125);
nand U4285 (N_4285,N_4096,N_4040);
or U4286 (N_4286,N_4144,N_4027);
nor U4287 (N_4287,N_4199,N_4156);
nand U4288 (N_4288,N_4080,N_4083);
and U4289 (N_4289,N_4117,N_4046);
nor U4290 (N_4290,N_4066,N_4130);
xor U4291 (N_4291,N_4140,N_4045);
and U4292 (N_4292,N_4052,N_4120);
nor U4293 (N_4293,N_4175,N_4034);
and U4294 (N_4294,N_4146,N_4007);
or U4295 (N_4295,N_4025,N_4002);
xnor U4296 (N_4296,N_4073,N_4112);
or U4297 (N_4297,N_4067,N_4031);
nand U4298 (N_4298,N_4084,N_4157);
xor U4299 (N_4299,N_4180,N_4012);
or U4300 (N_4300,N_4002,N_4015);
or U4301 (N_4301,N_4062,N_4025);
xor U4302 (N_4302,N_4112,N_4163);
xor U4303 (N_4303,N_4170,N_4094);
xor U4304 (N_4304,N_4193,N_4039);
nor U4305 (N_4305,N_4023,N_4177);
nor U4306 (N_4306,N_4001,N_4037);
xnor U4307 (N_4307,N_4116,N_4115);
nor U4308 (N_4308,N_4146,N_4014);
and U4309 (N_4309,N_4084,N_4096);
and U4310 (N_4310,N_4056,N_4160);
and U4311 (N_4311,N_4112,N_4127);
and U4312 (N_4312,N_4185,N_4176);
and U4313 (N_4313,N_4023,N_4136);
nand U4314 (N_4314,N_4010,N_4134);
nand U4315 (N_4315,N_4154,N_4065);
nor U4316 (N_4316,N_4138,N_4021);
nand U4317 (N_4317,N_4108,N_4161);
xnor U4318 (N_4318,N_4020,N_4144);
xnor U4319 (N_4319,N_4173,N_4180);
and U4320 (N_4320,N_4123,N_4122);
or U4321 (N_4321,N_4091,N_4135);
nor U4322 (N_4322,N_4087,N_4136);
nand U4323 (N_4323,N_4028,N_4137);
or U4324 (N_4324,N_4009,N_4179);
xor U4325 (N_4325,N_4063,N_4003);
and U4326 (N_4326,N_4065,N_4131);
xnor U4327 (N_4327,N_4100,N_4134);
nand U4328 (N_4328,N_4145,N_4093);
nor U4329 (N_4329,N_4130,N_4060);
nor U4330 (N_4330,N_4050,N_4139);
or U4331 (N_4331,N_4195,N_4068);
or U4332 (N_4332,N_4151,N_4002);
or U4333 (N_4333,N_4025,N_4032);
and U4334 (N_4334,N_4027,N_4035);
and U4335 (N_4335,N_4037,N_4194);
nand U4336 (N_4336,N_4128,N_4069);
nand U4337 (N_4337,N_4084,N_4068);
xnor U4338 (N_4338,N_4161,N_4064);
and U4339 (N_4339,N_4170,N_4077);
nand U4340 (N_4340,N_4167,N_4096);
and U4341 (N_4341,N_4190,N_4150);
or U4342 (N_4342,N_4038,N_4077);
nand U4343 (N_4343,N_4172,N_4192);
nand U4344 (N_4344,N_4132,N_4050);
nand U4345 (N_4345,N_4136,N_4191);
nor U4346 (N_4346,N_4184,N_4046);
or U4347 (N_4347,N_4093,N_4005);
xor U4348 (N_4348,N_4156,N_4180);
nor U4349 (N_4349,N_4132,N_4104);
or U4350 (N_4350,N_4186,N_4138);
xnor U4351 (N_4351,N_4166,N_4122);
nand U4352 (N_4352,N_4072,N_4136);
nor U4353 (N_4353,N_4007,N_4050);
nand U4354 (N_4354,N_4096,N_4120);
nor U4355 (N_4355,N_4050,N_4117);
or U4356 (N_4356,N_4157,N_4058);
nand U4357 (N_4357,N_4076,N_4045);
nand U4358 (N_4358,N_4043,N_4060);
nor U4359 (N_4359,N_4114,N_4127);
or U4360 (N_4360,N_4166,N_4181);
xor U4361 (N_4361,N_4176,N_4097);
nand U4362 (N_4362,N_4005,N_4078);
and U4363 (N_4363,N_4128,N_4153);
nor U4364 (N_4364,N_4054,N_4034);
nor U4365 (N_4365,N_4184,N_4063);
nor U4366 (N_4366,N_4063,N_4109);
nor U4367 (N_4367,N_4085,N_4111);
or U4368 (N_4368,N_4125,N_4097);
or U4369 (N_4369,N_4109,N_4075);
nand U4370 (N_4370,N_4155,N_4005);
or U4371 (N_4371,N_4146,N_4135);
nand U4372 (N_4372,N_4023,N_4133);
and U4373 (N_4373,N_4113,N_4107);
xor U4374 (N_4374,N_4027,N_4152);
or U4375 (N_4375,N_4137,N_4013);
nor U4376 (N_4376,N_4050,N_4027);
xnor U4377 (N_4377,N_4040,N_4012);
xnor U4378 (N_4378,N_4182,N_4185);
and U4379 (N_4379,N_4101,N_4094);
xnor U4380 (N_4380,N_4126,N_4140);
and U4381 (N_4381,N_4187,N_4102);
xnor U4382 (N_4382,N_4062,N_4035);
xor U4383 (N_4383,N_4191,N_4093);
or U4384 (N_4384,N_4066,N_4152);
and U4385 (N_4385,N_4165,N_4004);
nand U4386 (N_4386,N_4157,N_4021);
and U4387 (N_4387,N_4182,N_4054);
xnor U4388 (N_4388,N_4094,N_4077);
and U4389 (N_4389,N_4179,N_4068);
xor U4390 (N_4390,N_4139,N_4109);
and U4391 (N_4391,N_4147,N_4055);
or U4392 (N_4392,N_4175,N_4053);
nor U4393 (N_4393,N_4059,N_4041);
and U4394 (N_4394,N_4174,N_4150);
nor U4395 (N_4395,N_4152,N_4039);
or U4396 (N_4396,N_4032,N_4072);
nand U4397 (N_4397,N_4177,N_4172);
nand U4398 (N_4398,N_4163,N_4057);
xnor U4399 (N_4399,N_4078,N_4061);
and U4400 (N_4400,N_4283,N_4294);
xor U4401 (N_4401,N_4312,N_4353);
or U4402 (N_4402,N_4293,N_4340);
and U4403 (N_4403,N_4284,N_4245);
xor U4404 (N_4404,N_4205,N_4246);
nand U4405 (N_4405,N_4260,N_4285);
and U4406 (N_4406,N_4309,N_4269);
xnor U4407 (N_4407,N_4352,N_4335);
nand U4408 (N_4408,N_4262,N_4204);
nor U4409 (N_4409,N_4351,N_4314);
xnor U4410 (N_4410,N_4381,N_4265);
nand U4411 (N_4411,N_4344,N_4304);
nand U4412 (N_4412,N_4348,N_4208);
or U4413 (N_4413,N_4327,N_4364);
nor U4414 (N_4414,N_4261,N_4256);
nor U4415 (N_4415,N_4386,N_4207);
nand U4416 (N_4416,N_4393,N_4227);
xor U4417 (N_4417,N_4282,N_4221);
and U4418 (N_4418,N_4300,N_4303);
nand U4419 (N_4419,N_4358,N_4375);
nand U4420 (N_4420,N_4266,N_4232);
nand U4421 (N_4421,N_4373,N_4210);
xnor U4422 (N_4422,N_4224,N_4218);
nor U4423 (N_4423,N_4248,N_4363);
nor U4424 (N_4424,N_4330,N_4306);
and U4425 (N_4425,N_4298,N_4359);
xnor U4426 (N_4426,N_4339,N_4270);
nand U4427 (N_4427,N_4328,N_4349);
nor U4428 (N_4428,N_4380,N_4296);
and U4429 (N_4429,N_4288,N_4225);
nand U4430 (N_4430,N_4233,N_4377);
xor U4431 (N_4431,N_4313,N_4223);
xor U4432 (N_4432,N_4236,N_4372);
xor U4433 (N_4433,N_4329,N_4322);
nand U4434 (N_4434,N_4290,N_4215);
and U4435 (N_4435,N_4315,N_4280);
nand U4436 (N_4436,N_4244,N_4201);
xnor U4437 (N_4437,N_4354,N_4310);
or U4438 (N_4438,N_4365,N_4355);
or U4439 (N_4439,N_4239,N_4399);
nand U4440 (N_4440,N_4247,N_4252);
or U4441 (N_4441,N_4332,N_4389);
nor U4442 (N_4442,N_4211,N_4241);
or U4443 (N_4443,N_4240,N_4231);
nand U4444 (N_4444,N_4326,N_4324);
or U4445 (N_4445,N_4385,N_4297);
or U4446 (N_4446,N_4267,N_4273);
nor U4447 (N_4447,N_4311,N_4209);
or U4448 (N_4448,N_4230,N_4371);
xor U4449 (N_4449,N_4376,N_4243);
nand U4450 (N_4450,N_4219,N_4368);
nand U4451 (N_4451,N_4200,N_4337);
or U4452 (N_4452,N_4396,N_4361);
xnor U4453 (N_4453,N_4235,N_4369);
xor U4454 (N_4454,N_4391,N_4206);
nor U4455 (N_4455,N_4301,N_4387);
nand U4456 (N_4456,N_4341,N_4347);
xor U4457 (N_4457,N_4259,N_4217);
nor U4458 (N_4458,N_4258,N_4366);
nand U4459 (N_4459,N_4382,N_4251);
or U4460 (N_4460,N_4242,N_4220);
or U4461 (N_4461,N_4390,N_4238);
and U4462 (N_4462,N_4287,N_4374);
and U4463 (N_4463,N_4342,N_4289);
or U4464 (N_4464,N_4378,N_4305);
or U4465 (N_4465,N_4323,N_4222);
xor U4466 (N_4466,N_4255,N_4302);
nor U4467 (N_4467,N_4383,N_4321);
nor U4468 (N_4468,N_4271,N_4253);
xnor U4469 (N_4469,N_4367,N_4292);
or U4470 (N_4470,N_4319,N_4331);
nand U4471 (N_4471,N_4316,N_4237);
or U4472 (N_4472,N_4343,N_4263);
nor U4473 (N_4473,N_4398,N_4397);
xor U4474 (N_4474,N_4379,N_4249);
or U4475 (N_4475,N_4346,N_4272);
nor U4476 (N_4476,N_4338,N_4362);
nand U4477 (N_4477,N_4394,N_4216);
xor U4478 (N_4478,N_4357,N_4336);
xnor U4479 (N_4479,N_4279,N_4291);
or U4480 (N_4480,N_4234,N_4345);
xor U4481 (N_4481,N_4214,N_4299);
or U4482 (N_4482,N_4392,N_4274);
or U4483 (N_4483,N_4356,N_4333);
xnor U4484 (N_4484,N_4384,N_4307);
and U4485 (N_4485,N_4325,N_4295);
nor U4486 (N_4486,N_4212,N_4228);
nand U4487 (N_4487,N_4334,N_4388);
or U4488 (N_4488,N_4278,N_4360);
xor U4489 (N_4489,N_4370,N_4250);
xnor U4490 (N_4490,N_4202,N_4276);
nor U4491 (N_4491,N_4264,N_4317);
and U4492 (N_4492,N_4268,N_4254);
and U4493 (N_4493,N_4229,N_4350);
and U4494 (N_4494,N_4318,N_4226);
nor U4495 (N_4495,N_4275,N_4257);
and U4496 (N_4496,N_4286,N_4213);
and U4497 (N_4497,N_4308,N_4203);
and U4498 (N_4498,N_4320,N_4395);
nand U4499 (N_4499,N_4277,N_4281);
or U4500 (N_4500,N_4324,N_4348);
or U4501 (N_4501,N_4306,N_4360);
or U4502 (N_4502,N_4282,N_4330);
nand U4503 (N_4503,N_4262,N_4319);
xnor U4504 (N_4504,N_4301,N_4307);
or U4505 (N_4505,N_4246,N_4316);
nand U4506 (N_4506,N_4398,N_4260);
and U4507 (N_4507,N_4375,N_4203);
xnor U4508 (N_4508,N_4278,N_4235);
xor U4509 (N_4509,N_4342,N_4247);
nor U4510 (N_4510,N_4252,N_4225);
nand U4511 (N_4511,N_4393,N_4256);
or U4512 (N_4512,N_4246,N_4250);
nand U4513 (N_4513,N_4226,N_4235);
xnor U4514 (N_4514,N_4352,N_4366);
nor U4515 (N_4515,N_4289,N_4355);
nor U4516 (N_4516,N_4217,N_4288);
nand U4517 (N_4517,N_4357,N_4227);
and U4518 (N_4518,N_4332,N_4229);
or U4519 (N_4519,N_4364,N_4236);
nor U4520 (N_4520,N_4268,N_4322);
xnor U4521 (N_4521,N_4399,N_4394);
or U4522 (N_4522,N_4228,N_4256);
nand U4523 (N_4523,N_4397,N_4371);
and U4524 (N_4524,N_4339,N_4328);
or U4525 (N_4525,N_4309,N_4262);
or U4526 (N_4526,N_4375,N_4237);
or U4527 (N_4527,N_4238,N_4314);
and U4528 (N_4528,N_4368,N_4258);
nand U4529 (N_4529,N_4332,N_4209);
or U4530 (N_4530,N_4292,N_4362);
nand U4531 (N_4531,N_4373,N_4285);
or U4532 (N_4532,N_4351,N_4340);
and U4533 (N_4533,N_4350,N_4238);
nor U4534 (N_4534,N_4311,N_4293);
or U4535 (N_4535,N_4356,N_4311);
and U4536 (N_4536,N_4343,N_4237);
and U4537 (N_4537,N_4397,N_4300);
and U4538 (N_4538,N_4257,N_4315);
nand U4539 (N_4539,N_4360,N_4227);
or U4540 (N_4540,N_4316,N_4313);
nor U4541 (N_4541,N_4225,N_4220);
xor U4542 (N_4542,N_4388,N_4321);
nand U4543 (N_4543,N_4348,N_4259);
or U4544 (N_4544,N_4343,N_4392);
or U4545 (N_4545,N_4338,N_4269);
and U4546 (N_4546,N_4377,N_4365);
nor U4547 (N_4547,N_4376,N_4297);
or U4548 (N_4548,N_4248,N_4366);
and U4549 (N_4549,N_4312,N_4229);
or U4550 (N_4550,N_4305,N_4284);
or U4551 (N_4551,N_4211,N_4393);
nor U4552 (N_4552,N_4209,N_4335);
nand U4553 (N_4553,N_4267,N_4316);
nor U4554 (N_4554,N_4289,N_4374);
or U4555 (N_4555,N_4318,N_4263);
and U4556 (N_4556,N_4219,N_4397);
or U4557 (N_4557,N_4317,N_4283);
nor U4558 (N_4558,N_4254,N_4207);
xor U4559 (N_4559,N_4275,N_4298);
nand U4560 (N_4560,N_4300,N_4323);
nor U4561 (N_4561,N_4229,N_4355);
xor U4562 (N_4562,N_4236,N_4381);
xnor U4563 (N_4563,N_4272,N_4278);
xor U4564 (N_4564,N_4340,N_4316);
xor U4565 (N_4565,N_4286,N_4258);
nand U4566 (N_4566,N_4382,N_4202);
or U4567 (N_4567,N_4380,N_4204);
xnor U4568 (N_4568,N_4229,N_4248);
or U4569 (N_4569,N_4226,N_4338);
xor U4570 (N_4570,N_4358,N_4345);
and U4571 (N_4571,N_4202,N_4224);
nor U4572 (N_4572,N_4348,N_4366);
xor U4573 (N_4573,N_4244,N_4287);
nand U4574 (N_4574,N_4398,N_4203);
nand U4575 (N_4575,N_4237,N_4389);
xnor U4576 (N_4576,N_4288,N_4203);
nand U4577 (N_4577,N_4293,N_4270);
nor U4578 (N_4578,N_4206,N_4317);
nand U4579 (N_4579,N_4381,N_4386);
nand U4580 (N_4580,N_4219,N_4342);
and U4581 (N_4581,N_4207,N_4295);
or U4582 (N_4582,N_4211,N_4396);
xor U4583 (N_4583,N_4320,N_4263);
and U4584 (N_4584,N_4264,N_4382);
and U4585 (N_4585,N_4203,N_4293);
nor U4586 (N_4586,N_4276,N_4304);
nor U4587 (N_4587,N_4383,N_4264);
nor U4588 (N_4588,N_4288,N_4269);
or U4589 (N_4589,N_4385,N_4376);
and U4590 (N_4590,N_4226,N_4211);
xnor U4591 (N_4591,N_4318,N_4323);
or U4592 (N_4592,N_4302,N_4315);
or U4593 (N_4593,N_4273,N_4292);
xor U4594 (N_4594,N_4203,N_4286);
nand U4595 (N_4595,N_4200,N_4201);
or U4596 (N_4596,N_4291,N_4249);
nor U4597 (N_4597,N_4360,N_4224);
nor U4598 (N_4598,N_4312,N_4333);
nand U4599 (N_4599,N_4373,N_4268);
nor U4600 (N_4600,N_4591,N_4470);
nor U4601 (N_4601,N_4404,N_4459);
or U4602 (N_4602,N_4582,N_4583);
nand U4603 (N_4603,N_4532,N_4446);
or U4604 (N_4604,N_4478,N_4594);
or U4605 (N_4605,N_4505,N_4590);
or U4606 (N_4606,N_4529,N_4580);
and U4607 (N_4607,N_4595,N_4568);
nor U4608 (N_4608,N_4515,N_4474);
and U4609 (N_4609,N_4424,N_4488);
nand U4610 (N_4610,N_4442,N_4471);
nor U4611 (N_4611,N_4540,N_4422);
nand U4612 (N_4612,N_4517,N_4411);
and U4613 (N_4613,N_4425,N_4530);
and U4614 (N_4614,N_4581,N_4437);
or U4615 (N_4615,N_4562,N_4416);
nor U4616 (N_4616,N_4533,N_4509);
nand U4617 (N_4617,N_4447,N_4401);
nand U4618 (N_4618,N_4467,N_4545);
nor U4619 (N_4619,N_4445,N_4503);
nor U4620 (N_4620,N_4486,N_4405);
xnor U4621 (N_4621,N_4482,N_4454);
xor U4622 (N_4622,N_4520,N_4448);
nand U4623 (N_4623,N_4541,N_4599);
nand U4624 (N_4624,N_4436,N_4423);
and U4625 (N_4625,N_4500,N_4550);
and U4626 (N_4626,N_4563,N_4458);
and U4627 (N_4627,N_4496,N_4400);
xnor U4628 (N_4628,N_4477,N_4491);
and U4629 (N_4629,N_4483,N_4490);
xor U4630 (N_4630,N_4537,N_4434);
nor U4631 (N_4631,N_4465,N_4552);
nor U4632 (N_4632,N_4527,N_4410);
nand U4633 (N_4633,N_4456,N_4551);
nand U4634 (N_4634,N_4526,N_4484);
and U4635 (N_4635,N_4531,N_4572);
and U4636 (N_4636,N_4586,N_4507);
and U4637 (N_4637,N_4439,N_4455);
nand U4638 (N_4638,N_4579,N_4544);
nand U4639 (N_4639,N_4513,N_4564);
or U4640 (N_4640,N_4506,N_4501);
nand U4641 (N_4641,N_4460,N_4567);
nor U4642 (N_4642,N_4559,N_4539);
xor U4643 (N_4643,N_4556,N_4577);
and U4644 (N_4644,N_4548,N_4407);
nand U4645 (N_4645,N_4593,N_4438);
nand U4646 (N_4646,N_4421,N_4464);
and U4647 (N_4647,N_4596,N_4589);
and U4648 (N_4648,N_4479,N_4431);
and U4649 (N_4649,N_4440,N_4487);
xor U4650 (N_4650,N_4457,N_4419);
and U4651 (N_4651,N_4502,N_4511);
or U4652 (N_4652,N_4462,N_4555);
nor U4653 (N_4653,N_4558,N_4430);
or U4654 (N_4654,N_4578,N_4570);
nor U4655 (N_4655,N_4469,N_4554);
nor U4656 (N_4656,N_4480,N_4574);
and U4657 (N_4657,N_4566,N_4497);
xor U4658 (N_4658,N_4499,N_4519);
nor U4659 (N_4659,N_4587,N_4403);
xor U4660 (N_4660,N_4584,N_4553);
nand U4661 (N_4661,N_4476,N_4585);
and U4662 (N_4662,N_4489,N_4546);
nand U4663 (N_4663,N_4514,N_4535);
xor U4664 (N_4664,N_4523,N_4543);
or U4665 (N_4665,N_4576,N_4406);
nor U4666 (N_4666,N_4414,N_4557);
or U4667 (N_4667,N_4441,N_4598);
and U4668 (N_4668,N_4561,N_4536);
nor U4669 (N_4669,N_4463,N_4444);
nand U4670 (N_4670,N_4528,N_4592);
or U4671 (N_4671,N_4468,N_4418);
and U4672 (N_4672,N_4466,N_4426);
nand U4673 (N_4673,N_4573,N_4565);
nor U4674 (N_4674,N_4435,N_4473);
or U4675 (N_4675,N_4450,N_4415);
xor U4676 (N_4676,N_4485,N_4475);
or U4677 (N_4677,N_4472,N_4498);
nor U4678 (N_4678,N_4549,N_4510);
xnor U4679 (N_4679,N_4504,N_4518);
or U4680 (N_4680,N_4534,N_4453);
or U4681 (N_4681,N_4560,N_4508);
nor U4682 (N_4682,N_4588,N_4547);
or U4683 (N_4683,N_4516,N_4542);
xor U4684 (N_4684,N_4449,N_4495);
nor U4685 (N_4685,N_4494,N_4412);
and U4686 (N_4686,N_4417,N_4409);
nor U4687 (N_4687,N_4428,N_4432);
and U4688 (N_4688,N_4413,N_4521);
and U4689 (N_4689,N_4429,N_4492);
and U4690 (N_4690,N_4427,N_4408);
nand U4691 (N_4691,N_4538,N_4493);
or U4692 (N_4692,N_4569,N_4452);
or U4693 (N_4693,N_4597,N_4420);
nand U4694 (N_4694,N_4461,N_4522);
or U4695 (N_4695,N_4481,N_4433);
xnor U4696 (N_4696,N_4443,N_4525);
nor U4697 (N_4697,N_4524,N_4575);
xnor U4698 (N_4698,N_4512,N_4571);
nand U4699 (N_4699,N_4451,N_4402);
nor U4700 (N_4700,N_4459,N_4581);
or U4701 (N_4701,N_4472,N_4553);
or U4702 (N_4702,N_4467,N_4424);
xor U4703 (N_4703,N_4495,N_4563);
and U4704 (N_4704,N_4457,N_4524);
nor U4705 (N_4705,N_4546,N_4508);
nor U4706 (N_4706,N_4549,N_4470);
or U4707 (N_4707,N_4420,N_4522);
xnor U4708 (N_4708,N_4564,N_4524);
and U4709 (N_4709,N_4485,N_4454);
or U4710 (N_4710,N_4502,N_4406);
and U4711 (N_4711,N_4405,N_4494);
nand U4712 (N_4712,N_4536,N_4558);
or U4713 (N_4713,N_4440,N_4578);
or U4714 (N_4714,N_4499,N_4495);
nor U4715 (N_4715,N_4402,N_4459);
nor U4716 (N_4716,N_4411,N_4430);
or U4717 (N_4717,N_4428,N_4479);
and U4718 (N_4718,N_4559,N_4443);
nand U4719 (N_4719,N_4412,N_4574);
and U4720 (N_4720,N_4536,N_4404);
and U4721 (N_4721,N_4470,N_4582);
nor U4722 (N_4722,N_4523,N_4407);
and U4723 (N_4723,N_4599,N_4438);
xor U4724 (N_4724,N_4556,N_4490);
or U4725 (N_4725,N_4420,N_4598);
nor U4726 (N_4726,N_4405,N_4506);
xor U4727 (N_4727,N_4575,N_4415);
nor U4728 (N_4728,N_4574,N_4443);
xnor U4729 (N_4729,N_4565,N_4471);
nand U4730 (N_4730,N_4456,N_4444);
nand U4731 (N_4731,N_4546,N_4451);
xor U4732 (N_4732,N_4477,N_4411);
nand U4733 (N_4733,N_4573,N_4461);
and U4734 (N_4734,N_4531,N_4461);
or U4735 (N_4735,N_4469,N_4492);
nand U4736 (N_4736,N_4435,N_4555);
xnor U4737 (N_4737,N_4508,N_4520);
nand U4738 (N_4738,N_4561,N_4511);
xor U4739 (N_4739,N_4597,N_4512);
and U4740 (N_4740,N_4437,N_4504);
xor U4741 (N_4741,N_4567,N_4584);
xnor U4742 (N_4742,N_4437,N_4513);
nand U4743 (N_4743,N_4586,N_4562);
nand U4744 (N_4744,N_4551,N_4510);
nor U4745 (N_4745,N_4403,N_4482);
or U4746 (N_4746,N_4548,N_4531);
and U4747 (N_4747,N_4471,N_4425);
or U4748 (N_4748,N_4561,N_4406);
and U4749 (N_4749,N_4414,N_4576);
nor U4750 (N_4750,N_4427,N_4433);
and U4751 (N_4751,N_4593,N_4553);
nand U4752 (N_4752,N_4464,N_4598);
nor U4753 (N_4753,N_4405,N_4553);
and U4754 (N_4754,N_4438,N_4547);
and U4755 (N_4755,N_4415,N_4566);
or U4756 (N_4756,N_4407,N_4439);
nor U4757 (N_4757,N_4438,N_4597);
nand U4758 (N_4758,N_4485,N_4400);
nand U4759 (N_4759,N_4452,N_4481);
and U4760 (N_4760,N_4421,N_4561);
or U4761 (N_4761,N_4415,N_4419);
or U4762 (N_4762,N_4525,N_4502);
nand U4763 (N_4763,N_4597,N_4560);
nor U4764 (N_4764,N_4437,N_4572);
and U4765 (N_4765,N_4489,N_4427);
xnor U4766 (N_4766,N_4553,N_4541);
and U4767 (N_4767,N_4475,N_4443);
nand U4768 (N_4768,N_4520,N_4584);
nor U4769 (N_4769,N_4559,N_4536);
nor U4770 (N_4770,N_4558,N_4422);
nor U4771 (N_4771,N_4401,N_4494);
nand U4772 (N_4772,N_4580,N_4503);
xor U4773 (N_4773,N_4583,N_4460);
and U4774 (N_4774,N_4561,N_4403);
nor U4775 (N_4775,N_4525,N_4403);
or U4776 (N_4776,N_4477,N_4540);
nor U4777 (N_4777,N_4548,N_4536);
nor U4778 (N_4778,N_4541,N_4538);
or U4779 (N_4779,N_4400,N_4426);
and U4780 (N_4780,N_4408,N_4493);
or U4781 (N_4781,N_4582,N_4461);
nor U4782 (N_4782,N_4540,N_4563);
or U4783 (N_4783,N_4420,N_4511);
xnor U4784 (N_4784,N_4488,N_4475);
and U4785 (N_4785,N_4540,N_4471);
nand U4786 (N_4786,N_4583,N_4464);
or U4787 (N_4787,N_4500,N_4469);
nor U4788 (N_4788,N_4461,N_4403);
xnor U4789 (N_4789,N_4407,N_4512);
xnor U4790 (N_4790,N_4557,N_4436);
xnor U4791 (N_4791,N_4440,N_4401);
and U4792 (N_4792,N_4435,N_4416);
nor U4793 (N_4793,N_4593,N_4492);
nand U4794 (N_4794,N_4580,N_4402);
nand U4795 (N_4795,N_4560,N_4578);
or U4796 (N_4796,N_4556,N_4549);
nor U4797 (N_4797,N_4527,N_4438);
nand U4798 (N_4798,N_4477,N_4575);
and U4799 (N_4799,N_4410,N_4543);
and U4800 (N_4800,N_4733,N_4776);
nor U4801 (N_4801,N_4713,N_4684);
xor U4802 (N_4802,N_4793,N_4620);
and U4803 (N_4803,N_4685,N_4785);
xor U4804 (N_4804,N_4751,N_4702);
and U4805 (N_4805,N_4749,N_4689);
xor U4806 (N_4806,N_4732,N_4700);
xor U4807 (N_4807,N_4623,N_4681);
nor U4808 (N_4808,N_4647,N_4784);
xnor U4809 (N_4809,N_4614,N_4672);
or U4810 (N_4810,N_4731,N_4788);
nand U4811 (N_4811,N_4709,N_4797);
nor U4812 (N_4812,N_4634,N_4611);
xor U4813 (N_4813,N_4769,N_4730);
nand U4814 (N_4814,N_4682,N_4636);
and U4815 (N_4815,N_4716,N_4720);
nor U4816 (N_4816,N_4692,N_4632);
and U4817 (N_4817,N_4603,N_4798);
and U4818 (N_4818,N_4637,N_4640);
nand U4819 (N_4819,N_4646,N_4762);
xor U4820 (N_4820,N_4666,N_4626);
or U4821 (N_4821,N_4792,N_4653);
and U4822 (N_4822,N_4624,N_4693);
nor U4823 (N_4823,N_4704,N_4728);
nand U4824 (N_4824,N_4754,N_4606);
nand U4825 (N_4825,N_4764,N_4775);
and U4826 (N_4826,N_4694,N_4686);
xnor U4827 (N_4827,N_4605,N_4667);
or U4828 (N_4828,N_4711,N_4717);
or U4829 (N_4829,N_4616,N_4688);
and U4830 (N_4830,N_4691,N_4745);
xor U4831 (N_4831,N_4781,N_4744);
nand U4832 (N_4832,N_4604,N_4779);
and U4833 (N_4833,N_4673,N_4724);
nand U4834 (N_4834,N_4687,N_4789);
xor U4835 (N_4835,N_4786,N_4629);
nor U4836 (N_4836,N_4652,N_4655);
nand U4837 (N_4837,N_4639,N_4767);
xor U4838 (N_4838,N_4707,N_4755);
or U4839 (N_4839,N_4670,N_4746);
nand U4840 (N_4840,N_4770,N_4699);
or U4841 (N_4841,N_4662,N_4663);
and U4842 (N_4842,N_4703,N_4638);
nor U4843 (N_4843,N_4743,N_4738);
xnor U4844 (N_4844,N_4750,N_4665);
and U4845 (N_4845,N_4627,N_4787);
or U4846 (N_4846,N_4763,N_4772);
and U4847 (N_4847,N_4705,N_4610);
nor U4848 (N_4848,N_4613,N_4719);
and U4849 (N_4849,N_4674,N_4735);
or U4850 (N_4850,N_4773,N_4723);
xor U4851 (N_4851,N_4656,N_4630);
nand U4852 (N_4852,N_4664,N_4617);
xor U4853 (N_4853,N_4690,N_4759);
and U4854 (N_4854,N_4615,N_4718);
and U4855 (N_4855,N_4706,N_4601);
nor U4856 (N_4856,N_4635,N_4677);
nor U4857 (N_4857,N_4618,N_4651);
and U4858 (N_4858,N_4600,N_4714);
and U4859 (N_4859,N_4619,N_4696);
nor U4860 (N_4860,N_4780,N_4683);
nand U4861 (N_4861,N_4737,N_4660);
xnor U4862 (N_4862,N_4729,N_4649);
nand U4863 (N_4863,N_4625,N_4760);
nand U4864 (N_4864,N_4768,N_4771);
xnor U4865 (N_4865,N_4740,N_4607);
and U4866 (N_4866,N_4645,N_4680);
xor U4867 (N_4867,N_4722,N_4774);
and U4868 (N_4868,N_4658,N_4621);
nand U4869 (N_4869,N_4796,N_4777);
and U4870 (N_4870,N_4633,N_4650);
and U4871 (N_4871,N_4747,N_4758);
nand U4872 (N_4872,N_4783,N_4654);
nor U4873 (N_4873,N_4710,N_4695);
or U4874 (N_4874,N_4698,N_4753);
and U4875 (N_4875,N_4734,N_4679);
or U4876 (N_4876,N_4757,N_4712);
and U4877 (N_4877,N_4752,N_4657);
nand U4878 (N_4878,N_4741,N_4782);
xor U4879 (N_4879,N_4791,N_4678);
nand U4880 (N_4880,N_4622,N_4643);
nor U4881 (N_4881,N_4609,N_4676);
and U4882 (N_4882,N_4765,N_4794);
nor U4883 (N_4883,N_4612,N_4725);
nand U4884 (N_4884,N_4628,N_4790);
nor U4885 (N_4885,N_4608,N_4675);
nand U4886 (N_4886,N_4701,N_4671);
or U4887 (N_4887,N_4742,N_4659);
and U4888 (N_4888,N_4602,N_4726);
xnor U4889 (N_4889,N_4631,N_4748);
nor U4890 (N_4890,N_4727,N_4799);
nor U4891 (N_4891,N_4736,N_4715);
xor U4892 (N_4892,N_4661,N_4648);
xnor U4893 (N_4893,N_4668,N_4756);
nor U4894 (N_4894,N_4761,N_4739);
nor U4895 (N_4895,N_4669,N_4778);
nor U4896 (N_4896,N_4795,N_4641);
or U4897 (N_4897,N_4708,N_4697);
nand U4898 (N_4898,N_4644,N_4721);
nor U4899 (N_4899,N_4766,N_4642);
nor U4900 (N_4900,N_4680,N_4799);
or U4901 (N_4901,N_4614,N_4729);
nand U4902 (N_4902,N_4660,N_4739);
and U4903 (N_4903,N_4671,N_4711);
and U4904 (N_4904,N_4617,N_4736);
nand U4905 (N_4905,N_4717,N_4671);
and U4906 (N_4906,N_4647,N_4759);
nand U4907 (N_4907,N_4720,N_4690);
nand U4908 (N_4908,N_4744,N_4661);
nor U4909 (N_4909,N_4743,N_4655);
nand U4910 (N_4910,N_4786,N_4760);
nand U4911 (N_4911,N_4782,N_4674);
nor U4912 (N_4912,N_4630,N_4771);
or U4913 (N_4913,N_4650,N_4658);
or U4914 (N_4914,N_4729,N_4772);
nor U4915 (N_4915,N_4790,N_4755);
and U4916 (N_4916,N_4725,N_4702);
nand U4917 (N_4917,N_4607,N_4604);
nor U4918 (N_4918,N_4650,N_4717);
nor U4919 (N_4919,N_4733,N_4728);
nor U4920 (N_4920,N_4601,N_4786);
nand U4921 (N_4921,N_4750,N_4669);
and U4922 (N_4922,N_4748,N_4766);
nor U4923 (N_4923,N_4683,N_4629);
xor U4924 (N_4924,N_4699,N_4642);
or U4925 (N_4925,N_4744,N_4657);
xnor U4926 (N_4926,N_4704,N_4794);
or U4927 (N_4927,N_4605,N_4678);
and U4928 (N_4928,N_4602,N_4676);
nor U4929 (N_4929,N_4795,N_4624);
xnor U4930 (N_4930,N_4763,N_4677);
and U4931 (N_4931,N_4761,N_4741);
nand U4932 (N_4932,N_4620,N_4776);
and U4933 (N_4933,N_4786,N_4666);
xor U4934 (N_4934,N_4679,N_4648);
and U4935 (N_4935,N_4694,N_4653);
and U4936 (N_4936,N_4611,N_4761);
or U4937 (N_4937,N_4669,N_4606);
nor U4938 (N_4938,N_4781,N_4603);
xnor U4939 (N_4939,N_4730,N_4670);
nor U4940 (N_4940,N_4728,N_4722);
xnor U4941 (N_4941,N_4651,N_4705);
nand U4942 (N_4942,N_4790,N_4605);
xnor U4943 (N_4943,N_4756,N_4626);
or U4944 (N_4944,N_4749,N_4604);
nand U4945 (N_4945,N_4749,N_4607);
or U4946 (N_4946,N_4683,N_4675);
xnor U4947 (N_4947,N_4777,N_4676);
or U4948 (N_4948,N_4758,N_4611);
xor U4949 (N_4949,N_4730,N_4791);
nand U4950 (N_4950,N_4772,N_4730);
nand U4951 (N_4951,N_4781,N_4790);
xor U4952 (N_4952,N_4726,N_4783);
nand U4953 (N_4953,N_4727,N_4698);
xnor U4954 (N_4954,N_4620,N_4600);
and U4955 (N_4955,N_4600,N_4723);
xor U4956 (N_4956,N_4625,N_4601);
or U4957 (N_4957,N_4721,N_4624);
nand U4958 (N_4958,N_4795,N_4668);
and U4959 (N_4959,N_4730,N_4727);
nand U4960 (N_4960,N_4782,N_4622);
or U4961 (N_4961,N_4631,N_4625);
nor U4962 (N_4962,N_4601,N_4743);
nand U4963 (N_4963,N_4771,N_4795);
xnor U4964 (N_4964,N_4606,N_4694);
nand U4965 (N_4965,N_4779,N_4776);
or U4966 (N_4966,N_4641,N_4783);
nor U4967 (N_4967,N_4708,N_4790);
or U4968 (N_4968,N_4709,N_4663);
or U4969 (N_4969,N_4710,N_4704);
or U4970 (N_4970,N_4665,N_4659);
and U4971 (N_4971,N_4765,N_4775);
and U4972 (N_4972,N_4753,N_4705);
xnor U4973 (N_4973,N_4763,N_4786);
nor U4974 (N_4974,N_4767,N_4694);
and U4975 (N_4975,N_4640,N_4677);
nor U4976 (N_4976,N_4670,N_4631);
xor U4977 (N_4977,N_4626,N_4695);
or U4978 (N_4978,N_4682,N_4718);
or U4979 (N_4979,N_4727,N_4618);
and U4980 (N_4980,N_4734,N_4624);
nor U4981 (N_4981,N_4726,N_4604);
and U4982 (N_4982,N_4795,N_4689);
and U4983 (N_4983,N_4634,N_4715);
nand U4984 (N_4984,N_4641,N_4666);
nand U4985 (N_4985,N_4630,N_4658);
or U4986 (N_4986,N_4773,N_4604);
and U4987 (N_4987,N_4696,N_4685);
nor U4988 (N_4988,N_4722,N_4765);
xnor U4989 (N_4989,N_4631,N_4773);
or U4990 (N_4990,N_4623,N_4622);
nor U4991 (N_4991,N_4766,N_4781);
nor U4992 (N_4992,N_4708,N_4611);
nand U4993 (N_4993,N_4760,N_4793);
nor U4994 (N_4994,N_4644,N_4692);
nand U4995 (N_4995,N_4613,N_4630);
nor U4996 (N_4996,N_4673,N_4719);
nor U4997 (N_4997,N_4774,N_4741);
nor U4998 (N_4998,N_4617,N_4706);
and U4999 (N_4999,N_4705,N_4790);
nand U5000 (N_5000,N_4885,N_4957);
xnor U5001 (N_5001,N_4912,N_4925);
and U5002 (N_5002,N_4807,N_4984);
xnor U5003 (N_5003,N_4864,N_4820);
nand U5004 (N_5004,N_4859,N_4840);
xor U5005 (N_5005,N_4884,N_4891);
nand U5006 (N_5006,N_4968,N_4839);
and U5007 (N_5007,N_4818,N_4841);
or U5008 (N_5008,N_4961,N_4998);
nor U5009 (N_5009,N_4910,N_4836);
xor U5010 (N_5010,N_4953,N_4995);
and U5011 (N_5011,N_4861,N_4921);
xor U5012 (N_5012,N_4950,N_4846);
and U5013 (N_5013,N_4920,N_4808);
and U5014 (N_5014,N_4835,N_4972);
and U5015 (N_5015,N_4865,N_4863);
xnor U5016 (N_5016,N_4889,N_4928);
nand U5017 (N_5017,N_4978,N_4816);
nand U5018 (N_5018,N_4933,N_4958);
and U5019 (N_5019,N_4860,N_4855);
and U5020 (N_5020,N_4981,N_4952);
xnor U5021 (N_5021,N_4917,N_4869);
and U5022 (N_5022,N_4858,N_4913);
nand U5023 (N_5023,N_4943,N_4821);
xor U5024 (N_5024,N_4969,N_4923);
nand U5025 (N_5025,N_4862,N_4980);
or U5026 (N_5026,N_4976,N_4898);
and U5027 (N_5027,N_4954,N_4990);
xor U5028 (N_5028,N_4886,N_4809);
and U5029 (N_5029,N_4963,N_4938);
or U5030 (N_5030,N_4982,N_4825);
or U5031 (N_5031,N_4926,N_4986);
xor U5032 (N_5032,N_4962,N_4827);
or U5033 (N_5033,N_4879,N_4993);
xnor U5034 (N_5034,N_4823,N_4838);
nor U5035 (N_5035,N_4833,N_4922);
nor U5036 (N_5036,N_4892,N_4903);
and U5037 (N_5037,N_4966,N_4826);
and U5038 (N_5038,N_4882,N_4851);
and U5039 (N_5039,N_4974,N_4894);
nand U5040 (N_5040,N_4975,N_4899);
or U5041 (N_5041,N_4842,N_4955);
or U5042 (N_5042,N_4852,N_4812);
nand U5043 (N_5043,N_4927,N_4871);
and U5044 (N_5044,N_4802,N_4830);
nand U5045 (N_5045,N_4813,N_4960);
xnor U5046 (N_5046,N_4956,N_4902);
nor U5047 (N_5047,N_4931,N_4936);
or U5048 (N_5048,N_4867,N_4806);
and U5049 (N_5049,N_4985,N_4906);
nand U5050 (N_5050,N_4887,N_4843);
xor U5051 (N_5051,N_4991,N_4890);
xnor U5052 (N_5052,N_4992,N_4977);
and U5053 (N_5053,N_4949,N_4915);
and U5054 (N_5054,N_4944,N_4811);
xnor U5055 (N_5055,N_4937,N_4856);
nor U5056 (N_5056,N_4900,N_4848);
nor U5057 (N_5057,N_4803,N_4934);
xor U5058 (N_5058,N_4908,N_4911);
xor U5059 (N_5059,N_4929,N_4964);
or U5060 (N_5060,N_4942,N_4989);
or U5061 (N_5061,N_4904,N_4979);
nor U5062 (N_5062,N_4872,N_4951);
and U5063 (N_5063,N_4918,N_4849);
and U5064 (N_5064,N_4947,N_4994);
xnor U5065 (N_5065,N_4905,N_4845);
nand U5066 (N_5066,N_4895,N_4983);
or U5067 (N_5067,N_4907,N_4973);
nor U5068 (N_5068,N_4870,N_4854);
nand U5069 (N_5069,N_4805,N_4817);
nor U5070 (N_5070,N_4873,N_4901);
xor U5071 (N_5071,N_4834,N_4822);
nand U5072 (N_5072,N_4919,N_4819);
xnor U5073 (N_5073,N_4996,N_4829);
nand U5074 (N_5074,N_4814,N_4935);
and U5075 (N_5075,N_4815,N_4971);
nor U5076 (N_5076,N_4832,N_4850);
and U5077 (N_5077,N_4866,N_4857);
and U5078 (N_5078,N_4831,N_4941);
or U5079 (N_5079,N_4924,N_4837);
nor U5080 (N_5080,N_4868,N_4965);
nor U5081 (N_5081,N_4824,N_4930);
and U5082 (N_5082,N_4997,N_4878);
nand U5083 (N_5083,N_4970,N_4914);
nand U5084 (N_5084,N_4909,N_4946);
and U5085 (N_5085,N_4874,N_4853);
nand U5086 (N_5086,N_4987,N_4883);
nand U5087 (N_5087,N_4916,N_4844);
nand U5088 (N_5088,N_4932,N_4988);
xnor U5089 (N_5089,N_4967,N_4880);
xor U5090 (N_5090,N_4875,N_4847);
or U5091 (N_5091,N_4948,N_4876);
nor U5092 (N_5092,N_4801,N_4810);
xnor U5093 (N_5093,N_4940,N_4800);
or U5094 (N_5094,N_4877,N_4893);
and U5095 (N_5095,N_4804,N_4959);
nand U5096 (N_5096,N_4888,N_4896);
or U5097 (N_5097,N_4939,N_4897);
and U5098 (N_5098,N_4945,N_4999);
nor U5099 (N_5099,N_4828,N_4881);
nor U5100 (N_5100,N_4952,N_4905);
or U5101 (N_5101,N_4944,N_4882);
nand U5102 (N_5102,N_4871,N_4882);
xor U5103 (N_5103,N_4874,N_4999);
nand U5104 (N_5104,N_4901,N_4978);
nand U5105 (N_5105,N_4919,N_4895);
and U5106 (N_5106,N_4876,N_4819);
nand U5107 (N_5107,N_4994,N_4940);
nand U5108 (N_5108,N_4805,N_4831);
nor U5109 (N_5109,N_4914,N_4986);
or U5110 (N_5110,N_4983,N_4934);
nand U5111 (N_5111,N_4887,N_4911);
nand U5112 (N_5112,N_4913,N_4976);
and U5113 (N_5113,N_4994,N_4992);
xor U5114 (N_5114,N_4805,N_4971);
nand U5115 (N_5115,N_4998,N_4869);
nand U5116 (N_5116,N_4882,N_4931);
nand U5117 (N_5117,N_4945,N_4852);
or U5118 (N_5118,N_4942,N_4944);
xor U5119 (N_5119,N_4995,N_4917);
or U5120 (N_5120,N_4975,N_4953);
and U5121 (N_5121,N_4907,N_4931);
xor U5122 (N_5122,N_4807,N_4941);
or U5123 (N_5123,N_4887,N_4905);
xor U5124 (N_5124,N_4931,N_4895);
and U5125 (N_5125,N_4811,N_4947);
and U5126 (N_5126,N_4927,N_4821);
nor U5127 (N_5127,N_4896,N_4980);
xnor U5128 (N_5128,N_4939,N_4840);
xor U5129 (N_5129,N_4850,N_4978);
nor U5130 (N_5130,N_4846,N_4888);
nor U5131 (N_5131,N_4812,N_4826);
or U5132 (N_5132,N_4848,N_4871);
and U5133 (N_5133,N_4949,N_4828);
xor U5134 (N_5134,N_4964,N_4901);
or U5135 (N_5135,N_4890,N_4878);
or U5136 (N_5136,N_4881,N_4852);
nand U5137 (N_5137,N_4984,N_4819);
and U5138 (N_5138,N_4891,N_4882);
or U5139 (N_5139,N_4962,N_4977);
or U5140 (N_5140,N_4809,N_4861);
xor U5141 (N_5141,N_4881,N_4851);
or U5142 (N_5142,N_4871,N_4854);
and U5143 (N_5143,N_4830,N_4949);
nor U5144 (N_5144,N_4871,N_4831);
or U5145 (N_5145,N_4858,N_4904);
or U5146 (N_5146,N_4949,N_4976);
nor U5147 (N_5147,N_4865,N_4841);
or U5148 (N_5148,N_4934,N_4821);
and U5149 (N_5149,N_4877,N_4980);
or U5150 (N_5150,N_4846,N_4861);
nor U5151 (N_5151,N_4849,N_4836);
and U5152 (N_5152,N_4895,N_4894);
and U5153 (N_5153,N_4839,N_4805);
nand U5154 (N_5154,N_4989,N_4892);
xnor U5155 (N_5155,N_4967,N_4929);
or U5156 (N_5156,N_4862,N_4924);
nor U5157 (N_5157,N_4945,N_4827);
nand U5158 (N_5158,N_4834,N_4928);
nand U5159 (N_5159,N_4898,N_4859);
xnor U5160 (N_5160,N_4960,N_4864);
and U5161 (N_5161,N_4987,N_4821);
or U5162 (N_5162,N_4997,N_4979);
or U5163 (N_5163,N_4913,N_4961);
and U5164 (N_5164,N_4922,N_4835);
nand U5165 (N_5165,N_4935,N_4890);
and U5166 (N_5166,N_4825,N_4841);
or U5167 (N_5167,N_4810,N_4903);
or U5168 (N_5168,N_4835,N_4892);
or U5169 (N_5169,N_4909,N_4862);
and U5170 (N_5170,N_4843,N_4932);
and U5171 (N_5171,N_4819,N_4989);
nand U5172 (N_5172,N_4912,N_4842);
or U5173 (N_5173,N_4827,N_4805);
xnor U5174 (N_5174,N_4830,N_4968);
nand U5175 (N_5175,N_4804,N_4887);
nand U5176 (N_5176,N_4950,N_4860);
xnor U5177 (N_5177,N_4886,N_4845);
xor U5178 (N_5178,N_4844,N_4848);
nand U5179 (N_5179,N_4995,N_4973);
and U5180 (N_5180,N_4827,N_4966);
or U5181 (N_5181,N_4834,N_4800);
nor U5182 (N_5182,N_4996,N_4937);
or U5183 (N_5183,N_4905,N_4869);
and U5184 (N_5184,N_4928,N_4922);
nor U5185 (N_5185,N_4810,N_4805);
nor U5186 (N_5186,N_4959,N_4968);
nand U5187 (N_5187,N_4984,N_4904);
and U5188 (N_5188,N_4976,N_4888);
nand U5189 (N_5189,N_4926,N_4907);
xnor U5190 (N_5190,N_4852,N_4944);
and U5191 (N_5191,N_4986,N_4989);
xnor U5192 (N_5192,N_4958,N_4858);
nor U5193 (N_5193,N_4866,N_4954);
xor U5194 (N_5194,N_4953,N_4939);
and U5195 (N_5195,N_4861,N_4806);
and U5196 (N_5196,N_4948,N_4922);
nor U5197 (N_5197,N_4858,N_4946);
xnor U5198 (N_5198,N_4830,N_4989);
or U5199 (N_5199,N_4814,N_4866);
nor U5200 (N_5200,N_5068,N_5013);
nand U5201 (N_5201,N_5195,N_5040);
and U5202 (N_5202,N_5095,N_5113);
xnor U5203 (N_5203,N_5093,N_5119);
xnor U5204 (N_5204,N_5138,N_5059);
nor U5205 (N_5205,N_5014,N_5146);
nor U5206 (N_5206,N_5157,N_5151);
or U5207 (N_5207,N_5050,N_5159);
xnor U5208 (N_5208,N_5112,N_5190);
nor U5209 (N_5209,N_5103,N_5106);
nand U5210 (N_5210,N_5011,N_5169);
xnor U5211 (N_5211,N_5060,N_5006);
and U5212 (N_5212,N_5069,N_5086);
xor U5213 (N_5213,N_5049,N_5100);
or U5214 (N_5214,N_5188,N_5063);
nor U5215 (N_5215,N_5118,N_5134);
nor U5216 (N_5216,N_5171,N_5167);
nor U5217 (N_5217,N_5066,N_5038);
nor U5218 (N_5218,N_5192,N_5085);
or U5219 (N_5219,N_5012,N_5129);
nor U5220 (N_5220,N_5136,N_5065);
and U5221 (N_5221,N_5110,N_5022);
nand U5222 (N_5222,N_5116,N_5035);
and U5223 (N_5223,N_5015,N_5133);
nor U5224 (N_5224,N_5183,N_5185);
nor U5225 (N_5225,N_5073,N_5010);
or U5226 (N_5226,N_5178,N_5111);
and U5227 (N_5227,N_5021,N_5131);
and U5228 (N_5228,N_5024,N_5132);
or U5229 (N_5229,N_5028,N_5036);
nand U5230 (N_5230,N_5124,N_5117);
nand U5231 (N_5231,N_5142,N_5189);
nor U5232 (N_5232,N_5099,N_5109);
or U5233 (N_5233,N_5054,N_5091);
nor U5234 (N_5234,N_5139,N_5166);
xor U5235 (N_5235,N_5191,N_5017);
nand U5236 (N_5236,N_5078,N_5122);
and U5237 (N_5237,N_5046,N_5172);
xnor U5238 (N_5238,N_5016,N_5168);
and U5239 (N_5239,N_5061,N_5067);
nand U5240 (N_5240,N_5039,N_5076);
nand U5241 (N_5241,N_5077,N_5009);
nand U5242 (N_5242,N_5184,N_5026);
nand U5243 (N_5243,N_5080,N_5072);
or U5244 (N_5244,N_5096,N_5162);
nor U5245 (N_5245,N_5181,N_5030);
and U5246 (N_5246,N_5057,N_5175);
nand U5247 (N_5247,N_5186,N_5003);
nand U5248 (N_5248,N_5197,N_5149);
xnor U5249 (N_5249,N_5164,N_5165);
xnor U5250 (N_5250,N_5089,N_5156);
nand U5251 (N_5251,N_5051,N_5005);
or U5252 (N_5252,N_5135,N_5155);
and U5253 (N_5253,N_5092,N_5081);
and U5254 (N_5254,N_5043,N_5158);
nor U5255 (N_5255,N_5120,N_5031);
and U5256 (N_5256,N_5056,N_5048);
nand U5257 (N_5257,N_5034,N_5199);
xor U5258 (N_5258,N_5144,N_5102);
or U5259 (N_5259,N_5090,N_5071);
or U5260 (N_5260,N_5105,N_5141);
nor U5261 (N_5261,N_5152,N_5170);
xnor U5262 (N_5262,N_5115,N_5121);
nand U5263 (N_5263,N_5193,N_5196);
and U5264 (N_5264,N_5161,N_5033);
or U5265 (N_5265,N_5023,N_5198);
nand U5266 (N_5266,N_5020,N_5177);
or U5267 (N_5267,N_5176,N_5145);
or U5268 (N_5268,N_5107,N_5041);
and U5269 (N_5269,N_5008,N_5083);
nand U5270 (N_5270,N_5032,N_5174);
or U5271 (N_5271,N_5097,N_5148);
nor U5272 (N_5272,N_5094,N_5088);
or U5273 (N_5273,N_5001,N_5150);
or U5274 (N_5274,N_5182,N_5058);
nor U5275 (N_5275,N_5101,N_5163);
nor U5276 (N_5276,N_5128,N_5147);
nand U5277 (N_5277,N_5062,N_5153);
or U5278 (N_5278,N_5187,N_5127);
xor U5279 (N_5279,N_5037,N_5104);
and U5280 (N_5280,N_5087,N_5143);
xnor U5281 (N_5281,N_5052,N_5045);
and U5282 (N_5282,N_5194,N_5114);
or U5283 (N_5283,N_5018,N_5082);
nor U5284 (N_5284,N_5130,N_5098);
nor U5285 (N_5285,N_5004,N_5042);
or U5286 (N_5286,N_5173,N_5064);
and U5287 (N_5287,N_5084,N_5125);
or U5288 (N_5288,N_5027,N_5179);
nand U5289 (N_5289,N_5137,N_5070);
or U5290 (N_5290,N_5075,N_5029);
and U5291 (N_5291,N_5123,N_5180);
and U5292 (N_5292,N_5002,N_5055);
nand U5293 (N_5293,N_5019,N_5108);
nand U5294 (N_5294,N_5025,N_5000);
and U5295 (N_5295,N_5140,N_5044);
or U5296 (N_5296,N_5047,N_5160);
xnor U5297 (N_5297,N_5007,N_5053);
and U5298 (N_5298,N_5154,N_5079);
nor U5299 (N_5299,N_5074,N_5126);
or U5300 (N_5300,N_5082,N_5069);
xnor U5301 (N_5301,N_5184,N_5158);
nand U5302 (N_5302,N_5003,N_5085);
nand U5303 (N_5303,N_5086,N_5003);
nand U5304 (N_5304,N_5158,N_5055);
xnor U5305 (N_5305,N_5117,N_5173);
or U5306 (N_5306,N_5116,N_5164);
nand U5307 (N_5307,N_5103,N_5154);
xor U5308 (N_5308,N_5031,N_5194);
nor U5309 (N_5309,N_5107,N_5095);
xor U5310 (N_5310,N_5174,N_5144);
and U5311 (N_5311,N_5162,N_5041);
and U5312 (N_5312,N_5176,N_5118);
or U5313 (N_5313,N_5169,N_5080);
and U5314 (N_5314,N_5090,N_5150);
and U5315 (N_5315,N_5154,N_5077);
and U5316 (N_5316,N_5109,N_5174);
or U5317 (N_5317,N_5022,N_5178);
and U5318 (N_5318,N_5166,N_5046);
nand U5319 (N_5319,N_5182,N_5144);
nor U5320 (N_5320,N_5017,N_5057);
and U5321 (N_5321,N_5049,N_5174);
nor U5322 (N_5322,N_5170,N_5044);
nor U5323 (N_5323,N_5106,N_5014);
or U5324 (N_5324,N_5144,N_5087);
nand U5325 (N_5325,N_5111,N_5196);
or U5326 (N_5326,N_5025,N_5140);
and U5327 (N_5327,N_5164,N_5151);
or U5328 (N_5328,N_5070,N_5181);
xnor U5329 (N_5329,N_5005,N_5098);
nor U5330 (N_5330,N_5132,N_5058);
xnor U5331 (N_5331,N_5158,N_5136);
and U5332 (N_5332,N_5022,N_5040);
nor U5333 (N_5333,N_5135,N_5080);
xnor U5334 (N_5334,N_5125,N_5183);
xnor U5335 (N_5335,N_5196,N_5137);
nand U5336 (N_5336,N_5068,N_5175);
or U5337 (N_5337,N_5056,N_5176);
nor U5338 (N_5338,N_5118,N_5186);
nor U5339 (N_5339,N_5156,N_5193);
nor U5340 (N_5340,N_5104,N_5187);
nor U5341 (N_5341,N_5045,N_5147);
or U5342 (N_5342,N_5061,N_5108);
xor U5343 (N_5343,N_5072,N_5091);
xor U5344 (N_5344,N_5095,N_5022);
nand U5345 (N_5345,N_5094,N_5011);
or U5346 (N_5346,N_5054,N_5130);
nor U5347 (N_5347,N_5038,N_5157);
and U5348 (N_5348,N_5177,N_5161);
nor U5349 (N_5349,N_5011,N_5111);
xnor U5350 (N_5350,N_5063,N_5073);
and U5351 (N_5351,N_5096,N_5027);
nand U5352 (N_5352,N_5102,N_5170);
or U5353 (N_5353,N_5016,N_5160);
xor U5354 (N_5354,N_5100,N_5000);
nand U5355 (N_5355,N_5080,N_5079);
and U5356 (N_5356,N_5081,N_5197);
or U5357 (N_5357,N_5101,N_5074);
nand U5358 (N_5358,N_5069,N_5085);
nor U5359 (N_5359,N_5083,N_5197);
nor U5360 (N_5360,N_5013,N_5171);
nand U5361 (N_5361,N_5145,N_5153);
xnor U5362 (N_5362,N_5127,N_5145);
nor U5363 (N_5363,N_5138,N_5187);
or U5364 (N_5364,N_5159,N_5031);
nand U5365 (N_5365,N_5074,N_5149);
nor U5366 (N_5366,N_5072,N_5154);
xnor U5367 (N_5367,N_5131,N_5133);
and U5368 (N_5368,N_5004,N_5035);
xnor U5369 (N_5369,N_5026,N_5122);
or U5370 (N_5370,N_5039,N_5108);
or U5371 (N_5371,N_5074,N_5094);
nor U5372 (N_5372,N_5180,N_5155);
xor U5373 (N_5373,N_5028,N_5092);
and U5374 (N_5374,N_5078,N_5094);
or U5375 (N_5375,N_5092,N_5124);
and U5376 (N_5376,N_5048,N_5151);
and U5377 (N_5377,N_5102,N_5112);
or U5378 (N_5378,N_5046,N_5064);
or U5379 (N_5379,N_5146,N_5151);
xnor U5380 (N_5380,N_5175,N_5059);
nor U5381 (N_5381,N_5056,N_5059);
or U5382 (N_5382,N_5073,N_5091);
or U5383 (N_5383,N_5095,N_5059);
or U5384 (N_5384,N_5020,N_5134);
and U5385 (N_5385,N_5126,N_5168);
xnor U5386 (N_5386,N_5091,N_5140);
or U5387 (N_5387,N_5055,N_5106);
or U5388 (N_5388,N_5097,N_5150);
nand U5389 (N_5389,N_5159,N_5199);
and U5390 (N_5390,N_5153,N_5192);
nor U5391 (N_5391,N_5098,N_5096);
nand U5392 (N_5392,N_5151,N_5093);
or U5393 (N_5393,N_5189,N_5190);
or U5394 (N_5394,N_5057,N_5096);
and U5395 (N_5395,N_5057,N_5183);
xor U5396 (N_5396,N_5056,N_5026);
and U5397 (N_5397,N_5102,N_5008);
nor U5398 (N_5398,N_5180,N_5064);
xor U5399 (N_5399,N_5083,N_5109);
or U5400 (N_5400,N_5381,N_5325);
and U5401 (N_5401,N_5361,N_5277);
and U5402 (N_5402,N_5353,N_5370);
nor U5403 (N_5403,N_5318,N_5363);
and U5404 (N_5404,N_5305,N_5265);
and U5405 (N_5405,N_5299,N_5391);
nor U5406 (N_5406,N_5252,N_5220);
nor U5407 (N_5407,N_5234,N_5289);
nand U5408 (N_5408,N_5319,N_5328);
nor U5409 (N_5409,N_5254,N_5267);
xnor U5410 (N_5410,N_5323,N_5230);
and U5411 (N_5411,N_5285,N_5296);
and U5412 (N_5412,N_5287,N_5340);
xnor U5413 (N_5413,N_5205,N_5384);
and U5414 (N_5414,N_5348,N_5284);
or U5415 (N_5415,N_5240,N_5311);
nor U5416 (N_5416,N_5337,N_5209);
nor U5417 (N_5417,N_5207,N_5360);
or U5418 (N_5418,N_5236,N_5274);
and U5419 (N_5419,N_5359,N_5243);
xor U5420 (N_5420,N_5395,N_5259);
xor U5421 (N_5421,N_5344,N_5366);
xnor U5422 (N_5422,N_5333,N_5309);
nor U5423 (N_5423,N_5253,N_5354);
xor U5424 (N_5424,N_5387,N_5339);
nand U5425 (N_5425,N_5203,N_5390);
or U5426 (N_5426,N_5316,N_5281);
nor U5427 (N_5427,N_5373,N_5218);
or U5428 (N_5428,N_5292,N_5376);
and U5429 (N_5429,N_5394,N_5255);
and U5430 (N_5430,N_5330,N_5298);
nor U5431 (N_5431,N_5278,N_5239);
nor U5432 (N_5432,N_5269,N_5260);
xnor U5433 (N_5433,N_5283,N_5368);
xor U5434 (N_5434,N_5202,N_5241);
xor U5435 (N_5435,N_5228,N_5242);
nor U5436 (N_5436,N_5399,N_5335);
xnor U5437 (N_5437,N_5338,N_5379);
xnor U5438 (N_5438,N_5317,N_5237);
nand U5439 (N_5439,N_5273,N_5372);
and U5440 (N_5440,N_5275,N_5227);
nor U5441 (N_5441,N_5276,N_5225);
and U5442 (N_5442,N_5375,N_5272);
nor U5443 (N_5443,N_5336,N_5392);
nor U5444 (N_5444,N_5221,N_5223);
or U5445 (N_5445,N_5201,N_5343);
xor U5446 (N_5446,N_5367,N_5369);
xnor U5447 (N_5447,N_5219,N_5248);
xor U5448 (N_5448,N_5294,N_5385);
nand U5449 (N_5449,N_5374,N_5295);
nand U5450 (N_5450,N_5364,N_5261);
and U5451 (N_5451,N_5380,N_5245);
and U5452 (N_5452,N_5355,N_5263);
or U5453 (N_5453,N_5282,N_5382);
or U5454 (N_5454,N_5279,N_5217);
and U5455 (N_5455,N_5206,N_5347);
or U5456 (N_5456,N_5341,N_5280);
and U5457 (N_5457,N_5334,N_5352);
nand U5458 (N_5458,N_5329,N_5262);
or U5459 (N_5459,N_5350,N_5214);
and U5460 (N_5460,N_5371,N_5257);
and U5461 (N_5461,N_5356,N_5246);
nand U5462 (N_5462,N_5216,N_5320);
xnor U5463 (N_5463,N_5250,N_5268);
nand U5464 (N_5464,N_5291,N_5313);
and U5465 (N_5465,N_5212,N_5226);
nor U5466 (N_5466,N_5232,N_5393);
nor U5467 (N_5467,N_5321,N_5342);
or U5468 (N_5468,N_5210,N_5386);
or U5469 (N_5469,N_5271,N_5327);
or U5470 (N_5470,N_5208,N_5362);
or U5471 (N_5471,N_5358,N_5270);
and U5472 (N_5472,N_5301,N_5258);
or U5473 (N_5473,N_5286,N_5383);
and U5474 (N_5474,N_5247,N_5251);
nand U5475 (N_5475,N_5326,N_5332);
xnor U5476 (N_5476,N_5377,N_5244);
or U5477 (N_5477,N_5293,N_5231);
and U5478 (N_5478,N_5357,N_5314);
xor U5479 (N_5479,N_5398,N_5378);
xor U5480 (N_5480,N_5389,N_5264);
nor U5481 (N_5481,N_5351,N_5233);
nand U5482 (N_5482,N_5310,N_5229);
nand U5483 (N_5483,N_5324,N_5249);
or U5484 (N_5484,N_5256,N_5211);
nand U5485 (N_5485,N_5315,N_5204);
xnor U5486 (N_5486,N_5312,N_5307);
xnor U5487 (N_5487,N_5290,N_5235);
nor U5488 (N_5488,N_5345,N_5308);
nand U5489 (N_5489,N_5306,N_5297);
xnor U5490 (N_5490,N_5266,N_5331);
or U5491 (N_5491,N_5303,N_5388);
xor U5492 (N_5492,N_5346,N_5322);
xnor U5493 (N_5493,N_5300,N_5365);
nand U5494 (N_5494,N_5238,N_5222);
and U5495 (N_5495,N_5215,N_5288);
and U5496 (N_5496,N_5397,N_5302);
xnor U5497 (N_5497,N_5396,N_5213);
or U5498 (N_5498,N_5304,N_5349);
and U5499 (N_5499,N_5200,N_5224);
and U5500 (N_5500,N_5229,N_5240);
xor U5501 (N_5501,N_5256,N_5325);
and U5502 (N_5502,N_5390,N_5384);
or U5503 (N_5503,N_5282,N_5244);
xor U5504 (N_5504,N_5360,N_5314);
nor U5505 (N_5505,N_5298,N_5355);
nand U5506 (N_5506,N_5320,N_5361);
or U5507 (N_5507,N_5306,N_5288);
or U5508 (N_5508,N_5210,N_5207);
nor U5509 (N_5509,N_5200,N_5347);
and U5510 (N_5510,N_5268,N_5337);
xnor U5511 (N_5511,N_5304,N_5360);
or U5512 (N_5512,N_5235,N_5250);
or U5513 (N_5513,N_5269,N_5284);
nor U5514 (N_5514,N_5235,N_5207);
xor U5515 (N_5515,N_5295,N_5354);
and U5516 (N_5516,N_5380,N_5221);
nand U5517 (N_5517,N_5237,N_5377);
or U5518 (N_5518,N_5284,N_5253);
nor U5519 (N_5519,N_5390,N_5249);
or U5520 (N_5520,N_5304,N_5384);
and U5521 (N_5521,N_5311,N_5315);
xor U5522 (N_5522,N_5309,N_5290);
nor U5523 (N_5523,N_5365,N_5240);
nand U5524 (N_5524,N_5301,N_5352);
nor U5525 (N_5525,N_5302,N_5383);
or U5526 (N_5526,N_5245,N_5265);
nand U5527 (N_5527,N_5314,N_5239);
and U5528 (N_5528,N_5336,N_5396);
nor U5529 (N_5529,N_5367,N_5256);
and U5530 (N_5530,N_5224,N_5334);
nand U5531 (N_5531,N_5326,N_5288);
nand U5532 (N_5532,N_5232,N_5374);
and U5533 (N_5533,N_5253,N_5379);
and U5534 (N_5534,N_5232,N_5245);
and U5535 (N_5535,N_5203,N_5339);
xnor U5536 (N_5536,N_5376,N_5318);
xor U5537 (N_5537,N_5256,N_5329);
xor U5538 (N_5538,N_5311,N_5297);
and U5539 (N_5539,N_5215,N_5373);
xor U5540 (N_5540,N_5368,N_5261);
nor U5541 (N_5541,N_5289,N_5388);
and U5542 (N_5542,N_5301,N_5330);
or U5543 (N_5543,N_5234,N_5299);
and U5544 (N_5544,N_5303,N_5333);
nor U5545 (N_5545,N_5286,N_5222);
nand U5546 (N_5546,N_5337,N_5266);
and U5547 (N_5547,N_5220,N_5335);
nand U5548 (N_5548,N_5266,N_5305);
nand U5549 (N_5549,N_5381,N_5369);
or U5550 (N_5550,N_5299,N_5365);
or U5551 (N_5551,N_5216,N_5305);
nand U5552 (N_5552,N_5290,N_5276);
or U5553 (N_5553,N_5320,N_5232);
or U5554 (N_5554,N_5233,N_5256);
nor U5555 (N_5555,N_5326,N_5282);
nand U5556 (N_5556,N_5328,N_5356);
nor U5557 (N_5557,N_5314,N_5243);
xnor U5558 (N_5558,N_5326,N_5255);
and U5559 (N_5559,N_5218,N_5239);
xnor U5560 (N_5560,N_5249,N_5277);
nand U5561 (N_5561,N_5346,N_5327);
and U5562 (N_5562,N_5236,N_5206);
or U5563 (N_5563,N_5390,N_5381);
xnor U5564 (N_5564,N_5208,N_5348);
and U5565 (N_5565,N_5232,N_5312);
or U5566 (N_5566,N_5216,N_5399);
and U5567 (N_5567,N_5228,N_5249);
or U5568 (N_5568,N_5378,N_5250);
nand U5569 (N_5569,N_5299,N_5399);
xnor U5570 (N_5570,N_5316,N_5347);
xor U5571 (N_5571,N_5203,N_5270);
nor U5572 (N_5572,N_5203,N_5334);
nor U5573 (N_5573,N_5280,N_5268);
xnor U5574 (N_5574,N_5397,N_5206);
and U5575 (N_5575,N_5368,N_5222);
and U5576 (N_5576,N_5292,N_5314);
xor U5577 (N_5577,N_5308,N_5246);
and U5578 (N_5578,N_5217,N_5243);
and U5579 (N_5579,N_5297,N_5331);
nand U5580 (N_5580,N_5274,N_5279);
or U5581 (N_5581,N_5326,N_5388);
nor U5582 (N_5582,N_5274,N_5229);
or U5583 (N_5583,N_5228,N_5238);
nand U5584 (N_5584,N_5397,N_5211);
nand U5585 (N_5585,N_5311,N_5320);
xnor U5586 (N_5586,N_5262,N_5266);
xnor U5587 (N_5587,N_5304,N_5270);
xor U5588 (N_5588,N_5352,N_5306);
and U5589 (N_5589,N_5200,N_5220);
nand U5590 (N_5590,N_5361,N_5325);
and U5591 (N_5591,N_5386,N_5370);
or U5592 (N_5592,N_5322,N_5238);
xor U5593 (N_5593,N_5379,N_5231);
or U5594 (N_5594,N_5276,N_5210);
and U5595 (N_5595,N_5226,N_5245);
or U5596 (N_5596,N_5280,N_5331);
or U5597 (N_5597,N_5212,N_5325);
nor U5598 (N_5598,N_5237,N_5333);
xor U5599 (N_5599,N_5366,N_5236);
and U5600 (N_5600,N_5521,N_5538);
nor U5601 (N_5601,N_5465,N_5466);
xnor U5602 (N_5602,N_5586,N_5529);
xor U5603 (N_5603,N_5594,N_5578);
nand U5604 (N_5604,N_5432,N_5581);
or U5605 (N_5605,N_5498,N_5520);
or U5606 (N_5606,N_5468,N_5429);
nor U5607 (N_5607,N_5407,N_5588);
and U5608 (N_5608,N_5557,N_5572);
nand U5609 (N_5609,N_5471,N_5478);
xnor U5610 (N_5610,N_5585,N_5583);
xnor U5611 (N_5611,N_5590,N_5431);
nor U5612 (N_5612,N_5486,N_5411);
or U5613 (N_5613,N_5592,N_5462);
and U5614 (N_5614,N_5454,N_5460);
xor U5615 (N_5615,N_5464,N_5458);
and U5616 (N_5616,N_5563,N_5558);
nor U5617 (N_5617,N_5409,N_5435);
and U5618 (N_5618,N_5414,N_5404);
and U5619 (N_5619,N_5503,N_5548);
nand U5620 (N_5620,N_5472,N_5420);
nand U5621 (N_5621,N_5576,N_5449);
or U5622 (N_5622,N_5469,N_5412);
nand U5623 (N_5623,N_5452,N_5584);
or U5624 (N_5624,N_5425,N_5443);
xor U5625 (N_5625,N_5509,N_5540);
xor U5626 (N_5626,N_5505,N_5573);
and U5627 (N_5627,N_5568,N_5444);
and U5628 (N_5628,N_5428,N_5492);
and U5629 (N_5629,N_5554,N_5480);
and U5630 (N_5630,N_5457,N_5542);
xor U5631 (N_5631,N_5560,N_5489);
or U5632 (N_5632,N_5516,N_5439);
nor U5633 (N_5633,N_5456,N_5490);
or U5634 (N_5634,N_5528,N_5484);
nor U5635 (N_5635,N_5419,N_5418);
nand U5636 (N_5636,N_5559,N_5587);
nor U5637 (N_5637,N_5499,N_5427);
nand U5638 (N_5638,N_5546,N_5422);
and U5639 (N_5639,N_5589,N_5596);
and U5640 (N_5640,N_5524,N_5525);
or U5641 (N_5641,N_5481,N_5582);
xnor U5642 (N_5642,N_5562,N_5434);
or U5643 (N_5643,N_5436,N_5598);
nor U5644 (N_5644,N_5569,N_5544);
xor U5645 (N_5645,N_5593,N_5513);
xor U5646 (N_5646,N_5410,N_5580);
xor U5647 (N_5647,N_5566,N_5523);
or U5648 (N_5648,N_5553,N_5506);
or U5649 (N_5649,N_5597,N_5599);
and U5650 (N_5650,N_5496,N_5474);
nor U5651 (N_5651,N_5423,N_5522);
xor U5652 (N_5652,N_5406,N_5417);
and U5653 (N_5653,N_5438,N_5403);
nand U5654 (N_5654,N_5487,N_5441);
nand U5655 (N_5655,N_5477,N_5476);
or U5656 (N_5656,N_5530,N_5534);
nor U5657 (N_5657,N_5401,N_5470);
xnor U5658 (N_5658,N_5519,N_5459);
or U5659 (N_5659,N_5448,N_5555);
nor U5660 (N_5660,N_5400,N_5450);
or U5661 (N_5661,N_5491,N_5442);
nor U5662 (N_5662,N_5440,N_5446);
or U5663 (N_5663,N_5539,N_5531);
or U5664 (N_5664,N_5536,N_5543);
or U5665 (N_5665,N_5502,N_5550);
nand U5666 (N_5666,N_5433,N_5494);
nand U5667 (N_5667,N_5512,N_5493);
and U5668 (N_5668,N_5482,N_5416);
xnor U5669 (N_5669,N_5511,N_5475);
and U5670 (N_5670,N_5500,N_5445);
nor U5671 (N_5671,N_5527,N_5571);
nor U5672 (N_5672,N_5437,N_5415);
nand U5673 (N_5673,N_5561,N_5507);
nand U5674 (N_5674,N_5461,N_5495);
nand U5675 (N_5675,N_5537,N_5567);
or U5676 (N_5676,N_5575,N_5421);
nor U5677 (N_5677,N_5591,N_5552);
xnor U5678 (N_5678,N_5515,N_5579);
and U5679 (N_5679,N_5526,N_5453);
nand U5680 (N_5680,N_5564,N_5485);
or U5681 (N_5681,N_5405,N_5545);
or U5682 (N_5682,N_5547,N_5532);
nor U5683 (N_5683,N_5424,N_5501);
and U5684 (N_5684,N_5565,N_5463);
nand U5685 (N_5685,N_5549,N_5430);
or U5686 (N_5686,N_5504,N_5447);
nand U5687 (N_5687,N_5467,N_5426);
or U5688 (N_5688,N_5570,N_5556);
xor U5689 (N_5689,N_5517,N_5574);
nor U5690 (N_5690,N_5541,N_5535);
xor U5691 (N_5691,N_5408,N_5577);
and U5692 (N_5692,N_5455,N_5551);
nor U5693 (N_5693,N_5402,N_5595);
or U5694 (N_5694,N_5473,N_5488);
or U5695 (N_5695,N_5451,N_5533);
nor U5696 (N_5696,N_5514,N_5518);
or U5697 (N_5697,N_5479,N_5483);
nand U5698 (N_5698,N_5497,N_5413);
nand U5699 (N_5699,N_5508,N_5510);
and U5700 (N_5700,N_5433,N_5531);
xor U5701 (N_5701,N_5450,N_5465);
xor U5702 (N_5702,N_5462,N_5508);
and U5703 (N_5703,N_5528,N_5558);
nand U5704 (N_5704,N_5459,N_5497);
nor U5705 (N_5705,N_5428,N_5462);
nor U5706 (N_5706,N_5442,N_5544);
nand U5707 (N_5707,N_5456,N_5581);
or U5708 (N_5708,N_5573,N_5570);
nand U5709 (N_5709,N_5415,N_5502);
xnor U5710 (N_5710,N_5506,N_5411);
nor U5711 (N_5711,N_5526,N_5597);
nand U5712 (N_5712,N_5437,N_5470);
nand U5713 (N_5713,N_5469,N_5514);
xnor U5714 (N_5714,N_5416,N_5525);
and U5715 (N_5715,N_5527,N_5518);
and U5716 (N_5716,N_5526,N_5496);
or U5717 (N_5717,N_5446,N_5495);
or U5718 (N_5718,N_5402,N_5589);
xor U5719 (N_5719,N_5420,N_5419);
xnor U5720 (N_5720,N_5438,N_5597);
or U5721 (N_5721,N_5478,N_5465);
nor U5722 (N_5722,N_5583,N_5527);
and U5723 (N_5723,N_5507,N_5526);
xnor U5724 (N_5724,N_5474,N_5500);
or U5725 (N_5725,N_5541,N_5481);
and U5726 (N_5726,N_5425,N_5455);
and U5727 (N_5727,N_5457,N_5444);
nand U5728 (N_5728,N_5557,N_5548);
or U5729 (N_5729,N_5539,N_5589);
and U5730 (N_5730,N_5471,N_5429);
xnor U5731 (N_5731,N_5436,N_5553);
nor U5732 (N_5732,N_5504,N_5412);
xor U5733 (N_5733,N_5562,N_5487);
nand U5734 (N_5734,N_5511,N_5523);
or U5735 (N_5735,N_5501,N_5549);
or U5736 (N_5736,N_5582,N_5505);
nor U5737 (N_5737,N_5595,N_5561);
xnor U5738 (N_5738,N_5438,N_5583);
or U5739 (N_5739,N_5555,N_5540);
or U5740 (N_5740,N_5597,N_5489);
nand U5741 (N_5741,N_5403,N_5414);
nand U5742 (N_5742,N_5562,N_5479);
nor U5743 (N_5743,N_5573,N_5467);
or U5744 (N_5744,N_5424,N_5529);
or U5745 (N_5745,N_5466,N_5548);
nor U5746 (N_5746,N_5522,N_5462);
nor U5747 (N_5747,N_5577,N_5548);
nor U5748 (N_5748,N_5402,N_5554);
and U5749 (N_5749,N_5438,N_5468);
nand U5750 (N_5750,N_5449,N_5503);
nor U5751 (N_5751,N_5529,N_5499);
nor U5752 (N_5752,N_5572,N_5535);
xnor U5753 (N_5753,N_5544,N_5460);
or U5754 (N_5754,N_5501,N_5521);
nand U5755 (N_5755,N_5533,N_5437);
or U5756 (N_5756,N_5561,N_5543);
or U5757 (N_5757,N_5415,N_5511);
nor U5758 (N_5758,N_5564,N_5486);
nor U5759 (N_5759,N_5567,N_5578);
or U5760 (N_5760,N_5444,N_5410);
nor U5761 (N_5761,N_5478,N_5500);
xor U5762 (N_5762,N_5470,N_5504);
nor U5763 (N_5763,N_5411,N_5433);
or U5764 (N_5764,N_5440,N_5434);
and U5765 (N_5765,N_5556,N_5475);
or U5766 (N_5766,N_5501,N_5529);
or U5767 (N_5767,N_5555,N_5439);
xor U5768 (N_5768,N_5496,N_5448);
and U5769 (N_5769,N_5497,N_5487);
or U5770 (N_5770,N_5411,N_5521);
or U5771 (N_5771,N_5495,N_5468);
nor U5772 (N_5772,N_5402,N_5502);
or U5773 (N_5773,N_5425,N_5409);
nand U5774 (N_5774,N_5423,N_5513);
or U5775 (N_5775,N_5464,N_5489);
xnor U5776 (N_5776,N_5462,N_5582);
nand U5777 (N_5777,N_5419,N_5421);
nor U5778 (N_5778,N_5438,N_5542);
nor U5779 (N_5779,N_5529,N_5525);
or U5780 (N_5780,N_5511,N_5419);
xor U5781 (N_5781,N_5538,N_5465);
nand U5782 (N_5782,N_5568,N_5421);
xor U5783 (N_5783,N_5478,N_5486);
and U5784 (N_5784,N_5543,N_5504);
nor U5785 (N_5785,N_5491,N_5539);
nand U5786 (N_5786,N_5530,N_5478);
or U5787 (N_5787,N_5457,N_5536);
nand U5788 (N_5788,N_5536,N_5529);
nor U5789 (N_5789,N_5587,N_5504);
nand U5790 (N_5790,N_5494,N_5487);
or U5791 (N_5791,N_5514,N_5546);
nand U5792 (N_5792,N_5574,N_5459);
nand U5793 (N_5793,N_5457,N_5423);
nand U5794 (N_5794,N_5542,N_5524);
nand U5795 (N_5795,N_5549,N_5424);
nor U5796 (N_5796,N_5454,N_5597);
or U5797 (N_5797,N_5580,N_5587);
and U5798 (N_5798,N_5511,N_5553);
and U5799 (N_5799,N_5449,N_5509);
or U5800 (N_5800,N_5704,N_5649);
or U5801 (N_5801,N_5658,N_5625);
nand U5802 (N_5802,N_5700,N_5622);
or U5803 (N_5803,N_5641,N_5750);
nor U5804 (N_5804,N_5745,N_5682);
nor U5805 (N_5805,N_5733,N_5674);
xor U5806 (N_5806,N_5784,N_5762);
or U5807 (N_5807,N_5719,N_5794);
nand U5808 (N_5808,N_5611,N_5739);
nand U5809 (N_5809,N_5721,N_5787);
or U5810 (N_5810,N_5683,N_5647);
or U5811 (N_5811,N_5706,N_5650);
or U5812 (N_5812,N_5757,N_5747);
or U5813 (N_5813,N_5772,N_5723);
nor U5814 (N_5814,N_5636,N_5709);
or U5815 (N_5815,N_5640,N_5618);
or U5816 (N_5816,N_5604,N_5613);
and U5817 (N_5817,N_5761,N_5659);
and U5818 (N_5818,N_5755,N_5769);
nand U5819 (N_5819,N_5631,N_5705);
nor U5820 (N_5820,N_5616,N_5760);
xor U5821 (N_5821,N_5736,N_5718);
nor U5822 (N_5822,N_5672,N_5667);
or U5823 (N_5823,N_5766,N_5795);
and U5824 (N_5824,N_5738,N_5730);
nand U5825 (N_5825,N_5661,N_5741);
and U5826 (N_5826,N_5786,N_5715);
nand U5827 (N_5827,N_5644,N_5756);
nand U5828 (N_5828,N_5639,N_5782);
and U5829 (N_5829,N_5790,N_5798);
nand U5830 (N_5830,N_5792,N_5734);
nand U5831 (N_5831,N_5724,N_5701);
nor U5832 (N_5832,N_5785,N_5780);
nor U5833 (N_5833,N_5764,N_5679);
nor U5834 (N_5834,N_5702,N_5717);
and U5835 (N_5835,N_5758,N_5713);
or U5836 (N_5836,N_5686,N_5751);
xnor U5837 (N_5837,N_5694,N_5765);
nand U5838 (N_5838,N_5699,N_5778);
nor U5839 (N_5839,N_5633,N_5722);
xor U5840 (N_5840,N_5609,N_5742);
nand U5841 (N_5841,N_5793,N_5774);
nor U5842 (N_5842,N_5749,N_5768);
or U5843 (N_5843,N_5695,N_5729);
or U5844 (N_5844,N_5690,N_5720);
xor U5845 (N_5845,N_5703,N_5668);
and U5846 (N_5846,N_5692,N_5678);
nand U5847 (N_5847,N_5797,N_5681);
xnor U5848 (N_5848,N_5687,N_5677);
xor U5849 (N_5849,N_5624,N_5691);
nor U5850 (N_5850,N_5669,N_5771);
or U5851 (N_5851,N_5726,N_5783);
or U5852 (N_5852,N_5693,N_5752);
nand U5853 (N_5853,N_5642,N_5754);
nor U5854 (N_5854,N_5711,N_5608);
or U5855 (N_5855,N_5619,N_5653);
xor U5856 (N_5856,N_5728,N_5670);
xor U5857 (N_5857,N_5791,N_5666);
xnor U5858 (N_5858,N_5620,N_5732);
xnor U5859 (N_5859,N_5662,N_5621);
xor U5860 (N_5860,N_5708,N_5744);
nand U5861 (N_5861,N_5684,N_5646);
and U5862 (N_5862,N_5637,N_5656);
xnor U5863 (N_5863,N_5652,N_5660);
and U5864 (N_5864,N_5776,N_5602);
or U5865 (N_5865,N_5796,N_5601);
nand U5866 (N_5866,N_5731,N_5767);
xor U5867 (N_5867,N_5638,N_5688);
and U5868 (N_5868,N_5763,N_5696);
xor U5869 (N_5869,N_5770,N_5725);
nor U5870 (N_5870,N_5740,N_5712);
nor U5871 (N_5871,N_5676,N_5628);
and U5872 (N_5872,N_5735,N_5663);
xor U5873 (N_5873,N_5654,N_5675);
or U5874 (N_5874,N_5665,N_5603);
xnor U5875 (N_5875,N_5612,N_5707);
or U5876 (N_5876,N_5664,N_5775);
and U5877 (N_5877,N_5737,N_5610);
or U5878 (N_5878,N_5779,N_5788);
nor U5879 (N_5879,N_5629,N_5605);
or U5880 (N_5880,N_5689,N_5773);
nor U5881 (N_5881,N_5606,N_5748);
and U5882 (N_5882,N_5746,N_5607);
and U5883 (N_5883,N_5643,N_5671);
nor U5884 (N_5884,N_5685,N_5651);
xnor U5885 (N_5885,N_5645,N_5799);
nand U5886 (N_5886,N_5615,N_5714);
and U5887 (N_5887,N_5635,N_5634);
nand U5888 (N_5888,N_5743,N_5716);
nor U5889 (N_5889,N_5710,N_5680);
nand U5890 (N_5890,N_5626,N_5623);
and U5891 (N_5891,N_5753,N_5632);
or U5892 (N_5892,N_5614,N_5789);
or U5893 (N_5893,N_5698,N_5648);
or U5894 (N_5894,N_5600,N_5727);
nor U5895 (N_5895,N_5627,N_5617);
xor U5896 (N_5896,N_5655,N_5630);
nor U5897 (N_5897,N_5697,N_5673);
and U5898 (N_5898,N_5657,N_5777);
xnor U5899 (N_5899,N_5759,N_5781);
xor U5900 (N_5900,N_5686,N_5763);
or U5901 (N_5901,N_5749,N_5720);
or U5902 (N_5902,N_5652,N_5681);
xor U5903 (N_5903,N_5663,N_5706);
or U5904 (N_5904,N_5673,N_5713);
and U5905 (N_5905,N_5716,N_5663);
and U5906 (N_5906,N_5609,N_5795);
nand U5907 (N_5907,N_5642,N_5709);
and U5908 (N_5908,N_5739,N_5626);
nand U5909 (N_5909,N_5665,N_5664);
or U5910 (N_5910,N_5626,N_5704);
nand U5911 (N_5911,N_5778,N_5617);
nor U5912 (N_5912,N_5656,N_5619);
xor U5913 (N_5913,N_5723,N_5709);
xnor U5914 (N_5914,N_5618,N_5662);
nor U5915 (N_5915,N_5630,N_5738);
or U5916 (N_5916,N_5631,N_5657);
and U5917 (N_5917,N_5703,N_5701);
and U5918 (N_5918,N_5741,N_5787);
nor U5919 (N_5919,N_5685,N_5723);
and U5920 (N_5920,N_5655,N_5751);
and U5921 (N_5921,N_5700,N_5799);
and U5922 (N_5922,N_5794,N_5692);
and U5923 (N_5923,N_5635,N_5757);
and U5924 (N_5924,N_5645,N_5721);
nand U5925 (N_5925,N_5616,N_5788);
or U5926 (N_5926,N_5779,N_5654);
xor U5927 (N_5927,N_5766,N_5662);
or U5928 (N_5928,N_5712,N_5673);
or U5929 (N_5929,N_5704,N_5644);
nor U5930 (N_5930,N_5637,N_5676);
nand U5931 (N_5931,N_5705,N_5733);
nand U5932 (N_5932,N_5654,N_5612);
xnor U5933 (N_5933,N_5646,N_5782);
xnor U5934 (N_5934,N_5607,N_5720);
xnor U5935 (N_5935,N_5735,N_5658);
and U5936 (N_5936,N_5761,N_5627);
nand U5937 (N_5937,N_5680,N_5683);
and U5938 (N_5938,N_5688,N_5719);
or U5939 (N_5939,N_5742,N_5765);
nand U5940 (N_5940,N_5625,N_5731);
nand U5941 (N_5941,N_5696,N_5735);
nand U5942 (N_5942,N_5697,N_5775);
xnor U5943 (N_5943,N_5765,N_5696);
nor U5944 (N_5944,N_5650,N_5713);
or U5945 (N_5945,N_5704,N_5785);
or U5946 (N_5946,N_5719,N_5675);
or U5947 (N_5947,N_5641,N_5774);
nand U5948 (N_5948,N_5649,N_5695);
xor U5949 (N_5949,N_5617,N_5751);
nand U5950 (N_5950,N_5718,N_5627);
xnor U5951 (N_5951,N_5710,N_5672);
nor U5952 (N_5952,N_5729,N_5698);
or U5953 (N_5953,N_5657,N_5740);
xnor U5954 (N_5954,N_5601,N_5762);
nand U5955 (N_5955,N_5797,N_5673);
nor U5956 (N_5956,N_5654,N_5729);
xnor U5957 (N_5957,N_5602,N_5713);
and U5958 (N_5958,N_5633,N_5782);
nand U5959 (N_5959,N_5642,N_5669);
or U5960 (N_5960,N_5726,N_5681);
nor U5961 (N_5961,N_5681,N_5677);
xnor U5962 (N_5962,N_5739,N_5754);
nand U5963 (N_5963,N_5649,N_5779);
or U5964 (N_5964,N_5762,N_5677);
and U5965 (N_5965,N_5757,N_5655);
nand U5966 (N_5966,N_5627,N_5726);
or U5967 (N_5967,N_5607,N_5725);
nor U5968 (N_5968,N_5766,N_5703);
xnor U5969 (N_5969,N_5642,N_5665);
or U5970 (N_5970,N_5738,N_5722);
nor U5971 (N_5971,N_5687,N_5774);
or U5972 (N_5972,N_5698,N_5641);
xor U5973 (N_5973,N_5753,N_5703);
nor U5974 (N_5974,N_5714,N_5620);
xor U5975 (N_5975,N_5619,N_5731);
and U5976 (N_5976,N_5664,N_5694);
nand U5977 (N_5977,N_5755,N_5664);
nand U5978 (N_5978,N_5653,N_5648);
or U5979 (N_5979,N_5717,N_5730);
nor U5980 (N_5980,N_5792,N_5626);
xnor U5981 (N_5981,N_5730,N_5715);
and U5982 (N_5982,N_5761,N_5764);
and U5983 (N_5983,N_5703,N_5775);
nand U5984 (N_5984,N_5675,N_5680);
xnor U5985 (N_5985,N_5728,N_5687);
xor U5986 (N_5986,N_5613,N_5724);
or U5987 (N_5987,N_5698,N_5676);
nor U5988 (N_5988,N_5715,N_5699);
nor U5989 (N_5989,N_5612,N_5772);
nand U5990 (N_5990,N_5754,N_5648);
nor U5991 (N_5991,N_5740,N_5747);
and U5992 (N_5992,N_5768,N_5713);
nor U5993 (N_5993,N_5737,N_5724);
xnor U5994 (N_5994,N_5736,N_5633);
nand U5995 (N_5995,N_5782,N_5677);
or U5996 (N_5996,N_5612,N_5615);
nor U5997 (N_5997,N_5680,N_5657);
nor U5998 (N_5998,N_5756,N_5792);
and U5999 (N_5999,N_5611,N_5629);
or U6000 (N_6000,N_5928,N_5800);
xor U6001 (N_6001,N_5973,N_5916);
xnor U6002 (N_6002,N_5810,N_5837);
or U6003 (N_6003,N_5887,N_5962);
nand U6004 (N_6004,N_5840,N_5874);
and U6005 (N_6005,N_5885,N_5927);
and U6006 (N_6006,N_5960,N_5977);
and U6007 (N_6007,N_5950,N_5831);
and U6008 (N_6008,N_5917,N_5816);
nor U6009 (N_6009,N_5979,N_5937);
xnor U6010 (N_6010,N_5877,N_5825);
xnor U6011 (N_6011,N_5966,N_5861);
or U6012 (N_6012,N_5809,N_5978);
nand U6013 (N_6013,N_5867,N_5898);
and U6014 (N_6014,N_5870,N_5846);
nand U6015 (N_6015,N_5983,N_5972);
and U6016 (N_6016,N_5807,N_5866);
nand U6017 (N_6017,N_5872,N_5929);
or U6018 (N_6018,N_5985,N_5919);
xnor U6019 (N_6019,N_5882,N_5871);
nor U6020 (N_6020,N_5869,N_5967);
and U6021 (N_6021,N_5941,N_5942);
nor U6022 (N_6022,N_5976,N_5954);
and U6023 (N_6023,N_5895,N_5932);
nand U6024 (N_6024,N_5849,N_5828);
nor U6025 (N_6025,N_5819,N_5912);
and U6026 (N_6026,N_5860,N_5995);
xnor U6027 (N_6027,N_5990,N_5881);
or U6028 (N_6028,N_5875,N_5952);
nand U6029 (N_6029,N_5926,N_5832);
nand U6030 (N_6030,N_5879,N_5981);
nand U6031 (N_6031,N_5933,N_5843);
or U6032 (N_6032,N_5984,N_5925);
nand U6033 (N_6033,N_5915,N_5908);
or U6034 (N_6034,N_5901,N_5818);
or U6035 (N_6035,N_5914,N_5988);
and U6036 (N_6036,N_5975,N_5986);
or U6037 (N_6037,N_5913,N_5938);
and U6038 (N_6038,N_5851,N_5994);
and U6039 (N_6039,N_5905,N_5997);
and U6040 (N_6040,N_5808,N_5865);
nor U6041 (N_6041,N_5953,N_5923);
or U6042 (N_6042,N_5827,N_5823);
nor U6043 (N_6043,N_5876,N_5833);
nor U6044 (N_6044,N_5817,N_5811);
or U6045 (N_6045,N_5836,N_5924);
or U6046 (N_6046,N_5963,N_5965);
and U6047 (N_6047,N_5844,N_5884);
xor U6048 (N_6048,N_5839,N_5922);
and U6049 (N_6049,N_5873,N_5974);
nor U6050 (N_6050,N_5803,N_5902);
xnor U6051 (N_6051,N_5852,N_5951);
or U6052 (N_6052,N_5900,N_5920);
or U6053 (N_6053,N_5991,N_5918);
and U6054 (N_6054,N_5804,N_5864);
or U6055 (N_6055,N_5847,N_5940);
and U6056 (N_6056,N_5829,N_5863);
nand U6057 (N_6057,N_5883,N_5930);
nor U6058 (N_6058,N_5909,N_5821);
nor U6059 (N_6059,N_5968,N_5894);
xor U6060 (N_6060,N_5805,N_5957);
xor U6061 (N_6061,N_5959,N_5854);
and U6062 (N_6062,N_5945,N_5853);
or U6063 (N_6063,N_5886,N_5907);
xor U6064 (N_6064,N_5848,N_5834);
nand U6065 (N_6065,N_5862,N_5890);
nand U6066 (N_6066,N_5820,N_5931);
nand U6067 (N_6067,N_5955,N_5964);
and U6068 (N_6068,N_5857,N_5812);
nor U6069 (N_6069,N_5801,N_5856);
nand U6070 (N_6070,N_5893,N_5980);
nand U6071 (N_6071,N_5999,N_5822);
xnor U6072 (N_6072,N_5943,N_5802);
xor U6073 (N_6073,N_5838,N_5904);
xor U6074 (N_6074,N_5996,N_5888);
xnor U6075 (N_6075,N_5958,N_5970);
and U6076 (N_6076,N_5982,N_5992);
xor U6077 (N_6077,N_5998,N_5813);
nand U6078 (N_6078,N_5835,N_5993);
xnor U6079 (N_6079,N_5921,N_5815);
and U6080 (N_6080,N_5936,N_5845);
and U6081 (N_6081,N_5906,N_5910);
and U6082 (N_6082,N_5826,N_5858);
nand U6083 (N_6083,N_5850,N_5859);
nor U6084 (N_6084,N_5899,N_5989);
or U6085 (N_6085,N_5889,N_5903);
and U6086 (N_6086,N_5814,N_5911);
and U6087 (N_6087,N_5934,N_5841);
nand U6088 (N_6088,N_5971,N_5896);
nor U6089 (N_6089,N_5806,N_5891);
or U6090 (N_6090,N_5855,N_5947);
xnor U6091 (N_6091,N_5842,N_5987);
nor U6092 (N_6092,N_5824,N_5956);
nand U6093 (N_6093,N_5868,N_5878);
and U6094 (N_6094,N_5939,N_5949);
and U6095 (N_6095,N_5961,N_5830);
xnor U6096 (N_6096,N_5880,N_5969);
nor U6097 (N_6097,N_5897,N_5935);
and U6098 (N_6098,N_5892,N_5948);
xnor U6099 (N_6099,N_5944,N_5946);
xor U6100 (N_6100,N_5987,N_5997);
and U6101 (N_6101,N_5952,N_5937);
nand U6102 (N_6102,N_5987,N_5918);
nor U6103 (N_6103,N_5883,N_5915);
xnor U6104 (N_6104,N_5807,N_5819);
nor U6105 (N_6105,N_5823,N_5981);
xor U6106 (N_6106,N_5876,N_5845);
nand U6107 (N_6107,N_5905,N_5835);
nand U6108 (N_6108,N_5894,N_5929);
nand U6109 (N_6109,N_5977,N_5839);
and U6110 (N_6110,N_5805,N_5999);
or U6111 (N_6111,N_5815,N_5808);
and U6112 (N_6112,N_5855,N_5815);
nor U6113 (N_6113,N_5946,N_5864);
nand U6114 (N_6114,N_5902,N_5999);
and U6115 (N_6115,N_5947,N_5911);
nor U6116 (N_6116,N_5937,N_5864);
nand U6117 (N_6117,N_5816,N_5859);
or U6118 (N_6118,N_5952,N_5950);
nor U6119 (N_6119,N_5876,N_5852);
xor U6120 (N_6120,N_5824,N_5913);
xor U6121 (N_6121,N_5973,N_5929);
nand U6122 (N_6122,N_5935,N_5982);
nor U6123 (N_6123,N_5984,N_5964);
and U6124 (N_6124,N_5851,N_5950);
and U6125 (N_6125,N_5913,N_5981);
nand U6126 (N_6126,N_5816,N_5978);
xnor U6127 (N_6127,N_5941,N_5976);
and U6128 (N_6128,N_5864,N_5822);
nor U6129 (N_6129,N_5903,N_5807);
nand U6130 (N_6130,N_5862,N_5886);
xnor U6131 (N_6131,N_5815,N_5948);
or U6132 (N_6132,N_5998,N_5972);
nand U6133 (N_6133,N_5874,N_5979);
or U6134 (N_6134,N_5904,N_5901);
xnor U6135 (N_6135,N_5915,N_5854);
nor U6136 (N_6136,N_5988,N_5835);
nand U6137 (N_6137,N_5821,N_5933);
nor U6138 (N_6138,N_5827,N_5978);
and U6139 (N_6139,N_5907,N_5833);
or U6140 (N_6140,N_5964,N_5896);
nand U6141 (N_6141,N_5846,N_5873);
and U6142 (N_6142,N_5801,N_5923);
and U6143 (N_6143,N_5820,N_5968);
nand U6144 (N_6144,N_5908,N_5874);
and U6145 (N_6145,N_5938,N_5800);
nand U6146 (N_6146,N_5857,N_5972);
xor U6147 (N_6147,N_5919,N_5921);
or U6148 (N_6148,N_5933,N_5938);
nand U6149 (N_6149,N_5824,N_5847);
nor U6150 (N_6150,N_5972,N_5884);
and U6151 (N_6151,N_5873,N_5814);
nand U6152 (N_6152,N_5900,N_5853);
nor U6153 (N_6153,N_5895,N_5827);
nor U6154 (N_6154,N_5969,N_5937);
or U6155 (N_6155,N_5924,N_5803);
and U6156 (N_6156,N_5852,N_5815);
nor U6157 (N_6157,N_5822,N_5917);
and U6158 (N_6158,N_5847,N_5930);
nor U6159 (N_6159,N_5927,N_5847);
and U6160 (N_6160,N_5953,N_5859);
or U6161 (N_6161,N_5933,N_5819);
or U6162 (N_6162,N_5934,N_5847);
or U6163 (N_6163,N_5918,N_5875);
nand U6164 (N_6164,N_5943,N_5826);
or U6165 (N_6165,N_5861,N_5836);
nor U6166 (N_6166,N_5958,N_5981);
xnor U6167 (N_6167,N_5818,N_5874);
nand U6168 (N_6168,N_5824,N_5990);
xnor U6169 (N_6169,N_5912,N_5911);
nor U6170 (N_6170,N_5892,N_5931);
or U6171 (N_6171,N_5859,N_5887);
and U6172 (N_6172,N_5841,N_5950);
or U6173 (N_6173,N_5857,N_5951);
or U6174 (N_6174,N_5813,N_5800);
or U6175 (N_6175,N_5841,N_5884);
nor U6176 (N_6176,N_5840,N_5896);
nor U6177 (N_6177,N_5971,N_5819);
or U6178 (N_6178,N_5963,N_5852);
nand U6179 (N_6179,N_5846,N_5847);
and U6180 (N_6180,N_5928,N_5965);
xor U6181 (N_6181,N_5923,N_5818);
or U6182 (N_6182,N_5800,N_5989);
or U6183 (N_6183,N_5923,N_5886);
xor U6184 (N_6184,N_5817,N_5935);
xnor U6185 (N_6185,N_5811,N_5818);
nand U6186 (N_6186,N_5997,N_5809);
nor U6187 (N_6187,N_5805,N_5900);
nor U6188 (N_6188,N_5813,N_5940);
nand U6189 (N_6189,N_5815,N_5924);
xor U6190 (N_6190,N_5914,N_5926);
nor U6191 (N_6191,N_5909,N_5989);
or U6192 (N_6192,N_5864,N_5885);
xnor U6193 (N_6193,N_5986,N_5860);
xnor U6194 (N_6194,N_5995,N_5840);
or U6195 (N_6195,N_5942,N_5945);
and U6196 (N_6196,N_5966,N_5807);
or U6197 (N_6197,N_5949,N_5954);
nand U6198 (N_6198,N_5850,N_5939);
nor U6199 (N_6199,N_5940,N_5965);
or U6200 (N_6200,N_6066,N_6029);
and U6201 (N_6201,N_6039,N_6003);
or U6202 (N_6202,N_6069,N_6158);
and U6203 (N_6203,N_6088,N_6127);
xor U6204 (N_6204,N_6167,N_6084);
or U6205 (N_6205,N_6027,N_6095);
and U6206 (N_6206,N_6010,N_6021);
or U6207 (N_6207,N_6169,N_6179);
xnor U6208 (N_6208,N_6007,N_6079);
and U6209 (N_6209,N_6104,N_6163);
nor U6210 (N_6210,N_6112,N_6156);
and U6211 (N_6211,N_6030,N_6064);
nand U6212 (N_6212,N_6185,N_6159);
and U6213 (N_6213,N_6197,N_6001);
xor U6214 (N_6214,N_6195,N_6181);
xor U6215 (N_6215,N_6130,N_6170);
nor U6216 (N_6216,N_6124,N_6067);
nor U6217 (N_6217,N_6024,N_6113);
and U6218 (N_6218,N_6143,N_6171);
xor U6219 (N_6219,N_6140,N_6086);
or U6220 (N_6220,N_6090,N_6013);
nand U6221 (N_6221,N_6048,N_6191);
nor U6222 (N_6222,N_6133,N_6148);
or U6223 (N_6223,N_6154,N_6015);
nand U6224 (N_6224,N_6198,N_6135);
xnor U6225 (N_6225,N_6085,N_6151);
or U6226 (N_6226,N_6103,N_6105);
xnor U6227 (N_6227,N_6060,N_6132);
and U6228 (N_6228,N_6116,N_6111);
nand U6229 (N_6229,N_6155,N_6180);
nand U6230 (N_6230,N_6096,N_6117);
nor U6231 (N_6231,N_6054,N_6188);
xor U6232 (N_6232,N_6118,N_6074);
or U6233 (N_6233,N_6026,N_6087);
xnor U6234 (N_6234,N_6068,N_6196);
nor U6235 (N_6235,N_6102,N_6023);
nor U6236 (N_6236,N_6160,N_6098);
or U6237 (N_6237,N_6082,N_6081);
nor U6238 (N_6238,N_6194,N_6152);
xnor U6239 (N_6239,N_6093,N_6063);
nor U6240 (N_6240,N_6031,N_6182);
nor U6241 (N_6241,N_6009,N_6042);
xnor U6242 (N_6242,N_6134,N_6121);
nand U6243 (N_6243,N_6120,N_6002);
nor U6244 (N_6244,N_6149,N_6128);
xnor U6245 (N_6245,N_6162,N_6109);
or U6246 (N_6246,N_6036,N_6080);
and U6247 (N_6247,N_6173,N_6178);
and U6248 (N_6248,N_6164,N_6035);
nor U6249 (N_6249,N_6065,N_6061);
nand U6250 (N_6250,N_6083,N_6052);
nand U6251 (N_6251,N_6004,N_6174);
nand U6252 (N_6252,N_6183,N_6106);
and U6253 (N_6253,N_6005,N_6025);
and U6254 (N_6254,N_6016,N_6175);
and U6255 (N_6255,N_6168,N_6014);
or U6256 (N_6256,N_6020,N_6076);
nor U6257 (N_6257,N_6037,N_6141);
or U6258 (N_6258,N_6059,N_6049);
or U6259 (N_6259,N_6041,N_6097);
and U6260 (N_6260,N_6053,N_6012);
xor U6261 (N_6261,N_6000,N_6100);
or U6262 (N_6262,N_6040,N_6126);
and U6263 (N_6263,N_6033,N_6142);
and U6264 (N_6264,N_6115,N_6186);
or U6265 (N_6265,N_6139,N_6008);
xnor U6266 (N_6266,N_6073,N_6187);
xnor U6267 (N_6267,N_6125,N_6047);
xor U6268 (N_6268,N_6107,N_6190);
and U6269 (N_6269,N_6032,N_6192);
nor U6270 (N_6270,N_6157,N_6137);
xnor U6271 (N_6271,N_6094,N_6122);
nor U6272 (N_6272,N_6028,N_6058);
nor U6273 (N_6273,N_6044,N_6193);
nor U6274 (N_6274,N_6017,N_6131);
xnor U6275 (N_6275,N_6199,N_6123);
nor U6276 (N_6276,N_6108,N_6119);
xnor U6277 (N_6277,N_6144,N_6043);
nor U6278 (N_6278,N_6045,N_6150);
or U6279 (N_6279,N_6172,N_6091);
and U6280 (N_6280,N_6146,N_6184);
nor U6281 (N_6281,N_6055,N_6056);
and U6282 (N_6282,N_6099,N_6011);
nand U6283 (N_6283,N_6071,N_6189);
or U6284 (N_6284,N_6075,N_6147);
nand U6285 (N_6285,N_6176,N_6018);
xor U6286 (N_6286,N_6161,N_6019);
nor U6287 (N_6287,N_6166,N_6129);
or U6288 (N_6288,N_6110,N_6092);
or U6289 (N_6289,N_6057,N_6138);
or U6290 (N_6290,N_6136,N_6078);
nand U6291 (N_6291,N_6072,N_6051);
or U6292 (N_6292,N_6114,N_6077);
or U6293 (N_6293,N_6101,N_6145);
nor U6294 (N_6294,N_6022,N_6006);
xnor U6295 (N_6295,N_6034,N_6089);
and U6296 (N_6296,N_6177,N_6050);
or U6297 (N_6297,N_6038,N_6165);
or U6298 (N_6298,N_6046,N_6153);
nand U6299 (N_6299,N_6062,N_6070);
or U6300 (N_6300,N_6024,N_6197);
nor U6301 (N_6301,N_6062,N_6133);
and U6302 (N_6302,N_6034,N_6007);
nor U6303 (N_6303,N_6194,N_6098);
and U6304 (N_6304,N_6168,N_6120);
nor U6305 (N_6305,N_6070,N_6125);
or U6306 (N_6306,N_6103,N_6110);
nor U6307 (N_6307,N_6179,N_6079);
xnor U6308 (N_6308,N_6111,N_6035);
nor U6309 (N_6309,N_6174,N_6126);
or U6310 (N_6310,N_6130,N_6167);
nand U6311 (N_6311,N_6130,N_6094);
and U6312 (N_6312,N_6108,N_6121);
nand U6313 (N_6313,N_6123,N_6137);
or U6314 (N_6314,N_6026,N_6124);
and U6315 (N_6315,N_6016,N_6104);
or U6316 (N_6316,N_6013,N_6196);
xnor U6317 (N_6317,N_6085,N_6140);
and U6318 (N_6318,N_6115,N_6015);
or U6319 (N_6319,N_6185,N_6129);
nor U6320 (N_6320,N_6053,N_6026);
and U6321 (N_6321,N_6105,N_6021);
and U6322 (N_6322,N_6138,N_6072);
nor U6323 (N_6323,N_6037,N_6050);
nor U6324 (N_6324,N_6091,N_6140);
xnor U6325 (N_6325,N_6148,N_6012);
xnor U6326 (N_6326,N_6112,N_6196);
and U6327 (N_6327,N_6192,N_6147);
xnor U6328 (N_6328,N_6103,N_6087);
nand U6329 (N_6329,N_6143,N_6147);
and U6330 (N_6330,N_6102,N_6195);
nor U6331 (N_6331,N_6059,N_6105);
and U6332 (N_6332,N_6108,N_6131);
nand U6333 (N_6333,N_6040,N_6065);
nor U6334 (N_6334,N_6061,N_6125);
nor U6335 (N_6335,N_6177,N_6190);
and U6336 (N_6336,N_6066,N_6061);
xnor U6337 (N_6337,N_6032,N_6072);
nor U6338 (N_6338,N_6012,N_6122);
or U6339 (N_6339,N_6012,N_6074);
xor U6340 (N_6340,N_6064,N_6023);
nand U6341 (N_6341,N_6146,N_6017);
nor U6342 (N_6342,N_6020,N_6050);
xnor U6343 (N_6343,N_6003,N_6019);
nor U6344 (N_6344,N_6074,N_6169);
xor U6345 (N_6345,N_6164,N_6147);
or U6346 (N_6346,N_6157,N_6073);
and U6347 (N_6347,N_6157,N_6024);
or U6348 (N_6348,N_6033,N_6135);
nand U6349 (N_6349,N_6028,N_6005);
nor U6350 (N_6350,N_6167,N_6045);
and U6351 (N_6351,N_6065,N_6063);
xor U6352 (N_6352,N_6032,N_6074);
nor U6353 (N_6353,N_6154,N_6031);
nand U6354 (N_6354,N_6036,N_6070);
or U6355 (N_6355,N_6199,N_6105);
xor U6356 (N_6356,N_6056,N_6001);
and U6357 (N_6357,N_6160,N_6179);
xor U6358 (N_6358,N_6123,N_6190);
nand U6359 (N_6359,N_6047,N_6086);
nand U6360 (N_6360,N_6116,N_6166);
and U6361 (N_6361,N_6123,N_6023);
nor U6362 (N_6362,N_6012,N_6123);
xor U6363 (N_6363,N_6049,N_6056);
and U6364 (N_6364,N_6119,N_6027);
and U6365 (N_6365,N_6155,N_6003);
xor U6366 (N_6366,N_6054,N_6049);
and U6367 (N_6367,N_6090,N_6034);
xor U6368 (N_6368,N_6111,N_6090);
nand U6369 (N_6369,N_6098,N_6148);
nand U6370 (N_6370,N_6139,N_6134);
or U6371 (N_6371,N_6095,N_6017);
or U6372 (N_6372,N_6132,N_6120);
xnor U6373 (N_6373,N_6161,N_6097);
or U6374 (N_6374,N_6114,N_6014);
xnor U6375 (N_6375,N_6144,N_6120);
or U6376 (N_6376,N_6163,N_6142);
xnor U6377 (N_6377,N_6121,N_6011);
xor U6378 (N_6378,N_6180,N_6130);
nor U6379 (N_6379,N_6046,N_6132);
xor U6380 (N_6380,N_6072,N_6083);
and U6381 (N_6381,N_6015,N_6133);
and U6382 (N_6382,N_6073,N_6076);
or U6383 (N_6383,N_6057,N_6047);
and U6384 (N_6384,N_6043,N_6167);
or U6385 (N_6385,N_6187,N_6007);
and U6386 (N_6386,N_6184,N_6190);
nor U6387 (N_6387,N_6075,N_6172);
nand U6388 (N_6388,N_6157,N_6183);
or U6389 (N_6389,N_6079,N_6093);
nor U6390 (N_6390,N_6026,N_6031);
nor U6391 (N_6391,N_6135,N_6055);
or U6392 (N_6392,N_6187,N_6109);
or U6393 (N_6393,N_6119,N_6186);
nand U6394 (N_6394,N_6080,N_6037);
nand U6395 (N_6395,N_6019,N_6073);
xor U6396 (N_6396,N_6147,N_6065);
nand U6397 (N_6397,N_6054,N_6140);
or U6398 (N_6398,N_6198,N_6014);
or U6399 (N_6399,N_6052,N_6117);
nand U6400 (N_6400,N_6317,N_6311);
nor U6401 (N_6401,N_6372,N_6300);
nand U6402 (N_6402,N_6380,N_6282);
xor U6403 (N_6403,N_6378,N_6221);
or U6404 (N_6404,N_6234,N_6294);
or U6405 (N_6405,N_6379,N_6230);
and U6406 (N_6406,N_6212,N_6329);
and U6407 (N_6407,N_6307,N_6396);
nand U6408 (N_6408,N_6219,N_6354);
and U6409 (N_6409,N_6324,N_6328);
and U6410 (N_6410,N_6269,N_6224);
nand U6411 (N_6411,N_6263,N_6314);
nor U6412 (N_6412,N_6209,N_6323);
xnor U6413 (N_6413,N_6285,N_6281);
nor U6414 (N_6414,N_6290,N_6397);
xnor U6415 (N_6415,N_6249,N_6200);
nand U6416 (N_6416,N_6278,N_6312);
or U6417 (N_6417,N_6303,N_6393);
xor U6418 (N_6418,N_6360,N_6349);
xor U6419 (N_6419,N_6291,N_6231);
xor U6420 (N_6420,N_6277,N_6370);
nand U6421 (N_6421,N_6270,N_6255);
and U6422 (N_6422,N_6335,N_6220);
or U6423 (N_6423,N_6353,N_6222);
and U6424 (N_6424,N_6374,N_6348);
nor U6425 (N_6425,N_6326,N_6299);
nand U6426 (N_6426,N_6254,N_6388);
xnor U6427 (N_6427,N_6321,N_6384);
or U6428 (N_6428,N_6233,N_6286);
nand U6429 (N_6429,N_6252,N_6274);
xor U6430 (N_6430,N_6340,N_6295);
nand U6431 (N_6431,N_6346,N_6386);
nand U6432 (N_6432,N_6331,N_6256);
xor U6433 (N_6433,N_6245,N_6217);
or U6434 (N_6434,N_6330,N_6288);
nand U6435 (N_6435,N_6316,N_6351);
and U6436 (N_6436,N_6333,N_6336);
and U6437 (N_6437,N_6377,N_6342);
nand U6438 (N_6438,N_6392,N_6352);
or U6439 (N_6439,N_6215,N_6273);
nand U6440 (N_6440,N_6344,N_6244);
xnor U6441 (N_6441,N_6306,N_6240);
or U6442 (N_6442,N_6271,N_6243);
and U6443 (N_6443,N_6319,N_6225);
or U6444 (N_6444,N_6398,N_6226);
and U6445 (N_6445,N_6210,N_6339);
nand U6446 (N_6446,N_6357,N_6361);
nand U6447 (N_6447,N_6293,N_6204);
xor U6448 (N_6448,N_6223,N_6366);
and U6449 (N_6449,N_6202,N_6376);
xor U6450 (N_6450,N_6261,N_6262);
and U6451 (N_6451,N_6310,N_6399);
and U6452 (N_6452,N_6362,N_6375);
or U6453 (N_6453,N_6229,N_6216);
or U6454 (N_6454,N_6247,N_6395);
and U6455 (N_6455,N_6325,N_6350);
nor U6456 (N_6456,N_6371,N_6341);
nor U6457 (N_6457,N_6258,N_6365);
nand U6458 (N_6458,N_6283,N_6284);
nand U6459 (N_6459,N_6381,N_6242);
nor U6460 (N_6460,N_6238,N_6236);
nor U6461 (N_6461,N_6309,N_6382);
nand U6462 (N_6462,N_6389,N_6302);
or U6463 (N_6463,N_6265,N_6373);
or U6464 (N_6464,N_6235,N_6264);
and U6465 (N_6465,N_6218,N_6367);
xnor U6466 (N_6466,N_6248,N_6214);
or U6467 (N_6467,N_6227,N_6332);
nand U6468 (N_6468,N_6253,N_6205);
nand U6469 (N_6469,N_6390,N_6207);
and U6470 (N_6470,N_6298,N_6266);
nand U6471 (N_6471,N_6322,N_6211);
and U6472 (N_6472,N_6237,N_6347);
nor U6473 (N_6473,N_6267,N_6208);
nor U6474 (N_6474,N_6313,N_6391);
xnor U6475 (N_6475,N_6272,N_6287);
nor U6476 (N_6476,N_6368,N_6305);
xor U6477 (N_6477,N_6275,N_6345);
xnor U6478 (N_6478,N_6383,N_6296);
and U6479 (N_6479,N_6304,N_6358);
or U6480 (N_6480,N_6292,N_6280);
xnor U6481 (N_6481,N_6297,N_6246);
or U6482 (N_6482,N_6276,N_6363);
and U6483 (N_6483,N_6334,N_6369);
nor U6484 (N_6484,N_6228,N_6260);
or U6485 (N_6485,N_6232,N_6318);
or U6486 (N_6486,N_6327,N_6355);
xnor U6487 (N_6487,N_6203,N_6343);
nor U6488 (N_6488,N_6289,N_6250);
and U6489 (N_6489,N_6337,N_6279);
or U6490 (N_6490,N_6364,N_6356);
and U6491 (N_6491,N_6257,N_6251);
or U6492 (N_6492,N_6206,N_6241);
nor U6493 (N_6493,N_6308,N_6301);
and U6494 (N_6494,N_6213,N_6394);
and U6495 (N_6495,N_6201,N_6320);
nor U6496 (N_6496,N_6239,N_6315);
nor U6497 (N_6497,N_6338,N_6387);
xor U6498 (N_6498,N_6268,N_6385);
nor U6499 (N_6499,N_6359,N_6259);
xor U6500 (N_6500,N_6267,N_6247);
and U6501 (N_6501,N_6249,N_6240);
xor U6502 (N_6502,N_6291,N_6309);
and U6503 (N_6503,N_6387,N_6256);
nor U6504 (N_6504,N_6322,N_6386);
xor U6505 (N_6505,N_6220,N_6293);
nor U6506 (N_6506,N_6262,N_6311);
nand U6507 (N_6507,N_6209,N_6321);
xnor U6508 (N_6508,N_6205,N_6296);
or U6509 (N_6509,N_6275,N_6360);
or U6510 (N_6510,N_6358,N_6251);
or U6511 (N_6511,N_6263,N_6320);
and U6512 (N_6512,N_6319,N_6221);
and U6513 (N_6513,N_6385,N_6390);
or U6514 (N_6514,N_6204,N_6322);
and U6515 (N_6515,N_6347,N_6208);
and U6516 (N_6516,N_6322,N_6238);
and U6517 (N_6517,N_6337,N_6275);
nand U6518 (N_6518,N_6303,N_6360);
and U6519 (N_6519,N_6319,N_6282);
and U6520 (N_6520,N_6294,N_6356);
nor U6521 (N_6521,N_6317,N_6210);
xnor U6522 (N_6522,N_6292,N_6226);
nor U6523 (N_6523,N_6396,N_6384);
and U6524 (N_6524,N_6234,N_6302);
nand U6525 (N_6525,N_6340,N_6309);
nor U6526 (N_6526,N_6272,N_6232);
xor U6527 (N_6527,N_6281,N_6298);
or U6528 (N_6528,N_6375,N_6226);
or U6529 (N_6529,N_6230,N_6361);
nor U6530 (N_6530,N_6232,N_6239);
or U6531 (N_6531,N_6221,N_6326);
xnor U6532 (N_6532,N_6364,N_6240);
xnor U6533 (N_6533,N_6248,N_6247);
nand U6534 (N_6534,N_6288,N_6237);
or U6535 (N_6535,N_6361,N_6206);
or U6536 (N_6536,N_6224,N_6228);
nand U6537 (N_6537,N_6344,N_6216);
or U6538 (N_6538,N_6341,N_6271);
nor U6539 (N_6539,N_6237,N_6322);
xor U6540 (N_6540,N_6236,N_6241);
nor U6541 (N_6541,N_6311,N_6357);
nand U6542 (N_6542,N_6312,N_6233);
xor U6543 (N_6543,N_6266,N_6226);
nor U6544 (N_6544,N_6291,N_6391);
xor U6545 (N_6545,N_6220,N_6303);
or U6546 (N_6546,N_6363,N_6244);
nand U6547 (N_6547,N_6268,N_6289);
nand U6548 (N_6548,N_6209,N_6294);
or U6549 (N_6549,N_6357,N_6258);
xnor U6550 (N_6550,N_6399,N_6216);
nand U6551 (N_6551,N_6245,N_6262);
xnor U6552 (N_6552,N_6253,N_6310);
and U6553 (N_6553,N_6205,N_6254);
nand U6554 (N_6554,N_6266,N_6224);
xnor U6555 (N_6555,N_6277,N_6216);
xnor U6556 (N_6556,N_6398,N_6276);
or U6557 (N_6557,N_6333,N_6351);
or U6558 (N_6558,N_6360,N_6387);
xnor U6559 (N_6559,N_6394,N_6240);
and U6560 (N_6560,N_6326,N_6333);
and U6561 (N_6561,N_6363,N_6335);
nor U6562 (N_6562,N_6279,N_6238);
and U6563 (N_6563,N_6327,N_6220);
nor U6564 (N_6564,N_6223,N_6319);
nand U6565 (N_6565,N_6331,N_6212);
nor U6566 (N_6566,N_6396,N_6330);
and U6567 (N_6567,N_6334,N_6370);
and U6568 (N_6568,N_6396,N_6232);
nor U6569 (N_6569,N_6364,N_6282);
or U6570 (N_6570,N_6325,N_6268);
or U6571 (N_6571,N_6207,N_6384);
and U6572 (N_6572,N_6377,N_6310);
xnor U6573 (N_6573,N_6394,N_6343);
xor U6574 (N_6574,N_6280,N_6241);
or U6575 (N_6575,N_6241,N_6268);
nand U6576 (N_6576,N_6273,N_6297);
nand U6577 (N_6577,N_6319,N_6331);
xnor U6578 (N_6578,N_6265,N_6288);
xor U6579 (N_6579,N_6230,N_6307);
xor U6580 (N_6580,N_6233,N_6394);
and U6581 (N_6581,N_6380,N_6254);
nor U6582 (N_6582,N_6264,N_6383);
and U6583 (N_6583,N_6228,N_6345);
xnor U6584 (N_6584,N_6391,N_6344);
and U6585 (N_6585,N_6298,N_6333);
nor U6586 (N_6586,N_6219,N_6292);
nor U6587 (N_6587,N_6226,N_6252);
nor U6588 (N_6588,N_6314,N_6257);
nor U6589 (N_6589,N_6299,N_6335);
nor U6590 (N_6590,N_6309,N_6259);
or U6591 (N_6591,N_6251,N_6313);
xor U6592 (N_6592,N_6280,N_6348);
and U6593 (N_6593,N_6294,N_6371);
or U6594 (N_6594,N_6311,N_6221);
xor U6595 (N_6595,N_6279,N_6208);
xor U6596 (N_6596,N_6317,N_6303);
xor U6597 (N_6597,N_6215,N_6224);
or U6598 (N_6598,N_6303,N_6206);
nor U6599 (N_6599,N_6336,N_6383);
nor U6600 (N_6600,N_6529,N_6407);
nor U6601 (N_6601,N_6446,N_6582);
or U6602 (N_6602,N_6413,N_6577);
xor U6603 (N_6603,N_6593,N_6537);
nor U6604 (N_6604,N_6498,N_6426);
or U6605 (N_6605,N_6434,N_6559);
xnor U6606 (N_6606,N_6497,N_6552);
nand U6607 (N_6607,N_6538,N_6596);
nor U6608 (N_6608,N_6465,N_6578);
nor U6609 (N_6609,N_6534,N_6439);
xor U6610 (N_6610,N_6425,N_6525);
xnor U6611 (N_6611,N_6589,N_6503);
nor U6612 (N_6612,N_6493,N_6496);
nand U6613 (N_6613,N_6443,N_6526);
or U6614 (N_6614,N_6449,N_6447);
or U6615 (N_6615,N_6572,N_6504);
or U6616 (N_6616,N_6513,N_6468);
nand U6617 (N_6617,N_6528,N_6516);
nor U6618 (N_6618,N_6542,N_6597);
xnor U6619 (N_6619,N_6495,N_6514);
nor U6620 (N_6620,N_6583,N_6401);
nor U6621 (N_6621,N_6576,N_6424);
nor U6622 (N_6622,N_6400,N_6402);
or U6623 (N_6623,N_6432,N_6518);
or U6624 (N_6624,N_6460,N_6414);
nand U6625 (N_6625,N_6440,N_6483);
nand U6626 (N_6626,N_6508,N_6558);
nand U6627 (N_6627,N_6475,N_6410);
nor U6628 (N_6628,N_6455,N_6520);
or U6629 (N_6629,N_6442,N_6416);
or U6630 (N_6630,N_6458,N_6462);
and U6631 (N_6631,N_6501,N_6545);
nor U6632 (N_6632,N_6584,N_6421);
nor U6633 (N_6633,N_6482,N_6566);
and U6634 (N_6634,N_6444,N_6574);
or U6635 (N_6635,N_6419,N_6562);
xor U6636 (N_6636,N_6420,N_6565);
and U6637 (N_6637,N_6499,N_6480);
nand U6638 (N_6638,N_6463,N_6488);
nand U6639 (N_6639,N_6408,N_6599);
xnor U6640 (N_6640,N_6456,N_6473);
and U6641 (N_6641,N_6532,N_6595);
nand U6642 (N_6642,N_6587,N_6489);
and U6643 (N_6643,N_6411,N_6594);
and U6644 (N_6644,N_6575,N_6521);
xor U6645 (N_6645,N_6494,N_6539);
and U6646 (N_6646,N_6484,N_6487);
and U6647 (N_6647,N_6569,N_6452);
xnor U6648 (N_6648,N_6471,N_6469);
and U6649 (N_6649,N_6560,N_6580);
xnor U6650 (N_6650,N_6568,N_6547);
nand U6651 (N_6651,N_6409,N_6564);
or U6652 (N_6652,N_6586,N_6453);
or U6653 (N_6653,N_6567,N_6527);
or U6654 (N_6654,N_6429,N_6403);
xor U6655 (N_6655,N_6570,N_6445);
xnor U6656 (N_6656,N_6588,N_6512);
and U6657 (N_6657,N_6437,N_6492);
or U6658 (N_6658,N_6451,N_6491);
nor U6659 (N_6659,N_6517,N_6590);
xor U6660 (N_6660,N_6585,N_6427);
xor U6661 (N_6661,N_6511,N_6418);
xor U6662 (N_6662,N_6459,N_6486);
xor U6663 (N_6663,N_6598,N_6592);
xnor U6664 (N_6664,N_6441,N_6554);
and U6665 (N_6665,N_6573,N_6428);
nor U6666 (N_6666,N_6553,N_6404);
nor U6667 (N_6667,N_6506,N_6531);
or U6668 (N_6668,N_6519,N_6423);
xnor U6669 (N_6669,N_6454,N_6523);
or U6670 (N_6670,N_6481,N_6544);
or U6671 (N_6671,N_6417,N_6561);
nand U6672 (N_6672,N_6579,N_6464);
or U6673 (N_6673,N_6546,N_6466);
nand U6674 (N_6674,N_6479,N_6550);
xor U6675 (N_6675,N_6581,N_6556);
xor U6676 (N_6676,N_6540,N_6448);
xnor U6677 (N_6677,N_6461,N_6438);
and U6678 (N_6678,N_6549,N_6507);
or U6679 (N_6679,N_6415,N_6551);
nor U6680 (N_6680,N_6485,N_6535);
nand U6681 (N_6681,N_6490,N_6530);
nand U6682 (N_6682,N_6470,N_6515);
xnor U6683 (N_6683,N_6467,N_6541);
or U6684 (N_6684,N_6431,N_6543);
nand U6685 (N_6685,N_6412,N_6548);
xor U6686 (N_6686,N_6500,N_6436);
xor U6687 (N_6687,N_6555,N_6422);
nor U6688 (N_6688,N_6563,N_6533);
nand U6689 (N_6689,N_6591,N_6557);
xor U6690 (N_6690,N_6474,N_6524);
nor U6691 (N_6691,N_6536,N_6477);
and U6692 (N_6692,N_6406,N_6433);
and U6693 (N_6693,N_6430,N_6476);
xnor U6694 (N_6694,N_6502,N_6522);
xnor U6695 (N_6695,N_6510,N_6478);
and U6696 (N_6696,N_6472,N_6457);
and U6697 (N_6697,N_6571,N_6405);
and U6698 (N_6698,N_6435,N_6509);
nor U6699 (N_6699,N_6505,N_6450);
and U6700 (N_6700,N_6567,N_6560);
or U6701 (N_6701,N_6487,N_6545);
and U6702 (N_6702,N_6413,N_6510);
xor U6703 (N_6703,N_6483,N_6500);
or U6704 (N_6704,N_6599,N_6412);
nor U6705 (N_6705,N_6406,N_6576);
xor U6706 (N_6706,N_6485,N_6468);
xor U6707 (N_6707,N_6576,N_6542);
or U6708 (N_6708,N_6433,N_6520);
nand U6709 (N_6709,N_6472,N_6433);
or U6710 (N_6710,N_6407,N_6518);
xnor U6711 (N_6711,N_6445,N_6509);
xor U6712 (N_6712,N_6432,N_6585);
xnor U6713 (N_6713,N_6561,N_6501);
nor U6714 (N_6714,N_6547,N_6525);
xor U6715 (N_6715,N_6445,N_6549);
or U6716 (N_6716,N_6417,N_6434);
or U6717 (N_6717,N_6503,N_6595);
nand U6718 (N_6718,N_6594,N_6537);
xnor U6719 (N_6719,N_6591,N_6587);
nand U6720 (N_6720,N_6565,N_6553);
nand U6721 (N_6721,N_6443,N_6573);
nand U6722 (N_6722,N_6411,N_6567);
nor U6723 (N_6723,N_6485,N_6472);
nor U6724 (N_6724,N_6509,N_6441);
and U6725 (N_6725,N_6401,N_6451);
or U6726 (N_6726,N_6480,N_6550);
and U6727 (N_6727,N_6498,N_6468);
xnor U6728 (N_6728,N_6509,N_6583);
xor U6729 (N_6729,N_6455,N_6593);
or U6730 (N_6730,N_6420,N_6563);
and U6731 (N_6731,N_6585,N_6496);
nor U6732 (N_6732,N_6457,N_6475);
or U6733 (N_6733,N_6444,N_6492);
nor U6734 (N_6734,N_6424,N_6559);
or U6735 (N_6735,N_6443,N_6416);
or U6736 (N_6736,N_6528,N_6434);
nor U6737 (N_6737,N_6421,N_6429);
nor U6738 (N_6738,N_6542,N_6485);
nand U6739 (N_6739,N_6565,N_6430);
nand U6740 (N_6740,N_6426,N_6473);
and U6741 (N_6741,N_6476,N_6537);
or U6742 (N_6742,N_6599,N_6529);
nor U6743 (N_6743,N_6562,N_6446);
or U6744 (N_6744,N_6548,N_6552);
or U6745 (N_6745,N_6569,N_6511);
or U6746 (N_6746,N_6437,N_6513);
nand U6747 (N_6747,N_6491,N_6512);
xnor U6748 (N_6748,N_6500,N_6481);
xor U6749 (N_6749,N_6489,N_6410);
nand U6750 (N_6750,N_6436,N_6433);
and U6751 (N_6751,N_6453,N_6565);
xor U6752 (N_6752,N_6535,N_6589);
nor U6753 (N_6753,N_6485,N_6562);
and U6754 (N_6754,N_6456,N_6454);
nand U6755 (N_6755,N_6573,N_6412);
and U6756 (N_6756,N_6442,N_6407);
nand U6757 (N_6757,N_6439,N_6438);
nand U6758 (N_6758,N_6455,N_6546);
nand U6759 (N_6759,N_6549,N_6438);
nor U6760 (N_6760,N_6518,N_6586);
or U6761 (N_6761,N_6485,N_6511);
and U6762 (N_6762,N_6587,N_6564);
and U6763 (N_6763,N_6423,N_6547);
or U6764 (N_6764,N_6511,N_6430);
and U6765 (N_6765,N_6509,N_6528);
and U6766 (N_6766,N_6510,N_6425);
and U6767 (N_6767,N_6413,N_6555);
or U6768 (N_6768,N_6509,N_6450);
and U6769 (N_6769,N_6489,N_6566);
or U6770 (N_6770,N_6549,N_6471);
nor U6771 (N_6771,N_6447,N_6520);
nor U6772 (N_6772,N_6560,N_6464);
nor U6773 (N_6773,N_6546,N_6419);
nand U6774 (N_6774,N_6474,N_6405);
nor U6775 (N_6775,N_6458,N_6407);
or U6776 (N_6776,N_6559,N_6459);
xnor U6777 (N_6777,N_6481,N_6574);
nand U6778 (N_6778,N_6583,N_6486);
or U6779 (N_6779,N_6401,N_6478);
nor U6780 (N_6780,N_6464,N_6598);
nor U6781 (N_6781,N_6438,N_6410);
xnor U6782 (N_6782,N_6407,N_6448);
nand U6783 (N_6783,N_6479,N_6504);
and U6784 (N_6784,N_6576,N_6428);
and U6785 (N_6785,N_6445,N_6516);
or U6786 (N_6786,N_6577,N_6415);
xnor U6787 (N_6787,N_6581,N_6584);
nand U6788 (N_6788,N_6426,N_6587);
nor U6789 (N_6789,N_6434,N_6526);
nand U6790 (N_6790,N_6457,N_6596);
and U6791 (N_6791,N_6438,N_6525);
nor U6792 (N_6792,N_6427,N_6431);
or U6793 (N_6793,N_6514,N_6484);
nor U6794 (N_6794,N_6521,N_6415);
nor U6795 (N_6795,N_6555,N_6439);
and U6796 (N_6796,N_6495,N_6571);
xnor U6797 (N_6797,N_6502,N_6474);
or U6798 (N_6798,N_6456,N_6417);
nor U6799 (N_6799,N_6483,N_6572);
nor U6800 (N_6800,N_6616,N_6726);
nor U6801 (N_6801,N_6716,N_6650);
or U6802 (N_6802,N_6659,N_6733);
nor U6803 (N_6803,N_6731,N_6643);
xnor U6804 (N_6804,N_6718,N_6607);
and U6805 (N_6805,N_6720,N_6705);
nor U6806 (N_6806,N_6682,N_6656);
nor U6807 (N_6807,N_6722,N_6639);
xnor U6808 (N_6808,N_6793,N_6688);
and U6809 (N_6809,N_6623,N_6763);
or U6810 (N_6810,N_6781,N_6737);
xnor U6811 (N_6811,N_6640,N_6608);
xor U6812 (N_6812,N_6613,N_6695);
nor U6813 (N_6813,N_6666,N_6744);
and U6814 (N_6814,N_6645,N_6615);
nor U6815 (N_6815,N_6753,N_6784);
and U6816 (N_6816,N_6642,N_6738);
nand U6817 (N_6817,N_6755,N_6617);
or U6818 (N_6818,N_6783,N_6610);
nor U6819 (N_6819,N_6729,N_6631);
xnor U6820 (N_6820,N_6684,N_6609);
nand U6821 (N_6821,N_6652,N_6669);
or U6822 (N_6822,N_6795,N_6751);
xor U6823 (N_6823,N_6750,N_6638);
nor U6824 (N_6824,N_6633,N_6727);
xor U6825 (N_6825,N_6646,N_6620);
and U6826 (N_6826,N_6647,N_6797);
nand U6827 (N_6827,N_6754,N_6628);
or U6828 (N_6828,N_6779,N_6776);
or U6829 (N_6829,N_6758,N_6612);
and U6830 (N_6830,N_6704,N_6703);
or U6831 (N_6831,N_6680,N_6713);
and U6832 (N_6832,N_6799,N_6601);
and U6833 (N_6833,N_6604,N_6674);
and U6834 (N_6834,N_6707,N_6760);
nand U6835 (N_6835,N_6685,N_6603);
xor U6836 (N_6836,N_6723,N_6619);
xnor U6837 (N_6837,N_6699,N_6681);
nand U6838 (N_6838,N_6759,N_6622);
nand U6839 (N_6839,N_6766,N_6796);
nor U6840 (N_6840,N_6698,N_6664);
or U6841 (N_6841,N_6696,N_6630);
nand U6842 (N_6842,N_6732,N_6748);
and U6843 (N_6843,N_6730,N_6677);
or U6844 (N_6844,N_6670,N_6756);
nor U6845 (N_6845,N_6606,N_6773);
or U6846 (N_6846,N_6658,N_6675);
xnor U6847 (N_6847,N_6693,N_6767);
xor U6848 (N_6848,N_6626,N_6770);
and U6849 (N_6849,N_6788,N_6661);
and U6850 (N_6850,N_6761,N_6752);
nand U6851 (N_6851,N_6701,N_6663);
and U6852 (N_6852,N_6777,N_6746);
and U6853 (N_6853,N_6690,N_6605);
nand U6854 (N_6854,N_6787,N_6708);
xor U6855 (N_6855,N_6602,N_6673);
nand U6856 (N_6856,N_6764,N_6769);
xnor U6857 (N_6857,N_6653,N_6790);
nor U6858 (N_6858,N_6778,N_6772);
xnor U6859 (N_6859,N_6665,N_6749);
nor U6860 (N_6860,N_6710,N_6785);
or U6861 (N_6861,N_6637,N_6600);
or U6862 (N_6862,N_6644,N_6735);
nor U6863 (N_6863,N_6686,N_6614);
or U6864 (N_6864,N_6721,N_6629);
xnor U6865 (N_6865,N_6714,N_6678);
nand U6866 (N_6866,N_6741,N_6780);
nor U6867 (N_6867,N_6798,N_6743);
and U6868 (N_6868,N_6657,N_6655);
xor U6869 (N_6869,N_6757,N_6789);
and U6870 (N_6870,N_6660,N_6611);
nand U6871 (N_6871,N_6728,N_6689);
or U6872 (N_6872,N_6774,N_6668);
nor U6873 (N_6873,N_6676,N_6786);
and U6874 (N_6874,N_6687,N_6672);
nor U6875 (N_6875,N_6691,N_6671);
or U6876 (N_6876,N_6634,N_6649);
or U6877 (N_6877,N_6621,N_6702);
nor U6878 (N_6878,N_6791,N_6742);
xnor U6879 (N_6879,N_6662,N_6794);
nand U6880 (N_6880,N_6782,N_6768);
xor U6881 (N_6881,N_6709,N_6697);
and U6882 (N_6882,N_6627,N_6719);
nor U6883 (N_6883,N_6694,N_6736);
xnor U6884 (N_6884,N_6775,N_6711);
nand U6885 (N_6885,N_6717,N_6654);
xor U6886 (N_6886,N_6651,N_6618);
nor U6887 (N_6887,N_6667,N_6679);
and U6888 (N_6888,N_6648,N_6724);
nor U6889 (N_6889,N_6739,N_6771);
nand U6890 (N_6890,N_6625,N_6745);
and U6891 (N_6891,N_6762,N_6692);
nor U6892 (N_6892,N_6792,N_6636);
nor U6893 (N_6893,N_6706,N_6740);
xnor U6894 (N_6894,N_6715,N_6635);
xor U6895 (N_6895,N_6734,N_6747);
nand U6896 (N_6896,N_6765,N_6683);
or U6897 (N_6897,N_6641,N_6725);
xor U6898 (N_6898,N_6632,N_6624);
xor U6899 (N_6899,N_6700,N_6712);
nand U6900 (N_6900,N_6789,N_6675);
nor U6901 (N_6901,N_6781,N_6742);
xor U6902 (N_6902,N_6712,N_6691);
nor U6903 (N_6903,N_6634,N_6704);
xnor U6904 (N_6904,N_6710,N_6644);
nor U6905 (N_6905,N_6690,N_6726);
and U6906 (N_6906,N_6738,N_6704);
xor U6907 (N_6907,N_6617,N_6669);
and U6908 (N_6908,N_6608,N_6613);
nor U6909 (N_6909,N_6719,N_6704);
nand U6910 (N_6910,N_6659,N_6790);
or U6911 (N_6911,N_6602,N_6706);
nand U6912 (N_6912,N_6633,N_6622);
xnor U6913 (N_6913,N_6709,N_6606);
xnor U6914 (N_6914,N_6651,N_6641);
xnor U6915 (N_6915,N_6636,N_6793);
nor U6916 (N_6916,N_6748,N_6602);
nand U6917 (N_6917,N_6741,N_6691);
and U6918 (N_6918,N_6637,N_6709);
nor U6919 (N_6919,N_6698,N_6616);
and U6920 (N_6920,N_6703,N_6600);
nor U6921 (N_6921,N_6750,N_6683);
or U6922 (N_6922,N_6659,N_6666);
or U6923 (N_6923,N_6737,N_6798);
xnor U6924 (N_6924,N_6656,N_6705);
xnor U6925 (N_6925,N_6676,N_6730);
nand U6926 (N_6926,N_6695,N_6737);
and U6927 (N_6927,N_6658,N_6624);
or U6928 (N_6928,N_6785,N_6694);
and U6929 (N_6929,N_6712,N_6600);
nor U6930 (N_6930,N_6679,N_6687);
and U6931 (N_6931,N_6749,N_6792);
nand U6932 (N_6932,N_6724,N_6758);
nand U6933 (N_6933,N_6622,N_6617);
xor U6934 (N_6934,N_6616,N_6663);
and U6935 (N_6935,N_6632,N_6674);
nor U6936 (N_6936,N_6761,N_6631);
or U6937 (N_6937,N_6740,N_6607);
nand U6938 (N_6938,N_6672,N_6626);
nand U6939 (N_6939,N_6754,N_6693);
or U6940 (N_6940,N_6782,N_6715);
nand U6941 (N_6941,N_6719,N_6640);
or U6942 (N_6942,N_6739,N_6753);
or U6943 (N_6943,N_6718,N_6798);
xor U6944 (N_6944,N_6605,N_6667);
xnor U6945 (N_6945,N_6619,N_6776);
nor U6946 (N_6946,N_6640,N_6704);
and U6947 (N_6947,N_6797,N_6784);
xnor U6948 (N_6948,N_6623,N_6729);
xor U6949 (N_6949,N_6786,N_6627);
xor U6950 (N_6950,N_6678,N_6685);
xor U6951 (N_6951,N_6704,N_6632);
or U6952 (N_6952,N_6644,N_6712);
nand U6953 (N_6953,N_6764,N_6708);
nor U6954 (N_6954,N_6779,N_6632);
and U6955 (N_6955,N_6741,N_6732);
nor U6956 (N_6956,N_6758,N_6702);
and U6957 (N_6957,N_6650,N_6639);
and U6958 (N_6958,N_6687,N_6722);
xnor U6959 (N_6959,N_6612,N_6712);
or U6960 (N_6960,N_6677,N_6719);
or U6961 (N_6961,N_6608,N_6681);
nand U6962 (N_6962,N_6656,N_6607);
nand U6963 (N_6963,N_6685,N_6609);
xor U6964 (N_6964,N_6648,N_6722);
or U6965 (N_6965,N_6695,N_6660);
nor U6966 (N_6966,N_6767,N_6609);
nor U6967 (N_6967,N_6713,N_6645);
and U6968 (N_6968,N_6602,N_6636);
or U6969 (N_6969,N_6739,N_6721);
and U6970 (N_6970,N_6645,N_6723);
and U6971 (N_6971,N_6686,N_6618);
or U6972 (N_6972,N_6716,N_6770);
nor U6973 (N_6973,N_6773,N_6794);
or U6974 (N_6974,N_6624,N_6638);
or U6975 (N_6975,N_6770,N_6764);
or U6976 (N_6976,N_6682,N_6799);
and U6977 (N_6977,N_6749,N_6723);
and U6978 (N_6978,N_6655,N_6650);
and U6979 (N_6979,N_6743,N_6793);
and U6980 (N_6980,N_6778,N_6769);
and U6981 (N_6981,N_6628,N_6635);
nor U6982 (N_6982,N_6790,N_6736);
or U6983 (N_6983,N_6730,N_6673);
xor U6984 (N_6984,N_6766,N_6786);
nand U6985 (N_6985,N_6766,N_6734);
or U6986 (N_6986,N_6690,N_6677);
nor U6987 (N_6987,N_6725,N_6716);
xnor U6988 (N_6988,N_6690,N_6750);
xnor U6989 (N_6989,N_6729,N_6712);
xor U6990 (N_6990,N_6616,N_6624);
nor U6991 (N_6991,N_6672,N_6642);
nand U6992 (N_6992,N_6714,N_6647);
and U6993 (N_6993,N_6627,N_6756);
xor U6994 (N_6994,N_6686,N_6627);
nor U6995 (N_6995,N_6764,N_6739);
nand U6996 (N_6996,N_6785,N_6754);
nand U6997 (N_6997,N_6753,N_6674);
xnor U6998 (N_6998,N_6617,N_6732);
and U6999 (N_6999,N_6790,N_6687);
and U7000 (N_7000,N_6827,N_6873);
or U7001 (N_7001,N_6988,N_6830);
nor U7002 (N_7002,N_6979,N_6839);
nand U7003 (N_7003,N_6820,N_6965);
and U7004 (N_7004,N_6823,N_6958);
or U7005 (N_7005,N_6915,N_6859);
nor U7006 (N_7006,N_6886,N_6906);
nand U7007 (N_7007,N_6897,N_6922);
and U7008 (N_7008,N_6907,N_6815);
and U7009 (N_7009,N_6809,N_6831);
and U7010 (N_7010,N_6882,N_6801);
nor U7011 (N_7011,N_6876,N_6854);
nor U7012 (N_7012,N_6810,N_6819);
nand U7013 (N_7013,N_6804,N_6954);
nand U7014 (N_7014,N_6803,N_6864);
xnor U7015 (N_7015,N_6939,N_6805);
or U7016 (N_7016,N_6899,N_6868);
xnor U7017 (N_7017,N_6981,N_6877);
nand U7018 (N_7018,N_6937,N_6871);
nor U7019 (N_7019,N_6984,N_6977);
xnor U7020 (N_7020,N_6866,N_6829);
or U7021 (N_7021,N_6989,N_6942);
nor U7022 (N_7022,N_6843,N_6933);
or U7023 (N_7023,N_6817,N_6821);
or U7024 (N_7024,N_6930,N_6855);
and U7025 (N_7025,N_6881,N_6961);
nor U7026 (N_7026,N_6980,N_6901);
and U7027 (N_7027,N_6846,N_6992);
and U7028 (N_7028,N_6959,N_6875);
nor U7029 (N_7029,N_6894,N_6966);
nand U7030 (N_7030,N_6806,N_6970);
nor U7031 (N_7031,N_6945,N_6923);
nand U7032 (N_7032,N_6911,N_6816);
nand U7033 (N_7033,N_6925,N_6913);
nand U7034 (N_7034,N_6892,N_6990);
nor U7035 (N_7035,N_6946,N_6828);
xnor U7036 (N_7036,N_6953,N_6996);
nand U7037 (N_7037,N_6808,N_6999);
xnor U7038 (N_7038,N_6818,N_6916);
or U7039 (N_7039,N_6890,N_6902);
xnor U7040 (N_7040,N_6962,N_6924);
nor U7041 (N_7041,N_6834,N_6842);
nor U7042 (N_7042,N_6969,N_6857);
xor U7043 (N_7043,N_6949,N_6893);
nor U7044 (N_7044,N_6837,N_6974);
and U7045 (N_7045,N_6891,N_6975);
nor U7046 (N_7046,N_6870,N_6928);
nand U7047 (N_7047,N_6879,N_6950);
and U7048 (N_7048,N_6904,N_6967);
and U7049 (N_7049,N_6835,N_6921);
and U7050 (N_7050,N_6847,N_6919);
and U7051 (N_7051,N_6968,N_6940);
or U7052 (N_7052,N_6858,N_6938);
nand U7053 (N_7053,N_6912,N_6934);
or U7054 (N_7054,N_6995,N_6936);
and U7055 (N_7055,N_6872,N_6972);
or U7056 (N_7056,N_6991,N_6848);
and U7057 (N_7057,N_6852,N_6814);
nor U7058 (N_7058,N_6844,N_6856);
and U7059 (N_7059,N_6869,N_6983);
or U7060 (N_7060,N_6932,N_6960);
and U7061 (N_7061,N_6955,N_6833);
nor U7062 (N_7062,N_6917,N_6800);
xor U7063 (N_7063,N_6889,N_6998);
nor U7064 (N_7064,N_6822,N_6824);
or U7065 (N_7065,N_6941,N_6865);
xnor U7066 (N_7066,N_6929,N_6909);
nand U7067 (N_7067,N_6903,N_6931);
xnor U7068 (N_7068,N_6825,N_6896);
nand U7069 (N_7069,N_6914,N_6826);
and U7070 (N_7070,N_6811,N_6860);
and U7071 (N_7071,N_6982,N_6867);
nand U7072 (N_7072,N_6943,N_6905);
nand U7073 (N_7073,N_6812,N_6985);
nor U7074 (N_7074,N_6973,N_6807);
nand U7075 (N_7075,N_6987,N_6863);
and U7076 (N_7076,N_6845,N_6997);
nand U7077 (N_7077,N_6976,N_6840);
xnor U7078 (N_7078,N_6963,N_6957);
nor U7079 (N_7079,N_6898,N_6964);
nand U7080 (N_7080,N_6910,N_6885);
and U7081 (N_7081,N_6994,N_6813);
nor U7082 (N_7082,N_6927,N_6861);
xor U7083 (N_7083,N_6956,N_6850);
and U7084 (N_7084,N_6883,N_6895);
nor U7085 (N_7085,N_6947,N_6951);
and U7086 (N_7086,N_6900,N_6948);
xor U7087 (N_7087,N_6853,N_6971);
nand U7088 (N_7088,N_6920,N_6849);
nor U7089 (N_7089,N_6862,N_6851);
and U7090 (N_7090,N_6836,N_6874);
nor U7091 (N_7091,N_6838,N_6888);
xnor U7092 (N_7092,N_6944,N_6841);
nand U7093 (N_7093,N_6952,N_6908);
nand U7094 (N_7094,N_6880,N_6935);
and U7095 (N_7095,N_6986,N_6832);
xnor U7096 (N_7096,N_6993,N_6802);
and U7097 (N_7097,N_6884,N_6926);
or U7098 (N_7098,N_6918,N_6887);
nand U7099 (N_7099,N_6978,N_6878);
or U7100 (N_7100,N_6963,N_6936);
or U7101 (N_7101,N_6905,N_6876);
nand U7102 (N_7102,N_6998,N_6833);
xnor U7103 (N_7103,N_6984,N_6878);
nor U7104 (N_7104,N_6961,N_6885);
nand U7105 (N_7105,N_6901,N_6984);
and U7106 (N_7106,N_6902,N_6819);
or U7107 (N_7107,N_6896,N_6963);
xor U7108 (N_7108,N_6998,N_6849);
or U7109 (N_7109,N_6857,N_6973);
nor U7110 (N_7110,N_6880,N_6923);
or U7111 (N_7111,N_6936,N_6951);
nor U7112 (N_7112,N_6895,N_6826);
and U7113 (N_7113,N_6998,N_6980);
xor U7114 (N_7114,N_6899,N_6946);
and U7115 (N_7115,N_6957,N_6868);
nor U7116 (N_7116,N_6865,N_6807);
nand U7117 (N_7117,N_6850,N_6964);
or U7118 (N_7118,N_6929,N_6830);
and U7119 (N_7119,N_6883,N_6812);
and U7120 (N_7120,N_6946,N_6971);
nand U7121 (N_7121,N_6955,N_6801);
nand U7122 (N_7122,N_6890,N_6894);
or U7123 (N_7123,N_6955,N_6812);
nand U7124 (N_7124,N_6868,N_6998);
xnor U7125 (N_7125,N_6881,N_6840);
nand U7126 (N_7126,N_6843,N_6897);
nor U7127 (N_7127,N_6989,N_6886);
and U7128 (N_7128,N_6814,N_6968);
nand U7129 (N_7129,N_6930,N_6823);
xor U7130 (N_7130,N_6967,N_6919);
or U7131 (N_7131,N_6854,N_6932);
nor U7132 (N_7132,N_6820,N_6933);
or U7133 (N_7133,N_6952,N_6943);
or U7134 (N_7134,N_6961,N_6812);
nor U7135 (N_7135,N_6837,N_6922);
xor U7136 (N_7136,N_6936,N_6992);
nor U7137 (N_7137,N_6857,N_6903);
nand U7138 (N_7138,N_6938,N_6846);
and U7139 (N_7139,N_6864,N_6917);
xnor U7140 (N_7140,N_6896,N_6883);
nor U7141 (N_7141,N_6801,N_6976);
or U7142 (N_7142,N_6870,N_6813);
xor U7143 (N_7143,N_6881,N_6928);
nor U7144 (N_7144,N_6829,N_6978);
and U7145 (N_7145,N_6996,N_6853);
nand U7146 (N_7146,N_6874,N_6824);
or U7147 (N_7147,N_6987,N_6838);
nand U7148 (N_7148,N_6970,N_6930);
nor U7149 (N_7149,N_6939,N_6909);
nor U7150 (N_7150,N_6945,N_6992);
xnor U7151 (N_7151,N_6811,N_6963);
nor U7152 (N_7152,N_6880,N_6882);
xor U7153 (N_7153,N_6806,N_6837);
nand U7154 (N_7154,N_6862,N_6946);
or U7155 (N_7155,N_6936,N_6929);
xnor U7156 (N_7156,N_6859,N_6828);
and U7157 (N_7157,N_6861,N_6909);
nor U7158 (N_7158,N_6952,N_6936);
nor U7159 (N_7159,N_6860,N_6970);
nor U7160 (N_7160,N_6868,N_6893);
and U7161 (N_7161,N_6853,N_6908);
xor U7162 (N_7162,N_6832,N_6858);
and U7163 (N_7163,N_6947,N_6930);
and U7164 (N_7164,N_6897,N_6947);
or U7165 (N_7165,N_6888,N_6822);
or U7166 (N_7166,N_6973,N_6808);
or U7167 (N_7167,N_6959,N_6933);
and U7168 (N_7168,N_6825,N_6868);
or U7169 (N_7169,N_6887,N_6811);
or U7170 (N_7170,N_6953,N_6898);
and U7171 (N_7171,N_6962,N_6953);
xor U7172 (N_7172,N_6935,N_6854);
nand U7173 (N_7173,N_6899,N_6885);
nor U7174 (N_7174,N_6847,N_6839);
or U7175 (N_7175,N_6916,N_6982);
nor U7176 (N_7176,N_6940,N_6900);
and U7177 (N_7177,N_6907,N_6823);
nor U7178 (N_7178,N_6814,N_6969);
and U7179 (N_7179,N_6979,N_6832);
nand U7180 (N_7180,N_6934,N_6922);
xnor U7181 (N_7181,N_6872,N_6909);
nor U7182 (N_7182,N_6973,N_6899);
nor U7183 (N_7183,N_6816,N_6839);
xnor U7184 (N_7184,N_6828,N_6929);
and U7185 (N_7185,N_6904,N_6916);
and U7186 (N_7186,N_6906,N_6947);
xnor U7187 (N_7187,N_6962,N_6939);
xnor U7188 (N_7188,N_6902,N_6929);
or U7189 (N_7189,N_6935,N_6918);
and U7190 (N_7190,N_6803,N_6848);
or U7191 (N_7191,N_6951,N_6997);
nand U7192 (N_7192,N_6938,N_6915);
nor U7193 (N_7193,N_6886,N_6936);
and U7194 (N_7194,N_6956,N_6906);
xnor U7195 (N_7195,N_6876,N_6888);
or U7196 (N_7196,N_6993,N_6944);
and U7197 (N_7197,N_6934,N_6881);
nand U7198 (N_7198,N_6929,N_6968);
xnor U7199 (N_7199,N_6894,N_6816);
nand U7200 (N_7200,N_7013,N_7022);
and U7201 (N_7201,N_7136,N_7119);
or U7202 (N_7202,N_7091,N_7134);
nand U7203 (N_7203,N_7071,N_7129);
nand U7204 (N_7204,N_7076,N_7083);
and U7205 (N_7205,N_7020,N_7146);
nor U7206 (N_7206,N_7050,N_7128);
xnor U7207 (N_7207,N_7199,N_7040);
and U7208 (N_7208,N_7085,N_7008);
xnor U7209 (N_7209,N_7177,N_7080);
and U7210 (N_7210,N_7028,N_7142);
nor U7211 (N_7211,N_7035,N_7193);
nand U7212 (N_7212,N_7024,N_7059);
nand U7213 (N_7213,N_7079,N_7167);
and U7214 (N_7214,N_7141,N_7092);
and U7215 (N_7215,N_7086,N_7118);
nor U7216 (N_7216,N_7150,N_7117);
or U7217 (N_7217,N_7171,N_7123);
nand U7218 (N_7218,N_7164,N_7183);
and U7219 (N_7219,N_7007,N_7056);
or U7220 (N_7220,N_7127,N_7004);
or U7221 (N_7221,N_7166,N_7068);
and U7222 (N_7222,N_7095,N_7126);
nor U7223 (N_7223,N_7009,N_7017);
or U7224 (N_7224,N_7132,N_7006);
and U7225 (N_7225,N_7034,N_7151);
nand U7226 (N_7226,N_7075,N_7180);
nand U7227 (N_7227,N_7100,N_7072);
nand U7228 (N_7228,N_7157,N_7149);
nor U7229 (N_7229,N_7131,N_7098);
nor U7230 (N_7230,N_7053,N_7170);
xor U7231 (N_7231,N_7031,N_7172);
nand U7232 (N_7232,N_7154,N_7087);
nand U7233 (N_7233,N_7067,N_7042);
nor U7234 (N_7234,N_7001,N_7104);
nand U7235 (N_7235,N_7054,N_7137);
or U7236 (N_7236,N_7084,N_7069);
nor U7237 (N_7237,N_7182,N_7143);
or U7238 (N_7238,N_7195,N_7187);
xnor U7239 (N_7239,N_7070,N_7122);
or U7240 (N_7240,N_7046,N_7124);
nor U7241 (N_7241,N_7176,N_7152);
nand U7242 (N_7242,N_7185,N_7181);
xor U7243 (N_7243,N_7094,N_7074);
nand U7244 (N_7244,N_7153,N_7108);
nand U7245 (N_7245,N_7189,N_7144);
or U7246 (N_7246,N_7096,N_7038);
nor U7247 (N_7247,N_7110,N_7043);
and U7248 (N_7248,N_7049,N_7198);
or U7249 (N_7249,N_7058,N_7037);
nor U7250 (N_7250,N_7158,N_7130);
nand U7251 (N_7251,N_7111,N_7140);
xnor U7252 (N_7252,N_7121,N_7194);
xor U7253 (N_7253,N_7093,N_7101);
nor U7254 (N_7254,N_7168,N_7192);
nor U7255 (N_7255,N_7027,N_7191);
nand U7256 (N_7256,N_7016,N_7155);
xor U7257 (N_7257,N_7163,N_7148);
nor U7258 (N_7258,N_7173,N_7135);
and U7259 (N_7259,N_7109,N_7147);
or U7260 (N_7260,N_7179,N_7066);
nand U7261 (N_7261,N_7041,N_7023);
nor U7262 (N_7262,N_7052,N_7064);
or U7263 (N_7263,N_7169,N_7003);
nor U7264 (N_7264,N_7184,N_7051);
and U7265 (N_7265,N_7010,N_7145);
nor U7266 (N_7266,N_7099,N_7114);
nor U7267 (N_7267,N_7188,N_7113);
xor U7268 (N_7268,N_7107,N_7073);
nand U7269 (N_7269,N_7178,N_7062);
or U7270 (N_7270,N_7018,N_7160);
or U7271 (N_7271,N_7026,N_7036);
nand U7272 (N_7272,N_7048,N_7133);
nor U7273 (N_7273,N_7197,N_7138);
xor U7274 (N_7274,N_7000,N_7011);
xnor U7275 (N_7275,N_7047,N_7081);
nor U7276 (N_7276,N_7029,N_7057);
nand U7277 (N_7277,N_7186,N_7021);
xnor U7278 (N_7278,N_7175,N_7015);
xor U7279 (N_7279,N_7078,N_7165);
xor U7280 (N_7280,N_7102,N_7077);
nor U7281 (N_7281,N_7012,N_7044);
and U7282 (N_7282,N_7174,N_7033);
nor U7283 (N_7283,N_7082,N_7019);
and U7284 (N_7284,N_7159,N_7112);
or U7285 (N_7285,N_7030,N_7045);
nand U7286 (N_7286,N_7088,N_7055);
xnor U7287 (N_7287,N_7039,N_7125);
nor U7288 (N_7288,N_7005,N_7032);
xnor U7289 (N_7289,N_7065,N_7061);
or U7290 (N_7290,N_7025,N_7161);
or U7291 (N_7291,N_7105,N_7120);
nor U7292 (N_7292,N_7060,N_7116);
and U7293 (N_7293,N_7090,N_7002);
xnor U7294 (N_7294,N_7115,N_7196);
and U7295 (N_7295,N_7106,N_7014);
xnor U7296 (N_7296,N_7190,N_7103);
and U7297 (N_7297,N_7097,N_7156);
and U7298 (N_7298,N_7139,N_7162);
or U7299 (N_7299,N_7063,N_7089);
xor U7300 (N_7300,N_7004,N_7149);
or U7301 (N_7301,N_7188,N_7131);
nor U7302 (N_7302,N_7119,N_7105);
nor U7303 (N_7303,N_7170,N_7028);
xor U7304 (N_7304,N_7109,N_7054);
nand U7305 (N_7305,N_7195,N_7026);
xor U7306 (N_7306,N_7041,N_7112);
nor U7307 (N_7307,N_7159,N_7096);
nor U7308 (N_7308,N_7172,N_7077);
or U7309 (N_7309,N_7133,N_7180);
xnor U7310 (N_7310,N_7116,N_7143);
nor U7311 (N_7311,N_7095,N_7146);
nand U7312 (N_7312,N_7080,N_7139);
and U7313 (N_7313,N_7116,N_7179);
nand U7314 (N_7314,N_7190,N_7006);
xnor U7315 (N_7315,N_7000,N_7004);
xor U7316 (N_7316,N_7052,N_7031);
nor U7317 (N_7317,N_7192,N_7060);
xnor U7318 (N_7318,N_7066,N_7184);
nand U7319 (N_7319,N_7190,N_7030);
and U7320 (N_7320,N_7062,N_7094);
nor U7321 (N_7321,N_7170,N_7016);
and U7322 (N_7322,N_7021,N_7035);
nor U7323 (N_7323,N_7062,N_7120);
and U7324 (N_7324,N_7145,N_7123);
nor U7325 (N_7325,N_7078,N_7063);
nand U7326 (N_7326,N_7192,N_7144);
nor U7327 (N_7327,N_7026,N_7144);
nand U7328 (N_7328,N_7037,N_7147);
nand U7329 (N_7329,N_7051,N_7072);
or U7330 (N_7330,N_7141,N_7089);
xnor U7331 (N_7331,N_7007,N_7123);
nor U7332 (N_7332,N_7042,N_7144);
nand U7333 (N_7333,N_7125,N_7071);
nand U7334 (N_7334,N_7048,N_7183);
nand U7335 (N_7335,N_7090,N_7154);
nor U7336 (N_7336,N_7096,N_7178);
nand U7337 (N_7337,N_7139,N_7130);
xnor U7338 (N_7338,N_7115,N_7062);
or U7339 (N_7339,N_7185,N_7186);
nand U7340 (N_7340,N_7169,N_7011);
xnor U7341 (N_7341,N_7133,N_7119);
nand U7342 (N_7342,N_7078,N_7058);
nand U7343 (N_7343,N_7094,N_7135);
xnor U7344 (N_7344,N_7032,N_7147);
or U7345 (N_7345,N_7065,N_7076);
and U7346 (N_7346,N_7185,N_7059);
or U7347 (N_7347,N_7069,N_7067);
or U7348 (N_7348,N_7173,N_7182);
and U7349 (N_7349,N_7121,N_7154);
nand U7350 (N_7350,N_7038,N_7033);
nand U7351 (N_7351,N_7136,N_7156);
nand U7352 (N_7352,N_7033,N_7126);
xnor U7353 (N_7353,N_7116,N_7194);
xor U7354 (N_7354,N_7083,N_7053);
nor U7355 (N_7355,N_7122,N_7050);
or U7356 (N_7356,N_7095,N_7124);
and U7357 (N_7357,N_7024,N_7173);
nor U7358 (N_7358,N_7033,N_7113);
nand U7359 (N_7359,N_7156,N_7075);
and U7360 (N_7360,N_7165,N_7057);
xor U7361 (N_7361,N_7022,N_7015);
xnor U7362 (N_7362,N_7167,N_7065);
xor U7363 (N_7363,N_7064,N_7184);
or U7364 (N_7364,N_7101,N_7193);
xor U7365 (N_7365,N_7019,N_7007);
xor U7366 (N_7366,N_7089,N_7071);
nand U7367 (N_7367,N_7131,N_7125);
nand U7368 (N_7368,N_7100,N_7021);
xnor U7369 (N_7369,N_7182,N_7178);
nand U7370 (N_7370,N_7006,N_7052);
and U7371 (N_7371,N_7038,N_7143);
or U7372 (N_7372,N_7016,N_7004);
nor U7373 (N_7373,N_7106,N_7195);
nor U7374 (N_7374,N_7147,N_7121);
and U7375 (N_7375,N_7119,N_7058);
xor U7376 (N_7376,N_7178,N_7132);
nand U7377 (N_7377,N_7148,N_7076);
nand U7378 (N_7378,N_7012,N_7182);
nor U7379 (N_7379,N_7180,N_7125);
or U7380 (N_7380,N_7157,N_7069);
nor U7381 (N_7381,N_7040,N_7159);
nor U7382 (N_7382,N_7062,N_7105);
nand U7383 (N_7383,N_7091,N_7114);
and U7384 (N_7384,N_7098,N_7109);
and U7385 (N_7385,N_7141,N_7041);
nor U7386 (N_7386,N_7106,N_7136);
nor U7387 (N_7387,N_7109,N_7002);
nand U7388 (N_7388,N_7126,N_7195);
xnor U7389 (N_7389,N_7136,N_7079);
or U7390 (N_7390,N_7086,N_7111);
xnor U7391 (N_7391,N_7087,N_7070);
nand U7392 (N_7392,N_7041,N_7004);
nand U7393 (N_7393,N_7037,N_7073);
and U7394 (N_7394,N_7173,N_7011);
and U7395 (N_7395,N_7059,N_7099);
and U7396 (N_7396,N_7116,N_7184);
or U7397 (N_7397,N_7022,N_7146);
and U7398 (N_7398,N_7061,N_7135);
or U7399 (N_7399,N_7071,N_7010);
nor U7400 (N_7400,N_7373,N_7266);
and U7401 (N_7401,N_7284,N_7322);
nand U7402 (N_7402,N_7247,N_7232);
and U7403 (N_7403,N_7345,N_7319);
xor U7404 (N_7404,N_7375,N_7392);
xnor U7405 (N_7405,N_7391,N_7293);
and U7406 (N_7406,N_7395,N_7393);
nor U7407 (N_7407,N_7304,N_7353);
xor U7408 (N_7408,N_7294,N_7399);
or U7409 (N_7409,N_7372,N_7226);
nor U7410 (N_7410,N_7383,N_7338);
xnor U7411 (N_7411,N_7291,N_7370);
or U7412 (N_7412,N_7287,N_7268);
xor U7413 (N_7413,N_7346,N_7314);
nor U7414 (N_7414,N_7224,N_7295);
nor U7415 (N_7415,N_7364,N_7378);
xnor U7416 (N_7416,N_7317,N_7361);
or U7417 (N_7417,N_7258,N_7257);
nand U7418 (N_7418,N_7341,N_7242);
or U7419 (N_7419,N_7347,N_7313);
nand U7420 (N_7420,N_7329,N_7398);
and U7421 (N_7421,N_7262,N_7215);
or U7422 (N_7422,N_7396,N_7264);
nand U7423 (N_7423,N_7235,N_7323);
nand U7424 (N_7424,N_7212,N_7316);
xor U7425 (N_7425,N_7325,N_7385);
or U7426 (N_7426,N_7336,N_7282);
nor U7427 (N_7427,N_7277,N_7339);
nand U7428 (N_7428,N_7209,N_7203);
nand U7429 (N_7429,N_7220,N_7332);
and U7430 (N_7430,N_7222,N_7286);
nor U7431 (N_7431,N_7388,N_7279);
and U7432 (N_7432,N_7327,N_7250);
nor U7433 (N_7433,N_7248,N_7231);
xor U7434 (N_7434,N_7280,N_7324);
nor U7435 (N_7435,N_7254,N_7205);
xor U7436 (N_7436,N_7208,N_7267);
nor U7437 (N_7437,N_7227,N_7305);
or U7438 (N_7438,N_7320,N_7359);
or U7439 (N_7439,N_7350,N_7290);
xnor U7440 (N_7440,N_7334,N_7269);
nand U7441 (N_7441,N_7337,N_7261);
nor U7442 (N_7442,N_7251,N_7263);
and U7443 (N_7443,N_7328,N_7214);
xnor U7444 (N_7444,N_7223,N_7233);
and U7445 (N_7445,N_7265,N_7239);
or U7446 (N_7446,N_7238,N_7389);
xnor U7447 (N_7447,N_7240,N_7394);
or U7448 (N_7448,N_7342,N_7340);
and U7449 (N_7449,N_7360,N_7289);
and U7450 (N_7450,N_7285,N_7218);
or U7451 (N_7451,N_7253,N_7275);
and U7452 (N_7452,N_7245,N_7260);
or U7453 (N_7453,N_7366,N_7200);
nand U7454 (N_7454,N_7367,N_7374);
nand U7455 (N_7455,N_7343,N_7376);
and U7456 (N_7456,N_7234,N_7246);
or U7457 (N_7457,N_7216,N_7201);
and U7458 (N_7458,N_7241,N_7272);
or U7459 (N_7459,N_7217,N_7243);
and U7460 (N_7460,N_7335,N_7274);
or U7461 (N_7461,N_7352,N_7387);
nor U7462 (N_7462,N_7296,N_7380);
xnor U7463 (N_7463,N_7303,N_7278);
nor U7464 (N_7464,N_7377,N_7276);
xor U7465 (N_7465,N_7299,N_7281);
or U7466 (N_7466,N_7369,N_7207);
nand U7467 (N_7467,N_7315,N_7236);
nand U7468 (N_7468,N_7365,N_7382);
and U7469 (N_7469,N_7368,N_7219);
nand U7470 (N_7470,N_7386,N_7255);
and U7471 (N_7471,N_7306,N_7318);
xor U7472 (N_7472,N_7330,N_7356);
nor U7473 (N_7473,N_7206,N_7283);
nand U7474 (N_7474,N_7273,N_7308);
and U7475 (N_7475,N_7309,N_7326);
and U7476 (N_7476,N_7225,N_7259);
or U7477 (N_7477,N_7354,N_7362);
xnor U7478 (N_7478,N_7210,N_7348);
nand U7479 (N_7479,N_7331,N_7390);
nor U7480 (N_7480,N_7288,N_7307);
or U7481 (N_7481,N_7228,N_7298);
nor U7482 (N_7482,N_7351,N_7311);
nor U7483 (N_7483,N_7384,N_7256);
and U7484 (N_7484,N_7252,N_7371);
xor U7485 (N_7485,N_7211,N_7301);
nand U7486 (N_7486,N_7249,N_7237);
xnor U7487 (N_7487,N_7355,N_7292);
nor U7488 (N_7488,N_7381,N_7204);
and U7489 (N_7489,N_7397,N_7363);
nor U7490 (N_7490,N_7302,N_7333);
or U7491 (N_7491,N_7213,N_7221);
or U7492 (N_7492,N_7349,N_7300);
and U7493 (N_7493,N_7230,N_7344);
xnor U7494 (N_7494,N_7310,N_7358);
and U7495 (N_7495,N_7229,N_7202);
nor U7496 (N_7496,N_7379,N_7271);
or U7497 (N_7497,N_7270,N_7321);
xnor U7498 (N_7498,N_7244,N_7312);
nand U7499 (N_7499,N_7297,N_7357);
nor U7500 (N_7500,N_7364,N_7363);
nor U7501 (N_7501,N_7372,N_7224);
nor U7502 (N_7502,N_7265,N_7330);
xnor U7503 (N_7503,N_7355,N_7206);
nand U7504 (N_7504,N_7248,N_7233);
nor U7505 (N_7505,N_7319,N_7349);
nor U7506 (N_7506,N_7368,N_7283);
or U7507 (N_7507,N_7333,N_7280);
or U7508 (N_7508,N_7322,N_7398);
and U7509 (N_7509,N_7342,N_7220);
nand U7510 (N_7510,N_7349,N_7363);
xnor U7511 (N_7511,N_7239,N_7241);
or U7512 (N_7512,N_7286,N_7314);
xnor U7513 (N_7513,N_7250,N_7306);
xor U7514 (N_7514,N_7263,N_7365);
and U7515 (N_7515,N_7322,N_7285);
nor U7516 (N_7516,N_7387,N_7257);
nand U7517 (N_7517,N_7300,N_7348);
nor U7518 (N_7518,N_7349,N_7261);
xor U7519 (N_7519,N_7372,N_7258);
xnor U7520 (N_7520,N_7257,N_7370);
nand U7521 (N_7521,N_7310,N_7312);
and U7522 (N_7522,N_7324,N_7245);
nand U7523 (N_7523,N_7366,N_7205);
nor U7524 (N_7524,N_7340,N_7321);
nor U7525 (N_7525,N_7319,N_7272);
or U7526 (N_7526,N_7214,N_7365);
nand U7527 (N_7527,N_7218,N_7351);
and U7528 (N_7528,N_7301,N_7261);
nor U7529 (N_7529,N_7362,N_7296);
or U7530 (N_7530,N_7202,N_7313);
nand U7531 (N_7531,N_7238,N_7352);
or U7532 (N_7532,N_7355,N_7361);
nand U7533 (N_7533,N_7321,N_7360);
or U7534 (N_7534,N_7242,N_7318);
or U7535 (N_7535,N_7346,N_7386);
and U7536 (N_7536,N_7361,N_7302);
and U7537 (N_7537,N_7299,N_7265);
or U7538 (N_7538,N_7279,N_7256);
or U7539 (N_7539,N_7354,N_7372);
xor U7540 (N_7540,N_7253,N_7309);
nand U7541 (N_7541,N_7333,N_7242);
xor U7542 (N_7542,N_7290,N_7268);
xnor U7543 (N_7543,N_7378,N_7270);
and U7544 (N_7544,N_7244,N_7343);
nor U7545 (N_7545,N_7210,N_7376);
xnor U7546 (N_7546,N_7356,N_7387);
and U7547 (N_7547,N_7347,N_7220);
nand U7548 (N_7548,N_7291,N_7349);
or U7549 (N_7549,N_7260,N_7361);
or U7550 (N_7550,N_7202,N_7396);
nor U7551 (N_7551,N_7370,N_7299);
xnor U7552 (N_7552,N_7330,N_7390);
xor U7553 (N_7553,N_7284,N_7221);
nand U7554 (N_7554,N_7348,N_7250);
nor U7555 (N_7555,N_7393,N_7228);
or U7556 (N_7556,N_7212,N_7243);
or U7557 (N_7557,N_7204,N_7241);
and U7558 (N_7558,N_7356,N_7396);
nor U7559 (N_7559,N_7356,N_7267);
or U7560 (N_7560,N_7275,N_7241);
xnor U7561 (N_7561,N_7249,N_7214);
and U7562 (N_7562,N_7220,N_7395);
xor U7563 (N_7563,N_7224,N_7203);
xnor U7564 (N_7564,N_7306,N_7307);
and U7565 (N_7565,N_7384,N_7364);
or U7566 (N_7566,N_7261,N_7391);
xnor U7567 (N_7567,N_7255,N_7269);
xor U7568 (N_7568,N_7353,N_7273);
nor U7569 (N_7569,N_7316,N_7336);
xor U7570 (N_7570,N_7226,N_7202);
nand U7571 (N_7571,N_7337,N_7387);
and U7572 (N_7572,N_7265,N_7319);
and U7573 (N_7573,N_7274,N_7321);
xnor U7574 (N_7574,N_7264,N_7301);
nor U7575 (N_7575,N_7202,N_7365);
or U7576 (N_7576,N_7228,N_7213);
nand U7577 (N_7577,N_7202,N_7357);
xor U7578 (N_7578,N_7356,N_7295);
xnor U7579 (N_7579,N_7293,N_7365);
and U7580 (N_7580,N_7234,N_7255);
or U7581 (N_7581,N_7375,N_7325);
or U7582 (N_7582,N_7266,N_7369);
or U7583 (N_7583,N_7257,N_7369);
xnor U7584 (N_7584,N_7246,N_7296);
nor U7585 (N_7585,N_7201,N_7236);
or U7586 (N_7586,N_7377,N_7251);
nand U7587 (N_7587,N_7246,N_7226);
or U7588 (N_7588,N_7284,N_7259);
nor U7589 (N_7589,N_7380,N_7237);
and U7590 (N_7590,N_7336,N_7338);
nor U7591 (N_7591,N_7364,N_7399);
xor U7592 (N_7592,N_7397,N_7285);
and U7593 (N_7593,N_7368,N_7251);
nor U7594 (N_7594,N_7297,N_7321);
or U7595 (N_7595,N_7398,N_7332);
or U7596 (N_7596,N_7357,N_7377);
or U7597 (N_7597,N_7382,N_7359);
nand U7598 (N_7598,N_7324,N_7261);
nand U7599 (N_7599,N_7249,N_7291);
xor U7600 (N_7600,N_7462,N_7492);
or U7601 (N_7601,N_7576,N_7489);
nand U7602 (N_7602,N_7466,N_7404);
nand U7603 (N_7603,N_7516,N_7551);
nor U7604 (N_7604,N_7411,N_7465);
or U7605 (N_7605,N_7405,N_7568);
nor U7606 (N_7606,N_7580,N_7447);
nor U7607 (N_7607,N_7486,N_7517);
or U7608 (N_7608,N_7452,N_7490);
xor U7609 (N_7609,N_7400,N_7569);
nor U7610 (N_7610,N_7575,N_7547);
and U7611 (N_7611,N_7444,N_7485);
and U7612 (N_7612,N_7415,N_7564);
nor U7613 (N_7613,N_7480,N_7402);
and U7614 (N_7614,N_7457,N_7539);
nor U7615 (N_7615,N_7582,N_7599);
and U7616 (N_7616,N_7595,N_7474);
nand U7617 (N_7617,N_7530,N_7585);
nand U7618 (N_7618,N_7426,N_7560);
nand U7619 (N_7619,N_7546,N_7443);
xnor U7620 (N_7620,N_7430,N_7449);
nor U7621 (N_7621,N_7495,N_7418);
xnor U7622 (N_7622,N_7523,N_7482);
nor U7623 (N_7623,N_7409,N_7428);
xnor U7624 (N_7624,N_7519,N_7522);
and U7625 (N_7625,N_7534,N_7429);
or U7626 (N_7626,N_7521,N_7561);
xor U7627 (N_7627,N_7513,N_7417);
nor U7628 (N_7628,N_7571,N_7434);
nand U7629 (N_7629,N_7491,N_7461);
and U7630 (N_7630,N_7588,N_7496);
or U7631 (N_7631,N_7590,N_7422);
or U7632 (N_7632,N_7584,N_7552);
xnor U7633 (N_7633,N_7460,N_7532);
nand U7634 (N_7634,N_7459,N_7597);
nand U7635 (N_7635,N_7499,N_7541);
and U7636 (N_7636,N_7544,N_7515);
xnor U7637 (N_7637,N_7476,N_7529);
nor U7638 (N_7638,N_7470,N_7506);
nand U7639 (N_7639,N_7512,N_7567);
or U7640 (N_7640,N_7412,N_7554);
nand U7641 (N_7641,N_7410,N_7440);
nand U7642 (N_7642,N_7503,N_7500);
or U7643 (N_7643,N_7536,N_7596);
and U7644 (N_7644,N_7493,N_7494);
xnor U7645 (N_7645,N_7420,N_7583);
nand U7646 (N_7646,N_7487,N_7566);
nor U7647 (N_7647,N_7414,N_7558);
and U7648 (N_7648,N_7510,N_7454);
xnor U7649 (N_7649,N_7548,N_7555);
nor U7650 (N_7650,N_7403,N_7537);
nor U7651 (N_7651,N_7456,N_7436);
nand U7652 (N_7652,N_7498,N_7477);
or U7653 (N_7653,N_7526,N_7559);
nand U7654 (N_7654,N_7473,N_7464);
and U7655 (N_7655,N_7587,N_7531);
xnor U7656 (N_7656,N_7518,N_7545);
and U7657 (N_7657,N_7525,N_7455);
or U7658 (N_7658,N_7445,N_7549);
nor U7659 (N_7659,N_7591,N_7425);
and U7660 (N_7660,N_7586,N_7472);
nand U7661 (N_7661,N_7504,N_7432);
nor U7662 (N_7662,N_7535,N_7553);
xor U7663 (N_7663,N_7435,N_7488);
nor U7664 (N_7664,N_7484,N_7598);
nand U7665 (N_7665,N_7565,N_7446);
nor U7666 (N_7666,N_7514,N_7483);
or U7667 (N_7667,N_7448,N_7401);
nor U7668 (N_7668,N_7505,N_7594);
and U7669 (N_7669,N_7451,N_7556);
and U7670 (N_7670,N_7538,N_7507);
nand U7671 (N_7671,N_7543,N_7509);
and U7672 (N_7672,N_7562,N_7577);
nor U7673 (N_7673,N_7468,N_7406);
nand U7674 (N_7674,N_7592,N_7433);
nand U7675 (N_7675,N_7579,N_7475);
xor U7676 (N_7676,N_7502,N_7581);
nand U7677 (N_7677,N_7423,N_7478);
or U7678 (N_7678,N_7463,N_7557);
or U7679 (N_7679,N_7424,N_7408);
xnor U7680 (N_7680,N_7467,N_7453);
xnor U7681 (N_7681,N_7441,N_7550);
xnor U7682 (N_7682,N_7574,N_7578);
and U7683 (N_7683,N_7439,N_7407);
nor U7684 (N_7684,N_7442,N_7413);
or U7685 (N_7685,N_7416,N_7438);
or U7686 (N_7686,N_7508,N_7542);
or U7687 (N_7687,N_7427,N_7570);
nor U7688 (N_7688,N_7524,N_7419);
nand U7689 (N_7689,N_7501,N_7469);
nor U7690 (N_7690,N_7497,N_7572);
xor U7691 (N_7691,N_7573,N_7563);
and U7692 (N_7692,N_7431,N_7528);
nand U7693 (N_7693,N_7527,N_7511);
nor U7694 (N_7694,N_7533,N_7421);
nand U7695 (N_7695,N_7450,N_7471);
or U7696 (N_7696,N_7593,N_7540);
or U7697 (N_7697,N_7458,N_7437);
or U7698 (N_7698,N_7479,N_7481);
nor U7699 (N_7699,N_7520,N_7589);
nor U7700 (N_7700,N_7428,N_7416);
and U7701 (N_7701,N_7582,N_7451);
or U7702 (N_7702,N_7454,N_7410);
nor U7703 (N_7703,N_7499,N_7532);
and U7704 (N_7704,N_7447,N_7494);
xor U7705 (N_7705,N_7449,N_7472);
xor U7706 (N_7706,N_7478,N_7441);
nand U7707 (N_7707,N_7569,N_7444);
or U7708 (N_7708,N_7436,N_7538);
nand U7709 (N_7709,N_7504,N_7495);
and U7710 (N_7710,N_7476,N_7553);
xnor U7711 (N_7711,N_7450,N_7588);
and U7712 (N_7712,N_7411,N_7469);
and U7713 (N_7713,N_7527,N_7425);
and U7714 (N_7714,N_7488,N_7483);
and U7715 (N_7715,N_7475,N_7578);
nand U7716 (N_7716,N_7490,N_7485);
nor U7717 (N_7717,N_7497,N_7478);
nand U7718 (N_7718,N_7457,N_7581);
nor U7719 (N_7719,N_7505,N_7574);
or U7720 (N_7720,N_7523,N_7410);
nand U7721 (N_7721,N_7551,N_7456);
nor U7722 (N_7722,N_7463,N_7544);
or U7723 (N_7723,N_7504,N_7494);
nor U7724 (N_7724,N_7408,N_7565);
and U7725 (N_7725,N_7480,N_7446);
and U7726 (N_7726,N_7483,N_7577);
xnor U7727 (N_7727,N_7551,N_7468);
xor U7728 (N_7728,N_7575,N_7473);
nor U7729 (N_7729,N_7594,N_7410);
nor U7730 (N_7730,N_7465,N_7440);
nand U7731 (N_7731,N_7599,N_7534);
xor U7732 (N_7732,N_7403,N_7599);
and U7733 (N_7733,N_7511,N_7463);
nand U7734 (N_7734,N_7504,N_7468);
or U7735 (N_7735,N_7414,N_7483);
nand U7736 (N_7736,N_7423,N_7561);
nand U7737 (N_7737,N_7429,N_7508);
nand U7738 (N_7738,N_7500,N_7522);
and U7739 (N_7739,N_7481,N_7581);
nor U7740 (N_7740,N_7585,N_7406);
xnor U7741 (N_7741,N_7528,N_7474);
nor U7742 (N_7742,N_7420,N_7550);
or U7743 (N_7743,N_7464,N_7596);
xor U7744 (N_7744,N_7521,N_7527);
xor U7745 (N_7745,N_7455,N_7480);
xor U7746 (N_7746,N_7406,N_7586);
xnor U7747 (N_7747,N_7480,N_7560);
nor U7748 (N_7748,N_7562,N_7409);
nor U7749 (N_7749,N_7441,N_7500);
and U7750 (N_7750,N_7517,N_7463);
nand U7751 (N_7751,N_7520,N_7429);
xnor U7752 (N_7752,N_7515,N_7485);
and U7753 (N_7753,N_7533,N_7414);
nand U7754 (N_7754,N_7436,N_7588);
xor U7755 (N_7755,N_7532,N_7454);
nand U7756 (N_7756,N_7558,N_7508);
and U7757 (N_7757,N_7443,N_7456);
nand U7758 (N_7758,N_7445,N_7425);
or U7759 (N_7759,N_7482,N_7465);
nor U7760 (N_7760,N_7489,N_7587);
nand U7761 (N_7761,N_7523,N_7577);
or U7762 (N_7762,N_7449,N_7492);
xnor U7763 (N_7763,N_7489,N_7581);
nor U7764 (N_7764,N_7464,N_7562);
nor U7765 (N_7765,N_7429,N_7594);
xor U7766 (N_7766,N_7419,N_7523);
and U7767 (N_7767,N_7485,N_7577);
xnor U7768 (N_7768,N_7402,N_7462);
or U7769 (N_7769,N_7517,N_7548);
or U7770 (N_7770,N_7514,N_7448);
or U7771 (N_7771,N_7440,N_7472);
nand U7772 (N_7772,N_7436,N_7591);
nor U7773 (N_7773,N_7567,N_7456);
xnor U7774 (N_7774,N_7488,N_7431);
nor U7775 (N_7775,N_7520,N_7417);
xnor U7776 (N_7776,N_7552,N_7527);
xor U7777 (N_7777,N_7534,N_7551);
xor U7778 (N_7778,N_7430,N_7582);
nor U7779 (N_7779,N_7599,N_7419);
nand U7780 (N_7780,N_7468,N_7422);
and U7781 (N_7781,N_7460,N_7510);
and U7782 (N_7782,N_7417,N_7529);
nor U7783 (N_7783,N_7493,N_7578);
or U7784 (N_7784,N_7484,N_7490);
and U7785 (N_7785,N_7470,N_7423);
or U7786 (N_7786,N_7567,N_7511);
xor U7787 (N_7787,N_7523,N_7466);
nand U7788 (N_7788,N_7548,N_7497);
nand U7789 (N_7789,N_7406,N_7505);
nor U7790 (N_7790,N_7585,N_7575);
and U7791 (N_7791,N_7595,N_7442);
xnor U7792 (N_7792,N_7565,N_7430);
or U7793 (N_7793,N_7492,N_7446);
xnor U7794 (N_7794,N_7402,N_7456);
or U7795 (N_7795,N_7502,N_7582);
or U7796 (N_7796,N_7574,N_7528);
and U7797 (N_7797,N_7535,N_7408);
nor U7798 (N_7798,N_7551,N_7404);
xnor U7799 (N_7799,N_7469,N_7401);
nor U7800 (N_7800,N_7682,N_7698);
nor U7801 (N_7801,N_7726,N_7681);
and U7802 (N_7802,N_7624,N_7627);
nand U7803 (N_7803,N_7699,N_7655);
nor U7804 (N_7804,N_7664,N_7725);
xor U7805 (N_7805,N_7781,N_7622);
nand U7806 (N_7806,N_7694,N_7625);
nor U7807 (N_7807,N_7665,N_7678);
nor U7808 (N_7808,N_7673,N_7676);
xnor U7809 (N_7809,N_7734,N_7609);
or U7810 (N_7810,N_7789,N_7656);
nand U7811 (N_7811,N_7666,N_7718);
and U7812 (N_7812,N_7610,N_7631);
nor U7813 (N_7813,N_7707,N_7629);
and U7814 (N_7814,N_7604,N_7790);
nand U7815 (N_7815,N_7640,N_7647);
nor U7816 (N_7816,N_7763,N_7738);
and U7817 (N_7817,N_7689,N_7628);
and U7818 (N_7818,N_7639,N_7705);
xor U7819 (N_7819,N_7747,N_7688);
and U7820 (N_7820,N_7630,N_7772);
nand U7821 (N_7821,N_7644,N_7785);
xnor U7822 (N_7822,N_7691,N_7788);
xnor U7823 (N_7823,N_7633,N_7671);
or U7824 (N_7824,N_7617,N_7724);
nor U7825 (N_7825,N_7693,N_7708);
and U7826 (N_7826,N_7746,N_7775);
and U7827 (N_7827,N_7635,N_7687);
and U7828 (N_7828,N_7751,N_7715);
nand U7829 (N_7829,N_7607,N_7722);
nor U7830 (N_7830,N_7720,N_7713);
and U7831 (N_7831,N_7701,N_7748);
xor U7832 (N_7832,N_7677,N_7780);
and U7833 (N_7833,N_7754,N_7723);
and U7834 (N_7834,N_7762,N_7766);
or U7835 (N_7835,N_7768,N_7663);
and U7836 (N_7836,N_7615,N_7614);
and U7837 (N_7837,N_7741,N_7774);
nand U7838 (N_7838,N_7638,N_7618);
xor U7839 (N_7839,N_7733,N_7684);
or U7840 (N_7840,N_7773,N_7784);
and U7841 (N_7841,N_7795,N_7716);
nand U7842 (N_7842,N_7692,N_7658);
xor U7843 (N_7843,N_7645,N_7755);
nand U7844 (N_7844,N_7714,N_7674);
xor U7845 (N_7845,N_7745,N_7637);
and U7846 (N_7846,N_7744,N_7668);
or U7847 (N_7847,N_7728,N_7606);
xor U7848 (N_7848,N_7709,N_7632);
xnor U7849 (N_7849,N_7777,N_7753);
and U7850 (N_7850,N_7736,N_7662);
nand U7851 (N_7851,N_7605,N_7685);
nand U7852 (N_7852,N_7659,N_7739);
nand U7853 (N_7853,N_7634,N_7704);
nor U7854 (N_7854,N_7783,N_7752);
nor U7855 (N_7855,N_7670,N_7651);
nor U7856 (N_7856,N_7641,N_7727);
xnor U7857 (N_7857,N_7799,N_7697);
and U7858 (N_7858,N_7729,N_7760);
nand U7859 (N_7859,N_7652,N_7782);
xnor U7860 (N_7860,N_7616,N_7657);
or U7861 (N_7861,N_7761,N_7717);
nand U7862 (N_7862,N_7758,N_7667);
nand U7863 (N_7863,N_7711,N_7756);
xor U7864 (N_7864,N_7750,N_7740);
or U7865 (N_7865,N_7792,N_7643);
or U7866 (N_7866,N_7731,N_7686);
or U7867 (N_7867,N_7767,N_7742);
nand U7868 (N_7868,N_7675,N_7702);
xor U7869 (N_7869,N_7796,N_7703);
xnor U7870 (N_7870,N_7613,N_7710);
or U7871 (N_7871,N_7737,N_7769);
nand U7872 (N_7872,N_7778,N_7794);
nor U7873 (N_7873,N_7735,N_7650);
nand U7874 (N_7874,N_7621,N_7683);
nand U7875 (N_7875,N_7786,N_7636);
and U7876 (N_7876,N_7757,N_7672);
and U7877 (N_7877,N_7791,N_7603);
xnor U7878 (N_7878,N_7661,N_7743);
xor U7879 (N_7879,N_7770,N_7649);
nor U7880 (N_7880,N_7797,N_7660);
xnor U7881 (N_7881,N_7787,N_7700);
nand U7882 (N_7882,N_7653,N_7623);
or U7883 (N_7883,N_7669,N_7679);
and U7884 (N_7884,N_7619,N_7690);
nand U7885 (N_7885,N_7793,N_7732);
or U7886 (N_7886,N_7601,N_7608);
xnor U7887 (N_7887,N_7764,N_7654);
nand U7888 (N_7888,N_7730,N_7611);
or U7889 (N_7889,N_7759,N_7696);
xor U7890 (N_7890,N_7648,N_7642);
nor U7891 (N_7891,N_7646,N_7719);
nor U7892 (N_7892,N_7776,N_7680);
and U7893 (N_7893,N_7706,N_7695);
xnor U7894 (N_7894,N_7721,N_7749);
nand U7895 (N_7895,N_7602,N_7612);
and U7896 (N_7896,N_7626,N_7600);
xnor U7897 (N_7897,N_7765,N_7712);
xnor U7898 (N_7898,N_7779,N_7620);
and U7899 (N_7899,N_7798,N_7771);
or U7900 (N_7900,N_7759,N_7713);
or U7901 (N_7901,N_7792,N_7765);
nand U7902 (N_7902,N_7645,N_7641);
nor U7903 (N_7903,N_7688,N_7640);
nor U7904 (N_7904,N_7605,N_7643);
and U7905 (N_7905,N_7797,N_7637);
or U7906 (N_7906,N_7739,N_7784);
nand U7907 (N_7907,N_7733,N_7719);
or U7908 (N_7908,N_7791,N_7759);
and U7909 (N_7909,N_7619,N_7787);
xnor U7910 (N_7910,N_7646,N_7602);
and U7911 (N_7911,N_7719,N_7735);
xor U7912 (N_7912,N_7657,N_7776);
or U7913 (N_7913,N_7761,N_7770);
nor U7914 (N_7914,N_7675,N_7780);
xor U7915 (N_7915,N_7777,N_7669);
nand U7916 (N_7916,N_7618,N_7609);
or U7917 (N_7917,N_7799,N_7636);
and U7918 (N_7918,N_7690,N_7691);
and U7919 (N_7919,N_7680,N_7777);
and U7920 (N_7920,N_7797,N_7619);
nor U7921 (N_7921,N_7686,N_7751);
nand U7922 (N_7922,N_7762,N_7709);
and U7923 (N_7923,N_7714,N_7735);
nor U7924 (N_7924,N_7742,N_7776);
or U7925 (N_7925,N_7651,N_7671);
and U7926 (N_7926,N_7695,N_7691);
or U7927 (N_7927,N_7772,N_7681);
xor U7928 (N_7928,N_7765,N_7767);
nor U7929 (N_7929,N_7677,N_7711);
and U7930 (N_7930,N_7789,N_7630);
and U7931 (N_7931,N_7756,N_7701);
xor U7932 (N_7932,N_7653,N_7635);
and U7933 (N_7933,N_7719,N_7641);
or U7934 (N_7934,N_7688,N_7676);
nor U7935 (N_7935,N_7767,N_7645);
nand U7936 (N_7936,N_7600,N_7644);
nand U7937 (N_7937,N_7714,N_7739);
and U7938 (N_7938,N_7708,N_7721);
nor U7939 (N_7939,N_7773,N_7736);
nand U7940 (N_7940,N_7689,N_7730);
xor U7941 (N_7941,N_7635,N_7774);
nor U7942 (N_7942,N_7696,N_7698);
xor U7943 (N_7943,N_7626,N_7628);
and U7944 (N_7944,N_7673,N_7774);
nor U7945 (N_7945,N_7767,N_7789);
nor U7946 (N_7946,N_7700,N_7664);
and U7947 (N_7947,N_7775,N_7714);
nand U7948 (N_7948,N_7797,N_7603);
nor U7949 (N_7949,N_7768,N_7678);
xnor U7950 (N_7950,N_7650,N_7676);
and U7951 (N_7951,N_7784,N_7791);
nor U7952 (N_7952,N_7706,N_7631);
xor U7953 (N_7953,N_7663,N_7782);
and U7954 (N_7954,N_7725,N_7624);
and U7955 (N_7955,N_7681,N_7622);
nor U7956 (N_7956,N_7793,N_7703);
nor U7957 (N_7957,N_7779,N_7782);
nor U7958 (N_7958,N_7781,N_7668);
xnor U7959 (N_7959,N_7661,N_7713);
or U7960 (N_7960,N_7684,N_7742);
nor U7961 (N_7961,N_7754,N_7678);
or U7962 (N_7962,N_7755,N_7644);
and U7963 (N_7963,N_7694,N_7720);
or U7964 (N_7964,N_7754,N_7632);
nand U7965 (N_7965,N_7770,N_7781);
or U7966 (N_7966,N_7717,N_7684);
and U7967 (N_7967,N_7716,N_7624);
nor U7968 (N_7968,N_7739,N_7740);
nand U7969 (N_7969,N_7781,N_7783);
nor U7970 (N_7970,N_7734,N_7627);
or U7971 (N_7971,N_7718,N_7625);
or U7972 (N_7972,N_7735,N_7755);
nor U7973 (N_7973,N_7670,N_7729);
and U7974 (N_7974,N_7606,N_7652);
nand U7975 (N_7975,N_7690,N_7661);
nor U7976 (N_7976,N_7791,N_7643);
and U7977 (N_7977,N_7661,N_7609);
or U7978 (N_7978,N_7608,N_7688);
or U7979 (N_7979,N_7722,N_7625);
or U7980 (N_7980,N_7715,N_7606);
or U7981 (N_7981,N_7734,N_7712);
nor U7982 (N_7982,N_7682,N_7628);
xor U7983 (N_7983,N_7612,N_7755);
xor U7984 (N_7984,N_7732,N_7779);
or U7985 (N_7985,N_7724,N_7779);
or U7986 (N_7986,N_7673,N_7671);
nor U7987 (N_7987,N_7762,N_7727);
and U7988 (N_7988,N_7791,N_7622);
xor U7989 (N_7989,N_7643,N_7664);
and U7990 (N_7990,N_7688,N_7644);
and U7991 (N_7991,N_7617,N_7635);
nor U7992 (N_7992,N_7748,N_7796);
and U7993 (N_7993,N_7765,N_7745);
or U7994 (N_7994,N_7776,N_7672);
xor U7995 (N_7995,N_7669,N_7710);
xor U7996 (N_7996,N_7618,N_7669);
and U7997 (N_7997,N_7671,N_7601);
and U7998 (N_7998,N_7638,N_7726);
nand U7999 (N_7999,N_7690,N_7789);
nand U8000 (N_8000,N_7947,N_7943);
nor U8001 (N_8001,N_7906,N_7829);
and U8002 (N_8002,N_7806,N_7884);
xor U8003 (N_8003,N_7877,N_7814);
xnor U8004 (N_8004,N_7976,N_7842);
nor U8005 (N_8005,N_7846,N_7845);
or U8006 (N_8006,N_7808,N_7968);
nand U8007 (N_8007,N_7830,N_7953);
and U8008 (N_8008,N_7855,N_7997);
nand U8009 (N_8009,N_7853,N_7944);
xnor U8010 (N_8010,N_7983,N_7898);
nand U8011 (N_8011,N_7820,N_7990);
nand U8012 (N_8012,N_7979,N_7902);
xor U8013 (N_8013,N_7986,N_7818);
nor U8014 (N_8014,N_7803,N_7858);
and U8015 (N_8015,N_7825,N_7962);
nor U8016 (N_8016,N_7856,N_7913);
nand U8017 (N_8017,N_7907,N_7876);
or U8018 (N_8018,N_7920,N_7908);
or U8019 (N_8019,N_7927,N_7992);
and U8020 (N_8020,N_7926,N_7885);
xor U8021 (N_8021,N_7869,N_7859);
or U8022 (N_8022,N_7928,N_7975);
xor U8023 (N_8023,N_7958,N_7952);
and U8024 (N_8024,N_7994,N_7900);
xor U8025 (N_8025,N_7903,N_7981);
or U8026 (N_8026,N_7870,N_7833);
xnor U8027 (N_8027,N_7824,N_7939);
or U8028 (N_8028,N_7946,N_7888);
and U8029 (N_8029,N_7895,N_7923);
and U8030 (N_8030,N_7889,N_7977);
or U8031 (N_8031,N_7932,N_7973);
nor U8032 (N_8032,N_7937,N_7921);
or U8033 (N_8033,N_7866,N_7989);
nor U8034 (N_8034,N_7852,N_7960);
nor U8035 (N_8035,N_7998,N_7995);
and U8036 (N_8036,N_7987,N_7872);
nand U8037 (N_8037,N_7942,N_7816);
nor U8038 (N_8038,N_7822,N_7919);
nand U8039 (N_8039,N_7837,N_7864);
nor U8040 (N_8040,N_7810,N_7915);
nor U8041 (N_8041,N_7828,N_7894);
nand U8042 (N_8042,N_7867,N_7980);
or U8043 (N_8043,N_7911,N_7883);
or U8044 (N_8044,N_7967,N_7891);
or U8045 (N_8045,N_7925,N_7809);
nand U8046 (N_8046,N_7899,N_7938);
xnor U8047 (N_8047,N_7892,N_7933);
nor U8048 (N_8048,N_7914,N_7969);
nand U8049 (N_8049,N_7880,N_7811);
or U8050 (N_8050,N_7917,N_7812);
nand U8051 (N_8051,N_7916,N_7991);
nand U8052 (N_8052,N_7918,N_7924);
nand U8053 (N_8053,N_7861,N_7988);
nand U8054 (N_8054,N_7972,N_7857);
nor U8055 (N_8055,N_7959,N_7936);
or U8056 (N_8056,N_7881,N_7996);
nand U8057 (N_8057,N_7868,N_7948);
nor U8058 (N_8058,N_7865,N_7912);
nor U8059 (N_8059,N_7905,N_7887);
or U8060 (N_8060,N_7823,N_7854);
or U8061 (N_8061,N_7955,N_7984);
nor U8062 (N_8062,N_7974,N_7850);
nor U8063 (N_8063,N_7930,N_7807);
nand U8064 (N_8064,N_7843,N_7826);
or U8065 (N_8065,N_7831,N_7945);
or U8066 (N_8066,N_7954,N_7951);
and U8067 (N_8067,N_7805,N_7863);
nand U8068 (N_8068,N_7890,N_7878);
or U8069 (N_8069,N_7896,N_7874);
nor U8070 (N_8070,N_7931,N_7964);
nor U8071 (N_8071,N_7804,N_7886);
nand U8072 (N_8072,N_7978,N_7966);
nand U8073 (N_8073,N_7963,N_7838);
nor U8074 (N_8074,N_7839,N_7832);
xnor U8075 (N_8075,N_7834,N_7922);
or U8076 (N_8076,N_7909,N_7949);
nand U8077 (N_8077,N_7836,N_7844);
xor U8078 (N_8078,N_7848,N_7940);
or U8079 (N_8079,N_7815,N_7813);
xnor U8080 (N_8080,N_7819,N_7941);
nor U8081 (N_8081,N_7957,N_7851);
nand U8082 (N_8082,N_7901,N_7993);
nand U8083 (N_8083,N_7897,N_7882);
and U8084 (N_8084,N_7827,N_7934);
and U8085 (N_8085,N_7904,N_7802);
nor U8086 (N_8086,N_7879,N_7801);
nand U8087 (N_8087,N_7860,N_7817);
xnor U8088 (N_8088,N_7910,N_7961);
or U8089 (N_8089,N_7841,N_7935);
or U8090 (N_8090,N_7956,N_7982);
nand U8091 (N_8091,N_7950,N_7821);
xnor U8092 (N_8092,N_7971,N_7893);
nor U8093 (N_8093,N_7965,N_7835);
nand U8094 (N_8094,N_7873,N_7847);
nand U8095 (N_8095,N_7929,N_7875);
nor U8096 (N_8096,N_7970,N_7840);
and U8097 (N_8097,N_7985,N_7871);
nor U8098 (N_8098,N_7849,N_7800);
nand U8099 (N_8099,N_7862,N_7999);
nor U8100 (N_8100,N_7945,N_7908);
or U8101 (N_8101,N_7887,N_7809);
or U8102 (N_8102,N_7956,N_7892);
or U8103 (N_8103,N_7878,N_7853);
xnor U8104 (N_8104,N_7824,N_7991);
xnor U8105 (N_8105,N_7979,N_7915);
xor U8106 (N_8106,N_7995,N_7872);
and U8107 (N_8107,N_7971,N_7966);
or U8108 (N_8108,N_7884,N_7877);
xor U8109 (N_8109,N_7886,N_7806);
xnor U8110 (N_8110,N_7867,N_7806);
nor U8111 (N_8111,N_7800,N_7991);
nand U8112 (N_8112,N_7869,N_7940);
nand U8113 (N_8113,N_7848,N_7931);
nor U8114 (N_8114,N_7917,N_7925);
or U8115 (N_8115,N_7965,N_7841);
nor U8116 (N_8116,N_7966,N_7852);
and U8117 (N_8117,N_7906,N_7943);
or U8118 (N_8118,N_7818,N_7900);
nand U8119 (N_8119,N_7930,N_7887);
nor U8120 (N_8120,N_7842,N_7981);
or U8121 (N_8121,N_7938,N_7802);
or U8122 (N_8122,N_7861,N_7972);
nor U8123 (N_8123,N_7968,N_7805);
or U8124 (N_8124,N_7942,N_7940);
or U8125 (N_8125,N_7984,N_7895);
xor U8126 (N_8126,N_7943,N_7994);
or U8127 (N_8127,N_7852,N_7921);
xnor U8128 (N_8128,N_7929,N_7969);
or U8129 (N_8129,N_7875,N_7971);
or U8130 (N_8130,N_7851,N_7814);
or U8131 (N_8131,N_7957,N_7937);
xnor U8132 (N_8132,N_7879,N_7857);
nor U8133 (N_8133,N_7879,N_7968);
xor U8134 (N_8134,N_7923,N_7800);
nand U8135 (N_8135,N_7953,N_7871);
xor U8136 (N_8136,N_7871,N_7906);
and U8137 (N_8137,N_7996,N_7895);
nand U8138 (N_8138,N_7871,N_7813);
nor U8139 (N_8139,N_7830,N_7815);
xnor U8140 (N_8140,N_7865,N_7883);
or U8141 (N_8141,N_7881,N_7921);
xor U8142 (N_8142,N_7967,N_7853);
or U8143 (N_8143,N_7975,N_7968);
nor U8144 (N_8144,N_7840,N_7959);
nor U8145 (N_8145,N_7936,N_7852);
nor U8146 (N_8146,N_7861,N_7953);
xor U8147 (N_8147,N_7910,N_7835);
nand U8148 (N_8148,N_7911,N_7984);
nor U8149 (N_8149,N_7843,N_7828);
nor U8150 (N_8150,N_7918,N_7804);
and U8151 (N_8151,N_7828,N_7895);
and U8152 (N_8152,N_7892,N_7894);
and U8153 (N_8153,N_7872,N_7918);
and U8154 (N_8154,N_7948,N_7955);
and U8155 (N_8155,N_7845,N_7972);
and U8156 (N_8156,N_7848,N_7972);
or U8157 (N_8157,N_7923,N_7907);
or U8158 (N_8158,N_7881,N_7963);
xnor U8159 (N_8159,N_7996,N_7866);
nor U8160 (N_8160,N_7946,N_7940);
nand U8161 (N_8161,N_7833,N_7982);
or U8162 (N_8162,N_7852,N_7875);
or U8163 (N_8163,N_7908,N_7937);
or U8164 (N_8164,N_7958,N_7920);
or U8165 (N_8165,N_7944,N_7960);
xor U8166 (N_8166,N_7879,N_7945);
nand U8167 (N_8167,N_7824,N_7878);
nand U8168 (N_8168,N_7833,N_7925);
nand U8169 (N_8169,N_7896,N_7831);
or U8170 (N_8170,N_7961,N_7974);
nor U8171 (N_8171,N_7978,N_7869);
nor U8172 (N_8172,N_7863,N_7985);
and U8173 (N_8173,N_7830,N_7930);
xnor U8174 (N_8174,N_7907,N_7884);
and U8175 (N_8175,N_7801,N_7848);
nand U8176 (N_8176,N_7819,N_7861);
nor U8177 (N_8177,N_7986,N_7922);
nor U8178 (N_8178,N_7939,N_7881);
or U8179 (N_8179,N_7800,N_7911);
nand U8180 (N_8180,N_7983,N_7952);
xor U8181 (N_8181,N_7977,N_7916);
or U8182 (N_8182,N_7984,N_7963);
and U8183 (N_8183,N_7913,N_7847);
or U8184 (N_8184,N_7827,N_7992);
nand U8185 (N_8185,N_7903,N_7946);
nand U8186 (N_8186,N_7838,N_7879);
and U8187 (N_8187,N_7952,N_7828);
xnor U8188 (N_8188,N_7977,N_7972);
nand U8189 (N_8189,N_7963,N_7876);
and U8190 (N_8190,N_7980,N_7960);
and U8191 (N_8191,N_7958,N_7940);
xnor U8192 (N_8192,N_7944,N_7808);
xor U8193 (N_8193,N_7803,N_7990);
xnor U8194 (N_8194,N_7944,N_7846);
or U8195 (N_8195,N_7947,N_7912);
xor U8196 (N_8196,N_7822,N_7844);
or U8197 (N_8197,N_7945,N_7917);
nand U8198 (N_8198,N_7948,N_7869);
and U8199 (N_8199,N_7861,N_7964);
xnor U8200 (N_8200,N_8116,N_8042);
or U8201 (N_8201,N_8081,N_8144);
xnor U8202 (N_8202,N_8126,N_8095);
nor U8203 (N_8203,N_8053,N_8077);
nor U8204 (N_8204,N_8000,N_8115);
or U8205 (N_8205,N_8059,N_8114);
and U8206 (N_8206,N_8047,N_8195);
nand U8207 (N_8207,N_8036,N_8146);
and U8208 (N_8208,N_8045,N_8064);
nor U8209 (N_8209,N_8092,N_8039);
or U8210 (N_8210,N_8041,N_8100);
nand U8211 (N_8211,N_8179,N_8063);
and U8212 (N_8212,N_8139,N_8050);
nor U8213 (N_8213,N_8186,N_8178);
nor U8214 (N_8214,N_8133,N_8082);
xor U8215 (N_8215,N_8070,N_8005);
or U8216 (N_8216,N_8011,N_8072);
nand U8217 (N_8217,N_8054,N_8049);
xor U8218 (N_8218,N_8127,N_8198);
or U8219 (N_8219,N_8154,N_8008);
xnor U8220 (N_8220,N_8018,N_8019);
nor U8221 (N_8221,N_8128,N_8142);
and U8222 (N_8222,N_8194,N_8130);
nand U8223 (N_8223,N_8079,N_8105);
nand U8224 (N_8224,N_8062,N_8013);
xnor U8225 (N_8225,N_8057,N_8035);
and U8226 (N_8226,N_8102,N_8060);
and U8227 (N_8227,N_8086,N_8068);
or U8228 (N_8228,N_8046,N_8040);
nand U8229 (N_8229,N_8104,N_8058);
nand U8230 (N_8230,N_8074,N_8101);
and U8231 (N_8231,N_8165,N_8107);
and U8232 (N_8232,N_8141,N_8015);
or U8233 (N_8233,N_8123,N_8143);
or U8234 (N_8234,N_8112,N_8188);
and U8235 (N_8235,N_8038,N_8026);
and U8236 (N_8236,N_8106,N_8030);
and U8237 (N_8237,N_8012,N_8199);
xor U8238 (N_8238,N_8065,N_8134);
nand U8239 (N_8239,N_8177,N_8121);
or U8240 (N_8240,N_8187,N_8073);
or U8241 (N_8241,N_8191,N_8131);
xnor U8242 (N_8242,N_8003,N_8163);
or U8243 (N_8243,N_8006,N_8167);
or U8244 (N_8244,N_8031,N_8002);
xor U8245 (N_8245,N_8151,N_8009);
and U8246 (N_8246,N_8088,N_8025);
and U8247 (N_8247,N_8029,N_8098);
nand U8248 (N_8248,N_8111,N_8172);
and U8249 (N_8249,N_8132,N_8067);
nor U8250 (N_8250,N_8158,N_8166);
or U8251 (N_8251,N_8090,N_8093);
or U8252 (N_8252,N_8122,N_8148);
or U8253 (N_8253,N_8118,N_8007);
or U8254 (N_8254,N_8091,N_8022);
and U8255 (N_8255,N_8168,N_8159);
or U8256 (N_8256,N_8014,N_8017);
or U8257 (N_8257,N_8185,N_8021);
nor U8258 (N_8258,N_8169,N_8083);
and U8259 (N_8259,N_8028,N_8037);
xnor U8260 (N_8260,N_8197,N_8182);
xnor U8261 (N_8261,N_8135,N_8183);
or U8262 (N_8262,N_8066,N_8056);
or U8263 (N_8263,N_8173,N_8170);
nor U8264 (N_8264,N_8080,N_8193);
or U8265 (N_8265,N_8164,N_8103);
nor U8266 (N_8266,N_8150,N_8117);
nand U8267 (N_8267,N_8024,N_8157);
xor U8268 (N_8268,N_8156,N_8001);
and U8269 (N_8269,N_8153,N_8110);
nor U8270 (N_8270,N_8109,N_8181);
nand U8271 (N_8271,N_8180,N_8176);
or U8272 (N_8272,N_8147,N_8189);
or U8273 (N_8273,N_8087,N_8094);
nor U8274 (N_8274,N_8125,N_8078);
or U8275 (N_8275,N_8023,N_8033);
and U8276 (N_8276,N_8196,N_8108);
and U8277 (N_8277,N_8085,N_8138);
nor U8278 (N_8278,N_8145,N_8113);
or U8279 (N_8279,N_8099,N_8160);
xor U8280 (N_8280,N_8097,N_8010);
nand U8281 (N_8281,N_8152,N_8137);
or U8282 (N_8282,N_8192,N_8075);
nor U8283 (N_8283,N_8051,N_8061);
nand U8284 (N_8284,N_8120,N_8124);
and U8285 (N_8285,N_8076,N_8155);
nor U8286 (N_8286,N_8052,N_8044);
and U8287 (N_8287,N_8162,N_8184);
or U8288 (N_8288,N_8048,N_8055);
xor U8289 (N_8289,N_8027,N_8174);
and U8290 (N_8290,N_8190,N_8071);
nor U8291 (N_8291,N_8016,N_8096);
nand U8292 (N_8292,N_8175,N_8171);
nand U8293 (N_8293,N_8136,N_8089);
nand U8294 (N_8294,N_8069,N_8034);
nor U8295 (N_8295,N_8119,N_8129);
xor U8296 (N_8296,N_8140,N_8004);
and U8297 (N_8297,N_8149,N_8032);
or U8298 (N_8298,N_8161,N_8020);
nor U8299 (N_8299,N_8084,N_8043);
nand U8300 (N_8300,N_8150,N_8148);
xor U8301 (N_8301,N_8047,N_8184);
nor U8302 (N_8302,N_8026,N_8183);
nor U8303 (N_8303,N_8135,N_8165);
or U8304 (N_8304,N_8172,N_8031);
and U8305 (N_8305,N_8071,N_8023);
or U8306 (N_8306,N_8189,N_8054);
or U8307 (N_8307,N_8073,N_8027);
or U8308 (N_8308,N_8198,N_8011);
or U8309 (N_8309,N_8051,N_8083);
xnor U8310 (N_8310,N_8198,N_8154);
and U8311 (N_8311,N_8184,N_8137);
or U8312 (N_8312,N_8061,N_8093);
and U8313 (N_8313,N_8089,N_8083);
xor U8314 (N_8314,N_8012,N_8125);
nor U8315 (N_8315,N_8106,N_8176);
or U8316 (N_8316,N_8133,N_8045);
xnor U8317 (N_8317,N_8045,N_8162);
xnor U8318 (N_8318,N_8052,N_8033);
nand U8319 (N_8319,N_8045,N_8063);
xnor U8320 (N_8320,N_8098,N_8081);
nor U8321 (N_8321,N_8013,N_8180);
or U8322 (N_8322,N_8012,N_8194);
and U8323 (N_8323,N_8129,N_8000);
xnor U8324 (N_8324,N_8085,N_8119);
nand U8325 (N_8325,N_8109,N_8070);
and U8326 (N_8326,N_8175,N_8015);
or U8327 (N_8327,N_8104,N_8073);
and U8328 (N_8328,N_8063,N_8071);
nor U8329 (N_8329,N_8047,N_8125);
nor U8330 (N_8330,N_8046,N_8097);
nor U8331 (N_8331,N_8113,N_8199);
or U8332 (N_8332,N_8062,N_8120);
nor U8333 (N_8333,N_8032,N_8006);
or U8334 (N_8334,N_8140,N_8020);
xor U8335 (N_8335,N_8004,N_8031);
nand U8336 (N_8336,N_8151,N_8012);
nand U8337 (N_8337,N_8042,N_8077);
xor U8338 (N_8338,N_8028,N_8100);
xnor U8339 (N_8339,N_8088,N_8076);
nor U8340 (N_8340,N_8177,N_8153);
and U8341 (N_8341,N_8178,N_8049);
and U8342 (N_8342,N_8180,N_8189);
xnor U8343 (N_8343,N_8077,N_8006);
nand U8344 (N_8344,N_8087,N_8182);
nor U8345 (N_8345,N_8016,N_8144);
nor U8346 (N_8346,N_8017,N_8096);
nor U8347 (N_8347,N_8055,N_8184);
or U8348 (N_8348,N_8098,N_8064);
or U8349 (N_8349,N_8173,N_8084);
xnor U8350 (N_8350,N_8116,N_8104);
nand U8351 (N_8351,N_8164,N_8137);
nand U8352 (N_8352,N_8050,N_8081);
xor U8353 (N_8353,N_8010,N_8194);
xnor U8354 (N_8354,N_8026,N_8140);
or U8355 (N_8355,N_8025,N_8127);
and U8356 (N_8356,N_8156,N_8145);
nand U8357 (N_8357,N_8175,N_8131);
nor U8358 (N_8358,N_8117,N_8018);
or U8359 (N_8359,N_8092,N_8077);
xnor U8360 (N_8360,N_8072,N_8190);
and U8361 (N_8361,N_8157,N_8085);
and U8362 (N_8362,N_8007,N_8109);
nand U8363 (N_8363,N_8105,N_8156);
nand U8364 (N_8364,N_8127,N_8027);
nand U8365 (N_8365,N_8104,N_8153);
or U8366 (N_8366,N_8060,N_8093);
or U8367 (N_8367,N_8055,N_8043);
or U8368 (N_8368,N_8093,N_8184);
nor U8369 (N_8369,N_8042,N_8103);
xnor U8370 (N_8370,N_8073,N_8029);
xor U8371 (N_8371,N_8145,N_8043);
and U8372 (N_8372,N_8172,N_8089);
or U8373 (N_8373,N_8077,N_8103);
and U8374 (N_8374,N_8021,N_8105);
or U8375 (N_8375,N_8027,N_8056);
or U8376 (N_8376,N_8087,N_8050);
xor U8377 (N_8377,N_8094,N_8009);
or U8378 (N_8378,N_8152,N_8178);
xnor U8379 (N_8379,N_8056,N_8005);
nor U8380 (N_8380,N_8078,N_8027);
or U8381 (N_8381,N_8110,N_8154);
nand U8382 (N_8382,N_8067,N_8060);
nor U8383 (N_8383,N_8081,N_8095);
or U8384 (N_8384,N_8177,N_8023);
nor U8385 (N_8385,N_8160,N_8045);
xnor U8386 (N_8386,N_8012,N_8174);
nand U8387 (N_8387,N_8106,N_8123);
nor U8388 (N_8388,N_8184,N_8141);
or U8389 (N_8389,N_8191,N_8147);
and U8390 (N_8390,N_8009,N_8000);
nand U8391 (N_8391,N_8004,N_8190);
nor U8392 (N_8392,N_8053,N_8124);
nand U8393 (N_8393,N_8129,N_8089);
nor U8394 (N_8394,N_8136,N_8187);
or U8395 (N_8395,N_8068,N_8159);
nand U8396 (N_8396,N_8013,N_8000);
or U8397 (N_8397,N_8111,N_8070);
xor U8398 (N_8398,N_8174,N_8167);
or U8399 (N_8399,N_8194,N_8028);
nand U8400 (N_8400,N_8252,N_8243);
or U8401 (N_8401,N_8387,N_8211);
or U8402 (N_8402,N_8307,N_8316);
nor U8403 (N_8403,N_8291,N_8204);
or U8404 (N_8404,N_8358,N_8258);
or U8405 (N_8405,N_8317,N_8288);
nand U8406 (N_8406,N_8384,N_8236);
xnor U8407 (N_8407,N_8260,N_8386);
xnor U8408 (N_8408,N_8293,N_8329);
nand U8409 (N_8409,N_8349,N_8247);
or U8410 (N_8410,N_8360,N_8231);
xor U8411 (N_8411,N_8245,N_8394);
nand U8412 (N_8412,N_8265,N_8327);
xnor U8413 (N_8413,N_8262,N_8356);
or U8414 (N_8414,N_8223,N_8216);
nand U8415 (N_8415,N_8226,N_8283);
xor U8416 (N_8416,N_8361,N_8346);
xor U8417 (N_8417,N_8290,N_8220);
xnor U8418 (N_8418,N_8210,N_8305);
and U8419 (N_8419,N_8287,N_8397);
nand U8420 (N_8420,N_8271,N_8319);
nor U8421 (N_8421,N_8202,N_8269);
xor U8422 (N_8422,N_8344,N_8389);
or U8423 (N_8423,N_8294,N_8310);
or U8424 (N_8424,N_8372,N_8328);
nor U8425 (N_8425,N_8280,N_8311);
xnor U8426 (N_8426,N_8337,N_8266);
or U8427 (N_8427,N_8276,N_8268);
and U8428 (N_8428,N_8371,N_8335);
and U8429 (N_8429,N_8278,N_8395);
nand U8430 (N_8430,N_8214,N_8302);
nand U8431 (N_8431,N_8295,N_8355);
or U8432 (N_8432,N_8345,N_8208);
and U8433 (N_8433,N_8366,N_8264);
nor U8434 (N_8434,N_8279,N_8312);
xor U8435 (N_8435,N_8359,N_8378);
xor U8436 (N_8436,N_8207,N_8332);
xor U8437 (N_8437,N_8205,N_8336);
nand U8438 (N_8438,N_8370,N_8323);
nand U8439 (N_8439,N_8342,N_8314);
xor U8440 (N_8440,N_8206,N_8354);
or U8441 (N_8441,N_8390,N_8351);
xor U8442 (N_8442,N_8289,N_8224);
and U8443 (N_8443,N_8261,N_8237);
xnor U8444 (N_8444,N_8241,N_8242);
and U8445 (N_8445,N_8256,N_8201);
nor U8446 (N_8446,N_8347,N_8249);
or U8447 (N_8447,N_8213,N_8304);
and U8448 (N_8448,N_8298,N_8246);
nor U8449 (N_8449,N_8200,N_8373);
xor U8450 (N_8450,N_8353,N_8218);
xnor U8451 (N_8451,N_8250,N_8257);
nor U8452 (N_8452,N_8240,N_8393);
nor U8453 (N_8453,N_8263,N_8296);
xor U8454 (N_8454,N_8340,N_8374);
or U8455 (N_8455,N_8318,N_8232);
and U8456 (N_8456,N_8273,N_8322);
nor U8457 (N_8457,N_8320,N_8251);
or U8458 (N_8458,N_8338,N_8282);
xor U8459 (N_8459,N_8274,N_8308);
and U8460 (N_8460,N_8334,N_8253);
nand U8461 (N_8461,N_8248,N_8297);
and U8462 (N_8462,N_8330,N_8350);
or U8463 (N_8463,N_8300,N_8235);
xnor U8464 (N_8464,N_8369,N_8333);
xnor U8465 (N_8465,N_8233,N_8238);
xnor U8466 (N_8466,N_8267,N_8391);
xnor U8467 (N_8467,N_8382,N_8331);
nor U8468 (N_8468,N_8315,N_8244);
xnor U8469 (N_8469,N_8234,N_8217);
xnor U8470 (N_8470,N_8277,N_8396);
nand U8471 (N_8471,N_8381,N_8368);
nand U8472 (N_8472,N_8286,N_8398);
and U8473 (N_8473,N_8309,N_8301);
and U8474 (N_8474,N_8367,N_8219);
xnor U8475 (N_8475,N_8376,N_8399);
nor U8476 (N_8476,N_8324,N_8341);
and U8477 (N_8477,N_8222,N_8380);
or U8478 (N_8478,N_8348,N_8228);
nor U8479 (N_8479,N_8270,N_8385);
xor U8480 (N_8480,N_8362,N_8225);
xnor U8481 (N_8481,N_8255,N_8203);
and U8482 (N_8482,N_8227,N_8221);
nand U8483 (N_8483,N_8306,N_8379);
xnor U8484 (N_8484,N_8313,N_8212);
or U8485 (N_8485,N_8339,N_8365);
or U8486 (N_8486,N_8209,N_8352);
nor U8487 (N_8487,N_8254,N_8229);
and U8488 (N_8488,N_8357,N_8292);
and U8489 (N_8489,N_8215,N_8281);
or U8490 (N_8490,N_8272,N_8375);
xnor U8491 (N_8491,N_8363,N_8285);
xor U8492 (N_8492,N_8377,N_8383);
nand U8493 (N_8493,N_8388,N_8275);
or U8494 (N_8494,N_8326,N_8303);
xor U8495 (N_8495,N_8230,N_8364);
nor U8496 (N_8496,N_8299,N_8321);
nor U8497 (N_8497,N_8392,N_8325);
or U8498 (N_8498,N_8259,N_8343);
or U8499 (N_8499,N_8239,N_8284);
xnor U8500 (N_8500,N_8305,N_8283);
nand U8501 (N_8501,N_8350,N_8378);
and U8502 (N_8502,N_8247,N_8269);
nand U8503 (N_8503,N_8394,N_8234);
nand U8504 (N_8504,N_8382,N_8375);
nand U8505 (N_8505,N_8254,N_8328);
or U8506 (N_8506,N_8262,N_8359);
and U8507 (N_8507,N_8348,N_8245);
nor U8508 (N_8508,N_8330,N_8341);
or U8509 (N_8509,N_8334,N_8257);
nand U8510 (N_8510,N_8309,N_8300);
nand U8511 (N_8511,N_8263,N_8349);
nor U8512 (N_8512,N_8261,N_8294);
nand U8513 (N_8513,N_8329,N_8388);
xor U8514 (N_8514,N_8276,N_8298);
xnor U8515 (N_8515,N_8380,N_8363);
or U8516 (N_8516,N_8335,N_8326);
nand U8517 (N_8517,N_8313,N_8392);
xnor U8518 (N_8518,N_8292,N_8203);
and U8519 (N_8519,N_8321,N_8288);
nand U8520 (N_8520,N_8229,N_8316);
xnor U8521 (N_8521,N_8355,N_8212);
xnor U8522 (N_8522,N_8392,N_8331);
nor U8523 (N_8523,N_8204,N_8255);
or U8524 (N_8524,N_8232,N_8335);
or U8525 (N_8525,N_8349,N_8364);
or U8526 (N_8526,N_8240,N_8380);
nor U8527 (N_8527,N_8393,N_8243);
nor U8528 (N_8528,N_8264,N_8393);
nand U8529 (N_8529,N_8294,N_8239);
nor U8530 (N_8530,N_8292,N_8375);
nor U8531 (N_8531,N_8372,N_8319);
and U8532 (N_8532,N_8234,N_8360);
xor U8533 (N_8533,N_8268,N_8381);
and U8534 (N_8534,N_8350,N_8292);
nand U8535 (N_8535,N_8284,N_8318);
nor U8536 (N_8536,N_8331,N_8239);
nor U8537 (N_8537,N_8239,N_8299);
xor U8538 (N_8538,N_8249,N_8332);
xor U8539 (N_8539,N_8367,N_8212);
xnor U8540 (N_8540,N_8360,N_8311);
nand U8541 (N_8541,N_8353,N_8389);
nor U8542 (N_8542,N_8311,N_8316);
or U8543 (N_8543,N_8332,N_8299);
and U8544 (N_8544,N_8382,N_8380);
or U8545 (N_8545,N_8357,N_8240);
and U8546 (N_8546,N_8374,N_8254);
or U8547 (N_8547,N_8332,N_8252);
nor U8548 (N_8548,N_8347,N_8354);
and U8549 (N_8549,N_8263,N_8271);
nor U8550 (N_8550,N_8388,N_8246);
xor U8551 (N_8551,N_8227,N_8288);
nor U8552 (N_8552,N_8223,N_8328);
and U8553 (N_8553,N_8334,N_8370);
or U8554 (N_8554,N_8349,N_8254);
nand U8555 (N_8555,N_8279,N_8366);
nor U8556 (N_8556,N_8240,N_8353);
nand U8557 (N_8557,N_8322,N_8356);
nand U8558 (N_8558,N_8339,N_8222);
xnor U8559 (N_8559,N_8222,N_8351);
and U8560 (N_8560,N_8297,N_8353);
xor U8561 (N_8561,N_8228,N_8350);
and U8562 (N_8562,N_8235,N_8308);
nor U8563 (N_8563,N_8221,N_8327);
and U8564 (N_8564,N_8341,N_8334);
nand U8565 (N_8565,N_8291,N_8343);
xnor U8566 (N_8566,N_8214,N_8284);
xnor U8567 (N_8567,N_8237,N_8238);
xnor U8568 (N_8568,N_8314,N_8256);
nor U8569 (N_8569,N_8335,N_8353);
xnor U8570 (N_8570,N_8238,N_8243);
and U8571 (N_8571,N_8280,N_8390);
and U8572 (N_8572,N_8259,N_8287);
nor U8573 (N_8573,N_8383,N_8316);
or U8574 (N_8574,N_8342,N_8343);
xor U8575 (N_8575,N_8284,N_8268);
or U8576 (N_8576,N_8356,N_8215);
nor U8577 (N_8577,N_8386,N_8314);
nand U8578 (N_8578,N_8346,N_8347);
and U8579 (N_8579,N_8301,N_8211);
nand U8580 (N_8580,N_8327,N_8333);
and U8581 (N_8581,N_8325,N_8236);
nor U8582 (N_8582,N_8204,N_8327);
or U8583 (N_8583,N_8328,N_8330);
nor U8584 (N_8584,N_8343,N_8356);
nand U8585 (N_8585,N_8248,N_8295);
and U8586 (N_8586,N_8290,N_8259);
xnor U8587 (N_8587,N_8313,N_8329);
xor U8588 (N_8588,N_8271,N_8292);
nand U8589 (N_8589,N_8260,N_8257);
nand U8590 (N_8590,N_8355,N_8305);
and U8591 (N_8591,N_8321,N_8357);
nor U8592 (N_8592,N_8281,N_8302);
or U8593 (N_8593,N_8316,N_8300);
and U8594 (N_8594,N_8294,N_8235);
nor U8595 (N_8595,N_8322,N_8323);
or U8596 (N_8596,N_8218,N_8246);
and U8597 (N_8597,N_8377,N_8228);
nor U8598 (N_8598,N_8235,N_8345);
nand U8599 (N_8599,N_8283,N_8327);
nor U8600 (N_8600,N_8506,N_8492);
nor U8601 (N_8601,N_8471,N_8554);
xnor U8602 (N_8602,N_8484,N_8587);
xnor U8603 (N_8603,N_8421,N_8453);
xor U8604 (N_8604,N_8488,N_8594);
nor U8605 (N_8605,N_8412,N_8577);
nand U8606 (N_8606,N_8517,N_8450);
xnor U8607 (N_8607,N_8504,N_8520);
or U8608 (N_8608,N_8496,N_8523);
nand U8609 (N_8609,N_8475,N_8596);
nand U8610 (N_8610,N_8536,N_8442);
and U8611 (N_8611,N_8581,N_8550);
nor U8612 (N_8612,N_8534,N_8485);
nand U8613 (N_8613,N_8527,N_8589);
xor U8614 (N_8614,N_8528,N_8410);
and U8615 (N_8615,N_8538,N_8586);
xnor U8616 (N_8616,N_8499,N_8495);
xnor U8617 (N_8617,N_8459,N_8533);
nand U8618 (N_8618,N_8415,N_8432);
xor U8619 (N_8619,N_8401,N_8447);
and U8620 (N_8620,N_8456,N_8526);
nand U8621 (N_8621,N_8402,N_8487);
nor U8622 (N_8622,N_8409,N_8505);
and U8623 (N_8623,N_8564,N_8451);
and U8624 (N_8624,N_8572,N_8503);
and U8625 (N_8625,N_8413,N_8478);
or U8626 (N_8626,N_8429,N_8498);
or U8627 (N_8627,N_8420,N_8437);
xor U8628 (N_8628,N_8474,N_8560);
xor U8629 (N_8629,N_8508,N_8515);
nor U8630 (N_8630,N_8552,N_8571);
or U8631 (N_8631,N_8406,N_8425);
nand U8632 (N_8632,N_8449,N_8501);
xnor U8633 (N_8633,N_8584,N_8466);
xor U8634 (N_8634,N_8513,N_8588);
nand U8635 (N_8635,N_8422,N_8592);
nor U8636 (N_8636,N_8486,N_8511);
nor U8637 (N_8637,N_8482,N_8463);
xor U8638 (N_8638,N_8477,N_8404);
nor U8639 (N_8639,N_8539,N_8431);
or U8640 (N_8640,N_8507,N_8483);
or U8641 (N_8641,N_8597,N_8419);
nor U8642 (N_8642,N_8512,N_8480);
nand U8643 (N_8643,N_8531,N_8553);
xor U8644 (N_8644,N_8446,N_8583);
nor U8645 (N_8645,N_8433,N_8591);
xnor U8646 (N_8646,N_8549,N_8545);
nand U8647 (N_8647,N_8445,N_8521);
or U8648 (N_8648,N_8519,N_8590);
nor U8649 (N_8649,N_8541,N_8489);
xnor U8650 (N_8650,N_8472,N_8473);
xnor U8651 (N_8651,N_8563,N_8535);
and U8652 (N_8652,N_8467,N_8479);
or U8653 (N_8653,N_8497,N_8557);
or U8654 (N_8654,N_8522,N_8529);
or U8655 (N_8655,N_8408,N_8524);
or U8656 (N_8656,N_8417,N_8491);
or U8657 (N_8657,N_8414,N_8430);
nor U8658 (N_8658,N_8565,N_8464);
xor U8659 (N_8659,N_8540,N_8510);
xor U8660 (N_8660,N_8578,N_8407);
nand U8661 (N_8661,N_8559,N_8490);
or U8662 (N_8662,N_8461,N_8427);
nand U8663 (N_8663,N_8502,N_8454);
nor U8664 (N_8664,N_8562,N_8434);
nand U8665 (N_8665,N_8476,N_8544);
or U8666 (N_8666,N_8457,N_8452);
and U8667 (N_8667,N_8558,N_8569);
or U8668 (N_8668,N_8403,N_8424);
xnor U8669 (N_8669,N_8530,N_8469);
nand U8670 (N_8670,N_8460,N_8426);
nand U8671 (N_8671,N_8428,N_8574);
and U8672 (N_8672,N_8551,N_8448);
xnor U8673 (N_8673,N_8455,N_8547);
xor U8674 (N_8674,N_8438,N_8543);
nand U8675 (N_8675,N_8444,N_8436);
or U8676 (N_8676,N_8575,N_8400);
and U8677 (N_8677,N_8570,N_8439);
nand U8678 (N_8678,N_8405,N_8500);
and U8679 (N_8679,N_8418,N_8542);
xor U8680 (N_8680,N_8441,N_8567);
and U8681 (N_8681,N_8423,N_8585);
nor U8682 (N_8682,N_8537,N_8579);
xnor U8683 (N_8683,N_8555,N_8525);
xor U8684 (N_8684,N_8599,N_8493);
nand U8685 (N_8685,N_8416,N_8561);
or U8686 (N_8686,N_8516,N_8576);
xor U8687 (N_8687,N_8548,N_8481);
and U8688 (N_8688,N_8593,N_8514);
xnor U8689 (N_8689,N_8518,N_8595);
and U8690 (N_8690,N_8411,N_8598);
nor U8691 (N_8691,N_8462,N_8468);
xnor U8692 (N_8692,N_8440,N_8546);
and U8693 (N_8693,N_8465,N_8556);
or U8694 (N_8694,N_8582,N_8568);
and U8695 (N_8695,N_8580,N_8443);
or U8696 (N_8696,N_8509,N_8532);
or U8697 (N_8697,N_8435,N_8470);
and U8698 (N_8698,N_8573,N_8458);
nor U8699 (N_8699,N_8566,N_8494);
nand U8700 (N_8700,N_8596,N_8496);
nor U8701 (N_8701,N_8539,N_8453);
nand U8702 (N_8702,N_8490,N_8554);
and U8703 (N_8703,N_8546,N_8583);
nor U8704 (N_8704,N_8483,N_8564);
nand U8705 (N_8705,N_8526,N_8548);
nand U8706 (N_8706,N_8434,N_8436);
xnor U8707 (N_8707,N_8418,N_8558);
nor U8708 (N_8708,N_8406,N_8458);
xnor U8709 (N_8709,N_8581,N_8574);
nor U8710 (N_8710,N_8589,N_8486);
and U8711 (N_8711,N_8515,N_8597);
nand U8712 (N_8712,N_8439,N_8470);
nor U8713 (N_8713,N_8483,N_8419);
nor U8714 (N_8714,N_8574,N_8544);
nor U8715 (N_8715,N_8475,N_8400);
or U8716 (N_8716,N_8430,N_8504);
nor U8717 (N_8717,N_8422,N_8575);
nand U8718 (N_8718,N_8597,N_8530);
nor U8719 (N_8719,N_8516,N_8555);
and U8720 (N_8720,N_8510,N_8526);
nor U8721 (N_8721,N_8442,N_8403);
nor U8722 (N_8722,N_8595,N_8409);
nand U8723 (N_8723,N_8537,N_8464);
xor U8724 (N_8724,N_8572,N_8435);
and U8725 (N_8725,N_8580,N_8452);
and U8726 (N_8726,N_8421,N_8493);
and U8727 (N_8727,N_8516,N_8433);
or U8728 (N_8728,N_8457,N_8486);
nor U8729 (N_8729,N_8499,N_8567);
or U8730 (N_8730,N_8543,N_8545);
nand U8731 (N_8731,N_8436,N_8428);
and U8732 (N_8732,N_8432,N_8569);
or U8733 (N_8733,N_8497,N_8411);
nor U8734 (N_8734,N_8425,N_8585);
and U8735 (N_8735,N_8452,N_8426);
and U8736 (N_8736,N_8555,N_8496);
xor U8737 (N_8737,N_8420,N_8539);
and U8738 (N_8738,N_8463,N_8508);
nand U8739 (N_8739,N_8438,N_8468);
nand U8740 (N_8740,N_8426,N_8582);
or U8741 (N_8741,N_8573,N_8464);
nor U8742 (N_8742,N_8544,N_8502);
xor U8743 (N_8743,N_8466,N_8458);
xnor U8744 (N_8744,N_8460,N_8404);
nor U8745 (N_8745,N_8505,N_8444);
nand U8746 (N_8746,N_8423,N_8533);
nand U8747 (N_8747,N_8456,N_8477);
nand U8748 (N_8748,N_8508,N_8493);
xnor U8749 (N_8749,N_8407,N_8446);
nand U8750 (N_8750,N_8465,N_8426);
nor U8751 (N_8751,N_8465,N_8511);
xor U8752 (N_8752,N_8452,N_8444);
and U8753 (N_8753,N_8407,N_8484);
nand U8754 (N_8754,N_8467,N_8468);
or U8755 (N_8755,N_8457,N_8560);
xnor U8756 (N_8756,N_8553,N_8439);
nand U8757 (N_8757,N_8549,N_8538);
nand U8758 (N_8758,N_8489,N_8578);
or U8759 (N_8759,N_8494,N_8577);
and U8760 (N_8760,N_8528,N_8492);
or U8761 (N_8761,N_8582,N_8476);
nor U8762 (N_8762,N_8432,N_8436);
or U8763 (N_8763,N_8503,N_8531);
xnor U8764 (N_8764,N_8577,N_8482);
xor U8765 (N_8765,N_8502,N_8514);
nand U8766 (N_8766,N_8478,N_8450);
nand U8767 (N_8767,N_8452,N_8480);
nand U8768 (N_8768,N_8431,N_8403);
and U8769 (N_8769,N_8440,N_8411);
or U8770 (N_8770,N_8419,N_8530);
and U8771 (N_8771,N_8463,N_8481);
nand U8772 (N_8772,N_8439,N_8456);
xnor U8773 (N_8773,N_8553,N_8468);
nand U8774 (N_8774,N_8568,N_8525);
nand U8775 (N_8775,N_8559,N_8472);
nor U8776 (N_8776,N_8575,N_8562);
xor U8777 (N_8777,N_8403,N_8438);
and U8778 (N_8778,N_8496,N_8504);
or U8779 (N_8779,N_8521,N_8546);
or U8780 (N_8780,N_8436,N_8484);
nand U8781 (N_8781,N_8501,N_8537);
nand U8782 (N_8782,N_8484,N_8435);
and U8783 (N_8783,N_8535,N_8430);
or U8784 (N_8784,N_8589,N_8485);
nor U8785 (N_8785,N_8535,N_8412);
and U8786 (N_8786,N_8543,N_8526);
nor U8787 (N_8787,N_8481,N_8452);
or U8788 (N_8788,N_8584,N_8498);
or U8789 (N_8789,N_8517,N_8547);
xnor U8790 (N_8790,N_8431,N_8463);
xor U8791 (N_8791,N_8507,N_8574);
xor U8792 (N_8792,N_8569,N_8544);
xnor U8793 (N_8793,N_8439,N_8517);
or U8794 (N_8794,N_8496,N_8475);
nor U8795 (N_8795,N_8517,N_8525);
nand U8796 (N_8796,N_8541,N_8495);
xor U8797 (N_8797,N_8452,N_8532);
nor U8798 (N_8798,N_8536,N_8437);
and U8799 (N_8799,N_8474,N_8465);
and U8800 (N_8800,N_8695,N_8643);
xor U8801 (N_8801,N_8783,N_8715);
nand U8802 (N_8802,N_8778,N_8762);
or U8803 (N_8803,N_8752,N_8750);
or U8804 (N_8804,N_8768,N_8686);
and U8805 (N_8805,N_8667,N_8646);
or U8806 (N_8806,N_8690,N_8781);
or U8807 (N_8807,N_8617,N_8700);
xnor U8808 (N_8808,N_8738,N_8613);
xnor U8809 (N_8809,N_8641,N_8632);
or U8810 (N_8810,N_8602,N_8611);
or U8811 (N_8811,N_8769,N_8731);
or U8812 (N_8812,N_8794,N_8694);
xnor U8813 (N_8813,N_8718,N_8619);
or U8814 (N_8814,N_8708,N_8607);
nand U8815 (N_8815,N_8721,N_8797);
nand U8816 (N_8816,N_8622,N_8691);
or U8817 (N_8817,N_8680,N_8633);
or U8818 (N_8818,N_8628,N_8751);
xnor U8819 (N_8819,N_8760,N_8705);
xnor U8820 (N_8820,N_8712,N_8669);
or U8821 (N_8821,N_8727,N_8744);
nor U8822 (N_8822,N_8767,N_8650);
or U8823 (N_8823,N_8652,N_8735);
nor U8824 (N_8824,N_8638,N_8782);
nand U8825 (N_8825,N_8687,N_8625);
xor U8826 (N_8826,N_8726,N_8629);
nand U8827 (N_8827,N_8671,N_8634);
or U8828 (N_8828,N_8739,N_8615);
or U8829 (N_8829,N_8713,N_8761);
nand U8830 (N_8830,N_8606,N_8716);
xor U8831 (N_8831,N_8720,N_8658);
nand U8832 (N_8832,N_8732,N_8645);
nand U8833 (N_8833,N_8709,N_8688);
nor U8834 (N_8834,N_8777,N_8668);
or U8835 (N_8835,N_8722,N_8730);
and U8836 (N_8836,N_8770,N_8765);
xor U8837 (N_8837,N_8636,N_8654);
nand U8838 (N_8838,N_8746,N_8614);
or U8839 (N_8839,N_8662,N_8626);
and U8840 (N_8840,N_8784,N_8683);
xor U8841 (N_8841,N_8648,N_8754);
nand U8842 (N_8842,N_8651,N_8789);
nand U8843 (N_8843,N_8659,N_8656);
and U8844 (N_8844,N_8773,N_8657);
xor U8845 (N_8845,N_8664,N_8681);
nand U8846 (N_8846,N_8791,N_8729);
nand U8847 (N_8847,N_8660,N_8758);
nor U8848 (N_8848,N_8759,N_8601);
or U8849 (N_8849,N_8665,N_8792);
nand U8850 (N_8850,N_8741,N_8655);
or U8851 (N_8851,N_8749,N_8623);
and U8852 (N_8852,N_8701,N_8679);
or U8853 (N_8853,N_8685,N_8637);
and U8854 (N_8854,N_8764,N_8745);
nand U8855 (N_8855,N_8644,N_8672);
nand U8856 (N_8856,N_8639,N_8677);
xnor U8857 (N_8857,N_8661,N_8698);
nand U8858 (N_8858,N_8719,N_8670);
or U8859 (N_8859,N_8799,N_8734);
xnor U8860 (N_8860,N_8728,N_8620);
and U8861 (N_8861,N_8717,N_8774);
and U8862 (N_8862,N_8640,N_8616);
nand U8863 (N_8863,N_8725,N_8630);
nand U8864 (N_8864,N_8772,N_8674);
nand U8865 (N_8865,N_8743,N_8787);
nand U8866 (N_8866,N_8706,N_8723);
xnor U8867 (N_8867,N_8740,N_8757);
nor U8868 (N_8868,N_8699,N_8684);
xnor U8869 (N_8869,N_8714,N_8631);
nor U8870 (N_8870,N_8747,N_8775);
nand U8871 (N_8871,N_8600,N_8692);
or U8872 (N_8872,N_8793,N_8702);
xnor U8873 (N_8873,N_8693,N_8682);
nand U8874 (N_8874,N_8627,N_8755);
xnor U8875 (N_8875,N_8618,N_8642);
or U8876 (N_8876,N_8624,N_8776);
nor U8877 (N_8877,N_8647,N_8663);
and U8878 (N_8878,N_8710,N_8704);
nand U8879 (N_8879,N_8678,N_8610);
nor U8880 (N_8880,N_8753,N_8796);
nor U8881 (N_8881,N_8711,N_8766);
or U8882 (N_8882,N_8603,N_8635);
xnor U8883 (N_8883,N_8798,N_8795);
xor U8884 (N_8884,N_8608,N_8707);
and U8885 (N_8885,N_8786,N_8621);
or U8886 (N_8886,N_8748,N_8780);
and U8887 (N_8887,N_8779,N_8666);
xor U8888 (N_8888,N_8689,N_8612);
nor U8889 (N_8889,N_8697,N_8771);
and U8890 (N_8890,N_8609,N_8724);
nor U8891 (N_8891,N_8653,N_8676);
nand U8892 (N_8892,N_8605,N_8696);
nor U8893 (N_8893,N_8756,N_8649);
nor U8894 (N_8894,N_8763,N_8785);
and U8895 (N_8895,N_8673,N_8703);
and U8896 (N_8896,N_8733,N_8604);
or U8897 (N_8897,N_8788,N_8737);
nand U8898 (N_8898,N_8736,N_8742);
and U8899 (N_8899,N_8675,N_8790);
or U8900 (N_8900,N_8734,N_8657);
or U8901 (N_8901,N_8683,N_8760);
nand U8902 (N_8902,N_8733,N_8700);
nand U8903 (N_8903,N_8775,N_8720);
and U8904 (N_8904,N_8731,N_8789);
nand U8905 (N_8905,N_8639,N_8711);
and U8906 (N_8906,N_8616,N_8746);
xor U8907 (N_8907,N_8606,N_8727);
nor U8908 (N_8908,N_8609,N_8680);
or U8909 (N_8909,N_8796,N_8710);
nor U8910 (N_8910,N_8651,N_8795);
xnor U8911 (N_8911,N_8794,N_8671);
and U8912 (N_8912,N_8732,N_8622);
and U8913 (N_8913,N_8645,N_8633);
or U8914 (N_8914,N_8717,N_8631);
or U8915 (N_8915,N_8740,N_8673);
nor U8916 (N_8916,N_8681,N_8661);
xnor U8917 (N_8917,N_8688,N_8652);
nand U8918 (N_8918,N_8735,N_8695);
nand U8919 (N_8919,N_8717,N_8719);
and U8920 (N_8920,N_8731,N_8636);
nand U8921 (N_8921,N_8618,N_8689);
or U8922 (N_8922,N_8675,N_8647);
nor U8923 (N_8923,N_8629,N_8785);
nor U8924 (N_8924,N_8731,N_8691);
nor U8925 (N_8925,N_8739,N_8783);
or U8926 (N_8926,N_8744,N_8693);
or U8927 (N_8927,N_8753,N_8604);
or U8928 (N_8928,N_8796,N_8717);
nand U8929 (N_8929,N_8792,N_8722);
nor U8930 (N_8930,N_8606,N_8712);
xor U8931 (N_8931,N_8753,N_8650);
nand U8932 (N_8932,N_8709,N_8721);
nor U8933 (N_8933,N_8621,N_8713);
nand U8934 (N_8934,N_8612,N_8728);
nor U8935 (N_8935,N_8694,N_8666);
or U8936 (N_8936,N_8662,N_8770);
nor U8937 (N_8937,N_8794,N_8735);
nor U8938 (N_8938,N_8618,N_8747);
and U8939 (N_8939,N_8629,N_8671);
and U8940 (N_8940,N_8794,N_8624);
or U8941 (N_8941,N_8703,N_8612);
nor U8942 (N_8942,N_8674,N_8646);
and U8943 (N_8943,N_8706,N_8695);
xor U8944 (N_8944,N_8672,N_8641);
and U8945 (N_8945,N_8780,N_8643);
xor U8946 (N_8946,N_8611,N_8698);
or U8947 (N_8947,N_8683,N_8633);
xnor U8948 (N_8948,N_8740,N_8762);
nor U8949 (N_8949,N_8750,N_8669);
xnor U8950 (N_8950,N_8746,N_8627);
nor U8951 (N_8951,N_8721,N_8696);
and U8952 (N_8952,N_8720,N_8714);
xor U8953 (N_8953,N_8623,N_8637);
xnor U8954 (N_8954,N_8660,N_8712);
nand U8955 (N_8955,N_8662,N_8601);
and U8956 (N_8956,N_8626,N_8669);
xor U8957 (N_8957,N_8649,N_8786);
nand U8958 (N_8958,N_8603,N_8767);
xnor U8959 (N_8959,N_8738,N_8774);
nand U8960 (N_8960,N_8648,N_8772);
nand U8961 (N_8961,N_8624,N_8664);
and U8962 (N_8962,N_8694,N_8745);
nor U8963 (N_8963,N_8732,N_8650);
and U8964 (N_8964,N_8613,N_8785);
nor U8965 (N_8965,N_8799,N_8602);
or U8966 (N_8966,N_8719,N_8783);
and U8967 (N_8967,N_8668,N_8680);
nand U8968 (N_8968,N_8671,N_8725);
nand U8969 (N_8969,N_8754,N_8763);
nand U8970 (N_8970,N_8624,N_8798);
nor U8971 (N_8971,N_8717,N_8753);
or U8972 (N_8972,N_8777,N_8771);
and U8973 (N_8973,N_8740,N_8746);
or U8974 (N_8974,N_8713,N_8625);
xnor U8975 (N_8975,N_8784,N_8778);
nor U8976 (N_8976,N_8683,N_8607);
or U8977 (N_8977,N_8762,N_8728);
xnor U8978 (N_8978,N_8609,N_8702);
nor U8979 (N_8979,N_8772,N_8612);
xor U8980 (N_8980,N_8775,N_8622);
xor U8981 (N_8981,N_8645,N_8739);
and U8982 (N_8982,N_8768,N_8607);
nor U8983 (N_8983,N_8758,N_8751);
and U8984 (N_8984,N_8748,N_8711);
and U8985 (N_8985,N_8691,N_8770);
nand U8986 (N_8986,N_8704,N_8772);
or U8987 (N_8987,N_8738,N_8667);
nor U8988 (N_8988,N_8631,N_8735);
or U8989 (N_8989,N_8637,N_8746);
and U8990 (N_8990,N_8768,N_8795);
or U8991 (N_8991,N_8717,N_8775);
xnor U8992 (N_8992,N_8652,N_8619);
xor U8993 (N_8993,N_8694,N_8612);
or U8994 (N_8994,N_8784,N_8744);
xor U8995 (N_8995,N_8629,N_8653);
nand U8996 (N_8996,N_8740,N_8695);
or U8997 (N_8997,N_8713,N_8724);
nand U8998 (N_8998,N_8738,N_8610);
nand U8999 (N_8999,N_8712,N_8725);
xor U9000 (N_9000,N_8910,N_8868);
xnor U9001 (N_9001,N_8887,N_8993);
and U9002 (N_9002,N_8804,N_8862);
and U9003 (N_9003,N_8809,N_8982);
nand U9004 (N_9004,N_8896,N_8866);
nor U9005 (N_9005,N_8874,N_8994);
xor U9006 (N_9006,N_8856,N_8955);
and U9007 (N_9007,N_8941,N_8976);
xnor U9008 (N_9008,N_8915,N_8840);
nor U9009 (N_9009,N_8966,N_8892);
nand U9010 (N_9010,N_8968,N_8995);
nor U9011 (N_9011,N_8942,N_8878);
xnor U9012 (N_9012,N_8872,N_8836);
or U9013 (N_9013,N_8815,N_8826);
nand U9014 (N_9014,N_8842,N_8914);
nand U9015 (N_9015,N_8947,N_8900);
or U9016 (N_9016,N_8933,N_8908);
nand U9017 (N_9017,N_8898,N_8818);
xor U9018 (N_9018,N_8958,N_8880);
nor U9019 (N_9019,N_8823,N_8851);
or U9020 (N_9020,N_8960,N_8885);
nand U9021 (N_9021,N_8990,N_8889);
nor U9022 (N_9022,N_8894,N_8812);
nand U9023 (N_9023,N_8984,N_8903);
nor U9024 (N_9024,N_8803,N_8899);
and U9025 (N_9025,N_8972,N_8806);
nand U9026 (N_9026,N_8986,N_8992);
and U9027 (N_9027,N_8952,N_8813);
nor U9028 (N_9028,N_8913,N_8814);
or U9029 (N_9029,N_8817,N_8846);
or U9030 (N_9030,N_8882,N_8834);
xnor U9031 (N_9031,N_8877,N_8975);
xor U9032 (N_9032,N_8989,N_8860);
xnor U9033 (N_9033,N_8977,N_8978);
or U9034 (N_9034,N_8983,N_8996);
or U9035 (N_9035,N_8921,N_8839);
and U9036 (N_9036,N_8808,N_8871);
xor U9037 (N_9037,N_8861,N_8849);
nor U9038 (N_9038,N_8888,N_8931);
or U9039 (N_9039,N_8837,N_8829);
or U9040 (N_9040,N_8912,N_8890);
nand U9041 (N_9041,N_8841,N_8920);
nand U9042 (N_9042,N_8825,N_8924);
xor U9043 (N_9043,N_8820,N_8917);
nand U9044 (N_9044,N_8895,N_8897);
and U9045 (N_9045,N_8980,N_8843);
or U9046 (N_9046,N_8988,N_8922);
xnor U9047 (N_9047,N_8852,N_8985);
or U9048 (N_9048,N_8831,N_8893);
xor U9049 (N_9049,N_8954,N_8807);
or U9050 (N_9050,N_8802,N_8953);
nand U9051 (N_9051,N_8937,N_8821);
or U9052 (N_9052,N_8859,N_8881);
or U9053 (N_9053,N_8867,N_8800);
nand U9054 (N_9054,N_8963,N_8930);
or U9055 (N_9055,N_8883,N_8929);
or U9056 (N_9056,N_8876,N_8965);
nand U9057 (N_9057,N_8943,N_8999);
nor U9058 (N_9058,N_8944,N_8911);
nor U9059 (N_9059,N_8875,N_8835);
xor U9060 (N_9060,N_8950,N_8886);
or U9061 (N_9061,N_8819,N_8936);
nand U9062 (N_9062,N_8909,N_8961);
nor U9063 (N_9063,N_8906,N_8884);
xnor U9064 (N_9064,N_8970,N_8853);
nand U9065 (N_9065,N_8946,N_8901);
nor U9066 (N_9066,N_8870,N_8918);
nand U9067 (N_9067,N_8940,N_8832);
xnor U9068 (N_9068,N_8855,N_8948);
nand U9069 (N_9069,N_8971,N_8902);
and U9070 (N_9070,N_8848,N_8945);
and U9071 (N_9071,N_8951,N_8927);
nand U9072 (N_9072,N_8962,N_8907);
or U9073 (N_9073,N_8865,N_8830);
and U9074 (N_9074,N_8810,N_8838);
xnor U9075 (N_9075,N_8981,N_8905);
nor U9076 (N_9076,N_8857,N_8811);
or U9077 (N_9077,N_8987,N_8879);
xor U9078 (N_9078,N_8916,N_8844);
nor U9079 (N_9079,N_8938,N_8997);
and U9080 (N_9080,N_8919,N_8863);
xnor U9081 (N_9081,N_8967,N_8969);
nand U9082 (N_9082,N_8824,N_8923);
and U9083 (N_9083,N_8816,N_8959);
nor U9084 (N_9084,N_8850,N_8827);
and U9085 (N_9085,N_8932,N_8873);
xnor U9086 (N_9086,N_8847,N_8822);
and U9087 (N_9087,N_8991,N_8828);
or U9088 (N_9088,N_8925,N_8979);
or U9089 (N_9089,N_8928,N_8869);
xor U9090 (N_9090,N_8833,N_8964);
and U9091 (N_9091,N_8845,N_8926);
or U9092 (N_9092,N_8934,N_8864);
and U9093 (N_9093,N_8956,N_8935);
and U9094 (N_9094,N_8973,N_8891);
and U9095 (N_9095,N_8805,N_8939);
or U9096 (N_9096,N_8957,N_8858);
xnor U9097 (N_9097,N_8801,N_8998);
and U9098 (N_9098,N_8949,N_8904);
xnor U9099 (N_9099,N_8974,N_8854);
nor U9100 (N_9100,N_8925,N_8851);
and U9101 (N_9101,N_8803,N_8887);
or U9102 (N_9102,N_8979,N_8882);
nor U9103 (N_9103,N_8921,N_8945);
and U9104 (N_9104,N_8813,N_8897);
or U9105 (N_9105,N_8869,N_8845);
xor U9106 (N_9106,N_8875,N_8970);
or U9107 (N_9107,N_8996,N_8898);
or U9108 (N_9108,N_8805,N_8937);
and U9109 (N_9109,N_8846,N_8819);
and U9110 (N_9110,N_8902,N_8889);
xor U9111 (N_9111,N_8921,N_8803);
and U9112 (N_9112,N_8829,N_8926);
or U9113 (N_9113,N_8981,N_8921);
and U9114 (N_9114,N_8880,N_8911);
nand U9115 (N_9115,N_8827,N_8915);
xnor U9116 (N_9116,N_8810,N_8941);
and U9117 (N_9117,N_8879,N_8800);
nor U9118 (N_9118,N_8883,N_8912);
xor U9119 (N_9119,N_8948,N_8876);
or U9120 (N_9120,N_8968,N_8873);
and U9121 (N_9121,N_8997,N_8854);
xnor U9122 (N_9122,N_8889,N_8912);
nand U9123 (N_9123,N_8834,N_8850);
or U9124 (N_9124,N_8824,N_8805);
nand U9125 (N_9125,N_8954,N_8950);
and U9126 (N_9126,N_8968,N_8801);
xor U9127 (N_9127,N_8942,N_8822);
xnor U9128 (N_9128,N_8996,N_8864);
nand U9129 (N_9129,N_8800,N_8888);
nand U9130 (N_9130,N_8932,N_8941);
xnor U9131 (N_9131,N_8815,N_8825);
or U9132 (N_9132,N_8848,N_8973);
and U9133 (N_9133,N_8911,N_8920);
xor U9134 (N_9134,N_8902,N_8861);
or U9135 (N_9135,N_8869,N_8922);
nand U9136 (N_9136,N_8841,N_8918);
xnor U9137 (N_9137,N_8980,N_8904);
xnor U9138 (N_9138,N_8819,N_8948);
nor U9139 (N_9139,N_8953,N_8851);
nand U9140 (N_9140,N_8861,N_8890);
nand U9141 (N_9141,N_8919,N_8875);
or U9142 (N_9142,N_8954,N_8842);
or U9143 (N_9143,N_8825,N_8921);
nor U9144 (N_9144,N_8878,N_8972);
or U9145 (N_9145,N_8826,N_8925);
nor U9146 (N_9146,N_8986,N_8909);
xor U9147 (N_9147,N_8868,N_8933);
nor U9148 (N_9148,N_8940,N_8981);
nor U9149 (N_9149,N_8953,N_8985);
or U9150 (N_9150,N_8935,N_8922);
and U9151 (N_9151,N_8941,N_8937);
nand U9152 (N_9152,N_8822,N_8998);
nand U9153 (N_9153,N_8995,N_8882);
nor U9154 (N_9154,N_8966,N_8962);
or U9155 (N_9155,N_8865,N_8975);
nor U9156 (N_9156,N_8831,N_8807);
xnor U9157 (N_9157,N_8837,N_8848);
xnor U9158 (N_9158,N_8908,N_8855);
nand U9159 (N_9159,N_8812,N_8934);
nand U9160 (N_9160,N_8962,N_8976);
nor U9161 (N_9161,N_8905,N_8980);
or U9162 (N_9162,N_8916,N_8826);
nor U9163 (N_9163,N_8806,N_8931);
nand U9164 (N_9164,N_8904,N_8969);
nand U9165 (N_9165,N_8973,N_8969);
or U9166 (N_9166,N_8882,N_8878);
xor U9167 (N_9167,N_8867,N_8812);
and U9168 (N_9168,N_8894,N_8868);
nand U9169 (N_9169,N_8984,N_8850);
nand U9170 (N_9170,N_8893,N_8952);
xor U9171 (N_9171,N_8813,N_8851);
xor U9172 (N_9172,N_8969,N_8820);
xnor U9173 (N_9173,N_8909,N_8837);
or U9174 (N_9174,N_8885,N_8970);
xor U9175 (N_9175,N_8838,N_8832);
nor U9176 (N_9176,N_8851,N_8969);
and U9177 (N_9177,N_8916,N_8964);
nand U9178 (N_9178,N_8960,N_8959);
nor U9179 (N_9179,N_8904,N_8857);
nor U9180 (N_9180,N_8818,N_8876);
and U9181 (N_9181,N_8801,N_8868);
and U9182 (N_9182,N_8998,N_8970);
xor U9183 (N_9183,N_8920,N_8832);
xnor U9184 (N_9184,N_8969,N_8872);
xnor U9185 (N_9185,N_8900,N_8903);
xor U9186 (N_9186,N_8990,N_8968);
xor U9187 (N_9187,N_8834,N_8845);
nor U9188 (N_9188,N_8805,N_8823);
and U9189 (N_9189,N_8822,N_8855);
and U9190 (N_9190,N_8944,N_8991);
or U9191 (N_9191,N_8902,N_8838);
xor U9192 (N_9192,N_8982,N_8960);
and U9193 (N_9193,N_8997,N_8815);
and U9194 (N_9194,N_8934,N_8929);
and U9195 (N_9195,N_8895,N_8870);
or U9196 (N_9196,N_8935,N_8923);
or U9197 (N_9197,N_8905,N_8827);
nand U9198 (N_9198,N_8927,N_8813);
xnor U9199 (N_9199,N_8883,N_8904);
and U9200 (N_9200,N_9053,N_9015);
or U9201 (N_9201,N_9139,N_9011);
and U9202 (N_9202,N_9173,N_9178);
nand U9203 (N_9203,N_9128,N_9054);
xor U9204 (N_9204,N_9070,N_9004);
nor U9205 (N_9205,N_9078,N_9061);
nor U9206 (N_9206,N_9144,N_9026);
and U9207 (N_9207,N_9059,N_9046);
nand U9208 (N_9208,N_9083,N_9087);
or U9209 (N_9209,N_9131,N_9189);
xor U9210 (N_9210,N_9159,N_9077);
and U9211 (N_9211,N_9039,N_9142);
nor U9212 (N_9212,N_9064,N_9071);
xnor U9213 (N_9213,N_9063,N_9109);
xnor U9214 (N_9214,N_9097,N_9001);
nor U9215 (N_9215,N_9007,N_9075);
and U9216 (N_9216,N_9067,N_9110);
or U9217 (N_9217,N_9082,N_9132);
xnor U9218 (N_9218,N_9029,N_9050);
nor U9219 (N_9219,N_9151,N_9192);
nor U9220 (N_9220,N_9025,N_9080);
nand U9221 (N_9221,N_9008,N_9085);
and U9222 (N_9222,N_9197,N_9081);
or U9223 (N_9223,N_9092,N_9091);
or U9224 (N_9224,N_9003,N_9058);
nor U9225 (N_9225,N_9019,N_9006);
and U9226 (N_9226,N_9055,N_9045);
nand U9227 (N_9227,N_9073,N_9016);
nor U9228 (N_9228,N_9154,N_9105);
xnor U9229 (N_9229,N_9176,N_9130);
xnor U9230 (N_9230,N_9000,N_9168);
and U9231 (N_9231,N_9199,N_9122);
or U9232 (N_9232,N_9032,N_9021);
nor U9233 (N_9233,N_9191,N_9020);
and U9234 (N_9234,N_9079,N_9009);
xnor U9235 (N_9235,N_9171,N_9174);
nor U9236 (N_9236,N_9121,N_9177);
nor U9237 (N_9237,N_9194,N_9014);
xnor U9238 (N_9238,N_9187,N_9115);
nor U9239 (N_9239,N_9164,N_9153);
nand U9240 (N_9240,N_9072,N_9106);
nand U9241 (N_9241,N_9140,N_9036);
nor U9242 (N_9242,N_9038,N_9195);
and U9243 (N_9243,N_9134,N_9024);
or U9244 (N_9244,N_9012,N_9179);
xnor U9245 (N_9245,N_9137,N_9065);
nand U9246 (N_9246,N_9031,N_9028);
nor U9247 (N_9247,N_9126,N_9141);
or U9248 (N_9248,N_9102,N_9183);
and U9249 (N_9249,N_9107,N_9033);
nand U9250 (N_9250,N_9157,N_9166);
or U9251 (N_9251,N_9198,N_9129);
nor U9252 (N_9252,N_9049,N_9022);
nor U9253 (N_9253,N_9099,N_9018);
nand U9254 (N_9254,N_9051,N_9124);
nand U9255 (N_9255,N_9162,N_9196);
and U9256 (N_9256,N_9108,N_9098);
and U9257 (N_9257,N_9114,N_9069);
xnor U9258 (N_9258,N_9112,N_9090);
xnor U9259 (N_9259,N_9143,N_9182);
xnor U9260 (N_9260,N_9158,N_9044);
or U9261 (N_9261,N_9035,N_9120);
and U9262 (N_9262,N_9165,N_9042);
nor U9263 (N_9263,N_9167,N_9169);
xor U9264 (N_9264,N_9104,N_9181);
and U9265 (N_9265,N_9146,N_9040);
or U9266 (N_9266,N_9010,N_9180);
nand U9267 (N_9267,N_9093,N_9062);
nor U9268 (N_9268,N_9136,N_9086);
or U9269 (N_9269,N_9125,N_9094);
or U9270 (N_9270,N_9117,N_9103);
and U9271 (N_9271,N_9160,N_9100);
and U9272 (N_9272,N_9096,N_9152);
xnor U9273 (N_9273,N_9138,N_9052);
and U9274 (N_9274,N_9190,N_9041);
and U9275 (N_9275,N_9147,N_9101);
or U9276 (N_9276,N_9066,N_9060);
and U9277 (N_9277,N_9149,N_9023);
nand U9278 (N_9278,N_9047,N_9127);
nand U9279 (N_9279,N_9172,N_9186);
xor U9280 (N_9280,N_9005,N_9161);
nand U9281 (N_9281,N_9017,N_9056);
xor U9282 (N_9282,N_9193,N_9068);
nor U9283 (N_9283,N_9175,N_9111);
nor U9284 (N_9284,N_9116,N_9057);
xor U9285 (N_9285,N_9030,N_9145);
xor U9286 (N_9286,N_9156,N_9002);
xnor U9287 (N_9287,N_9170,N_9148);
nand U9288 (N_9288,N_9113,N_9188);
and U9289 (N_9289,N_9163,N_9037);
and U9290 (N_9290,N_9074,N_9013);
nor U9291 (N_9291,N_9118,N_9150);
nand U9292 (N_9292,N_9043,N_9185);
nand U9293 (N_9293,N_9119,N_9034);
nand U9294 (N_9294,N_9095,N_9135);
and U9295 (N_9295,N_9076,N_9027);
nand U9296 (N_9296,N_9133,N_9088);
nand U9297 (N_9297,N_9184,N_9084);
nor U9298 (N_9298,N_9048,N_9155);
nor U9299 (N_9299,N_9123,N_9089);
xnor U9300 (N_9300,N_9074,N_9075);
xnor U9301 (N_9301,N_9192,N_9168);
or U9302 (N_9302,N_9100,N_9011);
nand U9303 (N_9303,N_9024,N_9174);
and U9304 (N_9304,N_9073,N_9075);
or U9305 (N_9305,N_9041,N_9002);
or U9306 (N_9306,N_9059,N_9050);
and U9307 (N_9307,N_9073,N_9063);
nor U9308 (N_9308,N_9048,N_9049);
nand U9309 (N_9309,N_9181,N_9014);
or U9310 (N_9310,N_9137,N_9108);
and U9311 (N_9311,N_9134,N_9070);
nand U9312 (N_9312,N_9181,N_9199);
nand U9313 (N_9313,N_9062,N_9187);
xnor U9314 (N_9314,N_9177,N_9089);
and U9315 (N_9315,N_9196,N_9178);
nor U9316 (N_9316,N_9130,N_9140);
nand U9317 (N_9317,N_9063,N_9108);
nor U9318 (N_9318,N_9062,N_9009);
nand U9319 (N_9319,N_9190,N_9113);
nor U9320 (N_9320,N_9023,N_9055);
and U9321 (N_9321,N_9083,N_9044);
nor U9322 (N_9322,N_9090,N_9067);
and U9323 (N_9323,N_9097,N_9058);
nand U9324 (N_9324,N_9176,N_9061);
xnor U9325 (N_9325,N_9058,N_9139);
xnor U9326 (N_9326,N_9116,N_9140);
nand U9327 (N_9327,N_9025,N_9152);
nand U9328 (N_9328,N_9033,N_9069);
and U9329 (N_9329,N_9001,N_9170);
xor U9330 (N_9330,N_9195,N_9015);
and U9331 (N_9331,N_9051,N_9149);
and U9332 (N_9332,N_9161,N_9199);
xnor U9333 (N_9333,N_9007,N_9194);
nand U9334 (N_9334,N_9004,N_9198);
or U9335 (N_9335,N_9151,N_9129);
and U9336 (N_9336,N_9145,N_9130);
or U9337 (N_9337,N_9196,N_9161);
and U9338 (N_9338,N_9013,N_9088);
xor U9339 (N_9339,N_9052,N_9165);
xnor U9340 (N_9340,N_9105,N_9153);
and U9341 (N_9341,N_9137,N_9122);
xnor U9342 (N_9342,N_9037,N_9076);
nor U9343 (N_9343,N_9033,N_9131);
nand U9344 (N_9344,N_9094,N_9020);
or U9345 (N_9345,N_9102,N_9046);
and U9346 (N_9346,N_9081,N_9155);
nor U9347 (N_9347,N_9048,N_9043);
nand U9348 (N_9348,N_9008,N_9146);
xnor U9349 (N_9349,N_9013,N_9138);
xor U9350 (N_9350,N_9080,N_9152);
xnor U9351 (N_9351,N_9093,N_9157);
nand U9352 (N_9352,N_9148,N_9147);
nand U9353 (N_9353,N_9173,N_9086);
or U9354 (N_9354,N_9037,N_9166);
nand U9355 (N_9355,N_9130,N_9150);
and U9356 (N_9356,N_9176,N_9063);
and U9357 (N_9357,N_9180,N_9175);
nand U9358 (N_9358,N_9024,N_9199);
xor U9359 (N_9359,N_9181,N_9155);
nor U9360 (N_9360,N_9065,N_9028);
or U9361 (N_9361,N_9142,N_9125);
or U9362 (N_9362,N_9006,N_9111);
nand U9363 (N_9363,N_9087,N_9171);
xor U9364 (N_9364,N_9099,N_9078);
or U9365 (N_9365,N_9068,N_9037);
and U9366 (N_9366,N_9180,N_9055);
xnor U9367 (N_9367,N_9186,N_9080);
or U9368 (N_9368,N_9083,N_9110);
xnor U9369 (N_9369,N_9010,N_9183);
and U9370 (N_9370,N_9092,N_9140);
or U9371 (N_9371,N_9150,N_9068);
and U9372 (N_9372,N_9009,N_9073);
and U9373 (N_9373,N_9066,N_9052);
xor U9374 (N_9374,N_9109,N_9050);
nor U9375 (N_9375,N_9021,N_9148);
nand U9376 (N_9376,N_9166,N_9129);
nand U9377 (N_9377,N_9089,N_9108);
xnor U9378 (N_9378,N_9194,N_9076);
or U9379 (N_9379,N_9087,N_9125);
xor U9380 (N_9380,N_9072,N_9059);
and U9381 (N_9381,N_9107,N_9096);
nand U9382 (N_9382,N_9173,N_9194);
and U9383 (N_9383,N_9014,N_9129);
nor U9384 (N_9384,N_9195,N_9190);
or U9385 (N_9385,N_9012,N_9116);
xor U9386 (N_9386,N_9077,N_9093);
or U9387 (N_9387,N_9060,N_9033);
xor U9388 (N_9388,N_9164,N_9036);
nor U9389 (N_9389,N_9053,N_9108);
nand U9390 (N_9390,N_9140,N_9083);
or U9391 (N_9391,N_9161,N_9061);
nor U9392 (N_9392,N_9147,N_9189);
nand U9393 (N_9393,N_9030,N_9185);
nor U9394 (N_9394,N_9021,N_9049);
nor U9395 (N_9395,N_9050,N_9023);
xnor U9396 (N_9396,N_9190,N_9164);
or U9397 (N_9397,N_9011,N_9098);
xor U9398 (N_9398,N_9081,N_9175);
xor U9399 (N_9399,N_9000,N_9090);
or U9400 (N_9400,N_9225,N_9263);
and U9401 (N_9401,N_9237,N_9389);
nor U9402 (N_9402,N_9306,N_9255);
nor U9403 (N_9403,N_9229,N_9242);
nor U9404 (N_9404,N_9217,N_9369);
or U9405 (N_9405,N_9256,N_9208);
nor U9406 (N_9406,N_9399,N_9294);
nand U9407 (N_9407,N_9329,N_9298);
nand U9408 (N_9408,N_9388,N_9379);
or U9409 (N_9409,N_9380,N_9324);
and U9410 (N_9410,N_9233,N_9333);
and U9411 (N_9411,N_9232,N_9371);
nor U9412 (N_9412,N_9206,N_9349);
and U9413 (N_9413,N_9384,N_9363);
nand U9414 (N_9414,N_9243,N_9377);
nor U9415 (N_9415,N_9202,N_9330);
nand U9416 (N_9416,N_9374,N_9254);
and U9417 (N_9417,N_9266,N_9316);
and U9418 (N_9418,N_9343,N_9364);
xor U9419 (N_9419,N_9271,N_9297);
and U9420 (N_9420,N_9395,N_9270);
nand U9421 (N_9421,N_9317,N_9354);
or U9422 (N_9422,N_9279,N_9230);
or U9423 (N_9423,N_9296,N_9328);
or U9424 (N_9424,N_9258,N_9355);
and U9425 (N_9425,N_9285,N_9336);
or U9426 (N_9426,N_9340,N_9239);
nand U9427 (N_9427,N_9338,N_9325);
or U9428 (N_9428,N_9353,N_9261);
xor U9429 (N_9429,N_9334,N_9362);
or U9430 (N_9430,N_9396,N_9247);
and U9431 (N_9431,N_9284,N_9302);
and U9432 (N_9432,N_9245,N_9265);
or U9433 (N_9433,N_9273,N_9210);
xor U9434 (N_9434,N_9268,N_9342);
xor U9435 (N_9435,N_9360,N_9301);
xor U9436 (N_9436,N_9385,N_9226);
or U9437 (N_9437,N_9357,N_9201);
nor U9438 (N_9438,N_9394,N_9323);
nand U9439 (N_9439,N_9315,N_9378);
or U9440 (N_9440,N_9209,N_9308);
nand U9441 (N_9441,N_9344,N_9367);
xnor U9442 (N_9442,N_9234,N_9356);
and U9443 (N_9443,N_9332,N_9219);
nand U9444 (N_9444,N_9264,N_9224);
nand U9445 (N_9445,N_9321,N_9269);
and U9446 (N_9446,N_9267,N_9207);
nor U9447 (N_9447,N_9326,N_9337);
nor U9448 (N_9448,N_9276,N_9305);
and U9449 (N_9449,N_9278,N_9288);
nor U9450 (N_9450,N_9293,N_9299);
xor U9451 (N_9451,N_9303,N_9238);
nor U9452 (N_9452,N_9300,N_9223);
and U9453 (N_9453,N_9319,N_9291);
nor U9454 (N_9454,N_9331,N_9204);
or U9455 (N_9455,N_9352,N_9365);
xor U9456 (N_9456,N_9272,N_9236);
nand U9457 (N_9457,N_9398,N_9382);
nor U9458 (N_9458,N_9283,N_9213);
xnor U9459 (N_9459,N_9361,N_9281);
xnor U9460 (N_9460,N_9235,N_9347);
and U9461 (N_9461,N_9251,N_9220);
nor U9462 (N_9462,N_9366,N_9253);
or U9463 (N_9463,N_9375,N_9228);
and U9464 (N_9464,N_9327,N_9383);
and U9465 (N_9465,N_9368,N_9313);
and U9466 (N_9466,N_9386,N_9322);
and U9467 (N_9467,N_9295,N_9227);
xor U9468 (N_9468,N_9311,N_9318);
xor U9469 (N_9469,N_9200,N_9348);
nor U9470 (N_9470,N_9370,N_9359);
and U9471 (N_9471,N_9214,N_9351);
xor U9472 (N_9472,N_9393,N_9286);
and U9473 (N_9473,N_9335,N_9287);
or U9474 (N_9474,N_9222,N_9277);
or U9475 (N_9475,N_9376,N_9290);
nand U9476 (N_9476,N_9312,N_9275);
or U9477 (N_9477,N_9260,N_9387);
nand U9478 (N_9478,N_9346,N_9274);
or U9479 (N_9479,N_9216,N_9381);
nand U9480 (N_9480,N_9203,N_9309);
nor U9481 (N_9481,N_9205,N_9250);
nor U9482 (N_9482,N_9246,N_9231);
or U9483 (N_9483,N_9390,N_9341);
and U9484 (N_9484,N_9307,N_9304);
and U9485 (N_9485,N_9314,N_9211);
and U9486 (N_9486,N_9244,N_9259);
nand U9487 (N_9487,N_9350,N_9310);
or U9488 (N_9488,N_9373,N_9248);
nand U9489 (N_9489,N_9257,N_9221);
nand U9490 (N_9490,N_9320,N_9241);
nand U9491 (N_9491,N_9240,N_9339);
or U9492 (N_9492,N_9252,N_9372);
and U9493 (N_9493,N_9358,N_9212);
or U9494 (N_9494,N_9282,N_9391);
and U9495 (N_9495,N_9249,N_9289);
nand U9496 (N_9496,N_9218,N_9345);
nand U9497 (N_9497,N_9292,N_9397);
nor U9498 (N_9498,N_9392,N_9215);
and U9499 (N_9499,N_9280,N_9262);
or U9500 (N_9500,N_9213,N_9393);
xor U9501 (N_9501,N_9307,N_9231);
and U9502 (N_9502,N_9212,N_9352);
and U9503 (N_9503,N_9209,N_9342);
and U9504 (N_9504,N_9281,N_9327);
xor U9505 (N_9505,N_9273,N_9337);
or U9506 (N_9506,N_9287,N_9390);
nor U9507 (N_9507,N_9289,N_9371);
xnor U9508 (N_9508,N_9358,N_9315);
and U9509 (N_9509,N_9381,N_9203);
nor U9510 (N_9510,N_9333,N_9264);
xor U9511 (N_9511,N_9315,N_9329);
nor U9512 (N_9512,N_9385,N_9223);
nor U9513 (N_9513,N_9243,N_9266);
nand U9514 (N_9514,N_9376,N_9242);
and U9515 (N_9515,N_9226,N_9258);
or U9516 (N_9516,N_9229,N_9274);
xor U9517 (N_9517,N_9293,N_9280);
xor U9518 (N_9518,N_9256,N_9229);
and U9519 (N_9519,N_9364,N_9385);
nor U9520 (N_9520,N_9281,N_9362);
or U9521 (N_9521,N_9375,N_9212);
and U9522 (N_9522,N_9359,N_9278);
nand U9523 (N_9523,N_9211,N_9322);
or U9524 (N_9524,N_9292,N_9285);
and U9525 (N_9525,N_9334,N_9381);
or U9526 (N_9526,N_9375,N_9373);
nor U9527 (N_9527,N_9357,N_9295);
xor U9528 (N_9528,N_9382,N_9335);
or U9529 (N_9529,N_9302,N_9270);
nand U9530 (N_9530,N_9325,N_9260);
nand U9531 (N_9531,N_9373,N_9345);
or U9532 (N_9532,N_9274,N_9288);
and U9533 (N_9533,N_9374,N_9223);
nor U9534 (N_9534,N_9244,N_9345);
and U9535 (N_9535,N_9305,N_9257);
nand U9536 (N_9536,N_9317,N_9381);
nor U9537 (N_9537,N_9219,N_9323);
xor U9538 (N_9538,N_9353,N_9268);
and U9539 (N_9539,N_9270,N_9306);
xor U9540 (N_9540,N_9204,N_9371);
nor U9541 (N_9541,N_9319,N_9343);
xor U9542 (N_9542,N_9387,N_9219);
xor U9543 (N_9543,N_9312,N_9322);
xnor U9544 (N_9544,N_9210,N_9358);
or U9545 (N_9545,N_9273,N_9315);
nand U9546 (N_9546,N_9343,N_9384);
and U9547 (N_9547,N_9376,N_9227);
nand U9548 (N_9548,N_9304,N_9368);
and U9549 (N_9549,N_9368,N_9243);
or U9550 (N_9550,N_9276,N_9399);
or U9551 (N_9551,N_9213,N_9241);
nand U9552 (N_9552,N_9362,N_9346);
nor U9553 (N_9553,N_9369,N_9341);
and U9554 (N_9554,N_9320,N_9343);
nand U9555 (N_9555,N_9355,N_9254);
nor U9556 (N_9556,N_9322,N_9240);
and U9557 (N_9557,N_9239,N_9361);
and U9558 (N_9558,N_9315,N_9263);
nand U9559 (N_9559,N_9308,N_9280);
and U9560 (N_9560,N_9284,N_9242);
nor U9561 (N_9561,N_9335,N_9323);
nand U9562 (N_9562,N_9345,N_9391);
nor U9563 (N_9563,N_9322,N_9244);
xor U9564 (N_9564,N_9228,N_9220);
xnor U9565 (N_9565,N_9292,N_9239);
xnor U9566 (N_9566,N_9334,N_9231);
xnor U9567 (N_9567,N_9237,N_9354);
nand U9568 (N_9568,N_9338,N_9329);
nand U9569 (N_9569,N_9264,N_9330);
nor U9570 (N_9570,N_9318,N_9215);
or U9571 (N_9571,N_9201,N_9340);
nor U9572 (N_9572,N_9247,N_9375);
and U9573 (N_9573,N_9224,N_9222);
or U9574 (N_9574,N_9209,N_9253);
and U9575 (N_9575,N_9374,N_9306);
or U9576 (N_9576,N_9357,N_9315);
and U9577 (N_9577,N_9231,N_9284);
nand U9578 (N_9578,N_9345,N_9323);
xnor U9579 (N_9579,N_9307,N_9363);
xnor U9580 (N_9580,N_9235,N_9308);
nand U9581 (N_9581,N_9283,N_9309);
xor U9582 (N_9582,N_9238,N_9254);
and U9583 (N_9583,N_9266,N_9395);
nand U9584 (N_9584,N_9227,N_9344);
xnor U9585 (N_9585,N_9391,N_9250);
xnor U9586 (N_9586,N_9200,N_9393);
or U9587 (N_9587,N_9305,N_9230);
or U9588 (N_9588,N_9397,N_9275);
nand U9589 (N_9589,N_9291,N_9387);
or U9590 (N_9590,N_9399,N_9348);
nor U9591 (N_9591,N_9363,N_9232);
nor U9592 (N_9592,N_9206,N_9340);
xnor U9593 (N_9593,N_9216,N_9240);
xnor U9594 (N_9594,N_9340,N_9395);
or U9595 (N_9595,N_9230,N_9398);
nand U9596 (N_9596,N_9380,N_9372);
nand U9597 (N_9597,N_9377,N_9379);
and U9598 (N_9598,N_9398,N_9361);
and U9599 (N_9599,N_9363,N_9234);
nor U9600 (N_9600,N_9480,N_9565);
nand U9601 (N_9601,N_9502,N_9587);
xnor U9602 (N_9602,N_9520,N_9523);
or U9603 (N_9603,N_9521,N_9552);
nand U9604 (N_9604,N_9596,N_9514);
xor U9605 (N_9605,N_9487,N_9469);
xnor U9606 (N_9606,N_9586,N_9403);
nor U9607 (N_9607,N_9465,N_9434);
or U9608 (N_9608,N_9474,N_9462);
nor U9609 (N_9609,N_9575,N_9513);
or U9610 (N_9610,N_9582,N_9430);
nand U9611 (N_9611,N_9554,N_9570);
nand U9612 (N_9612,N_9432,N_9450);
xor U9613 (N_9613,N_9420,N_9553);
or U9614 (N_9614,N_9467,N_9549);
and U9615 (N_9615,N_9478,N_9519);
or U9616 (N_9616,N_9571,N_9441);
and U9617 (N_9617,N_9454,N_9561);
nand U9618 (N_9618,N_9557,N_9400);
or U9619 (N_9619,N_9529,N_9449);
nor U9620 (N_9620,N_9444,N_9483);
nand U9621 (N_9621,N_9528,N_9416);
and U9622 (N_9622,N_9488,N_9532);
or U9623 (N_9623,N_9564,N_9537);
or U9624 (N_9624,N_9579,N_9422);
nand U9625 (N_9625,N_9536,N_9563);
nor U9626 (N_9626,N_9473,N_9511);
xnor U9627 (N_9627,N_9481,N_9506);
and U9628 (N_9628,N_9461,N_9540);
nand U9629 (N_9629,N_9578,N_9541);
or U9630 (N_9630,N_9583,N_9494);
nand U9631 (N_9631,N_9415,N_9512);
or U9632 (N_9632,N_9452,N_9566);
nand U9633 (N_9633,N_9427,N_9475);
xnor U9634 (N_9634,N_9476,N_9484);
nand U9635 (N_9635,N_9580,N_9562);
xor U9636 (N_9636,N_9412,N_9567);
xor U9637 (N_9637,N_9477,N_9492);
nor U9638 (N_9638,N_9468,N_9401);
nor U9639 (N_9639,N_9515,N_9550);
nand U9640 (N_9640,N_9504,N_9471);
or U9641 (N_9641,N_9499,N_9414);
and U9642 (N_9642,N_9509,N_9581);
and U9643 (N_9643,N_9457,N_9518);
and U9644 (N_9644,N_9531,N_9428);
nand U9645 (N_9645,N_9507,N_9530);
nor U9646 (N_9646,N_9495,N_9417);
xnor U9647 (N_9647,N_9472,N_9439);
and U9648 (N_9648,N_9446,N_9524);
nand U9649 (N_9649,N_9542,N_9577);
xnor U9650 (N_9650,N_9595,N_9404);
nand U9651 (N_9651,N_9408,N_9493);
or U9652 (N_9652,N_9576,N_9589);
nor U9653 (N_9653,N_9546,N_9435);
xor U9654 (N_9654,N_9436,N_9497);
nand U9655 (N_9655,N_9501,N_9431);
xnor U9656 (N_9656,N_9433,N_9442);
or U9657 (N_9657,N_9545,N_9437);
nor U9658 (N_9658,N_9423,N_9426);
and U9659 (N_9659,N_9505,N_9558);
and U9660 (N_9660,N_9489,N_9503);
nor U9661 (N_9661,N_9419,N_9538);
nand U9662 (N_9662,N_9459,N_9555);
and U9663 (N_9663,N_9411,N_9539);
or U9664 (N_9664,N_9421,N_9598);
nand U9665 (N_9665,N_9445,N_9522);
or U9666 (N_9666,N_9405,N_9590);
and U9667 (N_9667,N_9424,N_9543);
or U9668 (N_9668,N_9479,N_9410);
or U9669 (N_9669,N_9486,N_9560);
or U9670 (N_9670,N_9517,N_9496);
nor U9671 (N_9671,N_9548,N_9406);
xor U9672 (N_9672,N_9547,N_9413);
nor U9673 (N_9673,N_9407,N_9568);
nand U9674 (N_9674,N_9510,N_9599);
nand U9675 (N_9675,N_9451,N_9429);
nor U9676 (N_9676,N_9491,N_9593);
and U9677 (N_9677,N_9490,N_9573);
or U9678 (N_9678,N_9470,N_9526);
nand U9679 (N_9679,N_9485,N_9588);
xor U9680 (N_9680,N_9500,N_9425);
nand U9681 (N_9681,N_9525,N_9440);
xor U9682 (N_9682,N_9533,N_9443);
and U9683 (N_9683,N_9458,N_9551);
and U9684 (N_9684,N_9402,N_9556);
or U9685 (N_9685,N_9527,N_9482);
nor U9686 (N_9686,N_9585,N_9455);
nor U9687 (N_9687,N_9409,N_9535);
nand U9688 (N_9688,N_9463,N_9447);
xor U9689 (N_9689,N_9448,N_9594);
and U9690 (N_9690,N_9534,N_9574);
and U9691 (N_9691,N_9453,N_9466);
and U9692 (N_9692,N_9572,N_9597);
or U9693 (N_9693,N_9498,N_9591);
nand U9694 (N_9694,N_9460,N_9508);
and U9695 (N_9695,N_9544,N_9584);
xor U9696 (N_9696,N_9464,N_9559);
and U9697 (N_9697,N_9418,N_9516);
or U9698 (N_9698,N_9456,N_9438);
xnor U9699 (N_9699,N_9569,N_9592);
nor U9700 (N_9700,N_9554,N_9451);
and U9701 (N_9701,N_9527,N_9469);
and U9702 (N_9702,N_9459,N_9449);
nor U9703 (N_9703,N_9583,N_9539);
nor U9704 (N_9704,N_9507,N_9469);
xor U9705 (N_9705,N_9535,N_9498);
nor U9706 (N_9706,N_9442,N_9587);
and U9707 (N_9707,N_9407,N_9553);
nand U9708 (N_9708,N_9407,N_9439);
xnor U9709 (N_9709,N_9429,N_9516);
nand U9710 (N_9710,N_9475,N_9486);
nor U9711 (N_9711,N_9533,N_9410);
nand U9712 (N_9712,N_9430,N_9459);
xor U9713 (N_9713,N_9562,N_9443);
nand U9714 (N_9714,N_9515,N_9540);
and U9715 (N_9715,N_9583,N_9438);
xor U9716 (N_9716,N_9409,N_9487);
xor U9717 (N_9717,N_9503,N_9586);
xor U9718 (N_9718,N_9526,N_9418);
and U9719 (N_9719,N_9419,N_9487);
or U9720 (N_9720,N_9505,N_9540);
xnor U9721 (N_9721,N_9432,N_9442);
and U9722 (N_9722,N_9423,N_9526);
nor U9723 (N_9723,N_9447,N_9477);
nor U9724 (N_9724,N_9449,N_9403);
nand U9725 (N_9725,N_9573,N_9463);
nor U9726 (N_9726,N_9475,N_9559);
or U9727 (N_9727,N_9508,N_9523);
and U9728 (N_9728,N_9505,N_9526);
xor U9729 (N_9729,N_9532,N_9452);
xor U9730 (N_9730,N_9501,N_9558);
xor U9731 (N_9731,N_9487,N_9544);
or U9732 (N_9732,N_9508,N_9527);
or U9733 (N_9733,N_9499,N_9430);
xor U9734 (N_9734,N_9534,N_9456);
or U9735 (N_9735,N_9567,N_9515);
nor U9736 (N_9736,N_9430,N_9502);
nand U9737 (N_9737,N_9560,N_9591);
nor U9738 (N_9738,N_9540,N_9431);
xnor U9739 (N_9739,N_9462,N_9504);
nor U9740 (N_9740,N_9518,N_9528);
xnor U9741 (N_9741,N_9427,N_9419);
xnor U9742 (N_9742,N_9503,N_9453);
nor U9743 (N_9743,N_9484,N_9448);
nand U9744 (N_9744,N_9513,N_9506);
or U9745 (N_9745,N_9599,N_9418);
or U9746 (N_9746,N_9418,N_9428);
nand U9747 (N_9747,N_9534,N_9419);
or U9748 (N_9748,N_9520,N_9419);
or U9749 (N_9749,N_9413,N_9485);
and U9750 (N_9750,N_9473,N_9449);
nor U9751 (N_9751,N_9597,N_9545);
and U9752 (N_9752,N_9492,N_9595);
nor U9753 (N_9753,N_9411,N_9502);
or U9754 (N_9754,N_9444,N_9419);
nand U9755 (N_9755,N_9558,N_9537);
nor U9756 (N_9756,N_9448,N_9568);
nand U9757 (N_9757,N_9523,N_9554);
xnor U9758 (N_9758,N_9498,N_9537);
nor U9759 (N_9759,N_9463,N_9589);
or U9760 (N_9760,N_9484,N_9478);
nor U9761 (N_9761,N_9543,N_9403);
xnor U9762 (N_9762,N_9579,N_9567);
or U9763 (N_9763,N_9469,N_9461);
or U9764 (N_9764,N_9516,N_9409);
nand U9765 (N_9765,N_9589,N_9598);
xnor U9766 (N_9766,N_9568,N_9518);
nor U9767 (N_9767,N_9413,N_9400);
or U9768 (N_9768,N_9405,N_9410);
xnor U9769 (N_9769,N_9499,N_9558);
nor U9770 (N_9770,N_9505,N_9545);
nor U9771 (N_9771,N_9505,N_9517);
or U9772 (N_9772,N_9580,N_9476);
nor U9773 (N_9773,N_9420,N_9552);
and U9774 (N_9774,N_9475,N_9431);
nand U9775 (N_9775,N_9409,N_9539);
xor U9776 (N_9776,N_9576,N_9499);
nand U9777 (N_9777,N_9477,N_9425);
nand U9778 (N_9778,N_9578,N_9428);
or U9779 (N_9779,N_9463,N_9472);
and U9780 (N_9780,N_9536,N_9498);
nor U9781 (N_9781,N_9405,N_9461);
xor U9782 (N_9782,N_9486,N_9439);
xnor U9783 (N_9783,N_9520,N_9492);
or U9784 (N_9784,N_9503,N_9418);
and U9785 (N_9785,N_9574,N_9531);
and U9786 (N_9786,N_9548,N_9451);
xor U9787 (N_9787,N_9503,N_9533);
nand U9788 (N_9788,N_9442,N_9514);
nor U9789 (N_9789,N_9553,N_9506);
or U9790 (N_9790,N_9575,N_9594);
nand U9791 (N_9791,N_9504,N_9570);
and U9792 (N_9792,N_9512,N_9448);
xnor U9793 (N_9793,N_9421,N_9565);
nand U9794 (N_9794,N_9423,N_9566);
xor U9795 (N_9795,N_9581,N_9579);
nor U9796 (N_9796,N_9495,N_9482);
and U9797 (N_9797,N_9563,N_9524);
nand U9798 (N_9798,N_9531,N_9421);
nor U9799 (N_9799,N_9510,N_9463);
nor U9800 (N_9800,N_9759,N_9707);
xor U9801 (N_9801,N_9696,N_9635);
nand U9802 (N_9802,N_9626,N_9723);
xnor U9803 (N_9803,N_9665,N_9602);
xnor U9804 (N_9804,N_9666,N_9603);
and U9805 (N_9805,N_9680,N_9640);
and U9806 (N_9806,N_9737,N_9623);
xnor U9807 (N_9807,N_9670,N_9650);
or U9808 (N_9808,N_9729,N_9649);
nor U9809 (N_9809,N_9761,N_9777);
nand U9810 (N_9810,N_9620,N_9714);
xor U9811 (N_9811,N_9719,N_9728);
xor U9812 (N_9812,N_9684,N_9645);
or U9813 (N_9813,N_9653,N_9746);
nor U9814 (N_9814,N_9648,N_9745);
nand U9815 (N_9815,N_9773,N_9789);
and U9816 (N_9816,N_9618,N_9630);
or U9817 (N_9817,N_9611,N_9652);
nor U9818 (N_9818,N_9796,N_9776);
xor U9819 (N_9819,N_9772,N_9739);
and U9820 (N_9820,N_9610,N_9664);
nand U9821 (N_9821,N_9685,N_9713);
nor U9822 (N_9822,N_9758,N_9643);
nor U9823 (N_9823,N_9724,N_9753);
or U9824 (N_9824,N_9614,N_9633);
xor U9825 (N_9825,N_9698,N_9711);
and U9826 (N_9826,N_9612,N_9693);
nor U9827 (N_9827,N_9625,N_9683);
and U9828 (N_9828,N_9712,N_9795);
or U9829 (N_9829,N_9629,N_9659);
xnor U9830 (N_9830,N_9688,N_9690);
nor U9831 (N_9831,N_9725,N_9654);
xnor U9832 (N_9832,N_9733,N_9646);
nand U9833 (N_9833,N_9669,N_9634);
and U9834 (N_9834,N_9744,N_9686);
and U9835 (N_9835,N_9655,N_9661);
xnor U9836 (N_9836,N_9624,N_9770);
xor U9837 (N_9837,N_9769,N_9700);
and U9838 (N_9838,N_9681,N_9720);
nor U9839 (N_9839,N_9619,N_9705);
nand U9840 (N_9840,N_9768,N_9793);
and U9841 (N_9841,N_9657,N_9798);
or U9842 (N_9842,N_9694,N_9775);
or U9843 (N_9843,N_9736,N_9703);
nor U9844 (N_9844,N_9609,N_9701);
nor U9845 (N_9845,N_9656,N_9721);
nand U9846 (N_9846,N_9794,N_9644);
or U9847 (N_9847,N_9667,N_9692);
nor U9848 (N_9848,N_9608,N_9740);
nand U9849 (N_9849,N_9735,N_9742);
and U9850 (N_9850,N_9651,N_9722);
nand U9851 (N_9851,N_9780,N_9781);
xor U9852 (N_9852,N_9731,N_9764);
xnor U9853 (N_9853,N_9615,N_9697);
xnor U9854 (N_9854,N_9734,N_9660);
nand U9855 (N_9855,N_9674,N_9787);
xnor U9856 (N_9856,N_9606,N_9658);
nand U9857 (N_9857,N_9704,N_9699);
nand U9858 (N_9858,N_9749,N_9671);
xnor U9859 (N_9859,N_9783,N_9799);
xnor U9860 (N_9860,N_9621,N_9617);
xnor U9861 (N_9861,N_9672,N_9767);
nand U9862 (N_9862,N_9689,N_9727);
or U9863 (N_9863,N_9771,N_9679);
xor U9864 (N_9864,N_9600,N_9791);
and U9865 (N_9865,N_9784,N_9642);
nand U9866 (N_9866,N_9718,N_9668);
and U9867 (N_9867,N_9748,N_9709);
and U9868 (N_9868,N_9639,N_9647);
or U9869 (N_9869,N_9779,N_9763);
or U9870 (N_9870,N_9687,N_9716);
nand U9871 (N_9871,N_9628,N_9604);
nand U9872 (N_9872,N_9663,N_9786);
nand U9873 (N_9873,N_9751,N_9662);
and U9874 (N_9874,N_9788,N_9706);
and U9875 (N_9875,N_9616,N_9778);
xor U9876 (N_9876,N_9797,N_9792);
nor U9877 (N_9877,N_9785,N_9677);
and U9878 (N_9878,N_9691,N_9607);
nor U9879 (N_9879,N_9782,N_9675);
xor U9880 (N_9880,N_9752,N_9710);
and U9881 (N_9881,N_9613,N_9765);
nand U9882 (N_9882,N_9638,N_9738);
xor U9883 (N_9883,N_9756,N_9743);
nand U9884 (N_9884,N_9766,N_9676);
and U9885 (N_9885,N_9702,N_9732);
xor U9886 (N_9886,N_9730,N_9622);
nand U9887 (N_9887,N_9673,N_9755);
nor U9888 (N_9888,N_9682,N_9695);
or U9889 (N_9889,N_9750,N_9741);
and U9890 (N_9890,N_9760,N_9637);
or U9891 (N_9891,N_9754,N_9726);
and U9892 (N_9892,N_9632,N_9708);
nor U9893 (N_9893,N_9678,N_9747);
nand U9894 (N_9894,N_9757,N_9762);
and U9895 (N_9895,N_9631,N_9790);
nor U9896 (N_9896,N_9605,N_9715);
nand U9897 (N_9897,N_9774,N_9641);
xnor U9898 (N_9898,N_9636,N_9627);
and U9899 (N_9899,N_9601,N_9717);
nor U9900 (N_9900,N_9799,N_9760);
and U9901 (N_9901,N_9699,N_9758);
and U9902 (N_9902,N_9735,N_9793);
nand U9903 (N_9903,N_9611,N_9793);
xnor U9904 (N_9904,N_9668,N_9776);
and U9905 (N_9905,N_9750,N_9742);
nor U9906 (N_9906,N_9700,N_9709);
nor U9907 (N_9907,N_9787,N_9688);
nor U9908 (N_9908,N_9706,N_9779);
xnor U9909 (N_9909,N_9704,N_9748);
nor U9910 (N_9910,N_9707,N_9679);
or U9911 (N_9911,N_9715,N_9791);
nor U9912 (N_9912,N_9748,N_9770);
and U9913 (N_9913,N_9760,N_9753);
or U9914 (N_9914,N_9622,N_9697);
nor U9915 (N_9915,N_9764,N_9758);
xor U9916 (N_9916,N_9603,N_9692);
nor U9917 (N_9917,N_9639,N_9697);
xor U9918 (N_9918,N_9672,N_9710);
or U9919 (N_9919,N_9689,N_9744);
xnor U9920 (N_9920,N_9717,N_9719);
nand U9921 (N_9921,N_9785,N_9601);
or U9922 (N_9922,N_9767,N_9648);
and U9923 (N_9923,N_9606,N_9733);
nor U9924 (N_9924,N_9794,N_9738);
and U9925 (N_9925,N_9747,N_9787);
or U9926 (N_9926,N_9620,N_9764);
or U9927 (N_9927,N_9736,N_9722);
and U9928 (N_9928,N_9646,N_9788);
or U9929 (N_9929,N_9718,N_9728);
and U9930 (N_9930,N_9703,N_9735);
nand U9931 (N_9931,N_9743,N_9689);
and U9932 (N_9932,N_9628,N_9676);
xor U9933 (N_9933,N_9695,N_9748);
nand U9934 (N_9934,N_9678,N_9688);
and U9935 (N_9935,N_9771,N_9614);
nor U9936 (N_9936,N_9674,N_9732);
or U9937 (N_9937,N_9649,N_9622);
nor U9938 (N_9938,N_9620,N_9706);
nor U9939 (N_9939,N_9734,N_9699);
or U9940 (N_9940,N_9785,N_9774);
nand U9941 (N_9941,N_9659,N_9670);
or U9942 (N_9942,N_9683,N_9719);
nand U9943 (N_9943,N_9789,N_9733);
or U9944 (N_9944,N_9734,N_9673);
or U9945 (N_9945,N_9628,N_9687);
nor U9946 (N_9946,N_9708,N_9747);
nor U9947 (N_9947,N_9675,N_9766);
xor U9948 (N_9948,N_9769,N_9656);
and U9949 (N_9949,N_9787,N_9720);
and U9950 (N_9950,N_9790,N_9614);
nand U9951 (N_9951,N_9758,N_9680);
nand U9952 (N_9952,N_9761,N_9633);
nor U9953 (N_9953,N_9703,N_9789);
nand U9954 (N_9954,N_9735,N_9731);
nor U9955 (N_9955,N_9776,N_9768);
xnor U9956 (N_9956,N_9630,N_9629);
xor U9957 (N_9957,N_9708,N_9720);
or U9958 (N_9958,N_9782,N_9705);
xnor U9959 (N_9959,N_9644,N_9770);
or U9960 (N_9960,N_9668,N_9664);
or U9961 (N_9961,N_9741,N_9677);
nand U9962 (N_9962,N_9603,N_9791);
xnor U9963 (N_9963,N_9774,N_9766);
or U9964 (N_9964,N_9600,N_9628);
nor U9965 (N_9965,N_9794,N_9746);
xnor U9966 (N_9966,N_9719,N_9729);
nor U9967 (N_9967,N_9634,N_9680);
xor U9968 (N_9968,N_9682,N_9606);
nand U9969 (N_9969,N_9656,N_9738);
nor U9970 (N_9970,N_9726,N_9713);
nand U9971 (N_9971,N_9783,N_9720);
xnor U9972 (N_9972,N_9699,N_9659);
nor U9973 (N_9973,N_9774,N_9602);
and U9974 (N_9974,N_9691,N_9780);
nand U9975 (N_9975,N_9608,N_9754);
xnor U9976 (N_9976,N_9735,N_9734);
nand U9977 (N_9977,N_9785,N_9783);
xnor U9978 (N_9978,N_9731,N_9639);
nand U9979 (N_9979,N_9783,N_9754);
nor U9980 (N_9980,N_9720,N_9731);
or U9981 (N_9981,N_9630,N_9678);
xor U9982 (N_9982,N_9763,N_9780);
and U9983 (N_9983,N_9712,N_9626);
or U9984 (N_9984,N_9656,N_9622);
or U9985 (N_9985,N_9765,N_9633);
nand U9986 (N_9986,N_9701,N_9759);
nand U9987 (N_9987,N_9628,N_9677);
and U9988 (N_9988,N_9635,N_9742);
and U9989 (N_9989,N_9740,N_9605);
or U9990 (N_9990,N_9708,N_9770);
xor U9991 (N_9991,N_9789,N_9661);
or U9992 (N_9992,N_9747,N_9609);
nand U9993 (N_9993,N_9710,N_9669);
or U9994 (N_9994,N_9777,N_9746);
or U9995 (N_9995,N_9738,N_9748);
and U9996 (N_9996,N_9703,N_9751);
nand U9997 (N_9997,N_9710,N_9742);
xnor U9998 (N_9998,N_9710,N_9620);
nor U9999 (N_9999,N_9722,N_9617);
and UO_0 (O_0,N_9847,N_9815);
xor UO_1 (O_1,N_9875,N_9800);
nand UO_2 (O_2,N_9839,N_9950);
xor UO_3 (O_3,N_9897,N_9860);
nor UO_4 (O_4,N_9862,N_9904);
xor UO_5 (O_5,N_9840,N_9980);
and UO_6 (O_6,N_9976,N_9983);
nand UO_7 (O_7,N_9825,N_9816);
or UO_8 (O_8,N_9932,N_9958);
and UO_9 (O_9,N_9898,N_9929);
and UO_10 (O_10,N_9977,N_9968);
xnor UO_11 (O_11,N_9824,N_9808);
and UO_12 (O_12,N_9827,N_9984);
and UO_13 (O_13,N_9996,N_9817);
nor UO_14 (O_14,N_9919,N_9835);
xor UO_15 (O_15,N_9990,N_9812);
xnor UO_16 (O_16,N_9991,N_9908);
nand UO_17 (O_17,N_9803,N_9972);
and UO_18 (O_18,N_9936,N_9969);
or UO_19 (O_19,N_9838,N_9842);
nor UO_20 (O_20,N_9918,N_9841);
nor UO_21 (O_21,N_9981,N_9818);
or UO_22 (O_22,N_9834,N_9831);
nand UO_23 (O_23,N_9924,N_9809);
nand UO_24 (O_24,N_9903,N_9952);
nor UO_25 (O_25,N_9870,N_9964);
nor UO_26 (O_26,N_9961,N_9883);
and UO_27 (O_27,N_9855,N_9999);
and UO_28 (O_28,N_9820,N_9994);
xnor UO_29 (O_29,N_9806,N_9829);
or UO_30 (O_30,N_9873,N_9985);
nand UO_31 (O_31,N_9998,N_9905);
nand UO_32 (O_32,N_9896,N_9988);
xnor UO_33 (O_33,N_9966,N_9975);
and UO_34 (O_34,N_9986,N_9931);
or UO_35 (O_35,N_9890,N_9844);
nand UO_36 (O_36,N_9913,N_9830);
nor UO_37 (O_37,N_9956,N_9833);
and UO_38 (O_38,N_9869,N_9902);
xnor UO_39 (O_39,N_9974,N_9849);
and UO_40 (O_40,N_9881,N_9948);
nand UO_41 (O_41,N_9911,N_9920);
and UO_42 (O_42,N_9843,N_9814);
or UO_43 (O_43,N_9861,N_9802);
or UO_44 (O_44,N_9947,N_9995);
and UO_45 (O_45,N_9971,N_9893);
nor UO_46 (O_46,N_9959,N_9876);
nor UO_47 (O_47,N_9993,N_9942);
nor UO_48 (O_48,N_9954,N_9805);
nor UO_49 (O_49,N_9845,N_9891);
and UO_50 (O_50,N_9933,N_9863);
and UO_51 (O_51,N_9851,N_9850);
xor UO_52 (O_52,N_9953,N_9865);
nor UO_53 (O_53,N_9997,N_9877);
nand UO_54 (O_54,N_9946,N_9941);
or UO_55 (O_55,N_9857,N_9982);
or UO_56 (O_56,N_9963,N_9852);
and UO_57 (O_57,N_9819,N_9837);
and UO_58 (O_58,N_9955,N_9979);
nor UO_59 (O_59,N_9895,N_9886);
nand UO_60 (O_60,N_9922,N_9872);
nand UO_61 (O_61,N_9810,N_9868);
nand UO_62 (O_62,N_9992,N_9879);
or UO_63 (O_63,N_9866,N_9889);
nand UO_64 (O_64,N_9871,N_9989);
and UO_65 (O_65,N_9951,N_9935);
nand UO_66 (O_66,N_9926,N_9848);
xor UO_67 (O_67,N_9928,N_9813);
nor UO_68 (O_68,N_9943,N_9965);
xnor UO_69 (O_69,N_9909,N_9960);
xor UO_70 (O_70,N_9970,N_9858);
and UO_71 (O_71,N_9957,N_9937);
nor UO_72 (O_72,N_9973,N_9804);
nor UO_73 (O_73,N_9912,N_9826);
xor UO_74 (O_74,N_9821,N_9828);
nand UO_75 (O_75,N_9940,N_9892);
and UO_76 (O_76,N_9944,N_9923);
or UO_77 (O_77,N_9894,N_9962);
and UO_78 (O_78,N_9885,N_9856);
or UO_79 (O_79,N_9811,N_9874);
nand UO_80 (O_80,N_9949,N_9906);
or UO_81 (O_81,N_9938,N_9859);
nor UO_82 (O_82,N_9880,N_9927);
or UO_83 (O_83,N_9884,N_9978);
nand UO_84 (O_84,N_9916,N_9939);
and UO_85 (O_85,N_9900,N_9930);
nor UO_86 (O_86,N_9823,N_9846);
and UO_87 (O_87,N_9832,N_9822);
nor UO_88 (O_88,N_9934,N_9914);
xnor UO_89 (O_89,N_9917,N_9864);
nand UO_90 (O_90,N_9899,N_9925);
and UO_91 (O_91,N_9807,N_9921);
or UO_92 (O_92,N_9867,N_9836);
nand UO_93 (O_93,N_9853,N_9854);
nand UO_94 (O_94,N_9901,N_9945);
or UO_95 (O_95,N_9801,N_9878);
xnor UO_96 (O_96,N_9907,N_9910);
nor UO_97 (O_97,N_9888,N_9887);
and UO_98 (O_98,N_9915,N_9987);
or UO_99 (O_99,N_9882,N_9967);
or UO_100 (O_100,N_9950,N_9964);
and UO_101 (O_101,N_9993,N_9826);
or UO_102 (O_102,N_9850,N_9820);
nor UO_103 (O_103,N_9977,N_9957);
and UO_104 (O_104,N_9819,N_9874);
and UO_105 (O_105,N_9827,N_9888);
nor UO_106 (O_106,N_9862,N_9832);
nand UO_107 (O_107,N_9978,N_9806);
and UO_108 (O_108,N_9876,N_9917);
xor UO_109 (O_109,N_9872,N_9998);
or UO_110 (O_110,N_9891,N_9951);
and UO_111 (O_111,N_9905,N_9825);
xor UO_112 (O_112,N_9996,N_9824);
nand UO_113 (O_113,N_9866,N_9884);
nor UO_114 (O_114,N_9921,N_9847);
and UO_115 (O_115,N_9884,N_9986);
xor UO_116 (O_116,N_9948,N_9897);
nand UO_117 (O_117,N_9990,N_9927);
and UO_118 (O_118,N_9930,N_9941);
and UO_119 (O_119,N_9804,N_9937);
nor UO_120 (O_120,N_9858,N_9954);
and UO_121 (O_121,N_9893,N_9881);
or UO_122 (O_122,N_9848,N_9822);
nor UO_123 (O_123,N_9972,N_9917);
nor UO_124 (O_124,N_9959,N_9840);
xnor UO_125 (O_125,N_9908,N_9912);
and UO_126 (O_126,N_9872,N_9833);
xnor UO_127 (O_127,N_9943,N_9870);
xor UO_128 (O_128,N_9850,N_9983);
and UO_129 (O_129,N_9881,N_9873);
xor UO_130 (O_130,N_9827,N_9900);
xnor UO_131 (O_131,N_9819,N_9906);
or UO_132 (O_132,N_9811,N_9897);
nor UO_133 (O_133,N_9984,N_9803);
xor UO_134 (O_134,N_9903,N_9858);
xor UO_135 (O_135,N_9898,N_9955);
nand UO_136 (O_136,N_9894,N_9807);
or UO_137 (O_137,N_9873,N_9854);
nor UO_138 (O_138,N_9986,N_9863);
nand UO_139 (O_139,N_9838,N_9986);
xor UO_140 (O_140,N_9829,N_9988);
xor UO_141 (O_141,N_9905,N_9832);
and UO_142 (O_142,N_9838,N_9905);
nor UO_143 (O_143,N_9814,N_9807);
and UO_144 (O_144,N_9904,N_9976);
nand UO_145 (O_145,N_9856,N_9888);
and UO_146 (O_146,N_9988,N_9905);
or UO_147 (O_147,N_9869,N_9930);
nand UO_148 (O_148,N_9925,N_9879);
and UO_149 (O_149,N_9975,N_9809);
and UO_150 (O_150,N_9802,N_9890);
or UO_151 (O_151,N_9843,N_9887);
nand UO_152 (O_152,N_9963,N_9930);
xor UO_153 (O_153,N_9825,N_9851);
or UO_154 (O_154,N_9873,N_9822);
nor UO_155 (O_155,N_9829,N_9945);
nand UO_156 (O_156,N_9832,N_9873);
and UO_157 (O_157,N_9953,N_9932);
nor UO_158 (O_158,N_9913,N_9927);
or UO_159 (O_159,N_9859,N_9906);
nor UO_160 (O_160,N_9807,N_9906);
xor UO_161 (O_161,N_9948,N_9858);
or UO_162 (O_162,N_9888,N_9897);
or UO_163 (O_163,N_9914,N_9926);
nand UO_164 (O_164,N_9895,N_9960);
nor UO_165 (O_165,N_9988,N_9820);
xor UO_166 (O_166,N_9815,N_9892);
or UO_167 (O_167,N_9815,N_9988);
xnor UO_168 (O_168,N_9879,N_9829);
nor UO_169 (O_169,N_9898,N_9932);
xor UO_170 (O_170,N_9986,N_9902);
xor UO_171 (O_171,N_9809,N_9972);
or UO_172 (O_172,N_9925,N_9910);
nand UO_173 (O_173,N_9934,N_9818);
nor UO_174 (O_174,N_9968,N_9829);
and UO_175 (O_175,N_9894,N_9869);
or UO_176 (O_176,N_9998,N_9915);
nor UO_177 (O_177,N_9907,N_9979);
or UO_178 (O_178,N_9941,N_9977);
nand UO_179 (O_179,N_9957,N_9834);
nand UO_180 (O_180,N_9833,N_9929);
nand UO_181 (O_181,N_9974,N_9883);
nor UO_182 (O_182,N_9987,N_9825);
or UO_183 (O_183,N_9886,N_9876);
or UO_184 (O_184,N_9872,N_9847);
nor UO_185 (O_185,N_9927,N_9960);
or UO_186 (O_186,N_9846,N_9943);
nor UO_187 (O_187,N_9843,N_9904);
and UO_188 (O_188,N_9811,N_9814);
nor UO_189 (O_189,N_9991,N_9804);
and UO_190 (O_190,N_9826,N_9960);
xor UO_191 (O_191,N_9906,N_9801);
nand UO_192 (O_192,N_9872,N_9897);
xnor UO_193 (O_193,N_9805,N_9808);
xor UO_194 (O_194,N_9974,N_9957);
nor UO_195 (O_195,N_9987,N_9974);
xor UO_196 (O_196,N_9882,N_9957);
or UO_197 (O_197,N_9857,N_9835);
and UO_198 (O_198,N_9853,N_9838);
nor UO_199 (O_199,N_9966,N_9912);
nand UO_200 (O_200,N_9951,N_9948);
and UO_201 (O_201,N_9937,N_9916);
xor UO_202 (O_202,N_9868,N_9825);
xnor UO_203 (O_203,N_9860,N_9821);
and UO_204 (O_204,N_9950,N_9937);
nor UO_205 (O_205,N_9821,N_9980);
and UO_206 (O_206,N_9813,N_9984);
xnor UO_207 (O_207,N_9963,N_9853);
or UO_208 (O_208,N_9823,N_9987);
and UO_209 (O_209,N_9860,N_9825);
xor UO_210 (O_210,N_9858,N_9975);
or UO_211 (O_211,N_9856,N_9971);
nand UO_212 (O_212,N_9915,N_9821);
xor UO_213 (O_213,N_9999,N_9857);
and UO_214 (O_214,N_9965,N_9927);
nor UO_215 (O_215,N_9932,N_9926);
nor UO_216 (O_216,N_9838,N_9911);
and UO_217 (O_217,N_9840,N_9961);
nand UO_218 (O_218,N_9912,N_9999);
nand UO_219 (O_219,N_9927,N_9872);
nor UO_220 (O_220,N_9944,N_9829);
nand UO_221 (O_221,N_9864,N_9955);
xnor UO_222 (O_222,N_9890,N_9948);
nor UO_223 (O_223,N_9961,N_9803);
xor UO_224 (O_224,N_9816,N_9916);
or UO_225 (O_225,N_9843,N_9833);
xor UO_226 (O_226,N_9952,N_9959);
nand UO_227 (O_227,N_9885,N_9973);
and UO_228 (O_228,N_9875,N_9948);
nor UO_229 (O_229,N_9881,N_9865);
or UO_230 (O_230,N_9837,N_9832);
and UO_231 (O_231,N_9858,N_9939);
and UO_232 (O_232,N_9855,N_9948);
xnor UO_233 (O_233,N_9871,N_9876);
or UO_234 (O_234,N_9815,N_9819);
and UO_235 (O_235,N_9932,N_9881);
xor UO_236 (O_236,N_9884,N_9993);
nand UO_237 (O_237,N_9837,N_9971);
or UO_238 (O_238,N_9939,N_9898);
and UO_239 (O_239,N_9978,N_9870);
and UO_240 (O_240,N_9873,N_9931);
nand UO_241 (O_241,N_9920,N_9936);
or UO_242 (O_242,N_9802,N_9838);
or UO_243 (O_243,N_9882,N_9917);
nand UO_244 (O_244,N_9888,N_9807);
xnor UO_245 (O_245,N_9827,N_9970);
xor UO_246 (O_246,N_9992,N_9875);
nor UO_247 (O_247,N_9801,N_9937);
nor UO_248 (O_248,N_9888,N_9857);
xor UO_249 (O_249,N_9944,N_9860);
nand UO_250 (O_250,N_9897,N_9884);
xnor UO_251 (O_251,N_9807,N_9915);
nor UO_252 (O_252,N_9935,N_9851);
or UO_253 (O_253,N_9979,N_9903);
xnor UO_254 (O_254,N_9878,N_9991);
and UO_255 (O_255,N_9987,N_9866);
nor UO_256 (O_256,N_9951,N_9949);
xnor UO_257 (O_257,N_9924,N_9810);
xnor UO_258 (O_258,N_9914,N_9941);
nor UO_259 (O_259,N_9931,N_9923);
nor UO_260 (O_260,N_9979,N_9895);
xnor UO_261 (O_261,N_9825,N_9889);
nand UO_262 (O_262,N_9980,N_9936);
and UO_263 (O_263,N_9934,N_9991);
nor UO_264 (O_264,N_9886,N_9951);
nor UO_265 (O_265,N_9905,N_9890);
nor UO_266 (O_266,N_9852,N_9905);
nor UO_267 (O_267,N_9872,N_9971);
or UO_268 (O_268,N_9962,N_9985);
nor UO_269 (O_269,N_9952,N_9823);
xnor UO_270 (O_270,N_9986,N_9889);
or UO_271 (O_271,N_9909,N_9927);
xnor UO_272 (O_272,N_9937,N_9889);
nand UO_273 (O_273,N_9866,N_9885);
nor UO_274 (O_274,N_9832,N_9860);
xor UO_275 (O_275,N_9894,N_9872);
or UO_276 (O_276,N_9832,N_9919);
and UO_277 (O_277,N_9878,N_9926);
xnor UO_278 (O_278,N_9893,N_9970);
xnor UO_279 (O_279,N_9950,N_9870);
and UO_280 (O_280,N_9965,N_9924);
nand UO_281 (O_281,N_9854,N_9817);
nor UO_282 (O_282,N_9858,N_9814);
or UO_283 (O_283,N_9969,N_9835);
and UO_284 (O_284,N_9940,N_9958);
nand UO_285 (O_285,N_9877,N_9805);
xnor UO_286 (O_286,N_9895,N_9835);
or UO_287 (O_287,N_9973,N_9955);
nor UO_288 (O_288,N_9924,N_9803);
nor UO_289 (O_289,N_9881,N_9943);
xor UO_290 (O_290,N_9820,N_9999);
nor UO_291 (O_291,N_9980,N_9876);
nor UO_292 (O_292,N_9956,N_9970);
nand UO_293 (O_293,N_9996,N_9881);
nor UO_294 (O_294,N_9916,N_9849);
and UO_295 (O_295,N_9887,N_9922);
and UO_296 (O_296,N_9995,N_9852);
and UO_297 (O_297,N_9884,N_9961);
nor UO_298 (O_298,N_9962,N_9858);
or UO_299 (O_299,N_9828,N_9918);
nand UO_300 (O_300,N_9909,N_9866);
xnor UO_301 (O_301,N_9987,N_9856);
xnor UO_302 (O_302,N_9958,N_9864);
or UO_303 (O_303,N_9929,N_9838);
nor UO_304 (O_304,N_9806,N_9944);
nor UO_305 (O_305,N_9862,N_9891);
nand UO_306 (O_306,N_9875,N_9820);
and UO_307 (O_307,N_9814,N_9864);
and UO_308 (O_308,N_9809,N_9917);
and UO_309 (O_309,N_9946,N_9966);
nand UO_310 (O_310,N_9910,N_9932);
or UO_311 (O_311,N_9800,N_9809);
and UO_312 (O_312,N_9810,N_9853);
and UO_313 (O_313,N_9842,N_9805);
nand UO_314 (O_314,N_9933,N_9867);
xnor UO_315 (O_315,N_9856,N_9994);
or UO_316 (O_316,N_9886,N_9919);
and UO_317 (O_317,N_9821,N_9853);
xor UO_318 (O_318,N_9922,N_9856);
nand UO_319 (O_319,N_9939,N_9848);
and UO_320 (O_320,N_9983,N_9880);
xor UO_321 (O_321,N_9907,N_9986);
nand UO_322 (O_322,N_9880,N_9862);
and UO_323 (O_323,N_9924,N_9954);
or UO_324 (O_324,N_9851,N_9905);
xnor UO_325 (O_325,N_9943,N_9810);
or UO_326 (O_326,N_9916,N_9981);
nand UO_327 (O_327,N_9867,N_9864);
and UO_328 (O_328,N_9967,N_9830);
or UO_329 (O_329,N_9974,N_9845);
and UO_330 (O_330,N_9858,N_9902);
nand UO_331 (O_331,N_9911,N_9852);
or UO_332 (O_332,N_9823,N_9985);
xnor UO_333 (O_333,N_9803,N_9926);
or UO_334 (O_334,N_9801,N_9871);
and UO_335 (O_335,N_9961,N_9951);
nand UO_336 (O_336,N_9950,N_9963);
and UO_337 (O_337,N_9818,N_9843);
nor UO_338 (O_338,N_9841,N_9998);
nor UO_339 (O_339,N_9927,N_9924);
nor UO_340 (O_340,N_9995,N_9980);
xnor UO_341 (O_341,N_9863,N_9885);
nand UO_342 (O_342,N_9909,N_9962);
xor UO_343 (O_343,N_9948,N_9893);
xor UO_344 (O_344,N_9871,N_9817);
xnor UO_345 (O_345,N_9883,N_9980);
and UO_346 (O_346,N_9829,N_9810);
nand UO_347 (O_347,N_9809,N_9885);
and UO_348 (O_348,N_9833,N_9909);
xor UO_349 (O_349,N_9884,N_9830);
and UO_350 (O_350,N_9809,N_9925);
xor UO_351 (O_351,N_9848,N_9973);
nand UO_352 (O_352,N_9976,N_9939);
or UO_353 (O_353,N_9904,N_9931);
nor UO_354 (O_354,N_9992,N_9801);
nor UO_355 (O_355,N_9859,N_9987);
or UO_356 (O_356,N_9947,N_9993);
or UO_357 (O_357,N_9980,N_9867);
nor UO_358 (O_358,N_9958,N_9946);
xnor UO_359 (O_359,N_9838,N_9854);
or UO_360 (O_360,N_9931,N_9897);
nand UO_361 (O_361,N_9812,N_9821);
nor UO_362 (O_362,N_9983,N_9815);
nand UO_363 (O_363,N_9856,N_9847);
nand UO_364 (O_364,N_9920,N_9800);
and UO_365 (O_365,N_9969,N_9820);
and UO_366 (O_366,N_9972,N_9993);
or UO_367 (O_367,N_9988,N_9985);
xor UO_368 (O_368,N_9957,N_9939);
nand UO_369 (O_369,N_9899,N_9836);
nor UO_370 (O_370,N_9817,N_9914);
xnor UO_371 (O_371,N_9935,N_9842);
or UO_372 (O_372,N_9991,N_9821);
nor UO_373 (O_373,N_9994,N_9878);
or UO_374 (O_374,N_9909,N_9817);
xor UO_375 (O_375,N_9982,N_9975);
and UO_376 (O_376,N_9901,N_9915);
nor UO_377 (O_377,N_9967,N_9954);
or UO_378 (O_378,N_9892,N_9919);
xnor UO_379 (O_379,N_9870,N_9961);
and UO_380 (O_380,N_9809,N_9968);
nand UO_381 (O_381,N_9841,N_9856);
xnor UO_382 (O_382,N_9913,N_9930);
nand UO_383 (O_383,N_9952,N_9907);
nand UO_384 (O_384,N_9895,N_9956);
nor UO_385 (O_385,N_9814,N_9817);
or UO_386 (O_386,N_9900,N_9810);
nor UO_387 (O_387,N_9964,N_9977);
xnor UO_388 (O_388,N_9894,N_9868);
nand UO_389 (O_389,N_9819,N_9839);
or UO_390 (O_390,N_9814,N_9865);
or UO_391 (O_391,N_9843,N_9926);
nor UO_392 (O_392,N_9811,N_9864);
nand UO_393 (O_393,N_9865,N_9993);
nor UO_394 (O_394,N_9892,N_9894);
xor UO_395 (O_395,N_9929,N_9985);
and UO_396 (O_396,N_9811,N_9932);
nor UO_397 (O_397,N_9912,N_9895);
or UO_398 (O_398,N_9893,N_9860);
xor UO_399 (O_399,N_9830,N_9821);
or UO_400 (O_400,N_9908,N_9938);
and UO_401 (O_401,N_9923,N_9909);
nor UO_402 (O_402,N_9831,N_9808);
xor UO_403 (O_403,N_9986,N_9873);
or UO_404 (O_404,N_9864,N_9919);
nor UO_405 (O_405,N_9998,N_9936);
and UO_406 (O_406,N_9937,N_9985);
and UO_407 (O_407,N_9942,N_9888);
or UO_408 (O_408,N_9899,N_9962);
or UO_409 (O_409,N_9900,N_9907);
and UO_410 (O_410,N_9938,N_9963);
nor UO_411 (O_411,N_9802,N_9811);
nand UO_412 (O_412,N_9901,N_9900);
or UO_413 (O_413,N_9862,N_9888);
nor UO_414 (O_414,N_9881,N_9998);
xor UO_415 (O_415,N_9875,N_9971);
nand UO_416 (O_416,N_9922,N_9803);
and UO_417 (O_417,N_9883,N_9928);
and UO_418 (O_418,N_9927,N_9925);
and UO_419 (O_419,N_9829,N_9820);
and UO_420 (O_420,N_9975,N_9996);
or UO_421 (O_421,N_9844,N_9860);
nor UO_422 (O_422,N_9970,N_9811);
nand UO_423 (O_423,N_9840,N_9800);
or UO_424 (O_424,N_9811,N_9919);
or UO_425 (O_425,N_9852,N_9808);
nand UO_426 (O_426,N_9943,N_9859);
xnor UO_427 (O_427,N_9897,N_9837);
xor UO_428 (O_428,N_9995,N_9816);
xor UO_429 (O_429,N_9910,N_9950);
nor UO_430 (O_430,N_9941,N_9806);
and UO_431 (O_431,N_9898,N_9961);
xnor UO_432 (O_432,N_9851,N_9896);
xor UO_433 (O_433,N_9862,N_9834);
and UO_434 (O_434,N_9863,N_9995);
nor UO_435 (O_435,N_9804,N_9965);
nor UO_436 (O_436,N_9802,N_9961);
xnor UO_437 (O_437,N_9916,N_9941);
or UO_438 (O_438,N_9874,N_9917);
nand UO_439 (O_439,N_9918,N_9824);
or UO_440 (O_440,N_9825,N_9940);
nand UO_441 (O_441,N_9849,N_9954);
nor UO_442 (O_442,N_9996,N_9916);
nand UO_443 (O_443,N_9869,N_9989);
nand UO_444 (O_444,N_9928,N_9926);
nor UO_445 (O_445,N_9861,N_9839);
nand UO_446 (O_446,N_9863,N_9922);
xor UO_447 (O_447,N_9863,N_9918);
nand UO_448 (O_448,N_9989,N_9802);
nand UO_449 (O_449,N_9872,N_9843);
nor UO_450 (O_450,N_9846,N_9898);
nor UO_451 (O_451,N_9974,N_9930);
and UO_452 (O_452,N_9805,N_9825);
and UO_453 (O_453,N_9873,N_9899);
nor UO_454 (O_454,N_9977,N_9980);
and UO_455 (O_455,N_9987,N_9890);
nand UO_456 (O_456,N_9992,N_9844);
nand UO_457 (O_457,N_9987,N_9800);
and UO_458 (O_458,N_9975,N_9886);
nor UO_459 (O_459,N_9809,N_9963);
xnor UO_460 (O_460,N_9957,N_9932);
nor UO_461 (O_461,N_9970,N_9873);
or UO_462 (O_462,N_9961,N_9916);
xnor UO_463 (O_463,N_9980,N_9967);
and UO_464 (O_464,N_9881,N_9899);
xnor UO_465 (O_465,N_9919,N_9839);
xor UO_466 (O_466,N_9833,N_9984);
or UO_467 (O_467,N_9890,N_9834);
xor UO_468 (O_468,N_9857,N_9885);
and UO_469 (O_469,N_9811,N_9940);
or UO_470 (O_470,N_9884,N_9816);
nor UO_471 (O_471,N_9852,N_9892);
nor UO_472 (O_472,N_9842,N_9911);
nor UO_473 (O_473,N_9988,N_9917);
nand UO_474 (O_474,N_9895,N_9899);
and UO_475 (O_475,N_9837,N_9933);
and UO_476 (O_476,N_9911,N_9882);
xnor UO_477 (O_477,N_9808,N_9943);
nor UO_478 (O_478,N_9832,N_9913);
nor UO_479 (O_479,N_9936,N_9959);
and UO_480 (O_480,N_9996,N_9844);
xor UO_481 (O_481,N_9991,N_9814);
xor UO_482 (O_482,N_9901,N_9808);
xor UO_483 (O_483,N_9926,N_9809);
nand UO_484 (O_484,N_9863,N_9818);
xnor UO_485 (O_485,N_9915,N_9814);
xor UO_486 (O_486,N_9837,N_9986);
nand UO_487 (O_487,N_9952,N_9902);
nand UO_488 (O_488,N_9807,N_9980);
nor UO_489 (O_489,N_9965,N_9964);
and UO_490 (O_490,N_9939,N_9983);
nor UO_491 (O_491,N_9974,N_9969);
nor UO_492 (O_492,N_9976,N_9910);
and UO_493 (O_493,N_9823,N_9821);
nand UO_494 (O_494,N_9917,N_9940);
and UO_495 (O_495,N_9902,N_9911);
or UO_496 (O_496,N_9814,N_9804);
xor UO_497 (O_497,N_9985,N_9871);
or UO_498 (O_498,N_9898,N_9819);
nor UO_499 (O_499,N_9887,N_9821);
nor UO_500 (O_500,N_9972,N_9923);
nor UO_501 (O_501,N_9924,N_9886);
or UO_502 (O_502,N_9975,N_9936);
and UO_503 (O_503,N_9862,N_9992);
and UO_504 (O_504,N_9916,N_9933);
nand UO_505 (O_505,N_9984,N_9960);
nor UO_506 (O_506,N_9888,N_9930);
nor UO_507 (O_507,N_9880,N_9849);
nand UO_508 (O_508,N_9984,N_9900);
xor UO_509 (O_509,N_9969,N_9883);
nor UO_510 (O_510,N_9852,N_9902);
nand UO_511 (O_511,N_9866,N_9916);
xor UO_512 (O_512,N_9928,N_9863);
or UO_513 (O_513,N_9880,N_9957);
xnor UO_514 (O_514,N_9824,N_9928);
xor UO_515 (O_515,N_9881,N_9977);
xnor UO_516 (O_516,N_9925,N_9922);
or UO_517 (O_517,N_9905,N_9950);
xnor UO_518 (O_518,N_9912,N_9935);
nor UO_519 (O_519,N_9860,N_9892);
nand UO_520 (O_520,N_9991,N_9807);
or UO_521 (O_521,N_9848,N_9827);
or UO_522 (O_522,N_9839,N_9969);
nand UO_523 (O_523,N_9929,N_9839);
nand UO_524 (O_524,N_9887,N_9952);
nand UO_525 (O_525,N_9877,N_9836);
nand UO_526 (O_526,N_9939,N_9844);
or UO_527 (O_527,N_9961,N_9881);
and UO_528 (O_528,N_9874,N_9993);
nor UO_529 (O_529,N_9991,N_9902);
or UO_530 (O_530,N_9968,N_9867);
and UO_531 (O_531,N_9929,N_9801);
xnor UO_532 (O_532,N_9801,N_9942);
nand UO_533 (O_533,N_9870,N_9939);
xor UO_534 (O_534,N_9954,N_9955);
or UO_535 (O_535,N_9984,N_9851);
or UO_536 (O_536,N_9989,N_9859);
nor UO_537 (O_537,N_9988,N_9929);
nand UO_538 (O_538,N_9833,N_9832);
nor UO_539 (O_539,N_9904,N_9927);
nor UO_540 (O_540,N_9830,N_9807);
nand UO_541 (O_541,N_9968,N_9882);
or UO_542 (O_542,N_9843,N_9804);
nor UO_543 (O_543,N_9937,N_9830);
nor UO_544 (O_544,N_9849,N_9995);
and UO_545 (O_545,N_9941,N_9928);
xor UO_546 (O_546,N_9927,N_9939);
nor UO_547 (O_547,N_9966,N_9863);
nand UO_548 (O_548,N_9826,N_9918);
or UO_549 (O_549,N_9979,N_9835);
and UO_550 (O_550,N_9876,N_9946);
or UO_551 (O_551,N_9928,N_9956);
xnor UO_552 (O_552,N_9934,N_9834);
and UO_553 (O_553,N_9919,N_9945);
or UO_554 (O_554,N_9990,N_9935);
nand UO_555 (O_555,N_9935,N_9861);
and UO_556 (O_556,N_9902,N_9849);
nor UO_557 (O_557,N_9868,N_9973);
and UO_558 (O_558,N_9986,N_9979);
nand UO_559 (O_559,N_9900,N_9886);
or UO_560 (O_560,N_9945,N_9878);
nand UO_561 (O_561,N_9870,N_9811);
xor UO_562 (O_562,N_9878,N_9853);
and UO_563 (O_563,N_9942,N_9827);
nand UO_564 (O_564,N_9879,N_9949);
nand UO_565 (O_565,N_9999,N_9961);
xor UO_566 (O_566,N_9992,N_9853);
or UO_567 (O_567,N_9901,N_9865);
and UO_568 (O_568,N_9851,N_9883);
nand UO_569 (O_569,N_9979,N_9959);
nor UO_570 (O_570,N_9892,N_9850);
nand UO_571 (O_571,N_9898,N_9908);
or UO_572 (O_572,N_9867,N_9993);
nand UO_573 (O_573,N_9857,N_9830);
and UO_574 (O_574,N_9804,N_9828);
nor UO_575 (O_575,N_9902,N_9838);
nor UO_576 (O_576,N_9985,N_9810);
or UO_577 (O_577,N_9972,N_9907);
xor UO_578 (O_578,N_9976,N_9875);
nand UO_579 (O_579,N_9955,N_9884);
xnor UO_580 (O_580,N_9911,N_9953);
xor UO_581 (O_581,N_9994,N_9912);
xor UO_582 (O_582,N_9868,N_9835);
and UO_583 (O_583,N_9854,N_9945);
xor UO_584 (O_584,N_9875,N_9956);
xnor UO_585 (O_585,N_9953,N_9809);
nand UO_586 (O_586,N_9829,N_9954);
xnor UO_587 (O_587,N_9843,N_9858);
and UO_588 (O_588,N_9845,N_9890);
nand UO_589 (O_589,N_9859,N_9804);
nand UO_590 (O_590,N_9859,N_9809);
xnor UO_591 (O_591,N_9832,N_9852);
and UO_592 (O_592,N_9816,N_9863);
nor UO_593 (O_593,N_9813,N_9920);
nand UO_594 (O_594,N_9979,N_9973);
and UO_595 (O_595,N_9923,N_9823);
nand UO_596 (O_596,N_9851,N_9992);
and UO_597 (O_597,N_9881,N_9854);
nand UO_598 (O_598,N_9948,N_9848);
or UO_599 (O_599,N_9807,N_9834);
and UO_600 (O_600,N_9961,N_9983);
or UO_601 (O_601,N_9870,N_9871);
xor UO_602 (O_602,N_9936,N_9955);
nor UO_603 (O_603,N_9816,N_9862);
and UO_604 (O_604,N_9980,N_9990);
nor UO_605 (O_605,N_9964,N_9929);
nor UO_606 (O_606,N_9947,N_9987);
nor UO_607 (O_607,N_9960,N_9989);
xnor UO_608 (O_608,N_9900,N_9970);
xnor UO_609 (O_609,N_9988,N_9951);
nand UO_610 (O_610,N_9884,N_9810);
and UO_611 (O_611,N_9897,N_9951);
nor UO_612 (O_612,N_9835,N_9841);
nor UO_613 (O_613,N_9928,N_9981);
and UO_614 (O_614,N_9828,N_9994);
xor UO_615 (O_615,N_9904,N_9903);
or UO_616 (O_616,N_9963,N_9811);
or UO_617 (O_617,N_9989,N_9986);
or UO_618 (O_618,N_9918,N_9995);
or UO_619 (O_619,N_9820,N_9839);
xnor UO_620 (O_620,N_9956,N_9941);
and UO_621 (O_621,N_9987,N_9850);
xnor UO_622 (O_622,N_9876,N_9867);
xor UO_623 (O_623,N_9957,N_9868);
nor UO_624 (O_624,N_9962,N_9848);
or UO_625 (O_625,N_9937,N_9932);
or UO_626 (O_626,N_9896,N_9897);
and UO_627 (O_627,N_9834,N_9938);
or UO_628 (O_628,N_9838,N_9801);
and UO_629 (O_629,N_9823,N_9835);
nand UO_630 (O_630,N_9963,N_9882);
and UO_631 (O_631,N_9891,N_9972);
nand UO_632 (O_632,N_9954,N_9898);
nand UO_633 (O_633,N_9994,N_9891);
xor UO_634 (O_634,N_9967,N_9970);
nor UO_635 (O_635,N_9842,N_9852);
xnor UO_636 (O_636,N_9885,N_9932);
and UO_637 (O_637,N_9940,N_9820);
xor UO_638 (O_638,N_9811,N_9885);
nand UO_639 (O_639,N_9812,N_9899);
and UO_640 (O_640,N_9832,N_9869);
nand UO_641 (O_641,N_9835,N_9972);
nor UO_642 (O_642,N_9842,N_9867);
and UO_643 (O_643,N_9932,N_9833);
and UO_644 (O_644,N_9906,N_9831);
nor UO_645 (O_645,N_9892,N_9842);
and UO_646 (O_646,N_9910,N_9862);
or UO_647 (O_647,N_9944,N_9823);
and UO_648 (O_648,N_9906,N_9886);
nand UO_649 (O_649,N_9955,N_9989);
nand UO_650 (O_650,N_9993,N_9971);
and UO_651 (O_651,N_9992,N_9961);
or UO_652 (O_652,N_9875,N_9964);
nand UO_653 (O_653,N_9837,N_9943);
or UO_654 (O_654,N_9992,N_9954);
nand UO_655 (O_655,N_9959,N_9802);
nor UO_656 (O_656,N_9926,N_9950);
nand UO_657 (O_657,N_9918,N_9885);
nor UO_658 (O_658,N_9875,N_9868);
nand UO_659 (O_659,N_9811,N_9848);
or UO_660 (O_660,N_9873,N_9908);
xor UO_661 (O_661,N_9907,N_9938);
and UO_662 (O_662,N_9840,N_9933);
nor UO_663 (O_663,N_9928,N_9915);
nor UO_664 (O_664,N_9829,N_9870);
or UO_665 (O_665,N_9821,N_9914);
xnor UO_666 (O_666,N_9924,N_9864);
nand UO_667 (O_667,N_9807,N_9987);
or UO_668 (O_668,N_9990,N_9842);
nor UO_669 (O_669,N_9979,N_9872);
and UO_670 (O_670,N_9958,N_9894);
nand UO_671 (O_671,N_9976,N_9818);
xnor UO_672 (O_672,N_9854,N_9919);
and UO_673 (O_673,N_9859,N_9909);
nor UO_674 (O_674,N_9821,N_9926);
xnor UO_675 (O_675,N_9886,N_9998);
or UO_676 (O_676,N_9886,N_9973);
or UO_677 (O_677,N_9995,N_9862);
and UO_678 (O_678,N_9970,N_9854);
xor UO_679 (O_679,N_9932,N_9938);
and UO_680 (O_680,N_9972,N_9834);
xor UO_681 (O_681,N_9836,N_9809);
xor UO_682 (O_682,N_9849,N_9858);
or UO_683 (O_683,N_9858,N_9862);
and UO_684 (O_684,N_9852,N_9868);
or UO_685 (O_685,N_9932,N_9802);
xor UO_686 (O_686,N_9910,N_9917);
nor UO_687 (O_687,N_9884,N_9856);
nand UO_688 (O_688,N_9920,N_9805);
nor UO_689 (O_689,N_9850,N_9837);
nand UO_690 (O_690,N_9887,N_9925);
and UO_691 (O_691,N_9887,N_9802);
xnor UO_692 (O_692,N_9964,N_9913);
nor UO_693 (O_693,N_9817,N_9828);
nor UO_694 (O_694,N_9947,N_9833);
and UO_695 (O_695,N_9877,N_9898);
or UO_696 (O_696,N_9972,N_9893);
nand UO_697 (O_697,N_9940,N_9823);
nand UO_698 (O_698,N_9975,N_9947);
xor UO_699 (O_699,N_9837,N_9921);
xnor UO_700 (O_700,N_9897,N_9827);
nor UO_701 (O_701,N_9860,N_9906);
xor UO_702 (O_702,N_9808,N_9926);
xnor UO_703 (O_703,N_9856,N_9946);
nor UO_704 (O_704,N_9950,N_9897);
xnor UO_705 (O_705,N_9820,N_9836);
nor UO_706 (O_706,N_9883,N_9881);
xnor UO_707 (O_707,N_9935,N_9980);
nor UO_708 (O_708,N_9966,N_9802);
nor UO_709 (O_709,N_9987,N_9877);
xnor UO_710 (O_710,N_9932,N_9879);
nand UO_711 (O_711,N_9860,N_9880);
nor UO_712 (O_712,N_9852,N_9858);
and UO_713 (O_713,N_9838,N_9873);
and UO_714 (O_714,N_9875,N_9951);
and UO_715 (O_715,N_9937,N_9908);
nor UO_716 (O_716,N_9910,N_9872);
nand UO_717 (O_717,N_9954,N_9897);
nand UO_718 (O_718,N_9981,N_9846);
or UO_719 (O_719,N_9946,N_9886);
nor UO_720 (O_720,N_9805,N_9956);
nand UO_721 (O_721,N_9970,N_9817);
and UO_722 (O_722,N_9888,N_9954);
and UO_723 (O_723,N_9985,N_9841);
nand UO_724 (O_724,N_9886,N_9932);
nor UO_725 (O_725,N_9945,N_9860);
and UO_726 (O_726,N_9943,N_9983);
nor UO_727 (O_727,N_9954,N_9808);
nor UO_728 (O_728,N_9983,N_9813);
or UO_729 (O_729,N_9937,N_9815);
nor UO_730 (O_730,N_9956,N_9962);
and UO_731 (O_731,N_9810,N_9945);
and UO_732 (O_732,N_9999,N_9886);
xnor UO_733 (O_733,N_9924,N_9911);
nand UO_734 (O_734,N_9817,N_9954);
nor UO_735 (O_735,N_9896,N_9914);
or UO_736 (O_736,N_9888,N_9838);
or UO_737 (O_737,N_9851,N_9915);
or UO_738 (O_738,N_9933,N_9930);
and UO_739 (O_739,N_9992,N_9983);
nand UO_740 (O_740,N_9823,N_9885);
nor UO_741 (O_741,N_9994,N_9998);
nor UO_742 (O_742,N_9967,N_9904);
or UO_743 (O_743,N_9995,N_9973);
xor UO_744 (O_744,N_9840,N_9904);
xnor UO_745 (O_745,N_9970,N_9882);
nand UO_746 (O_746,N_9891,N_9942);
and UO_747 (O_747,N_9960,N_9862);
and UO_748 (O_748,N_9802,N_9839);
or UO_749 (O_749,N_9896,N_9847);
or UO_750 (O_750,N_9814,N_9833);
nand UO_751 (O_751,N_9809,N_9921);
and UO_752 (O_752,N_9900,N_9809);
xnor UO_753 (O_753,N_9870,N_9878);
xnor UO_754 (O_754,N_9987,N_9889);
nor UO_755 (O_755,N_9964,N_9914);
xnor UO_756 (O_756,N_9952,N_9988);
or UO_757 (O_757,N_9915,N_9989);
nor UO_758 (O_758,N_9967,N_9955);
and UO_759 (O_759,N_9980,N_9956);
or UO_760 (O_760,N_9946,N_9917);
xnor UO_761 (O_761,N_9929,N_9847);
nand UO_762 (O_762,N_9813,N_9823);
nand UO_763 (O_763,N_9814,N_9840);
xor UO_764 (O_764,N_9853,N_9886);
or UO_765 (O_765,N_9835,N_9836);
nand UO_766 (O_766,N_9997,N_9950);
and UO_767 (O_767,N_9885,N_9965);
nand UO_768 (O_768,N_9967,N_9834);
nand UO_769 (O_769,N_9934,N_9920);
or UO_770 (O_770,N_9838,N_9837);
and UO_771 (O_771,N_9869,N_9844);
and UO_772 (O_772,N_9832,N_9894);
nand UO_773 (O_773,N_9804,N_9961);
and UO_774 (O_774,N_9822,N_9929);
nor UO_775 (O_775,N_9917,N_9943);
and UO_776 (O_776,N_9925,N_9961);
nand UO_777 (O_777,N_9811,N_9873);
and UO_778 (O_778,N_9918,N_9871);
xor UO_779 (O_779,N_9847,N_9931);
xnor UO_780 (O_780,N_9994,N_9975);
nand UO_781 (O_781,N_9920,N_9890);
and UO_782 (O_782,N_9823,N_9989);
or UO_783 (O_783,N_9805,N_9832);
nand UO_784 (O_784,N_9903,N_9802);
nand UO_785 (O_785,N_9909,N_9839);
nor UO_786 (O_786,N_9864,N_9999);
nand UO_787 (O_787,N_9940,N_9947);
xor UO_788 (O_788,N_9922,N_9938);
nor UO_789 (O_789,N_9888,N_9909);
and UO_790 (O_790,N_9849,N_9980);
xor UO_791 (O_791,N_9966,N_9845);
nand UO_792 (O_792,N_9904,N_9835);
nor UO_793 (O_793,N_9944,N_9903);
or UO_794 (O_794,N_9835,N_9842);
nand UO_795 (O_795,N_9886,N_9836);
xor UO_796 (O_796,N_9878,N_9937);
and UO_797 (O_797,N_9826,N_9943);
or UO_798 (O_798,N_9870,N_9860);
nand UO_799 (O_799,N_9913,N_9848);
nand UO_800 (O_800,N_9811,N_9872);
and UO_801 (O_801,N_9930,N_9836);
xor UO_802 (O_802,N_9900,N_9828);
xor UO_803 (O_803,N_9936,N_9919);
or UO_804 (O_804,N_9997,N_9813);
xnor UO_805 (O_805,N_9992,N_9979);
or UO_806 (O_806,N_9996,N_9999);
nand UO_807 (O_807,N_9953,N_9893);
xor UO_808 (O_808,N_9825,N_9950);
nor UO_809 (O_809,N_9866,N_9822);
nand UO_810 (O_810,N_9863,N_9834);
or UO_811 (O_811,N_9890,N_9897);
nor UO_812 (O_812,N_9932,N_9991);
and UO_813 (O_813,N_9968,N_9993);
nor UO_814 (O_814,N_9876,N_9942);
nor UO_815 (O_815,N_9948,N_9916);
nand UO_816 (O_816,N_9928,N_9985);
or UO_817 (O_817,N_9833,N_9954);
xor UO_818 (O_818,N_9821,N_9832);
and UO_819 (O_819,N_9887,N_9905);
nor UO_820 (O_820,N_9848,N_9800);
or UO_821 (O_821,N_9873,N_9942);
and UO_822 (O_822,N_9884,N_9867);
xor UO_823 (O_823,N_9989,N_9877);
or UO_824 (O_824,N_9975,N_9930);
xnor UO_825 (O_825,N_9804,N_9959);
or UO_826 (O_826,N_9929,N_9818);
xor UO_827 (O_827,N_9902,N_9994);
xnor UO_828 (O_828,N_9923,N_9900);
xor UO_829 (O_829,N_9830,N_9969);
or UO_830 (O_830,N_9974,N_9871);
nand UO_831 (O_831,N_9851,N_9816);
nand UO_832 (O_832,N_9846,N_9873);
and UO_833 (O_833,N_9910,N_9979);
nand UO_834 (O_834,N_9923,N_9991);
or UO_835 (O_835,N_9932,N_9978);
xor UO_836 (O_836,N_9944,N_9975);
nor UO_837 (O_837,N_9939,N_9999);
nor UO_838 (O_838,N_9986,N_9872);
and UO_839 (O_839,N_9982,N_9825);
or UO_840 (O_840,N_9846,N_9867);
and UO_841 (O_841,N_9968,N_9951);
nor UO_842 (O_842,N_9812,N_9871);
nand UO_843 (O_843,N_9915,N_9927);
nand UO_844 (O_844,N_9907,N_9992);
xor UO_845 (O_845,N_9870,N_9848);
or UO_846 (O_846,N_9930,N_9825);
xor UO_847 (O_847,N_9997,N_9927);
nand UO_848 (O_848,N_9933,N_9870);
nor UO_849 (O_849,N_9808,N_9829);
and UO_850 (O_850,N_9908,N_9855);
xor UO_851 (O_851,N_9911,N_9929);
or UO_852 (O_852,N_9866,N_9897);
xor UO_853 (O_853,N_9820,N_9800);
or UO_854 (O_854,N_9823,N_9825);
or UO_855 (O_855,N_9973,N_9989);
or UO_856 (O_856,N_9994,N_9933);
nand UO_857 (O_857,N_9931,N_9971);
xor UO_858 (O_858,N_9976,N_9913);
xor UO_859 (O_859,N_9896,N_9939);
xor UO_860 (O_860,N_9887,N_9842);
and UO_861 (O_861,N_9895,N_9879);
or UO_862 (O_862,N_9974,N_9945);
and UO_863 (O_863,N_9913,N_9803);
xnor UO_864 (O_864,N_9821,N_9813);
and UO_865 (O_865,N_9888,N_9978);
nand UO_866 (O_866,N_9815,N_9998);
nand UO_867 (O_867,N_9830,N_9994);
xnor UO_868 (O_868,N_9973,N_9872);
or UO_869 (O_869,N_9872,N_9983);
nor UO_870 (O_870,N_9952,N_9947);
and UO_871 (O_871,N_9854,N_9804);
or UO_872 (O_872,N_9981,N_9870);
and UO_873 (O_873,N_9964,N_9843);
xnor UO_874 (O_874,N_9874,N_9882);
nor UO_875 (O_875,N_9901,N_9914);
nor UO_876 (O_876,N_9873,N_9979);
and UO_877 (O_877,N_9919,N_9827);
nor UO_878 (O_878,N_9876,N_9923);
and UO_879 (O_879,N_9856,N_9897);
and UO_880 (O_880,N_9892,N_9971);
nor UO_881 (O_881,N_9826,N_9843);
or UO_882 (O_882,N_9884,N_9845);
or UO_883 (O_883,N_9919,N_9842);
nand UO_884 (O_884,N_9804,N_9860);
nor UO_885 (O_885,N_9858,N_9881);
and UO_886 (O_886,N_9831,N_9820);
nand UO_887 (O_887,N_9935,N_9849);
and UO_888 (O_888,N_9914,N_9980);
or UO_889 (O_889,N_9862,N_9908);
nand UO_890 (O_890,N_9979,N_9962);
nor UO_891 (O_891,N_9970,N_9908);
nor UO_892 (O_892,N_9801,N_9966);
nor UO_893 (O_893,N_9986,N_9875);
nor UO_894 (O_894,N_9923,N_9903);
nand UO_895 (O_895,N_9874,N_9923);
nand UO_896 (O_896,N_9953,N_9859);
nor UO_897 (O_897,N_9882,N_9897);
and UO_898 (O_898,N_9986,N_9980);
nand UO_899 (O_899,N_9873,N_9872);
nand UO_900 (O_900,N_9934,N_9974);
nor UO_901 (O_901,N_9907,N_9816);
nor UO_902 (O_902,N_9831,N_9922);
or UO_903 (O_903,N_9833,N_9906);
xnor UO_904 (O_904,N_9873,N_9945);
and UO_905 (O_905,N_9946,N_9811);
nand UO_906 (O_906,N_9843,N_9840);
nand UO_907 (O_907,N_9925,N_9972);
nand UO_908 (O_908,N_9905,N_9995);
or UO_909 (O_909,N_9834,N_9928);
xor UO_910 (O_910,N_9903,N_9897);
or UO_911 (O_911,N_9988,N_9966);
or UO_912 (O_912,N_9954,N_9977);
and UO_913 (O_913,N_9883,N_9936);
nor UO_914 (O_914,N_9832,N_9997);
nor UO_915 (O_915,N_9896,N_9838);
and UO_916 (O_916,N_9897,N_9921);
nand UO_917 (O_917,N_9924,N_9976);
or UO_918 (O_918,N_9976,N_9922);
and UO_919 (O_919,N_9891,N_9802);
nor UO_920 (O_920,N_9951,N_9898);
and UO_921 (O_921,N_9830,N_9829);
nand UO_922 (O_922,N_9959,N_9847);
nor UO_923 (O_923,N_9936,N_9856);
and UO_924 (O_924,N_9915,N_9868);
or UO_925 (O_925,N_9883,N_9958);
and UO_926 (O_926,N_9815,N_9981);
xor UO_927 (O_927,N_9876,N_9852);
nor UO_928 (O_928,N_9843,N_9941);
and UO_929 (O_929,N_9956,N_9827);
nor UO_930 (O_930,N_9860,N_9989);
or UO_931 (O_931,N_9832,N_9812);
and UO_932 (O_932,N_9861,N_9862);
and UO_933 (O_933,N_9977,N_9958);
nor UO_934 (O_934,N_9813,N_9810);
nand UO_935 (O_935,N_9827,N_9947);
and UO_936 (O_936,N_9886,N_9824);
nor UO_937 (O_937,N_9912,N_9904);
nor UO_938 (O_938,N_9937,N_9970);
and UO_939 (O_939,N_9982,N_9936);
or UO_940 (O_940,N_9992,N_9930);
and UO_941 (O_941,N_9909,N_9838);
nor UO_942 (O_942,N_9868,N_9897);
nor UO_943 (O_943,N_9958,N_9982);
or UO_944 (O_944,N_9812,N_9860);
nand UO_945 (O_945,N_9980,N_9809);
and UO_946 (O_946,N_9997,N_9847);
xor UO_947 (O_947,N_9992,N_9817);
xnor UO_948 (O_948,N_9800,N_9908);
xor UO_949 (O_949,N_9953,N_9913);
xor UO_950 (O_950,N_9826,N_9818);
and UO_951 (O_951,N_9808,N_9922);
nand UO_952 (O_952,N_9909,N_9821);
or UO_953 (O_953,N_9888,N_9999);
nand UO_954 (O_954,N_9827,N_9910);
xnor UO_955 (O_955,N_9975,N_9968);
and UO_956 (O_956,N_9848,N_9996);
and UO_957 (O_957,N_9824,N_9828);
and UO_958 (O_958,N_9919,N_9878);
or UO_959 (O_959,N_9817,N_9938);
and UO_960 (O_960,N_9935,N_9895);
or UO_961 (O_961,N_9976,N_9889);
nor UO_962 (O_962,N_9967,N_9979);
nor UO_963 (O_963,N_9870,N_9980);
or UO_964 (O_964,N_9941,N_9981);
nor UO_965 (O_965,N_9883,N_9874);
xor UO_966 (O_966,N_9876,N_9849);
nor UO_967 (O_967,N_9906,N_9983);
or UO_968 (O_968,N_9821,N_9994);
nor UO_969 (O_969,N_9858,N_9925);
or UO_970 (O_970,N_9960,N_9991);
nor UO_971 (O_971,N_9993,N_9891);
nor UO_972 (O_972,N_9852,N_9984);
nand UO_973 (O_973,N_9815,N_9933);
and UO_974 (O_974,N_9816,N_9964);
nor UO_975 (O_975,N_9861,N_9925);
nand UO_976 (O_976,N_9874,N_9957);
nand UO_977 (O_977,N_9844,N_9815);
and UO_978 (O_978,N_9970,N_9828);
xor UO_979 (O_979,N_9953,N_9925);
nand UO_980 (O_980,N_9866,N_9925);
and UO_981 (O_981,N_9925,N_9915);
nand UO_982 (O_982,N_9980,N_9822);
xor UO_983 (O_983,N_9815,N_9886);
and UO_984 (O_984,N_9961,N_9946);
nand UO_985 (O_985,N_9968,N_9978);
and UO_986 (O_986,N_9926,N_9958);
or UO_987 (O_987,N_9856,N_9876);
nor UO_988 (O_988,N_9815,N_9934);
and UO_989 (O_989,N_9820,N_9986);
or UO_990 (O_990,N_9912,N_9825);
nand UO_991 (O_991,N_9817,N_9912);
and UO_992 (O_992,N_9929,N_9850);
nand UO_993 (O_993,N_9992,N_9953);
or UO_994 (O_994,N_9946,N_9907);
nand UO_995 (O_995,N_9884,N_9998);
or UO_996 (O_996,N_9851,N_9801);
or UO_997 (O_997,N_9846,N_9994);
nand UO_998 (O_998,N_9850,N_9818);
nand UO_999 (O_999,N_9965,N_9905);
nor UO_1000 (O_1000,N_9878,N_9924);
nor UO_1001 (O_1001,N_9899,N_9852);
nor UO_1002 (O_1002,N_9955,N_9844);
nor UO_1003 (O_1003,N_9998,N_9917);
or UO_1004 (O_1004,N_9847,N_9986);
nor UO_1005 (O_1005,N_9949,N_9836);
and UO_1006 (O_1006,N_9990,N_9960);
or UO_1007 (O_1007,N_9823,N_9832);
and UO_1008 (O_1008,N_9899,N_9933);
nand UO_1009 (O_1009,N_9829,N_9868);
nor UO_1010 (O_1010,N_9818,N_9807);
nor UO_1011 (O_1011,N_9976,N_9811);
or UO_1012 (O_1012,N_9854,N_9832);
xor UO_1013 (O_1013,N_9900,N_9987);
nor UO_1014 (O_1014,N_9881,N_9892);
or UO_1015 (O_1015,N_9807,N_9989);
nand UO_1016 (O_1016,N_9938,N_9905);
nand UO_1017 (O_1017,N_9964,N_9976);
and UO_1018 (O_1018,N_9820,N_9978);
nand UO_1019 (O_1019,N_9948,N_9904);
and UO_1020 (O_1020,N_9891,N_9937);
and UO_1021 (O_1021,N_9851,N_9906);
or UO_1022 (O_1022,N_9966,N_9810);
nand UO_1023 (O_1023,N_9990,N_9983);
and UO_1024 (O_1024,N_9997,N_9939);
xor UO_1025 (O_1025,N_9970,N_9918);
or UO_1026 (O_1026,N_9994,N_9995);
nor UO_1027 (O_1027,N_9934,N_9936);
xnor UO_1028 (O_1028,N_9830,N_9900);
or UO_1029 (O_1029,N_9881,N_9931);
and UO_1030 (O_1030,N_9909,N_9928);
or UO_1031 (O_1031,N_9917,N_9866);
xnor UO_1032 (O_1032,N_9952,N_9829);
xnor UO_1033 (O_1033,N_9909,N_9879);
or UO_1034 (O_1034,N_9824,N_9947);
nor UO_1035 (O_1035,N_9885,N_9933);
xnor UO_1036 (O_1036,N_9914,N_9822);
and UO_1037 (O_1037,N_9900,N_9840);
nor UO_1038 (O_1038,N_9819,N_9808);
or UO_1039 (O_1039,N_9887,N_9955);
or UO_1040 (O_1040,N_9867,N_9893);
or UO_1041 (O_1041,N_9846,N_9970);
xnor UO_1042 (O_1042,N_9858,N_9853);
or UO_1043 (O_1043,N_9862,N_9875);
or UO_1044 (O_1044,N_9992,N_9987);
nor UO_1045 (O_1045,N_9973,N_9943);
and UO_1046 (O_1046,N_9824,N_9994);
xnor UO_1047 (O_1047,N_9984,N_9903);
and UO_1048 (O_1048,N_9860,N_9898);
and UO_1049 (O_1049,N_9992,N_9815);
nand UO_1050 (O_1050,N_9856,N_9964);
nand UO_1051 (O_1051,N_9903,N_9819);
or UO_1052 (O_1052,N_9883,N_9800);
and UO_1053 (O_1053,N_9957,N_9990);
nand UO_1054 (O_1054,N_9856,N_9981);
nor UO_1055 (O_1055,N_9952,N_9989);
nor UO_1056 (O_1056,N_9964,N_9987);
nand UO_1057 (O_1057,N_9988,N_9959);
and UO_1058 (O_1058,N_9828,N_9863);
nor UO_1059 (O_1059,N_9973,N_9883);
and UO_1060 (O_1060,N_9898,N_9956);
nand UO_1061 (O_1061,N_9982,N_9887);
and UO_1062 (O_1062,N_9931,N_9814);
nor UO_1063 (O_1063,N_9859,N_9837);
xnor UO_1064 (O_1064,N_9906,N_9813);
and UO_1065 (O_1065,N_9958,N_9804);
nor UO_1066 (O_1066,N_9993,N_9825);
nor UO_1067 (O_1067,N_9899,N_9880);
nor UO_1068 (O_1068,N_9845,N_9864);
or UO_1069 (O_1069,N_9995,N_9853);
or UO_1070 (O_1070,N_9848,N_9903);
nor UO_1071 (O_1071,N_9908,N_9922);
nor UO_1072 (O_1072,N_9877,N_9834);
and UO_1073 (O_1073,N_9943,N_9868);
nand UO_1074 (O_1074,N_9816,N_9952);
and UO_1075 (O_1075,N_9825,N_9996);
or UO_1076 (O_1076,N_9809,N_9964);
and UO_1077 (O_1077,N_9888,N_9921);
nor UO_1078 (O_1078,N_9937,N_9892);
nand UO_1079 (O_1079,N_9928,N_9984);
or UO_1080 (O_1080,N_9828,N_9809);
nand UO_1081 (O_1081,N_9840,N_9838);
nor UO_1082 (O_1082,N_9802,N_9917);
and UO_1083 (O_1083,N_9883,N_9954);
xnor UO_1084 (O_1084,N_9806,N_9908);
or UO_1085 (O_1085,N_9930,N_9880);
xor UO_1086 (O_1086,N_9838,N_9858);
or UO_1087 (O_1087,N_9913,N_9840);
nand UO_1088 (O_1088,N_9868,N_9986);
or UO_1089 (O_1089,N_9969,N_9998);
xor UO_1090 (O_1090,N_9855,N_9927);
nor UO_1091 (O_1091,N_9850,N_9944);
nor UO_1092 (O_1092,N_9802,N_9925);
or UO_1093 (O_1093,N_9818,N_9952);
or UO_1094 (O_1094,N_9981,N_9825);
nand UO_1095 (O_1095,N_9942,N_9811);
or UO_1096 (O_1096,N_9920,N_9976);
or UO_1097 (O_1097,N_9974,N_9972);
or UO_1098 (O_1098,N_9816,N_9837);
and UO_1099 (O_1099,N_9998,N_9837);
nand UO_1100 (O_1100,N_9842,N_9811);
nand UO_1101 (O_1101,N_9847,N_9835);
or UO_1102 (O_1102,N_9885,N_9869);
nor UO_1103 (O_1103,N_9986,N_9928);
or UO_1104 (O_1104,N_9987,N_9962);
nor UO_1105 (O_1105,N_9956,N_9834);
or UO_1106 (O_1106,N_9971,N_9883);
nand UO_1107 (O_1107,N_9958,N_9852);
nor UO_1108 (O_1108,N_9981,N_9847);
nand UO_1109 (O_1109,N_9832,N_9943);
or UO_1110 (O_1110,N_9812,N_9965);
nand UO_1111 (O_1111,N_9842,N_9817);
nand UO_1112 (O_1112,N_9964,N_9807);
and UO_1113 (O_1113,N_9849,N_9878);
nand UO_1114 (O_1114,N_9972,N_9992);
xnor UO_1115 (O_1115,N_9834,N_9883);
or UO_1116 (O_1116,N_9993,N_9875);
nor UO_1117 (O_1117,N_9953,N_9831);
or UO_1118 (O_1118,N_9930,N_9934);
nor UO_1119 (O_1119,N_9872,N_9890);
nor UO_1120 (O_1120,N_9921,N_9857);
nand UO_1121 (O_1121,N_9829,N_9995);
and UO_1122 (O_1122,N_9938,N_9844);
nand UO_1123 (O_1123,N_9852,N_9934);
and UO_1124 (O_1124,N_9833,N_9982);
nor UO_1125 (O_1125,N_9810,N_9845);
nor UO_1126 (O_1126,N_9915,N_9862);
nor UO_1127 (O_1127,N_9832,N_9801);
nor UO_1128 (O_1128,N_9916,N_9860);
and UO_1129 (O_1129,N_9891,N_9900);
nor UO_1130 (O_1130,N_9860,N_9822);
nor UO_1131 (O_1131,N_9873,N_9886);
or UO_1132 (O_1132,N_9943,N_9934);
xor UO_1133 (O_1133,N_9881,N_9840);
xor UO_1134 (O_1134,N_9930,N_9961);
xor UO_1135 (O_1135,N_9919,N_9933);
nand UO_1136 (O_1136,N_9829,N_9929);
or UO_1137 (O_1137,N_9977,N_9959);
xor UO_1138 (O_1138,N_9811,N_9827);
and UO_1139 (O_1139,N_9850,N_9817);
and UO_1140 (O_1140,N_9803,N_9982);
xnor UO_1141 (O_1141,N_9920,N_9886);
nand UO_1142 (O_1142,N_9972,N_9942);
xnor UO_1143 (O_1143,N_9807,N_9910);
or UO_1144 (O_1144,N_9917,N_9919);
nor UO_1145 (O_1145,N_9811,N_9951);
nand UO_1146 (O_1146,N_9834,N_9913);
xor UO_1147 (O_1147,N_9940,N_9826);
or UO_1148 (O_1148,N_9882,N_9865);
xnor UO_1149 (O_1149,N_9885,N_9982);
and UO_1150 (O_1150,N_9947,N_9976);
and UO_1151 (O_1151,N_9849,N_9807);
or UO_1152 (O_1152,N_9801,N_9945);
xnor UO_1153 (O_1153,N_9824,N_9821);
xnor UO_1154 (O_1154,N_9887,N_9883);
and UO_1155 (O_1155,N_9845,N_9883);
nand UO_1156 (O_1156,N_9877,N_9839);
nand UO_1157 (O_1157,N_9960,N_9944);
xor UO_1158 (O_1158,N_9987,N_9985);
xnor UO_1159 (O_1159,N_9885,N_9882);
and UO_1160 (O_1160,N_9903,N_9963);
or UO_1161 (O_1161,N_9972,N_9989);
and UO_1162 (O_1162,N_9960,N_9880);
and UO_1163 (O_1163,N_9948,N_9991);
nand UO_1164 (O_1164,N_9842,N_9894);
and UO_1165 (O_1165,N_9953,N_9900);
and UO_1166 (O_1166,N_9941,N_9825);
or UO_1167 (O_1167,N_9919,N_9939);
nor UO_1168 (O_1168,N_9806,N_9903);
and UO_1169 (O_1169,N_9845,N_9906);
nand UO_1170 (O_1170,N_9967,N_9837);
or UO_1171 (O_1171,N_9883,N_9979);
and UO_1172 (O_1172,N_9811,N_9823);
nor UO_1173 (O_1173,N_9925,N_9957);
nand UO_1174 (O_1174,N_9938,N_9918);
nand UO_1175 (O_1175,N_9953,N_9828);
nor UO_1176 (O_1176,N_9922,N_9968);
nor UO_1177 (O_1177,N_9847,N_9970);
and UO_1178 (O_1178,N_9859,N_9923);
nor UO_1179 (O_1179,N_9854,N_9993);
xnor UO_1180 (O_1180,N_9828,N_9938);
or UO_1181 (O_1181,N_9902,N_9906);
or UO_1182 (O_1182,N_9906,N_9975);
and UO_1183 (O_1183,N_9822,N_9890);
nor UO_1184 (O_1184,N_9812,N_9841);
nor UO_1185 (O_1185,N_9820,N_9832);
or UO_1186 (O_1186,N_9989,N_9814);
nand UO_1187 (O_1187,N_9874,N_9848);
nand UO_1188 (O_1188,N_9888,N_9989);
nor UO_1189 (O_1189,N_9900,N_9972);
nand UO_1190 (O_1190,N_9894,N_9946);
xnor UO_1191 (O_1191,N_9998,N_9964);
and UO_1192 (O_1192,N_9974,N_9904);
or UO_1193 (O_1193,N_9845,N_9932);
nand UO_1194 (O_1194,N_9962,N_9977);
xor UO_1195 (O_1195,N_9866,N_9895);
and UO_1196 (O_1196,N_9953,N_9820);
or UO_1197 (O_1197,N_9989,N_9903);
or UO_1198 (O_1198,N_9953,N_9823);
xor UO_1199 (O_1199,N_9912,N_9857);
xnor UO_1200 (O_1200,N_9839,N_9906);
or UO_1201 (O_1201,N_9914,N_9985);
xor UO_1202 (O_1202,N_9878,N_9825);
nand UO_1203 (O_1203,N_9932,N_9968);
or UO_1204 (O_1204,N_9851,N_9970);
nand UO_1205 (O_1205,N_9857,N_9974);
and UO_1206 (O_1206,N_9996,N_9898);
nand UO_1207 (O_1207,N_9940,N_9893);
or UO_1208 (O_1208,N_9920,N_9839);
xor UO_1209 (O_1209,N_9809,N_9849);
or UO_1210 (O_1210,N_9916,N_9931);
xor UO_1211 (O_1211,N_9961,N_9926);
and UO_1212 (O_1212,N_9825,N_9850);
nand UO_1213 (O_1213,N_9927,N_9810);
xnor UO_1214 (O_1214,N_9823,N_9984);
xor UO_1215 (O_1215,N_9902,N_9978);
nor UO_1216 (O_1216,N_9822,N_9818);
and UO_1217 (O_1217,N_9961,N_9975);
nand UO_1218 (O_1218,N_9855,N_9841);
xor UO_1219 (O_1219,N_9936,N_9880);
xnor UO_1220 (O_1220,N_9937,N_9886);
and UO_1221 (O_1221,N_9988,N_9941);
nand UO_1222 (O_1222,N_9851,N_9847);
xor UO_1223 (O_1223,N_9911,N_9857);
nor UO_1224 (O_1224,N_9978,N_9931);
and UO_1225 (O_1225,N_9937,N_9964);
nand UO_1226 (O_1226,N_9886,N_9904);
xnor UO_1227 (O_1227,N_9836,N_9917);
and UO_1228 (O_1228,N_9879,N_9834);
and UO_1229 (O_1229,N_9975,N_9872);
xnor UO_1230 (O_1230,N_9823,N_9920);
or UO_1231 (O_1231,N_9977,N_9981);
and UO_1232 (O_1232,N_9992,N_9838);
nor UO_1233 (O_1233,N_9960,N_9997);
xor UO_1234 (O_1234,N_9900,N_9927);
nand UO_1235 (O_1235,N_9881,N_9898);
nand UO_1236 (O_1236,N_9891,N_9807);
and UO_1237 (O_1237,N_9956,N_9845);
xor UO_1238 (O_1238,N_9800,N_9994);
and UO_1239 (O_1239,N_9960,N_9872);
xnor UO_1240 (O_1240,N_9956,N_9894);
and UO_1241 (O_1241,N_9801,N_9903);
xnor UO_1242 (O_1242,N_9940,N_9849);
and UO_1243 (O_1243,N_9809,N_9841);
xor UO_1244 (O_1244,N_9843,N_9968);
and UO_1245 (O_1245,N_9998,N_9834);
and UO_1246 (O_1246,N_9894,N_9987);
nor UO_1247 (O_1247,N_9965,N_9981);
nand UO_1248 (O_1248,N_9849,N_9817);
xor UO_1249 (O_1249,N_9945,N_9895);
nor UO_1250 (O_1250,N_9838,N_9857);
nand UO_1251 (O_1251,N_9906,N_9853);
nand UO_1252 (O_1252,N_9999,N_9978);
or UO_1253 (O_1253,N_9825,N_9861);
and UO_1254 (O_1254,N_9875,N_9822);
nor UO_1255 (O_1255,N_9893,N_9892);
nand UO_1256 (O_1256,N_9812,N_9877);
nand UO_1257 (O_1257,N_9866,N_9903);
nor UO_1258 (O_1258,N_9914,N_9972);
xor UO_1259 (O_1259,N_9836,N_9814);
or UO_1260 (O_1260,N_9915,N_9870);
nor UO_1261 (O_1261,N_9977,N_9802);
nand UO_1262 (O_1262,N_9966,N_9832);
or UO_1263 (O_1263,N_9955,N_9995);
nand UO_1264 (O_1264,N_9911,N_9936);
xor UO_1265 (O_1265,N_9989,N_9833);
nor UO_1266 (O_1266,N_9949,N_9962);
and UO_1267 (O_1267,N_9965,N_9893);
nand UO_1268 (O_1268,N_9814,N_9999);
nor UO_1269 (O_1269,N_9891,N_9980);
nand UO_1270 (O_1270,N_9827,N_9825);
nor UO_1271 (O_1271,N_9887,N_9927);
nand UO_1272 (O_1272,N_9868,N_9809);
nand UO_1273 (O_1273,N_9833,N_9925);
nand UO_1274 (O_1274,N_9863,N_9870);
nor UO_1275 (O_1275,N_9964,N_9993);
or UO_1276 (O_1276,N_9839,N_9852);
nor UO_1277 (O_1277,N_9938,N_9802);
or UO_1278 (O_1278,N_9913,N_9891);
and UO_1279 (O_1279,N_9982,N_9813);
nor UO_1280 (O_1280,N_9803,N_9942);
nor UO_1281 (O_1281,N_9843,N_9802);
nand UO_1282 (O_1282,N_9928,N_9882);
nand UO_1283 (O_1283,N_9905,N_9923);
and UO_1284 (O_1284,N_9800,N_9990);
or UO_1285 (O_1285,N_9875,N_9991);
nor UO_1286 (O_1286,N_9945,N_9971);
nand UO_1287 (O_1287,N_9855,N_9868);
xor UO_1288 (O_1288,N_9810,N_9973);
xnor UO_1289 (O_1289,N_9964,N_9830);
and UO_1290 (O_1290,N_9982,N_9983);
nand UO_1291 (O_1291,N_9951,N_9813);
xnor UO_1292 (O_1292,N_9883,N_9871);
nand UO_1293 (O_1293,N_9998,N_9973);
nor UO_1294 (O_1294,N_9922,N_9956);
and UO_1295 (O_1295,N_9825,N_9896);
nor UO_1296 (O_1296,N_9835,N_9838);
and UO_1297 (O_1297,N_9989,N_9934);
nand UO_1298 (O_1298,N_9838,N_9859);
nand UO_1299 (O_1299,N_9938,N_9959);
and UO_1300 (O_1300,N_9959,N_9937);
nand UO_1301 (O_1301,N_9822,N_9809);
xnor UO_1302 (O_1302,N_9867,N_9939);
or UO_1303 (O_1303,N_9828,N_9813);
xor UO_1304 (O_1304,N_9821,N_9900);
xor UO_1305 (O_1305,N_9929,N_9975);
and UO_1306 (O_1306,N_9988,N_9999);
xor UO_1307 (O_1307,N_9807,N_9926);
or UO_1308 (O_1308,N_9949,N_9905);
xnor UO_1309 (O_1309,N_9834,N_9810);
and UO_1310 (O_1310,N_9931,N_9968);
nand UO_1311 (O_1311,N_9930,N_9916);
and UO_1312 (O_1312,N_9837,N_9938);
xnor UO_1313 (O_1313,N_9919,N_9823);
nor UO_1314 (O_1314,N_9949,N_9999);
xor UO_1315 (O_1315,N_9975,N_9893);
and UO_1316 (O_1316,N_9811,N_9961);
xnor UO_1317 (O_1317,N_9949,N_9994);
and UO_1318 (O_1318,N_9843,N_9998);
and UO_1319 (O_1319,N_9811,N_9910);
or UO_1320 (O_1320,N_9879,N_9873);
nor UO_1321 (O_1321,N_9865,N_9908);
nor UO_1322 (O_1322,N_9960,N_9935);
nand UO_1323 (O_1323,N_9858,N_9993);
nor UO_1324 (O_1324,N_9839,N_9828);
or UO_1325 (O_1325,N_9992,N_9986);
nor UO_1326 (O_1326,N_9810,N_9823);
nor UO_1327 (O_1327,N_9977,N_9963);
nand UO_1328 (O_1328,N_9919,N_9928);
and UO_1329 (O_1329,N_9987,N_9997);
xnor UO_1330 (O_1330,N_9916,N_9867);
xnor UO_1331 (O_1331,N_9910,N_9858);
xor UO_1332 (O_1332,N_9987,N_9805);
nand UO_1333 (O_1333,N_9953,N_9845);
nor UO_1334 (O_1334,N_9818,N_9908);
nor UO_1335 (O_1335,N_9904,N_9810);
xor UO_1336 (O_1336,N_9872,N_9996);
or UO_1337 (O_1337,N_9927,N_9860);
or UO_1338 (O_1338,N_9950,N_9954);
nor UO_1339 (O_1339,N_9832,N_9847);
nor UO_1340 (O_1340,N_9931,N_9906);
and UO_1341 (O_1341,N_9845,N_9836);
or UO_1342 (O_1342,N_9873,N_9930);
and UO_1343 (O_1343,N_9870,N_9809);
and UO_1344 (O_1344,N_9963,N_9818);
xnor UO_1345 (O_1345,N_9805,N_9986);
and UO_1346 (O_1346,N_9976,N_9895);
xnor UO_1347 (O_1347,N_9888,N_9922);
or UO_1348 (O_1348,N_9880,N_9891);
and UO_1349 (O_1349,N_9928,N_9995);
or UO_1350 (O_1350,N_9831,N_9994);
xor UO_1351 (O_1351,N_9870,N_9849);
nand UO_1352 (O_1352,N_9853,N_9957);
or UO_1353 (O_1353,N_9880,N_9955);
nand UO_1354 (O_1354,N_9861,N_9904);
or UO_1355 (O_1355,N_9882,N_9991);
nor UO_1356 (O_1356,N_9807,N_9919);
xor UO_1357 (O_1357,N_9855,N_9859);
nor UO_1358 (O_1358,N_9938,N_9953);
xor UO_1359 (O_1359,N_9848,N_9944);
and UO_1360 (O_1360,N_9835,N_9866);
nand UO_1361 (O_1361,N_9994,N_9809);
nand UO_1362 (O_1362,N_9977,N_9828);
or UO_1363 (O_1363,N_9890,N_9952);
xnor UO_1364 (O_1364,N_9892,N_9829);
nor UO_1365 (O_1365,N_9842,N_9854);
or UO_1366 (O_1366,N_9842,N_9863);
xnor UO_1367 (O_1367,N_9819,N_9968);
nor UO_1368 (O_1368,N_9897,N_9902);
nor UO_1369 (O_1369,N_9849,N_9815);
or UO_1370 (O_1370,N_9956,N_9989);
and UO_1371 (O_1371,N_9872,N_9943);
nand UO_1372 (O_1372,N_9952,N_9847);
and UO_1373 (O_1373,N_9809,N_9950);
xnor UO_1374 (O_1374,N_9849,N_9958);
or UO_1375 (O_1375,N_9807,N_9925);
or UO_1376 (O_1376,N_9816,N_9975);
or UO_1377 (O_1377,N_9899,N_9875);
and UO_1378 (O_1378,N_9853,N_9846);
nor UO_1379 (O_1379,N_9802,N_9806);
or UO_1380 (O_1380,N_9921,N_9822);
nor UO_1381 (O_1381,N_9869,N_9962);
xnor UO_1382 (O_1382,N_9814,N_9854);
nand UO_1383 (O_1383,N_9911,N_9923);
nand UO_1384 (O_1384,N_9891,N_9861);
xor UO_1385 (O_1385,N_9862,N_9871);
xor UO_1386 (O_1386,N_9890,N_9887);
or UO_1387 (O_1387,N_9853,N_9934);
nand UO_1388 (O_1388,N_9808,N_9906);
xnor UO_1389 (O_1389,N_9812,N_9837);
nor UO_1390 (O_1390,N_9893,N_9939);
nand UO_1391 (O_1391,N_9949,N_9834);
nor UO_1392 (O_1392,N_9836,N_9881);
and UO_1393 (O_1393,N_9842,N_9847);
and UO_1394 (O_1394,N_9808,N_9945);
nor UO_1395 (O_1395,N_9905,N_9913);
and UO_1396 (O_1396,N_9807,N_9815);
nor UO_1397 (O_1397,N_9846,N_9931);
nor UO_1398 (O_1398,N_9801,N_9829);
or UO_1399 (O_1399,N_9906,N_9850);
or UO_1400 (O_1400,N_9909,N_9830);
and UO_1401 (O_1401,N_9937,N_9967);
nor UO_1402 (O_1402,N_9961,N_9865);
or UO_1403 (O_1403,N_9957,N_9936);
and UO_1404 (O_1404,N_9953,N_9931);
xor UO_1405 (O_1405,N_9886,N_9921);
or UO_1406 (O_1406,N_9824,N_9873);
nor UO_1407 (O_1407,N_9978,N_9886);
nor UO_1408 (O_1408,N_9840,N_9901);
nand UO_1409 (O_1409,N_9924,N_9980);
nand UO_1410 (O_1410,N_9915,N_9907);
xor UO_1411 (O_1411,N_9912,N_9959);
xor UO_1412 (O_1412,N_9841,N_9819);
and UO_1413 (O_1413,N_9832,N_9983);
or UO_1414 (O_1414,N_9808,N_9803);
nor UO_1415 (O_1415,N_9914,N_9967);
nand UO_1416 (O_1416,N_9855,N_9809);
nand UO_1417 (O_1417,N_9862,N_9839);
xor UO_1418 (O_1418,N_9905,N_9967);
xor UO_1419 (O_1419,N_9882,N_9929);
and UO_1420 (O_1420,N_9892,N_9873);
xor UO_1421 (O_1421,N_9893,N_9850);
xor UO_1422 (O_1422,N_9916,N_9940);
nor UO_1423 (O_1423,N_9948,N_9865);
nor UO_1424 (O_1424,N_9809,N_9933);
or UO_1425 (O_1425,N_9953,N_9903);
and UO_1426 (O_1426,N_9921,N_9875);
and UO_1427 (O_1427,N_9967,N_9869);
nand UO_1428 (O_1428,N_9957,N_9847);
xor UO_1429 (O_1429,N_9944,N_9958);
or UO_1430 (O_1430,N_9843,N_9961);
and UO_1431 (O_1431,N_9934,N_9841);
nand UO_1432 (O_1432,N_9991,N_9817);
nor UO_1433 (O_1433,N_9838,N_9864);
nor UO_1434 (O_1434,N_9828,N_9950);
or UO_1435 (O_1435,N_9832,N_9875);
nand UO_1436 (O_1436,N_9901,N_9823);
nand UO_1437 (O_1437,N_9817,N_9893);
nand UO_1438 (O_1438,N_9987,N_9981);
and UO_1439 (O_1439,N_9931,N_9893);
nor UO_1440 (O_1440,N_9883,N_9843);
or UO_1441 (O_1441,N_9921,N_9832);
nand UO_1442 (O_1442,N_9977,N_9897);
or UO_1443 (O_1443,N_9904,N_9845);
or UO_1444 (O_1444,N_9838,N_9872);
xnor UO_1445 (O_1445,N_9840,N_9833);
nor UO_1446 (O_1446,N_9976,N_9876);
xnor UO_1447 (O_1447,N_9991,N_9871);
nor UO_1448 (O_1448,N_9949,N_9979);
nand UO_1449 (O_1449,N_9978,N_9860);
nand UO_1450 (O_1450,N_9921,N_9830);
nand UO_1451 (O_1451,N_9911,N_9974);
and UO_1452 (O_1452,N_9919,N_9948);
or UO_1453 (O_1453,N_9881,N_9920);
xor UO_1454 (O_1454,N_9825,N_9927);
and UO_1455 (O_1455,N_9986,N_9958);
nor UO_1456 (O_1456,N_9938,N_9995);
or UO_1457 (O_1457,N_9972,N_9967);
or UO_1458 (O_1458,N_9835,N_9876);
nand UO_1459 (O_1459,N_9848,N_9869);
or UO_1460 (O_1460,N_9889,N_9915);
nand UO_1461 (O_1461,N_9812,N_9938);
nor UO_1462 (O_1462,N_9917,N_9823);
xor UO_1463 (O_1463,N_9897,N_9976);
xnor UO_1464 (O_1464,N_9917,N_9833);
nand UO_1465 (O_1465,N_9807,N_9805);
and UO_1466 (O_1466,N_9837,N_9979);
or UO_1467 (O_1467,N_9978,N_9901);
nand UO_1468 (O_1468,N_9984,N_9848);
xor UO_1469 (O_1469,N_9855,N_9850);
and UO_1470 (O_1470,N_9818,N_9986);
and UO_1471 (O_1471,N_9854,N_9958);
or UO_1472 (O_1472,N_9874,N_9800);
xnor UO_1473 (O_1473,N_9960,N_9959);
xor UO_1474 (O_1474,N_9918,N_9876);
nand UO_1475 (O_1475,N_9945,N_9892);
or UO_1476 (O_1476,N_9852,N_9926);
and UO_1477 (O_1477,N_9982,N_9829);
nand UO_1478 (O_1478,N_9898,N_9855);
or UO_1479 (O_1479,N_9912,N_9909);
nand UO_1480 (O_1480,N_9911,N_9820);
xnor UO_1481 (O_1481,N_9928,N_9884);
nor UO_1482 (O_1482,N_9906,N_9827);
nor UO_1483 (O_1483,N_9947,N_9979);
nor UO_1484 (O_1484,N_9875,N_9841);
and UO_1485 (O_1485,N_9863,N_9886);
nor UO_1486 (O_1486,N_9839,N_9992);
xor UO_1487 (O_1487,N_9936,N_9809);
nand UO_1488 (O_1488,N_9890,N_9816);
or UO_1489 (O_1489,N_9965,N_9822);
nor UO_1490 (O_1490,N_9847,N_9880);
nor UO_1491 (O_1491,N_9997,N_9853);
or UO_1492 (O_1492,N_9810,N_9856);
nand UO_1493 (O_1493,N_9999,N_9922);
xnor UO_1494 (O_1494,N_9861,N_9976);
or UO_1495 (O_1495,N_9938,N_9878);
xnor UO_1496 (O_1496,N_9922,N_9862);
xnor UO_1497 (O_1497,N_9837,N_9903);
nand UO_1498 (O_1498,N_9820,N_9807);
and UO_1499 (O_1499,N_9920,N_9904);
endmodule