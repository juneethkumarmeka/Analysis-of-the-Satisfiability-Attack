module basic_500_3000_500_50_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_237,In_176);
nand U1 (N_1,In_457,In_443);
or U2 (N_2,In_140,In_487);
nand U3 (N_3,In_298,In_67);
nor U4 (N_4,In_185,In_432);
and U5 (N_5,In_1,In_453);
or U6 (N_6,In_472,In_198);
and U7 (N_7,In_106,In_256);
nand U8 (N_8,In_409,In_143);
or U9 (N_9,In_440,In_356);
xnor U10 (N_10,In_192,In_167);
or U11 (N_11,In_184,In_32);
nor U12 (N_12,In_364,In_423);
xor U13 (N_13,In_310,In_374);
or U14 (N_14,In_29,In_157);
nand U15 (N_15,In_244,In_53);
or U16 (N_16,In_387,In_332);
nor U17 (N_17,In_40,In_367);
or U18 (N_18,In_324,In_64);
xor U19 (N_19,In_58,In_283);
nand U20 (N_20,In_411,In_18);
or U21 (N_21,In_236,In_100);
nand U22 (N_22,In_149,In_249);
nand U23 (N_23,In_52,In_109);
xor U24 (N_24,In_57,In_240);
nor U25 (N_25,In_144,In_10);
nand U26 (N_26,In_59,In_239);
nand U27 (N_27,In_172,In_295);
and U28 (N_28,In_320,In_258);
nand U29 (N_29,In_325,In_415);
nor U30 (N_30,In_391,In_372);
xor U31 (N_31,In_86,In_70);
nand U32 (N_32,In_75,In_102);
or U33 (N_33,In_322,In_107);
and U34 (N_34,In_412,In_476);
or U35 (N_35,In_279,In_395);
nand U36 (N_36,In_284,In_273);
xnor U37 (N_37,In_403,In_229);
and U38 (N_38,In_141,In_68);
or U39 (N_39,In_19,In_0);
nand U40 (N_40,In_301,In_282);
nand U41 (N_41,In_478,In_93);
and U42 (N_42,In_352,In_340);
or U43 (N_43,In_145,In_254);
or U44 (N_44,In_365,In_385);
or U45 (N_45,In_116,In_264);
or U46 (N_46,In_309,In_71);
or U47 (N_47,In_490,In_384);
or U48 (N_48,In_233,In_499);
xnor U49 (N_49,In_307,In_248);
nand U50 (N_50,In_416,In_47);
nand U51 (N_51,In_326,In_419);
nor U52 (N_52,In_246,In_481);
or U53 (N_53,In_261,In_111);
nand U54 (N_54,In_468,In_306);
nor U55 (N_55,In_427,In_35);
or U56 (N_56,In_96,In_190);
nor U57 (N_57,In_91,In_422);
nand U58 (N_58,In_55,In_54);
xor U59 (N_59,In_438,In_449);
nand U60 (N_60,In_245,In_327);
xor U61 (N_61,In_413,In_117);
and U62 (N_62,In_424,In_114);
or U63 (N_63,N_40,In_80);
and U64 (N_64,In_253,In_483);
nand U65 (N_65,N_17,In_497);
and U66 (N_66,In_134,In_473);
xor U67 (N_67,In_436,In_5);
xnor U68 (N_68,In_126,In_381);
xor U69 (N_69,In_397,In_66);
and U70 (N_70,N_9,In_337);
nor U71 (N_71,In_353,In_4);
and U72 (N_72,In_418,In_90);
xor U73 (N_73,In_269,In_130);
nand U74 (N_74,In_101,In_450);
nand U75 (N_75,In_146,In_189);
nand U76 (N_76,In_319,N_15);
and U77 (N_77,N_8,In_376);
and U78 (N_78,In_44,In_88);
nand U79 (N_79,In_348,In_294);
and U80 (N_80,In_179,In_346);
or U81 (N_81,In_17,In_458);
and U82 (N_82,In_203,In_159);
nor U83 (N_83,In_426,In_128);
xnor U84 (N_84,In_170,In_97);
and U85 (N_85,N_7,N_54);
xnor U86 (N_86,N_38,In_160);
nand U87 (N_87,In_286,In_480);
and U88 (N_88,In_123,In_370);
nand U89 (N_89,In_386,In_194);
xor U90 (N_90,In_217,In_69);
xnor U91 (N_91,In_489,In_461);
or U92 (N_92,In_414,In_43);
nand U93 (N_93,In_174,In_357);
xnor U94 (N_94,In_323,In_243);
nand U95 (N_95,In_389,In_108);
and U96 (N_96,In_292,In_31);
nor U97 (N_97,N_37,In_135);
nor U98 (N_98,In_485,In_496);
or U99 (N_99,In_475,In_308);
or U100 (N_100,In_118,In_467);
nand U101 (N_101,In_474,In_77);
nand U102 (N_102,In_333,N_52);
and U103 (N_103,In_50,N_12);
nor U104 (N_104,In_216,In_488);
nor U105 (N_105,In_434,In_293);
xnor U106 (N_106,N_36,In_56);
nor U107 (N_107,In_345,In_288);
nand U108 (N_108,In_13,In_15);
nand U109 (N_109,In_166,In_359);
nor U110 (N_110,In_417,In_347);
nor U111 (N_111,In_178,In_151);
xnor U112 (N_112,N_23,In_173);
nor U113 (N_113,In_451,In_460);
xor U114 (N_114,N_31,In_22);
and U115 (N_115,In_393,N_42);
or U116 (N_116,In_287,In_277);
or U117 (N_117,In_49,In_428);
xor U118 (N_118,In_42,In_36);
nor U119 (N_119,In_180,In_156);
nor U120 (N_120,In_281,In_343);
nor U121 (N_121,In_289,In_390);
xnor U122 (N_122,N_20,In_268);
nor U123 (N_123,In_41,N_57);
nor U124 (N_124,N_77,In_441);
xor U125 (N_125,In_181,In_379);
and U126 (N_126,In_247,N_14);
or U127 (N_127,In_259,In_495);
or U128 (N_128,In_163,N_11);
nand U129 (N_129,In_230,N_58);
nand U130 (N_130,In_20,In_38);
nand U131 (N_131,In_368,In_152);
nand U132 (N_132,In_271,N_92);
or U133 (N_133,In_182,In_155);
or U134 (N_134,N_82,In_342);
or U135 (N_135,In_350,In_177);
and U136 (N_136,In_272,In_24);
or U137 (N_137,In_215,In_331);
or U138 (N_138,N_116,In_459);
xor U139 (N_139,N_21,In_48);
nor U140 (N_140,In_291,In_99);
and U141 (N_141,In_299,In_329);
or U142 (N_142,N_47,In_211);
nor U143 (N_143,In_388,In_78);
and U144 (N_144,In_242,N_63);
xnor U145 (N_145,In_12,In_471);
xor U146 (N_146,In_104,In_11);
or U147 (N_147,In_314,In_164);
and U148 (N_148,In_456,In_371);
or U149 (N_149,N_85,N_118);
nor U150 (N_150,In_39,In_447);
nand U151 (N_151,In_321,In_112);
or U152 (N_152,In_7,In_197);
and U153 (N_153,N_45,N_93);
xor U154 (N_154,In_410,In_122);
and U155 (N_155,N_43,N_114);
xnor U156 (N_156,N_74,In_65);
xor U157 (N_157,In_191,N_102);
nand U158 (N_158,N_81,In_300);
nand U159 (N_159,N_33,N_72);
xnor U160 (N_160,In_85,In_439);
nor U161 (N_161,In_187,In_51);
nor U162 (N_162,In_399,N_24);
xor U163 (N_163,In_125,In_74);
and U164 (N_164,N_65,In_201);
and U165 (N_165,N_22,N_28);
or U166 (N_166,In_14,In_354);
nor U167 (N_167,In_218,In_105);
nor U168 (N_168,In_26,N_73);
xnor U169 (N_169,In_231,In_338);
and U170 (N_170,N_119,N_111);
nor U171 (N_171,In_142,In_455);
nor U172 (N_172,In_82,In_366);
xnor U173 (N_173,N_75,In_133);
or U174 (N_174,N_35,In_304);
nand U175 (N_175,In_30,In_33);
xor U176 (N_176,In_330,In_328);
nor U177 (N_177,In_206,N_68);
xnor U178 (N_178,N_97,In_437);
and U179 (N_179,In_260,In_165);
nor U180 (N_180,In_95,N_34);
or U181 (N_181,In_336,N_178);
xnor U182 (N_182,In_219,In_339);
nand U183 (N_183,In_498,In_225);
nor U184 (N_184,In_110,N_138);
nand U185 (N_185,In_252,In_6);
and U186 (N_186,N_4,N_25);
xor U187 (N_187,In_463,In_37);
nand U188 (N_188,N_71,In_265);
or U189 (N_189,N_151,In_394);
and U190 (N_190,In_241,In_27);
nand U191 (N_191,N_148,In_311);
xnor U192 (N_192,In_195,In_210);
nor U193 (N_193,In_358,N_165);
or U194 (N_194,N_103,In_316);
or U195 (N_195,N_99,In_169);
nand U196 (N_196,In_200,N_56);
nand U197 (N_197,In_266,In_83);
nor U198 (N_198,In_161,N_113);
or U199 (N_199,In_486,N_130);
nand U200 (N_200,In_94,In_84);
or U201 (N_201,N_123,N_125);
nand U202 (N_202,In_290,N_160);
and U203 (N_203,N_5,In_214);
xnor U204 (N_204,In_238,In_45);
nand U205 (N_205,N_144,In_318);
nand U206 (N_206,In_405,In_25);
and U207 (N_207,N_3,N_46);
or U208 (N_208,N_100,In_262);
or U209 (N_209,In_213,N_149);
xnor U210 (N_210,In_34,In_382);
or U211 (N_211,In_362,N_1);
and U212 (N_212,In_223,In_76);
or U213 (N_213,In_482,N_59);
xnor U214 (N_214,In_147,In_396);
nor U215 (N_215,In_484,In_81);
or U216 (N_216,In_171,In_369);
xor U217 (N_217,In_61,N_115);
nand U218 (N_218,In_400,In_380);
nand U219 (N_219,In_129,In_98);
nor U220 (N_220,In_444,N_61);
nand U221 (N_221,N_139,In_16);
nand U222 (N_222,In_404,In_355);
and U223 (N_223,N_166,N_95);
nand U224 (N_224,N_88,In_115);
and U225 (N_225,N_163,N_129);
nand U226 (N_226,In_232,In_392);
xnor U227 (N_227,In_87,In_148);
or U228 (N_228,In_280,N_13);
or U229 (N_229,N_16,N_169);
and U230 (N_230,In_28,N_156);
xor U231 (N_231,N_137,N_49);
nor U232 (N_232,In_278,N_170);
and U233 (N_233,In_446,N_29);
or U234 (N_234,N_91,N_18);
nand U235 (N_235,In_469,N_19);
nor U236 (N_236,N_155,In_464);
or U237 (N_237,N_50,N_161);
or U238 (N_238,N_69,In_344);
nand U239 (N_239,In_183,N_76);
xnor U240 (N_240,In_274,In_479);
or U241 (N_241,In_21,N_172);
and U242 (N_242,In_162,In_8);
nor U243 (N_243,N_110,N_101);
nor U244 (N_244,N_229,In_120);
and U245 (N_245,In_360,N_146);
or U246 (N_246,N_141,N_159);
xor U247 (N_247,N_233,In_131);
and U248 (N_248,In_378,In_430);
nor U249 (N_249,In_138,N_112);
and U250 (N_250,N_51,In_9);
nor U251 (N_251,N_128,N_217);
xnor U252 (N_252,N_173,N_193);
or U253 (N_253,In_63,In_46);
nand U254 (N_254,In_226,N_30);
and U255 (N_255,In_234,In_150);
xor U256 (N_256,In_212,In_207);
nor U257 (N_257,N_124,N_218);
and U258 (N_258,In_462,N_236);
or U259 (N_259,N_191,N_201);
nand U260 (N_260,N_192,N_222);
or U261 (N_261,In_373,N_184);
and U262 (N_262,N_224,N_108);
and U263 (N_263,In_221,N_239);
nand U264 (N_264,N_10,N_190);
nand U265 (N_265,N_80,N_98);
and U266 (N_266,N_136,N_6);
and U267 (N_267,N_117,N_231);
nand U268 (N_268,In_435,N_223);
nand U269 (N_269,N_135,N_86);
and U270 (N_270,N_232,N_41);
nand U271 (N_271,In_466,N_79);
nand U272 (N_272,In_407,In_72);
or U273 (N_273,In_383,N_145);
or U274 (N_274,In_477,N_168);
and U275 (N_275,In_296,N_187);
nor U276 (N_276,In_401,In_205);
nor U277 (N_277,N_126,In_493);
xnor U278 (N_278,N_228,N_132);
and U279 (N_279,In_452,N_96);
nand U280 (N_280,In_60,In_153);
or U281 (N_281,N_26,N_104);
nor U282 (N_282,N_39,In_334);
and U283 (N_283,In_408,In_158);
nand U284 (N_284,In_62,N_109);
nor U285 (N_285,In_270,N_158);
xor U286 (N_286,In_494,In_285);
and U287 (N_287,N_121,N_188);
nand U288 (N_288,N_62,In_421);
nand U289 (N_289,N_230,N_122);
nand U290 (N_290,N_70,In_2);
nand U291 (N_291,N_176,N_162);
and U292 (N_292,In_137,N_66);
xor U293 (N_293,In_208,N_106);
or U294 (N_294,N_189,N_212);
or U295 (N_295,N_198,In_250);
nor U296 (N_296,N_181,In_276);
and U297 (N_297,In_433,In_315);
and U298 (N_298,N_48,In_23);
and U299 (N_299,N_142,N_226);
and U300 (N_300,N_246,N_55);
nor U301 (N_301,N_143,N_237);
xnor U302 (N_302,In_168,In_375);
and U303 (N_303,In_127,N_200);
or U304 (N_304,In_431,N_195);
nor U305 (N_305,N_133,In_235);
nor U306 (N_306,In_445,N_153);
xor U307 (N_307,N_183,In_402);
nor U308 (N_308,N_157,In_204);
nor U309 (N_309,N_258,In_351);
or U310 (N_310,N_298,N_127);
nand U311 (N_311,N_154,N_207);
nor U312 (N_312,N_78,N_260);
and U313 (N_313,N_261,N_175);
nand U314 (N_314,N_250,N_244);
nand U315 (N_315,In_263,N_214);
or U316 (N_316,In_425,In_257);
or U317 (N_317,In_303,In_361);
nand U318 (N_318,N_167,N_281);
or U319 (N_319,In_92,N_251);
nand U320 (N_320,N_257,In_227);
nor U321 (N_321,In_124,In_139);
or U322 (N_322,In_113,In_406);
nor U323 (N_323,N_248,N_253);
and U324 (N_324,In_251,N_271);
or U325 (N_325,N_262,N_289);
and U326 (N_326,N_60,N_2);
xnor U327 (N_327,In_448,N_284);
nand U328 (N_328,N_270,In_297);
and U329 (N_329,N_209,N_265);
or U330 (N_330,In_3,N_287);
or U331 (N_331,N_89,N_147);
nor U332 (N_332,N_254,N_131);
and U333 (N_333,In_267,In_196);
xnor U334 (N_334,N_105,In_255);
and U335 (N_335,N_216,In_199);
xor U336 (N_336,N_243,In_228);
nand U337 (N_337,In_188,N_295);
and U338 (N_338,N_264,N_290);
and U339 (N_339,In_175,N_185);
and U340 (N_340,N_291,N_220);
nand U341 (N_341,N_225,N_275);
or U342 (N_342,In_79,N_150);
nand U343 (N_343,N_182,N_87);
and U344 (N_344,N_179,N_276);
and U345 (N_345,N_277,N_293);
xnor U346 (N_346,In_442,N_296);
or U347 (N_347,In_119,N_134);
nand U348 (N_348,In_335,In_220);
xnor U349 (N_349,N_202,In_186);
and U350 (N_350,In_103,N_273);
nor U351 (N_351,In_465,N_206);
or U352 (N_352,N_180,N_279);
nor U353 (N_353,N_186,N_215);
or U354 (N_354,N_249,N_285);
xor U355 (N_355,N_247,N_238);
or U356 (N_356,N_252,N_84);
nand U357 (N_357,In_454,N_242);
nand U358 (N_358,In_193,In_492);
nor U359 (N_359,N_196,N_299);
and U360 (N_360,N_67,N_268);
or U361 (N_361,N_338,In_202);
and U362 (N_362,N_342,N_314);
xor U363 (N_363,N_340,N_319);
xor U364 (N_364,N_211,N_213);
xnor U365 (N_365,In_317,N_323);
nand U366 (N_366,N_234,N_140);
xnor U367 (N_367,N_269,N_345);
nor U368 (N_368,N_318,N_341);
xor U369 (N_369,N_107,N_307);
or U370 (N_370,N_309,In_121);
and U371 (N_371,In_222,N_219);
xnor U372 (N_372,In_349,N_351);
xor U373 (N_373,N_272,N_292);
or U374 (N_374,N_359,N_0);
nor U375 (N_375,N_320,N_325);
xor U376 (N_376,N_245,N_171);
or U377 (N_377,N_316,N_280);
and U378 (N_378,N_241,N_294);
nand U379 (N_379,In_470,N_355);
or U380 (N_380,N_331,N_339);
nor U381 (N_381,In_89,In_209);
nor U382 (N_382,N_199,N_348);
or U383 (N_383,In_302,N_308);
or U384 (N_384,N_210,N_297);
nor U385 (N_385,N_357,N_263);
or U386 (N_386,N_327,N_90);
and U387 (N_387,N_27,N_358);
nand U388 (N_388,N_266,In_341);
nand U389 (N_389,N_310,In_420);
and U390 (N_390,In_313,N_259);
and U391 (N_391,N_177,N_83);
or U392 (N_392,N_335,N_356);
and U393 (N_393,In_398,N_311);
and U394 (N_394,In_305,N_152);
xor U395 (N_395,N_255,In_136);
and U396 (N_396,In_224,N_344);
xnor U397 (N_397,In_154,N_64);
xnor U398 (N_398,N_350,N_286);
xor U399 (N_399,N_347,N_203);
and U400 (N_400,N_204,N_256);
nor U401 (N_401,N_282,N_120);
or U402 (N_402,N_235,N_32);
or U403 (N_403,N_283,N_334);
xnor U404 (N_404,N_44,N_315);
or U405 (N_405,N_205,N_53);
or U406 (N_406,N_321,N_337);
nor U407 (N_407,N_343,N_300);
and U408 (N_408,N_312,N_302);
or U409 (N_409,N_332,N_324);
or U410 (N_410,N_94,N_330);
nor U411 (N_411,In_429,N_301);
xnor U412 (N_412,N_329,N_326);
xnor U413 (N_413,N_208,N_227);
or U414 (N_414,In_363,N_240);
nand U415 (N_415,N_304,N_303);
nor U416 (N_416,N_333,N_174);
xnor U417 (N_417,N_267,N_274);
nor U418 (N_418,N_322,In_377);
nand U419 (N_419,N_278,N_164);
nor U420 (N_420,N_409,N_403);
or U421 (N_421,N_395,N_360);
xnor U422 (N_422,N_407,N_418);
nor U423 (N_423,N_390,N_373);
xnor U424 (N_424,N_387,N_346);
xnor U425 (N_425,N_393,N_349);
and U426 (N_426,N_366,N_353);
nand U427 (N_427,N_365,N_377);
nand U428 (N_428,N_381,N_383);
nor U429 (N_429,N_404,N_392);
or U430 (N_430,N_369,N_382);
or U431 (N_431,N_397,N_415);
and U432 (N_432,N_197,N_394);
and U433 (N_433,N_405,N_379);
and U434 (N_434,N_419,In_132);
and U435 (N_435,N_354,In_73);
nand U436 (N_436,N_367,N_414);
nand U437 (N_437,N_194,N_386);
nand U438 (N_438,N_388,N_378);
nand U439 (N_439,N_402,N_389);
nor U440 (N_440,N_368,N_413);
nand U441 (N_441,In_312,N_396);
nand U442 (N_442,N_305,N_370);
or U443 (N_443,N_391,N_221);
nor U444 (N_444,N_317,N_364);
or U445 (N_445,N_416,N_336);
and U446 (N_446,N_406,N_412);
nor U447 (N_447,In_491,N_313);
nor U448 (N_448,N_288,N_380);
or U449 (N_449,N_352,N_385);
xor U450 (N_450,N_328,N_410);
nor U451 (N_451,N_375,N_411);
nand U452 (N_452,N_417,N_372);
and U453 (N_453,N_371,N_374);
nor U454 (N_454,In_275,N_363);
xor U455 (N_455,N_400,N_398);
xor U456 (N_456,N_361,N_384);
or U457 (N_457,N_408,N_362);
or U458 (N_458,N_306,N_376);
nand U459 (N_459,N_399,N_401);
nand U460 (N_460,N_364,N_363);
or U461 (N_461,N_402,N_367);
nor U462 (N_462,N_393,N_376);
nor U463 (N_463,N_362,N_336);
nand U464 (N_464,N_390,N_364);
or U465 (N_465,N_409,N_410);
nor U466 (N_466,N_375,N_396);
and U467 (N_467,N_378,In_73);
xnor U468 (N_468,N_385,N_401);
nor U469 (N_469,N_391,N_349);
or U470 (N_470,N_328,N_367);
xnor U471 (N_471,N_394,N_366);
xnor U472 (N_472,N_394,N_372);
nand U473 (N_473,N_405,N_382);
xor U474 (N_474,N_349,N_328);
nand U475 (N_475,N_361,N_395);
nor U476 (N_476,N_313,N_397);
nor U477 (N_477,N_197,N_375);
or U478 (N_478,N_411,N_317);
xor U479 (N_479,N_362,N_418);
nand U480 (N_480,N_458,N_425);
or U481 (N_481,N_466,N_424);
nor U482 (N_482,N_477,N_446);
xor U483 (N_483,N_448,N_433);
nand U484 (N_484,N_431,N_462);
nor U485 (N_485,N_423,N_451);
and U486 (N_486,N_421,N_464);
and U487 (N_487,N_465,N_430);
nor U488 (N_488,N_468,N_445);
xor U489 (N_489,N_471,N_453);
and U490 (N_490,N_478,N_460);
xor U491 (N_491,N_447,N_475);
xor U492 (N_492,N_436,N_476);
and U493 (N_493,N_434,N_428);
nor U494 (N_494,N_459,N_473);
xnor U495 (N_495,N_449,N_463);
and U496 (N_496,N_432,N_455);
xor U497 (N_497,N_450,N_422);
nor U498 (N_498,N_444,N_469);
or U499 (N_499,N_443,N_470);
xnor U500 (N_500,N_441,N_474);
nor U501 (N_501,N_472,N_442);
nor U502 (N_502,N_479,N_439);
nand U503 (N_503,N_435,N_429);
nor U504 (N_504,N_461,N_438);
nand U505 (N_505,N_457,N_420);
or U506 (N_506,N_427,N_437);
xor U507 (N_507,N_426,N_440);
nand U508 (N_508,N_467,N_454);
and U509 (N_509,N_452,N_456);
nand U510 (N_510,N_473,N_467);
nor U511 (N_511,N_437,N_421);
xnor U512 (N_512,N_432,N_426);
or U513 (N_513,N_458,N_439);
and U514 (N_514,N_457,N_469);
or U515 (N_515,N_451,N_455);
nand U516 (N_516,N_442,N_475);
nor U517 (N_517,N_449,N_441);
nand U518 (N_518,N_467,N_453);
or U519 (N_519,N_451,N_433);
nand U520 (N_520,N_459,N_453);
nand U521 (N_521,N_426,N_456);
nor U522 (N_522,N_445,N_471);
nor U523 (N_523,N_454,N_461);
nand U524 (N_524,N_422,N_456);
xor U525 (N_525,N_471,N_470);
nand U526 (N_526,N_435,N_427);
nand U527 (N_527,N_428,N_443);
and U528 (N_528,N_447,N_422);
nor U529 (N_529,N_431,N_452);
nor U530 (N_530,N_479,N_469);
nor U531 (N_531,N_432,N_430);
nand U532 (N_532,N_438,N_472);
and U533 (N_533,N_424,N_464);
or U534 (N_534,N_443,N_451);
or U535 (N_535,N_422,N_466);
xnor U536 (N_536,N_475,N_466);
and U537 (N_537,N_436,N_421);
or U538 (N_538,N_468,N_477);
and U539 (N_539,N_477,N_475);
or U540 (N_540,N_483,N_505);
nor U541 (N_541,N_520,N_510);
xor U542 (N_542,N_490,N_516);
nand U543 (N_543,N_498,N_504);
nand U544 (N_544,N_493,N_482);
nand U545 (N_545,N_508,N_537);
nand U546 (N_546,N_536,N_529);
nor U547 (N_547,N_488,N_486);
or U548 (N_548,N_538,N_533);
nor U549 (N_549,N_514,N_524);
or U550 (N_550,N_535,N_500);
or U551 (N_551,N_526,N_484);
or U552 (N_552,N_502,N_480);
or U553 (N_553,N_492,N_511);
or U554 (N_554,N_501,N_517);
and U555 (N_555,N_531,N_489);
and U556 (N_556,N_539,N_525);
or U557 (N_557,N_523,N_532);
and U558 (N_558,N_491,N_487);
nand U559 (N_559,N_522,N_499);
nor U560 (N_560,N_519,N_513);
nand U561 (N_561,N_527,N_512);
or U562 (N_562,N_518,N_534);
nand U563 (N_563,N_521,N_496);
and U564 (N_564,N_485,N_509);
nor U565 (N_565,N_528,N_530);
and U566 (N_566,N_494,N_495);
and U567 (N_567,N_481,N_503);
xnor U568 (N_568,N_515,N_507);
and U569 (N_569,N_506,N_497);
and U570 (N_570,N_510,N_506);
or U571 (N_571,N_485,N_517);
nor U572 (N_572,N_527,N_497);
and U573 (N_573,N_512,N_501);
and U574 (N_574,N_504,N_495);
nand U575 (N_575,N_528,N_518);
or U576 (N_576,N_489,N_480);
xnor U577 (N_577,N_510,N_508);
xnor U578 (N_578,N_504,N_483);
xor U579 (N_579,N_527,N_514);
nand U580 (N_580,N_492,N_508);
nor U581 (N_581,N_485,N_527);
or U582 (N_582,N_534,N_489);
and U583 (N_583,N_536,N_490);
nor U584 (N_584,N_521,N_501);
xnor U585 (N_585,N_516,N_525);
and U586 (N_586,N_506,N_499);
and U587 (N_587,N_493,N_511);
and U588 (N_588,N_525,N_496);
nand U589 (N_589,N_522,N_510);
and U590 (N_590,N_535,N_487);
and U591 (N_591,N_490,N_538);
or U592 (N_592,N_491,N_481);
nand U593 (N_593,N_485,N_504);
xnor U594 (N_594,N_517,N_506);
xnor U595 (N_595,N_518,N_482);
and U596 (N_596,N_515,N_531);
nand U597 (N_597,N_510,N_513);
nand U598 (N_598,N_482,N_531);
and U599 (N_599,N_505,N_499);
and U600 (N_600,N_574,N_580);
or U601 (N_601,N_563,N_586);
xnor U602 (N_602,N_579,N_540);
xor U603 (N_603,N_558,N_561);
nor U604 (N_604,N_587,N_544);
nor U605 (N_605,N_584,N_598);
xor U606 (N_606,N_557,N_552);
and U607 (N_607,N_549,N_590);
xnor U608 (N_608,N_577,N_589);
and U609 (N_609,N_548,N_553);
xor U610 (N_610,N_592,N_560);
nor U611 (N_611,N_576,N_596);
and U612 (N_612,N_581,N_543);
nand U613 (N_613,N_568,N_541);
and U614 (N_614,N_591,N_550);
or U615 (N_615,N_585,N_567);
xnor U616 (N_616,N_572,N_545);
and U617 (N_617,N_597,N_555);
nand U618 (N_618,N_547,N_565);
xor U619 (N_619,N_546,N_556);
nor U620 (N_620,N_588,N_599);
xor U621 (N_621,N_582,N_559);
or U622 (N_622,N_554,N_569);
nand U623 (N_623,N_570,N_594);
nor U624 (N_624,N_593,N_573);
xnor U625 (N_625,N_575,N_578);
nor U626 (N_626,N_542,N_562);
xor U627 (N_627,N_571,N_583);
xor U628 (N_628,N_595,N_564);
and U629 (N_629,N_551,N_566);
xor U630 (N_630,N_588,N_569);
or U631 (N_631,N_575,N_597);
xnor U632 (N_632,N_564,N_563);
xor U633 (N_633,N_570,N_552);
or U634 (N_634,N_558,N_547);
or U635 (N_635,N_599,N_597);
and U636 (N_636,N_590,N_572);
nand U637 (N_637,N_586,N_576);
xor U638 (N_638,N_576,N_591);
nor U639 (N_639,N_569,N_552);
nand U640 (N_640,N_548,N_543);
and U641 (N_641,N_561,N_573);
nor U642 (N_642,N_550,N_584);
nor U643 (N_643,N_597,N_562);
and U644 (N_644,N_559,N_586);
nand U645 (N_645,N_551,N_547);
or U646 (N_646,N_547,N_582);
and U647 (N_647,N_596,N_572);
and U648 (N_648,N_552,N_574);
and U649 (N_649,N_597,N_596);
nor U650 (N_650,N_565,N_554);
or U651 (N_651,N_541,N_592);
nand U652 (N_652,N_542,N_540);
or U653 (N_653,N_592,N_582);
nor U654 (N_654,N_590,N_562);
or U655 (N_655,N_566,N_596);
or U656 (N_656,N_568,N_578);
or U657 (N_657,N_577,N_584);
nor U658 (N_658,N_593,N_579);
and U659 (N_659,N_543,N_594);
xnor U660 (N_660,N_632,N_605);
and U661 (N_661,N_619,N_636);
nand U662 (N_662,N_655,N_626);
nand U663 (N_663,N_640,N_650);
and U664 (N_664,N_609,N_628);
or U665 (N_665,N_615,N_630);
xnor U666 (N_666,N_651,N_631);
and U667 (N_667,N_603,N_618);
nor U668 (N_668,N_638,N_656);
nand U669 (N_669,N_622,N_606);
and U670 (N_670,N_652,N_635);
xnor U671 (N_671,N_627,N_653);
and U672 (N_672,N_624,N_600);
xor U673 (N_673,N_602,N_647);
xnor U674 (N_674,N_648,N_629);
and U675 (N_675,N_659,N_633);
xor U676 (N_676,N_614,N_613);
and U677 (N_677,N_641,N_644);
or U678 (N_678,N_611,N_645);
xor U679 (N_679,N_646,N_616);
and U680 (N_680,N_654,N_639);
or U681 (N_681,N_607,N_623);
and U682 (N_682,N_601,N_658);
nand U683 (N_683,N_610,N_634);
and U684 (N_684,N_637,N_649);
nor U685 (N_685,N_620,N_625);
or U686 (N_686,N_617,N_643);
nor U687 (N_687,N_657,N_621);
or U688 (N_688,N_612,N_608);
xnor U689 (N_689,N_642,N_604);
nand U690 (N_690,N_643,N_629);
xor U691 (N_691,N_604,N_620);
or U692 (N_692,N_601,N_636);
nor U693 (N_693,N_652,N_637);
xnor U694 (N_694,N_648,N_626);
or U695 (N_695,N_632,N_638);
and U696 (N_696,N_641,N_627);
nand U697 (N_697,N_626,N_651);
or U698 (N_698,N_610,N_633);
nand U699 (N_699,N_611,N_630);
nor U700 (N_700,N_624,N_637);
or U701 (N_701,N_608,N_643);
or U702 (N_702,N_658,N_644);
and U703 (N_703,N_659,N_647);
nor U704 (N_704,N_614,N_627);
xor U705 (N_705,N_640,N_627);
or U706 (N_706,N_656,N_644);
xor U707 (N_707,N_635,N_641);
and U708 (N_708,N_653,N_658);
nor U709 (N_709,N_656,N_602);
or U710 (N_710,N_627,N_618);
and U711 (N_711,N_652,N_627);
and U712 (N_712,N_648,N_618);
nand U713 (N_713,N_635,N_631);
and U714 (N_714,N_618,N_638);
xor U715 (N_715,N_659,N_642);
and U716 (N_716,N_640,N_607);
or U717 (N_717,N_604,N_603);
xor U718 (N_718,N_609,N_616);
nand U719 (N_719,N_629,N_605);
and U720 (N_720,N_706,N_677);
or U721 (N_721,N_699,N_681);
and U722 (N_722,N_661,N_688);
nor U723 (N_723,N_695,N_703);
xor U724 (N_724,N_672,N_684);
nor U725 (N_725,N_712,N_664);
and U726 (N_726,N_718,N_680);
xor U727 (N_727,N_669,N_711);
or U728 (N_728,N_704,N_679);
or U729 (N_729,N_668,N_689);
xnor U730 (N_730,N_690,N_675);
xor U731 (N_731,N_665,N_696);
nand U732 (N_732,N_694,N_691);
nor U733 (N_733,N_663,N_698);
nand U734 (N_734,N_713,N_697);
xor U735 (N_735,N_671,N_674);
and U736 (N_736,N_715,N_673);
xor U737 (N_737,N_719,N_714);
and U738 (N_738,N_683,N_676);
and U739 (N_739,N_682,N_700);
nand U740 (N_740,N_702,N_670);
and U741 (N_741,N_667,N_708);
or U742 (N_742,N_660,N_705);
nor U743 (N_743,N_687,N_685);
or U744 (N_744,N_701,N_693);
nor U745 (N_745,N_717,N_678);
nand U746 (N_746,N_710,N_709);
or U747 (N_747,N_707,N_686);
xnor U748 (N_748,N_662,N_716);
and U749 (N_749,N_666,N_692);
xor U750 (N_750,N_690,N_660);
nor U751 (N_751,N_689,N_686);
nand U752 (N_752,N_663,N_690);
or U753 (N_753,N_694,N_703);
and U754 (N_754,N_718,N_686);
xor U755 (N_755,N_703,N_669);
nand U756 (N_756,N_675,N_672);
or U757 (N_757,N_661,N_685);
nor U758 (N_758,N_667,N_670);
nand U759 (N_759,N_682,N_684);
and U760 (N_760,N_709,N_668);
xnor U761 (N_761,N_683,N_709);
and U762 (N_762,N_662,N_669);
and U763 (N_763,N_714,N_717);
or U764 (N_764,N_669,N_709);
nand U765 (N_765,N_714,N_693);
or U766 (N_766,N_689,N_688);
or U767 (N_767,N_681,N_710);
nand U768 (N_768,N_696,N_666);
or U769 (N_769,N_693,N_676);
xnor U770 (N_770,N_667,N_682);
and U771 (N_771,N_680,N_715);
xor U772 (N_772,N_691,N_684);
or U773 (N_773,N_697,N_669);
nor U774 (N_774,N_698,N_677);
and U775 (N_775,N_698,N_678);
nand U776 (N_776,N_703,N_676);
nor U777 (N_777,N_704,N_703);
or U778 (N_778,N_660,N_685);
and U779 (N_779,N_670,N_669);
nor U780 (N_780,N_763,N_733);
and U781 (N_781,N_768,N_731);
or U782 (N_782,N_726,N_746);
and U783 (N_783,N_752,N_744);
xor U784 (N_784,N_740,N_749);
xnor U785 (N_785,N_779,N_754);
nor U786 (N_786,N_753,N_720);
and U787 (N_787,N_771,N_747);
nor U788 (N_788,N_769,N_727);
xor U789 (N_789,N_761,N_766);
or U790 (N_790,N_732,N_739);
xor U791 (N_791,N_728,N_765);
and U792 (N_792,N_721,N_722);
nor U793 (N_793,N_730,N_778);
nand U794 (N_794,N_774,N_729);
or U795 (N_795,N_757,N_742);
nand U796 (N_796,N_737,N_735);
xor U797 (N_797,N_762,N_748);
and U798 (N_798,N_751,N_741);
and U799 (N_799,N_777,N_755);
and U800 (N_800,N_745,N_738);
nor U801 (N_801,N_770,N_734);
nor U802 (N_802,N_723,N_760);
nor U803 (N_803,N_736,N_759);
nand U804 (N_804,N_750,N_772);
and U805 (N_805,N_758,N_764);
xor U806 (N_806,N_756,N_725);
and U807 (N_807,N_767,N_773);
or U808 (N_808,N_775,N_743);
or U809 (N_809,N_776,N_724);
nor U810 (N_810,N_744,N_735);
and U811 (N_811,N_772,N_729);
and U812 (N_812,N_767,N_750);
or U813 (N_813,N_779,N_730);
nor U814 (N_814,N_749,N_750);
nand U815 (N_815,N_774,N_771);
xnor U816 (N_816,N_742,N_747);
or U817 (N_817,N_777,N_724);
xor U818 (N_818,N_777,N_764);
and U819 (N_819,N_737,N_771);
and U820 (N_820,N_732,N_735);
or U821 (N_821,N_727,N_756);
xor U822 (N_822,N_735,N_741);
nand U823 (N_823,N_771,N_750);
nand U824 (N_824,N_752,N_758);
or U825 (N_825,N_748,N_767);
nand U826 (N_826,N_772,N_767);
xnor U827 (N_827,N_738,N_758);
and U828 (N_828,N_755,N_754);
xor U829 (N_829,N_759,N_722);
or U830 (N_830,N_747,N_725);
nand U831 (N_831,N_777,N_734);
nor U832 (N_832,N_747,N_770);
nand U833 (N_833,N_778,N_761);
nor U834 (N_834,N_757,N_723);
and U835 (N_835,N_772,N_773);
nand U836 (N_836,N_752,N_771);
and U837 (N_837,N_750,N_759);
and U838 (N_838,N_766,N_768);
and U839 (N_839,N_730,N_758);
xor U840 (N_840,N_803,N_825);
nand U841 (N_841,N_836,N_826);
xnor U842 (N_842,N_786,N_805);
and U843 (N_843,N_820,N_785);
and U844 (N_844,N_821,N_819);
or U845 (N_845,N_822,N_817);
and U846 (N_846,N_839,N_797);
nand U847 (N_847,N_827,N_832);
xor U848 (N_848,N_837,N_795);
nor U849 (N_849,N_815,N_824);
and U850 (N_850,N_781,N_816);
and U851 (N_851,N_799,N_809);
nand U852 (N_852,N_788,N_814);
and U853 (N_853,N_835,N_838);
xor U854 (N_854,N_806,N_828);
and U855 (N_855,N_801,N_780);
xnor U856 (N_856,N_782,N_796);
nand U857 (N_857,N_810,N_798);
nand U858 (N_858,N_792,N_789);
xor U859 (N_859,N_812,N_823);
nor U860 (N_860,N_831,N_834);
nor U861 (N_861,N_818,N_833);
and U862 (N_862,N_790,N_784);
nand U863 (N_863,N_787,N_802);
or U864 (N_864,N_808,N_830);
or U865 (N_865,N_800,N_794);
nand U866 (N_866,N_804,N_829);
or U867 (N_867,N_793,N_813);
and U868 (N_868,N_783,N_811);
and U869 (N_869,N_807,N_791);
or U870 (N_870,N_799,N_837);
and U871 (N_871,N_783,N_793);
nor U872 (N_872,N_825,N_813);
nand U873 (N_873,N_796,N_791);
nor U874 (N_874,N_816,N_817);
and U875 (N_875,N_780,N_799);
nand U876 (N_876,N_832,N_783);
xor U877 (N_877,N_798,N_838);
nand U878 (N_878,N_811,N_838);
nand U879 (N_879,N_805,N_796);
and U880 (N_880,N_832,N_786);
or U881 (N_881,N_797,N_818);
nor U882 (N_882,N_796,N_820);
nor U883 (N_883,N_820,N_824);
or U884 (N_884,N_793,N_830);
nand U885 (N_885,N_827,N_788);
and U886 (N_886,N_806,N_802);
xnor U887 (N_887,N_818,N_809);
or U888 (N_888,N_811,N_801);
xnor U889 (N_889,N_820,N_809);
nor U890 (N_890,N_789,N_798);
or U891 (N_891,N_837,N_794);
xnor U892 (N_892,N_836,N_825);
nor U893 (N_893,N_820,N_795);
and U894 (N_894,N_797,N_786);
nor U895 (N_895,N_815,N_823);
nand U896 (N_896,N_795,N_794);
xnor U897 (N_897,N_832,N_831);
nand U898 (N_898,N_782,N_830);
or U899 (N_899,N_836,N_828);
or U900 (N_900,N_881,N_878);
nor U901 (N_901,N_841,N_870);
nor U902 (N_902,N_890,N_854);
or U903 (N_903,N_883,N_855);
or U904 (N_904,N_869,N_895);
nand U905 (N_905,N_893,N_849);
xor U906 (N_906,N_867,N_894);
nor U907 (N_907,N_860,N_866);
nor U908 (N_908,N_880,N_885);
xnor U909 (N_909,N_899,N_858);
and U910 (N_910,N_877,N_852);
xor U911 (N_911,N_874,N_850);
or U912 (N_912,N_896,N_882);
and U913 (N_913,N_856,N_861);
or U914 (N_914,N_862,N_851);
or U915 (N_915,N_891,N_842);
xor U916 (N_916,N_884,N_892);
nand U917 (N_917,N_865,N_889);
and U918 (N_918,N_875,N_873);
or U919 (N_919,N_876,N_848);
and U920 (N_920,N_898,N_853);
or U921 (N_921,N_845,N_887);
nand U922 (N_922,N_846,N_859);
nor U923 (N_923,N_844,N_872);
nand U924 (N_924,N_840,N_864);
and U925 (N_925,N_863,N_871);
xnor U926 (N_926,N_879,N_857);
or U927 (N_927,N_897,N_888);
nor U928 (N_928,N_886,N_847);
and U929 (N_929,N_843,N_868);
nor U930 (N_930,N_899,N_875);
xnor U931 (N_931,N_872,N_851);
nand U932 (N_932,N_884,N_893);
nand U933 (N_933,N_862,N_893);
nor U934 (N_934,N_882,N_856);
nand U935 (N_935,N_873,N_842);
xnor U936 (N_936,N_857,N_851);
or U937 (N_937,N_850,N_842);
nand U938 (N_938,N_874,N_897);
and U939 (N_939,N_867,N_881);
and U940 (N_940,N_899,N_844);
or U941 (N_941,N_892,N_855);
xnor U942 (N_942,N_895,N_899);
nand U943 (N_943,N_899,N_866);
nor U944 (N_944,N_898,N_867);
xor U945 (N_945,N_841,N_862);
nand U946 (N_946,N_845,N_868);
nor U947 (N_947,N_892,N_850);
nor U948 (N_948,N_866,N_873);
xnor U949 (N_949,N_862,N_868);
xnor U950 (N_950,N_858,N_854);
and U951 (N_951,N_889,N_846);
and U952 (N_952,N_842,N_896);
xor U953 (N_953,N_847,N_896);
xor U954 (N_954,N_898,N_845);
nor U955 (N_955,N_861,N_896);
nor U956 (N_956,N_884,N_890);
or U957 (N_957,N_864,N_883);
xnor U958 (N_958,N_896,N_853);
and U959 (N_959,N_841,N_840);
and U960 (N_960,N_944,N_912);
nand U961 (N_961,N_920,N_947);
nor U962 (N_962,N_907,N_911);
or U963 (N_963,N_948,N_945);
and U964 (N_964,N_932,N_942);
and U965 (N_965,N_923,N_949);
nand U966 (N_966,N_951,N_917);
and U967 (N_967,N_904,N_933);
xnor U968 (N_968,N_936,N_924);
or U969 (N_969,N_938,N_902);
and U970 (N_970,N_929,N_910);
nor U971 (N_971,N_928,N_931);
or U972 (N_972,N_952,N_939);
and U973 (N_973,N_941,N_921);
nand U974 (N_974,N_903,N_913);
and U975 (N_975,N_909,N_927);
nor U976 (N_976,N_956,N_926);
and U977 (N_977,N_916,N_919);
nand U978 (N_978,N_958,N_901);
xnor U979 (N_979,N_950,N_957);
xnor U980 (N_980,N_937,N_915);
and U981 (N_981,N_934,N_908);
and U982 (N_982,N_959,N_930);
or U983 (N_983,N_905,N_922);
xor U984 (N_984,N_935,N_953);
or U985 (N_985,N_918,N_955);
xnor U986 (N_986,N_943,N_946);
xor U987 (N_987,N_900,N_940);
xnor U988 (N_988,N_954,N_925);
or U989 (N_989,N_914,N_906);
nand U990 (N_990,N_904,N_925);
or U991 (N_991,N_902,N_907);
nand U992 (N_992,N_936,N_902);
xor U993 (N_993,N_917,N_947);
or U994 (N_994,N_932,N_907);
and U995 (N_995,N_929,N_941);
or U996 (N_996,N_918,N_944);
nand U997 (N_997,N_901,N_947);
nand U998 (N_998,N_903,N_916);
and U999 (N_999,N_954,N_947);
nand U1000 (N_1000,N_911,N_919);
nor U1001 (N_1001,N_915,N_909);
nor U1002 (N_1002,N_919,N_921);
xnor U1003 (N_1003,N_955,N_920);
nor U1004 (N_1004,N_937,N_946);
xnor U1005 (N_1005,N_947,N_949);
or U1006 (N_1006,N_927,N_940);
nor U1007 (N_1007,N_903,N_910);
nand U1008 (N_1008,N_932,N_952);
or U1009 (N_1009,N_938,N_905);
xor U1010 (N_1010,N_946,N_957);
and U1011 (N_1011,N_933,N_928);
or U1012 (N_1012,N_917,N_914);
or U1013 (N_1013,N_944,N_954);
or U1014 (N_1014,N_919,N_940);
nor U1015 (N_1015,N_918,N_928);
or U1016 (N_1016,N_927,N_955);
nand U1017 (N_1017,N_955,N_901);
and U1018 (N_1018,N_944,N_916);
nand U1019 (N_1019,N_921,N_940);
or U1020 (N_1020,N_980,N_1007);
xnor U1021 (N_1021,N_977,N_975);
and U1022 (N_1022,N_1015,N_967);
nand U1023 (N_1023,N_1012,N_1011);
and U1024 (N_1024,N_1000,N_1010);
or U1025 (N_1025,N_1004,N_983);
nor U1026 (N_1026,N_1017,N_1013);
or U1027 (N_1027,N_963,N_976);
or U1028 (N_1028,N_970,N_972);
or U1029 (N_1029,N_996,N_987);
nand U1030 (N_1030,N_1005,N_999);
and U1031 (N_1031,N_968,N_960);
nor U1032 (N_1032,N_1008,N_962);
and U1033 (N_1033,N_973,N_988);
and U1034 (N_1034,N_1009,N_1001);
nand U1035 (N_1035,N_997,N_979);
xnor U1036 (N_1036,N_990,N_989);
nor U1037 (N_1037,N_1014,N_1018);
nor U1038 (N_1038,N_1019,N_994);
and U1039 (N_1039,N_971,N_985);
or U1040 (N_1040,N_995,N_961);
and U1041 (N_1041,N_978,N_1016);
and U1042 (N_1042,N_982,N_965);
or U1043 (N_1043,N_966,N_992);
nor U1044 (N_1044,N_984,N_1003);
or U1045 (N_1045,N_991,N_1002);
nor U1046 (N_1046,N_986,N_964);
nor U1047 (N_1047,N_1006,N_969);
and U1048 (N_1048,N_998,N_993);
nand U1049 (N_1049,N_981,N_974);
nor U1050 (N_1050,N_985,N_966);
or U1051 (N_1051,N_1009,N_965);
nand U1052 (N_1052,N_1016,N_983);
nor U1053 (N_1053,N_1009,N_994);
nand U1054 (N_1054,N_993,N_1001);
nor U1055 (N_1055,N_1019,N_1000);
or U1056 (N_1056,N_988,N_982);
xor U1057 (N_1057,N_988,N_966);
xor U1058 (N_1058,N_982,N_996);
nand U1059 (N_1059,N_997,N_1008);
nor U1060 (N_1060,N_985,N_1002);
nor U1061 (N_1061,N_963,N_982);
nor U1062 (N_1062,N_973,N_962);
nand U1063 (N_1063,N_964,N_1009);
xor U1064 (N_1064,N_975,N_1011);
xor U1065 (N_1065,N_982,N_995);
or U1066 (N_1066,N_976,N_987);
or U1067 (N_1067,N_998,N_1015);
or U1068 (N_1068,N_973,N_991);
xnor U1069 (N_1069,N_993,N_974);
and U1070 (N_1070,N_960,N_974);
nor U1071 (N_1071,N_966,N_1008);
xnor U1072 (N_1072,N_992,N_995);
and U1073 (N_1073,N_967,N_979);
nor U1074 (N_1074,N_995,N_1002);
nor U1075 (N_1075,N_995,N_1015);
nand U1076 (N_1076,N_971,N_994);
or U1077 (N_1077,N_961,N_988);
nor U1078 (N_1078,N_973,N_990);
or U1079 (N_1079,N_987,N_1011);
nand U1080 (N_1080,N_1056,N_1067);
nor U1081 (N_1081,N_1065,N_1041);
xnor U1082 (N_1082,N_1060,N_1029);
nor U1083 (N_1083,N_1059,N_1020);
nor U1084 (N_1084,N_1068,N_1055);
nand U1085 (N_1085,N_1043,N_1039);
or U1086 (N_1086,N_1047,N_1053);
nor U1087 (N_1087,N_1036,N_1042);
xnor U1088 (N_1088,N_1038,N_1069);
nor U1089 (N_1089,N_1050,N_1037);
or U1090 (N_1090,N_1048,N_1044);
and U1091 (N_1091,N_1070,N_1028);
nand U1092 (N_1092,N_1025,N_1063);
or U1093 (N_1093,N_1064,N_1058);
nand U1094 (N_1094,N_1021,N_1062);
nand U1095 (N_1095,N_1045,N_1040);
and U1096 (N_1096,N_1074,N_1054);
and U1097 (N_1097,N_1066,N_1073);
and U1098 (N_1098,N_1061,N_1023);
or U1099 (N_1099,N_1079,N_1052);
nand U1100 (N_1100,N_1051,N_1075);
or U1101 (N_1101,N_1030,N_1077);
or U1102 (N_1102,N_1026,N_1033);
and U1103 (N_1103,N_1049,N_1022);
or U1104 (N_1104,N_1027,N_1031);
xnor U1105 (N_1105,N_1032,N_1072);
or U1106 (N_1106,N_1034,N_1046);
nor U1107 (N_1107,N_1057,N_1078);
or U1108 (N_1108,N_1024,N_1035);
or U1109 (N_1109,N_1076,N_1071);
or U1110 (N_1110,N_1067,N_1059);
nand U1111 (N_1111,N_1054,N_1034);
xnor U1112 (N_1112,N_1028,N_1047);
nor U1113 (N_1113,N_1029,N_1038);
or U1114 (N_1114,N_1063,N_1046);
xor U1115 (N_1115,N_1062,N_1046);
and U1116 (N_1116,N_1021,N_1037);
and U1117 (N_1117,N_1025,N_1035);
xor U1118 (N_1118,N_1021,N_1057);
or U1119 (N_1119,N_1077,N_1060);
xor U1120 (N_1120,N_1063,N_1072);
and U1121 (N_1121,N_1032,N_1054);
or U1122 (N_1122,N_1067,N_1051);
nor U1123 (N_1123,N_1027,N_1074);
xor U1124 (N_1124,N_1068,N_1030);
nand U1125 (N_1125,N_1053,N_1052);
xnor U1126 (N_1126,N_1052,N_1074);
nor U1127 (N_1127,N_1069,N_1031);
xnor U1128 (N_1128,N_1036,N_1043);
nor U1129 (N_1129,N_1069,N_1075);
xor U1130 (N_1130,N_1074,N_1069);
xor U1131 (N_1131,N_1023,N_1032);
and U1132 (N_1132,N_1030,N_1023);
nand U1133 (N_1133,N_1065,N_1025);
and U1134 (N_1134,N_1064,N_1044);
or U1135 (N_1135,N_1029,N_1020);
xor U1136 (N_1136,N_1023,N_1046);
and U1137 (N_1137,N_1063,N_1054);
nor U1138 (N_1138,N_1022,N_1034);
xnor U1139 (N_1139,N_1024,N_1025);
or U1140 (N_1140,N_1086,N_1112);
nor U1141 (N_1141,N_1114,N_1089);
nor U1142 (N_1142,N_1120,N_1087);
xnor U1143 (N_1143,N_1136,N_1085);
nor U1144 (N_1144,N_1097,N_1138);
or U1145 (N_1145,N_1101,N_1110);
or U1146 (N_1146,N_1129,N_1081);
or U1147 (N_1147,N_1119,N_1105);
nor U1148 (N_1148,N_1118,N_1133);
nand U1149 (N_1149,N_1109,N_1082);
and U1150 (N_1150,N_1093,N_1092);
nand U1151 (N_1151,N_1100,N_1080);
xor U1152 (N_1152,N_1139,N_1131);
nand U1153 (N_1153,N_1083,N_1121);
nand U1154 (N_1154,N_1132,N_1095);
and U1155 (N_1155,N_1125,N_1135);
xnor U1156 (N_1156,N_1134,N_1107);
or U1157 (N_1157,N_1106,N_1096);
and U1158 (N_1158,N_1116,N_1108);
or U1159 (N_1159,N_1130,N_1102);
xnor U1160 (N_1160,N_1111,N_1137);
xnor U1161 (N_1161,N_1123,N_1088);
or U1162 (N_1162,N_1128,N_1127);
or U1163 (N_1163,N_1099,N_1124);
or U1164 (N_1164,N_1122,N_1103);
nor U1165 (N_1165,N_1094,N_1126);
nor U1166 (N_1166,N_1091,N_1113);
or U1167 (N_1167,N_1090,N_1115);
or U1168 (N_1168,N_1084,N_1117);
nand U1169 (N_1169,N_1098,N_1104);
nand U1170 (N_1170,N_1109,N_1126);
xor U1171 (N_1171,N_1099,N_1135);
nor U1172 (N_1172,N_1128,N_1133);
nor U1173 (N_1173,N_1129,N_1125);
or U1174 (N_1174,N_1104,N_1100);
or U1175 (N_1175,N_1082,N_1136);
and U1176 (N_1176,N_1134,N_1115);
xnor U1177 (N_1177,N_1131,N_1111);
nand U1178 (N_1178,N_1098,N_1094);
and U1179 (N_1179,N_1101,N_1133);
or U1180 (N_1180,N_1125,N_1130);
xnor U1181 (N_1181,N_1110,N_1095);
xor U1182 (N_1182,N_1131,N_1136);
nor U1183 (N_1183,N_1089,N_1092);
or U1184 (N_1184,N_1128,N_1103);
nand U1185 (N_1185,N_1122,N_1115);
xnor U1186 (N_1186,N_1135,N_1121);
nor U1187 (N_1187,N_1103,N_1084);
and U1188 (N_1188,N_1133,N_1116);
xnor U1189 (N_1189,N_1083,N_1098);
and U1190 (N_1190,N_1093,N_1094);
nor U1191 (N_1191,N_1115,N_1104);
xor U1192 (N_1192,N_1086,N_1133);
or U1193 (N_1193,N_1109,N_1112);
or U1194 (N_1194,N_1120,N_1104);
nand U1195 (N_1195,N_1129,N_1080);
nand U1196 (N_1196,N_1106,N_1139);
or U1197 (N_1197,N_1107,N_1103);
nand U1198 (N_1198,N_1133,N_1105);
nor U1199 (N_1199,N_1103,N_1081);
and U1200 (N_1200,N_1198,N_1149);
and U1201 (N_1201,N_1154,N_1160);
nor U1202 (N_1202,N_1159,N_1170);
nand U1203 (N_1203,N_1178,N_1163);
and U1204 (N_1204,N_1153,N_1181);
nor U1205 (N_1205,N_1188,N_1140);
xnor U1206 (N_1206,N_1175,N_1151);
xnor U1207 (N_1207,N_1187,N_1141);
nand U1208 (N_1208,N_1145,N_1165);
and U1209 (N_1209,N_1157,N_1176);
and U1210 (N_1210,N_1180,N_1189);
and U1211 (N_1211,N_1174,N_1155);
or U1212 (N_1212,N_1168,N_1150);
or U1213 (N_1213,N_1190,N_1185);
xor U1214 (N_1214,N_1143,N_1142);
or U1215 (N_1215,N_1177,N_1172);
and U1216 (N_1216,N_1152,N_1183);
or U1217 (N_1217,N_1147,N_1173);
or U1218 (N_1218,N_1146,N_1166);
or U1219 (N_1219,N_1192,N_1169);
or U1220 (N_1220,N_1148,N_1191);
nor U1221 (N_1221,N_1182,N_1158);
nand U1222 (N_1222,N_1164,N_1199);
nand U1223 (N_1223,N_1195,N_1171);
xnor U1224 (N_1224,N_1186,N_1194);
and U1225 (N_1225,N_1193,N_1197);
and U1226 (N_1226,N_1184,N_1167);
nor U1227 (N_1227,N_1196,N_1161);
and U1228 (N_1228,N_1179,N_1144);
nand U1229 (N_1229,N_1162,N_1156);
xor U1230 (N_1230,N_1141,N_1146);
or U1231 (N_1231,N_1192,N_1187);
and U1232 (N_1232,N_1195,N_1192);
and U1233 (N_1233,N_1163,N_1185);
and U1234 (N_1234,N_1148,N_1163);
or U1235 (N_1235,N_1161,N_1167);
and U1236 (N_1236,N_1172,N_1155);
nand U1237 (N_1237,N_1152,N_1143);
or U1238 (N_1238,N_1176,N_1168);
and U1239 (N_1239,N_1178,N_1188);
and U1240 (N_1240,N_1199,N_1168);
xor U1241 (N_1241,N_1188,N_1180);
and U1242 (N_1242,N_1174,N_1146);
nand U1243 (N_1243,N_1182,N_1190);
and U1244 (N_1244,N_1151,N_1196);
or U1245 (N_1245,N_1152,N_1166);
nor U1246 (N_1246,N_1195,N_1176);
or U1247 (N_1247,N_1165,N_1188);
or U1248 (N_1248,N_1171,N_1165);
xor U1249 (N_1249,N_1193,N_1194);
nor U1250 (N_1250,N_1180,N_1187);
nor U1251 (N_1251,N_1172,N_1178);
xor U1252 (N_1252,N_1172,N_1141);
and U1253 (N_1253,N_1191,N_1179);
and U1254 (N_1254,N_1179,N_1168);
nand U1255 (N_1255,N_1175,N_1145);
nor U1256 (N_1256,N_1162,N_1196);
nor U1257 (N_1257,N_1160,N_1166);
nor U1258 (N_1258,N_1189,N_1196);
nor U1259 (N_1259,N_1175,N_1141);
nand U1260 (N_1260,N_1237,N_1218);
nand U1261 (N_1261,N_1249,N_1231);
or U1262 (N_1262,N_1251,N_1222);
xor U1263 (N_1263,N_1203,N_1255);
nor U1264 (N_1264,N_1239,N_1235);
or U1265 (N_1265,N_1240,N_1246);
or U1266 (N_1266,N_1209,N_1210);
nand U1267 (N_1267,N_1259,N_1213);
nand U1268 (N_1268,N_1225,N_1254);
nand U1269 (N_1269,N_1205,N_1232);
nor U1270 (N_1270,N_1212,N_1221);
nand U1271 (N_1271,N_1217,N_1236);
and U1272 (N_1272,N_1211,N_1223);
nand U1273 (N_1273,N_1238,N_1248);
or U1274 (N_1274,N_1252,N_1202);
nor U1275 (N_1275,N_1207,N_1220);
and U1276 (N_1276,N_1206,N_1253);
xnor U1277 (N_1277,N_1226,N_1219);
nor U1278 (N_1278,N_1204,N_1214);
and U1279 (N_1279,N_1208,N_1234);
xnor U1280 (N_1280,N_1215,N_1233);
or U1281 (N_1281,N_1228,N_1229);
and U1282 (N_1282,N_1227,N_1216);
or U1283 (N_1283,N_1256,N_1224);
xor U1284 (N_1284,N_1244,N_1200);
or U1285 (N_1285,N_1243,N_1245);
nor U1286 (N_1286,N_1250,N_1247);
nand U1287 (N_1287,N_1201,N_1242);
nor U1288 (N_1288,N_1241,N_1230);
xor U1289 (N_1289,N_1257,N_1258);
nand U1290 (N_1290,N_1250,N_1257);
xor U1291 (N_1291,N_1204,N_1244);
nand U1292 (N_1292,N_1246,N_1251);
or U1293 (N_1293,N_1248,N_1250);
and U1294 (N_1294,N_1212,N_1230);
and U1295 (N_1295,N_1206,N_1238);
nor U1296 (N_1296,N_1237,N_1239);
nand U1297 (N_1297,N_1243,N_1246);
nor U1298 (N_1298,N_1252,N_1216);
xor U1299 (N_1299,N_1254,N_1242);
and U1300 (N_1300,N_1213,N_1239);
xnor U1301 (N_1301,N_1254,N_1226);
nor U1302 (N_1302,N_1209,N_1204);
or U1303 (N_1303,N_1200,N_1251);
or U1304 (N_1304,N_1225,N_1257);
xor U1305 (N_1305,N_1215,N_1252);
xor U1306 (N_1306,N_1217,N_1226);
or U1307 (N_1307,N_1251,N_1239);
or U1308 (N_1308,N_1202,N_1253);
nor U1309 (N_1309,N_1237,N_1227);
nor U1310 (N_1310,N_1220,N_1236);
xor U1311 (N_1311,N_1249,N_1212);
xnor U1312 (N_1312,N_1237,N_1222);
xnor U1313 (N_1313,N_1202,N_1217);
nor U1314 (N_1314,N_1228,N_1256);
or U1315 (N_1315,N_1207,N_1212);
nor U1316 (N_1316,N_1232,N_1235);
nor U1317 (N_1317,N_1217,N_1200);
or U1318 (N_1318,N_1249,N_1208);
or U1319 (N_1319,N_1203,N_1256);
or U1320 (N_1320,N_1311,N_1272);
nand U1321 (N_1321,N_1264,N_1276);
and U1322 (N_1322,N_1290,N_1315);
xor U1323 (N_1323,N_1288,N_1306);
nand U1324 (N_1324,N_1261,N_1267);
xnor U1325 (N_1325,N_1287,N_1294);
and U1326 (N_1326,N_1309,N_1291);
xor U1327 (N_1327,N_1282,N_1275);
or U1328 (N_1328,N_1295,N_1273);
or U1329 (N_1329,N_1317,N_1293);
or U1330 (N_1330,N_1319,N_1266);
and U1331 (N_1331,N_1303,N_1296);
xor U1332 (N_1332,N_1299,N_1292);
or U1333 (N_1333,N_1314,N_1298);
nand U1334 (N_1334,N_1274,N_1278);
xnor U1335 (N_1335,N_1260,N_1286);
xnor U1336 (N_1336,N_1289,N_1270);
nor U1337 (N_1337,N_1302,N_1269);
or U1338 (N_1338,N_1310,N_1300);
and U1339 (N_1339,N_1304,N_1316);
nand U1340 (N_1340,N_1279,N_1265);
nor U1341 (N_1341,N_1312,N_1284);
and U1342 (N_1342,N_1285,N_1297);
or U1343 (N_1343,N_1263,N_1280);
and U1344 (N_1344,N_1307,N_1318);
nand U1345 (N_1345,N_1313,N_1308);
xnor U1346 (N_1346,N_1281,N_1271);
xnor U1347 (N_1347,N_1283,N_1301);
or U1348 (N_1348,N_1305,N_1268);
and U1349 (N_1349,N_1262,N_1277);
and U1350 (N_1350,N_1299,N_1293);
xnor U1351 (N_1351,N_1293,N_1273);
xor U1352 (N_1352,N_1315,N_1273);
and U1353 (N_1353,N_1266,N_1265);
or U1354 (N_1354,N_1277,N_1289);
or U1355 (N_1355,N_1308,N_1309);
xnor U1356 (N_1356,N_1291,N_1285);
nor U1357 (N_1357,N_1292,N_1267);
nor U1358 (N_1358,N_1286,N_1290);
or U1359 (N_1359,N_1303,N_1312);
or U1360 (N_1360,N_1276,N_1275);
xor U1361 (N_1361,N_1305,N_1265);
and U1362 (N_1362,N_1267,N_1284);
nor U1363 (N_1363,N_1313,N_1311);
and U1364 (N_1364,N_1314,N_1283);
and U1365 (N_1365,N_1294,N_1293);
nand U1366 (N_1366,N_1291,N_1302);
nand U1367 (N_1367,N_1274,N_1284);
nand U1368 (N_1368,N_1268,N_1304);
or U1369 (N_1369,N_1308,N_1284);
nor U1370 (N_1370,N_1264,N_1297);
nand U1371 (N_1371,N_1285,N_1278);
nand U1372 (N_1372,N_1297,N_1298);
or U1373 (N_1373,N_1278,N_1312);
nor U1374 (N_1374,N_1287,N_1312);
nand U1375 (N_1375,N_1303,N_1311);
nor U1376 (N_1376,N_1278,N_1303);
xor U1377 (N_1377,N_1298,N_1290);
nor U1378 (N_1378,N_1277,N_1317);
or U1379 (N_1379,N_1311,N_1305);
or U1380 (N_1380,N_1347,N_1352);
nand U1381 (N_1381,N_1338,N_1369);
and U1382 (N_1382,N_1328,N_1366);
or U1383 (N_1383,N_1374,N_1348);
and U1384 (N_1384,N_1327,N_1376);
xor U1385 (N_1385,N_1365,N_1337);
xor U1386 (N_1386,N_1379,N_1344);
nor U1387 (N_1387,N_1377,N_1364);
nand U1388 (N_1388,N_1362,N_1346);
and U1389 (N_1389,N_1368,N_1371);
and U1390 (N_1390,N_1378,N_1326);
xnor U1391 (N_1391,N_1329,N_1343);
nand U1392 (N_1392,N_1320,N_1330);
xor U1393 (N_1393,N_1357,N_1321);
and U1394 (N_1394,N_1353,N_1360);
or U1395 (N_1395,N_1367,N_1332);
nand U1396 (N_1396,N_1345,N_1331);
nand U1397 (N_1397,N_1372,N_1333);
or U1398 (N_1398,N_1325,N_1342);
or U1399 (N_1399,N_1361,N_1340);
and U1400 (N_1400,N_1335,N_1373);
and U1401 (N_1401,N_1323,N_1334);
nand U1402 (N_1402,N_1370,N_1339);
nor U1403 (N_1403,N_1355,N_1358);
xor U1404 (N_1404,N_1375,N_1359);
and U1405 (N_1405,N_1356,N_1351);
nand U1406 (N_1406,N_1350,N_1341);
and U1407 (N_1407,N_1324,N_1363);
xnor U1408 (N_1408,N_1354,N_1322);
xor U1409 (N_1409,N_1336,N_1349);
or U1410 (N_1410,N_1359,N_1367);
or U1411 (N_1411,N_1376,N_1360);
xor U1412 (N_1412,N_1377,N_1338);
xnor U1413 (N_1413,N_1328,N_1362);
and U1414 (N_1414,N_1320,N_1359);
nor U1415 (N_1415,N_1349,N_1358);
or U1416 (N_1416,N_1329,N_1358);
or U1417 (N_1417,N_1323,N_1345);
and U1418 (N_1418,N_1360,N_1340);
xnor U1419 (N_1419,N_1345,N_1340);
and U1420 (N_1420,N_1377,N_1359);
xnor U1421 (N_1421,N_1358,N_1351);
nor U1422 (N_1422,N_1353,N_1365);
nor U1423 (N_1423,N_1361,N_1372);
and U1424 (N_1424,N_1337,N_1357);
and U1425 (N_1425,N_1369,N_1339);
xor U1426 (N_1426,N_1337,N_1368);
nor U1427 (N_1427,N_1333,N_1355);
and U1428 (N_1428,N_1344,N_1329);
nor U1429 (N_1429,N_1377,N_1332);
xor U1430 (N_1430,N_1338,N_1330);
nand U1431 (N_1431,N_1349,N_1343);
and U1432 (N_1432,N_1327,N_1348);
nor U1433 (N_1433,N_1354,N_1321);
or U1434 (N_1434,N_1362,N_1322);
and U1435 (N_1435,N_1356,N_1331);
or U1436 (N_1436,N_1362,N_1337);
or U1437 (N_1437,N_1325,N_1321);
xor U1438 (N_1438,N_1322,N_1343);
nand U1439 (N_1439,N_1324,N_1332);
and U1440 (N_1440,N_1432,N_1386);
nand U1441 (N_1441,N_1381,N_1435);
xor U1442 (N_1442,N_1404,N_1416);
and U1443 (N_1443,N_1439,N_1427);
xnor U1444 (N_1444,N_1420,N_1383);
or U1445 (N_1445,N_1385,N_1419);
and U1446 (N_1446,N_1423,N_1396);
or U1447 (N_1447,N_1399,N_1407);
and U1448 (N_1448,N_1411,N_1390);
and U1449 (N_1449,N_1394,N_1410);
or U1450 (N_1450,N_1418,N_1406);
and U1451 (N_1451,N_1391,N_1433);
xor U1452 (N_1452,N_1438,N_1403);
nand U1453 (N_1453,N_1436,N_1387);
nand U1454 (N_1454,N_1429,N_1389);
and U1455 (N_1455,N_1398,N_1428);
xor U1456 (N_1456,N_1425,N_1424);
nor U1457 (N_1457,N_1405,N_1414);
or U1458 (N_1458,N_1400,N_1437);
and U1459 (N_1459,N_1392,N_1413);
and U1460 (N_1460,N_1393,N_1401);
nand U1461 (N_1461,N_1430,N_1384);
nor U1462 (N_1462,N_1395,N_1380);
nor U1463 (N_1463,N_1408,N_1397);
xnor U1464 (N_1464,N_1412,N_1426);
nor U1465 (N_1465,N_1431,N_1415);
and U1466 (N_1466,N_1382,N_1434);
nor U1467 (N_1467,N_1422,N_1409);
or U1468 (N_1468,N_1388,N_1421);
nand U1469 (N_1469,N_1417,N_1402);
nor U1470 (N_1470,N_1391,N_1413);
or U1471 (N_1471,N_1418,N_1380);
nor U1472 (N_1472,N_1413,N_1411);
and U1473 (N_1473,N_1439,N_1430);
or U1474 (N_1474,N_1431,N_1395);
and U1475 (N_1475,N_1414,N_1415);
nand U1476 (N_1476,N_1417,N_1431);
nand U1477 (N_1477,N_1383,N_1402);
nand U1478 (N_1478,N_1400,N_1407);
or U1479 (N_1479,N_1406,N_1384);
xnor U1480 (N_1480,N_1399,N_1418);
xnor U1481 (N_1481,N_1406,N_1383);
xnor U1482 (N_1482,N_1436,N_1393);
nand U1483 (N_1483,N_1403,N_1406);
nor U1484 (N_1484,N_1396,N_1427);
nor U1485 (N_1485,N_1423,N_1436);
or U1486 (N_1486,N_1382,N_1380);
xor U1487 (N_1487,N_1408,N_1413);
nor U1488 (N_1488,N_1419,N_1408);
xor U1489 (N_1489,N_1414,N_1406);
and U1490 (N_1490,N_1426,N_1417);
xor U1491 (N_1491,N_1420,N_1405);
xor U1492 (N_1492,N_1411,N_1436);
nand U1493 (N_1493,N_1418,N_1423);
nand U1494 (N_1494,N_1429,N_1438);
or U1495 (N_1495,N_1384,N_1426);
or U1496 (N_1496,N_1408,N_1401);
and U1497 (N_1497,N_1392,N_1407);
xnor U1498 (N_1498,N_1399,N_1401);
nor U1499 (N_1499,N_1415,N_1389);
and U1500 (N_1500,N_1451,N_1474);
and U1501 (N_1501,N_1456,N_1492);
nor U1502 (N_1502,N_1482,N_1472);
xnor U1503 (N_1503,N_1449,N_1480);
or U1504 (N_1504,N_1445,N_1459);
or U1505 (N_1505,N_1442,N_1447);
nor U1506 (N_1506,N_1462,N_1479);
nor U1507 (N_1507,N_1494,N_1481);
and U1508 (N_1508,N_1477,N_1478);
and U1509 (N_1509,N_1499,N_1453);
and U1510 (N_1510,N_1448,N_1469);
or U1511 (N_1511,N_1443,N_1496);
or U1512 (N_1512,N_1486,N_1490);
nand U1513 (N_1513,N_1452,N_1497);
nand U1514 (N_1514,N_1457,N_1441);
nor U1515 (N_1515,N_1475,N_1468);
and U1516 (N_1516,N_1489,N_1467);
or U1517 (N_1517,N_1493,N_1440);
nor U1518 (N_1518,N_1458,N_1495);
or U1519 (N_1519,N_1444,N_1476);
or U1520 (N_1520,N_1488,N_1471);
xnor U1521 (N_1521,N_1485,N_1460);
nor U1522 (N_1522,N_1498,N_1450);
xor U1523 (N_1523,N_1464,N_1470);
nand U1524 (N_1524,N_1463,N_1484);
xor U1525 (N_1525,N_1491,N_1461);
nor U1526 (N_1526,N_1455,N_1454);
nand U1527 (N_1527,N_1483,N_1487);
or U1528 (N_1528,N_1446,N_1473);
nand U1529 (N_1529,N_1465,N_1466);
nor U1530 (N_1530,N_1497,N_1445);
or U1531 (N_1531,N_1490,N_1461);
nand U1532 (N_1532,N_1455,N_1479);
xor U1533 (N_1533,N_1471,N_1440);
nand U1534 (N_1534,N_1461,N_1464);
and U1535 (N_1535,N_1441,N_1469);
or U1536 (N_1536,N_1456,N_1468);
or U1537 (N_1537,N_1440,N_1458);
xor U1538 (N_1538,N_1479,N_1468);
xnor U1539 (N_1539,N_1490,N_1499);
nor U1540 (N_1540,N_1442,N_1498);
xnor U1541 (N_1541,N_1456,N_1491);
nor U1542 (N_1542,N_1477,N_1442);
xor U1543 (N_1543,N_1473,N_1443);
nand U1544 (N_1544,N_1442,N_1467);
xnor U1545 (N_1545,N_1466,N_1489);
and U1546 (N_1546,N_1468,N_1442);
nor U1547 (N_1547,N_1487,N_1479);
or U1548 (N_1548,N_1448,N_1450);
or U1549 (N_1549,N_1476,N_1449);
or U1550 (N_1550,N_1469,N_1475);
nor U1551 (N_1551,N_1482,N_1481);
nand U1552 (N_1552,N_1469,N_1472);
xor U1553 (N_1553,N_1487,N_1470);
nand U1554 (N_1554,N_1446,N_1482);
nand U1555 (N_1555,N_1496,N_1475);
nor U1556 (N_1556,N_1449,N_1481);
or U1557 (N_1557,N_1443,N_1490);
xnor U1558 (N_1558,N_1498,N_1481);
nand U1559 (N_1559,N_1441,N_1463);
and U1560 (N_1560,N_1506,N_1514);
nand U1561 (N_1561,N_1510,N_1550);
or U1562 (N_1562,N_1555,N_1558);
xnor U1563 (N_1563,N_1539,N_1549);
or U1564 (N_1564,N_1552,N_1518);
nor U1565 (N_1565,N_1544,N_1532);
or U1566 (N_1566,N_1526,N_1504);
xor U1567 (N_1567,N_1540,N_1547);
and U1568 (N_1568,N_1507,N_1538);
or U1569 (N_1569,N_1522,N_1503);
and U1570 (N_1570,N_1529,N_1533);
xor U1571 (N_1571,N_1545,N_1548);
nor U1572 (N_1572,N_1517,N_1505);
nor U1573 (N_1573,N_1534,N_1536);
and U1574 (N_1574,N_1501,N_1537);
xor U1575 (N_1575,N_1520,N_1541);
nor U1576 (N_1576,N_1551,N_1500);
or U1577 (N_1577,N_1508,N_1509);
or U1578 (N_1578,N_1511,N_1516);
nor U1579 (N_1579,N_1528,N_1535);
xor U1580 (N_1580,N_1527,N_1530);
nand U1581 (N_1581,N_1542,N_1553);
nor U1582 (N_1582,N_1546,N_1502);
nor U1583 (N_1583,N_1556,N_1557);
nand U1584 (N_1584,N_1513,N_1519);
and U1585 (N_1585,N_1554,N_1559);
nor U1586 (N_1586,N_1524,N_1523);
xor U1587 (N_1587,N_1525,N_1512);
and U1588 (N_1588,N_1543,N_1515);
xnor U1589 (N_1589,N_1521,N_1531);
nor U1590 (N_1590,N_1508,N_1533);
or U1591 (N_1591,N_1509,N_1544);
nor U1592 (N_1592,N_1536,N_1517);
or U1593 (N_1593,N_1554,N_1531);
nor U1594 (N_1594,N_1502,N_1500);
and U1595 (N_1595,N_1543,N_1502);
or U1596 (N_1596,N_1524,N_1532);
and U1597 (N_1597,N_1557,N_1551);
and U1598 (N_1598,N_1549,N_1524);
nand U1599 (N_1599,N_1505,N_1544);
or U1600 (N_1600,N_1550,N_1532);
nor U1601 (N_1601,N_1515,N_1522);
and U1602 (N_1602,N_1548,N_1534);
or U1603 (N_1603,N_1504,N_1556);
nand U1604 (N_1604,N_1527,N_1547);
nand U1605 (N_1605,N_1503,N_1512);
or U1606 (N_1606,N_1545,N_1518);
and U1607 (N_1607,N_1503,N_1511);
or U1608 (N_1608,N_1556,N_1555);
xnor U1609 (N_1609,N_1521,N_1553);
and U1610 (N_1610,N_1544,N_1548);
nor U1611 (N_1611,N_1509,N_1525);
nor U1612 (N_1612,N_1511,N_1544);
or U1613 (N_1613,N_1503,N_1528);
or U1614 (N_1614,N_1507,N_1550);
nand U1615 (N_1615,N_1544,N_1500);
nand U1616 (N_1616,N_1543,N_1545);
or U1617 (N_1617,N_1505,N_1532);
xor U1618 (N_1618,N_1547,N_1545);
nor U1619 (N_1619,N_1531,N_1520);
xor U1620 (N_1620,N_1613,N_1582);
nor U1621 (N_1621,N_1604,N_1574);
nor U1622 (N_1622,N_1594,N_1569);
or U1623 (N_1623,N_1596,N_1581);
xnor U1624 (N_1624,N_1571,N_1560);
nor U1625 (N_1625,N_1602,N_1576);
nor U1626 (N_1626,N_1609,N_1587);
xor U1627 (N_1627,N_1589,N_1591);
nand U1628 (N_1628,N_1585,N_1603);
nand U1629 (N_1629,N_1617,N_1605);
nor U1630 (N_1630,N_1598,N_1599);
nor U1631 (N_1631,N_1597,N_1606);
and U1632 (N_1632,N_1612,N_1563);
xnor U1633 (N_1633,N_1567,N_1570);
or U1634 (N_1634,N_1595,N_1607);
xnor U1635 (N_1635,N_1565,N_1566);
nor U1636 (N_1636,N_1601,N_1615);
xor U1637 (N_1637,N_1618,N_1561);
nand U1638 (N_1638,N_1580,N_1592);
or U1639 (N_1639,N_1575,N_1590);
xnor U1640 (N_1640,N_1614,N_1588);
nor U1641 (N_1641,N_1579,N_1568);
and U1642 (N_1642,N_1573,N_1583);
nand U1643 (N_1643,N_1610,N_1562);
or U1644 (N_1644,N_1616,N_1600);
nor U1645 (N_1645,N_1584,N_1611);
nor U1646 (N_1646,N_1577,N_1586);
xnor U1647 (N_1647,N_1564,N_1572);
nor U1648 (N_1648,N_1578,N_1593);
or U1649 (N_1649,N_1608,N_1619);
and U1650 (N_1650,N_1602,N_1575);
xnor U1651 (N_1651,N_1589,N_1572);
nand U1652 (N_1652,N_1609,N_1611);
and U1653 (N_1653,N_1578,N_1605);
xnor U1654 (N_1654,N_1587,N_1602);
nor U1655 (N_1655,N_1576,N_1578);
nand U1656 (N_1656,N_1615,N_1597);
nand U1657 (N_1657,N_1565,N_1596);
and U1658 (N_1658,N_1596,N_1609);
nand U1659 (N_1659,N_1588,N_1603);
nor U1660 (N_1660,N_1619,N_1591);
nor U1661 (N_1661,N_1592,N_1573);
nor U1662 (N_1662,N_1584,N_1598);
and U1663 (N_1663,N_1607,N_1593);
nand U1664 (N_1664,N_1614,N_1580);
and U1665 (N_1665,N_1576,N_1619);
and U1666 (N_1666,N_1606,N_1611);
xor U1667 (N_1667,N_1611,N_1589);
xor U1668 (N_1668,N_1616,N_1578);
or U1669 (N_1669,N_1603,N_1605);
or U1670 (N_1670,N_1613,N_1578);
xor U1671 (N_1671,N_1562,N_1611);
or U1672 (N_1672,N_1583,N_1588);
nand U1673 (N_1673,N_1580,N_1603);
or U1674 (N_1674,N_1597,N_1572);
or U1675 (N_1675,N_1586,N_1578);
nor U1676 (N_1676,N_1612,N_1588);
xnor U1677 (N_1677,N_1564,N_1591);
and U1678 (N_1678,N_1573,N_1562);
nand U1679 (N_1679,N_1573,N_1563);
and U1680 (N_1680,N_1621,N_1677);
xor U1681 (N_1681,N_1676,N_1623);
and U1682 (N_1682,N_1674,N_1653);
and U1683 (N_1683,N_1652,N_1630);
xnor U1684 (N_1684,N_1631,N_1679);
nand U1685 (N_1685,N_1647,N_1661);
nor U1686 (N_1686,N_1642,N_1669);
nand U1687 (N_1687,N_1646,N_1651);
and U1688 (N_1688,N_1626,N_1672);
and U1689 (N_1689,N_1633,N_1657);
nor U1690 (N_1690,N_1649,N_1643);
nor U1691 (N_1691,N_1666,N_1671);
nand U1692 (N_1692,N_1629,N_1665);
nor U1693 (N_1693,N_1662,N_1628);
or U1694 (N_1694,N_1659,N_1620);
xor U1695 (N_1695,N_1678,N_1660);
or U1696 (N_1696,N_1639,N_1637);
and U1697 (N_1697,N_1624,N_1638);
or U1698 (N_1698,N_1675,N_1634);
nor U1699 (N_1699,N_1632,N_1667);
xnor U1700 (N_1700,N_1648,N_1627);
nor U1701 (N_1701,N_1645,N_1655);
nor U1702 (N_1702,N_1622,N_1670);
or U1703 (N_1703,N_1625,N_1650);
xnor U1704 (N_1704,N_1636,N_1635);
xor U1705 (N_1705,N_1668,N_1656);
nand U1706 (N_1706,N_1654,N_1641);
nand U1707 (N_1707,N_1644,N_1663);
xor U1708 (N_1708,N_1640,N_1673);
nand U1709 (N_1709,N_1658,N_1664);
and U1710 (N_1710,N_1622,N_1639);
nor U1711 (N_1711,N_1659,N_1634);
nand U1712 (N_1712,N_1637,N_1642);
xnor U1713 (N_1713,N_1655,N_1657);
nand U1714 (N_1714,N_1622,N_1626);
or U1715 (N_1715,N_1647,N_1649);
and U1716 (N_1716,N_1626,N_1655);
and U1717 (N_1717,N_1679,N_1633);
xnor U1718 (N_1718,N_1671,N_1625);
nand U1719 (N_1719,N_1663,N_1624);
nor U1720 (N_1720,N_1639,N_1661);
or U1721 (N_1721,N_1675,N_1649);
and U1722 (N_1722,N_1627,N_1674);
and U1723 (N_1723,N_1651,N_1657);
xnor U1724 (N_1724,N_1675,N_1625);
or U1725 (N_1725,N_1662,N_1671);
nand U1726 (N_1726,N_1654,N_1630);
or U1727 (N_1727,N_1642,N_1651);
or U1728 (N_1728,N_1626,N_1657);
or U1729 (N_1729,N_1676,N_1675);
nor U1730 (N_1730,N_1660,N_1676);
xor U1731 (N_1731,N_1671,N_1636);
and U1732 (N_1732,N_1623,N_1624);
or U1733 (N_1733,N_1661,N_1628);
nand U1734 (N_1734,N_1625,N_1634);
xnor U1735 (N_1735,N_1628,N_1633);
nor U1736 (N_1736,N_1637,N_1660);
xnor U1737 (N_1737,N_1670,N_1655);
nand U1738 (N_1738,N_1677,N_1659);
and U1739 (N_1739,N_1632,N_1640);
and U1740 (N_1740,N_1708,N_1735);
or U1741 (N_1741,N_1686,N_1706);
or U1742 (N_1742,N_1728,N_1702);
or U1743 (N_1743,N_1725,N_1685);
nor U1744 (N_1744,N_1721,N_1704);
nand U1745 (N_1745,N_1682,N_1699);
nand U1746 (N_1746,N_1734,N_1738);
nand U1747 (N_1747,N_1698,N_1707);
nor U1748 (N_1748,N_1695,N_1692);
xor U1749 (N_1749,N_1694,N_1689);
nor U1750 (N_1750,N_1723,N_1693);
and U1751 (N_1751,N_1729,N_1705);
nand U1752 (N_1752,N_1700,N_1711);
xnor U1753 (N_1753,N_1736,N_1731);
nand U1754 (N_1754,N_1720,N_1733);
xnor U1755 (N_1755,N_1701,N_1710);
nand U1756 (N_1756,N_1696,N_1709);
nor U1757 (N_1757,N_1739,N_1718);
nand U1758 (N_1758,N_1714,N_1715);
xnor U1759 (N_1759,N_1730,N_1690);
or U1760 (N_1760,N_1697,N_1703);
and U1761 (N_1761,N_1737,N_1688);
and U1762 (N_1762,N_1683,N_1712);
nor U1763 (N_1763,N_1726,N_1719);
and U1764 (N_1764,N_1724,N_1680);
or U1765 (N_1765,N_1713,N_1722);
nand U1766 (N_1766,N_1684,N_1687);
nand U1767 (N_1767,N_1681,N_1727);
nand U1768 (N_1768,N_1716,N_1691);
nor U1769 (N_1769,N_1717,N_1732);
and U1770 (N_1770,N_1680,N_1694);
nand U1771 (N_1771,N_1731,N_1726);
or U1772 (N_1772,N_1710,N_1708);
nand U1773 (N_1773,N_1715,N_1721);
and U1774 (N_1774,N_1734,N_1720);
nand U1775 (N_1775,N_1680,N_1712);
or U1776 (N_1776,N_1730,N_1694);
nor U1777 (N_1777,N_1719,N_1680);
nand U1778 (N_1778,N_1724,N_1690);
xnor U1779 (N_1779,N_1703,N_1732);
nand U1780 (N_1780,N_1685,N_1692);
and U1781 (N_1781,N_1682,N_1695);
nand U1782 (N_1782,N_1687,N_1704);
or U1783 (N_1783,N_1711,N_1689);
nor U1784 (N_1784,N_1728,N_1717);
and U1785 (N_1785,N_1708,N_1697);
or U1786 (N_1786,N_1691,N_1730);
nor U1787 (N_1787,N_1712,N_1695);
or U1788 (N_1788,N_1688,N_1728);
nor U1789 (N_1789,N_1721,N_1716);
and U1790 (N_1790,N_1697,N_1734);
xnor U1791 (N_1791,N_1710,N_1704);
and U1792 (N_1792,N_1728,N_1729);
or U1793 (N_1793,N_1698,N_1706);
nand U1794 (N_1794,N_1690,N_1680);
and U1795 (N_1795,N_1687,N_1737);
and U1796 (N_1796,N_1713,N_1714);
xor U1797 (N_1797,N_1701,N_1705);
and U1798 (N_1798,N_1731,N_1685);
nor U1799 (N_1799,N_1732,N_1692);
nand U1800 (N_1800,N_1783,N_1784);
nor U1801 (N_1801,N_1794,N_1756);
xnor U1802 (N_1802,N_1785,N_1742);
nor U1803 (N_1803,N_1768,N_1757);
nor U1804 (N_1804,N_1795,N_1771);
nand U1805 (N_1805,N_1760,N_1797);
nor U1806 (N_1806,N_1767,N_1751);
nor U1807 (N_1807,N_1799,N_1777);
nor U1808 (N_1808,N_1745,N_1779);
or U1809 (N_1809,N_1781,N_1793);
and U1810 (N_1810,N_1749,N_1778);
nor U1811 (N_1811,N_1765,N_1762);
nor U1812 (N_1812,N_1755,N_1753);
and U1813 (N_1813,N_1741,N_1740);
and U1814 (N_1814,N_1774,N_1789);
or U1815 (N_1815,N_1792,N_1796);
and U1816 (N_1816,N_1759,N_1769);
nand U1817 (N_1817,N_1752,N_1791);
nor U1818 (N_1818,N_1750,N_1770);
xnor U1819 (N_1819,N_1754,N_1748);
nor U1820 (N_1820,N_1758,N_1772);
or U1821 (N_1821,N_1788,N_1764);
or U1822 (N_1822,N_1780,N_1746);
nor U1823 (N_1823,N_1775,N_1786);
nor U1824 (N_1824,N_1773,N_1744);
and U1825 (N_1825,N_1766,N_1763);
nand U1826 (N_1826,N_1761,N_1798);
nand U1827 (N_1827,N_1747,N_1776);
xor U1828 (N_1828,N_1787,N_1782);
and U1829 (N_1829,N_1743,N_1790);
nor U1830 (N_1830,N_1764,N_1742);
nand U1831 (N_1831,N_1793,N_1782);
xor U1832 (N_1832,N_1768,N_1767);
and U1833 (N_1833,N_1790,N_1774);
nand U1834 (N_1834,N_1788,N_1772);
nor U1835 (N_1835,N_1762,N_1787);
nand U1836 (N_1836,N_1786,N_1752);
nor U1837 (N_1837,N_1778,N_1755);
nor U1838 (N_1838,N_1766,N_1764);
nand U1839 (N_1839,N_1743,N_1746);
and U1840 (N_1840,N_1741,N_1749);
xnor U1841 (N_1841,N_1751,N_1794);
or U1842 (N_1842,N_1759,N_1742);
xnor U1843 (N_1843,N_1795,N_1781);
nor U1844 (N_1844,N_1771,N_1765);
and U1845 (N_1845,N_1757,N_1786);
and U1846 (N_1846,N_1795,N_1785);
and U1847 (N_1847,N_1799,N_1788);
nand U1848 (N_1848,N_1788,N_1747);
or U1849 (N_1849,N_1767,N_1749);
or U1850 (N_1850,N_1786,N_1784);
or U1851 (N_1851,N_1768,N_1766);
and U1852 (N_1852,N_1767,N_1798);
nand U1853 (N_1853,N_1746,N_1757);
nand U1854 (N_1854,N_1759,N_1743);
nor U1855 (N_1855,N_1749,N_1799);
xnor U1856 (N_1856,N_1763,N_1788);
or U1857 (N_1857,N_1783,N_1792);
or U1858 (N_1858,N_1772,N_1774);
or U1859 (N_1859,N_1781,N_1746);
nand U1860 (N_1860,N_1849,N_1835);
nor U1861 (N_1861,N_1818,N_1857);
or U1862 (N_1862,N_1814,N_1847);
nor U1863 (N_1863,N_1824,N_1810);
nor U1864 (N_1864,N_1805,N_1856);
or U1865 (N_1865,N_1833,N_1832);
and U1866 (N_1866,N_1840,N_1811);
nor U1867 (N_1867,N_1841,N_1853);
and U1868 (N_1868,N_1844,N_1808);
nand U1869 (N_1869,N_1801,N_1826);
or U1870 (N_1870,N_1851,N_1804);
xnor U1871 (N_1871,N_1825,N_1854);
and U1872 (N_1872,N_1842,N_1828);
nand U1873 (N_1873,N_1839,N_1850);
nand U1874 (N_1874,N_1829,N_1803);
nor U1875 (N_1875,N_1831,N_1816);
nor U1876 (N_1876,N_1830,N_1813);
and U1877 (N_1877,N_1843,N_1838);
nor U1878 (N_1878,N_1852,N_1817);
xnor U1879 (N_1879,N_1819,N_1858);
and U1880 (N_1880,N_1821,N_1800);
or U1881 (N_1881,N_1809,N_1855);
nor U1882 (N_1882,N_1827,N_1823);
and U1883 (N_1883,N_1846,N_1820);
nor U1884 (N_1884,N_1859,N_1845);
nor U1885 (N_1885,N_1822,N_1815);
xnor U1886 (N_1886,N_1837,N_1834);
and U1887 (N_1887,N_1807,N_1812);
nand U1888 (N_1888,N_1848,N_1806);
or U1889 (N_1889,N_1836,N_1802);
xor U1890 (N_1890,N_1831,N_1828);
nand U1891 (N_1891,N_1844,N_1826);
xor U1892 (N_1892,N_1852,N_1824);
and U1893 (N_1893,N_1831,N_1839);
and U1894 (N_1894,N_1816,N_1855);
and U1895 (N_1895,N_1845,N_1821);
nor U1896 (N_1896,N_1802,N_1827);
and U1897 (N_1897,N_1858,N_1820);
xor U1898 (N_1898,N_1859,N_1856);
nor U1899 (N_1899,N_1842,N_1845);
or U1900 (N_1900,N_1804,N_1801);
nor U1901 (N_1901,N_1818,N_1836);
or U1902 (N_1902,N_1817,N_1838);
xnor U1903 (N_1903,N_1823,N_1830);
nor U1904 (N_1904,N_1841,N_1839);
nand U1905 (N_1905,N_1839,N_1825);
or U1906 (N_1906,N_1827,N_1844);
or U1907 (N_1907,N_1843,N_1831);
or U1908 (N_1908,N_1821,N_1831);
or U1909 (N_1909,N_1846,N_1838);
xor U1910 (N_1910,N_1810,N_1825);
nand U1911 (N_1911,N_1835,N_1827);
nand U1912 (N_1912,N_1819,N_1856);
and U1913 (N_1913,N_1815,N_1839);
nand U1914 (N_1914,N_1817,N_1801);
or U1915 (N_1915,N_1822,N_1840);
or U1916 (N_1916,N_1808,N_1811);
and U1917 (N_1917,N_1826,N_1812);
and U1918 (N_1918,N_1820,N_1808);
nor U1919 (N_1919,N_1821,N_1830);
xor U1920 (N_1920,N_1880,N_1867);
or U1921 (N_1921,N_1883,N_1884);
and U1922 (N_1922,N_1892,N_1903);
nand U1923 (N_1923,N_1909,N_1870);
or U1924 (N_1924,N_1876,N_1910);
or U1925 (N_1925,N_1899,N_1887);
nor U1926 (N_1926,N_1906,N_1898);
nand U1927 (N_1927,N_1917,N_1860);
and U1928 (N_1928,N_1911,N_1919);
and U1929 (N_1929,N_1863,N_1913);
or U1930 (N_1930,N_1864,N_1885);
and U1931 (N_1931,N_1894,N_1895);
nand U1932 (N_1932,N_1877,N_1879);
xnor U1933 (N_1933,N_1886,N_1914);
and U1934 (N_1934,N_1908,N_1900);
xnor U1935 (N_1935,N_1874,N_1878);
nand U1936 (N_1936,N_1868,N_1897);
nor U1937 (N_1937,N_1875,N_1893);
nand U1938 (N_1938,N_1861,N_1888);
or U1939 (N_1939,N_1916,N_1872);
xnor U1940 (N_1940,N_1873,N_1866);
xnor U1941 (N_1941,N_1896,N_1912);
and U1942 (N_1942,N_1862,N_1890);
or U1943 (N_1943,N_1905,N_1907);
nor U1944 (N_1944,N_1871,N_1918);
nand U1945 (N_1945,N_1902,N_1901);
xnor U1946 (N_1946,N_1869,N_1904);
and U1947 (N_1947,N_1915,N_1891);
nor U1948 (N_1948,N_1882,N_1881);
and U1949 (N_1949,N_1889,N_1865);
xor U1950 (N_1950,N_1895,N_1908);
or U1951 (N_1951,N_1904,N_1875);
nor U1952 (N_1952,N_1909,N_1919);
or U1953 (N_1953,N_1914,N_1901);
and U1954 (N_1954,N_1903,N_1901);
nand U1955 (N_1955,N_1885,N_1893);
xnor U1956 (N_1956,N_1919,N_1915);
and U1957 (N_1957,N_1910,N_1904);
nand U1958 (N_1958,N_1890,N_1885);
nand U1959 (N_1959,N_1908,N_1915);
or U1960 (N_1960,N_1864,N_1919);
nand U1961 (N_1961,N_1889,N_1905);
nor U1962 (N_1962,N_1878,N_1914);
xnor U1963 (N_1963,N_1873,N_1906);
nor U1964 (N_1964,N_1881,N_1911);
xor U1965 (N_1965,N_1898,N_1873);
or U1966 (N_1966,N_1912,N_1877);
or U1967 (N_1967,N_1874,N_1891);
or U1968 (N_1968,N_1899,N_1868);
and U1969 (N_1969,N_1863,N_1862);
xor U1970 (N_1970,N_1880,N_1862);
or U1971 (N_1971,N_1902,N_1906);
nor U1972 (N_1972,N_1878,N_1889);
nor U1973 (N_1973,N_1897,N_1915);
nor U1974 (N_1974,N_1906,N_1871);
or U1975 (N_1975,N_1902,N_1870);
nor U1976 (N_1976,N_1892,N_1889);
or U1977 (N_1977,N_1869,N_1887);
xor U1978 (N_1978,N_1864,N_1879);
or U1979 (N_1979,N_1885,N_1904);
nand U1980 (N_1980,N_1953,N_1934);
nand U1981 (N_1981,N_1966,N_1931);
and U1982 (N_1982,N_1962,N_1975);
nor U1983 (N_1983,N_1948,N_1963);
or U1984 (N_1984,N_1923,N_1951);
nand U1985 (N_1985,N_1946,N_1921);
nand U1986 (N_1986,N_1969,N_1936);
nand U1987 (N_1987,N_1973,N_1943);
nand U1988 (N_1988,N_1935,N_1949);
nand U1989 (N_1989,N_1957,N_1945);
nand U1990 (N_1990,N_1937,N_1942);
and U1991 (N_1991,N_1979,N_1968);
nand U1992 (N_1992,N_1932,N_1956);
and U1993 (N_1993,N_1955,N_1933);
nand U1994 (N_1994,N_1950,N_1960);
nand U1995 (N_1995,N_1972,N_1967);
and U1996 (N_1996,N_1971,N_1924);
nor U1997 (N_1997,N_1925,N_1939);
nor U1998 (N_1998,N_1964,N_1940);
or U1999 (N_1999,N_1961,N_1970);
and U2000 (N_2000,N_1954,N_1976);
nand U2001 (N_2001,N_1938,N_1926);
nand U2002 (N_2002,N_1977,N_1965);
nand U2003 (N_2003,N_1929,N_1920);
nor U2004 (N_2004,N_1941,N_1952);
or U2005 (N_2005,N_1927,N_1922);
and U2006 (N_2006,N_1978,N_1974);
or U2007 (N_2007,N_1958,N_1959);
nor U2008 (N_2008,N_1928,N_1944);
nor U2009 (N_2009,N_1930,N_1947);
nand U2010 (N_2010,N_1977,N_1966);
nor U2011 (N_2011,N_1949,N_1920);
and U2012 (N_2012,N_1941,N_1924);
xor U2013 (N_2013,N_1958,N_1963);
nand U2014 (N_2014,N_1929,N_1923);
and U2015 (N_2015,N_1922,N_1936);
or U2016 (N_2016,N_1931,N_1963);
nor U2017 (N_2017,N_1979,N_1955);
nor U2018 (N_2018,N_1959,N_1962);
or U2019 (N_2019,N_1949,N_1926);
and U2020 (N_2020,N_1973,N_1970);
nor U2021 (N_2021,N_1920,N_1937);
or U2022 (N_2022,N_1945,N_1943);
or U2023 (N_2023,N_1941,N_1935);
and U2024 (N_2024,N_1935,N_1958);
or U2025 (N_2025,N_1961,N_1920);
xor U2026 (N_2026,N_1921,N_1964);
nor U2027 (N_2027,N_1937,N_1941);
and U2028 (N_2028,N_1979,N_1948);
nand U2029 (N_2029,N_1953,N_1956);
xnor U2030 (N_2030,N_1960,N_1976);
and U2031 (N_2031,N_1943,N_1923);
nor U2032 (N_2032,N_1954,N_1929);
nor U2033 (N_2033,N_1931,N_1948);
nand U2034 (N_2034,N_1921,N_1929);
or U2035 (N_2035,N_1957,N_1976);
nor U2036 (N_2036,N_1952,N_1950);
and U2037 (N_2037,N_1921,N_1923);
or U2038 (N_2038,N_1956,N_1923);
or U2039 (N_2039,N_1934,N_1975);
xor U2040 (N_2040,N_1991,N_2014);
and U2041 (N_2041,N_1981,N_1997);
nand U2042 (N_2042,N_2034,N_1982);
and U2043 (N_2043,N_2010,N_1984);
xor U2044 (N_2044,N_2007,N_2033);
nor U2045 (N_2045,N_1980,N_2018);
and U2046 (N_2046,N_2038,N_2026);
nor U2047 (N_2047,N_1989,N_2005);
nand U2048 (N_2048,N_2022,N_1995);
nor U2049 (N_2049,N_2000,N_2012);
and U2050 (N_2050,N_2025,N_2006);
xnor U2051 (N_2051,N_1998,N_2023);
or U2052 (N_2052,N_2016,N_2001);
or U2053 (N_2053,N_2037,N_2011);
nand U2054 (N_2054,N_2024,N_2039);
or U2055 (N_2055,N_1999,N_2015);
nor U2056 (N_2056,N_1983,N_2020);
nand U2057 (N_2057,N_1988,N_2013);
nor U2058 (N_2058,N_1996,N_2017);
nor U2059 (N_2059,N_2030,N_1994);
nand U2060 (N_2060,N_1986,N_2028);
and U2061 (N_2061,N_2035,N_2003);
and U2062 (N_2062,N_2009,N_2031);
xor U2063 (N_2063,N_1987,N_2027);
xor U2064 (N_2064,N_1992,N_2002);
nor U2065 (N_2065,N_1990,N_2036);
xor U2066 (N_2066,N_2008,N_1993);
xor U2067 (N_2067,N_2021,N_2029);
nor U2068 (N_2068,N_2004,N_2019);
nor U2069 (N_2069,N_2032,N_1985);
or U2070 (N_2070,N_2012,N_2025);
and U2071 (N_2071,N_2001,N_1993);
nand U2072 (N_2072,N_2009,N_2015);
and U2073 (N_2073,N_1989,N_1987);
nand U2074 (N_2074,N_2026,N_2000);
xor U2075 (N_2075,N_2020,N_2027);
nor U2076 (N_2076,N_2000,N_2022);
nand U2077 (N_2077,N_1982,N_2038);
or U2078 (N_2078,N_2030,N_2024);
or U2079 (N_2079,N_1990,N_2031);
nand U2080 (N_2080,N_2037,N_2029);
and U2081 (N_2081,N_2022,N_2016);
nor U2082 (N_2082,N_2024,N_2010);
nand U2083 (N_2083,N_2025,N_1999);
or U2084 (N_2084,N_1997,N_2003);
nor U2085 (N_2085,N_2029,N_2005);
and U2086 (N_2086,N_1997,N_2008);
and U2087 (N_2087,N_1988,N_1989);
nand U2088 (N_2088,N_2009,N_2035);
nand U2089 (N_2089,N_1990,N_2012);
xor U2090 (N_2090,N_2005,N_1995);
xnor U2091 (N_2091,N_2001,N_2011);
nor U2092 (N_2092,N_2029,N_2009);
and U2093 (N_2093,N_1987,N_2007);
nand U2094 (N_2094,N_2004,N_2038);
nor U2095 (N_2095,N_1980,N_1999);
nand U2096 (N_2096,N_1987,N_1980);
or U2097 (N_2097,N_1998,N_2003);
nor U2098 (N_2098,N_2028,N_1981);
nand U2099 (N_2099,N_1991,N_2038);
nor U2100 (N_2100,N_2083,N_2055);
nand U2101 (N_2101,N_2053,N_2092);
nor U2102 (N_2102,N_2080,N_2089);
and U2103 (N_2103,N_2078,N_2071);
and U2104 (N_2104,N_2094,N_2043);
and U2105 (N_2105,N_2048,N_2047);
nor U2106 (N_2106,N_2077,N_2065);
xnor U2107 (N_2107,N_2091,N_2067);
or U2108 (N_2108,N_2050,N_2098);
and U2109 (N_2109,N_2052,N_2061);
and U2110 (N_2110,N_2049,N_2044);
or U2111 (N_2111,N_2046,N_2070);
and U2112 (N_2112,N_2074,N_2085);
or U2113 (N_2113,N_2099,N_2097);
xnor U2114 (N_2114,N_2086,N_2090);
nand U2115 (N_2115,N_2054,N_2076);
nor U2116 (N_2116,N_2045,N_2075);
xor U2117 (N_2117,N_2064,N_2068);
and U2118 (N_2118,N_2096,N_2084);
and U2119 (N_2119,N_2069,N_2072);
or U2120 (N_2120,N_2040,N_2079);
or U2121 (N_2121,N_2087,N_2062);
or U2122 (N_2122,N_2088,N_2063);
and U2123 (N_2123,N_2095,N_2042);
or U2124 (N_2124,N_2058,N_2041);
nor U2125 (N_2125,N_2066,N_2073);
and U2126 (N_2126,N_2056,N_2051);
xnor U2127 (N_2127,N_2060,N_2093);
xor U2128 (N_2128,N_2081,N_2082);
nand U2129 (N_2129,N_2059,N_2057);
or U2130 (N_2130,N_2065,N_2046);
or U2131 (N_2131,N_2089,N_2098);
or U2132 (N_2132,N_2050,N_2075);
nand U2133 (N_2133,N_2079,N_2075);
nand U2134 (N_2134,N_2046,N_2081);
xnor U2135 (N_2135,N_2042,N_2040);
nor U2136 (N_2136,N_2065,N_2089);
nor U2137 (N_2137,N_2070,N_2041);
nand U2138 (N_2138,N_2045,N_2099);
nand U2139 (N_2139,N_2058,N_2051);
nor U2140 (N_2140,N_2093,N_2042);
and U2141 (N_2141,N_2068,N_2047);
nor U2142 (N_2142,N_2049,N_2040);
xor U2143 (N_2143,N_2089,N_2084);
xnor U2144 (N_2144,N_2078,N_2055);
and U2145 (N_2145,N_2074,N_2077);
nand U2146 (N_2146,N_2097,N_2062);
nor U2147 (N_2147,N_2086,N_2066);
or U2148 (N_2148,N_2070,N_2074);
and U2149 (N_2149,N_2051,N_2049);
and U2150 (N_2150,N_2079,N_2088);
and U2151 (N_2151,N_2079,N_2052);
nand U2152 (N_2152,N_2085,N_2070);
and U2153 (N_2153,N_2087,N_2048);
nor U2154 (N_2154,N_2067,N_2063);
or U2155 (N_2155,N_2063,N_2066);
nor U2156 (N_2156,N_2089,N_2067);
or U2157 (N_2157,N_2064,N_2084);
nand U2158 (N_2158,N_2087,N_2097);
nand U2159 (N_2159,N_2097,N_2061);
or U2160 (N_2160,N_2148,N_2135);
xor U2161 (N_2161,N_2105,N_2112);
nand U2162 (N_2162,N_2104,N_2110);
or U2163 (N_2163,N_2152,N_2142);
and U2164 (N_2164,N_2114,N_2131);
or U2165 (N_2165,N_2119,N_2113);
or U2166 (N_2166,N_2146,N_2134);
nand U2167 (N_2167,N_2137,N_2138);
nor U2168 (N_2168,N_2120,N_2107);
and U2169 (N_2169,N_2147,N_2151);
xnor U2170 (N_2170,N_2144,N_2106);
xnor U2171 (N_2171,N_2121,N_2141);
nand U2172 (N_2172,N_2133,N_2132);
and U2173 (N_2173,N_2108,N_2154);
nor U2174 (N_2174,N_2101,N_2128);
nor U2175 (N_2175,N_2149,N_2115);
nor U2176 (N_2176,N_2140,N_2118);
or U2177 (N_2177,N_2111,N_2156);
nor U2178 (N_2178,N_2117,N_2100);
or U2179 (N_2179,N_2159,N_2155);
or U2180 (N_2180,N_2123,N_2157);
xnor U2181 (N_2181,N_2153,N_2129);
nand U2182 (N_2182,N_2143,N_2125);
or U2183 (N_2183,N_2130,N_2158);
nor U2184 (N_2184,N_2127,N_2139);
and U2185 (N_2185,N_2124,N_2109);
or U2186 (N_2186,N_2126,N_2103);
and U2187 (N_2187,N_2122,N_2145);
nand U2188 (N_2188,N_2150,N_2116);
or U2189 (N_2189,N_2102,N_2136);
or U2190 (N_2190,N_2136,N_2107);
nor U2191 (N_2191,N_2156,N_2140);
or U2192 (N_2192,N_2112,N_2154);
or U2193 (N_2193,N_2141,N_2115);
nor U2194 (N_2194,N_2128,N_2155);
nor U2195 (N_2195,N_2130,N_2116);
nand U2196 (N_2196,N_2155,N_2142);
nor U2197 (N_2197,N_2104,N_2157);
or U2198 (N_2198,N_2128,N_2135);
xnor U2199 (N_2199,N_2151,N_2119);
nand U2200 (N_2200,N_2151,N_2156);
or U2201 (N_2201,N_2121,N_2131);
xnor U2202 (N_2202,N_2103,N_2122);
xnor U2203 (N_2203,N_2120,N_2100);
nand U2204 (N_2204,N_2149,N_2151);
and U2205 (N_2205,N_2141,N_2117);
xor U2206 (N_2206,N_2120,N_2158);
nand U2207 (N_2207,N_2115,N_2145);
or U2208 (N_2208,N_2108,N_2152);
or U2209 (N_2209,N_2103,N_2108);
and U2210 (N_2210,N_2136,N_2112);
nand U2211 (N_2211,N_2142,N_2107);
nor U2212 (N_2212,N_2120,N_2101);
xor U2213 (N_2213,N_2151,N_2138);
or U2214 (N_2214,N_2138,N_2158);
xnor U2215 (N_2215,N_2142,N_2104);
nand U2216 (N_2216,N_2133,N_2134);
nor U2217 (N_2217,N_2128,N_2151);
and U2218 (N_2218,N_2158,N_2107);
nand U2219 (N_2219,N_2158,N_2127);
xnor U2220 (N_2220,N_2215,N_2197);
and U2221 (N_2221,N_2182,N_2199);
or U2222 (N_2222,N_2168,N_2164);
nand U2223 (N_2223,N_2176,N_2190);
or U2224 (N_2224,N_2178,N_2196);
and U2225 (N_2225,N_2179,N_2167);
nor U2226 (N_2226,N_2188,N_2162);
or U2227 (N_2227,N_2214,N_2213);
xnor U2228 (N_2228,N_2217,N_2206);
nand U2229 (N_2229,N_2191,N_2174);
nor U2230 (N_2230,N_2187,N_2210);
and U2231 (N_2231,N_2181,N_2186);
or U2232 (N_2232,N_2160,N_2192);
or U2233 (N_2233,N_2208,N_2211);
nor U2234 (N_2234,N_2201,N_2202);
xor U2235 (N_2235,N_2180,N_2207);
or U2236 (N_2236,N_2219,N_2198);
or U2237 (N_2237,N_2194,N_2200);
nor U2238 (N_2238,N_2209,N_2173);
and U2239 (N_2239,N_2177,N_2195);
and U2240 (N_2240,N_2204,N_2183);
nand U2241 (N_2241,N_2166,N_2185);
xor U2242 (N_2242,N_2212,N_2218);
and U2243 (N_2243,N_2170,N_2172);
nand U2244 (N_2244,N_2216,N_2189);
xor U2245 (N_2245,N_2161,N_2193);
xnor U2246 (N_2246,N_2184,N_2171);
nor U2247 (N_2247,N_2205,N_2169);
and U2248 (N_2248,N_2203,N_2163);
and U2249 (N_2249,N_2175,N_2165);
nor U2250 (N_2250,N_2207,N_2174);
or U2251 (N_2251,N_2195,N_2168);
nand U2252 (N_2252,N_2163,N_2178);
or U2253 (N_2253,N_2165,N_2168);
or U2254 (N_2254,N_2181,N_2204);
or U2255 (N_2255,N_2172,N_2176);
and U2256 (N_2256,N_2211,N_2206);
nand U2257 (N_2257,N_2193,N_2184);
or U2258 (N_2258,N_2167,N_2160);
nor U2259 (N_2259,N_2204,N_2212);
nand U2260 (N_2260,N_2165,N_2162);
nor U2261 (N_2261,N_2190,N_2162);
nor U2262 (N_2262,N_2168,N_2186);
nand U2263 (N_2263,N_2193,N_2216);
nor U2264 (N_2264,N_2211,N_2191);
nand U2265 (N_2265,N_2172,N_2178);
nand U2266 (N_2266,N_2180,N_2208);
nand U2267 (N_2267,N_2183,N_2164);
nor U2268 (N_2268,N_2184,N_2208);
nor U2269 (N_2269,N_2177,N_2188);
xor U2270 (N_2270,N_2207,N_2167);
nand U2271 (N_2271,N_2200,N_2216);
nor U2272 (N_2272,N_2176,N_2175);
nor U2273 (N_2273,N_2173,N_2188);
nand U2274 (N_2274,N_2180,N_2218);
xnor U2275 (N_2275,N_2194,N_2188);
nor U2276 (N_2276,N_2161,N_2198);
xnor U2277 (N_2277,N_2212,N_2216);
nor U2278 (N_2278,N_2193,N_2214);
nor U2279 (N_2279,N_2199,N_2200);
xor U2280 (N_2280,N_2262,N_2225);
or U2281 (N_2281,N_2229,N_2221);
or U2282 (N_2282,N_2233,N_2259);
nor U2283 (N_2283,N_2232,N_2230);
or U2284 (N_2284,N_2236,N_2245);
nand U2285 (N_2285,N_2263,N_2258);
xnor U2286 (N_2286,N_2265,N_2249);
or U2287 (N_2287,N_2275,N_2248);
xnor U2288 (N_2288,N_2240,N_2279);
nor U2289 (N_2289,N_2252,N_2244);
and U2290 (N_2290,N_2256,N_2276);
or U2291 (N_2291,N_2273,N_2250);
xor U2292 (N_2292,N_2220,N_2264);
xnor U2293 (N_2293,N_2274,N_2271);
nand U2294 (N_2294,N_2228,N_2231);
nor U2295 (N_2295,N_2246,N_2239);
or U2296 (N_2296,N_2255,N_2268);
nand U2297 (N_2297,N_2237,N_2261);
or U2298 (N_2298,N_2267,N_2223);
xnor U2299 (N_2299,N_2253,N_2247);
or U2300 (N_2300,N_2257,N_2238);
nor U2301 (N_2301,N_2272,N_2243);
xnor U2302 (N_2302,N_2266,N_2222);
nor U2303 (N_2303,N_2241,N_2269);
nand U2304 (N_2304,N_2277,N_2251);
xor U2305 (N_2305,N_2224,N_2278);
nor U2306 (N_2306,N_2226,N_2227);
or U2307 (N_2307,N_2235,N_2254);
and U2308 (N_2308,N_2270,N_2260);
nand U2309 (N_2309,N_2234,N_2242);
nand U2310 (N_2310,N_2265,N_2279);
or U2311 (N_2311,N_2258,N_2271);
or U2312 (N_2312,N_2222,N_2271);
nand U2313 (N_2313,N_2229,N_2259);
and U2314 (N_2314,N_2267,N_2235);
nand U2315 (N_2315,N_2262,N_2265);
xor U2316 (N_2316,N_2242,N_2226);
or U2317 (N_2317,N_2264,N_2245);
and U2318 (N_2318,N_2229,N_2252);
or U2319 (N_2319,N_2228,N_2221);
or U2320 (N_2320,N_2220,N_2246);
nand U2321 (N_2321,N_2238,N_2250);
nor U2322 (N_2322,N_2254,N_2239);
nor U2323 (N_2323,N_2268,N_2266);
xor U2324 (N_2324,N_2258,N_2275);
nor U2325 (N_2325,N_2245,N_2228);
nor U2326 (N_2326,N_2225,N_2224);
or U2327 (N_2327,N_2241,N_2233);
or U2328 (N_2328,N_2269,N_2270);
and U2329 (N_2329,N_2275,N_2242);
and U2330 (N_2330,N_2266,N_2257);
xnor U2331 (N_2331,N_2242,N_2266);
and U2332 (N_2332,N_2273,N_2233);
xnor U2333 (N_2333,N_2251,N_2241);
xor U2334 (N_2334,N_2247,N_2254);
xnor U2335 (N_2335,N_2262,N_2242);
nor U2336 (N_2336,N_2262,N_2248);
nor U2337 (N_2337,N_2252,N_2273);
nand U2338 (N_2338,N_2259,N_2249);
or U2339 (N_2339,N_2258,N_2233);
nand U2340 (N_2340,N_2338,N_2301);
nor U2341 (N_2341,N_2295,N_2317);
nor U2342 (N_2342,N_2291,N_2282);
xor U2343 (N_2343,N_2334,N_2314);
nor U2344 (N_2344,N_2300,N_2287);
xnor U2345 (N_2345,N_2330,N_2335);
nand U2346 (N_2346,N_2288,N_2310);
xnor U2347 (N_2347,N_2322,N_2307);
and U2348 (N_2348,N_2297,N_2308);
or U2349 (N_2349,N_2284,N_2309);
xor U2350 (N_2350,N_2304,N_2323);
and U2351 (N_2351,N_2281,N_2305);
or U2352 (N_2352,N_2303,N_2327);
xor U2353 (N_2353,N_2312,N_2336);
and U2354 (N_2354,N_2299,N_2293);
nor U2355 (N_2355,N_2331,N_2339);
nor U2356 (N_2356,N_2329,N_2326);
xor U2357 (N_2357,N_2290,N_2328);
or U2358 (N_2358,N_2306,N_2313);
nor U2359 (N_2359,N_2296,N_2321);
nand U2360 (N_2360,N_2337,N_2318);
or U2361 (N_2361,N_2302,N_2298);
or U2362 (N_2362,N_2324,N_2289);
nand U2363 (N_2363,N_2283,N_2333);
and U2364 (N_2364,N_2285,N_2325);
xnor U2365 (N_2365,N_2332,N_2315);
or U2366 (N_2366,N_2292,N_2320);
or U2367 (N_2367,N_2311,N_2294);
and U2368 (N_2368,N_2280,N_2319);
nand U2369 (N_2369,N_2286,N_2316);
and U2370 (N_2370,N_2335,N_2319);
nand U2371 (N_2371,N_2317,N_2305);
or U2372 (N_2372,N_2324,N_2301);
nor U2373 (N_2373,N_2329,N_2310);
nand U2374 (N_2374,N_2327,N_2329);
and U2375 (N_2375,N_2297,N_2327);
or U2376 (N_2376,N_2327,N_2331);
and U2377 (N_2377,N_2324,N_2310);
nor U2378 (N_2378,N_2297,N_2328);
xor U2379 (N_2379,N_2333,N_2298);
and U2380 (N_2380,N_2287,N_2283);
nand U2381 (N_2381,N_2299,N_2337);
nand U2382 (N_2382,N_2335,N_2299);
nor U2383 (N_2383,N_2283,N_2317);
or U2384 (N_2384,N_2286,N_2289);
nand U2385 (N_2385,N_2309,N_2297);
nand U2386 (N_2386,N_2287,N_2321);
nand U2387 (N_2387,N_2291,N_2327);
nor U2388 (N_2388,N_2300,N_2305);
nand U2389 (N_2389,N_2314,N_2339);
xnor U2390 (N_2390,N_2326,N_2298);
nand U2391 (N_2391,N_2324,N_2311);
or U2392 (N_2392,N_2282,N_2281);
or U2393 (N_2393,N_2306,N_2323);
nand U2394 (N_2394,N_2322,N_2306);
nor U2395 (N_2395,N_2317,N_2314);
xor U2396 (N_2396,N_2285,N_2336);
or U2397 (N_2397,N_2300,N_2331);
or U2398 (N_2398,N_2312,N_2331);
and U2399 (N_2399,N_2301,N_2334);
nand U2400 (N_2400,N_2367,N_2399);
nand U2401 (N_2401,N_2374,N_2382);
nand U2402 (N_2402,N_2363,N_2356);
nor U2403 (N_2403,N_2381,N_2359);
nand U2404 (N_2404,N_2375,N_2358);
nand U2405 (N_2405,N_2391,N_2373);
nand U2406 (N_2406,N_2378,N_2379);
nand U2407 (N_2407,N_2355,N_2365);
xor U2408 (N_2408,N_2353,N_2361);
or U2409 (N_2409,N_2341,N_2390);
nor U2410 (N_2410,N_2397,N_2396);
nor U2411 (N_2411,N_2393,N_2394);
or U2412 (N_2412,N_2350,N_2366);
nor U2413 (N_2413,N_2342,N_2398);
nor U2414 (N_2414,N_2369,N_2352);
or U2415 (N_2415,N_2380,N_2357);
and U2416 (N_2416,N_2368,N_2371);
and U2417 (N_2417,N_2387,N_2388);
and U2418 (N_2418,N_2351,N_2376);
nand U2419 (N_2419,N_2362,N_2354);
and U2420 (N_2420,N_2395,N_2346);
nand U2421 (N_2421,N_2348,N_2385);
nand U2422 (N_2422,N_2360,N_2343);
nand U2423 (N_2423,N_2349,N_2392);
xnor U2424 (N_2424,N_2383,N_2372);
xor U2425 (N_2425,N_2386,N_2389);
or U2426 (N_2426,N_2345,N_2370);
xor U2427 (N_2427,N_2377,N_2344);
or U2428 (N_2428,N_2384,N_2364);
or U2429 (N_2429,N_2340,N_2347);
nand U2430 (N_2430,N_2363,N_2365);
and U2431 (N_2431,N_2377,N_2343);
xnor U2432 (N_2432,N_2369,N_2390);
and U2433 (N_2433,N_2358,N_2394);
nor U2434 (N_2434,N_2376,N_2388);
and U2435 (N_2435,N_2374,N_2395);
nand U2436 (N_2436,N_2347,N_2397);
xnor U2437 (N_2437,N_2368,N_2352);
nor U2438 (N_2438,N_2395,N_2392);
xor U2439 (N_2439,N_2392,N_2393);
nor U2440 (N_2440,N_2376,N_2385);
and U2441 (N_2441,N_2357,N_2343);
nor U2442 (N_2442,N_2392,N_2399);
nand U2443 (N_2443,N_2391,N_2378);
and U2444 (N_2444,N_2354,N_2398);
xnor U2445 (N_2445,N_2397,N_2391);
nor U2446 (N_2446,N_2369,N_2398);
nor U2447 (N_2447,N_2385,N_2379);
or U2448 (N_2448,N_2361,N_2394);
and U2449 (N_2449,N_2396,N_2388);
nor U2450 (N_2450,N_2397,N_2357);
or U2451 (N_2451,N_2361,N_2381);
nand U2452 (N_2452,N_2391,N_2341);
or U2453 (N_2453,N_2343,N_2347);
nand U2454 (N_2454,N_2382,N_2352);
nand U2455 (N_2455,N_2353,N_2398);
or U2456 (N_2456,N_2392,N_2390);
nand U2457 (N_2457,N_2394,N_2351);
nand U2458 (N_2458,N_2340,N_2360);
nand U2459 (N_2459,N_2389,N_2399);
nor U2460 (N_2460,N_2443,N_2428);
xnor U2461 (N_2461,N_2450,N_2424);
xor U2462 (N_2462,N_2452,N_2455);
nor U2463 (N_2463,N_2416,N_2437);
nand U2464 (N_2464,N_2447,N_2411);
nand U2465 (N_2465,N_2453,N_2404);
nand U2466 (N_2466,N_2448,N_2426);
or U2467 (N_2467,N_2435,N_2413);
nor U2468 (N_2468,N_2421,N_2442);
or U2469 (N_2469,N_2436,N_2439);
nand U2470 (N_2470,N_2418,N_2415);
and U2471 (N_2471,N_2427,N_2451);
or U2472 (N_2472,N_2456,N_2440);
xnor U2473 (N_2473,N_2449,N_2405);
and U2474 (N_2474,N_2441,N_2429);
nand U2475 (N_2475,N_2432,N_2407);
and U2476 (N_2476,N_2412,N_2400);
and U2477 (N_2477,N_2457,N_2408);
xnor U2478 (N_2478,N_2420,N_2430);
nor U2479 (N_2479,N_2419,N_2446);
nor U2480 (N_2480,N_2403,N_2459);
xnor U2481 (N_2481,N_2444,N_2433);
and U2482 (N_2482,N_2410,N_2409);
xor U2483 (N_2483,N_2402,N_2431);
and U2484 (N_2484,N_2406,N_2417);
nor U2485 (N_2485,N_2414,N_2434);
or U2486 (N_2486,N_2454,N_2422);
nand U2487 (N_2487,N_2401,N_2438);
and U2488 (N_2488,N_2423,N_2425);
nor U2489 (N_2489,N_2458,N_2445);
and U2490 (N_2490,N_2448,N_2449);
or U2491 (N_2491,N_2432,N_2403);
nand U2492 (N_2492,N_2445,N_2450);
nor U2493 (N_2493,N_2430,N_2449);
nor U2494 (N_2494,N_2452,N_2446);
nor U2495 (N_2495,N_2415,N_2405);
nor U2496 (N_2496,N_2440,N_2436);
and U2497 (N_2497,N_2407,N_2416);
or U2498 (N_2498,N_2426,N_2434);
and U2499 (N_2499,N_2408,N_2456);
and U2500 (N_2500,N_2431,N_2405);
nor U2501 (N_2501,N_2411,N_2440);
xnor U2502 (N_2502,N_2456,N_2420);
xor U2503 (N_2503,N_2448,N_2441);
nor U2504 (N_2504,N_2412,N_2451);
xnor U2505 (N_2505,N_2414,N_2437);
nand U2506 (N_2506,N_2438,N_2449);
and U2507 (N_2507,N_2444,N_2404);
and U2508 (N_2508,N_2427,N_2405);
and U2509 (N_2509,N_2403,N_2423);
nand U2510 (N_2510,N_2443,N_2440);
and U2511 (N_2511,N_2440,N_2417);
nor U2512 (N_2512,N_2445,N_2443);
or U2513 (N_2513,N_2402,N_2413);
or U2514 (N_2514,N_2400,N_2417);
nand U2515 (N_2515,N_2420,N_2411);
nand U2516 (N_2516,N_2410,N_2448);
and U2517 (N_2517,N_2449,N_2444);
nand U2518 (N_2518,N_2400,N_2421);
nor U2519 (N_2519,N_2436,N_2450);
and U2520 (N_2520,N_2481,N_2510);
or U2521 (N_2521,N_2469,N_2504);
nand U2522 (N_2522,N_2482,N_2498);
nor U2523 (N_2523,N_2484,N_2506);
and U2524 (N_2524,N_2509,N_2463);
xor U2525 (N_2525,N_2477,N_2465);
or U2526 (N_2526,N_2467,N_2483);
nand U2527 (N_2527,N_2472,N_2495);
xor U2528 (N_2528,N_2489,N_2488);
nor U2529 (N_2529,N_2513,N_2496);
or U2530 (N_2530,N_2479,N_2497);
nand U2531 (N_2531,N_2475,N_2515);
xor U2532 (N_2532,N_2501,N_2508);
or U2533 (N_2533,N_2461,N_2468);
xnor U2534 (N_2534,N_2503,N_2516);
and U2535 (N_2535,N_2462,N_2490);
and U2536 (N_2536,N_2499,N_2466);
nor U2537 (N_2537,N_2517,N_2518);
xnor U2538 (N_2538,N_2493,N_2485);
and U2539 (N_2539,N_2480,N_2478);
or U2540 (N_2540,N_2507,N_2514);
xnor U2541 (N_2541,N_2492,N_2464);
xnor U2542 (N_2542,N_2505,N_2487);
nor U2543 (N_2543,N_2519,N_2474);
or U2544 (N_2544,N_2473,N_2460);
or U2545 (N_2545,N_2512,N_2502);
xnor U2546 (N_2546,N_2500,N_2471);
or U2547 (N_2547,N_2470,N_2486);
nand U2548 (N_2548,N_2511,N_2491);
and U2549 (N_2549,N_2476,N_2494);
and U2550 (N_2550,N_2469,N_2484);
xnor U2551 (N_2551,N_2509,N_2468);
nor U2552 (N_2552,N_2514,N_2494);
nor U2553 (N_2553,N_2494,N_2496);
xnor U2554 (N_2554,N_2513,N_2460);
and U2555 (N_2555,N_2478,N_2496);
and U2556 (N_2556,N_2506,N_2508);
or U2557 (N_2557,N_2498,N_2474);
nor U2558 (N_2558,N_2501,N_2494);
or U2559 (N_2559,N_2503,N_2462);
or U2560 (N_2560,N_2501,N_2519);
nor U2561 (N_2561,N_2493,N_2469);
xnor U2562 (N_2562,N_2514,N_2511);
or U2563 (N_2563,N_2492,N_2493);
xnor U2564 (N_2564,N_2515,N_2517);
nand U2565 (N_2565,N_2509,N_2508);
nand U2566 (N_2566,N_2481,N_2507);
nor U2567 (N_2567,N_2510,N_2507);
xnor U2568 (N_2568,N_2516,N_2487);
xnor U2569 (N_2569,N_2519,N_2516);
or U2570 (N_2570,N_2478,N_2490);
nor U2571 (N_2571,N_2513,N_2502);
nand U2572 (N_2572,N_2488,N_2463);
nand U2573 (N_2573,N_2473,N_2462);
and U2574 (N_2574,N_2484,N_2461);
xor U2575 (N_2575,N_2468,N_2517);
nor U2576 (N_2576,N_2466,N_2511);
or U2577 (N_2577,N_2471,N_2478);
and U2578 (N_2578,N_2502,N_2468);
nor U2579 (N_2579,N_2494,N_2497);
or U2580 (N_2580,N_2566,N_2559);
nand U2581 (N_2581,N_2525,N_2563);
xnor U2582 (N_2582,N_2560,N_2557);
and U2583 (N_2583,N_2533,N_2529);
nor U2584 (N_2584,N_2541,N_2542);
nand U2585 (N_2585,N_2555,N_2554);
nor U2586 (N_2586,N_2552,N_2538);
and U2587 (N_2587,N_2547,N_2548);
xor U2588 (N_2588,N_2532,N_2569);
or U2589 (N_2589,N_2536,N_2537);
xnor U2590 (N_2590,N_2568,N_2531);
nand U2591 (N_2591,N_2553,N_2523);
nor U2592 (N_2592,N_2575,N_2579);
or U2593 (N_2593,N_2540,N_2522);
and U2594 (N_2594,N_2545,N_2539);
xor U2595 (N_2595,N_2573,N_2527);
or U2596 (N_2596,N_2546,N_2530);
xor U2597 (N_2597,N_2558,N_2526);
xnor U2598 (N_2598,N_2577,N_2556);
or U2599 (N_2599,N_2544,N_2571);
and U2600 (N_2600,N_2524,N_2561);
or U2601 (N_2601,N_2549,N_2578);
and U2602 (N_2602,N_2534,N_2551);
or U2603 (N_2603,N_2520,N_2564);
nand U2604 (N_2604,N_2565,N_2562);
xnor U2605 (N_2605,N_2572,N_2528);
xor U2606 (N_2606,N_2574,N_2535);
or U2607 (N_2607,N_2567,N_2543);
or U2608 (N_2608,N_2521,N_2570);
nor U2609 (N_2609,N_2550,N_2576);
nand U2610 (N_2610,N_2556,N_2521);
or U2611 (N_2611,N_2542,N_2526);
and U2612 (N_2612,N_2536,N_2552);
and U2613 (N_2613,N_2523,N_2538);
xor U2614 (N_2614,N_2538,N_2528);
xnor U2615 (N_2615,N_2528,N_2579);
nor U2616 (N_2616,N_2547,N_2571);
and U2617 (N_2617,N_2543,N_2527);
xor U2618 (N_2618,N_2546,N_2544);
or U2619 (N_2619,N_2540,N_2555);
nand U2620 (N_2620,N_2538,N_2567);
xor U2621 (N_2621,N_2553,N_2538);
and U2622 (N_2622,N_2529,N_2574);
or U2623 (N_2623,N_2556,N_2558);
nor U2624 (N_2624,N_2577,N_2567);
and U2625 (N_2625,N_2533,N_2527);
xor U2626 (N_2626,N_2568,N_2544);
or U2627 (N_2627,N_2540,N_2543);
or U2628 (N_2628,N_2557,N_2525);
nor U2629 (N_2629,N_2542,N_2566);
xor U2630 (N_2630,N_2575,N_2545);
nand U2631 (N_2631,N_2560,N_2555);
and U2632 (N_2632,N_2560,N_2563);
and U2633 (N_2633,N_2551,N_2544);
or U2634 (N_2634,N_2568,N_2574);
or U2635 (N_2635,N_2564,N_2533);
nand U2636 (N_2636,N_2521,N_2548);
or U2637 (N_2637,N_2574,N_2577);
or U2638 (N_2638,N_2535,N_2562);
nand U2639 (N_2639,N_2569,N_2523);
xnor U2640 (N_2640,N_2584,N_2589);
nor U2641 (N_2641,N_2592,N_2605);
xor U2642 (N_2642,N_2585,N_2613);
xor U2643 (N_2643,N_2639,N_2630);
or U2644 (N_2644,N_2594,N_2618);
nand U2645 (N_2645,N_2590,N_2595);
xor U2646 (N_2646,N_2601,N_2608);
nor U2647 (N_2647,N_2596,N_2612);
nor U2648 (N_2648,N_2616,N_2623);
nor U2649 (N_2649,N_2600,N_2634);
or U2650 (N_2650,N_2598,N_2617);
xnor U2651 (N_2651,N_2636,N_2614);
xnor U2652 (N_2652,N_2620,N_2581);
xnor U2653 (N_2653,N_2619,N_2624);
and U2654 (N_2654,N_2631,N_2615);
xor U2655 (N_2655,N_2604,N_2583);
and U2656 (N_2656,N_2627,N_2588);
and U2657 (N_2657,N_2603,N_2606);
and U2658 (N_2658,N_2621,N_2628);
nor U2659 (N_2659,N_2611,N_2602);
and U2660 (N_2660,N_2638,N_2580);
nor U2661 (N_2661,N_2626,N_2587);
xor U2662 (N_2662,N_2633,N_2609);
and U2663 (N_2663,N_2625,N_2629);
xnor U2664 (N_2664,N_2622,N_2635);
xor U2665 (N_2665,N_2582,N_2632);
nand U2666 (N_2666,N_2586,N_2607);
nor U2667 (N_2667,N_2610,N_2637);
nor U2668 (N_2668,N_2599,N_2591);
or U2669 (N_2669,N_2597,N_2593);
or U2670 (N_2670,N_2616,N_2614);
nand U2671 (N_2671,N_2583,N_2607);
nor U2672 (N_2672,N_2589,N_2614);
or U2673 (N_2673,N_2584,N_2624);
or U2674 (N_2674,N_2594,N_2584);
and U2675 (N_2675,N_2596,N_2582);
nand U2676 (N_2676,N_2588,N_2611);
and U2677 (N_2677,N_2588,N_2616);
nand U2678 (N_2678,N_2621,N_2588);
or U2679 (N_2679,N_2580,N_2626);
nor U2680 (N_2680,N_2603,N_2635);
nand U2681 (N_2681,N_2620,N_2587);
or U2682 (N_2682,N_2599,N_2597);
and U2683 (N_2683,N_2593,N_2614);
and U2684 (N_2684,N_2611,N_2634);
nor U2685 (N_2685,N_2635,N_2601);
and U2686 (N_2686,N_2607,N_2581);
and U2687 (N_2687,N_2599,N_2587);
nor U2688 (N_2688,N_2600,N_2616);
or U2689 (N_2689,N_2618,N_2589);
and U2690 (N_2690,N_2602,N_2598);
xnor U2691 (N_2691,N_2591,N_2632);
and U2692 (N_2692,N_2633,N_2626);
nand U2693 (N_2693,N_2636,N_2595);
nand U2694 (N_2694,N_2639,N_2580);
nand U2695 (N_2695,N_2588,N_2636);
and U2696 (N_2696,N_2612,N_2602);
nor U2697 (N_2697,N_2580,N_2602);
nor U2698 (N_2698,N_2588,N_2624);
or U2699 (N_2699,N_2629,N_2612);
xnor U2700 (N_2700,N_2662,N_2684);
nand U2701 (N_2701,N_2673,N_2659);
or U2702 (N_2702,N_2680,N_2652);
xnor U2703 (N_2703,N_2648,N_2690);
xnor U2704 (N_2704,N_2663,N_2694);
xnor U2705 (N_2705,N_2645,N_2679);
or U2706 (N_2706,N_2675,N_2671);
xnor U2707 (N_2707,N_2693,N_2678);
xnor U2708 (N_2708,N_2649,N_2661);
xor U2709 (N_2709,N_2651,N_2676);
nor U2710 (N_2710,N_2646,N_2665);
or U2711 (N_2711,N_2643,N_2685);
xor U2712 (N_2712,N_2667,N_2656);
or U2713 (N_2713,N_2647,N_2689);
and U2714 (N_2714,N_2660,N_2695);
nand U2715 (N_2715,N_2640,N_2674);
and U2716 (N_2716,N_2697,N_2669);
nand U2717 (N_2717,N_2654,N_2677);
or U2718 (N_2718,N_2687,N_2691);
nand U2719 (N_2719,N_2655,N_2683);
xnor U2720 (N_2720,N_2642,N_2657);
and U2721 (N_2721,N_2650,N_2644);
xnor U2722 (N_2722,N_2672,N_2681);
or U2723 (N_2723,N_2653,N_2699);
nand U2724 (N_2724,N_2668,N_2682);
nand U2725 (N_2725,N_2658,N_2698);
nor U2726 (N_2726,N_2686,N_2696);
nor U2727 (N_2727,N_2670,N_2664);
nor U2728 (N_2728,N_2641,N_2692);
nand U2729 (N_2729,N_2688,N_2666);
and U2730 (N_2730,N_2695,N_2661);
and U2731 (N_2731,N_2694,N_2673);
or U2732 (N_2732,N_2695,N_2680);
or U2733 (N_2733,N_2653,N_2660);
xnor U2734 (N_2734,N_2641,N_2678);
nand U2735 (N_2735,N_2662,N_2698);
xnor U2736 (N_2736,N_2647,N_2697);
and U2737 (N_2737,N_2660,N_2699);
xnor U2738 (N_2738,N_2680,N_2681);
xor U2739 (N_2739,N_2672,N_2693);
nand U2740 (N_2740,N_2692,N_2670);
nor U2741 (N_2741,N_2667,N_2669);
and U2742 (N_2742,N_2652,N_2693);
nand U2743 (N_2743,N_2643,N_2647);
nand U2744 (N_2744,N_2678,N_2696);
nand U2745 (N_2745,N_2680,N_2679);
nor U2746 (N_2746,N_2663,N_2649);
xor U2747 (N_2747,N_2680,N_2669);
or U2748 (N_2748,N_2680,N_2661);
or U2749 (N_2749,N_2674,N_2660);
or U2750 (N_2750,N_2647,N_2652);
xor U2751 (N_2751,N_2670,N_2660);
nand U2752 (N_2752,N_2642,N_2655);
nor U2753 (N_2753,N_2657,N_2658);
or U2754 (N_2754,N_2675,N_2697);
nor U2755 (N_2755,N_2645,N_2693);
nor U2756 (N_2756,N_2667,N_2642);
xor U2757 (N_2757,N_2668,N_2647);
xor U2758 (N_2758,N_2642,N_2689);
nor U2759 (N_2759,N_2668,N_2656);
xor U2760 (N_2760,N_2750,N_2743);
nand U2761 (N_2761,N_2731,N_2720);
nand U2762 (N_2762,N_2709,N_2757);
and U2763 (N_2763,N_2718,N_2732);
nand U2764 (N_2764,N_2746,N_2725);
xnor U2765 (N_2765,N_2704,N_2728);
and U2766 (N_2766,N_2724,N_2702);
or U2767 (N_2767,N_2715,N_2745);
and U2768 (N_2768,N_2753,N_2736);
nor U2769 (N_2769,N_2716,N_2735);
or U2770 (N_2770,N_2711,N_2713);
and U2771 (N_2771,N_2710,N_2708);
xor U2772 (N_2772,N_2754,N_2707);
and U2773 (N_2773,N_2712,N_2717);
or U2774 (N_2774,N_2749,N_2756);
xnor U2775 (N_2775,N_2734,N_2747);
nor U2776 (N_2776,N_2714,N_2723);
xnor U2777 (N_2777,N_2726,N_2706);
or U2778 (N_2778,N_2744,N_2759);
and U2779 (N_2779,N_2727,N_2701);
and U2780 (N_2780,N_2752,N_2721);
or U2781 (N_2781,N_2700,N_2741);
and U2782 (N_2782,N_2705,N_2733);
or U2783 (N_2783,N_2737,N_2742);
nor U2784 (N_2784,N_2719,N_2730);
nand U2785 (N_2785,N_2758,N_2748);
and U2786 (N_2786,N_2755,N_2739);
or U2787 (N_2787,N_2722,N_2738);
or U2788 (N_2788,N_2751,N_2729);
xnor U2789 (N_2789,N_2740,N_2703);
nor U2790 (N_2790,N_2746,N_2733);
xor U2791 (N_2791,N_2744,N_2700);
and U2792 (N_2792,N_2740,N_2748);
xor U2793 (N_2793,N_2706,N_2719);
or U2794 (N_2794,N_2736,N_2722);
nand U2795 (N_2795,N_2743,N_2723);
nand U2796 (N_2796,N_2718,N_2715);
and U2797 (N_2797,N_2720,N_2738);
and U2798 (N_2798,N_2744,N_2708);
and U2799 (N_2799,N_2723,N_2728);
and U2800 (N_2800,N_2719,N_2701);
and U2801 (N_2801,N_2754,N_2744);
or U2802 (N_2802,N_2713,N_2707);
nor U2803 (N_2803,N_2734,N_2737);
xnor U2804 (N_2804,N_2738,N_2713);
and U2805 (N_2805,N_2759,N_2717);
nand U2806 (N_2806,N_2717,N_2721);
or U2807 (N_2807,N_2755,N_2716);
nand U2808 (N_2808,N_2746,N_2706);
and U2809 (N_2809,N_2726,N_2704);
and U2810 (N_2810,N_2725,N_2743);
or U2811 (N_2811,N_2742,N_2713);
or U2812 (N_2812,N_2750,N_2715);
xnor U2813 (N_2813,N_2735,N_2737);
and U2814 (N_2814,N_2735,N_2723);
nor U2815 (N_2815,N_2732,N_2715);
nand U2816 (N_2816,N_2724,N_2753);
xor U2817 (N_2817,N_2715,N_2754);
and U2818 (N_2818,N_2737,N_2729);
nor U2819 (N_2819,N_2722,N_2741);
and U2820 (N_2820,N_2795,N_2789);
or U2821 (N_2821,N_2819,N_2772);
and U2822 (N_2822,N_2764,N_2776);
nor U2823 (N_2823,N_2790,N_2817);
nand U2824 (N_2824,N_2779,N_2783);
nand U2825 (N_2825,N_2800,N_2811);
xnor U2826 (N_2826,N_2786,N_2807);
nor U2827 (N_2827,N_2814,N_2797);
nor U2828 (N_2828,N_2768,N_2815);
xor U2829 (N_2829,N_2784,N_2810);
nor U2830 (N_2830,N_2796,N_2793);
or U2831 (N_2831,N_2782,N_2778);
xnor U2832 (N_2832,N_2762,N_2812);
xor U2833 (N_2833,N_2794,N_2801);
nand U2834 (N_2834,N_2798,N_2774);
nand U2835 (N_2835,N_2799,N_2760);
or U2836 (N_2836,N_2771,N_2769);
or U2837 (N_2837,N_2802,N_2765);
xnor U2838 (N_2838,N_2767,N_2818);
and U2839 (N_2839,N_2770,N_2816);
and U2840 (N_2840,N_2777,N_2808);
or U2841 (N_2841,N_2803,N_2809);
or U2842 (N_2842,N_2761,N_2773);
and U2843 (N_2843,N_2763,N_2806);
xnor U2844 (N_2844,N_2780,N_2804);
nand U2845 (N_2845,N_2787,N_2791);
nor U2846 (N_2846,N_2813,N_2766);
and U2847 (N_2847,N_2775,N_2792);
nor U2848 (N_2848,N_2805,N_2785);
or U2849 (N_2849,N_2788,N_2781);
or U2850 (N_2850,N_2793,N_2784);
nor U2851 (N_2851,N_2795,N_2761);
or U2852 (N_2852,N_2810,N_2797);
nand U2853 (N_2853,N_2791,N_2767);
nand U2854 (N_2854,N_2789,N_2777);
nor U2855 (N_2855,N_2786,N_2813);
and U2856 (N_2856,N_2786,N_2780);
xor U2857 (N_2857,N_2771,N_2787);
xnor U2858 (N_2858,N_2805,N_2812);
and U2859 (N_2859,N_2793,N_2809);
nor U2860 (N_2860,N_2786,N_2806);
and U2861 (N_2861,N_2788,N_2767);
or U2862 (N_2862,N_2784,N_2773);
or U2863 (N_2863,N_2814,N_2765);
xor U2864 (N_2864,N_2801,N_2784);
xor U2865 (N_2865,N_2785,N_2777);
and U2866 (N_2866,N_2782,N_2779);
nor U2867 (N_2867,N_2765,N_2788);
or U2868 (N_2868,N_2814,N_2794);
and U2869 (N_2869,N_2819,N_2765);
nor U2870 (N_2870,N_2799,N_2803);
xor U2871 (N_2871,N_2795,N_2781);
and U2872 (N_2872,N_2766,N_2764);
and U2873 (N_2873,N_2815,N_2787);
and U2874 (N_2874,N_2818,N_2789);
or U2875 (N_2875,N_2764,N_2800);
and U2876 (N_2876,N_2781,N_2780);
and U2877 (N_2877,N_2785,N_2791);
nor U2878 (N_2878,N_2773,N_2777);
nand U2879 (N_2879,N_2815,N_2809);
nor U2880 (N_2880,N_2827,N_2822);
or U2881 (N_2881,N_2866,N_2835);
xor U2882 (N_2882,N_2869,N_2834);
nand U2883 (N_2883,N_2851,N_2837);
nand U2884 (N_2884,N_2870,N_2845);
nor U2885 (N_2885,N_2873,N_2833);
or U2886 (N_2886,N_2828,N_2841);
or U2887 (N_2887,N_2847,N_2856);
xnor U2888 (N_2888,N_2854,N_2857);
or U2889 (N_2889,N_2860,N_2824);
and U2890 (N_2890,N_2864,N_2871);
nor U2891 (N_2891,N_2836,N_2862);
nand U2892 (N_2892,N_2820,N_2829);
nand U2893 (N_2893,N_2861,N_2843);
or U2894 (N_2894,N_2838,N_2872);
nand U2895 (N_2895,N_2842,N_2863);
xnor U2896 (N_2896,N_2853,N_2823);
nand U2897 (N_2897,N_2865,N_2849);
or U2898 (N_2898,N_2876,N_2840);
and U2899 (N_2899,N_2858,N_2850);
and U2900 (N_2900,N_2826,N_2832);
and U2901 (N_2901,N_2825,N_2830);
or U2902 (N_2902,N_2868,N_2879);
nor U2903 (N_2903,N_2821,N_2867);
nor U2904 (N_2904,N_2875,N_2855);
or U2905 (N_2905,N_2877,N_2878);
nor U2906 (N_2906,N_2859,N_2852);
nor U2907 (N_2907,N_2831,N_2846);
and U2908 (N_2908,N_2839,N_2844);
xor U2909 (N_2909,N_2848,N_2874);
and U2910 (N_2910,N_2844,N_2879);
or U2911 (N_2911,N_2878,N_2857);
xor U2912 (N_2912,N_2874,N_2878);
nor U2913 (N_2913,N_2825,N_2836);
and U2914 (N_2914,N_2875,N_2858);
nand U2915 (N_2915,N_2845,N_2839);
nor U2916 (N_2916,N_2867,N_2859);
xnor U2917 (N_2917,N_2852,N_2876);
or U2918 (N_2918,N_2875,N_2870);
nand U2919 (N_2919,N_2857,N_2862);
nand U2920 (N_2920,N_2854,N_2860);
or U2921 (N_2921,N_2855,N_2837);
nand U2922 (N_2922,N_2834,N_2847);
nand U2923 (N_2923,N_2872,N_2835);
nand U2924 (N_2924,N_2839,N_2830);
nor U2925 (N_2925,N_2855,N_2822);
nor U2926 (N_2926,N_2848,N_2855);
and U2927 (N_2927,N_2833,N_2875);
and U2928 (N_2928,N_2820,N_2864);
or U2929 (N_2929,N_2862,N_2867);
nor U2930 (N_2930,N_2870,N_2820);
or U2931 (N_2931,N_2846,N_2858);
xor U2932 (N_2932,N_2850,N_2860);
nor U2933 (N_2933,N_2833,N_2824);
and U2934 (N_2934,N_2828,N_2821);
xor U2935 (N_2935,N_2832,N_2852);
xor U2936 (N_2936,N_2853,N_2878);
and U2937 (N_2937,N_2866,N_2847);
nor U2938 (N_2938,N_2839,N_2857);
xor U2939 (N_2939,N_2820,N_2823);
nand U2940 (N_2940,N_2880,N_2938);
or U2941 (N_2941,N_2920,N_2928);
xor U2942 (N_2942,N_2898,N_2939);
nor U2943 (N_2943,N_2893,N_2884);
nand U2944 (N_2944,N_2929,N_2885);
xnor U2945 (N_2945,N_2933,N_2913);
or U2946 (N_2946,N_2908,N_2905);
nand U2947 (N_2947,N_2889,N_2922);
and U2948 (N_2948,N_2912,N_2917);
nor U2949 (N_2949,N_2886,N_2881);
and U2950 (N_2950,N_2918,N_2909);
xor U2951 (N_2951,N_2931,N_2923);
xnor U2952 (N_2952,N_2924,N_2911);
nand U2953 (N_2953,N_2934,N_2899);
nand U2954 (N_2954,N_2891,N_2914);
nor U2955 (N_2955,N_2883,N_2892);
nand U2956 (N_2956,N_2907,N_2921);
xor U2957 (N_2957,N_2925,N_2937);
or U2958 (N_2958,N_2890,N_2910);
nand U2959 (N_2959,N_2903,N_2935);
xnor U2960 (N_2960,N_2906,N_2882);
or U2961 (N_2961,N_2915,N_2936);
nand U2962 (N_2962,N_2896,N_2930);
xnor U2963 (N_2963,N_2901,N_2895);
or U2964 (N_2964,N_2900,N_2897);
nand U2965 (N_2965,N_2887,N_2904);
xor U2966 (N_2966,N_2932,N_2926);
xnor U2967 (N_2967,N_2916,N_2902);
or U2968 (N_2968,N_2888,N_2927);
and U2969 (N_2969,N_2894,N_2919);
xor U2970 (N_2970,N_2918,N_2912);
or U2971 (N_2971,N_2888,N_2885);
and U2972 (N_2972,N_2911,N_2903);
or U2973 (N_2973,N_2902,N_2894);
xnor U2974 (N_2974,N_2916,N_2931);
xor U2975 (N_2975,N_2917,N_2899);
nor U2976 (N_2976,N_2898,N_2906);
xnor U2977 (N_2977,N_2918,N_2886);
xor U2978 (N_2978,N_2926,N_2913);
nand U2979 (N_2979,N_2886,N_2903);
or U2980 (N_2980,N_2882,N_2884);
or U2981 (N_2981,N_2904,N_2889);
nor U2982 (N_2982,N_2903,N_2938);
nand U2983 (N_2983,N_2909,N_2935);
nor U2984 (N_2984,N_2922,N_2912);
nor U2985 (N_2985,N_2892,N_2899);
or U2986 (N_2986,N_2926,N_2900);
and U2987 (N_2987,N_2891,N_2885);
and U2988 (N_2988,N_2895,N_2903);
or U2989 (N_2989,N_2919,N_2912);
and U2990 (N_2990,N_2880,N_2884);
nor U2991 (N_2991,N_2919,N_2884);
and U2992 (N_2992,N_2903,N_2921);
nor U2993 (N_2993,N_2882,N_2932);
and U2994 (N_2994,N_2880,N_2933);
or U2995 (N_2995,N_2911,N_2880);
xnor U2996 (N_2996,N_2900,N_2919);
or U2997 (N_2997,N_2899,N_2900);
xnor U2998 (N_2998,N_2891,N_2915);
nand U2999 (N_2999,N_2926,N_2888);
or UO_0 (O_0,N_2966,N_2984);
nor UO_1 (O_1,N_2977,N_2982);
and UO_2 (O_2,N_2954,N_2959);
nand UO_3 (O_3,N_2965,N_2979);
and UO_4 (O_4,N_2940,N_2957);
xor UO_5 (O_5,N_2955,N_2986);
xnor UO_6 (O_6,N_2951,N_2950);
nor UO_7 (O_7,N_2996,N_2948);
or UO_8 (O_8,N_2997,N_2941);
nand UO_9 (O_9,N_2945,N_2998);
and UO_10 (O_10,N_2953,N_2992);
nand UO_11 (O_11,N_2949,N_2989);
xnor UO_12 (O_12,N_2968,N_2981);
nor UO_13 (O_13,N_2962,N_2964);
nand UO_14 (O_14,N_2994,N_2991);
or UO_15 (O_15,N_2972,N_2960);
or UO_16 (O_16,N_2983,N_2975);
nand UO_17 (O_17,N_2952,N_2967);
nand UO_18 (O_18,N_2944,N_2980);
nand UO_19 (O_19,N_2990,N_2963);
nand UO_20 (O_20,N_2969,N_2946);
nor UO_21 (O_21,N_2956,N_2958);
nand UO_22 (O_22,N_2970,N_2987);
or UO_23 (O_23,N_2995,N_2988);
and UO_24 (O_24,N_2943,N_2961);
nor UO_25 (O_25,N_2947,N_2999);
nor UO_26 (O_26,N_2973,N_2978);
xnor UO_27 (O_27,N_2993,N_2942);
nor UO_28 (O_28,N_2985,N_2971);
or UO_29 (O_29,N_2976,N_2974);
or UO_30 (O_30,N_2944,N_2940);
nor UO_31 (O_31,N_2978,N_2958);
xor UO_32 (O_32,N_2978,N_2990);
and UO_33 (O_33,N_2956,N_2961);
nand UO_34 (O_34,N_2977,N_2971);
nor UO_35 (O_35,N_2947,N_2993);
nor UO_36 (O_36,N_2972,N_2962);
xnor UO_37 (O_37,N_2969,N_2949);
xnor UO_38 (O_38,N_2948,N_2990);
xor UO_39 (O_39,N_2988,N_2942);
xor UO_40 (O_40,N_2992,N_2973);
nand UO_41 (O_41,N_2957,N_2941);
nand UO_42 (O_42,N_2999,N_2978);
xor UO_43 (O_43,N_2949,N_2990);
xor UO_44 (O_44,N_2947,N_2960);
and UO_45 (O_45,N_2978,N_2995);
nand UO_46 (O_46,N_2944,N_2974);
nand UO_47 (O_47,N_2998,N_2983);
and UO_48 (O_48,N_2985,N_2945);
nand UO_49 (O_49,N_2997,N_2954);
xor UO_50 (O_50,N_2981,N_2977);
nor UO_51 (O_51,N_2990,N_2951);
nor UO_52 (O_52,N_2950,N_2986);
nand UO_53 (O_53,N_2995,N_2955);
xnor UO_54 (O_54,N_2984,N_2953);
xnor UO_55 (O_55,N_2990,N_2952);
or UO_56 (O_56,N_2962,N_2991);
xor UO_57 (O_57,N_2988,N_2998);
and UO_58 (O_58,N_2980,N_2970);
nor UO_59 (O_59,N_2951,N_2980);
or UO_60 (O_60,N_2950,N_2984);
nand UO_61 (O_61,N_2969,N_2966);
nor UO_62 (O_62,N_2965,N_2940);
xnor UO_63 (O_63,N_2944,N_2998);
xnor UO_64 (O_64,N_2986,N_2961);
nand UO_65 (O_65,N_2961,N_2964);
xor UO_66 (O_66,N_2961,N_2985);
and UO_67 (O_67,N_2981,N_2998);
nor UO_68 (O_68,N_2989,N_2975);
xor UO_69 (O_69,N_2956,N_2960);
or UO_70 (O_70,N_2996,N_2993);
or UO_71 (O_71,N_2985,N_2975);
nor UO_72 (O_72,N_2964,N_2948);
nor UO_73 (O_73,N_2966,N_2972);
nand UO_74 (O_74,N_2951,N_2956);
nand UO_75 (O_75,N_2997,N_2976);
nand UO_76 (O_76,N_2948,N_2983);
or UO_77 (O_77,N_2974,N_2994);
nor UO_78 (O_78,N_2951,N_2992);
or UO_79 (O_79,N_2991,N_2980);
xnor UO_80 (O_80,N_2981,N_2988);
or UO_81 (O_81,N_2998,N_2985);
or UO_82 (O_82,N_2957,N_2988);
nand UO_83 (O_83,N_2992,N_2987);
nor UO_84 (O_84,N_2972,N_2949);
and UO_85 (O_85,N_2984,N_2945);
nor UO_86 (O_86,N_2947,N_2979);
xor UO_87 (O_87,N_2945,N_2977);
nand UO_88 (O_88,N_2946,N_2970);
or UO_89 (O_89,N_2974,N_2941);
nor UO_90 (O_90,N_2955,N_2957);
nor UO_91 (O_91,N_2952,N_2974);
xor UO_92 (O_92,N_2948,N_2997);
xnor UO_93 (O_93,N_2983,N_2949);
or UO_94 (O_94,N_2980,N_2967);
nor UO_95 (O_95,N_2988,N_2968);
nand UO_96 (O_96,N_2954,N_2994);
or UO_97 (O_97,N_2940,N_2958);
or UO_98 (O_98,N_2952,N_2959);
and UO_99 (O_99,N_2941,N_2998);
and UO_100 (O_100,N_2992,N_2999);
or UO_101 (O_101,N_2964,N_2979);
nor UO_102 (O_102,N_2964,N_2991);
nand UO_103 (O_103,N_2947,N_2975);
xnor UO_104 (O_104,N_2969,N_2993);
nand UO_105 (O_105,N_2950,N_2992);
nor UO_106 (O_106,N_2958,N_2996);
nor UO_107 (O_107,N_2958,N_2952);
nor UO_108 (O_108,N_2942,N_2956);
xnor UO_109 (O_109,N_2967,N_2953);
and UO_110 (O_110,N_2951,N_2971);
and UO_111 (O_111,N_2963,N_2958);
nand UO_112 (O_112,N_2961,N_2982);
xnor UO_113 (O_113,N_2970,N_2949);
and UO_114 (O_114,N_2996,N_2951);
or UO_115 (O_115,N_2983,N_2996);
nor UO_116 (O_116,N_2986,N_2951);
xor UO_117 (O_117,N_2989,N_2959);
nor UO_118 (O_118,N_2965,N_2950);
or UO_119 (O_119,N_2959,N_2964);
or UO_120 (O_120,N_2987,N_2983);
or UO_121 (O_121,N_2962,N_2987);
xnor UO_122 (O_122,N_2958,N_2945);
xor UO_123 (O_123,N_2997,N_2974);
nand UO_124 (O_124,N_2942,N_2992);
and UO_125 (O_125,N_2979,N_2997);
or UO_126 (O_126,N_2944,N_2979);
or UO_127 (O_127,N_2942,N_2978);
or UO_128 (O_128,N_2973,N_2993);
and UO_129 (O_129,N_2970,N_2979);
nand UO_130 (O_130,N_2940,N_2946);
and UO_131 (O_131,N_2993,N_2986);
nand UO_132 (O_132,N_2984,N_2972);
or UO_133 (O_133,N_2987,N_2966);
and UO_134 (O_134,N_2979,N_2992);
nor UO_135 (O_135,N_2968,N_2996);
xnor UO_136 (O_136,N_2979,N_2957);
xnor UO_137 (O_137,N_2977,N_2986);
nor UO_138 (O_138,N_2987,N_2946);
nand UO_139 (O_139,N_2950,N_2941);
or UO_140 (O_140,N_2946,N_2955);
nor UO_141 (O_141,N_2969,N_2991);
and UO_142 (O_142,N_2979,N_2961);
nor UO_143 (O_143,N_2952,N_2986);
nor UO_144 (O_144,N_2985,N_2940);
xor UO_145 (O_145,N_2963,N_2973);
nor UO_146 (O_146,N_2971,N_2997);
or UO_147 (O_147,N_2983,N_2953);
xnor UO_148 (O_148,N_2976,N_2956);
or UO_149 (O_149,N_2997,N_2955);
or UO_150 (O_150,N_2971,N_2946);
or UO_151 (O_151,N_2953,N_2990);
xor UO_152 (O_152,N_2963,N_2983);
nor UO_153 (O_153,N_2991,N_2955);
and UO_154 (O_154,N_2942,N_2941);
nand UO_155 (O_155,N_2948,N_2942);
nor UO_156 (O_156,N_2957,N_2999);
and UO_157 (O_157,N_2950,N_2987);
nand UO_158 (O_158,N_2948,N_2944);
nor UO_159 (O_159,N_2992,N_2956);
xnor UO_160 (O_160,N_2962,N_2995);
and UO_161 (O_161,N_2997,N_2977);
xnor UO_162 (O_162,N_2959,N_2974);
or UO_163 (O_163,N_2946,N_2967);
xnor UO_164 (O_164,N_2993,N_2960);
or UO_165 (O_165,N_2984,N_2943);
and UO_166 (O_166,N_2948,N_2940);
or UO_167 (O_167,N_2945,N_2953);
or UO_168 (O_168,N_2970,N_2955);
and UO_169 (O_169,N_2981,N_2945);
nor UO_170 (O_170,N_2963,N_2976);
nor UO_171 (O_171,N_2947,N_2973);
and UO_172 (O_172,N_2974,N_2947);
or UO_173 (O_173,N_2962,N_2996);
or UO_174 (O_174,N_2996,N_2997);
nand UO_175 (O_175,N_2954,N_2964);
nand UO_176 (O_176,N_2963,N_2972);
or UO_177 (O_177,N_2989,N_2940);
nand UO_178 (O_178,N_2993,N_2951);
and UO_179 (O_179,N_2999,N_2940);
nand UO_180 (O_180,N_2977,N_2940);
and UO_181 (O_181,N_2971,N_2957);
nor UO_182 (O_182,N_2984,N_2949);
and UO_183 (O_183,N_2944,N_2947);
or UO_184 (O_184,N_2973,N_2954);
and UO_185 (O_185,N_2957,N_2965);
and UO_186 (O_186,N_2980,N_2948);
or UO_187 (O_187,N_2985,N_2948);
nand UO_188 (O_188,N_2970,N_2974);
or UO_189 (O_189,N_2991,N_2966);
nand UO_190 (O_190,N_2967,N_2973);
or UO_191 (O_191,N_2985,N_2987);
and UO_192 (O_192,N_2961,N_2992);
xnor UO_193 (O_193,N_2963,N_2956);
nor UO_194 (O_194,N_2979,N_2981);
nand UO_195 (O_195,N_2965,N_2982);
nor UO_196 (O_196,N_2949,N_2940);
or UO_197 (O_197,N_2953,N_2999);
xnor UO_198 (O_198,N_2982,N_2978);
xnor UO_199 (O_199,N_2994,N_2944);
or UO_200 (O_200,N_2967,N_2996);
or UO_201 (O_201,N_2969,N_2948);
or UO_202 (O_202,N_2989,N_2974);
and UO_203 (O_203,N_2960,N_2989);
nand UO_204 (O_204,N_2948,N_2991);
nand UO_205 (O_205,N_2982,N_2942);
or UO_206 (O_206,N_2973,N_2946);
nor UO_207 (O_207,N_2965,N_2984);
nor UO_208 (O_208,N_2966,N_2962);
and UO_209 (O_209,N_2959,N_2948);
nor UO_210 (O_210,N_2963,N_2970);
nor UO_211 (O_211,N_2993,N_2984);
nand UO_212 (O_212,N_2988,N_2989);
xor UO_213 (O_213,N_2963,N_2969);
or UO_214 (O_214,N_2958,N_2951);
and UO_215 (O_215,N_2960,N_2946);
or UO_216 (O_216,N_2953,N_2991);
or UO_217 (O_217,N_2985,N_2988);
and UO_218 (O_218,N_2953,N_2966);
nor UO_219 (O_219,N_2966,N_2951);
nor UO_220 (O_220,N_2960,N_2948);
nor UO_221 (O_221,N_2987,N_2978);
nand UO_222 (O_222,N_2961,N_2995);
nor UO_223 (O_223,N_2962,N_2999);
or UO_224 (O_224,N_2944,N_2960);
nor UO_225 (O_225,N_2943,N_2949);
nor UO_226 (O_226,N_2973,N_2988);
nor UO_227 (O_227,N_2943,N_2948);
nor UO_228 (O_228,N_2943,N_2993);
nor UO_229 (O_229,N_2961,N_2974);
and UO_230 (O_230,N_2946,N_2948);
and UO_231 (O_231,N_2981,N_2978);
nor UO_232 (O_232,N_2979,N_2975);
nand UO_233 (O_233,N_2941,N_2973);
xnor UO_234 (O_234,N_2955,N_2959);
and UO_235 (O_235,N_2991,N_2959);
nor UO_236 (O_236,N_2986,N_2941);
xnor UO_237 (O_237,N_2951,N_2944);
or UO_238 (O_238,N_2949,N_2964);
nand UO_239 (O_239,N_2956,N_2983);
or UO_240 (O_240,N_2984,N_2971);
and UO_241 (O_241,N_2950,N_2975);
or UO_242 (O_242,N_2940,N_2967);
nor UO_243 (O_243,N_2981,N_2975);
nand UO_244 (O_244,N_2992,N_2989);
xnor UO_245 (O_245,N_2944,N_2986);
or UO_246 (O_246,N_2946,N_2990);
or UO_247 (O_247,N_2983,N_2950);
nand UO_248 (O_248,N_2985,N_2982);
nand UO_249 (O_249,N_2962,N_2941);
nor UO_250 (O_250,N_2951,N_2960);
xnor UO_251 (O_251,N_2999,N_2952);
xor UO_252 (O_252,N_2980,N_2963);
or UO_253 (O_253,N_2943,N_2946);
nor UO_254 (O_254,N_2945,N_2990);
xor UO_255 (O_255,N_2944,N_2942);
xor UO_256 (O_256,N_2992,N_2947);
and UO_257 (O_257,N_2999,N_2987);
and UO_258 (O_258,N_2949,N_2951);
and UO_259 (O_259,N_2958,N_2991);
and UO_260 (O_260,N_2979,N_2950);
xnor UO_261 (O_261,N_2959,N_2986);
nand UO_262 (O_262,N_2998,N_2940);
nor UO_263 (O_263,N_2998,N_2950);
nand UO_264 (O_264,N_2977,N_2999);
or UO_265 (O_265,N_2981,N_2963);
or UO_266 (O_266,N_2981,N_2972);
or UO_267 (O_267,N_2955,N_2982);
nor UO_268 (O_268,N_2968,N_2957);
and UO_269 (O_269,N_2961,N_2959);
or UO_270 (O_270,N_2961,N_2977);
xor UO_271 (O_271,N_2951,N_2968);
xnor UO_272 (O_272,N_2943,N_2955);
nand UO_273 (O_273,N_2945,N_2955);
or UO_274 (O_274,N_2961,N_2944);
or UO_275 (O_275,N_2959,N_2984);
and UO_276 (O_276,N_2958,N_2987);
or UO_277 (O_277,N_2970,N_2953);
and UO_278 (O_278,N_2970,N_2981);
or UO_279 (O_279,N_2981,N_2951);
nand UO_280 (O_280,N_2963,N_2943);
nor UO_281 (O_281,N_2970,N_2959);
nor UO_282 (O_282,N_2996,N_2989);
or UO_283 (O_283,N_2951,N_2994);
nor UO_284 (O_284,N_2993,N_2945);
and UO_285 (O_285,N_2943,N_2999);
nand UO_286 (O_286,N_2973,N_2990);
xor UO_287 (O_287,N_2971,N_2942);
nand UO_288 (O_288,N_2972,N_2970);
and UO_289 (O_289,N_2989,N_2993);
nor UO_290 (O_290,N_2982,N_2945);
nor UO_291 (O_291,N_2945,N_2950);
nor UO_292 (O_292,N_2942,N_2997);
xnor UO_293 (O_293,N_2970,N_2943);
nand UO_294 (O_294,N_2985,N_2950);
nand UO_295 (O_295,N_2993,N_2990);
or UO_296 (O_296,N_2983,N_2985);
or UO_297 (O_297,N_2950,N_2981);
nand UO_298 (O_298,N_2954,N_2948);
nor UO_299 (O_299,N_2946,N_2997);
xnor UO_300 (O_300,N_2947,N_2988);
or UO_301 (O_301,N_2997,N_2975);
or UO_302 (O_302,N_2976,N_2968);
nand UO_303 (O_303,N_2966,N_2958);
nand UO_304 (O_304,N_2979,N_2955);
nand UO_305 (O_305,N_2964,N_2978);
nand UO_306 (O_306,N_2978,N_2991);
nor UO_307 (O_307,N_2999,N_2960);
xor UO_308 (O_308,N_2995,N_2971);
or UO_309 (O_309,N_2964,N_2990);
xor UO_310 (O_310,N_2949,N_2968);
nor UO_311 (O_311,N_2978,N_2984);
or UO_312 (O_312,N_2967,N_2959);
xor UO_313 (O_313,N_2954,N_2998);
nor UO_314 (O_314,N_2976,N_2987);
xor UO_315 (O_315,N_2980,N_2978);
nand UO_316 (O_316,N_2976,N_2967);
nand UO_317 (O_317,N_2976,N_2996);
nand UO_318 (O_318,N_2988,N_2945);
or UO_319 (O_319,N_2964,N_2960);
nor UO_320 (O_320,N_2978,N_2969);
nand UO_321 (O_321,N_2973,N_2965);
or UO_322 (O_322,N_2963,N_2984);
or UO_323 (O_323,N_2970,N_2950);
or UO_324 (O_324,N_2965,N_2958);
and UO_325 (O_325,N_2972,N_2969);
and UO_326 (O_326,N_2980,N_2974);
xnor UO_327 (O_327,N_2956,N_2948);
or UO_328 (O_328,N_2999,N_2966);
nor UO_329 (O_329,N_2991,N_2942);
xnor UO_330 (O_330,N_2983,N_2945);
and UO_331 (O_331,N_2963,N_2975);
and UO_332 (O_332,N_2954,N_2956);
or UO_333 (O_333,N_2966,N_2996);
nand UO_334 (O_334,N_2945,N_2963);
or UO_335 (O_335,N_2981,N_2992);
xor UO_336 (O_336,N_2962,N_2978);
xnor UO_337 (O_337,N_2996,N_2952);
or UO_338 (O_338,N_2946,N_2947);
or UO_339 (O_339,N_2978,N_2993);
nor UO_340 (O_340,N_2977,N_2995);
nand UO_341 (O_341,N_2993,N_2977);
and UO_342 (O_342,N_2944,N_2950);
and UO_343 (O_343,N_2989,N_2977);
and UO_344 (O_344,N_2991,N_2995);
and UO_345 (O_345,N_2984,N_2956);
nand UO_346 (O_346,N_2958,N_2970);
xor UO_347 (O_347,N_2948,N_2984);
and UO_348 (O_348,N_2988,N_2944);
nand UO_349 (O_349,N_2946,N_2983);
and UO_350 (O_350,N_2953,N_2976);
or UO_351 (O_351,N_2995,N_2946);
nor UO_352 (O_352,N_2977,N_2969);
xor UO_353 (O_353,N_2971,N_2993);
xor UO_354 (O_354,N_2961,N_2966);
or UO_355 (O_355,N_2996,N_2944);
xnor UO_356 (O_356,N_2995,N_2969);
and UO_357 (O_357,N_2985,N_2981);
nor UO_358 (O_358,N_2962,N_2988);
nand UO_359 (O_359,N_2952,N_2945);
nand UO_360 (O_360,N_2953,N_2942);
nand UO_361 (O_361,N_2972,N_2940);
or UO_362 (O_362,N_2949,N_2985);
nand UO_363 (O_363,N_2994,N_2957);
xor UO_364 (O_364,N_2979,N_2943);
nand UO_365 (O_365,N_2996,N_2995);
and UO_366 (O_366,N_2962,N_2979);
and UO_367 (O_367,N_2995,N_2982);
xor UO_368 (O_368,N_2965,N_2972);
nor UO_369 (O_369,N_2967,N_2984);
nor UO_370 (O_370,N_2970,N_2964);
or UO_371 (O_371,N_2962,N_2970);
nand UO_372 (O_372,N_2974,N_2990);
nand UO_373 (O_373,N_2974,N_2963);
or UO_374 (O_374,N_2970,N_2965);
nand UO_375 (O_375,N_2982,N_2941);
xnor UO_376 (O_376,N_2969,N_2940);
nor UO_377 (O_377,N_2963,N_2965);
nand UO_378 (O_378,N_2992,N_2945);
nand UO_379 (O_379,N_2996,N_2979);
or UO_380 (O_380,N_2940,N_2980);
xnor UO_381 (O_381,N_2998,N_2953);
nor UO_382 (O_382,N_2988,N_2980);
and UO_383 (O_383,N_2981,N_2948);
nor UO_384 (O_384,N_2984,N_2951);
xor UO_385 (O_385,N_2967,N_2986);
nand UO_386 (O_386,N_2989,N_2943);
and UO_387 (O_387,N_2987,N_2968);
nor UO_388 (O_388,N_2974,N_2965);
nand UO_389 (O_389,N_2983,N_2992);
or UO_390 (O_390,N_2982,N_2973);
nand UO_391 (O_391,N_2959,N_2992);
nor UO_392 (O_392,N_2996,N_2956);
or UO_393 (O_393,N_2993,N_2979);
nor UO_394 (O_394,N_2978,N_2957);
nand UO_395 (O_395,N_2956,N_2945);
and UO_396 (O_396,N_2948,N_2987);
xnor UO_397 (O_397,N_2962,N_2957);
and UO_398 (O_398,N_2952,N_2981);
nor UO_399 (O_399,N_2967,N_2985);
or UO_400 (O_400,N_2978,N_2988);
nor UO_401 (O_401,N_2951,N_2945);
and UO_402 (O_402,N_2973,N_2951);
xor UO_403 (O_403,N_2970,N_2975);
or UO_404 (O_404,N_2952,N_2991);
xor UO_405 (O_405,N_2957,N_2982);
nor UO_406 (O_406,N_2975,N_2952);
xnor UO_407 (O_407,N_2952,N_2971);
and UO_408 (O_408,N_2990,N_2988);
nand UO_409 (O_409,N_2969,N_2998);
xnor UO_410 (O_410,N_2941,N_2959);
nor UO_411 (O_411,N_2941,N_2940);
and UO_412 (O_412,N_2949,N_2966);
nand UO_413 (O_413,N_2997,N_2952);
or UO_414 (O_414,N_2967,N_2966);
or UO_415 (O_415,N_2993,N_2985);
or UO_416 (O_416,N_2970,N_2995);
and UO_417 (O_417,N_2958,N_2967);
xnor UO_418 (O_418,N_2998,N_2946);
and UO_419 (O_419,N_2947,N_2991);
nand UO_420 (O_420,N_2954,N_2988);
nor UO_421 (O_421,N_2954,N_2992);
xnor UO_422 (O_422,N_2958,N_2995);
or UO_423 (O_423,N_2968,N_2984);
nor UO_424 (O_424,N_2988,N_2969);
or UO_425 (O_425,N_2998,N_2996);
nor UO_426 (O_426,N_2940,N_2994);
xor UO_427 (O_427,N_2986,N_2962);
nor UO_428 (O_428,N_2966,N_2976);
xnor UO_429 (O_429,N_2992,N_2997);
or UO_430 (O_430,N_2976,N_2950);
nand UO_431 (O_431,N_2963,N_2977);
nor UO_432 (O_432,N_2951,N_2976);
nand UO_433 (O_433,N_2943,N_2994);
xor UO_434 (O_434,N_2949,N_2980);
or UO_435 (O_435,N_2990,N_2944);
xnor UO_436 (O_436,N_2976,N_2962);
or UO_437 (O_437,N_2995,N_2940);
xor UO_438 (O_438,N_2971,N_2972);
xor UO_439 (O_439,N_2969,N_2974);
and UO_440 (O_440,N_2980,N_2998);
or UO_441 (O_441,N_2950,N_2969);
xnor UO_442 (O_442,N_2964,N_2965);
xnor UO_443 (O_443,N_2999,N_2949);
xnor UO_444 (O_444,N_2960,N_2943);
nand UO_445 (O_445,N_2943,N_2951);
nor UO_446 (O_446,N_2982,N_2962);
or UO_447 (O_447,N_2953,N_2989);
nand UO_448 (O_448,N_2941,N_2945);
nor UO_449 (O_449,N_2995,N_2960);
and UO_450 (O_450,N_2948,N_2976);
xnor UO_451 (O_451,N_2978,N_2971);
and UO_452 (O_452,N_2966,N_2978);
nor UO_453 (O_453,N_2941,N_2963);
or UO_454 (O_454,N_2952,N_2948);
xor UO_455 (O_455,N_2977,N_2996);
nor UO_456 (O_456,N_2951,N_2974);
nand UO_457 (O_457,N_2989,N_2961);
nand UO_458 (O_458,N_2986,N_2960);
nand UO_459 (O_459,N_2972,N_2980);
and UO_460 (O_460,N_2988,N_2996);
and UO_461 (O_461,N_2942,N_2945);
nor UO_462 (O_462,N_2973,N_2945);
nand UO_463 (O_463,N_2944,N_2970);
nand UO_464 (O_464,N_2952,N_2963);
nor UO_465 (O_465,N_2946,N_2965);
xnor UO_466 (O_466,N_2961,N_2975);
nor UO_467 (O_467,N_2964,N_2973);
and UO_468 (O_468,N_2941,N_2994);
or UO_469 (O_469,N_2951,N_2978);
or UO_470 (O_470,N_2970,N_2947);
xnor UO_471 (O_471,N_2971,N_2948);
nand UO_472 (O_472,N_2999,N_2969);
nor UO_473 (O_473,N_2983,N_2944);
nand UO_474 (O_474,N_2953,N_2997);
and UO_475 (O_475,N_2977,N_2944);
or UO_476 (O_476,N_2976,N_2984);
or UO_477 (O_477,N_2978,N_2974);
or UO_478 (O_478,N_2947,N_2966);
and UO_479 (O_479,N_2967,N_2947);
or UO_480 (O_480,N_2956,N_2990);
or UO_481 (O_481,N_2982,N_2953);
xnor UO_482 (O_482,N_2987,N_2991);
nand UO_483 (O_483,N_2995,N_2979);
nor UO_484 (O_484,N_2952,N_2964);
or UO_485 (O_485,N_2940,N_2959);
nor UO_486 (O_486,N_2985,N_2947);
nor UO_487 (O_487,N_2992,N_2943);
xor UO_488 (O_488,N_2968,N_2979);
or UO_489 (O_489,N_2989,N_2966);
or UO_490 (O_490,N_2967,N_2969);
nand UO_491 (O_491,N_2941,N_2960);
or UO_492 (O_492,N_2944,N_2965);
xnor UO_493 (O_493,N_2987,N_2949);
xnor UO_494 (O_494,N_2988,N_2983);
and UO_495 (O_495,N_2985,N_2966);
xor UO_496 (O_496,N_2979,N_2988);
nand UO_497 (O_497,N_2955,N_2988);
nand UO_498 (O_498,N_2942,N_2965);
nand UO_499 (O_499,N_2989,N_2980);
endmodule