module basic_750_5000_1000_5_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_229,In_85);
nor U1 (N_1,In_200,In_430);
nor U2 (N_2,In_723,In_24);
nor U3 (N_3,In_467,In_80);
and U4 (N_4,In_511,In_523);
or U5 (N_5,In_233,In_259);
nor U6 (N_6,In_337,In_654);
or U7 (N_7,In_600,In_57);
and U8 (N_8,In_694,In_652);
nor U9 (N_9,In_223,In_577);
nor U10 (N_10,In_52,In_714);
and U11 (N_11,In_417,In_580);
nand U12 (N_12,In_28,In_728);
and U13 (N_13,In_552,In_492);
or U14 (N_14,In_746,In_373);
nand U15 (N_15,In_571,In_644);
or U16 (N_16,In_206,In_634);
or U17 (N_17,In_579,In_367);
nor U18 (N_18,In_357,In_463);
nor U19 (N_19,In_385,In_231);
nand U20 (N_20,In_667,In_697);
and U21 (N_21,In_464,In_447);
nand U22 (N_22,In_480,In_213);
and U23 (N_23,In_736,In_685);
or U24 (N_24,In_732,In_387);
nor U25 (N_25,In_225,In_495);
or U26 (N_26,In_699,In_614);
or U27 (N_27,In_638,In_451);
and U28 (N_28,In_674,In_731);
or U29 (N_29,In_352,In_1);
or U30 (N_30,In_358,In_635);
nor U31 (N_31,In_339,In_219);
or U32 (N_32,In_345,In_419);
nor U33 (N_33,In_221,In_60);
or U34 (N_34,In_74,In_163);
nand U35 (N_35,In_636,In_709);
nor U36 (N_36,In_598,In_449);
nand U37 (N_37,In_499,In_216);
and U38 (N_38,In_741,In_621);
nand U39 (N_39,In_313,In_136);
and U40 (N_40,In_536,In_189);
nor U41 (N_41,In_659,In_502);
nand U42 (N_42,In_76,In_214);
nand U43 (N_43,In_331,In_38);
nor U44 (N_44,In_174,In_362);
nor U45 (N_45,In_164,In_545);
nor U46 (N_46,In_128,In_663);
or U47 (N_47,In_627,In_186);
nor U48 (N_48,In_75,In_330);
and U49 (N_49,In_108,In_440);
nand U50 (N_50,In_435,In_386);
and U51 (N_51,In_530,In_183);
and U52 (N_52,In_281,In_326);
or U53 (N_53,In_733,In_740);
or U54 (N_54,In_743,In_411);
or U55 (N_55,In_261,In_372);
nand U56 (N_56,In_171,In_623);
nand U57 (N_57,In_524,In_309);
and U58 (N_58,In_421,In_143);
and U59 (N_59,In_263,In_528);
and U60 (N_60,In_209,In_490);
nor U61 (N_61,In_278,In_275);
xor U62 (N_62,In_413,In_248);
nand U63 (N_63,In_302,In_356);
or U64 (N_64,In_703,In_376);
or U65 (N_65,In_744,In_283);
or U66 (N_66,In_30,In_42);
nor U67 (N_67,In_119,In_153);
nand U68 (N_68,In_62,In_101);
or U69 (N_69,In_624,In_25);
and U70 (N_70,In_486,In_519);
nor U71 (N_71,In_604,In_154);
nand U72 (N_72,In_525,In_71);
nand U73 (N_73,In_178,In_110);
and U74 (N_74,In_250,In_687);
and U75 (N_75,In_144,In_498);
and U76 (N_76,In_238,In_12);
and U77 (N_77,In_43,In_48);
and U78 (N_78,In_518,In_510);
or U79 (N_79,In_246,In_645);
and U80 (N_80,In_488,In_64);
nand U81 (N_81,In_179,In_120);
or U82 (N_82,In_400,In_290);
nor U83 (N_83,In_658,In_734);
nor U84 (N_84,In_70,In_137);
nand U85 (N_85,In_68,In_454);
nand U86 (N_86,In_550,In_701);
nor U87 (N_87,In_90,In_425);
nor U88 (N_88,In_141,In_155);
nand U89 (N_89,In_148,In_93);
nor U90 (N_90,In_226,In_91);
nand U91 (N_91,In_202,In_256);
nor U92 (N_92,In_49,In_513);
nand U93 (N_93,In_472,In_465);
and U94 (N_94,In_737,In_404);
nand U95 (N_95,In_279,In_514);
nand U96 (N_96,In_210,In_505);
nand U97 (N_97,In_460,In_265);
nor U98 (N_98,In_98,In_158);
nor U99 (N_99,In_424,In_170);
xor U100 (N_100,In_156,In_615);
and U101 (N_101,In_506,In_77);
or U102 (N_102,In_686,In_132);
or U103 (N_103,In_348,In_271);
and U104 (N_104,In_560,In_18);
and U105 (N_105,In_642,In_34);
nand U106 (N_106,In_33,In_551);
nand U107 (N_107,In_471,In_570);
nand U108 (N_108,In_707,In_704);
nand U109 (N_109,In_36,In_359);
nor U110 (N_110,In_181,In_720);
nand U111 (N_111,In_347,In_626);
nand U112 (N_112,In_520,In_608);
nand U113 (N_113,In_415,In_201);
or U114 (N_114,In_702,In_205);
or U115 (N_115,In_602,In_355);
or U116 (N_116,In_344,In_211);
or U117 (N_117,In_380,In_241);
nand U118 (N_118,In_9,In_393);
nand U119 (N_119,In_187,In_611);
or U120 (N_120,In_239,In_478);
nor U121 (N_121,In_630,In_321);
or U122 (N_122,In_595,In_215);
nor U123 (N_123,In_522,In_414);
nand U124 (N_124,In_657,In_185);
or U125 (N_125,In_546,In_81);
nand U126 (N_126,In_294,In_289);
or U127 (N_127,In_117,In_199);
nor U128 (N_128,In_377,In_27);
nor U129 (N_129,In_473,In_656);
or U130 (N_130,In_675,In_484);
nand U131 (N_131,In_257,In_39);
nor U132 (N_132,In_323,In_103);
nor U133 (N_133,In_287,In_169);
nor U134 (N_134,In_547,In_455);
or U135 (N_135,In_274,In_721);
or U136 (N_136,In_237,In_182);
and U137 (N_137,In_651,In_742);
nor U138 (N_138,In_708,In_613);
or U139 (N_139,In_135,In_670);
or U140 (N_140,In_422,In_403);
or U141 (N_141,In_353,In_44);
or U142 (N_142,In_224,In_63);
or U143 (N_143,In_553,In_268);
and U144 (N_144,In_418,In_692);
and U145 (N_145,In_253,In_409);
nand U146 (N_146,In_612,In_240);
or U147 (N_147,In_647,In_264);
nor U148 (N_148,In_269,In_462);
xor U149 (N_149,In_105,In_625);
and U150 (N_150,In_533,In_21);
nor U151 (N_151,In_705,In_310);
and U152 (N_152,In_254,In_456);
nand U153 (N_153,In_540,In_561);
or U154 (N_154,In_354,In_138);
nor U155 (N_155,In_503,In_94);
nor U156 (N_156,In_730,In_47);
nand U157 (N_157,In_679,In_690);
nor U158 (N_158,In_102,In_333);
and U159 (N_159,In_350,In_107);
and U160 (N_160,In_361,In_84);
nor U161 (N_161,In_207,In_433);
or U162 (N_162,In_660,In_485);
nand U163 (N_163,In_575,In_459);
nor U164 (N_164,In_682,In_437);
nor U165 (N_165,In_191,In_335);
or U166 (N_166,In_678,In_672);
nor U167 (N_167,In_517,In_639);
and U168 (N_168,In_100,In_125);
xor U169 (N_169,In_583,In_17);
nand U170 (N_170,In_481,In_710);
nor U171 (N_171,In_311,In_655);
nor U172 (N_172,In_222,In_130);
nor U173 (N_173,In_662,In_606);
nand U174 (N_174,In_266,In_516);
and U175 (N_175,In_726,In_369);
nor U176 (N_176,In_487,In_439);
and U177 (N_177,In_35,In_477);
nor U178 (N_178,In_747,In_695);
or U179 (N_179,In_244,In_434);
nand U180 (N_180,In_578,In_151);
nand U181 (N_181,In_104,In_234);
nand U182 (N_182,In_51,In_431);
nand U183 (N_183,In_436,In_122);
and U184 (N_184,In_383,In_500);
and U185 (N_185,In_166,In_304);
and U186 (N_186,In_297,In_748);
and U187 (N_187,In_296,In_509);
and U188 (N_188,In_328,In_563);
or U189 (N_189,In_150,In_251);
nor U190 (N_190,In_474,In_618);
or U191 (N_191,In_194,In_295);
nand U192 (N_192,In_394,In_568);
nor U193 (N_193,In_89,In_458);
nand U194 (N_194,In_360,In_581);
and U195 (N_195,In_32,In_681);
or U196 (N_196,In_452,In_307);
nor U197 (N_197,In_589,In_529);
or U198 (N_198,In_527,In_649);
or U199 (N_199,In_338,In_446);
and U200 (N_200,In_212,In_515);
or U201 (N_201,In_72,In_537);
nor U202 (N_202,In_305,In_620);
nor U203 (N_203,In_468,In_343);
and U204 (N_204,In_466,In_719);
nor U205 (N_205,In_31,In_558);
or U206 (N_206,In_322,In_97);
nand U207 (N_207,In_725,In_26);
nor U208 (N_208,In_83,In_324);
nor U209 (N_209,In_41,In_508);
or U210 (N_210,In_374,In_147);
nor U211 (N_211,In_738,In_381);
nor U212 (N_212,In_13,In_395);
and U213 (N_213,In_448,In_10);
nor U214 (N_214,In_650,In_96);
and U215 (N_215,In_316,In_365);
and U216 (N_216,In_111,In_619);
or U217 (N_217,In_562,In_628);
nand U218 (N_218,In_450,In_469);
and U219 (N_219,In_364,In_689);
and U220 (N_220,In_121,In_521);
nor U221 (N_221,In_665,In_482);
nor U222 (N_222,In_228,In_336);
and U223 (N_223,In_476,In_190);
and U224 (N_224,In_493,In_483);
and U225 (N_225,In_584,In_198);
and U226 (N_226,In_539,In_693);
nor U227 (N_227,In_175,In_286);
or U228 (N_228,In_315,In_673);
and U229 (N_229,In_66,In_292);
and U230 (N_230,In_716,In_291);
nand U231 (N_231,In_272,In_165);
nor U232 (N_232,In_669,In_507);
nor U233 (N_233,In_88,In_573);
and U234 (N_234,In_399,In_340);
or U235 (N_235,In_14,In_59);
and U236 (N_236,In_423,In_20);
and U237 (N_237,In_653,In_327);
and U238 (N_238,In_270,In_582);
or U239 (N_239,In_129,In_236);
and U240 (N_240,In_549,In_177);
or U241 (N_241,In_16,In_162);
nor U242 (N_242,In_371,In_384);
nand U243 (N_243,In_306,In_643);
nand U244 (N_244,In_410,In_366);
nand U245 (N_245,In_109,In_401);
and U246 (N_246,In_173,In_123);
and U247 (N_247,In_574,In_11);
and U248 (N_248,In_61,In_632);
or U249 (N_249,In_140,In_646);
nand U250 (N_250,In_739,In_588);
nor U251 (N_251,In_698,In_176);
or U252 (N_252,In_641,In_79);
or U253 (N_253,In_406,In_334);
and U254 (N_254,In_443,In_0);
nand U255 (N_255,In_392,In_255);
nor U256 (N_256,In_599,In_408);
or U257 (N_257,In_260,In_548);
and U258 (N_258,In_696,In_388);
or U259 (N_259,In_55,In_567);
or U260 (N_260,In_161,In_616);
or U261 (N_261,In_479,In_149);
nor U262 (N_262,In_727,In_622);
nand U263 (N_263,In_368,In_609);
nor U264 (N_264,In_19,In_273);
nand U265 (N_265,In_203,In_557);
xor U266 (N_266,In_3,In_92);
and U267 (N_267,In_106,In_113);
nor U268 (N_268,In_501,In_197);
nor U269 (N_269,In_188,In_142);
or U270 (N_270,In_40,In_133);
or U271 (N_271,In_668,In_314);
nand U272 (N_272,In_543,In_299);
nand U273 (N_273,In_717,In_412);
nand U274 (N_274,In_526,In_489);
and U275 (N_275,In_5,In_230);
or U276 (N_276,In_405,In_45);
nand U277 (N_277,In_438,In_308);
or U278 (N_278,In_95,In_576);
nand U279 (N_279,In_82,In_683);
or U280 (N_280,In_303,In_564);
or U281 (N_281,In_131,In_217);
or U282 (N_282,In_29,In_535);
or U283 (N_283,In_73,In_8);
or U284 (N_284,In_99,In_470);
and U285 (N_285,In_134,In_218);
or U286 (N_286,In_2,In_6);
nand U287 (N_287,In_152,In_288);
or U288 (N_288,In_724,In_637);
nand U289 (N_289,In_592,In_688);
nor U290 (N_290,In_23,In_204);
nand U291 (N_291,In_180,In_69);
nor U292 (N_292,In_341,In_318);
nor U293 (N_293,In_594,In_370);
nand U294 (N_294,In_745,In_284);
nor U295 (N_295,In_749,In_713);
or U296 (N_296,In_596,In_684);
or U297 (N_297,In_160,In_661);
nand U298 (N_298,In_512,In_116);
and U299 (N_299,In_37,In_46);
nand U300 (N_300,In_53,In_559);
or U301 (N_301,In_245,In_262);
or U302 (N_302,In_54,In_7);
or U303 (N_303,In_428,In_610);
nor U304 (N_304,In_67,In_544);
nand U305 (N_305,In_640,In_398);
nor U306 (N_306,In_249,In_617);
or U307 (N_307,In_633,In_298);
nor U308 (N_308,In_396,In_232);
nor U309 (N_309,In_711,In_397);
and U310 (N_310,In_461,In_700);
and U311 (N_311,In_587,In_677);
nor U312 (N_312,In_591,In_208);
or U313 (N_313,In_597,In_293);
nor U314 (N_314,In_127,In_494);
nand U315 (N_315,In_607,In_715);
nand U316 (N_316,In_300,In_504);
or U317 (N_317,In_534,In_15);
or U318 (N_318,In_325,In_402);
and U319 (N_319,In_301,In_554);
or U320 (N_320,In_58,In_193);
or U321 (N_321,In_195,In_735);
nand U322 (N_322,In_168,In_227);
nand U323 (N_323,In_457,In_220);
and U324 (N_324,In_247,In_124);
nor U325 (N_325,In_192,In_382);
and U326 (N_326,In_444,In_680);
or U327 (N_327,In_442,In_429);
and U328 (N_328,In_565,In_349);
nor U329 (N_329,In_729,In_586);
nand U330 (N_330,In_541,In_605);
and U331 (N_331,In_242,In_351);
nor U332 (N_332,In_139,In_426);
and U333 (N_333,In_258,In_555);
and U334 (N_334,In_78,In_390);
nand U335 (N_335,In_445,In_332);
and U336 (N_336,In_648,In_346);
nor U337 (N_337,In_496,In_664);
nor U338 (N_338,In_391,In_722);
nand U339 (N_339,In_432,In_172);
nor U340 (N_340,In_497,In_556);
nor U341 (N_341,In_112,In_718);
or U342 (N_342,In_407,In_319);
and U343 (N_343,In_629,In_569);
or U344 (N_344,In_56,In_566);
or U345 (N_345,In_671,In_65);
nand U346 (N_346,In_375,In_243);
nor U347 (N_347,In_196,In_542);
nor U348 (N_348,In_691,In_593);
nand U349 (N_349,In_145,In_538);
and U350 (N_350,In_666,In_453);
or U351 (N_351,In_416,In_475);
and U352 (N_352,In_267,In_276);
and U353 (N_353,In_378,In_157);
or U354 (N_354,In_4,In_320);
nand U355 (N_355,In_631,In_572);
nand U356 (N_356,In_342,In_585);
nor U357 (N_357,In_252,In_118);
and U358 (N_358,In_285,In_427);
nand U359 (N_359,In_184,In_676);
and U360 (N_360,In_532,In_235);
or U361 (N_361,In_420,In_50);
nor U362 (N_362,In_87,In_22);
nor U363 (N_363,In_706,In_167);
nand U364 (N_364,In_126,In_590);
or U365 (N_365,In_282,In_379);
or U366 (N_366,In_146,In_329);
or U367 (N_367,In_317,In_389);
nand U368 (N_368,In_86,In_159);
nor U369 (N_369,In_114,In_603);
nor U370 (N_370,In_363,In_280);
nor U371 (N_371,In_712,In_441);
and U372 (N_372,In_277,In_115);
nor U373 (N_373,In_312,In_491);
or U374 (N_374,In_531,In_601);
and U375 (N_375,In_353,In_698);
or U376 (N_376,In_44,In_573);
and U377 (N_377,In_81,In_87);
or U378 (N_378,In_56,In_188);
and U379 (N_379,In_627,In_143);
or U380 (N_380,In_23,In_340);
nand U381 (N_381,In_427,In_336);
nand U382 (N_382,In_566,In_457);
nor U383 (N_383,In_611,In_480);
and U384 (N_384,In_490,In_523);
nor U385 (N_385,In_483,In_723);
nand U386 (N_386,In_443,In_376);
nand U387 (N_387,In_348,In_243);
and U388 (N_388,In_43,In_504);
or U389 (N_389,In_56,In_730);
and U390 (N_390,In_249,In_388);
or U391 (N_391,In_495,In_478);
and U392 (N_392,In_282,In_622);
and U393 (N_393,In_485,In_691);
nand U394 (N_394,In_104,In_144);
nor U395 (N_395,In_179,In_225);
nor U396 (N_396,In_601,In_460);
and U397 (N_397,In_547,In_305);
or U398 (N_398,In_182,In_118);
nor U399 (N_399,In_51,In_136);
nor U400 (N_400,In_449,In_342);
and U401 (N_401,In_352,In_709);
nand U402 (N_402,In_603,In_594);
nand U403 (N_403,In_2,In_400);
nor U404 (N_404,In_667,In_76);
or U405 (N_405,In_622,In_479);
and U406 (N_406,In_688,In_11);
nor U407 (N_407,In_698,In_161);
nand U408 (N_408,In_356,In_238);
nand U409 (N_409,In_658,In_630);
nand U410 (N_410,In_325,In_563);
nand U411 (N_411,In_298,In_392);
or U412 (N_412,In_465,In_390);
and U413 (N_413,In_447,In_413);
or U414 (N_414,In_541,In_378);
or U415 (N_415,In_405,In_598);
nor U416 (N_416,In_734,In_718);
nand U417 (N_417,In_372,In_560);
or U418 (N_418,In_601,In_713);
or U419 (N_419,In_168,In_357);
or U420 (N_420,In_484,In_649);
nor U421 (N_421,In_556,In_244);
nor U422 (N_422,In_693,In_84);
or U423 (N_423,In_632,In_469);
or U424 (N_424,In_191,In_274);
nand U425 (N_425,In_701,In_78);
nor U426 (N_426,In_264,In_506);
or U427 (N_427,In_385,In_500);
nor U428 (N_428,In_145,In_363);
nor U429 (N_429,In_541,In_232);
nor U430 (N_430,In_588,In_518);
and U431 (N_431,In_691,In_138);
nand U432 (N_432,In_429,In_113);
nor U433 (N_433,In_366,In_353);
or U434 (N_434,In_142,In_384);
nand U435 (N_435,In_240,In_206);
nand U436 (N_436,In_557,In_693);
nor U437 (N_437,In_87,In_49);
or U438 (N_438,In_389,In_716);
nor U439 (N_439,In_131,In_510);
nor U440 (N_440,In_562,In_533);
nor U441 (N_441,In_298,In_464);
or U442 (N_442,In_740,In_435);
or U443 (N_443,In_284,In_308);
nor U444 (N_444,In_739,In_137);
xnor U445 (N_445,In_359,In_320);
nor U446 (N_446,In_218,In_417);
nand U447 (N_447,In_264,In_156);
and U448 (N_448,In_326,In_705);
nor U449 (N_449,In_644,In_297);
nor U450 (N_450,In_665,In_556);
nand U451 (N_451,In_309,In_721);
nand U452 (N_452,In_204,In_457);
and U453 (N_453,In_663,In_355);
or U454 (N_454,In_741,In_195);
nor U455 (N_455,In_276,In_363);
nand U456 (N_456,In_231,In_473);
nand U457 (N_457,In_173,In_262);
and U458 (N_458,In_10,In_598);
or U459 (N_459,In_88,In_399);
nand U460 (N_460,In_449,In_520);
or U461 (N_461,In_311,In_274);
nor U462 (N_462,In_515,In_719);
nor U463 (N_463,In_69,In_576);
or U464 (N_464,In_74,In_608);
xor U465 (N_465,In_545,In_748);
nand U466 (N_466,In_633,In_377);
nor U467 (N_467,In_230,In_584);
or U468 (N_468,In_600,In_592);
nand U469 (N_469,In_477,In_478);
or U470 (N_470,In_194,In_569);
and U471 (N_471,In_364,In_430);
nor U472 (N_472,In_503,In_676);
nand U473 (N_473,In_205,In_226);
or U474 (N_474,In_5,In_731);
nand U475 (N_475,In_566,In_365);
nand U476 (N_476,In_545,In_438);
nand U477 (N_477,In_4,In_145);
and U478 (N_478,In_265,In_727);
nor U479 (N_479,In_316,In_592);
and U480 (N_480,In_115,In_322);
and U481 (N_481,In_648,In_228);
nand U482 (N_482,In_309,In_98);
nand U483 (N_483,In_536,In_97);
nand U484 (N_484,In_419,In_369);
nor U485 (N_485,In_527,In_56);
and U486 (N_486,In_568,In_526);
or U487 (N_487,In_640,In_452);
nor U488 (N_488,In_414,In_163);
nand U489 (N_489,In_552,In_712);
or U490 (N_490,In_315,In_728);
nand U491 (N_491,In_60,In_257);
nand U492 (N_492,In_491,In_38);
nor U493 (N_493,In_289,In_472);
nor U494 (N_494,In_391,In_96);
or U495 (N_495,In_89,In_474);
or U496 (N_496,In_617,In_209);
and U497 (N_497,In_640,In_62);
nand U498 (N_498,In_628,In_484);
or U499 (N_499,In_657,In_178);
nand U500 (N_500,In_456,In_638);
nand U501 (N_501,In_185,In_243);
and U502 (N_502,In_447,In_192);
or U503 (N_503,In_439,In_468);
nand U504 (N_504,In_19,In_15);
or U505 (N_505,In_346,In_345);
and U506 (N_506,In_549,In_33);
nand U507 (N_507,In_121,In_691);
nand U508 (N_508,In_715,In_653);
nand U509 (N_509,In_500,In_710);
nor U510 (N_510,In_248,In_653);
nor U511 (N_511,In_176,In_528);
nor U512 (N_512,In_84,In_290);
and U513 (N_513,In_336,In_475);
nor U514 (N_514,In_581,In_69);
and U515 (N_515,In_597,In_414);
and U516 (N_516,In_675,In_25);
and U517 (N_517,In_725,In_138);
and U518 (N_518,In_91,In_523);
nand U519 (N_519,In_76,In_631);
nor U520 (N_520,In_467,In_670);
nor U521 (N_521,In_684,In_474);
or U522 (N_522,In_210,In_629);
nor U523 (N_523,In_635,In_561);
nand U524 (N_524,In_682,In_314);
or U525 (N_525,In_604,In_677);
and U526 (N_526,In_432,In_725);
nor U527 (N_527,In_131,In_155);
nand U528 (N_528,In_105,In_49);
and U529 (N_529,In_647,In_533);
nand U530 (N_530,In_746,In_717);
nor U531 (N_531,In_56,In_66);
nor U532 (N_532,In_143,In_492);
nor U533 (N_533,In_6,In_575);
or U534 (N_534,In_162,In_179);
or U535 (N_535,In_296,In_488);
or U536 (N_536,In_258,In_29);
nor U537 (N_537,In_384,In_114);
xnor U538 (N_538,In_365,In_563);
nand U539 (N_539,In_373,In_179);
xnor U540 (N_540,In_574,In_133);
and U541 (N_541,In_323,In_532);
or U542 (N_542,In_239,In_53);
or U543 (N_543,In_95,In_63);
or U544 (N_544,In_200,In_616);
and U545 (N_545,In_193,In_464);
or U546 (N_546,In_317,In_552);
or U547 (N_547,In_586,In_5);
or U548 (N_548,In_654,In_631);
nand U549 (N_549,In_736,In_178);
and U550 (N_550,In_63,In_606);
nor U551 (N_551,In_562,In_426);
nor U552 (N_552,In_69,In_299);
nor U553 (N_553,In_724,In_326);
and U554 (N_554,In_578,In_660);
nor U555 (N_555,In_216,In_159);
or U556 (N_556,In_298,In_570);
nand U557 (N_557,In_247,In_717);
or U558 (N_558,In_284,In_435);
xor U559 (N_559,In_720,In_599);
or U560 (N_560,In_296,In_732);
and U561 (N_561,In_579,In_166);
or U562 (N_562,In_688,In_63);
nor U563 (N_563,In_392,In_368);
or U564 (N_564,In_148,In_310);
and U565 (N_565,In_255,In_446);
and U566 (N_566,In_502,In_154);
nor U567 (N_567,In_411,In_549);
nor U568 (N_568,In_199,In_599);
and U569 (N_569,In_242,In_392);
nand U570 (N_570,In_247,In_359);
or U571 (N_571,In_51,In_484);
or U572 (N_572,In_721,In_164);
nand U573 (N_573,In_91,In_418);
nand U574 (N_574,In_514,In_107);
and U575 (N_575,In_196,In_651);
nor U576 (N_576,In_654,In_743);
or U577 (N_577,In_127,In_42);
nor U578 (N_578,In_329,In_642);
nor U579 (N_579,In_301,In_56);
nand U580 (N_580,In_480,In_40);
and U581 (N_581,In_455,In_656);
or U582 (N_582,In_1,In_651);
nand U583 (N_583,In_492,In_645);
nand U584 (N_584,In_491,In_64);
or U585 (N_585,In_182,In_134);
nor U586 (N_586,In_553,In_626);
nor U587 (N_587,In_613,In_469);
and U588 (N_588,In_278,In_347);
or U589 (N_589,In_367,In_551);
nand U590 (N_590,In_368,In_432);
nand U591 (N_591,In_656,In_347);
nand U592 (N_592,In_665,In_325);
and U593 (N_593,In_311,In_668);
or U594 (N_594,In_247,In_600);
or U595 (N_595,In_584,In_464);
or U596 (N_596,In_212,In_645);
and U597 (N_597,In_349,In_145);
nand U598 (N_598,In_637,In_211);
and U599 (N_599,In_36,In_60);
nand U600 (N_600,In_153,In_137);
and U601 (N_601,In_269,In_711);
and U602 (N_602,In_588,In_452);
and U603 (N_603,In_250,In_117);
nand U604 (N_604,In_684,In_122);
and U605 (N_605,In_475,In_579);
nor U606 (N_606,In_498,In_30);
nand U607 (N_607,In_562,In_400);
nand U608 (N_608,In_280,In_701);
nor U609 (N_609,In_413,In_568);
and U610 (N_610,In_249,In_106);
and U611 (N_611,In_413,In_238);
nor U612 (N_612,In_478,In_130);
and U613 (N_613,In_128,In_286);
or U614 (N_614,In_630,In_661);
and U615 (N_615,In_525,In_183);
nand U616 (N_616,In_104,In_244);
nor U617 (N_617,In_283,In_712);
nand U618 (N_618,In_398,In_84);
nor U619 (N_619,In_84,In_296);
or U620 (N_620,In_68,In_717);
nor U621 (N_621,In_465,In_200);
nand U622 (N_622,In_507,In_461);
or U623 (N_623,In_676,In_660);
nor U624 (N_624,In_481,In_549);
and U625 (N_625,In_260,In_228);
or U626 (N_626,In_716,In_256);
nor U627 (N_627,In_408,In_276);
nand U628 (N_628,In_521,In_488);
nand U629 (N_629,In_368,In_55);
nor U630 (N_630,In_438,In_144);
nand U631 (N_631,In_80,In_268);
nor U632 (N_632,In_416,In_253);
nor U633 (N_633,In_432,In_207);
nand U634 (N_634,In_440,In_697);
nand U635 (N_635,In_100,In_433);
or U636 (N_636,In_203,In_573);
and U637 (N_637,In_509,In_630);
and U638 (N_638,In_12,In_606);
nor U639 (N_639,In_206,In_632);
nand U640 (N_640,In_80,In_11);
nand U641 (N_641,In_597,In_722);
nand U642 (N_642,In_576,In_595);
xor U643 (N_643,In_541,In_594);
nand U644 (N_644,In_704,In_385);
and U645 (N_645,In_280,In_29);
nand U646 (N_646,In_712,In_26);
and U647 (N_647,In_630,In_671);
nand U648 (N_648,In_151,In_404);
or U649 (N_649,In_354,In_459);
or U650 (N_650,In_279,In_200);
nor U651 (N_651,In_202,In_583);
nor U652 (N_652,In_491,In_298);
or U653 (N_653,In_555,In_564);
nor U654 (N_654,In_335,In_21);
and U655 (N_655,In_180,In_85);
nor U656 (N_656,In_291,In_1);
or U657 (N_657,In_653,In_719);
and U658 (N_658,In_418,In_656);
and U659 (N_659,In_144,In_279);
or U660 (N_660,In_422,In_11);
nand U661 (N_661,In_531,In_108);
nand U662 (N_662,In_238,In_409);
or U663 (N_663,In_129,In_614);
or U664 (N_664,In_598,In_713);
nor U665 (N_665,In_137,In_31);
nand U666 (N_666,In_576,In_457);
nand U667 (N_667,In_347,In_648);
nor U668 (N_668,In_36,In_377);
nor U669 (N_669,In_591,In_164);
and U670 (N_670,In_616,In_7);
and U671 (N_671,In_350,In_439);
nand U672 (N_672,In_400,In_154);
and U673 (N_673,In_20,In_330);
nor U674 (N_674,In_162,In_135);
and U675 (N_675,In_341,In_264);
or U676 (N_676,In_653,In_521);
nand U677 (N_677,In_412,In_655);
and U678 (N_678,In_55,In_619);
and U679 (N_679,In_540,In_252);
and U680 (N_680,In_562,In_93);
nor U681 (N_681,In_351,In_724);
nor U682 (N_682,In_304,In_424);
xor U683 (N_683,In_590,In_556);
nor U684 (N_684,In_506,In_193);
nand U685 (N_685,In_682,In_706);
nand U686 (N_686,In_598,In_215);
nand U687 (N_687,In_557,In_154);
nor U688 (N_688,In_696,In_731);
or U689 (N_689,In_287,In_422);
nand U690 (N_690,In_246,In_601);
and U691 (N_691,In_579,In_528);
and U692 (N_692,In_367,In_276);
nand U693 (N_693,In_622,In_48);
nor U694 (N_694,In_21,In_643);
or U695 (N_695,In_409,In_437);
nand U696 (N_696,In_553,In_709);
nor U697 (N_697,In_478,In_156);
or U698 (N_698,In_470,In_511);
nor U699 (N_699,In_453,In_524);
nor U700 (N_700,In_280,In_313);
nand U701 (N_701,In_460,In_715);
nand U702 (N_702,In_31,In_436);
or U703 (N_703,In_141,In_701);
nor U704 (N_704,In_233,In_470);
or U705 (N_705,In_77,In_136);
or U706 (N_706,In_3,In_710);
nand U707 (N_707,In_570,In_379);
nand U708 (N_708,In_210,In_521);
nand U709 (N_709,In_315,In_292);
and U710 (N_710,In_517,In_514);
and U711 (N_711,In_469,In_16);
or U712 (N_712,In_77,In_441);
or U713 (N_713,In_431,In_401);
and U714 (N_714,In_319,In_535);
and U715 (N_715,In_493,In_264);
and U716 (N_716,In_660,In_621);
nand U717 (N_717,In_241,In_398);
nand U718 (N_718,In_286,In_445);
nor U719 (N_719,In_626,In_8);
and U720 (N_720,In_744,In_230);
or U721 (N_721,In_652,In_418);
or U722 (N_722,In_329,In_456);
and U723 (N_723,In_34,In_77);
nand U724 (N_724,In_574,In_421);
nand U725 (N_725,In_81,In_655);
or U726 (N_726,In_124,In_120);
nor U727 (N_727,In_681,In_371);
or U728 (N_728,In_164,In_391);
nand U729 (N_729,In_615,In_503);
and U730 (N_730,In_607,In_550);
or U731 (N_731,In_382,In_101);
nor U732 (N_732,In_320,In_411);
nand U733 (N_733,In_535,In_177);
or U734 (N_734,In_441,In_103);
and U735 (N_735,In_92,In_222);
nand U736 (N_736,In_105,In_119);
nand U737 (N_737,In_525,In_456);
or U738 (N_738,In_0,In_543);
nand U739 (N_739,In_504,In_352);
nand U740 (N_740,In_128,In_476);
nor U741 (N_741,In_383,In_72);
xor U742 (N_742,In_28,In_459);
or U743 (N_743,In_103,In_294);
nand U744 (N_744,In_379,In_515);
nor U745 (N_745,In_312,In_45);
or U746 (N_746,In_564,In_172);
nor U747 (N_747,In_747,In_361);
nor U748 (N_748,In_544,In_86);
or U749 (N_749,In_510,In_514);
or U750 (N_750,In_506,In_424);
and U751 (N_751,In_143,In_736);
or U752 (N_752,In_458,In_717);
or U753 (N_753,In_235,In_460);
nor U754 (N_754,In_77,In_226);
nor U755 (N_755,In_433,In_167);
nor U756 (N_756,In_567,In_514);
and U757 (N_757,In_231,In_151);
or U758 (N_758,In_483,In_243);
nor U759 (N_759,In_528,In_181);
and U760 (N_760,In_486,In_496);
or U761 (N_761,In_342,In_695);
nor U762 (N_762,In_568,In_675);
or U763 (N_763,In_293,In_709);
nor U764 (N_764,In_356,In_2);
nand U765 (N_765,In_121,In_175);
nand U766 (N_766,In_81,In_742);
or U767 (N_767,In_421,In_236);
nand U768 (N_768,In_24,In_348);
or U769 (N_769,In_693,In_396);
or U770 (N_770,In_58,In_498);
and U771 (N_771,In_687,In_402);
or U772 (N_772,In_161,In_467);
nand U773 (N_773,In_205,In_736);
or U774 (N_774,In_453,In_185);
or U775 (N_775,In_110,In_352);
and U776 (N_776,In_502,In_697);
or U777 (N_777,In_187,In_711);
or U778 (N_778,In_149,In_228);
or U779 (N_779,In_602,In_167);
nor U780 (N_780,In_127,In_70);
or U781 (N_781,In_538,In_552);
xor U782 (N_782,In_69,In_409);
nor U783 (N_783,In_73,In_149);
nor U784 (N_784,In_49,In_473);
nand U785 (N_785,In_191,In_294);
and U786 (N_786,In_737,In_268);
nand U787 (N_787,In_502,In_661);
or U788 (N_788,In_747,In_709);
and U789 (N_789,In_572,In_625);
nand U790 (N_790,In_650,In_507);
and U791 (N_791,In_598,In_521);
nand U792 (N_792,In_327,In_572);
nand U793 (N_793,In_609,In_201);
and U794 (N_794,In_169,In_328);
and U795 (N_795,In_200,In_543);
nand U796 (N_796,In_66,In_611);
or U797 (N_797,In_221,In_600);
nand U798 (N_798,In_447,In_269);
or U799 (N_799,In_639,In_280);
or U800 (N_800,In_502,In_642);
nor U801 (N_801,In_300,In_439);
nand U802 (N_802,In_652,In_37);
or U803 (N_803,In_545,In_377);
and U804 (N_804,In_600,In_187);
and U805 (N_805,In_633,In_144);
or U806 (N_806,In_549,In_659);
and U807 (N_807,In_608,In_529);
nor U808 (N_808,In_472,In_684);
or U809 (N_809,In_291,In_308);
nand U810 (N_810,In_256,In_116);
or U811 (N_811,In_596,In_339);
and U812 (N_812,In_123,In_376);
nand U813 (N_813,In_481,In_676);
nand U814 (N_814,In_422,In_262);
nor U815 (N_815,In_347,In_688);
and U816 (N_816,In_490,In_615);
nand U817 (N_817,In_77,In_537);
nor U818 (N_818,In_433,In_208);
nand U819 (N_819,In_332,In_508);
and U820 (N_820,In_650,In_304);
nand U821 (N_821,In_358,In_65);
nand U822 (N_822,In_715,In_159);
or U823 (N_823,In_555,In_429);
nand U824 (N_824,In_125,In_608);
nand U825 (N_825,In_311,In_152);
nand U826 (N_826,In_558,In_183);
nand U827 (N_827,In_442,In_125);
nand U828 (N_828,In_168,In_741);
nand U829 (N_829,In_329,In_108);
nand U830 (N_830,In_21,In_184);
or U831 (N_831,In_655,In_563);
nor U832 (N_832,In_334,In_443);
or U833 (N_833,In_446,In_283);
nor U834 (N_834,In_288,In_575);
or U835 (N_835,In_74,In_524);
nand U836 (N_836,In_632,In_616);
and U837 (N_837,In_459,In_694);
nand U838 (N_838,In_299,In_617);
or U839 (N_839,In_507,In_355);
nor U840 (N_840,In_563,In_302);
nor U841 (N_841,In_62,In_405);
and U842 (N_842,In_483,In_402);
nand U843 (N_843,In_243,In_269);
or U844 (N_844,In_336,In_170);
and U845 (N_845,In_578,In_282);
nor U846 (N_846,In_726,In_52);
or U847 (N_847,In_176,In_646);
or U848 (N_848,In_513,In_620);
nand U849 (N_849,In_347,In_493);
and U850 (N_850,In_466,In_435);
nor U851 (N_851,In_537,In_389);
nand U852 (N_852,In_467,In_104);
or U853 (N_853,In_3,In_89);
nand U854 (N_854,In_17,In_166);
nand U855 (N_855,In_302,In_492);
or U856 (N_856,In_266,In_578);
nor U857 (N_857,In_495,In_309);
or U858 (N_858,In_642,In_364);
and U859 (N_859,In_236,In_570);
or U860 (N_860,In_286,In_547);
nand U861 (N_861,In_182,In_587);
nor U862 (N_862,In_361,In_666);
or U863 (N_863,In_94,In_256);
and U864 (N_864,In_389,In_698);
nand U865 (N_865,In_287,In_646);
or U866 (N_866,In_539,In_54);
or U867 (N_867,In_495,In_589);
nand U868 (N_868,In_686,In_731);
or U869 (N_869,In_492,In_458);
and U870 (N_870,In_640,In_241);
nor U871 (N_871,In_682,In_211);
nand U872 (N_872,In_345,In_719);
nand U873 (N_873,In_377,In_157);
nor U874 (N_874,In_481,In_125);
nor U875 (N_875,In_31,In_682);
nor U876 (N_876,In_169,In_360);
nand U877 (N_877,In_267,In_33);
nor U878 (N_878,In_378,In_253);
nor U879 (N_879,In_652,In_546);
nor U880 (N_880,In_717,In_461);
nand U881 (N_881,In_479,In_550);
nand U882 (N_882,In_6,In_600);
or U883 (N_883,In_588,In_399);
and U884 (N_884,In_231,In_548);
and U885 (N_885,In_688,In_720);
and U886 (N_886,In_646,In_676);
nor U887 (N_887,In_713,In_36);
and U888 (N_888,In_125,In_354);
nand U889 (N_889,In_87,In_477);
nor U890 (N_890,In_394,In_627);
and U891 (N_891,In_142,In_44);
nor U892 (N_892,In_501,In_663);
xor U893 (N_893,In_398,In_535);
nor U894 (N_894,In_469,In_136);
nand U895 (N_895,In_656,In_500);
or U896 (N_896,In_660,In_642);
nand U897 (N_897,In_293,In_741);
nand U898 (N_898,In_158,In_57);
nor U899 (N_899,In_68,In_571);
or U900 (N_900,In_518,In_28);
nor U901 (N_901,In_371,In_158);
or U902 (N_902,In_729,In_404);
or U903 (N_903,In_726,In_181);
nor U904 (N_904,In_40,In_216);
and U905 (N_905,In_732,In_289);
or U906 (N_906,In_702,In_289);
or U907 (N_907,In_562,In_627);
nor U908 (N_908,In_640,In_54);
and U909 (N_909,In_599,In_175);
or U910 (N_910,In_470,In_735);
or U911 (N_911,In_453,In_342);
nand U912 (N_912,In_711,In_383);
nand U913 (N_913,In_351,In_137);
nor U914 (N_914,In_451,In_668);
and U915 (N_915,In_180,In_668);
and U916 (N_916,In_337,In_646);
and U917 (N_917,In_732,In_680);
and U918 (N_918,In_358,In_50);
nor U919 (N_919,In_136,In_361);
nand U920 (N_920,In_83,In_310);
nor U921 (N_921,In_155,In_388);
or U922 (N_922,In_441,In_620);
nand U923 (N_923,In_282,In_225);
or U924 (N_924,In_231,In_626);
nor U925 (N_925,In_85,In_657);
or U926 (N_926,In_137,In_532);
and U927 (N_927,In_445,In_335);
nor U928 (N_928,In_405,In_537);
and U929 (N_929,In_436,In_5);
and U930 (N_930,In_452,In_540);
and U931 (N_931,In_514,In_286);
nand U932 (N_932,In_593,In_556);
and U933 (N_933,In_215,In_477);
and U934 (N_934,In_204,In_235);
nor U935 (N_935,In_580,In_168);
nand U936 (N_936,In_406,In_52);
or U937 (N_937,In_142,In_439);
nor U938 (N_938,In_744,In_476);
and U939 (N_939,In_422,In_335);
nand U940 (N_940,In_156,In_425);
nor U941 (N_941,In_668,In_606);
or U942 (N_942,In_317,In_295);
nor U943 (N_943,In_583,In_228);
nand U944 (N_944,In_284,In_579);
nor U945 (N_945,In_420,In_484);
nand U946 (N_946,In_253,In_656);
and U947 (N_947,In_422,In_503);
nand U948 (N_948,In_36,In_167);
nor U949 (N_949,In_36,In_678);
nor U950 (N_950,In_665,In_609);
nand U951 (N_951,In_329,In_475);
and U952 (N_952,In_673,In_448);
and U953 (N_953,In_68,In_568);
nand U954 (N_954,In_489,In_249);
nand U955 (N_955,In_174,In_618);
nor U956 (N_956,In_324,In_572);
nor U957 (N_957,In_48,In_522);
nand U958 (N_958,In_297,In_110);
nor U959 (N_959,In_389,In_308);
nand U960 (N_960,In_440,In_356);
nor U961 (N_961,In_466,In_6);
nand U962 (N_962,In_631,In_688);
or U963 (N_963,In_464,In_328);
nor U964 (N_964,In_327,In_636);
nand U965 (N_965,In_489,In_124);
and U966 (N_966,In_636,In_278);
nand U967 (N_967,In_130,In_1);
nor U968 (N_968,In_222,In_52);
or U969 (N_969,In_378,In_551);
nor U970 (N_970,In_152,In_54);
and U971 (N_971,In_434,In_356);
nor U972 (N_972,In_8,In_576);
and U973 (N_973,In_512,In_235);
nand U974 (N_974,In_731,In_156);
nand U975 (N_975,In_506,In_705);
nand U976 (N_976,In_400,In_94);
and U977 (N_977,In_626,In_68);
and U978 (N_978,In_29,In_230);
and U979 (N_979,In_106,In_520);
nand U980 (N_980,In_422,In_175);
and U981 (N_981,In_636,In_569);
nor U982 (N_982,In_223,In_116);
or U983 (N_983,In_528,In_272);
and U984 (N_984,In_84,In_313);
and U985 (N_985,In_113,In_28);
nor U986 (N_986,In_501,In_740);
nor U987 (N_987,In_160,In_183);
nand U988 (N_988,In_461,In_561);
nor U989 (N_989,In_444,In_251);
nor U990 (N_990,In_72,In_675);
and U991 (N_991,In_494,In_712);
or U992 (N_992,In_295,In_151);
or U993 (N_993,In_732,In_324);
nand U994 (N_994,In_607,In_256);
or U995 (N_995,In_499,In_239);
nand U996 (N_996,In_155,In_298);
nand U997 (N_997,In_597,In_738);
or U998 (N_998,In_383,In_55);
nor U999 (N_999,In_538,In_642);
nand U1000 (N_1000,N_326,N_583);
and U1001 (N_1001,N_467,N_417);
nand U1002 (N_1002,N_157,N_948);
nor U1003 (N_1003,N_932,N_660);
nor U1004 (N_1004,N_77,N_139);
xnor U1005 (N_1005,N_974,N_679);
nand U1006 (N_1006,N_671,N_686);
nor U1007 (N_1007,N_711,N_20);
nand U1008 (N_1008,N_296,N_619);
nor U1009 (N_1009,N_60,N_668);
nand U1010 (N_1010,N_859,N_167);
nor U1011 (N_1011,N_726,N_198);
nand U1012 (N_1012,N_216,N_897);
and U1013 (N_1013,N_873,N_485);
nor U1014 (N_1014,N_757,N_881);
nor U1015 (N_1015,N_913,N_165);
xnor U1016 (N_1016,N_459,N_779);
nand U1017 (N_1017,N_43,N_407);
nand U1018 (N_1018,N_237,N_310);
and U1019 (N_1019,N_273,N_602);
and U1020 (N_1020,N_240,N_737);
nor U1021 (N_1021,N_155,N_458);
nor U1022 (N_1022,N_82,N_730);
and U1023 (N_1023,N_276,N_341);
nand U1024 (N_1024,N_521,N_518);
and U1025 (N_1025,N_76,N_205);
nor U1026 (N_1026,N_256,N_912);
nand U1027 (N_1027,N_338,N_742);
nand U1028 (N_1028,N_93,N_332);
or U1029 (N_1029,N_851,N_741);
nor U1030 (N_1030,N_836,N_911);
nor U1031 (N_1031,N_158,N_69);
and U1032 (N_1032,N_544,N_937);
and U1033 (N_1033,N_150,N_192);
nand U1034 (N_1034,N_65,N_784);
and U1035 (N_1035,N_768,N_705);
nand U1036 (N_1036,N_294,N_747);
nand U1037 (N_1037,N_123,N_795);
nand U1038 (N_1038,N_412,N_709);
nand U1039 (N_1039,N_370,N_56);
nand U1040 (N_1040,N_290,N_342);
nand U1041 (N_1041,N_390,N_439);
nand U1042 (N_1042,N_535,N_207);
and U1043 (N_1043,N_440,N_788);
nor U1044 (N_1044,N_415,N_499);
or U1045 (N_1045,N_110,N_526);
or U1046 (N_1046,N_70,N_218);
and U1047 (N_1047,N_409,N_917);
nand U1048 (N_1048,N_21,N_186);
nor U1049 (N_1049,N_680,N_542);
nor U1050 (N_1050,N_11,N_166);
xnor U1051 (N_1051,N_66,N_532);
and U1052 (N_1052,N_714,N_80);
or U1053 (N_1053,N_630,N_580);
nor U1054 (N_1054,N_272,N_608);
nand U1055 (N_1055,N_41,N_321);
and U1056 (N_1056,N_175,N_945);
nor U1057 (N_1057,N_793,N_72);
and U1058 (N_1058,N_772,N_177);
and U1059 (N_1059,N_129,N_212);
and U1060 (N_1060,N_57,N_910);
or U1061 (N_1061,N_364,N_946);
and U1062 (N_1062,N_716,N_403);
or U1063 (N_1063,N_410,N_696);
or U1064 (N_1064,N_10,N_830);
or U1065 (N_1065,N_646,N_694);
nand U1066 (N_1066,N_1,N_800);
and U1067 (N_1067,N_581,N_151);
nand U1068 (N_1068,N_187,N_664);
or U1069 (N_1069,N_960,N_547);
nand U1070 (N_1070,N_37,N_810);
and U1071 (N_1071,N_239,N_40);
nand U1072 (N_1072,N_445,N_801);
or U1073 (N_1073,N_840,N_433);
and U1074 (N_1074,N_796,N_427);
nand U1075 (N_1075,N_394,N_847);
or U1076 (N_1076,N_63,N_24);
nand U1077 (N_1077,N_325,N_402);
and U1078 (N_1078,N_260,N_598);
and U1079 (N_1079,N_924,N_670);
nor U1080 (N_1080,N_751,N_429);
and U1081 (N_1081,N_822,N_382);
or U1082 (N_1082,N_791,N_6);
or U1083 (N_1083,N_597,N_49);
nand U1084 (N_1084,N_414,N_301);
or U1085 (N_1085,N_416,N_323);
nor U1086 (N_1086,N_389,N_564);
nor U1087 (N_1087,N_700,N_968);
and U1088 (N_1088,N_100,N_484);
nand U1089 (N_1089,N_718,N_208);
and U1090 (N_1090,N_826,N_928);
nand U1091 (N_1091,N_54,N_963);
or U1092 (N_1092,N_343,N_510);
nand U1093 (N_1093,N_136,N_969);
nor U1094 (N_1094,N_657,N_566);
and U1095 (N_1095,N_504,N_233);
nor U1096 (N_1096,N_536,N_42);
nor U1097 (N_1097,N_87,N_819);
and U1098 (N_1098,N_367,N_661);
or U1099 (N_1099,N_669,N_586);
nor U1100 (N_1100,N_620,N_243);
nand U1101 (N_1101,N_617,N_935);
nand U1102 (N_1102,N_629,N_677);
or U1103 (N_1103,N_380,N_555);
nand U1104 (N_1104,N_965,N_610);
nand U1105 (N_1105,N_302,N_854);
and U1106 (N_1106,N_713,N_16);
nor U1107 (N_1107,N_644,N_875);
nand U1108 (N_1108,N_97,N_456);
or U1109 (N_1109,N_393,N_199);
and U1110 (N_1110,N_856,N_430);
nand U1111 (N_1111,N_271,N_31);
nand U1112 (N_1112,N_297,N_340);
or U1113 (N_1113,N_571,N_156);
nor U1114 (N_1114,N_247,N_446);
and U1115 (N_1115,N_865,N_319);
and U1116 (N_1116,N_920,N_210);
nand U1117 (N_1117,N_453,N_170);
or U1118 (N_1118,N_786,N_162);
nor U1119 (N_1119,N_373,N_512);
nand U1120 (N_1120,N_607,N_314);
and U1121 (N_1121,N_584,N_251);
nand U1122 (N_1122,N_47,N_143);
nor U1123 (N_1123,N_463,N_209);
nand U1124 (N_1124,N_211,N_611);
or U1125 (N_1125,N_493,N_435);
and U1126 (N_1126,N_352,N_88);
or U1127 (N_1127,N_64,N_944);
nand U1128 (N_1128,N_33,N_426);
and U1129 (N_1129,N_995,N_472);
or U1130 (N_1130,N_196,N_188);
and U1131 (N_1131,N_73,N_213);
nor U1132 (N_1132,N_889,N_137);
and U1133 (N_1133,N_992,N_245);
or U1134 (N_1134,N_725,N_940);
and U1135 (N_1135,N_519,N_75);
and U1136 (N_1136,N_448,N_823);
nor U1137 (N_1137,N_874,N_640);
nand U1138 (N_1138,N_490,N_503);
or U1139 (N_1139,N_400,N_558);
nand U1140 (N_1140,N_527,N_220);
nor U1141 (N_1141,N_587,N_180);
or U1142 (N_1142,N_295,N_281);
nor U1143 (N_1143,N_612,N_766);
or U1144 (N_1144,N_534,N_293);
nand U1145 (N_1145,N_565,N_386);
nor U1146 (N_1146,N_728,N_720);
or U1147 (N_1147,N_591,N_746);
or U1148 (N_1148,N_219,N_684);
nand U1149 (N_1149,N_486,N_891);
nor U1150 (N_1150,N_770,N_86);
and U1151 (N_1151,N_886,N_357);
and U1152 (N_1152,N_857,N_45);
nand U1153 (N_1153,N_999,N_13);
and U1154 (N_1154,N_561,N_594);
or U1155 (N_1155,N_114,N_698);
nor U1156 (N_1156,N_471,N_708);
nor U1157 (N_1157,N_717,N_805);
nand U1158 (N_1158,N_572,N_933);
and U1159 (N_1159,N_115,N_998);
and U1160 (N_1160,N_579,N_515);
or U1161 (N_1161,N_487,N_539);
nand U1162 (N_1162,N_809,N_821);
or U1163 (N_1163,N_52,N_773);
nor U1164 (N_1164,N_868,N_756);
nand U1165 (N_1165,N_553,N_74);
nor U1166 (N_1166,N_596,N_530);
or U1167 (N_1167,N_739,N_906);
nor U1168 (N_1168,N_287,N_743);
nor U1169 (N_1169,N_91,N_622);
nor U1170 (N_1170,N_799,N_614);
nor U1171 (N_1171,N_349,N_436);
or U1172 (N_1172,N_964,N_627);
and U1173 (N_1173,N_423,N_844);
nand U1174 (N_1174,N_108,N_880);
nor U1175 (N_1175,N_22,N_329);
xnor U1176 (N_1176,N_588,N_953);
nor U1177 (N_1177,N_852,N_653);
nand U1178 (N_1178,N_624,N_548);
nand U1179 (N_1179,N_284,N_29);
and U1180 (N_1180,N_523,N_447);
xnor U1181 (N_1181,N_385,N_185);
or U1182 (N_1182,N_226,N_263);
nand U1183 (N_1183,N_887,N_904);
and U1184 (N_1184,N_28,N_422);
or U1185 (N_1185,N_674,N_497);
or U1186 (N_1186,N_921,N_438);
nand U1187 (N_1187,N_3,N_862);
nor U1188 (N_1188,N_505,N_330);
and U1189 (N_1189,N_842,N_817);
nand U1190 (N_1190,N_78,N_853);
or U1191 (N_1191,N_25,N_984);
and U1192 (N_1192,N_182,N_101);
nor U1193 (N_1193,N_549,N_864);
and U1194 (N_1194,N_238,N_976);
or U1195 (N_1195,N_845,N_356);
nor U1196 (N_1196,N_763,N_981);
nand U1197 (N_1197,N_59,N_543);
and U1198 (N_1198,N_361,N_815);
nand U1199 (N_1199,N_996,N_383);
and U1200 (N_1200,N_126,N_280);
nor U1201 (N_1201,N_408,N_424);
nand U1202 (N_1202,N_153,N_916);
nor U1203 (N_1203,N_592,N_971);
and U1204 (N_1204,N_923,N_362);
nor U1205 (N_1205,N_601,N_970);
nor U1206 (N_1206,N_303,N_79);
and U1207 (N_1207,N_236,N_480);
nor U1208 (N_1208,N_368,N_520);
nand U1209 (N_1209,N_344,N_152);
and U1210 (N_1210,N_305,N_811);
xnor U1211 (N_1211,N_222,N_972);
nand U1212 (N_1212,N_178,N_589);
and U1213 (N_1213,N_837,N_687);
nor U1214 (N_1214,N_681,N_89);
nor U1215 (N_1215,N_81,N_395);
or U1216 (N_1216,N_161,N_533);
and U1217 (N_1217,N_355,N_632);
or U1218 (N_1218,N_197,N_599);
nor U1219 (N_1219,N_789,N_869);
nand U1220 (N_1220,N_899,N_7);
and U1221 (N_1221,N_384,N_313);
nand U1222 (N_1222,N_248,N_903);
and U1223 (N_1223,N_255,N_203);
or U1224 (N_1224,N_306,N_160);
and U1225 (N_1225,N_292,N_229);
nand U1226 (N_1226,N_466,N_979);
nor U1227 (N_1227,N_846,N_217);
nand U1228 (N_1228,N_437,N_164);
or U1229 (N_1229,N_973,N_298);
or U1230 (N_1230,N_360,N_790);
and U1231 (N_1231,N_537,N_849);
and U1232 (N_1232,N_744,N_418);
and U1233 (N_1233,N_442,N_637);
nor U1234 (N_1234,N_309,N_39);
or U1235 (N_1235,N_96,N_254);
nor U1236 (N_1236,N_154,N_922);
and U1237 (N_1237,N_328,N_26);
or U1238 (N_1238,N_347,N_107);
and U1239 (N_1239,N_991,N_32);
nand U1240 (N_1240,N_371,N_605);
or U1241 (N_1241,N_753,N_896);
nor U1242 (N_1242,N_501,N_246);
or U1243 (N_1243,N_939,N_122);
and U1244 (N_1244,N_189,N_813);
nor U1245 (N_1245,N_618,N_884);
or U1246 (N_1246,N_324,N_118);
nand U1247 (N_1247,N_633,N_378);
xor U1248 (N_1248,N_638,N_643);
nor U1249 (N_1249,N_17,N_712);
nand U1250 (N_1250,N_265,N_787);
xor U1251 (N_1251,N_270,N_376);
and U1252 (N_1252,N_975,N_759);
and U1253 (N_1253,N_812,N_914);
or U1254 (N_1254,N_682,N_898);
or U1255 (N_1255,N_483,N_958);
nor U1256 (N_1256,N_365,N_286);
nand U1257 (N_1257,N_102,N_522);
or U1258 (N_1258,N_194,N_715);
or U1259 (N_1259,N_655,N_659);
and U1260 (N_1260,N_574,N_431);
nand U1261 (N_1261,N_0,N_835);
nor U1262 (N_1262,N_761,N_142);
and U1263 (N_1263,N_421,N_333);
nor U1264 (N_1264,N_145,N_289);
or U1265 (N_1265,N_44,N_2);
nor U1266 (N_1266,N_806,N_559);
nand U1267 (N_1267,N_235,N_545);
nor U1268 (N_1268,N_274,N_702);
nand U1269 (N_1269,N_938,N_802);
nor U1270 (N_1270,N_710,N_117);
nand U1271 (N_1271,N_754,N_513);
nand U1272 (N_1272,N_375,N_782);
or U1273 (N_1273,N_264,N_749);
and U1274 (N_1274,N_244,N_762);
nand U1275 (N_1275,N_936,N_267);
nor U1276 (N_1276,N_697,N_92);
nand U1277 (N_1277,N_650,N_475);
and U1278 (N_1278,N_954,N_401);
nand U1279 (N_1279,N_441,N_279);
nand U1280 (N_1280,N_103,N_541);
nor U1281 (N_1281,N_652,N_168);
nand U1282 (N_1282,N_259,N_308);
and U1283 (N_1283,N_363,N_723);
or U1284 (N_1284,N_146,N_269);
nor U1285 (N_1285,N_890,N_867);
nand U1286 (N_1286,N_311,N_36);
and U1287 (N_1287,N_734,N_95);
or U1288 (N_1288,N_691,N_200);
nor U1289 (N_1289,N_183,N_201);
nor U1290 (N_1290,N_516,N_832);
nor U1291 (N_1291,N_955,N_993);
nand U1292 (N_1292,N_531,N_777);
and U1293 (N_1293,N_818,N_977);
nand U1294 (N_1294,N_870,N_635);
or U1295 (N_1295,N_464,N_647);
nor U1296 (N_1296,N_797,N_927);
nor U1297 (N_1297,N_252,N_125);
or U1298 (N_1298,N_174,N_135);
and U1299 (N_1299,N_595,N_962);
nor U1300 (N_1300,N_663,N_651);
or U1301 (N_1301,N_420,N_227);
nor U1302 (N_1302,N_508,N_808);
and U1303 (N_1303,N_481,N_514);
nor U1304 (N_1304,N_834,N_642);
nor U1305 (N_1305,N_479,N_369);
or U1306 (N_1306,N_299,N_358);
or U1307 (N_1307,N_404,N_735);
or U1308 (N_1308,N_397,N_951);
nor U1309 (N_1309,N_132,N_179);
or U1310 (N_1310,N_989,N_570);
and U1311 (N_1311,N_335,N_947);
nor U1312 (N_1312,N_434,N_562);
or U1313 (N_1313,N_625,N_133);
or U1314 (N_1314,N_320,N_858);
nand U1315 (N_1315,N_98,N_727);
nand U1316 (N_1316,N_606,N_477);
or U1317 (N_1317,N_454,N_752);
and U1318 (N_1318,N_517,N_474);
or U1319 (N_1319,N_672,N_473);
or U1320 (N_1320,N_528,N_68);
nand U1321 (N_1321,N_334,N_55);
nor U1322 (N_1322,N_931,N_345);
nor U1323 (N_1323,N_764,N_169);
nor U1324 (N_1324,N_231,N_171);
nand U1325 (N_1325,N_776,N_814);
nand U1326 (N_1326,N_656,N_695);
and U1327 (N_1327,N_172,N_492);
nand U1328 (N_1328,N_678,N_683);
and U1329 (N_1329,N_980,N_860);
nand U1330 (N_1330,N_5,N_994);
and U1331 (N_1331,N_90,N_816);
nor U1332 (N_1332,N_224,N_736);
or U1333 (N_1333,N_144,N_673);
nor U1334 (N_1334,N_51,N_824);
nand U1335 (N_1335,N_148,N_99);
and U1336 (N_1336,N_491,N_291);
and U1337 (N_1337,N_496,N_755);
nor U1338 (N_1338,N_892,N_506);
nand U1339 (N_1339,N_841,N_988);
nor U1340 (N_1340,N_949,N_950);
and U1341 (N_1341,N_590,N_740);
or U1342 (N_1342,N_925,N_722);
and U1343 (N_1343,N_387,N_379);
and U1344 (N_1344,N_419,N_266);
or U1345 (N_1345,N_374,N_658);
and U1346 (N_1346,N_745,N_621);
nand U1347 (N_1347,N_825,N_985);
nor U1348 (N_1348,N_879,N_190);
or U1349 (N_1349,N_557,N_649);
and U1350 (N_1350,N_285,N_894);
and U1351 (N_1351,N_234,N_568);
and U1352 (N_1352,N_4,N_760);
and U1353 (N_1353,N_62,N_71);
nand U1354 (N_1354,N_863,N_27);
nor U1355 (N_1355,N_468,N_885);
or U1356 (N_1356,N_413,N_915);
nand U1357 (N_1357,N_986,N_907);
nand U1358 (N_1358,N_83,N_675);
or U1359 (N_1359,N_214,N_443);
or U1360 (N_1360,N_609,N_769);
nand U1361 (N_1361,N_366,N_843);
nand U1362 (N_1362,N_8,N_104);
nand U1363 (N_1363,N_317,N_478);
nand U1364 (N_1364,N_253,N_469);
or U1365 (N_1365,N_631,N_893);
nor U1366 (N_1366,N_833,N_38);
nand U1367 (N_1367,N_941,N_803);
nand U1368 (N_1368,N_871,N_829);
or U1369 (N_1369,N_706,N_14);
nor U1370 (N_1370,N_278,N_396);
or U1371 (N_1371,N_388,N_926);
and U1372 (N_1372,N_451,N_987);
or U1373 (N_1373,N_134,N_327);
and U1374 (N_1374,N_34,N_550);
xnor U1375 (N_1375,N_353,N_354);
and U1376 (N_1376,N_943,N_839);
and U1377 (N_1377,N_50,N_215);
nor U1378 (N_1378,N_902,N_575);
nand U1379 (N_1379,N_665,N_567);
nor U1380 (N_1380,N_85,N_53);
nand U1381 (N_1381,N_450,N_457);
nor U1382 (N_1382,N_577,N_952);
nor U1383 (N_1383,N_750,N_193);
or U1384 (N_1384,N_876,N_507);
and U1385 (N_1385,N_249,N_556);
nand U1386 (N_1386,N_112,N_318);
nand U1387 (N_1387,N_449,N_771);
or U1388 (N_1388,N_288,N_452);
nor U1389 (N_1389,N_666,N_67);
nor U1390 (N_1390,N_131,N_19);
nor U1391 (N_1391,N_578,N_639);
or U1392 (N_1392,N_322,N_560);
or U1393 (N_1393,N_498,N_827);
nor U1394 (N_1394,N_315,N_127);
nand U1395 (N_1395,N_552,N_465);
and U1396 (N_1396,N_982,N_688);
or U1397 (N_1397,N_774,N_147);
nand U1398 (N_1398,N_524,N_241);
nor U1399 (N_1399,N_721,N_628);
and U1400 (N_1400,N_304,N_654);
nand U1401 (N_1401,N_202,N_406);
and U1402 (N_1402,N_511,N_569);
nand U1403 (N_1403,N_563,N_111);
and U1404 (N_1404,N_94,N_351);
or U1405 (N_1405,N_540,N_173);
xnor U1406 (N_1406,N_106,N_381);
or U1407 (N_1407,N_277,N_121);
nor U1408 (N_1408,N_767,N_58);
and U1409 (N_1409,N_163,N_159);
nor U1410 (N_1410,N_616,N_119);
and U1411 (N_1411,N_900,N_391);
or U1412 (N_1412,N_895,N_109);
and U1413 (N_1413,N_444,N_861);
nor U1414 (N_1414,N_585,N_476);
and U1415 (N_1415,N_724,N_872);
nand U1416 (N_1416,N_411,N_206);
nor U1417 (N_1417,N_662,N_500);
or U1418 (N_1418,N_905,N_918);
nand U1419 (N_1419,N_804,N_758);
nor U1420 (N_1420,N_909,N_733);
nand U1421 (N_1421,N_719,N_48);
nand U1422 (N_1422,N_828,N_120);
nor U1423 (N_1423,N_645,N_783);
nor U1424 (N_1424,N_228,N_855);
and U1425 (N_1425,N_257,N_30);
nor U1426 (N_1426,N_838,N_221);
nor U1427 (N_1427,N_350,N_901);
nand U1428 (N_1428,N_593,N_250);
nor U1429 (N_1429,N_258,N_613);
nand U1430 (N_1430,N_701,N_554);
and U1431 (N_1431,N_392,N_703);
nand U1432 (N_1432,N_693,N_648);
and U1433 (N_1433,N_18,N_223);
and U1434 (N_1434,N_748,N_337);
nand U1435 (N_1435,N_399,N_883);
or U1436 (N_1436,N_957,N_495);
and U1437 (N_1437,N_372,N_798);
nand U1438 (N_1438,N_929,N_262);
or U1439 (N_1439,N_934,N_966);
or U1440 (N_1440,N_636,N_983);
and U1441 (N_1441,N_331,N_105);
nand U1442 (N_1442,N_494,N_312);
nor U1443 (N_1443,N_780,N_502);
and U1444 (N_1444,N_432,N_283);
or U1445 (N_1445,N_959,N_181);
nand U1446 (N_1446,N_990,N_731);
nand U1447 (N_1447,N_775,N_738);
nor U1448 (N_1448,N_140,N_781);
and U1449 (N_1449,N_919,N_184);
nand U1450 (N_1450,N_425,N_124);
and U1451 (N_1451,N_462,N_128);
and U1452 (N_1452,N_908,N_232);
and U1453 (N_1453,N_778,N_346);
nor U1454 (N_1454,N_12,N_690);
and U1455 (N_1455,N_23,N_667);
nand U1456 (N_1456,N_641,N_626);
nand U1457 (N_1457,N_546,N_978);
nor U1458 (N_1458,N_176,N_461);
nand U1459 (N_1459,N_398,N_191);
and U1460 (N_1460,N_138,N_615);
and U1461 (N_1461,N_488,N_878);
nor U1462 (N_1462,N_225,N_623);
or U1463 (N_1463,N_888,N_489);
nand U1464 (N_1464,N_634,N_807);
and U1465 (N_1465,N_428,N_15);
nor U1466 (N_1466,N_689,N_307);
nor U1467 (N_1467,N_538,N_692);
nor U1468 (N_1468,N_300,N_9);
and U1469 (N_1469,N_866,N_348);
nor U1470 (N_1470,N_470,N_46);
and U1471 (N_1471,N_130,N_997);
and U1472 (N_1472,N_359,N_942);
and U1473 (N_1473,N_460,N_230);
and U1474 (N_1474,N_482,N_956);
and U1475 (N_1475,N_676,N_704);
or U1476 (N_1476,N_377,N_967);
nand U1477 (N_1477,N_785,N_509);
nand U1478 (N_1478,N_405,N_282);
and U1479 (N_1479,N_699,N_268);
or U1480 (N_1480,N_84,N_765);
nor U1481 (N_1481,N_116,N_604);
nand U1482 (N_1482,N_582,N_707);
nand U1483 (N_1483,N_455,N_831);
nor U1484 (N_1484,N_275,N_204);
and U1485 (N_1485,N_792,N_529);
nor U1486 (N_1486,N_35,N_848);
or U1487 (N_1487,N_877,N_113);
nand U1488 (N_1488,N_732,N_61);
xor U1489 (N_1489,N_820,N_685);
nor U1490 (N_1490,N_930,N_573);
nand U1491 (N_1491,N_149,N_551);
nand U1492 (N_1492,N_576,N_729);
and U1493 (N_1493,N_850,N_195);
nor U1494 (N_1494,N_882,N_600);
or U1495 (N_1495,N_603,N_339);
nand U1496 (N_1496,N_961,N_242);
nor U1497 (N_1497,N_525,N_261);
or U1498 (N_1498,N_316,N_794);
or U1499 (N_1499,N_336,N_141);
or U1500 (N_1500,N_894,N_490);
nand U1501 (N_1501,N_672,N_897);
and U1502 (N_1502,N_763,N_697);
nand U1503 (N_1503,N_423,N_365);
or U1504 (N_1504,N_180,N_219);
and U1505 (N_1505,N_423,N_152);
nor U1506 (N_1506,N_552,N_468);
and U1507 (N_1507,N_727,N_645);
nor U1508 (N_1508,N_957,N_633);
or U1509 (N_1509,N_640,N_404);
or U1510 (N_1510,N_371,N_466);
nor U1511 (N_1511,N_580,N_715);
nand U1512 (N_1512,N_189,N_914);
nand U1513 (N_1513,N_98,N_593);
nor U1514 (N_1514,N_174,N_802);
nand U1515 (N_1515,N_732,N_464);
nand U1516 (N_1516,N_842,N_247);
and U1517 (N_1517,N_26,N_450);
or U1518 (N_1518,N_864,N_505);
nand U1519 (N_1519,N_203,N_569);
or U1520 (N_1520,N_305,N_326);
nor U1521 (N_1521,N_817,N_848);
nand U1522 (N_1522,N_487,N_589);
or U1523 (N_1523,N_304,N_20);
nand U1524 (N_1524,N_817,N_727);
nor U1525 (N_1525,N_463,N_994);
or U1526 (N_1526,N_953,N_51);
nor U1527 (N_1527,N_325,N_408);
xor U1528 (N_1528,N_156,N_94);
or U1529 (N_1529,N_29,N_20);
or U1530 (N_1530,N_499,N_100);
or U1531 (N_1531,N_963,N_0);
and U1532 (N_1532,N_4,N_441);
nand U1533 (N_1533,N_105,N_70);
nand U1534 (N_1534,N_736,N_77);
and U1535 (N_1535,N_205,N_870);
and U1536 (N_1536,N_797,N_430);
nand U1537 (N_1537,N_100,N_72);
nor U1538 (N_1538,N_816,N_759);
and U1539 (N_1539,N_197,N_893);
and U1540 (N_1540,N_913,N_403);
nor U1541 (N_1541,N_52,N_133);
or U1542 (N_1542,N_878,N_261);
and U1543 (N_1543,N_251,N_569);
and U1544 (N_1544,N_911,N_418);
nor U1545 (N_1545,N_918,N_433);
and U1546 (N_1546,N_374,N_405);
and U1547 (N_1547,N_748,N_326);
nand U1548 (N_1548,N_262,N_934);
xnor U1549 (N_1549,N_29,N_988);
or U1550 (N_1550,N_894,N_901);
nor U1551 (N_1551,N_22,N_856);
or U1552 (N_1552,N_156,N_633);
or U1553 (N_1553,N_107,N_873);
nor U1554 (N_1554,N_921,N_991);
nand U1555 (N_1555,N_838,N_677);
nand U1556 (N_1556,N_431,N_875);
or U1557 (N_1557,N_768,N_810);
and U1558 (N_1558,N_447,N_209);
and U1559 (N_1559,N_893,N_838);
nor U1560 (N_1560,N_526,N_899);
and U1561 (N_1561,N_784,N_589);
nand U1562 (N_1562,N_559,N_595);
and U1563 (N_1563,N_693,N_731);
nand U1564 (N_1564,N_288,N_781);
and U1565 (N_1565,N_451,N_651);
nand U1566 (N_1566,N_6,N_225);
and U1567 (N_1567,N_596,N_534);
or U1568 (N_1568,N_91,N_199);
nand U1569 (N_1569,N_525,N_605);
xor U1570 (N_1570,N_45,N_214);
nand U1571 (N_1571,N_161,N_496);
and U1572 (N_1572,N_393,N_273);
nor U1573 (N_1573,N_208,N_595);
and U1574 (N_1574,N_914,N_689);
and U1575 (N_1575,N_413,N_126);
nor U1576 (N_1576,N_623,N_76);
nand U1577 (N_1577,N_321,N_525);
nor U1578 (N_1578,N_78,N_344);
xor U1579 (N_1579,N_58,N_975);
nor U1580 (N_1580,N_465,N_76);
nand U1581 (N_1581,N_603,N_119);
nand U1582 (N_1582,N_212,N_965);
or U1583 (N_1583,N_898,N_416);
and U1584 (N_1584,N_849,N_13);
or U1585 (N_1585,N_434,N_523);
xor U1586 (N_1586,N_835,N_344);
nand U1587 (N_1587,N_559,N_300);
nor U1588 (N_1588,N_711,N_511);
and U1589 (N_1589,N_623,N_798);
and U1590 (N_1590,N_1,N_492);
or U1591 (N_1591,N_527,N_663);
or U1592 (N_1592,N_585,N_323);
nand U1593 (N_1593,N_261,N_366);
and U1594 (N_1594,N_985,N_912);
nor U1595 (N_1595,N_790,N_926);
nand U1596 (N_1596,N_14,N_286);
and U1597 (N_1597,N_583,N_498);
nand U1598 (N_1598,N_321,N_518);
or U1599 (N_1599,N_930,N_911);
nand U1600 (N_1600,N_821,N_867);
and U1601 (N_1601,N_140,N_975);
nand U1602 (N_1602,N_745,N_104);
nand U1603 (N_1603,N_383,N_873);
and U1604 (N_1604,N_3,N_150);
nand U1605 (N_1605,N_493,N_162);
nand U1606 (N_1606,N_303,N_242);
nand U1607 (N_1607,N_403,N_183);
and U1608 (N_1608,N_693,N_781);
nor U1609 (N_1609,N_225,N_296);
nand U1610 (N_1610,N_232,N_406);
or U1611 (N_1611,N_739,N_827);
or U1612 (N_1612,N_629,N_375);
or U1613 (N_1613,N_860,N_239);
nor U1614 (N_1614,N_561,N_207);
nand U1615 (N_1615,N_726,N_193);
nor U1616 (N_1616,N_710,N_905);
nand U1617 (N_1617,N_603,N_492);
nand U1618 (N_1618,N_743,N_11);
nand U1619 (N_1619,N_4,N_526);
and U1620 (N_1620,N_864,N_798);
nor U1621 (N_1621,N_725,N_2);
or U1622 (N_1622,N_215,N_349);
or U1623 (N_1623,N_404,N_283);
nor U1624 (N_1624,N_933,N_280);
nand U1625 (N_1625,N_572,N_252);
nand U1626 (N_1626,N_427,N_463);
nand U1627 (N_1627,N_635,N_142);
nand U1628 (N_1628,N_289,N_121);
and U1629 (N_1629,N_174,N_368);
or U1630 (N_1630,N_176,N_72);
nand U1631 (N_1631,N_562,N_632);
and U1632 (N_1632,N_157,N_360);
and U1633 (N_1633,N_20,N_940);
or U1634 (N_1634,N_80,N_534);
nor U1635 (N_1635,N_72,N_210);
nand U1636 (N_1636,N_768,N_786);
nand U1637 (N_1637,N_646,N_713);
nand U1638 (N_1638,N_844,N_101);
xor U1639 (N_1639,N_439,N_843);
or U1640 (N_1640,N_802,N_459);
or U1641 (N_1641,N_112,N_579);
nor U1642 (N_1642,N_488,N_775);
and U1643 (N_1643,N_971,N_640);
nor U1644 (N_1644,N_305,N_677);
nand U1645 (N_1645,N_987,N_6);
xnor U1646 (N_1646,N_775,N_292);
nor U1647 (N_1647,N_502,N_836);
and U1648 (N_1648,N_592,N_734);
or U1649 (N_1649,N_543,N_580);
or U1650 (N_1650,N_450,N_204);
nor U1651 (N_1651,N_912,N_51);
xor U1652 (N_1652,N_776,N_459);
and U1653 (N_1653,N_438,N_193);
nand U1654 (N_1654,N_444,N_1);
or U1655 (N_1655,N_392,N_356);
nor U1656 (N_1656,N_57,N_839);
or U1657 (N_1657,N_90,N_936);
or U1658 (N_1658,N_695,N_244);
or U1659 (N_1659,N_732,N_517);
nor U1660 (N_1660,N_468,N_665);
nand U1661 (N_1661,N_864,N_371);
nor U1662 (N_1662,N_468,N_590);
or U1663 (N_1663,N_962,N_699);
and U1664 (N_1664,N_722,N_182);
or U1665 (N_1665,N_222,N_830);
nor U1666 (N_1666,N_448,N_389);
nand U1667 (N_1667,N_876,N_880);
nor U1668 (N_1668,N_354,N_779);
or U1669 (N_1669,N_514,N_747);
nand U1670 (N_1670,N_599,N_760);
nor U1671 (N_1671,N_250,N_716);
or U1672 (N_1672,N_21,N_258);
nand U1673 (N_1673,N_497,N_70);
nand U1674 (N_1674,N_210,N_782);
nor U1675 (N_1675,N_979,N_378);
nand U1676 (N_1676,N_37,N_961);
or U1677 (N_1677,N_247,N_401);
nor U1678 (N_1678,N_983,N_561);
and U1679 (N_1679,N_963,N_163);
and U1680 (N_1680,N_918,N_681);
nand U1681 (N_1681,N_621,N_134);
or U1682 (N_1682,N_300,N_445);
and U1683 (N_1683,N_490,N_146);
or U1684 (N_1684,N_183,N_409);
nor U1685 (N_1685,N_328,N_914);
nor U1686 (N_1686,N_48,N_196);
and U1687 (N_1687,N_752,N_821);
and U1688 (N_1688,N_808,N_485);
nand U1689 (N_1689,N_769,N_6);
and U1690 (N_1690,N_387,N_806);
and U1691 (N_1691,N_397,N_315);
or U1692 (N_1692,N_707,N_827);
and U1693 (N_1693,N_72,N_984);
xor U1694 (N_1694,N_373,N_417);
nand U1695 (N_1695,N_240,N_112);
nor U1696 (N_1696,N_112,N_132);
nor U1697 (N_1697,N_428,N_939);
nor U1698 (N_1698,N_857,N_558);
and U1699 (N_1699,N_44,N_498);
and U1700 (N_1700,N_283,N_92);
xor U1701 (N_1701,N_947,N_157);
nor U1702 (N_1702,N_82,N_161);
and U1703 (N_1703,N_303,N_188);
nor U1704 (N_1704,N_959,N_832);
nand U1705 (N_1705,N_992,N_715);
nand U1706 (N_1706,N_968,N_5);
and U1707 (N_1707,N_262,N_642);
or U1708 (N_1708,N_512,N_697);
nor U1709 (N_1709,N_415,N_431);
nand U1710 (N_1710,N_541,N_525);
or U1711 (N_1711,N_953,N_151);
nand U1712 (N_1712,N_522,N_587);
and U1713 (N_1713,N_18,N_607);
or U1714 (N_1714,N_809,N_627);
nor U1715 (N_1715,N_479,N_884);
and U1716 (N_1716,N_356,N_195);
or U1717 (N_1717,N_382,N_701);
nand U1718 (N_1718,N_810,N_999);
nand U1719 (N_1719,N_325,N_752);
or U1720 (N_1720,N_441,N_349);
or U1721 (N_1721,N_172,N_632);
nand U1722 (N_1722,N_476,N_643);
or U1723 (N_1723,N_690,N_910);
nand U1724 (N_1724,N_714,N_606);
nand U1725 (N_1725,N_683,N_947);
nor U1726 (N_1726,N_454,N_990);
and U1727 (N_1727,N_93,N_448);
nand U1728 (N_1728,N_94,N_339);
nand U1729 (N_1729,N_381,N_204);
nand U1730 (N_1730,N_393,N_626);
or U1731 (N_1731,N_968,N_95);
nor U1732 (N_1732,N_973,N_880);
or U1733 (N_1733,N_52,N_113);
nor U1734 (N_1734,N_290,N_82);
or U1735 (N_1735,N_812,N_999);
and U1736 (N_1736,N_210,N_794);
nor U1737 (N_1737,N_575,N_797);
nand U1738 (N_1738,N_97,N_672);
or U1739 (N_1739,N_442,N_16);
and U1740 (N_1740,N_969,N_902);
or U1741 (N_1741,N_746,N_509);
nor U1742 (N_1742,N_583,N_852);
nor U1743 (N_1743,N_663,N_472);
nor U1744 (N_1744,N_2,N_265);
nor U1745 (N_1745,N_940,N_931);
nand U1746 (N_1746,N_242,N_259);
and U1747 (N_1747,N_855,N_325);
and U1748 (N_1748,N_131,N_403);
nor U1749 (N_1749,N_41,N_975);
and U1750 (N_1750,N_30,N_966);
xnor U1751 (N_1751,N_488,N_294);
or U1752 (N_1752,N_985,N_489);
or U1753 (N_1753,N_1,N_448);
and U1754 (N_1754,N_914,N_756);
nor U1755 (N_1755,N_987,N_264);
nor U1756 (N_1756,N_284,N_303);
and U1757 (N_1757,N_311,N_306);
nand U1758 (N_1758,N_685,N_562);
nand U1759 (N_1759,N_639,N_635);
and U1760 (N_1760,N_276,N_647);
nor U1761 (N_1761,N_522,N_365);
xor U1762 (N_1762,N_192,N_18);
nor U1763 (N_1763,N_543,N_338);
nand U1764 (N_1764,N_693,N_973);
nand U1765 (N_1765,N_131,N_37);
nor U1766 (N_1766,N_191,N_266);
nor U1767 (N_1767,N_723,N_9);
nand U1768 (N_1768,N_216,N_981);
nand U1769 (N_1769,N_493,N_878);
and U1770 (N_1770,N_350,N_354);
and U1771 (N_1771,N_915,N_486);
or U1772 (N_1772,N_108,N_237);
nand U1773 (N_1773,N_1,N_37);
or U1774 (N_1774,N_921,N_768);
or U1775 (N_1775,N_546,N_238);
nor U1776 (N_1776,N_255,N_264);
nor U1777 (N_1777,N_334,N_330);
or U1778 (N_1778,N_128,N_360);
nand U1779 (N_1779,N_632,N_76);
and U1780 (N_1780,N_910,N_480);
nand U1781 (N_1781,N_149,N_161);
and U1782 (N_1782,N_646,N_832);
or U1783 (N_1783,N_383,N_953);
nand U1784 (N_1784,N_82,N_258);
or U1785 (N_1785,N_438,N_608);
nor U1786 (N_1786,N_781,N_861);
nor U1787 (N_1787,N_896,N_473);
and U1788 (N_1788,N_690,N_785);
nor U1789 (N_1789,N_877,N_324);
nand U1790 (N_1790,N_597,N_226);
and U1791 (N_1791,N_677,N_332);
or U1792 (N_1792,N_475,N_716);
or U1793 (N_1793,N_241,N_858);
nor U1794 (N_1794,N_239,N_153);
and U1795 (N_1795,N_910,N_958);
and U1796 (N_1796,N_828,N_465);
nor U1797 (N_1797,N_893,N_69);
or U1798 (N_1798,N_783,N_887);
nor U1799 (N_1799,N_48,N_681);
or U1800 (N_1800,N_24,N_292);
nand U1801 (N_1801,N_107,N_687);
or U1802 (N_1802,N_306,N_893);
nor U1803 (N_1803,N_445,N_579);
and U1804 (N_1804,N_824,N_635);
nand U1805 (N_1805,N_441,N_213);
nor U1806 (N_1806,N_367,N_761);
nand U1807 (N_1807,N_191,N_830);
and U1808 (N_1808,N_822,N_831);
and U1809 (N_1809,N_425,N_669);
and U1810 (N_1810,N_233,N_782);
or U1811 (N_1811,N_492,N_500);
or U1812 (N_1812,N_597,N_307);
nand U1813 (N_1813,N_153,N_615);
and U1814 (N_1814,N_626,N_209);
and U1815 (N_1815,N_883,N_853);
or U1816 (N_1816,N_659,N_607);
or U1817 (N_1817,N_172,N_770);
or U1818 (N_1818,N_670,N_335);
or U1819 (N_1819,N_113,N_916);
and U1820 (N_1820,N_260,N_792);
nand U1821 (N_1821,N_928,N_621);
nor U1822 (N_1822,N_84,N_287);
nand U1823 (N_1823,N_784,N_814);
or U1824 (N_1824,N_923,N_438);
and U1825 (N_1825,N_361,N_396);
and U1826 (N_1826,N_128,N_488);
nand U1827 (N_1827,N_630,N_993);
or U1828 (N_1828,N_846,N_965);
nor U1829 (N_1829,N_120,N_986);
and U1830 (N_1830,N_31,N_267);
or U1831 (N_1831,N_123,N_953);
nor U1832 (N_1832,N_523,N_201);
and U1833 (N_1833,N_238,N_65);
and U1834 (N_1834,N_680,N_414);
nand U1835 (N_1835,N_235,N_516);
and U1836 (N_1836,N_637,N_312);
nand U1837 (N_1837,N_770,N_686);
and U1838 (N_1838,N_347,N_871);
nor U1839 (N_1839,N_43,N_567);
or U1840 (N_1840,N_851,N_706);
or U1841 (N_1841,N_341,N_924);
and U1842 (N_1842,N_478,N_642);
and U1843 (N_1843,N_427,N_235);
nor U1844 (N_1844,N_250,N_26);
and U1845 (N_1845,N_956,N_790);
or U1846 (N_1846,N_40,N_735);
nand U1847 (N_1847,N_440,N_70);
nor U1848 (N_1848,N_566,N_830);
or U1849 (N_1849,N_352,N_783);
and U1850 (N_1850,N_212,N_530);
nand U1851 (N_1851,N_189,N_514);
and U1852 (N_1852,N_221,N_960);
xor U1853 (N_1853,N_128,N_795);
nand U1854 (N_1854,N_730,N_351);
or U1855 (N_1855,N_317,N_792);
nand U1856 (N_1856,N_740,N_622);
and U1857 (N_1857,N_715,N_672);
nand U1858 (N_1858,N_931,N_862);
nor U1859 (N_1859,N_912,N_944);
and U1860 (N_1860,N_80,N_609);
nor U1861 (N_1861,N_93,N_904);
or U1862 (N_1862,N_705,N_114);
nand U1863 (N_1863,N_89,N_115);
and U1864 (N_1864,N_387,N_114);
or U1865 (N_1865,N_563,N_884);
and U1866 (N_1866,N_442,N_327);
or U1867 (N_1867,N_618,N_689);
nand U1868 (N_1868,N_597,N_55);
nand U1869 (N_1869,N_640,N_298);
or U1870 (N_1870,N_387,N_601);
nand U1871 (N_1871,N_650,N_242);
nor U1872 (N_1872,N_21,N_579);
and U1873 (N_1873,N_267,N_558);
or U1874 (N_1874,N_727,N_44);
and U1875 (N_1875,N_744,N_252);
nor U1876 (N_1876,N_133,N_243);
nor U1877 (N_1877,N_32,N_93);
nand U1878 (N_1878,N_232,N_532);
nor U1879 (N_1879,N_225,N_53);
nand U1880 (N_1880,N_669,N_142);
or U1881 (N_1881,N_766,N_460);
nor U1882 (N_1882,N_183,N_30);
nor U1883 (N_1883,N_300,N_486);
nand U1884 (N_1884,N_300,N_81);
and U1885 (N_1885,N_24,N_918);
and U1886 (N_1886,N_731,N_668);
and U1887 (N_1887,N_669,N_127);
or U1888 (N_1888,N_731,N_562);
nand U1889 (N_1889,N_858,N_461);
nor U1890 (N_1890,N_590,N_995);
nor U1891 (N_1891,N_510,N_370);
nor U1892 (N_1892,N_47,N_646);
nor U1893 (N_1893,N_305,N_29);
and U1894 (N_1894,N_765,N_719);
or U1895 (N_1895,N_206,N_808);
nor U1896 (N_1896,N_710,N_968);
or U1897 (N_1897,N_845,N_689);
and U1898 (N_1898,N_476,N_504);
or U1899 (N_1899,N_528,N_105);
nand U1900 (N_1900,N_651,N_296);
nand U1901 (N_1901,N_899,N_344);
nor U1902 (N_1902,N_243,N_368);
and U1903 (N_1903,N_365,N_842);
xnor U1904 (N_1904,N_695,N_718);
nor U1905 (N_1905,N_358,N_367);
nor U1906 (N_1906,N_585,N_358);
and U1907 (N_1907,N_629,N_4);
or U1908 (N_1908,N_705,N_993);
nor U1909 (N_1909,N_615,N_633);
nor U1910 (N_1910,N_731,N_653);
and U1911 (N_1911,N_173,N_267);
nor U1912 (N_1912,N_154,N_662);
nand U1913 (N_1913,N_495,N_947);
nand U1914 (N_1914,N_266,N_150);
nand U1915 (N_1915,N_10,N_265);
and U1916 (N_1916,N_285,N_168);
nor U1917 (N_1917,N_185,N_449);
nand U1918 (N_1918,N_988,N_289);
nor U1919 (N_1919,N_819,N_22);
nand U1920 (N_1920,N_297,N_227);
nor U1921 (N_1921,N_82,N_175);
or U1922 (N_1922,N_267,N_702);
xor U1923 (N_1923,N_349,N_965);
and U1924 (N_1924,N_578,N_218);
nor U1925 (N_1925,N_355,N_209);
nand U1926 (N_1926,N_786,N_467);
nor U1927 (N_1927,N_9,N_959);
or U1928 (N_1928,N_808,N_292);
or U1929 (N_1929,N_46,N_441);
and U1930 (N_1930,N_859,N_894);
and U1931 (N_1931,N_1,N_874);
and U1932 (N_1932,N_552,N_895);
nand U1933 (N_1933,N_342,N_208);
nand U1934 (N_1934,N_548,N_963);
nand U1935 (N_1935,N_331,N_117);
or U1936 (N_1936,N_819,N_270);
and U1937 (N_1937,N_1,N_616);
nand U1938 (N_1938,N_567,N_769);
nand U1939 (N_1939,N_200,N_926);
nor U1940 (N_1940,N_277,N_978);
nand U1941 (N_1941,N_201,N_196);
nand U1942 (N_1942,N_626,N_521);
or U1943 (N_1943,N_152,N_621);
nand U1944 (N_1944,N_292,N_268);
nand U1945 (N_1945,N_47,N_391);
or U1946 (N_1946,N_87,N_571);
or U1947 (N_1947,N_582,N_525);
nand U1948 (N_1948,N_373,N_457);
xor U1949 (N_1949,N_400,N_248);
and U1950 (N_1950,N_721,N_307);
nor U1951 (N_1951,N_426,N_898);
nor U1952 (N_1952,N_804,N_425);
and U1953 (N_1953,N_575,N_199);
nor U1954 (N_1954,N_706,N_401);
and U1955 (N_1955,N_636,N_687);
or U1956 (N_1956,N_344,N_100);
nor U1957 (N_1957,N_944,N_465);
or U1958 (N_1958,N_359,N_84);
or U1959 (N_1959,N_957,N_762);
nand U1960 (N_1960,N_920,N_215);
and U1961 (N_1961,N_106,N_866);
nand U1962 (N_1962,N_936,N_859);
and U1963 (N_1963,N_925,N_183);
nor U1964 (N_1964,N_582,N_779);
or U1965 (N_1965,N_606,N_588);
or U1966 (N_1966,N_422,N_167);
nand U1967 (N_1967,N_378,N_780);
and U1968 (N_1968,N_725,N_652);
and U1969 (N_1969,N_818,N_690);
nand U1970 (N_1970,N_420,N_295);
and U1971 (N_1971,N_547,N_458);
nand U1972 (N_1972,N_528,N_873);
or U1973 (N_1973,N_822,N_863);
nor U1974 (N_1974,N_442,N_701);
and U1975 (N_1975,N_489,N_478);
or U1976 (N_1976,N_605,N_53);
or U1977 (N_1977,N_772,N_65);
nor U1978 (N_1978,N_968,N_875);
nor U1979 (N_1979,N_850,N_712);
and U1980 (N_1980,N_454,N_834);
nand U1981 (N_1981,N_354,N_740);
nand U1982 (N_1982,N_465,N_224);
nand U1983 (N_1983,N_928,N_946);
and U1984 (N_1984,N_556,N_166);
or U1985 (N_1985,N_722,N_682);
nand U1986 (N_1986,N_793,N_494);
or U1987 (N_1987,N_234,N_97);
and U1988 (N_1988,N_639,N_708);
and U1989 (N_1989,N_96,N_617);
or U1990 (N_1990,N_59,N_32);
nand U1991 (N_1991,N_694,N_188);
or U1992 (N_1992,N_574,N_423);
nor U1993 (N_1993,N_39,N_229);
nor U1994 (N_1994,N_727,N_301);
and U1995 (N_1995,N_557,N_767);
nand U1996 (N_1996,N_993,N_750);
nand U1997 (N_1997,N_800,N_354);
nor U1998 (N_1998,N_107,N_745);
and U1999 (N_1999,N_372,N_955);
nand U2000 (N_2000,N_1846,N_1158);
or U2001 (N_2001,N_1693,N_1476);
or U2002 (N_2002,N_1123,N_1606);
and U2003 (N_2003,N_1442,N_1874);
and U2004 (N_2004,N_1230,N_1330);
or U2005 (N_2005,N_1720,N_1459);
nand U2006 (N_2006,N_1537,N_1660);
nor U2007 (N_2007,N_1178,N_1722);
nand U2008 (N_2008,N_1916,N_1010);
nor U2009 (N_2009,N_1822,N_1550);
or U2010 (N_2010,N_1472,N_1908);
or U2011 (N_2011,N_1321,N_1081);
and U2012 (N_2012,N_1807,N_1617);
nor U2013 (N_2013,N_1160,N_1124);
nor U2014 (N_2014,N_1818,N_1083);
or U2015 (N_2015,N_1862,N_1892);
nor U2016 (N_2016,N_1518,N_1740);
or U2017 (N_2017,N_1630,N_1483);
nor U2018 (N_2018,N_1618,N_1546);
and U2019 (N_2019,N_1153,N_1134);
and U2020 (N_2020,N_1547,N_1402);
and U2021 (N_2021,N_1070,N_1551);
and U2022 (N_2022,N_1917,N_1837);
or U2023 (N_2023,N_1888,N_1405);
and U2024 (N_2024,N_1261,N_1318);
and U2025 (N_2025,N_1562,N_1161);
or U2026 (N_2026,N_1190,N_1085);
and U2027 (N_2027,N_1785,N_1584);
and U2028 (N_2028,N_1163,N_1866);
and U2029 (N_2029,N_1924,N_1912);
or U2030 (N_2030,N_1151,N_1231);
and U2031 (N_2031,N_1713,N_1854);
nor U2032 (N_2032,N_1669,N_1305);
nor U2033 (N_2033,N_1703,N_1358);
or U2034 (N_2034,N_1801,N_1991);
nor U2035 (N_2035,N_1401,N_1209);
nand U2036 (N_2036,N_1355,N_1212);
or U2037 (N_2037,N_1378,N_1311);
or U2038 (N_2038,N_1580,N_1296);
nor U2039 (N_2039,N_1838,N_1457);
and U2040 (N_2040,N_1569,N_1181);
and U2041 (N_2041,N_1220,N_1269);
or U2042 (N_2042,N_1666,N_1725);
and U2043 (N_2043,N_1205,N_1564);
and U2044 (N_2044,N_1880,N_1006);
or U2045 (N_2045,N_1646,N_1023);
and U2046 (N_2046,N_1492,N_1348);
nand U2047 (N_2047,N_1977,N_1688);
nand U2048 (N_2048,N_1030,N_1601);
nor U2049 (N_2049,N_1497,N_1040);
and U2050 (N_2050,N_1978,N_1241);
nor U2051 (N_2051,N_1967,N_1399);
nand U2052 (N_2052,N_1239,N_1450);
nor U2053 (N_2053,N_1806,N_1117);
xnor U2054 (N_2054,N_1841,N_1025);
or U2055 (N_2055,N_1088,N_1037);
and U2056 (N_2056,N_1288,N_1101);
nor U2057 (N_2057,N_1131,N_1108);
or U2058 (N_2058,N_1850,N_1571);
nor U2059 (N_2059,N_1326,N_1460);
and U2060 (N_2060,N_1298,N_1169);
nand U2061 (N_2061,N_1988,N_1707);
nor U2062 (N_2062,N_1835,N_1183);
nor U2063 (N_2063,N_1449,N_1334);
nor U2064 (N_2064,N_1362,N_1572);
or U2065 (N_2065,N_1777,N_1929);
nor U2066 (N_2066,N_1769,N_1337);
and U2067 (N_2067,N_1204,N_1155);
nor U2068 (N_2068,N_1346,N_1448);
nand U2069 (N_2069,N_1965,N_1727);
and U2070 (N_2070,N_1675,N_1258);
nand U2071 (N_2071,N_1671,N_1622);
nor U2072 (N_2072,N_1074,N_1097);
and U2073 (N_2073,N_1146,N_1833);
and U2074 (N_2074,N_1895,N_1637);
nor U2075 (N_2075,N_1726,N_1691);
or U2076 (N_2076,N_1628,N_1508);
and U2077 (N_2077,N_1073,N_1237);
nand U2078 (N_2078,N_1975,N_1232);
nand U2079 (N_2079,N_1772,N_1594);
nand U2080 (N_2080,N_1186,N_1779);
nand U2081 (N_2081,N_1263,N_1007);
or U2082 (N_2082,N_1044,N_1118);
or U2083 (N_2083,N_1271,N_1918);
and U2084 (N_2084,N_1620,N_1351);
and U2085 (N_2085,N_1819,N_1605);
and U2086 (N_2086,N_1940,N_1328);
and U2087 (N_2087,N_1112,N_1133);
and U2088 (N_2088,N_1008,N_1043);
nand U2089 (N_2089,N_1927,N_1453);
and U2090 (N_2090,N_1955,N_1140);
or U2091 (N_2091,N_1739,N_1150);
nand U2092 (N_2092,N_1502,N_1694);
and U2093 (N_2093,N_1934,N_1238);
and U2094 (N_2094,N_1111,N_1737);
nor U2095 (N_2095,N_1379,N_1214);
and U2096 (N_2096,N_1501,N_1811);
and U2097 (N_2097,N_1782,N_1469);
or U2098 (N_2098,N_1603,N_1657);
nand U2099 (N_2099,N_1122,N_1272);
and U2100 (N_2100,N_1254,N_1643);
nand U2101 (N_2101,N_1445,N_1413);
nand U2102 (N_2102,N_1059,N_1091);
nor U2103 (N_2103,N_1886,N_1555);
nor U2104 (N_2104,N_1522,N_1266);
nand U2105 (N_2105,N_1847,N_1187);
and U2106 (N_2106,N_1390,N_1909);
nor U2107 (N_2107,N_1233,N_1915);
nor U2108 (N_2108,N_1798,N_1937);
or U2109 (N_2109,N_1670,N_1293);
and U2110 (N_2110,N_1294,N_1487);
nand U2111 (N_2111,N_1260,N_1170);
and U2112 (N_2112,N_1574,N_1273);
and U2113 (N_2113,N_1535,N_1129);
nor U2114 (N_2114,N_1395,N_1333);
and U2115 (N_2115,N_1864,N_1175);
nand U2116 (N_2116,N_1229,N_1621);
or U2117 (N_2117,N_1114,N_1022);
or U2118 (N_2118,N_1996,N_1331);
or U2119 (N_2119,N_1945,N_1386);
or U2120 (N_2120,N_1180,N_1375);
nor U2121 (N_2121,N_1724,N_1468);
nor U2122 (N_2122,N_1394,N_1608);
and U2123 (N_2123,N_1455,N_1000);
nor U2124 (N_2124,N_1039,N_1141);
nor U2125 (N_2125,N_1932,N_1859);
nand U2126 (N_2126,N_1310,N_1420);
or U2127 (N_2127,N_1100,N_1877);
and U2128 (N_2128,N_1791,N_1650);
nor U2129 (N_2129,N_1174,N_1661);
nor U2130 (N_2130,N_1685,N_1454);
nor U2131 (N_2131,N_1905,N_1145);
and U2132 (N_2132,N_1464,N_1813);
nand U2133 (N_2133,N_1885,N_1890);
nand U2134 (N_2134,N_1686,N_1255);
nand U2135 (N_2135,N_1031,N_1887);
nor U2136 (N_2136,N_1611,N_1659);
xor U2137 (N_2137,N_1061,N_1530);
nand U2138 (N_2138,N_1494,N_1216);
or U2139 (N_2139,N_1075,N_1356);
nor U2140 (N_2140,N_1775,N_1166);
nand U2141 (N_2141,N_1200,N_1383);
nor U2142 (N_2142,N_1176,N_1964);
nand U2143 (N_2143,N_1997,N_1147);
nor U2144 (N_2144,N_1935,N_1849);
nand U2145 (N_2145,N_1519,N_1414);
nand U2146 (N_2146,N_1665,N_1540);
or U2147 (N_2147,N_1802,N_1872);
or U2148 (N_2148,N_1466,N_1552);
nor U2149 (N_2149,N_1962,N_1634);
and U2150 (N_2150,N_1322,N_1132);
nor U2151 (N_2151,N_1403,N_1089);
nand U2152 (N_2152,N_1753,N_1712);
and U2153 (N_2153,N_1277,N_1848);
nor U2154 (N_2154,N_1981,N_1461);
or U2155 (N_2155,N_1195,N_1647);
nand U2156 (N_2156,N_1409,N_1370);
or U2157 (N_2157,N_1248,N_1570);
nand U2158 (N_2158,N_1171,N_1065);
or U2159 (N_2159,N_1789,N_1870);
and U2160 (N_2160,N_1788,N_1361);
nand U2161 (N_2161,N_1165,N_1032);
nor U2162 (N_2162,N_1246,N_1878);
nor U2163 (N_2163,N_1410,N_1307);
nor U2164 (N_2164,N_1716,N_1920);
nor U2165 (N_2165,N_1289,N_1047);
or U2166 (N_2166,N_1808,N_1323);
and U2167 (N_2167,N_1583,N_1208);
or U2168 (N_2168,N_1076,N_1768);
nand U2169 (N_2169,N_1319,N_1149);
nand U2170 (N_2170,N_1324,N_1306);
and U2171 (N_2171,N_1327,N_1979);
nand U2172 (N_2172,N_1049,N_1910);
nand U2173 (N_2173,N_1938,N_1418);
or U2174 (N_2174,N_1470,N_1095);
nor U2175 (N_2175,N_1861,N_1704);
or U2176 (N_2176,N_1786,N_1179);
xor U2177 (N_2177,N_1268,N_1948);
and U2178 (N_2178,N_1335,N_1653);
or U2179 (N_2179,N_1684,N_1824);
nor U2180 (N_2180,N_1014,N_1343);
nand U2181 (N_2181,N_1471,N_1626);
or U2182 (N_2182,N_1731,N_1612);
or U2183 (N_2183,N_1677,N_1314);
nand U2184 (N_2184,N_1227,N_1102);
and U2185 (N_2185,N_1425,N_1009);
nor U2186 (N_2186,N_1104,N_1714);
or U2187 (N_2187,N_1667,N_1698);
nand U2188 (N_2188,N_1651,N_1780);
nand U2189 (N_2189,N_1052,N_1729);
or U2190 (N_2190,N_1096,N_1631);
nand U2191 (N_2191,N_1106,N_1435);
or U2192 (N_2192,N_1538,N_1863);
nor U2193 (N_2193,N_1919,N_1718);
and U2194 (N_2194,N_1963,N_1749);
or U2195 (N_2195,N_1893,N_1115);
nor U2196 (N_2196,N_1814,N_1256);
or U2197 (N_2197,N_1172,N_1773);
nand U2198 (N_2198,N_1527,N_1488);
and U2199 (N_2199,N_1350,N_1734);
nor U2200 (N_2200,N_1743,N_1816);
or U2201 (N_2201,N_1676,N_1558);
nand U2202 (N_2202,N_1090,N_1354);
nand U2203 (N_2203,N_1529,N_1914);
and U2204 (N_2204,N_1820,N_1856);
nand U2205 (N_2205,N_1315,N_1697);
nor U2206 (N_2206,N_1778,N_1826);
nor U2207 (N_2207,N_1093,N_1774);
nor U2208 (N_2208,N_1201,N_1286);
or U2209 (N_2209,N_1803,N_1048);
and U2210 (N_2210,N_1673,N_1719);
and U2211 (N_2211,N_1904,N_1994);
and U2212 (N_2212,N_1595,N_1028);
nor U2213 (N_2213,N_1462,N_1748);
nor U2214 (N_2214,N_1800,N_1236);
nor U2215 (N_2215,N_1336,N_1064);
nand U2216 (N_2216,N_1280,N_1591);
nand U2217 (N_2217,N_1264,N_1221);
nand U2218 (N_2218,N_1197,N_1278);
nand U2219 (N_2219,N_1687,N_1711);
nor U2220 (N_2220,N_1329,N_1270);
nor U2221 (N_2221,N_1983,N_1843);
nor U2222 (N_2222,N_1051,N_1559);
or U2223 (N_2223,N_1980,N_1013);
nand U2224 (N_2224,N_1341,N_1510);
nand U2225 (N_2225,N_1004,N_1512);
nor U2226 (N_2226,N_1185,N_1876);
nor U2227 (N_2227,N_1436,N_1489);
nor U2228 (N_2228,N_1478,N_1860);
nand U2229 (N_2229,N_1135,N_1344);
nand U2230 (N_2230,N_1762,N_1906);
nand U2231 (N_2231,N_1105,N_1857);
or U2232 (N_2232,N_1563,N_1079);
and U2233 (N_2233,N_1672,N_1641);
or U2234 (N_2234,N_1509,N_1827);
nand U2235 (N_2235,N_1444,N_1162);
and U2236 (N_2236,N_1257,N_1137);
nor U2237 (N_2237,N_1058,N_1451);
or U2238 (N_2238,N_1573,N_1223);
xor U2239 (N_2239,N_1506,N_1525);
or U2240 (N_2240,N_1923,N_1276);
nand U2241 (N_2241,N_1925,N_1053);
and U2242 (N_2242,N_1957,N_1699);
nand U2243 (N_2243,N_1426,N_1486);
nand U2244 (N_2244,N_1610,N_1654);
or U2245 (N_2245,N_1349,N_1359);
and U2246 (N_2246,N_1226,N_1655);
nor U2247 (N_2247,N_1407,N_1645);
nor U2248 (N_2248,N_1623,N_1730);
nor U2249 (N_2249,N_1871,N_1302);
nor U2250 (N_2250,N_1473,N_1602);
nor U2251 (N_2251,N_1303,N_1944);
nand U2252 (N_2252,N_1869,N_1928);
nor U2253 (N_2253,N_1590,N_1369);
or U2254 (N_2254,N_1222,N_1320);
nand U2255 (N_2255,N_1130,N_1228);
xnor U2256 (N_2256,N_1883,N_1950);
or U2257 (N_2257,N_1182,N_1732);
or U2258 (N_2258,N_1974,N_1365);
nand U2259 (N_2259,N_1971,N_1891);
nor U2260 (N_2260,N_1292,N_1556);
nor U2261 (N_2261,N_1968,N_1998);
or U2262 (N_2262,N_1879,N_1038);
and U2263 (N_2263,N_1882,N_1138);
nor U2264 (N_2264,N_1642,N_1560);
nor U2265 (N_2265,N_1250,N_1275);
or U2266 (N_2266,N_1218,N_1143);
nand U2267 (N_2267,N_1585,N_1252);
xnor U2268 (N_2268,N_1127,N_1274);
nor U2269 (N_2269,N_1939,N_1027);
nor U2270 (N_2270,N_1066,N_1215);
nand U2271 (N_2271,N_1219,N_1592);
xnor U2272 (N_2272,N_1682,N_1380);
and U2273 (N_2273,N_1279,N_1398);
nand U2274 (N_2274,N_1760,N_1858);
or U2275 (N_2275,N_1467,N_1553);
or U2276 (N_2276,N_1709,N_1986);
nor U2277 (N_2277,N_1763,N_1982);
and U2278 (N_2278,N_1363,N_1382);
nor U2279 (N_2279,N_1504,N_1701);
and U2280 (N_2280,N_1217,N_1539);
or U2281 (N_2281,N_1071,N_1679);
nand U2282 (N_2282,N_1507,N_1285);
or U2283 (N_2283,N_1596,N_1514);
and U2284 (N_2284,N_1723,N_1804);
nor U2285 (N_2285,N_1068,N_1050);
xnor U2286 (N_2286,N_1317,N_1851);
nor U2287 (N_2287,N_1126,N_1735);
nor U2288 (N_2288,N_1951,N_1521);
nor U2289 (N_2289,N_1503,N_1253);
or U2290 (N_2290,N_1958,N_1441);
xor U2291 (N_2291,N_1831,N_1084);
xor U2292 (N_2292,N_1003,N_1531);
nand U2293 (N_2293,N_1644,N_1404);
or U2294 (N_2294,N_1598,N_1913);
nor U2295 (N_2295,N_1568,N_1954);
or U2296 (N_2296,N_1830,N_1304);
and U2297 (N_2297,N_1588,N_1211);
or U2298 (N_2298,N_1392,N_1192);
and U2299 (N_2299,N_1309,N_1867);
or U2300 (N_2300,N_1198,N_1668);
nor U2301 (N_2301,N_1832,N_1548);
and U2302 (N_2302,N_1952,N_1943);
nor U2303 (N_2303,N_1931,N_1499);
nand U2304 (N_2304,N_1406,N_1247);
nand U2305 (N_2305,N_1136,N_1479);
nand U2306 (N_2306,N_1312,N_1125);
and U2307 (N_2307,N_1225,N_1812);
and U2308 (N_2308,N_1224,N_1751);
or U2309 (N_2309,N_1056,N_1528);
nand U2310 (N_2310,N_1689,N_1029);
and U2311 (N_2311,N_1235,N_1947);
and U2312 (N_2312,N_1578,N_1002);
nor U2313 (N_2313,N_1416,N_1152);
or U2314 (N_2314,N_1034,N_1524);
nor U2315 (N_2315,N_1385,N_1475);
or U2316 (N_2316,N_1234,N_1616);
nor U2317 (N_2317,N_1244,N_1098);
and U2318 (N_2318,N_1092,N_1485);
nor U2319 (N_2319,N_1062,N_1443);
nor U2320 (N_2320,N_1364,N_1120);
or U2321 (N_2321,N_1770,N_1961);
nor U2322 (N_2322,N_1993,N_1700);
nand U2323 (N_2323,N_1884,N_1301);
nand U2324 (N_2324,N_1297,N_1020);
nor U2325 (N_2325,N_1017,N_1173);
or U2326 (N_2326,N_1683,N_1526);
or U2327 (N_2327,N_1889,N_1121);
or U2328 (N_2328,N_1805,N_1565);
nand U2329 (N_2329,N_1295,N_1128);
and U2330 (N_2330,N_1432,N_1855);
nor U2331 (N_2331,N_1078,N_1755);
and U2332 (N_2332,N_1463,N_1313);
and U2333 (N_2333,N_1781,N_1619);
nand U2334 (N_2334,N_1391,N_1408);
and U2335 (N_2335,N_1823,N_1139);
and U2336 (N_2336,N_1992,N_1148);
nor U2337 (N_2337,N_1873,N_1894);
and U2338 (N_2338,N_1541,N_1576);
and U2339 (N_2339,N_1439,N_1377);
nor U2340 (N_2340,N_1899,N_1692);
nor U2341 (N_2341,N_1845,N_1946);
or U2342 (N_2342,N_1784,N_1374);
and U2343 (N_2343,N_1103,N_1629);
and U2344 (N_2344,N_1157,N_1953);
and U2345 (N_2345,N_1736,N_1480);
or U2346 (N_2346,N_1520,N_1533);
and U2347 (N_2347,N_1373,N_1505);
or U2348 (N_2348,N_1119,N_1368);
nor U2349 (N_2349,N_1465,N_1156);
nor U2350 (N_2350,N_1767,N_1396);
nor U2351 (N_2351,N_1761,N_1589);
and U2352 (N_2352,N_1082,N_1168);
or U2353 (N_2353,N_1949,N_1633);
and U2354 (N_2354,N_1787,N_1393);
nand U2355 (N_2355,N_1005,N_1290);
or U2356 (N_2356,N_1352,N_1754);
or U2357 (N_2357,N_1207,N_1911);
and U2358 (N_2358,N_1376,N_1663);
or U2359 (N_2359,N_1999,N_1747);
nand U2360 (N_2360,N_1844,N_1446);
or U2361 (N_2361,N_1639,N_1387);
nor U2362 (N_2362,N_1721,N_1021);
or U2363 (N_2363,N_1708,N_1842);
or U2364 (N_2364,N_1243,N_1345);
nand U2365 (N_2365,N_1907,N_1680);
nor U2366 (N_2366,N_1177,N_1976);
nor U2367 (N_2367,N_1245,N_1771);
or U2368 (N_2368,N_1422,N_1549);
or U2369 (N_2369,N_1417,N_1500);
nor U2370 (N_2370,N_1491,N_1933);
nor U2371 (N_2371,N_1636,N_1566);
or U2372 (N_2372,N_1960,N_1203);
nor U2373 (N_2373,N_1109,N_1752);
or U2374 (N_2374,N_1926,N_1498);
nor U2375 (N_2375,N_1340,N_1710);
or U2376 (N_2376,N_1715,N_1069);
nand U2377 (N_2377,N_1759,N_1440);
xor U2378 (N_2378,N_1447,N_1625);
or U2379 (N_2379,N_1490,N_1987);
and U2380 (N_2380,N_1875,N_1678);
nand U2381 (N_2381,N_1430,N_1116);
and U2382 (N_2382,N_1587,N_1696);
nand U2383 (N_2383,N_1371,N_1632);
or U2384 (N_2384,N_1366,N_1903);
nand U2385 (N_2385,N_1901,N_1164);
nand U2386 (N_2386,N_1015,N_1188);
nor U2387 (N_2387,N_1597,N_1193);
and U2388 (N_2388,N_1431,N_1249);
nor U2389 (N_2389,N_1766,N_1989);
and U2390 (N_2390,N_1742,N_1966);
or U2391 (N_2391,N_1154,N_1419);
nand U2392 (N_2392,N_1536,N_1615);
nor U2393 (N_2393,N_1389,N_1400);
or U2394 (N_2394,N_1360,N_1900);
nor U2395 (N_2395,N_1199,N_1339);
nand U2396 (N_2396,N_1438,N_1144);
or U2397 (N_2397,N_1815,N_1080);
or U2398 (N_2398,N_1458,N_1757);
nor U2399 (N_2399,N_1744,N_1575);
nor U2400 (N_2400,N_1746,N_1242);
nand U2401 (N_2401,N_1086,N_1959);
or U2402 (N_2402,N_1415,N_1424);
nand U2403 (N_2403,N_1695,N_1561);
or U2404 (N_2404,N_1107,N_1809);
nand U2405 (N_2405,N_1523,N_1299);
nor U2406 (N_2406,N_1113,N_1664);
nand U2407 (N_2407,N_1018,N_1702);
or U2408 (N_2408,N_1033,N_1593);
and U2409 (N_2409,N_1388,N_1011);
nand U2410 (N_2410,N_1790,N_1493);
nand U2411 (N_2411,N_1300,N_1110);
xnor U2412 (N_2412,N_1001,N_1599);
nor U2413 (N_2413,N_1936,N_1482);
and U2414 (N_2414,N_1036,N_1452);
and U2415 (N_2415,N_1706,N_1542);
or U2416 (N_2416,N_1793,N_1338);
nand U2417 (N_2417,N_1184,N_1159);
or U2418 (N_2418,N_1434,N_1627);
or U2419 (N_2419,N_1969,N_1072);
or U2420 (N_2420,N_1635,N_1705);
and U2421 (N_2421,N_1828,N_1477);
nor U2422 (N_2422,N_1972,N_1532);
or U2423 (N_2423,N_1194,N_1956);
nand U2424 (N_2424,N_1821,N_1412);
and U2425 (N_2425,N_1041,N_1579);
and U2426 (N_2426,N_1662,N_1087);
or U2427 (N_2427,N_1984,N_1829);
nand U2428 (N_2428,N_1191,N_1674);
nor U2429 (N_2429,N_1795,N_1853);
and U2430 (N_2430,N_1019,N_1045);
and U2431 (N_2431,N_1796,N_1728);
or U2432 (N_2432,N_1985,N_1638);
and U2433 (N_2433,N_1604,N_1291);
nand U2434 (N_2434,N_1557,N_1429);
nor U2435 (N_2435,N_1681,N_1240);
nor U2436 (N_2436,N_1783,N_1516);
or U2437 (N_2437,N_1517,N_1267);
nand U2438 (N_2438,N_1411,N_1776);
and U2439 (N_2439,N_1834,N_1745);
and U2440 (N_2440,N_1099,N_1836);
and U2441 (N_2441,N_1283,N_1658);
nor U2442 (N_2442,N_1024,N_1582);
and U2443 (N_2443,N_1060,N_1481);
nand U2444 (N_2444,N_1428,N_1012);
and U2445 (N_2445,N_1281,N_1750);
or U2446 (N_2446,N_1995,N_1534);
or U2447 (N_2447,N_1921,N_1973);
or U2448 (N_2448,N_1262,N_1554);
nor U2449 (N_2449,N_1251,N_1758);
and U2450 (N_2450,N_1213,N_1941);
nand U2451 (N_2451,N_1581,N_1607);
and U2452 (N_2452,N_1067,N_1733);
and U2453 (N_2453,N_1035,N_1545);
or U2454 (N_2454,N_1189,N_1543);
nor U2455 (N_2455,N_1840,N_1042);
nor U2456 (N_2456,N_1342,N_1839);
or U2457 (N_2457,N_1325,N_1496);
or U2458 (N_2458,N_1797,N_1613);
nor U2459 (N_2459,N_1384,N_1609);
nand U2460 (N_2460,N_1624,N_1421);
and U2461 (N_2461,N_1817,N_1765);
or U2462 (N_2462,N_1054,N_1942);
and U2463 (N_2463,N_1756,N_1287);
and U2464 (N_2464,N_1614,N_1196);
nand U2465 (N_2465,N_1852,N_1437);
or U2466 (N_2466,N_1881,N_1764);
nor U2467 (N_2467,N_1922,N_1717);
and U2468 (N_2468,N_1094,N_1577);
nand U2469 (N_2469,N_1427,N_1690);
and U2470 (N_2470,N_1738,N_1026);
nand U2471 (N_2471,N_1057,N_1741);
and U2472 (N_2472,N_1357,N_1896);
or U2473 (N_2473,N_1077,N_1381);
and U2474 (N_2474,N_1586,N_1474);
or U2475 (N_2475,N_1063,N_1799);
nor U2476 (N_2476,N_1016,N_1810);
nor U2477 (N_2477,N_1046,N_1332);
nand U2478 (N_2478,N_1656,N_1456);
and U2479 (N_2479,N_1897,N_1640);
and U2480 (N_2480,N_1794,N_1423);
or U2481 (N_2481,N_1353,N_1649);
or U2482 (N_2482,N_1868,N_1515);
xnor U2483 (N_2483,N_1347,N_1167);
and U2484 (N_2484,N_1544,N_1206);
nor U2485 (N_2485,N_1600,N_1652);
or U2486 (N_2486,N_1567,N_1259);
or U2487 (N_2487,N_1825,N_1511);
and U2488 (N_2488,N_1055,N_1433);
nand U2489 (N_2489,N_1202,N_1990);
and U2490 (N_2490,N_1648,N_1284);
and U2491 (N_2491,N_1282,N_1367);
nor U2492 (N_2492,N_1265,N_1142);
or U2493 (N_2493,N_1484,N_1898);
nand U2494 (N_2494,N_1513,N_1930);
or U2495 (N_2495,N_1210,N_1902);
or U2496 (N_2496,N_1316,N_1792);
and U2497 (N_2497,N_1970,N_1308);
nor U2498 (N_2498,N_1372,N_1865);
nor U2499 (N_2499,N_1397,N_1495);
or U2500 (N_2500,N_1602,N_1028);
and U2501 (N_2501,N_1782,N_1984);
and U2502 (N_2502,N_1597,N_1636);
nor U2503 (N_2503,N_1570,N_1400);
and U2504 (N_2504,N_1224,N_1740);
nand U2505 (N_2505,N_1088,N_1189);
and U2506 (N_2506,N_1533,N_1039);
nor U2507 (N_2507,N_1477,N_1478);
nor U2508 (N_2508,N_1050,N_1957);
nor U2509 (N_2509,N_1712,N_1090);
nand U2510 (N_2510,N_1558,N_1885);
nand U2511 (N_2511,N_1098,N_1254);
nand U2512 (N_2512,N_1629,N_1058);
or U2513 (N_2513,N_1507,N_1007);
and U2514 (N_2514,N_1849,N_1752);
or U2515 (N_2515,N_1882,N_1742);
or U2516 (N_2516,N_1884,N_1380);
nor U2517 (N_2517,N_1748,N_1877);
or U2518 (N_2518,N_1581,N_1494);
or U2519 (N_2519,N_1467,N_1854);
nor U2520 (N_2520,N_1571,N_1218);
nor U2521 (N_2521,N_1894,N_1342);
and U2522 (N_2522,N_1770,N_1527);
nand U2523 (N_2523,N_1335,N_1478);
and U2524 (N_2524,N_1576,N_1826);
or U2525 (N_2525,N_1891,N_1220);
xor U2526 (N_2526,N_1124,N_1440);
or U2527 (N_2527,N_1880,N_1336);
nor U2528 (N_2528,N_1990,N_1429);
and U2529 (N_2529,N_1329,N_1064);
and U2530 (N_2530,N_1122,N_1521);
nand U2531 (N_2531,N_1808,N_1612);
and U2532 (N_2532,N_1820,N_1091);
nor U2533 (N_2533,N_1680,N_1374);
nor U2534 (N_2534,N_1118,N_1976);
nor U2535 (N_2535,N_1530,N_1383);
or U2536 (N_2536,N_1534,N_1544);
nor U2537 (N_2537,N_1963,N_1494);
and U2538 (N_2538,N_1509,N_1830);
and U2539 (N_2539,N_1561,N_1067);
nor U2540 (N_2540,N_1441,N_1308);
or U2541 (N_2541,N_1562,N_1258);
nand U2542 (N_2542,N_1193,N_1678);
and U2543 (N_2543,N_1422,N_1044);
nor U2544 (N_2544,N_1751,N_1095);
nand U2545 (N_2545,N_1320,N_1728);
nand U2546 (N_2546,N_1030,N_1542);
and U2547 (N_2547,N_1658,N_1023);
nand U2548 (N_2548,N_1524,N_1473);
nor U2549 (N_2549,N_1642,N_1715);
and U2550 (N_2550,N_1104,N_1581);
and U2551 (N_2551,N_1614,N_1848);
and U2552 (N_2552,N_1757,N_1871);
and U2553 (N_2553,N_1372,N_1288);
nor U2554 (N_2554,N_1443,N_1633);
or U2555 (N_2555,N_1081,N_1238);
nand U2556 (N_2556,N_1619,N_1519);
and U2557 (N_2557,N_1085,N_1054);
nor U2558 (N_2558,N_1316,N_1379);
and U2559 (N_2559,N_1492,N_1330);
and U2560 (N_2560,N_1560,N_1578);
or U2561 (N_2561,N_1541,N_1353);
nor U2562 (N_2562,N_1356,N_1030);
or U2563 (N_2563,N_1632,N_1271);
or U2564 (N_2564,N_1099,N_1750);
xor U2565 (N_2565,N_1264,N_1686);
nand U2566 (N_2566,N_1752,N_1357);
nor U2567 (N_2567,N_1211,N_1621);
or U2568 (N_2568,N_1730,N_1722);
xnor U2569 (N_2569,N_1154,N_1608);
nand U2570 (N_2570,N_1481,N_1242);
nand U2571 (N_2571,N_1906,N_1367);
nor U2572 (N_2572,N_1924,N_1155);
nand U2573 (N_2573,N_1876,N_1242);
nand U2574 (N_2574,N_1085,N_1158);
and U2575 (N_2575,N_1365,N_1515);
and U2576 (N_2576,N_1252,N_1123);
and U2577 (N_2577,N_1938,N_1899);
and U2578 (N_2578,N_1351,N_1693);
nor U2579 (N_2579,N_1211,N_1134);
nor U2580 (N_2580,N_1537,N_1816);
or U2581 (N_2581,N_1768,N_1213);
or U2582 (N_2582,N_1831,N_1670);
nand U2583 (N_2583,N_1982,N_1130);
nand U2584 (N_2584,N_1779,N_1912);
or U2585 (N_2585,N_1896,N_1141);
or U2586 (N_2586,N_1224,N_1282);
nand U2587 (N_2587,N_1625,N_1380);
nand U2588 (N_2588,N_1720,N_1147);
or U2589 (N_2589,N_1098,N_1300);
or U2590 (N_2590,N_1560,N_1712);
nor U2591 (N_2591,N_1454,N_1279);
nor U2592 (N_2592,N_1041,N_1163);
or U2593 (N_2593,N_1158,N_1714);
or U2594 (N_2594,N_1401,N_1247);
or U2595 (N_2595,N_1082,N_1248);
nand U2596 (N_2596,N_1089,N_1629);
or U2597 (N_2597,N_1788,N_1100);
or U2598 (N_2598,N_1058,N_1182);
nand U2599 (N_2599,N_1264,N_1676);
nor U2600 (N_2600,N_1104,N_1169);
and U2601 (N_2601,N_1150,N_1163);
nor U2602 (N_2602,N_1939,N_1703);
nor U2603 (N_2603,N_1022,N_1509);
nor U2604 (N_2604,N_1841,N_1690);
nor U2605 (N_2605,N_1010,N_1499);
or U2606 (N_2606,N_1662,N_1120);
or U2607 (N_2607,N_1628,N_1637);
nor U2608 (N_2608,N_1222,N_1849);
nand U2609 (N_2609,N_1563,N_1817);
nor U2610 (N_2610,N_1511,N_1391);
nand U2611 (N_2611,N_1702,N_1680);
nor U2612 (N_2612,N_1649,N_1999);
nor U2613 (N_2613,N_1005,N_1807);
nor U2614 (N_2614,N_1223,N_1689);
or U2615 (N_2615,N_1199,N_1311);
and U2616 (N_2616,N_1723,N_1156);
and U2617 (N_2617,N_1893,N_1842);
nand U2618 (N_2618,N_1230,N_1463);
nand U2619 (N_2619,N_1942,N_1880);
and U2620 (N_2620,N_1858,N_1964);
or U2621 (N_2621,N_1022,N_1903);
nor U2622 (N_2622,N_1352,N_1955);
nand U2623 (N_2623,N_1843,N_1063);
or U2624 (N_2624,N_1008,N_1857);
nor U2625 (N_2625,N_1038,N_1876);
nand U2626 (N_2626,N_1092,N_1244);
and U2627 (N_2627,N_1868,N_1398);
nand U2628 (N_2628,N_1058,N_1620);
or U2629 (N_2629,N_1514,N_1834);
or U2630 (N_2630,N_1718,N_1374);
and U2631 (N_2631,N_1670,N_1356);
and U2632 (N_2632,N_1035,N_1440);
and U2633 (N_2633,N_1703,N_1768);
xnor U2634 (N_2634,N_1189,N_1682);
nor U2635 (N_2635,N_1207,N_1419);
or U2636 (N_2636,N_1314,N_1383);
and U2637 (N_2637,N_1801,N_1911);
nor U2638 (N_2638,N_1751,N_1445);
nor U2639 (N_2639,N_1553,N_1299);
and U2640 (N_2640,N_1348,N_1541);
or U2641 (N_2641,N_1106,N_1814);
or U2642 (N_2642,N_1217,N_1202);
or U2643 (N_2643,N_1904,N_1337);
nand U2644 (N_2644,N_1574,N_1399);
nand U2645 (N_2645,N_1703,N_1384);
nand U2646 (N_2646,N_1784,N_1383);
and U2647 (N_2647,N_1033,N_1937);
nor U2648 (N_2648,N_1630,N_1735);
nand U2649 (N_2649,N_1421,N_1899);
or U2650 (N_2650,N_1807,N_1514);
or U2651 (N_2651,N_1132,N_1588);
xnor U2652 (N_2652,N_1652,N_1358);
or U2653 (N_2653,N_1020,N_1110);
nor U2654 (N_2654,N_1601,N_1063);
nor U2655 (N_2655,N_1708,N_1392);
nor U2656 (N_2656,N_1866,N_1903);
or U2657 (N_2657,N_1858,N_1674);
nor U2658 (N_2658,N_1001,N_1948);
nand U2659 (N_2659,N_1422,N_1264);
nor U2660 (N_2660,N_1629,N_1808);
nor U2661 (N_2661,N_1248,N_1635);
or U2662 (N_2662,N_1101,N_1516);
nand U2663 (N_2663,N_1407,N_1824);
and U2664 (N_2664,N_1072,N_1192);
nor U2665 (N_2665,N_1413,N_1786);
nor U2666 (N_2666,N_1139,N_1790);
nand U2667 (N_2667,N_1735,N_1594);
or U2668 (N_2668,N_1914,N_1118);
nor U2669 (N_2669,N_1325,N_1725);
or U2670 (N_2670,N_1714,N_1880);
nand U2671 (N_2671,N_1116,N_1340);
nor U2672 (N_2672,N_1046,N_1580);
or U2673 (N_2673,N_1538,N_1752);
or U2674 (N_2674,N_1996,N_1566);
nor U2675 (N_2675,N_1849,N_1692);
or U2676 (N_2676,N_1149,N_1474);
and U2677 (N_2677,N_1826,N_1629);
nor U2678 (N_2678,N_1861,N_1558);
or U2679 (N_2679,N_1551,N_1473);
nor U2680 (N_2680,N_1403,N_1133);
or U2681 (N_2681,N_1703,N_1447);
or U2682 (N_2682,N_1039,N_1562);
nor U2683 (N_2683,N_1668,N_1492);
or U2684 (N_2684,N_1751,N_1315);
xnor U2685 (N_2685,N_1217,N_1974);
nor U2686 (N_2686,N_1601,N_1715);
and U2687 (N_2687,N_1639,N_1452);
nand U2688 (N_2688,N_1146,N_1768);
nand U2689 (N_2689,N_1045,N_1905);
nand U2690 (N_2690,N_1752,N_1497);
nand U2691 (N_2691,N_1970,N_1856);
and U2692 (N_2692,N_1466,N_1599);
nand U2693 (N_2693,N_1255,N_1195);
or U2694 (N_2694,N_1761,N_1595);
or U2695 (N_2695,N_1403,N_1584);
nor U2696 (N_2696,N_1728,N_1810);
and U2697 (N_2697,N_1532,N_1943);
or U2698 (N_2698,N_1989,N_1081);
nor U2699 (N_2699,N_1721,N_1684);
or U2700 (N_2700,N_1951,N_1608);
or U2701 (N_2701,N_1940,N_1538);
or U2702 (N_2702,N_1491,N_1714);
and U2703 (N_2703,N_1608,N_1508);
nand U2704 (N_2704,N_1866,N_1139);
and U2705 (N_2705,N_1612,N_1084);
or U2706 (N_2706,N_1907,N_1594);
nor U2707 (N_2707,N_1785,N_1374);
and U2708 (N_2708,N_1100,N_1319);
nand U2709 (N_2709,N_1748,N_1230);
nor U2710 (N_2710,N_1460,N_1396);
nand U2711 (N_2711,N_1109,N_1025);
or U2712 (N_2712,N_1042,N_1640);
or U2713 (N_2713,N_1728,N_1011);
or U2714 (N_2714,N_1250,N_1269);
or U2715 (N_2715,N_1708,N_1138);
and U2716 (N_2716,N_1987,N_1345);
or U2717 (N_2717,N_1108,N_1506);
nand U2718 (N_2718,N_1523,N_1422);
or U2719 (N_2719,N_1824,N_1857);
nand U2720 (N_2720,N_1573,N_1398);
xnor U2721 (N_2721,N_1914,N_1188);
nand U2722 (N_2722,N_1515,N_1691);
nor U2723 (N_2723,N_1347,N_1149);
and U2724 (N_2724,N_1746,N_1444);
nor U2725 (N_2725,N_1177,N_1270);
and U2726 (N_2726,N_1611,N_1779);
nor U2727 (N_2727,N_1846,N_1234);
nand U2728 (N_2728,N_1467,N_1471);
or U2729 (N_2729,N_1836,N_1938);
nor U2730 (N_2730,N_1361,N_1427);
or U2731 (N_2731,N_1947,N_1517);
and U2732 (N_2732,N_1241,N_1064);
nor U2733 (N_2733,N_1512,N_1647);
nand U2734 (N_2734,N_1020,N_1097);
nand U2735 (N_2735,N_1106,N_1191);
or U2736 (N_2736,N_1010,N_1344);
and U2737 (N_2737,N_1408,N_1029);
nand U2738 (N_2738,N_1245,N_1015);
and U2739 (N_2739,N_1652,N_1898);
nand U2740 (N_2740,N_1671,N_1281);
nand U2741 (N_2741,N_1628,N_1877);
nor U2742 (N_2742,N_1604,N_1276);
nand U2743 (N_2743,N_1717,N_1510);
nor U2744 (N_2744,N_1662,N_1146);
nand U2745 (N_2745,N_1118,N_1912);
nand U2746 (N_2746,N_1805,N_1966);
or U2747 (N_2747,N_1577,N_1848);
nor U2748 (N_2748,N_1234,N_1547);
nand U2749 (N_2749,N_1700,N_1072);
nor U2750 (N_2750,N_1991,N_1075);
or U2751 (N_2751,N_1746,N_1363);
nand U2752 (N_2752,N_1367,N_1416);
nand U2753 (N_2753,N_1169,N_1891);
nand U2754 (N_2754,N_1471,N_1096);
nor U2755 (N_2755,N_1275,N_1329);
and U2756 (N_2756,N_1171,N_1718);
and U2757 (N_2757,N_1471,N_1684);
xor U2758 (N_2758,N_1115,N_1660);
and U2759 (N_2759,N_1778,N_1179);
or U2760 (N_2760,N_1467,N_1912);
or U2761 (N_2761,N_1997,N_1743);
and U2762 (N_2762,N_1893,N_1301);
and U2763 (N_2763,N_1630,N_1568);
or U2764 (N_2764,N_1057,N_1560);
or U2765 (N_2765,N_1880,N_1345);
nand U2766 (N_2766,N_1818,N_1485);
nor U2767 (N_2767,N_1166,N_1248);
nand U2768 (N_2768,N_1811,N_1424);
or U2769 (N_2769,N_1462,N_1400);
or U2770 (N_2770,N_1521,N_1959);
nand U2771 (N_2771,N_1363,N_1010);
and U2772 (N_2772,N_1617,N_1194);
or U2773 (N_2773,N_1003,N_1894);
or U2774 (N_2774,N_1345,N_1959);
nand U2775 (N_2775,N_1482,N_1131);
nor U2776 (N_2776,N_1760,N_1184);
or U2777 (N_2777,N_1648,N_1289);
and U2778 (N_2778,N_1016,N_1000);
and U2779 (N_2779,N_1598,N_1528);
and U2780 (N_2780,N_1312,N_1788);
nand U2781 (N_2781,N_1218,N_1813);
nor U2782 (N_2782,N_1585,N_1364);
nand U2783 (N_2783,N_1831,N_1610);
and U2784 (N_2784,N_1408,N_1483);
or U2785 (N_2785,N_1527,N_1410);
and U2786 (N_2786,N_1293,N_1376);
and U2787 (N_2787,N_1421,N_1765);
nor U2788 (N_2788,N_1501,N_1009);
or U2789 (N_2789,N_1892,N_1283);
or U2790 (N_2790,N_1251,N_1075);
nand U2791 (N_2791,N_1739,N_1470);
nand U2792 (N_2792,N_1267,N_1760);
and U2793 (N_2793,N_1085,N_1569);
and U2794 (N_2794,N_1054,N_1161);
nand U2795 (N_2795,N_1996,N_1787);
nor U2796 (N_2796,N_1511,N_1086);
and U2797 (N_2797,N_1396,N_1005);
nand U2798 (N_2798,N_1626,N_1208);
nor U2799 (N_2799,N_1697,N_1746);
nor U2800 (N_2800,N_1971,N_1814);
nand U2801 (N_2801,N_1110,N_1509);
nand U2802 (N_2802,N_1310,N_1529);
nor U2803 (N_2803,N_1243,N_1514);
nand U2804 (N_2804,N_1811,N_1319);
or U2805 (N_2805,N_1269,N_1845);
nor U2806 (N_2806,N_1186,N_1791);
or U2807 (N_2807,N_1567,N_1281);
and U2808 (N_2808,N_1110,N_1606);
nor U2809 (N_2809,N_1533,N_1963);
nand U2810 (N_2810,N_1015,N_1737);
or U2811 (N_2811,N_1345,N_1118);
nor U2812 (N_2812,N_1892,N_1572);
nand U2813 (N_2813,N_1938,N_1799);
or U2814 (N_2814,N_1612,N_1184);
and U2815 (N_2815,N_1033,N_1556);
and U2816 (N_2816,N_1583,N_1062);
nor U2817 (N_2817,N_1787,N_1872);
nor U2818 (N_2818,N_1153,N_1218);
nor U2819 (N_2819,N_1852,N_1965);
nand U2820 (N_2820,N_1942,N_1706);
or U2821 (N_2821,N_1474,N_1516);
and U2822 (N_2822,N_1626,N_1916);
nor U2823 (N_2823,N_1685,N_1562);
nor U2824 (N_2824,N_1528,N_1814);
or U2825 (N_2825,N_1324,N_1077);
nor U2826 (N_2826,N_1451,N_1756);
nand U2827 (N_2827,N_1158,N_1432);
nor U2828 (N_2828,N_1769,N_1361);
nand U2829 (N_2829,N_1382,N_1074);
or U2830 (N_2830,N_1498,N_1334);
or U2831 (N_2831,N_1415,N_1790);
and U2832 (N_2832,N_1917,N_1707);
or U2833 (N_2833,N_1936,N_1996);
nand U2834 (N_2834,N_1207,N_1591);
and U2835 (N_2835,N_1466,N_1227);
and U2836 (N_2836,N_1863,N_1555);
nand U2837 (N_2837,N_1195,N_1734);
xnor U2838 (N_2838,N_1937,N_1179);
nand U2839 (N_2839,N_1039,N_1302);
nand U2840 (N_2840,N_1791,N_1616);
and U2841 (N_2841,N_1722,N_1034);
or U2842 (N_2842,N_1455,N_1610);
or U2843 (N_2843,N_1253,N_1897);
or U2844 (N_2844,N_1678,N_1815);
nand U2845 (N_2845,N_1836,N_1718);
and U2846 (N_2846,N_1974,N_1422);
nand U2847 (N_2847,N_1268,N_1742);
nand U2848 (N_2848,N_1837,N_1971);
nand U2849 (N_2849,N_1215,N_1112);
nor U2850 (N_2850,N_1390,N_1075);
nand U2851 (N_2851,N_1608,N_1909);
and U2852 (N_2852,N_1496,N_1918);
nand U2853 (N_2853,N_1617,N_1584);
and U2854 (N_2854,N_1416,N_1753);
nor U2855 (N_2855,N_1573,N_1463);
and U2856 (N_2856,N_1443,N_1828);
or U2857 (N_2857,N_1337,N_1401);
nand U2858 (N_2858,N_1672,N_1778);
or U2859 (N_2859,N_1963,N_1064);
or U2860 (N_2860,N_1232,N_1517);
or U2861 (N_2861,N_1341,N_1416);
nor U2862 (N_2862,N_1061,N_1328);
nor U2863 (N_2863,N_1926,N_1920);
nand U2864 (N_2864,N_1646,N_1672);
and U2865 (N_2865,N_1670,N_1039);
nand U2866 (N_2866,N_1938,N_1557);
nor U2867 (N_2867,N_1443,N_1882);
or U2868 (N_2868,N_1670,N_1315);
nand U2869 (N_2869,N_1384,N_1318);
nor U2870 (N_2870,N_1432,N_1662);
and U2871 (N_2871,N_1463,N_1196);
or U2872 (N_2872,N_1302,N_1541);
or U2873 (N_2873,N_1832,N_1075);
nand U2874 (N_2874,N_1001,N_1277);
or U2875 (N_2875,N_1410,N_1848);
or U2876 (N_2876,N_1582,N_1344);
nand U2877 (N_2877,N_1912,N_1539);
and U2878 (N_2878,N_1703,N_1274);
nor U2879 (N_2879,N_1607,N_1944);
and U2880 (N_2880,N_1078,N_1494);
or U2881 (N_2881,N_1545,N_1749);
or U2882 (N_2882,N_1994,N_1033);
and U2883 (N_2883,N_1551,N_1326);
and U2884 (N_2884,N_1693,N_1799);
and U2885 (N_2885,N_1122,N_1003);
xnor U2886 (N_2886,N_1507,N_1657);
nor U2887 (N_2887,N_1564,N_1033);
nand U2888 (N_2888,N_1792,N_1769);
and U2889 (N_2889,N_1274,N_1103);
nor U2890 (N_2890,N_1822,N_1623);
nand U2891 (N_2891,N_1718,N_1562);
and U2892 (N_2892,N_1618,N_1276);
or U2893 (N_2893,N_1747,N_1372);
or U2894 (N_2894,N_1600,N_1190);
nand U2895 (N_2895,N_1629,N_1935);
nor U2896 (N_2896,N_1808,N_1099);
nand U2897 (N_2897,N_1658,N_1074);
and U2898 (N_2898,N_1170,N_1291);
or U2899 (N_2899,N_1001,N_1270);
or U2900 (N_2900,N_1595,N_1600);
or U2901 (N_2901,N_1507,N_1096);
and U2902 (N_2902,N_1332,N_1457);
or U2903 (N_2903,N_1407,N_1199);
or U2904 (N_2904,N_1987,N_1650);
nor U2905 (N_2905,N_1072,N_1335);
and U2906 (N_2906,N_1226,N_1840);
or U2907 (N_2907,N_1907,N_1425);
nand U2908 (N_2908,N_1226,N_1995);
nand U2909 (N_2909,N_1311,N_1852);
or U2910 (N_2910,N_1139,N_1044);
nand U2911 (N_2911,N_1328,N_1990);
and U2912 (N_2912,N_1866,N_1364);
nor U2913 (N_2913,N_1329,N_1392);
nor U2914 (N_2914,N_1248,N_1116);
nand U2915 (N_2915,N_1006,N_1248);
nor U2916 (N_2916,N_1970,N_1236);
and U2917 (N_2917,N_1152,N_1347);
and U2918 (N_2918,N_1659,N_1472);
nor U2919 (N_2919,N_1847,N_1517);
nand U2920 (N_2920,N_1805,N_1707);
or U2921 (N_2921,N_1404,N_1343);
or U2922 (N_2922,N_1786,N_1175);
and U2923 (N_2923,N_1326,N_1689);
and U2924 (N_2924,N_1908,N_1107);
nor U2925 (N_2925,N_1598,N_1696);
nor U2926 (N_2926,N_1392,N_1127);
xnor U2927 (N_2927,N_1774,N_1233);
and U2928 (N_2928,N_1065,N_1408);
or U2929 (N_2929,N_1011,N_1636);
nor U2930 (N_2930,N_1019,N_1520);
or U2931 (N_2931,N_1059,N_1241);
and U2932 (N_2932,N_1041,N_1923);
and U2933 (N_2933,N_1906,N_1626);
nand U2934 (N_2934,N_1205,N_1892);
and U2935 (N_2935,N_1746,N_1717);
nand U2936 (N_2936,N_1720,N_1380);
and U2937 (N_2937,N_1421,N_1597);
and U2938 (N_2938,N_1107,N_1993);
and U2939 (N_2939,N_1355,N_1699);
or U2940 (N_2940,N_1559,N_1605);
nand U2941 (N_2941,N_1709,N_1747);
nor U2942 (N_2942,N_1269,N_1653);
nor U2943 (N_2943,N_1307,N_1062);
or U2944 (N_2944,N_1306,N_1456);
nor U2945 (N_2945,N_1014,N_1180);
nand U2946 (N_2946,N_1513,N_1918);
nor U2947 (N_2947,N_1970,N_1697);
nand U2948 (N_2948,N_1695,N_1991);
nor U2949 (N_2949,N_1909,N_1631);
or U2950 (N_2950,N_1500,N_1669);
or U2951 (N_2951,N_1183,N_1969);
nor U2952 (N_2952,N_1883,N_1845);
or U2953 (N_2953,N_1375,N_1737);
or U2954 (N_2954,N_1096,N_1602);
nand U2955 (N_2955,N_1487,N_1552);
nand U2956 (N_2956,N_1249,N_1506);
nor U2957 (N_2957,N_1350,N_1452);
or U2958 (N_2958,N_1739,N_1923);
and U2959 (N_2959,N_1609,N_1667);
and U2960 (N_2960,N_1601,N_1504);
nor U2961 (N_2961,N_1206,N_1490);
and U2962 (N_2962,N_1127,N_1892);
nor U2963 (N_2963,N_1997,N_1222);
nor U2964 (N_2964,N_1824,N_1713);
and U2965 (N_2965,N_1060,N_1721);
and U2966 (N_2966,N_1913,N_1837);
or U2967 (N_2967,N_1229,N_1036);
or U2968 (N_2968,N_1840,N_1536);
nand U2969 (N_2969,N_1726,N_1360);
and U2970 (N_2970,N_1431,N_1303);
or U2971 (N_2971,N_1995,N_1381);
nand U2972 (N_2972,N_1882,N_1280);
and U2973 (N_2973,N_1782,N_1427);
and U2974 (N_2974,N_1538,N_1688);
and U2975 (N_2975,N_1765,N_1515);
nor U2976 (N_2976,N_1317,N_1573);
and U2977 (N_2977,N_1290,N_1994);
nand U2978 (N_2978,N_1358,N_1448);
or U2979 (N_2979,N_1162,N_1704);
and U2980 (N_2980,N_1768,N_1224);
or U2981 (N_2981,N_1014,N_1364);
nor U2982 (N_2982,N_1521,N_1459);
nor U2983 (N_2983,N_1600,N_1883);
nand U2984 (N_2984,N_1447,N_1594);
and U2985 (N_2985,N_1201,N_1182);
or U2986 (N_2986,N_1784,N_1953);
nand U2987 (N_2987,N_1820,N_1273);
and U2988 (N_2988,N_1190,N_1703);
nand U2989 (N_2989,N_1706,N_1866);
or U2990 (N_2990,N_1152,N_1687);
nand U2991 (N_2991,N_1224,N_1898);
and U2992 (N_2992,N_1224,N_1408);
and U2993 (N_2993,N_1465,N_1496);
nand U2994 (N_2994,N_1964,N_1770);
or U2995 (N_2995,N_1421,N_1944);
or U2996 (N_2996,N_1484,N_1990);
or U2997 (N_2997,N_1782,N_1656);
nor U2998 (N_2998,N_1262,N_1319);
or U2999 (N_2999,N_1039,N_1813);
or U3000 (N_3000,N_2374,N_2377);
and U3001 (N_3001,N_2217,N_2950);
nand U3002 (N_3002,N_2668,N_2077);
nor U3003 (N_3003,N_2144,N_2656);
nand U3004 (N_3004,N_2400,N_2323);
and U3005 (N_3005,N_2011,N_2650);
nor U3006 (N_3006,N_2168,N_2004);
nand U3007 (N_3007,N_2551,N_2170);
nor U3008 (N_3008,N_2878,N_2625);
xor U3009 (N_3009,N_2387,N_2651);
and U3010 (N_3010,N_2403,N_2489);
and U3011 (N_3011,N_2269,N_2791);
or U3012 (N_3012,N_2775,N_2352);
or U3013 (N_3013,N_2951,N_2568);
or U3014 (N_3014,N_2390,N_2894);
and U3015 (N_3015,N_2702,N_2541);
nand U3016 (N_3016,N_2421,N_2980);
or U3017 (N_3017,N_2443,N_2293);
nand U3018 (N_3018,N_2198,N_2175);
or U3019 (N_3019,N_2115,N_2823);
nor U3020 (N_3020,N_2076,N_2417);
nand U3021 (N_3021,N_2895,N_2666);
nand U3022 (N_3022,N_2462,N_2092);
and U3023 (N_3023,N_2189,N_2552);
and U3024 (N_3024,N_2863,N_2550);
nand U3025 (N_3025,N_2407,N_2978);
or U3026 (N_3026,N_2506,N_2670);
or U3027 (N_3027,N_2799,N_2086);
nor U3028 (N_3028,N_2990,N_2467);
and U3029 (N_3029,N_2380,N_2735);
and U3030 (N_3030,N_2594,N_2820);
or U3031 (N_3031,N_2697,N_2674);
nor U3032 (N_3032,N_2662,N_2285);
or U3033 (N_3033,N_2491,N_2796);
and U3034 (N_3034,N_2910,N_2525);
and U3035 (N_3035,N_2185,N_2871);
nor U3036 (N_3036,N_2671,N_2391);
or U3037 (N_3037,N_2729,N_2898);
and U3038 (N_3038,N_2954,N_2437);
nor U3039 (N_3039,N_2628,N_2381);
and U3040 (N_3040,N_2335,N_2104);
and U3041 (N_3041,N_2184,N_2366);
nor U3042 (N_3042,N_2777,N_2100);
nand U3043 (N_3043,N_2485,N_2250);
or U3044 (N_3044,N_2635,N_2499);
or U3045 (N_3045,N_2096,N_2789);
or U3046 (N_3046,N_2722,N_2794);
nand U3047 (N_3047,N_2340,N_2152);
and U3048 (N_3048,N_2923,N_2606);
or U3049 (N_3049,N_2422,N_2030);
nand U3050 (N_3050,N_2345,N_2476);
nand U3051 (N_3051,N_2306,N_2002);
nand U3052 (N_3052,N_2474,N_2557);
nand U3053 (N_3053,N_2042,N_2637);
and U3054 (N_3054,N_2725,N_2734);
or U3055 (N_3055,N_2605,N_2431);
nand U3056 (N_3056,N_2194,N_2530);
nor U3057 (N_3057,N_2800,N_2051);
or U3058 (N_3058,N_2012,N_2532);
or U3059 (N_3059,N_2483,N_2511);
nor U3060 (N_3060,N_2498,N_2522);
and U3061 (N_3061,N_2825,N_2634);
nand U3062 (N_3062,N_2717,N_2669);
nand U3063 (N_3063,N_2037,N_2101);
and U3064 (N_3064,N_2533,N_2346);
or U3065 (N_3065,N_2221,N_2079);
or U3066 (N_3066,N_2319,N_2049);
nor U3067 (N_3067,N_2881,N_2755);
and U3068 (N_3068,N_2518,N_2035);
nor U3069 (N_3069,N_2317,N_2428);
and U3070 (N_3070,N_2276,N_2015);
nand U3071 (N_3071,N_2828,N_2583);
nor U3072 (N_3072,N_2700,N_2942);
and U3073 (N_3073,N_2266,N_2413);
or U3074 (N_3074,N_2703,N_2418);
and U3075 (N_3075,N_2062,N_2438);
nand U3076 (N_3076,N_2989,N_2386);
nor U3077 (N_3077,N_2385,N_2563);
and U3078 (N_3078,N_2404,N_2248);
nor U3079 (N_3079,N_2075,N_2844);
xnor U3080 (N_3080,N_2135,N_2369);
or U3081 (N_3081,N_2507,N_2621);
nand U3082 (N_3082,N_2764,N_2026);
and U3083 (N_3083,N_2225,N_2274);
nor U3084 (N_3084,N_2003,N_2624);
nor U3085 (N_3085,N_2497,N_2016);
nand U3086 (N_3086,N_2932,N_2208);
nand U3087 (N_3087,N_2553,N_2398);
and U3088 (N_3088,N_2861,N_2787);
nand U3089 (N_3089,N_2239,N_2173);
or U3090 (N_3090,N_2257,N_2840);
and U3091 (N_3091,N_2542,N_2087);
nor U3092 (N_3092,N_2287,N_2920);
nor U3093 (N_3093,N_2432,N_2569);
or U3094 (N_3094,N_2401,N_2653);
or U3095 (N_3095,N_2707,N_2986);
and U3096 (N_3096,N_2639,N_2988);
or U3097 (N_3097,N_2661,N_2744);
and U3098 (N_3098,N_2054,N_2929);
or U3099 (N_3099,N_2236,N_2575);
nor U3100 (N_3100,N_2596,N_2275);
or U3101 (N_3101,N_2307,N_2685);
and U3102 (N_3102,N_2433,N_2640);
nor U3103 (N_3103,N_2000,N_2351);
and U3104 (N_3104,N_2905,N_2372);
nor U3105 (N_3105,N_2140,N_2448);
nand U3106 (N_3106,N_2979,N_2113);
nor U3107 (N_3107,N_2399,N_2893);
nor U3108 (N_3108,N_2290,N_2122);
xor U3109 (N_3109,N_2995,N_2009);
or U3110 (N_3110,N_2921,N_2589);
or U3111 (N_3111,N_2342,N_2870);
nand U3112 (N_3112,N_2373,N_2544);
or U3113 (N_3113,N_2367,N_2570);
nor U3114 (N_3114,N_2021,N_2998);
nand U3115 (N_3115,N_2136,N_2604);
or U3116 (N_3116,N_2996,N_2089);
nor U3117 (N_3117,N_2383,N_2419);
and U3118 (N_3118,N_2658,N_2592);
nand U3119 (N_3119,N_2028,N_2769);
nand U3120 (N_3120,N_2244,N_2896);
nand U3121 (N_3121,N_2712,N_2254);
nor U3122 (N_3122,N_2412,N_2649);
or U3123 (N_3123,N_2526,N_2962);
nand U3124 (N_3124,N_2022,N_2229);
nand U3125 (N_3125,N_2333,N_2698);
nand U3126 (N_3126,N_2129,N_2065);
nand U3127 (N_3127,N_2607,N_2316);
xnor U3128 (N_3128,N_2363,N_2311);
xnor U3129 (N_3129,N_2180,N_2106);
nand U3130 (N_3130,N_2176,N_2629);
or U3131 (N_3131,N_2482,N_2167);
nor U3132 (N_3132,N_2536,N_2534);
nand U3133 (N_3133,N_2681,N_2865);
nor U3134 (N_3134,N_2687,N_2574);
and U3135 (N_3135,N_2601,N_2975);
nand U3136 (N_3136,N_2020,N_2732);
nand U3137 (N_3137,N_2852,N_2321);
nor U3138 (N_3138,N_2141,N_2660);
nor U3139 (N_3139,N_2093,N_2528);
nand U3140 (N_3140,N_2127,N_2832);
or U3141 (N_3141,N_2750,N_2636);
nor U3142 (N_3142,N_2328,N_2466);
nand U3143 (N_3143,N_2108,N_2918);
nor U3144 (N_3144,N_2235,N_2361);
nand U3145 (N_3145,N_2934,N_2281);
and U3146 (N_3146,N_2183,N_2156);
nor U3147 (N_3147,N_2255,N_2118);
and U3148 (N_3148,N_2810,N_2925);
nand U3149 (N_3149,N_2326,N_2468);
or U3150 (N_3150,N_2405,N_2416);
and U3151 (N_3151,N_2831,N_2347);
or U3152 (N_3152,N_2580,N_2784);
or U3153 (N_3153,N_2465,N_2222);
nor U3154 (N_3154,N_2676,N_2296);
or U3155 (N_3155,N_2237,N_2360);
and U3156 (N_3156,N_2973,N_2720);
and U3157 (N_3157,N_2056,N_2778);
and U3158 (N_3158,N_2642,N_2402);
and U3159 (N_3159,N_2726,N_2821);
or U3160 (N_3160,N_2904,N_2450);
and U3161 (N_3161,N_2776,N_2880);
and U3162 (N_3162,N_2916,N_2758);
and U3163 (N_3163,N_2415,N_2302);
nand U3164 (N_3164,N_2699,N_2159);
and U3165 (N_3165,N_2546,N_2472);
xor U3166 (N_3166,N_2588,N_2627);
or U3167 (N_3167,N_2036,N_2782);
and U3168 (N_3168,N_2259,N_2233);
or U3169 (N_3169,N_2851,N_2610);
or U3170 (N_3170,N_2731,N_2907);
or U3171 (N_3171,N_2139,N_2046);
or U3172 (N_3172,N_2434,N_2945);
nand U3173 (N_3173,N_2130,N_2102);
xor U3174 (N_3174,N_2953,N_2967);
nand U3175 (N_3175,N_2862,N_2795);
nand U3176 (N_3176,N_2256,N_2430);
and U3177 (N_3177,N_2488,N_2158);
and U3178 (N_3178,N_2358,N_2204);
and U3179 (N_3179,N_2696,N_2460);
nor U3180 (N_3180,N_2667,N_2368);
and U3181 (N_3181,N_2120,N_2082);
or U3182 (N_3182,N_2423,N_2454);
and U3183 (N_3183,N_2767,N_2278);
xnor U3184 (N_3184,N_2309,N_2449);
nor U3185 (N_3185,N_2252,N_2126);
or U3186 (N_3186,N_2853,N_2154);
and U3187 (N_3187,N_2869,N_2582);
nand U3188 (N_3188,N_2470,N_2587);
nor U3189 (N_3189,N_2344,N_2301);
or U3190 (N_3190,N_2559,N_2691);
and U3191 (N_3191,N_2492,N_2043);
nor U3192 (N_3192,N_2505,N_2494);
and U3193 (N_3193,N_2091,N_2609);
nor U3194 (N_3194,N_2191,N_2850);
nand U3195 (N_3195,N_2859,N_2960);
and U3196 (N_3196,N_2745,N_2458);
and U3197 (N_3197,N_2786,N_2188);
and U3198 (N_3198,N_2708,N_2477);
and U3199 (N_3199,N_2186,N_2187);
nor U3200 (N_3200,N_2740,N_2811);
and U3201 (N_3201,N_2562,N_2213);
nand U3202 (N_3202,N_2531,N_2284);
nor U3203 (N_3203,N_2214,N_2375);
nor U3204 (N_3204,N_2827,N_2919);
nand U3205 (N_3205,N_2064,N_2959);
nor U3206 (N_3206,N_2496,N_2109);
or U3207 (N_3207,N_2084,N_2924);
xor U3208 (N_3208,N_2199,N_2288);
and U3209 (N_3209,N_2339,N_2913);
or U3210 (N_3210,N_2648,N_2812);
nor U3211 (N_3211,N_2085,N_2614);
nand U3212 (N_3212,N_2618,N_2993);
or U3213 (N_3213,N_2713,N_2890);
nor U3214 (N_3214,N_2451,N_2909);
nor U3215 (N_3215,N_2163,N_2888);
nor U3216 (N_3216,N_2055,N_2090);
or U3217 (N_3217,N_2209,N_2985);
nor U3218 (N_3218,N_2877,N_2216);
nor U3219 (N_3219,N_2930,N_2195);
or U3220 (N_3220,N_2479,N_2142);
nand U3221 (N_3221,N_2078,N_2882);
and U3222 (N_3222,N_2539,N_2463);
and U3223 (N_3223,N_2974,N_2689);
or U3224 (N_3224,N_2389,N_2561);
or U3225 (N_3225,N_2071,N_2972);
or U3226 (N_3226,N_2410,N_2040);
nor U3227 (N_3227,N_2297,N_2107);
or U3228 (N_3228,N_2314,N_2220);
nor U3229 (N_3229,N_2267,N_2982);
or U3230 (N_3230,N_2873,N_2709);
and U3231 (N_3231,N_2409,N_2517);
nand U3232 (N_3232,N_2718,N_2420);
nand U3233 (N_3233,N_2804,N_2271);
or U3234 (N_3234,N_2193,N_2073);
and U3235 (N_3235,N_2747,N_2338);
or U3236 (N_3236,N_2631,N_2359);
nor U3237 (N_3237,N_2817,N_2956);
nand U3238 (N_3238,N_2138,N_2590);
nor U3239 (N_3239,N_2652,N_2058);
and U3240 (N_3240,N_2567,N_2081);
and U3241 (N_3241,N_2223,N_2875);
or U3242 (N_3242,N_2461,N_2860);
nor U3243 (N_3243,N_2886,N_2663);
nor U3244 (N_3244,N_2439,N_2232);
nand U3245 (N_3245,N_2008,N_2838);
and U3246 (N_3246,N_2349,N_2478);
and U3247 (N_3247,N_2889,N_2149);
and U3248 (N_3248,N_2608,N_2356);
nand U3249 (N_3249,N_2493,N_2839);
or U3250 (N_3250,N_2645,N_2282);
or U3251 (N_3251,N_2125,N_2200);
nand U3252 (N_3252,N_2514,N_2900);
nor U3253 (N_3253,N_2510,N_2277);
nor U3254 (N_3254,N_2211,N_2023);
nand U3255 (N_3255,N_2955,N_2068);
nand U3256 (N_3256,N_2080,N_2445);
nand U3257 (N_3257,N_2251,N_2917);
and U3258 (N_3258,N_2751,N_2947);
or U3259 (N_3259,N_2205,N_2384);
and U3260 (N_3260,N_2411,N_2694);
nand U3261 (N_3261,N_2834,N_2521);
and U3262 (N_3262,N_2683,N_2396);
nand U3263 (N_3263,N_2513,N_2746);
nor U3264 (N_3264,N_2543,N_2704);
nor U3265 (N_3265,N_2006,N_2031);
nand U3266 (N_3266,N_2155,N_2981);
nand U3267 (N_3267,N_2868,N_2774);
and U3268 (N_3268,N_2987,N_2805);
nand U3269 (N_3269,N_2201,N_2171);
nand U3270 (N_3270,N_2435,N_2964);
nor U3271 (N_3271,N_2772,N_2265);
nor U3272 (N_3272,N_2727,N_2595);
or U3273 (N_3273,N_2944,N_2573);
and U3274 (N_3274,N_2710,N_2464);
nor U3275 (N_3275,N_2885,N_2379);
or U3276 (N_3276,N_2591,N_2884);
nand U3277 (N_3277,N_2847,N_2766);
and U3278 (N_3278,N_2447,N_2858);
nor U3279 (N_3279,N_2382,N_2779);
nand U3280 (N_3280,N_2957,N_2938);
and U3281 (N_3281,N_2145,N_2655);
or U3282 (N_3282,N_2295,N_2586);
or U3283 (N_3283,N_2341,N_2711);
or U3284 (N_3284,N_2516,N_2593);
and U3285 (N_3285,N_2728,N_2688);
nor U3286 (N_3286,N_2057,N_2270);
and U3287 (N_3287,N_2792,N_2902);
nand U3288 (N_3288,N_2647,N_2952);
nand U3289 (N_3289,N_2315,N_2268);
or U3290 (N_3290,N_2939,N_2114);
nor U3291 (N_3291,N_2376,N_2822);
nor U3292 (N_3292,N_2406,N_2181);
or U3293 (N_3293,N_2025,N_2121);
nand U3294 (N_3294,N_2897,N_2312);
nor U3295 (N_3295,N_2684,N_2749);
nor U3296 (N_3296,N_2283,N_2219);
or U3297 (N_3297,N_2809,N_2842);
nand U3298 (N_3298,N_2240,N_2322);
or U3299 (N_3299,N_2041,N_2701);
or U3300 (N_3300,N_2739,N_2619);
or U3301 (N_3301,N_2061,N_2940);
nor U3302 (N_3302,N_2337,N_2835);
nor U3303 (N_3303,N_2414,N_2680);
nand U3304 (N_3304,N_2949,N_2612);
and U3305 (N_3305,N_2289,N_2304);
or U3306 (N_3306,N_2992,N_2197);
nand U3307 (N_3307,N_2754,N_2446);
and U3308 (N_3308,N_2034,N_2578);
nand U3309 (N_3309,N_2598,N_2833);
nand U3310 (N_3310,N_2849,N_2966);
and U3311 (N_3311,N_2300,N_2816);
nand U3312 (N_3312,N_2741,N_2846);
nor U3313 (N_3313,N_2001,N_2500);
nand U3314 (N_3314,N_2440,N_2620);
nand U3315 (N_3315,N_2693,N_2394);
nand U3316 (N_3316,N_2753,N_2370);
nand U3317 (N_3317,N_2160,N_2018);
nand U3318 (N_3318,N_2164,N_2050);
or U3319 (N_3319,N_2174,N_2558);
nor U3320 (N_3320,N_2556,N_2124);
or U3321 (N_3321,N_2010,N_2581);
nor U3322 (N_3322,N_2502,N_2752);
nor U3323 (N_3323,N_2742,N_2958);
nor U3324 (N_3324,N_2123,N_2308);
nand U3325 (N_3325,N_2203,N_2576);
nor U3326 (N_3326,N_2157,N_2501);
and U3327 (N_3327,N_2272,N_2017);
and U3328 (N_3328,N_2357,N_2935);
or U3329 (N_3329,N_2686,N_2524);
or U3330 (N_3330,N_2790,N_2768);
or U3331 (N_3331,N_2603,N_2294);
nor U3332 (N_3332,N_2117,N_2819);
nand U3333 (N_3333,N_2705,N_2879);
or U3334 (N_3334,N_2161,N_2657);
nor U3335 (N_3335,N_2549,N_2179);
or U3336 (N_3336,N_2914,N_2095);
and U3337 (N_3337,N_2318,N_2814);
nor U3338 (N_3338,N_2146,N_2325);
nor U3339 (N_3339,N_2748,N_2780);
and U3340 (N_3340,N_2585,N_2429);
and U3341 (N_3341,N_2737,N_2757);
and U3342 (N_3342,N_2436,N_2560);
nand U3343 (N_3343,N_2310,N_2977);
or U3344 (N_3344,N_2716,N_2867);
nor U3345 (N_3345,N_2444,N_2110);
nand U3346 (N_3346,N_2353,N_2013);
or U3347 (N_3347,N_2706,N_2103);
or U3348 (N_3348,N_2969,N_2999);
or U3349 (N_3349,N_2623,N_2024);
nor U3350 (N_3350,N_2630,N_2857);
nor U3351 (N_3351,N_2770,N_2971);
or U3352 (N_3352,N_2088,N_2983);
or U3353 (N_3353,N_2646,N_2946);
nand U3354 (N_3354,N_2364,N_2771);
and U3355 (N_3355,N_2169,N_2843);
nand U3356 (N_3356,N_2230,N_2509);
nand U3357 (N_3357,N_2218,N_2459);
or U3358 (N_3358,N_2441,N_2943);
nand U3359 (N_3359,N_2392,N_2961);
and U3360 (N_3360,N_2053,N_2371);
nor U3361 (N_3361,N_2094,N_2519);
nor U3362 (N_3362,N_2298,N_2690);
and U3363 (N_3363,N_2622,N_2565);
and U3364 (N_3364,N_2566,N_2597);
nand U3365 (N_3365,N_2785,N_2119);
and U3366 (N_3366,N_2926,N_2872);
or U3367 (N_3367,N_2190,N_2329);
or U3368 (N_3368,N_2452,N_2249);
nor U3369 (N_3369,N_2664,N_2234);
nand U3370 (N_3370,N_2486,N_2207);
nand U3371 (N_3371,N_2348,N_2602);
nand U3372 (N_3372,N_2343,N_2279);
and U3373 (N_3373,N_2759,N_2836);
nand U3374 (N_3374,N_2762,N_2891);
or U3375 (N_3375,N_2480,N_2291);
nand U3376 (N_3376,N_2273,N_2111);
nand U3377 (N_3377,N_2245,N_2783);
nor U3378 (N_3378,N_2241,N_2427);
nor U3379 (N_3379,N_2854,N_2965);
or U3380 (N_3380,N_2131,N_2455);
nand U3381 (N_3381,N_2679,N_2143);
and U3382 (N_3382,N_2571,N_2538);
nor U3383 (N_3383,N_2292,N_2876);
nand U3384 (N_3384,N_2948,N_2334);
or U3385 (N_3385,N_2147,N_2045);
or U3386 (N_3386,N_2997,N_2231);
and U3387 (N_3387,N_2641,N_2616);
nand U3388 (N_3388,N_2763,N_2927);
or U3389 (N_3389,N_2063,N_2931);
nor U3390 (N_3390,N_2572,N_2243);
nor U3391 (N_3391,N_2584,N_2069);
nor U3392 (N_3392,N_2453,N_2765);
and U3393 (N_3393,N_2378,N_2475);
and U3394 (N_3394,N_2247,N_2678);
or U3395 (N_3395,N_2903,N_2970);
and U3396 (N_3396,N_2912,N_2781);
or U3397 (N_3397,N_2365,N_2756);
nand U3398 (N_3398,N_2611,N_2354);
nand U3399 (N_3399,N_2677,N_2537);
or U3400 (N_3400,N_2826,N_2866);
and U3401 (N_3401,N_2724,N_2901);
nand U3402 (N_3402,N_2038,N_2504);
nand U3403 (N_3403,N_2261,N_2801);
or U3404 (N_3404,N_2215,N_2773);
nor U3405 (N_3405,N_2665,N_2803);
xnor U3406 (N_3406,N_2227,N_2264);
and U3407 (N_3407,N_2471,N_2099);
or U3408 (N_3408,N_2824,N_2074);
nand U3409 (N_3409,N_2760,N_2070);
and U3410 (N_3410,N_2761,N_2808);
or U3411 (N_3411,N_2564,N_2617);
nor U3412 (N_3412,N_2523,N_2719);
or U3413 (N_3413,N_2172,N_2928);
nor U3414 (N_3414,N_2991,N_2856);
or U3415 (N_3415,N_2736,N_2487);
or U3416 (N_3416,N_2490,N_2330);
and U3417 (N_3417,N_2675,N_2484);
nor U3418 (N_3418,N_2128,N_2029);
and U3419 (N_3419,N_2798,N_2738);
and U3420 (N_3420,N_2848,N_2224);
and U3421 (N_3421,N_2915,N_2133);
nand U3422 (N_3422,N_2473,N_2730);
nor U3423 (N_3423,N_2829,N_2554);
nand U3424 (N_3424,N_2841,N_2280);
or U3425 (N_3425,N_2112,N_2864);
nor U3426 (N_3426,N_2132,N_2540);
nand U3427 (N_3427,N_2545,N_2052);
and U3428 (N_3428,N_2815,N_2984);
and U3429 (N_3429,N_2469,N_2350);
nand U3430 (N_3430,N_2723,N_2097);
nor U3431 (N_3431,N_2395,N_2892);
nor U3432 (N_3432,N_2263,N_2246);
or U3433 (N_3433,N_2626,N_2908);
nor U3434 (N_3434,N_2615,N_2408);
and U3435 (N_3435,N_2260,N_2941);
or U3436 (N_3436,N_2495,N_2633);
nor U3437 (N_3437,N_2936,N_2242);
nor U3438 (N_3438,N_2555,N_2442);
and U3439 (N_3439,N_2134,N_2512);
nor U3440 (N_3440,N_2212,N_2855);
nand U3441 (N_3441,N_2994,N_2547);
nor U3442 (N_3442,N_2067,N_2238);
nand U3443 (N_3443,N_2072,N_2032);
and U3444 (N_3444,N_2048,N_2425);
nor U3445 (N_3445,N_2286,N_2643);
or U3446 (N_3446,N_2911,N_2715);
nand U3447 (N_3447,N_2039,N_2105);
or U3448 (N_3448,N_2393,N_2520);
or U3449 (N_3449,N_2210,N_2743);
or U3450 (N_3450,N_2151,N_2424);
nor U3451 (N_3451,N_2638,N_2083);
or U3452 (N_3452,N_2682,N_2793);
nor U3453 (N_3453,N_2253,N_2883);
and U3454 (N_3454,N_2226,N_2033);
nor U3455 (N_3455,N_2692,N_2673);
and U3456 (N_3456,N_2327,N_2116);
nor U3457 (N_3457,N_2515,N_2874);
nor U3458 (N_3458,N_2019,N_2922);
and U3459 (N_3459,N_2299,N_2202);
nor U3460 (N_3460,N_2906,N_2837);
nor U3461 (N_3461,N_2005,N_2137);
nand U3462 (N_3462,N_2066,N_2027);
nor U3463 (N_3463,N_2899,N_2654);
nor U3464 (N_3464,N_2426,N_2228);
nand U3465 (N_3465,N_2044,N_2887);
nor U3466 (N_3466,N_2481,N_2508);
nor U3467 (N_3467,N_2320,N_2192);
and U3468 (N_3468,N_2457,N_2007);
and U3469 (N_3469,N_2178,N_2599);
or U3470 (N_3470,N_2659,N_2830);
or U3471 (N_3471,N_2177,N_2721);
and U3472 (N_3472,N_2548,N_2845);
and U3473 (N_3473,N_2672,N_2060);
nor U3474 (N_3474,N_2355,N_2262);
and U3475 (N_3475,N_2047,N_2529);
and U3476 (N_3476,N_2332,N_2362);
or U3477 (N_3477,N_2976,N_2331);
and U3478 (N_3478,N_2695,N_2162);
nor U3479 (N_3479,N_2336,N_2806);
or U3480 (N_3480,N_2098,N_2182);
nand U3481 (N_3481,N_2324,N_2014);
nor U3482 (N_3482,N_2963,N_2305);
nor U3483 (N_3483,N_2797,N_2968);
or U3484 (N_3484,N_2313,N_2733);
and U3485 (N_3485,N_2527,N_2714);
nand U3486 (N_3486,N_2788,N_2802);
and U3487 (N_3487,N_2937,N_2600);
and U3488 (N_3488,N_2206,N_2613);
or U3489 (N_3489,N_2150,N_2148);
and U3490 (N_3490,N_2303,N_2933);
nand U3491 (N_3491,N_2807,N_2397);
nand U3492 (N_3492,N_2644,N_2535);
or U3493 (N_3493,N_2165,N_2813);
and U3494 (N_3494,N_2196,N_2153);
and U3495 (N_3495,N_2632,N_2059);
and U3496 (N_3496,N_2579,N_2818);
nor U3497 (N_3497,N_2258,N_2577);
nand U3498 (N_3498,N_2456,N_2388);
and U3499 (N_3499,N_2503,N_2166);
nor U3500 (N_3500,N_2534,N_2913);
or U3501 (N_3501,N_2521,N_2849);
nor U3502 (N_3502,N_2183,N_2953);
or U3503 (N_3503,N_2723,N_2225);
nand U3504 (N_3504,N_2418,N_2210);
nor U3505 (N_3505,N_2972,N_2509);
and U3506 (N_3506,N_2596,N_2481);
and U3507 (N_3507,N_2727,N_2867);
and U3508 (N_3508,N_2659,N_2917);
nand U3509 (N_3509,N_2938,N_2670);
or U3510 (N_3510,N_2499,N_2426);
nor U3511 (N_3511,N_2736,N_2032);
nand U3512 (N_3512,N_2700,N_2546);
and U3513 (N_3513,N_2188,N_2121);
nand U3514 (N_3514,N_2925,N_2204);
nand U3515 (N_3515,N_2338,N_2065);
nor U3516 (N_3516,N_2952,N_2207);
or U3517 (N_3517,N_2579,N_2668);
nor U3518 (N_3518,N_2940,N_2695);
or U3519 (N_3519,N_2076,N_2058);
nand U3520 (N_3520,N_2828,N_2431);
and U3521 (N_3521,N_2379,N_2509);
nor U3522 (N_3522,N_2667,N_2030);
nand U3523 (N_3523,N_2605,N_2461);
xor U3524 (N_3524,N_2643,N_2737);
or U3525 (N_3525,N_2943,N_2226);
or U3526 (N_3526,N_2944,N_2775);
and U3527 (N_3527,N_2235,N_2569);
nand U3528 (N_3528,N_2583,N_2920);
nand U3529 (N_3529,N_2521,N_2505);
nor U3530 (N_3530,N_2734,N_2208);
and U3531 (N_3531,N_2275,N_2713);
nand U3532 (N_3532,N_2836,N_2755);
nor U3533 (N_3533,N_2175,N_2072);
xor U3534 (N_3534,N_2610,N_2142);
and U3535 (N_3535,N_2596,N_2723);
or U3536 (N_3536,N_2850,N_2863);
and U3537 (N_3537,N_2682,N_2184);
nor U3538 (N_3538,N_2708,N_2551);
or U3539 (N_3539,N_2704,N_2980);
or U3540 (N_3540,N_2622,N_2566);
nor U3541 (N_3541,N_2818,N_2541);
nand U3542 (N_3542,N_2554,N_2661);
and U3543 (N_3543,N_2987,N_2712);
or U3544 (N_3544,N_2847,N_2905);
or U3545 (N_3545,N_2079,N_2782);
nand U3546 (N_3546,N_2469,N_2203);
nor U3547 (N_3547,N_2052,N_2135);
nor U3548 (N_3548,N_2400,N_2150);
and U3549 (N_3549,N_2575,N_2424);
nand U3550 (N_3550,N_2010,N_2937);
or U3551 (N_3551,N_2322,N_2267);
nor U3552 (N_3552,N_2126,N_2611);
or U3553 (N_3553,N_2758,N_2718);
or U3554 (N_3554,N_2913,N_2161);
and U3555 (N_3555,N_2000,N_2892);
or U3556 (N_3556,N_2115,N_2409);
nor U3557 (N_3557,N_2657,N_2475);
nand U3558 (N_3558,N_2931,N_2844);
nor U3559 (N_3559,N_2081,N_2951);
nor U3560 (N_3560,N_2591,N_2925);
or U3561 (N_3561,N_2999,N_2610);
and U3562 (N_3562,N_2110,N_2649);
and U3563 (N_3563,N_2914,N_2501);
and U3564 (N_3564,N_2426,N_2861);
nand U3565 (N_3565,N_2834,N_2209);
or U3566 (N_3566,N_2058,N_2985);
nand U3567 (N_3567,N_2983,N_2682);
nand U3568 (N_3568,N_2467,N_2317);
and U3569 (N_3569,N_2704,N_2626);
or U3570 (N_3570,N_2254,N_2741);
and U3571 (N_3571,N_2483,N_2635);
or U3572 (N_3572,N_2752,N_2256);
nor U3573 (N_3573,N_2256,N_2810);
and U3574 (N_3574,N_2559,N_2142);
nor U3575 (N_3575,N_2544,N_2102);
and U3576 (N_3576,N_2988,N_2209);
nor U3577 (N_3577,N_2120,N_2996);
or U3578 (N_3578,N_2080,N_2041);
and U3579 (N_3579,N_2702,N_2636);
nand U3580 (N_3580,N_2668,N_2004);
nand U3581 (N_3581,N_2757,N_2416);
nor U3582 (N_3582,N_2673,N_2909);
nor U3583 (N_3583,N_2450,N_2752);
or U3584 (N_3584,N_2062,N_2641);
nor U3585 (N_3585,N_2852,N_2402);
and U3586 (N_3586,N_2218,N_2971);
or U3587 (N_3587,N_2767,N_2609);
and U3588 (N_3588,N_2954,N_2782);
nor U3589 (N_3589,N_2271,N_2721);
nand U3590 (N_3590,N_2894,N_2904);
nand U3591 (N_3591,N_2295,N_2171);
nand U3592 (N_3592,N_2045,N_2482);
and U3593 (N_3593,N_2736,N_2296);
and U3594 (N_3594,N_2077,N_2430);
nor U3595 (N_3595,N_2244,N_2021);
and U3596 (N_3596,N_2974,N_2675);
and U3597 (N_3597,N_2633,N_2757);
or U3598 (N_3598,N_2117,N_2717);
nand U3599 (N_3599,N_2395,N_2806);
nand U3600 (N_3600,N_2700,N_2782);
nand U3601 (N_3601,N_2149,N_2334);
nand U3602 (N_3602,N_2679,N_2272);
and U3603 (N_3603,N_2095,N_2096);
or U3604 (N_3604,N_2243,N_2399);
and U3605 (N_3605,N_2317,N_2662);
and U3606 (N_3606,N_2400,N_2408);
and U3607 (N_3607,N_2179,N_2199);
or U3608 (N_3608,N_2100,N_2547);
or U3609 (N_3609,N_2776,N_2658);
nor U3610 (N_3610,N_2345,N_2821);
nor U3611 (N_3611,N_2536,N_2157);
nand U3612 (N_3612,N_2263,N_2270);
or U3613 (N_3613,N_2657,N_2116);
and U3614 (N_3614,N_2887,N_2673);
nor U3615 (N_3615,N_2927,N_2364);
or U3616 (N_3616,N_2065,N_2269);
nand U3617 (N_3617,N_2213,N_2054);
nand U3618 (N_3618,N_2066,N_2090);
xor U3619 (N_3619,N_2804,N_2639);
and U3620 (N_3620,N_2584,N_2680);
and U3621 (N_3621,N_2571,N_2918);
and U3622 (N_3622,N_2910,N_2814);
nor U3623 (N_3623,N_2693,N_2011);
nand U3624 (N_3624,N_2842,N_2399);
or U3625 (N_3625,N_2039,N_2366);
and U3626 (N_3626,N_2813,N_2763);
nand U3627 (N_3627,N_2599,N_2888);
nand U3628 (N_3628,N_2769,N_2709);
or U3629 (N_3629,N_2021,N_2803);
nand U3630 (N_3630,N_2092,N_2178);
and U3631 (N_3631,N_2187,N_2638);
or U3632 (N_3632,N_2592,N_2851);
or U3633 (N_3633,N_2719,N_2542);
or U3634 (N_3634,N_2394,N_2579);
and U3635 (N_3635,N_2405,N_2852);
and U3636 (N_3636,N_2080,N_2889);
nor U3637 (N_3637,N_2678,N_2175);
nand U3638 (N_3638,N_2842,N_2447);
and U3639 (N_3639,N_2760,N_2022);
xnor U3640 (N_3640,N_2712,N_2681);
nand U3641 (N_3641,N_2878,N_2994);
or U3642 (N_3642,N_2116,N_2345);
nor U3643 (N_3643,N_2899,N_2770);
or U3644 (N_3644,N_2943,N_2426);
or U3645 (N_3645,N_2467,N_2508);
nand U3646 (N_3646,N_2194,N_2630);
or U3647 (N_3647,N_2035,N_2848);
or U3648 (N_3648,N_2955,N_2924);
and U3649 (N_3649,N_2142,N_2373);
nor U3650 (N_3650,N_2106,N_2350);
or U3651 (N_3651,N_2685,N_2116);
nor U3652 (N_3652,N_2078,N_2736);
and U3653 (N_3653,N_2282,N_2082);
or U3654 (N_3654,N_2009,N_2558);
and U3655 (N_3655,N_2792,N_2372);
nand U3656 (N_3656,N_2338,N_2034);
nand U3657 (N_3657,N_2366,N_2514);
or U3658 (N_3658,N_2525,N_2701);
nor U3659 (N_3659,N_2931,N_2756);
nor U3660 (N_3660,N_2477,N_2178);
nor U3661 (N_3661,N_2596,N_2931);
nor U3662 (N_3662,N_2309,N_2530);
nand U3663 (N_3663,N_2994,N_2222);
nand U3664 (N_3664,N_2364,N_2414);
or U3665 (N_3665,N_2433,N_2414);
or U3666 (N_3666,N_2211,N_2798);
nor U3667 (N_3667,N_2790,N_2908);
and U3668 (N_3668,N_2308,N_2488);
nor U3669 (N_3669,N_2489,N_2233);
nor U3670 (N_3670,N_2659,N_2150);
nor U3671 (N_3671,N_2792,N_2130);
xnor U3672 (N_3672,N_2443,N_2212);
nor U3673 (N_3673,N_2973,N_2486);
and U3674 (N_3674,N_2684,N_2269);
nor U3675 (N_3675,N_2226,N_2790);
and U3676 (N_3676,N_2079,N_2038);
nor U3677 (N_3677,N_2090,N_2103);
nand U3678 (N_3678,N_2878,N_2009);
nor U3679 (N_3679,N_2774,N_2730);
and U3680 (N_3680,N_2595,N_2709);
nand U3681 (N_3681,N_2818,N_2524);
or U3682 (N_3682,N_2654,N_2619);
nor U3683 (N_3683,N_2587,N_2681);
nor U3684 (N_3684,N_2750,N_2967);
nor U3685 (N_3685,N_2480,N_2598);
or U3686 (N_3686,N_2827,N_2200);
or U3687 (N_3687,N_2710,N_2286);
or U3688 (N_3688,N_2735,N_2368);
nor U3689 (N_3689,N_2787,N_2203);
nand U3690 (N_3690,N_2464,N_2923);
nand U3691 (N_3691,N_2433,N_2794);
or U3692 (N_3692,N_2957,N_2345);
or U3693 (N_3693,N_2738,N_2810);
nand U3694 (N_3694,N_2401,N_2559);
nor U3695 (N_3695,N_2086,N_2202);
and U3696 (N_3696,N_2684,N_2733);
and U3697 (N_3697,N_2865,N_2329);
nor U3698 (N_3698,N_2121,N_2336);
and U3699 (N_3699,N_2336,N_2739);
nand U3700 (N_3700,N_2892,N_2535);
and U3701 (N_3701,N_2143,N_2397);
nor U3702 (N_3702,N_2081,N_2245);
and U3703 (N_3703,N_2135,N_2837);
nor U3704 (N_3704,N_2532,N_2656);
nor U3705 (N_3705,N_2343,N_2589);
and U3706 (N_3706,N_2443,N_2154);
and U3707 (N_3707,N_2146,N_2647);
nor U3708 (N_3708,N_2046,N_2890);
nor U3709 (N_3709,N_2407,N_2664);
nor U3710 (N_3710,N_2498,N_2061);
or U3711 (N_3711,N_2591,N_2855);
xnor U3712 (N_3712,N_2378,N_2796);
and U3713 (N_3713,N_2733,N_2366);
nand U3714 (N_3714,N_2048,N_2412);
nand U3715 (N_3715,N_2146,N_2339);
nor U3716 (N_3716,N_2224,N_2334);
nand U3717 (N_3717,N_2824,N_2795);
and U3718 (N_3718,N_2676,N_2608);
xnor U3719 (N_3719,N_2958,N_2147);
or U3720 (N_3720,N_2155,N_2948);
xor U3721 (N_3721,N_2168,N_2536);
and U3722 (N_3722,N_2276,N_2609);
and U3723 (N_3723,N_2451,N_2386);
nor U3724 (N_3724,N_2265,N_2080);
or U3725 (N_3725,N_2954,N_2542);
or U3726 (N_3726,N_2334,N_2860);
nor U3727 (N_3727,N_2166,N_2255);
or U3728 (N_3728,N_2003,N_2707);
xor U3729 (N_3729,N_2660,N_2922);
nor U3730 (N_3730,N_2905,N_2621);
nor U3731 (N_3731,N_2774,N_2000);
nor U3732 (N_3732,N_2723,N_2786);
nand U3733 (N_3733,N_2391,N_2754);
nand U3734 (N_3734,N_2113,N_2126);
and U3735 (N_3735,N_2868,N_2486);
or U3736 (N_3736,N_2883,N_2329);
nand U3737 (N_3737,N_2643,N_2291);
nor U3738 (N_3738,N_2251,N_2669);
and U3739 (N_3739,N_2022,N_2350);
or U3740 (N_3740,N_2185,N_2069);
nand U3741 (N_3741,N_2162,N_2845);
nand U3742 (N_3742,N_2494,N_2610);
nand U3743 (N_3743,N_2706,N_2471);
and U3744 (N_3744,N_2225,N_2616);
or U3745 (N_3745,N_2117,N_2610);
nand U3746 (N_3746,N_2584,N_2931);
or U3747 (N_3747,N_2192,N_2123);
and U3748 (N_3748,N_2627,N_2763);
nor U3749 (N_3749,N_2231,N_2661);
nor U3750 (N_3750,N_2632,N_2237);
or U3751 (N_3751,N_2456,N_2259);
or U3752 (N_3752,N_2951,N_2518);
nand U3753 (N_3753,N_2652,N_2036);
nor U3754 (N_3754,N_2959,N_2216);
nand U3755 (N_3755,N_2154,N_2758);
nand U3756 (N_3756,N_2180,N_2426);
nor U3757 (N_3757,N_2504,N_2946);
nor U3758 (N_3758,N_2532,N_2306);
nand U3759 (N_3759,N_2612,N_2533);
nor U3760 (N_3760,N_2010,N_2257);
or U3761 (N_3761,N_2853,N_2881);
nor U3762 (N_3762,N_2005,N_2980);
or U3763 (N_3763,N_2123,N_2332);
nor U3764 (N_3764,N_2566,N_2023);
nor U3765 (N_3765,N_2099,N_2369);
and U3766 (N_3766,N_2435,N_2927);
and U3767 (N_3767,N_2712,N_2075);
and U3768 (N_3768,N_2601,N_2250);
or U3769 (N_3769,N_2143,N_2970);
nand U3770 (N_3770,N_2921,N_2772);
nand U3771 (N_3771,N_2396,N_2685);
and U3772 (N_3772,N_2674,N_2411);
nand U3773 (N_3773,N_2921,N_2375);
nor U3774 (N_3774,N_2204,N_2717);
or U3775 (N_3775,N_2653,N_2533);
nor U3776 (N_3776,N_2451,N_2775);
or U3777 (N_3777,N_2080,N_2636);
nand U3778 (N_3778,N_2715,N_2271);
nor U3779 (N_3779,N_2255,N_2340);
or U3780 (N_3780,N_2328,N_2244);
or U3781 (N_3781,N_2004,N_2361);
nor U3782 (N_3782,N_2734,N_2540);
nand U3783 (N_3783,N_2147,N_2051);
and U3784 (N_3784,N_2599,N_2346);
or U3785 (N_3785,N_2341,N_2019);
nand U3786 (N_3786,N_2007,N_2740);
and U3787 (N_3787,N_2711,N_2679);
and U3788 (N_3788,N_2570,N_2580);
nor U3789 (N_3789,N_2347,N_2245);
and U3790 (N_3790,N_2797,N_2680);
nor U3791 (N_3791,N_2095,N_2250);
and U3792 (N_3792,N_2047,N_2728);
or U3793 (N_3793,N_2511,N_2183);
or U3794 (N_3794,N_2428,N_2323);
nor U3795 (N_3795,N_2834,N_2634);
nand U3796 (N_3796,N_2594,N_2935);
nand U3797 (N_3797,N_2163,N_2513);
and U3798 (N_3798,N_2907,N_2516);
or U3799 (N_3799,N_2509,N_2555);
nor U3800 (N_3800,N_2503,N_2341);
or U3801 (N_3801,N_2898,N_2281);
or U3802 (N_3802,N_2486,N_2535);
and U3803 (N_3803,N_2546,N_2113);
or U3804 (N_3804,N_2718,N_2796);
or U3805 (N_3805,N_2234,N_2697);
and U3806 (N_3806,N_2076,N_2372);
or U3807 (N_3807,N_2047,N_2471);
or U3808 (N_3808,N_2108,N_2357);
nand U3809 (N_3809,N_2302,N_2492);
nand U3810 (N_3810,N_2798,N_2680);
or U3811 (N_3811,N_2633,N_2369);
nor U3812 (N_3812,N_2225,N_2124);
and U3813 (N_3813,N_2575,N_2413);
nor U3814 (N_3814,N_2461,N_2717);
and U3815 (N_3815,N_2702,N_2444);
nand U3816 (N_3816,N_2117,N_2746);
or U3817 (N_3817,N_2970,N_2038);
nor U3818 (N_3818,N_2000,N_2175);
or U3819 (N_3819,N_2039,N_2183);
or U3820 (N_3820,N_2712,N_2443);
nand U3821 (N_3821,N_2919,N_2126);
and U3822 (N_3822,N_2603,N_2923);
nor U3823 (N_3823,N_2332,N_2289);
or U3824 (N_3824,N_2749,N_2212);
or U3825 (N_3825,N_2940,N_2122);
nor U3826 (N_3826,N_2379,N_2382);
and U3827 (N_3827,N_2535,N_2617);
nor U3828 (N_3828,N_2958,N_2945);
nor U3829 (N_3829,N_2544,N_2562);
and U3830 (N_3830,N_2872,N_2948);
nor U3831 (N_3831,N_2632,N_2066);
and U3832 (N_3832,N_2781,N_2488);
nor U3833 (N_3833,N_2181,N_2944);
or U3834 (N_3834,N_2212,N_2932);
or U3835 (N_3835,N_2802,N_2360);
and U3836 (N_3836,N_2817,N_2075);
nand U3837 (N_3837,N_2030,N_2782);
nand U3838 (N_3838,N_2301,N_2046);
and U3839 (N_3839,N_2532,N_2664);
nand U3840 (N_3840,N_2073,N_2584);
nor U3841 (N_3841,N_2985,N_2261);
and U3842 (N_3842,N_2119,N_2579);
and U3843 (N_3843,N_2703,N_2032);
or U3844 (N_3844,N_2016,N_2097);
nand U3845 (N_3845,N_2845,N_2044);
or U3846 (N_3846,N_2433,N_2243);
xnor U3847 (N_3847,N_2890,N_2414);
nand U3848 (N_3848,N_2991,N_2734);
and U3849 (N_3849,N_2091,N_2472);
nor U3850 (N_3850,N_2687,N_2773);
nand U3851 (N_3851,N_2413,N_2580);
or U3852 (N_3852,N_2523,N_2121);
nor U3853 (N_3853,N_2489,N_2877);
nor U3854 (N_3854,N_2530,N_2050);
nor U3855 (N_3855,N_2110,N_2392);
and U3856 (N_3856,N_2295,N_2210);
or U3857 (N_3857,N_2481,N_2751);
nand U3858 (N_3858,N_2885,N_2475);
nor U3859 (N_3859,N_2908,N_2279);
nand U3860 (N_3860,N_2726,N_2520);
or U3861 (N_3861,N_2983,N_2136);
or U3862 (N_3862,N_2132,N_2618);
and U3863 (N_3863,N_2713,N_2934);
and U3864 (N_3864,N_2641,N_2819);
nand U3865 (N_3865,N_2389,N_2359);
nand U3866 (N_3866,N_2935,N_2403);
nor U3867 (N_3867,N_2726,N_2870);
and U3868 (N_3868,N_2451,N_2581);
nand U3869 (N_3869,N_2474,N_2056);
or U3870 (N_3870,N_2238,N_2858);
nor U3871 (N_3871,N_2314,N_2565);
and U3872 (N_3872,N_2570,N_2524);
nand U3873 (N_3873,N_2725,N_2504);
and U3874 (N_3874,N_2572,N_2830);
or U3875 (N_3875,N_2737,N_2171);
nor U3876 (N_3876,N_2410,N_2230);
and U3877 (N_3877,N_2351,N_2137);
nand U3878 (N_3878,N_2144,N_2105);
or U3879 (N_3879,N_2153,N_2343);
and U3880 (N_3880,N_2990,N_2087);
nand U3881 (N_3881,N_2210,N_2829);
nand U3882 (N_3882,N_2815,N_2747);
nand U3883 (N_3883,N_2102,N_2021);
nand U3884 (N_3884,N_2431,N_2259);
and U3885 (N_3885,N_2341,N_2559);
or U3886 (N_3886,N_2773,N_2673);
nor U3887 (N_3887,N_2586,N_2013);
and U3888 (N_3888,N_2603,N_2930);
nand U3889 (N_3889,N_2077,N_2694);
nand U3890 (N_3890,N_2257,N_2983);
or U3891 (N_3891,N_2725,N_2961);
nor U3892 (N_3892,N_2772,N_2492);
nand U3893 (N_3893,N_2478,N_2990);
or U3894 (N_3894,N_2313,N_2616);
or U3895 (N_3895,N_2396,N_2363);
or U3896 (N_3896,N_2100,N_2727);
nand U3897 (N_3897,N_2023,N_2458);
or U3898 (N_3898,N_2832,N_2954);
nand U3899 (N_3899,N_2023,N_2947);
nand U3900 (N_3900,N_2563,N_2142);
nor U3901 (N_3901,N_2420,N_2147);
and U3902 (N_3902,N_2590,N_2199);
and U3903 (N_3903,N_2475,N_2751);
or U3904 (N_3904,N_2743,N_2201);
or U3905 (N_3905,N_2685,N_2448);
or U3906 (N_3906,N_2952,N_2963);
nand U3907 (N_3907,N_2010,N_2125);
nand U3908 (N_3908,N_2396,N_2969);
and U3909 (N_3909,N_2104,N_2881);
nand U3910 (N_3910,N_2059,N_2027);
nand U3911 (N_3911,N_2086,N_2896);
nor U3912 (N_3912,N_2373,N_2032);
or U3913 (N_3913,N_2686,N_2225);
and U3914 (N_3914,N_2551,N_2948);
nand U3915 (N_3915,N_2360,N_2078);
or U3916 (N_3916,N_2700,N_2850);
nand U3917 (N_3917,N_2076,N_2825);
or U3918 (N_3918,N_2031,N_2851);
or U3919 (N_3919,N_2718,N_2194);
nor U3920 (N_3920,N_2023,N_2319);
nand U3921 (N_3921,N_2255,N_2927);
nand U3922 (N_3922,N_2212,N_2752);
nand U3923 (N_3923,N_2514,N_2538);
or U3924 (N_3924,N_2604,N_2582);
nor U3925 (N_3925,N_2727,N_2065);
nor U3926 (N_3926,N_2885,N_2448);
or U3927 (N_3927,N_2226,N_2327);
xnor U3928 (N_3928,N_2831,N_2709);
nand U3929 (N_3929,N_2827,N_2850);
and U3930 (N_3930,N_2967,N_2883);
and U3931 (N_3931,N_2956,N_2737);
nand U3932 (N_3932,N_2537,N_2016);
and U3933 (N_3933,N_2397,N_2174);
and U3934 (N_3934,N_2941,N_2603);
nand U3935 (N_3935,N_2005,N_2628);
and U3936 (N_3936,N_2121,N_2455);
nor U3937 (N_3937,N_2941,N_2704);
nor U3938 (N_3938,N_2340,N_2338);
and U3939 (N_3939,N_2022,N_2838);
or U3940 (N_3940,N_2318,N_2256);
or U3941 (N_3941,N_2982,N_2332);
nand U3942 (N_3942,N_2174,N_2250);
and U3943 (N_3943,N_2437,N_2509);
or U3944 (N_3944,N_2252,N_2047);
or U3945 (N_3945,N_2876,N_2018);
nand U3946 (N_3946,N_2609,N_2909);
nand U3947 (N_3947,N_2883,N_2857);
and U3948 (N_3948,N_2834,N_2422);
nor U3949 (N_3949,N_2097,N_2415);
nand U3950 (N_3950,N_2024,N_2287);
nand U3951 (N_3951,N_2862,N_2930);
and U3952 (N_3952,N_2080,N_2060);
or U3953 (N_3953,N_2091,N_2002);
and U3954 (N_3954,N_2263,N_2256);
nor U3955 (N_3955,N_2692,N_2874);
or U3956 (N_3956,N_2314,N_2222);
or U3957 (N_3957,N_2959,N_2969);
or U3958 (N_3958,N_2614,N_2721);
nor U3959 (N_3959,N_2006,N_2091);
or U3960 (N_3960,N_2239,N_2796);
or U3961 (N_3961,N_2260,N_2825);
nand U3962 (N_3962,N_2930,N_2437);
or U3963 (N_3963,N_2148,N_2320);
and U3964 (N_3964,N_2265,N_2646);
or U3965 (N_3965,N_2062,N_2985);
and U3966 (N_3966,N_2995,N_2656);
or U3967 (N_3967,N_2134,N_2644);
nand U3968 (N_3968,N_2816,N_2419);
nand U3969 (N_3969,N_2905,N_2762);
nor U3970 (N_3970,N_2623,N_2936);
nand U3971 (N_3971,N_2762,N_2965);
and U3972 (N_3972,N_2425,N_2334);
or U3973 (N_3973,N_2103,N_2832);
or U3974 (N_3974,N_2057,N_2416);
nor U3975 (N_3975,N_2339,N_2532);
and U3976 (N_3976,N_2643,N_2946);
or U3977 (N_3977,N_2455,N_2913);
nor U3978 (N_3978,N_2082,N_2494);
nor U3979 (N_3979,N_2079,N_2908);
or U3980 (N_3980,N_2264,N_2371);
nor U3981 (N_3981,N_2701,N_2725);
and U3982 (N_3982,N_2046,N_2583);
and U3983 (N_3983,N_2253,N_2306);
and U3984 (N_3984,N_2546,N_2593);
and U3985 (N_3985,N_2272,N_2143);
nor U3986 (N_3986,N_2977,N_2817);
or U3987 (N_3987,N_2654,N_2188);
or U3988 (N_3988,N_2154,N_2462);
nand U3989 (N_3989,N_2540,N_2662);
or U3990 (N_3990,N_2735,N_2412);
and U3991 (N_3991,N_2182,N_2185);
or U3992 (N_3992,N_2494,N_2938);
or U3993 (N_3993,N_2654,N_2935);
and U3994 (N_3994,N_2013,N_2543);
and U3995 (N_3995,N_2007,N_2894);
or U3996 (N_3996,N_2103,N_2122);
nor U3997 (N_3997,N_2507,N_2769);
nand U3998 (N_3998,N_2933,N_2757);
and U3999 (N_3999,N_2278,N_2258);
nor U4000 (N_4000,N_3380,N_3693);
and U4001 (N_4001,N_3867,N_3407);
nand U4002 (N_4002,N_3032,N_3153);
or U4003 (N_4003,N_3151,N_3599);
nand U4004 (N_4004,N_3976,N_3019);
nor U4005 (N_4005,N_3240,N_3885);
and U4006 (N_4006,N_3812,N_3262);
nand U4007 (N_4007,N_3639,N_3426);
or U4008 (N_4008,N_3642,N_3524);
and U4009 (N_4009,N_3231,N_3542);
and U4010 (N_4010,N_3418,N_3598);
nor U4011 (N_4011,N_3543,N_3601);
nand U4012 (N_4012,N_3286,N_3908);
nand U4013 (N_4013,N_3981,N_3261);
nor U4014 (N_4014,N_3587,N_3945);
and U4015 (N_4015,N_3849,N_3409);
nand U4016 (N_4016,N_3149,N_3910);
nor U4017 (N_4017,N_3205,N_3438);
nor U4018 (N_4018,N_3004,N_3566);
and U4019 (N_4019,N_3169,N_3027);
or U4020 (N_4020,N_3898,N_3485);
nor U4021 (N_4021,N_3682,N_3051);
nand U4022 (N_4022,N_3241,N_3395);
and U4023 (N_4023,N_3099,N_3412);
and U4024 (N_4024,N_3069,N_3697);
and U4025 (N_4025,N_3436,N_3500);
or U4026 (N_4026,N_3525,N_3788);
nand U4027 (N_4027,N_3683,N_3091);
or U4028 (N_4028,N_3203,N_3522);
nor U4029 (N_4029,N_3771,N_3660);
and U4030 (N_4030,N_3467,N_3012);
or U4031 (N_4031,N_3825,N_3057);
or U4032 (N_4032,N_3476,N_3782);
nor U4033 (N_4033,N_3650,N_3954);
or U4034 (N_4034,N_3165,N_3884);
and U4035 (N_4035,N_3483,N_3690);
nand U4036 (N_4036,N_3439,N_3901);
nor U4037 (N_4037,N_3523,N_3341);
nor U4038 (N_4038,N_3507,N_3211);
or U4039 (N_4039,N_3181,N_3818);
nor U4040 (N_4040,N_3506,N_3900);
or U4041 (N_4041,N_3848,N_3625);
or U4042 (N_4042,N_3389,N_3223);
nor U4043 (N_4043,N_3368,N_3662);
nor U4044 (N_4044,N_3556,N_3846);
and U4045 (N_4045,N_3580,N_3617);
and U4046 (N_4046,N_3646,N_3873);
or U4047 (N_4047,N_3768,N_3674);
nand U4048 (N_4048,N_3759,N_3354);
nand U4049 (N_4049,N_3992,N_3209);
nand U4050 (N_4050,N_3411,N_3727);
nand U4051 (N_4051,N_3943,N_3877);
nor U4052 (N_4052,N_3445,N_3535);
or U4053 (N_4053,N_3173,N_3538);
nand U4054 (N_4054,N_3725,N_3699);
or U4055 (N_4055,N_3750,N_3925);
or U4056 (N_4056,N_3276,N_3932);
nand U4057 (N_4057,N_3079,N_3317);
nand U4058 (N_4058,N_3893,N_3802);
and U4059 (N_4059,N_3675,N_3633);
and U4060 (N_4060,N_3859,N_3066);
and U4061 (N_4061,N_3422,N_3244);
nor U4062 (N_4062,N_3225,N_3794);
and U4063 (N_4063,N_3095,N_3050);
nor U4064 (N_4064,N_3297,N_3551);
nand U4065 (N_4065,N_3540,N_3872);
nand U4066 (N_4066,N_3714,N_3061);
or U4067 (N_4067,N_3432,N_3147);
or U4068 (N_4068,N_3894,N_3941);
nor U4069 (N_4069,N_3738,N_3928);
nand U4070 (N_4070,N_3776,N_3191);
nor U4071 (N_4071,N_3408,N_3037);
and U4072 (N_4072,N_3356,N_3573);
and U4073 (N_4073,N_3347,N_3806);
nor U4074 (N_4074,N_3866,N_3008);
or U4075 (N_4075,N_3454,N_3936);
nor U4076 (N_4076,N_3074,N_3114);
nand U4077 (N_4077,N_3083,N_3450);
nor U4078 (N_4078,N_3632,N_3670);
nor U4079 (N_4079,N_3529,N_3357);
nand U4080 (N_4080,N_3108,N_3072);
or U4081 (N_4081,N_3391,N_3327);
or U4082 (N_4082,N_3111,N_3162);
nor U4083 (N_4083,N_3552,N_3914);
nand U4084 (N_4084,N_3889,N_3420);
nand U4085 (N_4085,N_3772,N_3948);
or U4086 (N_4086,N_3284,N_3596);
and U4087 (N_4087,N_3110,N_3249);
nor U4088 (N_4088,N_3770,N_3927);
nor U4089 (N_4089,N_3311,N_3344);
nand U4090 (N_4090,N_3164,N_3453);
and U4091 (N_4091,N_3801,N_3196);
nand U4092 (N_4092,N_3030,N_3152);
nand U4093 (N_4093,N_3490,N_3055);
and U4094 (N_4094,N_3629,N_3621);
or U4095 (N_4095,N_3360,N_3237);
and U4096 (N_4096,N_3497,N_3526);
and U4097 (N_4097,N_3938,N_3329);
nor U4098 (N_4098,N_3748,N_3434);
nor U4099 (N_4099,N_3620,N_3955);
nand U4100 (N_4100,N_3602,N_3571);
and U4101 (N_4101,N_3081,N_3805);
and U4102 (N_4102,N_3475,N_3367);
or U4103 (N_4103,N_3887,N_3554);
nor U4104 (N_4104,N_3509,N_3847);
nor U4105 (N_4105,N_3879,N_3774);
and U4106 (N_4106,N_3605,N_3820);
nor U4107 (N_4107,N_3555,N_3519);
nand U4108 (N_4108,N_3756,N_3085);
nor U4109 (N_4109,N_3217,N_3113);
nor U4110 (N_4110,N_3006,N_3664);
or U4111 (N_4111,N_3935,N_3514);
and U4112 (N_4112,N_3864,N_3129);
and U4113 (N_4113,N_3843,N_3220);
and U4114 (N_4114,N_3906,N_3627);
nor U4115 (N_4115,N_3861,N_3919);
or U4116 (N_4116,N_3752,N_3251);
nand U4117 (N_4117,N_3075,N_3126);
or U4118 (N_4118,N_3597,N_3484);
or U4119 (N_4119,N_3589,N_3054);
nor U4120 (N_4120,N_3946,N_3604);
nand U4121 (N_4121,N_3857,N_3248);
and U4122 (N_4122,N_3973,N_3235);
or U4123 (N_4123,N_3266,N_3799);
nor U4124 (N_4124,N_3371,N_3315);
nand U4125 (N_4125,N_3860,N_3005);
nor U4126 (N_4126,N_3060,N_3379);
nand U4127 (N_4127,N_3708,N_3953);
and U4128 (N_4128,N_3146,N_3562);
and U4129 (N_4129,N_3364,N_3661);
nand U4130 (N_4130,N_3647,N_3133);
nand U4131 (N_4131,N_3268,N_3994);
or U4132 (N_4132,N_3545,N_3728);
or U4133 (N_4133,N_3871,N_3583);
or U4134 (N_4134,N_3876,N_3024);
or U4135 (N_4135,N_3840,N_3365);
nand U4136 (N_4136,N_3150,N_3491);
nor U4137 (N_4137,N_3437,N_3218);
and U4138 (N_4138,N_3308,N_3988);
and U4139 (N_4139,N_3299,N_3143);
or U4140 (N_4140,N_3844,N_3245);
or U4141 (N_4141,N_3691,N_3735);
and U4142 (N_4142,N_3335,N_3760);
nand U4143 (N_4143,N_3531,N_3301);
nand U4144 (N_4144,N_3737,N_3657);
nand U4145 (N_4145,N_3983,N_3707);
or U4146 (N_4146,N_3195,N_3731);
or U4147 (N_4147,N_3283,N_3440);
nand U4148 (N_4148,N_3912,N_3212);
nand U4149 (N_4149,N_3716,N_3744);
nor U4150 (N_4150,N_3534,N_3086);
nor U4151 (N_4151,N_3351,N_3918);
nor U4152 (N_4152,N_3082,N_3781);
nor U4153 (N_4153,N_3696,N_3194);
and U4154 (N_4154,N_3607,N_3681);
nor U4155 (N_4155,N_3732,N_3140);
and U4156 (N_4156,N_3511,N_3611);
nand U4157 (N_4157,N_3934,N_3119);
or U4158 (N_4158,N_3558,N_3667);
or U4159 (N_4159,N_3544,N_3274);
nand U4160 (N_4160,N_3285,N_3780);
nor U4161 (N_4161,N_3291,N_3975);
nor U4162 (N_4162,N_3922,N_3659);
nor U4163 (N_4163,N_3466,N_3362);
nor U4164 (N_4164,N_3905,N_3213);
nor U4165 (N_4165,N_3447,N_3115);
and U4166 (N_4166,N_3280,N_3512);
and U4167 (N_4167,N_3797,N_3779);
nand U4168 (N_4168,N_3159,N_3778);
and U4169 (N_4169,N_3459,N_3666);
and U4170 (N_4170,N_3487,N_3845);
nand U4171 (N_4171,N_3987,N_3855);
nand U4172 (N_4172,N_3997,N_3001);
nand U4173 (N_4173,N_3640,N_3678);
and U4174 (N_4174,N_3415,N_3383);
nand U4175 (N_4175,N_3036,N_3586);
nor U4176 (N_4176,N_3498,N_3403);
nand U4177 (N_4177,N_3479,N_3265);
or U4178 (N_4178,N_3536,N_3856);
and U4179 (N_4179,N_3594,N_3321);
nor U4180 (N_4180,N_3862,N_3182);
nand U4181 (N_4181,N_3273,N_3964);
or U4182 (N_4182,N_3713,N_3577);
nor U4183 (N_4183,N_3722,N_3931);
nand U4184 (N_4184,N_3710,N_3148);
nand U4185 (N_4185,N_3185,N_3814);
nand U4186 (N_4186,N_3482,N_3052);
and U4187 (N_4187,N_3917,N_3010);
nand U4188 (N_4188,N_3569,N_3764);
or U4189 (N_4189,N_3798,N_3104);
nor U4190 (N_4190,N_3769,N_3869);
nor U4191 (N_4191,N_3279,N_3324);
nor U4192 (N_4192,N_3358,N_3221);
and U4193 (N_4193,N_3292,N_3790);
and U4194 (N_4194,N_3401,N_3048);
nor U4195 (N_4195,N_3219,N_3773);
nor U4196 (N_4196,N_3747,N_3749);
nand U4197 (N_4197,N_3441,N_3309);
or U4198 (N_4198,N_3921,N_3891);
and U4199 (N_4199,N_3326,N_3736);
nor U4200 (N_4200,N_3503,N_3892);
or U4201 (N_4201,N_3207,N_3090);
nor U4202 (N_4202,N_3168,N_3363);
or U4203 (N_4203,N_3340,N_3916);
nor U4204 (N_4204,N_3288,N_3591);
nand U4205 (N_4205,N_3668,N_3250);
nor U4206 (N_4206,N_3811,N_3680);
and U4207 (N_4207,N_3016,N_3350);
or U4208 (N_4208,N_3800,N_3775);
or U4209 (N_4209,N_3791,N_3305);
or U4210 (N_4210,N_3031,N_3890);
nor U4211 (N_4211,N_3527,N_3157);
nor U4212 (N_4212,N_3565,N_3333);
and U4213 (N_4213,N_3582,N_3508);
nand U4214 (N_4214,N_3575,N_3457);
and U4215 (N_4215,N_3242,N_3015);
nor U4216 (N_4216,N_3971,N_3121);
nor U4217 (N_4217,N_3677,N_3355);
nor U4218 (N_4218,N_3648,N_3658);
nand U4219 (N_4219,N_3841,N_3112);
and U4220 (N_4220,N_3183,N_3366);
or U4221 (N_4221,N_3269,N_3167);
and U4222 (N_4222,N_3762,N_3455);
nor U4223 (N_4223,N_3703,N_3399);
nand U4224 (N_4224,N_3603,N_3043);
nand U4225 (N_4225,N_3089,N_3499);
and U4226 (N_4226,N_3331,N_3247);
and U4227 (N_4227,N_3613,N_3949);
or U4228 (N_4228,N_3616,N_3888);
or U4229 (N_4229,N_3413,N_3233);
nor U4230 (N_4230,N_3076,N_3763);
or U4231 (N_4231,N_3328,N_3128);
or U4232 (N_4232,N_3745,N_3130);
and U4233 (N_4233,N_3372,N_3809);
or U4234 (N_4234,N_3734,N_3641);
and U4235 (N_4235,N_3539,N_3828);
nand U4236 (N_4236,N_3883,N_3042);
or U4237 (N_4237,N_3468,N_3989);
nor U4238 (N_4238,N_3568,N_3614);
and U4239 (N_4239,N_3824,N_3094);
nand U4240 (N_4240,N_3706,N_3807);
nor U4241 (N_4241,N_3702,N_3784);
nor U4242 (N_4242,N_3480,N_3793);
nand U4243 (N_4243,N_3314,N_3656);
and U4244 (N_4244,N_3202,N_3170);
nand U4245 (N_4245,N_3230,N_3720);
or U4246 (N_4246,N_3816,N_3623);
nand U4247 (N_4247,N_3302,N_3904);
and U4248 (N_4248,N_3007,N_3442);
or U4249 (N_4249,N_3258,N_3117);
and U4250 (N_4250,N_3068,N_3836);
nand U4251 (N_4251,N_3990,N_3100);
nor U4252 (N_4252,N_3899,N_3215);
and U4253 (N_4253,N_3572,N_3915);
nand U4254 (N_4254,N_3502,N_3909);
nor U4255 (N_4255,N_3685,N_3272);
nand U4256 (N_4256,N_3561,N_3320);
nor U4257 (N_4257,N_3619,N_3044);
nor U4258 (N_4258,N_3187,N_3406);
and U4259 (N_4259,N_3197,N_3319);
or U4260 (N_4260,N_3939,N_3739);
or U4261 (N_4261,N_3626,N_3281);
nand U4262 (N_4262,N_3505,N_3330);
nor U4263 (N_4263,N_3142,N_3393);
and U4264 (N_4264,N_3684,N_3312);
nand U4265 (N_4265,N_3429,N_3049);
and U4266 (N_4266,N_3131,N_3200);
nand U4267 (N_4267,N_3743,N_3995);
and U4268 (N_4268,N_3070,N_3238);
and U4269 (N_4269,N_3831,N_3137);
nor U4270 (N_4270,N_3622,N_3966);
nand U4271 (N_4271,N_3277,N_3723);
xor U4272 (N_4272,N_3567,N_3926);
and U4273 (N_4273,N_3023,N_3676);
and U4274 (N_4274,N_3645,N_3789);
or U4275 (N_4275,N_3528,N_3134);
nand U4276 (N_4276,N_3106,N_3610);
and U4277 (N_4277,N_3496,N_3854);
and U4278 (N_4278,N_3397,N_3832);
or U4279 (N_4279,N_3753,N_3853);
nand U4280 (N_4280,N_3222,N_3259);
or U4281 (N_4281,N_3155,N_3880);
or U4282 (N_4282,N_3803,N_3998);
nor U4283 (N_4283,N_3882,N_3246);
or U4284 (N_4284,N_3851,N_3991);
nor U4285 (N_4285,N_3040,N_3039);
and U4286 (N_4286,N_3570,N_3107);
and U4287 (N_4287,N_3318,N_3557);
and U4288 (N_4288,N_3996,N_3180);
nand U4289 (N_4289,N_3102,N_3951);
and U4290 (N_4290,N_3630,N_3464);
and U4291 (N_4291,N_3414,N_3494);
nand U4292 (N_4292,N_3135,N_3388);
nor U4293 (N_4293,N_3838,N_3473);
nand U4294 (N_4294,N_3171,N_3352);
and U4295 (N_4295,N_3201,N_3374);
and U4296 (N_4296,N_3576,N_3673);
nor U4297 (N_4297,N_3638,N_3158);
or U4298 (N_4298,N_3672,N_3870);
or U4299 (N_4299,N_3829,N_3385);
nand U4300 (N_4300,N_3698,N_3785);
nand U4301 (N_4301,N_3537,N_3255);
nand U4302 (N_4302,N_3634,N_3033);
nor U4303 (N_4303,N_3977,N_3606);
nand U4304 (N_4304,N_3345,N_3087);
nand U4305 (N_4305,N_3216,N_3993);
or U4306 (N_4306,N_3270,N_3184);
or U4307 (N_4307,N_3028,N_3011);
and U4308 (N_4308,N_3489,N_3177);
nand U4309 (N_4309,N_3254,N_3637);
and U4310 (N_4310,N_3740,N_3236);
nor U4311 (N_4311,N_3593,N_3353);
nor U4312 (N_4312,N_3493,N_3175);
or U4313 (N_4313,N_3751,N_3433);
nand U4314 (N_4314,N_3176,N_3103);
nor U4315 (N_4315,N_3029,N_3478);
and U4316 (N_4316,N_3695,N_3116);
and U4317 (N_4317,N_3755,N_3822);
nor U4318 (N_4318,N_3260,N_3078);
and U4319 (N_4319,N_3190,N_3592);
nand U4320 (N_4320,N_3118,N_3654);
or U4321 (N_4321,N_3448,N_3423);
nand U4322 (N_4322,N_3313,N_3618);
nor U4323 (N_4323,N_3017,N_3850);
or U4324 (N_4324,N_3726,N_3777);
nand U4325 (N_4325,N_3073,N_3549);
or U4326 (N_4326,N_3020,N_3275);
and U4327 (N_4327,N_3421,N_3766);
nand U4328 (N_4328,N_3343,N_3961);
nand U4329 (N_4329,N_3141,N_3224);
or U4330 (N_4330,N_3923,N_3972);
nand U4331 (N_4331,N_3410,N_3821);
nand U4332 (N_4332,N_3227,N_3096);
nand U4333 (N_4333,N_3404,N_3390);
and U4334 (N_4334,N_3669,N_3127);
or U4335 (N_4335,N_3306,N_3842);
and U4336 (N_4336,N_3907,N_3584);
or U4337 (N_4337,N_3346,N_3446);
and U4338 (N_4338,N_3930,N_3635);
and U4339 (N_4339,N_3144,N_3746);
nand U4340 (N_4340,N_3449,N_3548);
or U4341 (N_4341,N_3210,N_3122);
or U4342 (N_4342,N_3174,N_3644);
nor U4343 (N_4343,N_3982,N_3192);
nand U4344 (N_4344,N_3896,N_3088);
and U4345 (N_4345,N_3590,N_3396);
and U4346 (N_4346,N_3694,N_3229);
or U4347 (N_4347,N_3375,N_3711);
nor U4348 (N_4348,N_3047,N_3679);
nor U4349 (N_4349,N_3163,N_3402);
and U4350 (N_4350,N_3232,N_3067);
nor U4351 (N_4351,N_3348,N_3692);
nand U4352 (N_4352,N_3959,N_3462);
nor U4353 (N_4353,N_3826,N_3428);
and U4354 (N_4354,N_3166,N_3098);
nand U4355 (N_4355,N_3701,N_3071);
nand U4356 (N_4356,N_3405,N_3295);
nand U4357 (N_4357,N_3792,N_3724);
and U4358 (N_4358,N_3257,N_3460);
nor U4359 (N_4359,N_3189,N_3895);
nor U4360 (N_4360,N_3835,N_3062);
nand U4361 (N_4361,N_3541,N_3600);
nor U4362 (N_4362,N_3733,N_3980);
or U4363 (N_4363,N_3026,N_3819);
nor U4364 (N_4364,N_3451,N_3712);
nor U4365 (N_4365,N_3704,N_3581);
or U4366 (N_4366,N_3278,N_3056);
and U4367 (N_4367,N_3517,N_3160);
or U4368 (N_4368,N_3786,N_3655);
and U4369 (N_4369,N_3530,N_3628);
nand U4370 (N_4370,N_3435,N_3969);
or U4371 (N_4371,N_3382,N_3559);
nor U4372 (N_4372,N_3014,N_3962);
or U4373 (N_4373,N_3136,N_3105);
and U4374 (N_4374,N_3443,N_3761);
and U4375 (N_4375,N_3120,N_3178);
nor U4376 (N_4376,N_3837,N_3214);
xnor U4377 (N_4377,N_3501,N_3471);
or U4378 (N_4378,N_3765,N_3332);
and U4379 (N_4379,N_3902,N_3767);
nor U4380 (N_4380,N_3974,N_3521);
or U4381 (N_4381,N_3717,N_3394);
or U4382 (N_4382,N_3316,N_3700);
nor U4383 (N_4383,N_3595,N_3349);
nor U4384 (N_4384,N_3193,N_3123);
nand U4385 (N_4385,N_3470,N_3874);
or U4386 (N_4386,N_3243,N_3359);
or U4387 (N_4387,N_3563,N_3481);
nand U4388 (N_4388,N_3553,N_3579);
or U4389 (N_4389,N_3000,N_3924);
nor U4390 (N_4390,N_3064,N_3560);
nand U4391 (N_4391,N_3294,N_3381);
nand U4392 (N_4392,N_3839,N_3077);
and U4393 (N_4393,N_3336,N_3377);
or U4394 (N_4394,N_3392,N_3533);
or U4395 (N_4395,N_3387,N_3665);
nor U4396 (N_4396,N_3817,N_3933);
nor U4397 (N_4397,N_3034,N_3296);
or U4398 (N_4398,N_3132,N_3156);
nor U4399 (N_4399,N_3172,N_3021);
nor U4400 (N_4400,N_3585,N_3041);
or U4401 (N_4401,N_3093,N_3609);
or U4402 (N_4402,N_3234,N_3287);
nand U4403 (N_4403,N_3881,N_3504);
or U4404 (N_4404,N_3431,N_3477);
nand U4405 (N_4405,N_3636,N_3124);
nor U4406 (N_4406,N_3532,N_3513);
nand U4407 (N_4407,N_3025,N_3199);
nor U4408 (N_4408,N_3686,N_3022);
nor U4409 (N_4409,N_3186,N_3038);
nand U4410 (N_4410,N_3084,N_3430);
and U4411 (N_4411,N_3474,N_3937);
nand U4412 (N_4412,N_3425,N_3378);
or U4413 (N_4413,N_3065,N_3687);
nor U4414 (N_4414,N_3967,N_3458);
nor U4415 (N_4415,N_3652,N_3952);
and U4416 (N_4416,N_3546,N_3960);
nor U4417 (N_4417,N_3444,N_3886);
nand U4418 (N_4418,N_3911,N_3092);
or U4419 (N_4419,N_3188,N_3263);
and U4420 (N_4420,N_3827,N_3719);
nor U4421 (N_4421,N_3649,N_3834);
nand U4422 (N_4422,N_3588,N_3520);
nand U4423 (N_4423,N_3957,N_3058);
nand U4424 (N_4424,N_3865,N_3304);
or U4425 (N_4425,N_3461,N_3754);
or U4426 (N_4426,N_3653,N_3705);
or U4427 (N_4427,N_3465,N_3045);
nor U4428 (N_4428,N_3109,N_3958);
xnor U4429 (N_4429,N_3804,N_3495);
or U4430 (N_4430,N_3239,N_3986);
or U4431 (N_4431,N_3944,N_3940);
and U4432 (N_4432,N_3267,N_3709);
nor U4433 (N_4433,N_3833,N_3950);
and U4434 (N_4434,N_3053,N_3264);
or U4435 (N_4435,N_3298,N_3985);
and U4436 (N_4436,N_3271,N_3968);
and U4437 (N_4437,N_3486,N_3424);
nor U4438 (N_4438,N_3035,N_3290);
or U4439 (N_4439,N_3742,N_3920);
or U4440 (N_4440,N_3965,N_3863);
nor U4441 (N_4441,N_3730,N_3325);
nand U4442 (N_4442,N_3868,N_3080);
or U4443 (N_4443,N_3417,N_3813);
nand U4444 (N_4444,N_3386,N_3456);
or U4445 (N_4445,N_3852,N_3013);
nand U4446 (N_4446,N_3956,N_3878);
nand U4447 (N_4447,N_3518,N_3472);
xor U4448 (N_4448,N_3289,N_3337);
nor U4449 (N_4449,N_3721,N_3550);
and U4450 (N_4450,N_3310,N_3663);
and U4451 (N_4451,N_3463,N_3615);
nor U4452 (N_4452,N_3063,N_3624);
nor U4453 (N_4453,N_3947,N_3161);
nor U4454 (N_4454,N_3469,N_3204);
and U4455 (N_4455,N_3758,N_3688);
or U4456 (N_4456,N_3370,N_3307);
or U4457 (N_4457,N_3979,N_3398);
and U4458 (N_4458,N_3003,N_3376);
and U4459 (N_4459,N_3198,N_3715);
nor U4460 (N_4460,N_3154,N_3515);
nand U4461 (N_4461,N_3046,N_3823);
nor U4462 (N_4462,N_3547,N_3815);
nand U4463 (N_4463,N_3903,N_3369);
or U4464 (N_4464,N_3009,N_3631);
nor U4465 (N_4465,N_3783,N_3795);
and U4466 (N_4466,N_3718,N_3139);
or U4467 (N_4467,N_3206,N_3018);
and U4468 (N_4468,N_3875,N_3138);
or U4469 (N_4469,N_3059,N_3897);
or U4470 (N_4470,N_3179,N_3810);
nand U4471 (N_4471,N_3427,N_3929);
or U4472 (N_4472,N_3145,N_3651);
nor U4473 (N_4473,N_3002,N_3578);
or U4474 (N_4474,N_3300,N_3612);
nor U4475 (N_4475,N_3339,N_3256);
and U4476 (N_4476,N_3338,N_3858);
nor U4477 (N_4477,N_3729,N_3978);
nand U4478 (N_4478,N_3322,N_3787);
and U4479 (N_4479,N_3913,N_3323);
nand U4480 (N_4480,N_3671,N_3419);
xnor U4481 (N_4481,N_3416,N_3999);
and U4482 (N_4482,N_3293,N_3334);
nor U4483 (N_4483,N_3564,N_3796);
nand U4484 (N_4484,N_3488,N_3361);
and U4485 (N_4485,N_3516,N_3574);
nand U4486 (N_4486,N_3643,N_3282);
and U4487 (N_4487,N_3510,N_3228);
and U4488 (N_4488,N_3608,N_3373);
nand U4489 (N_4489,N_3252,N_3808);
nand U4490 (N_4490,N_3963,N_3984);
or U4491 (N_4491,N_3830,N_3689);
or U4492 (N_4492,N_3342,N_3125);
nor U4493 (N_4493,N_3400,N_3253);
and U4494 (N_4494,N_3970,N_3097);
or U4495 (N_4495,N_3757,N_3942);
and U4496 (N_4496,N_3741,N_3101);
or U4497 (N_4497,N_3208,N_3303);
nor U4498 (N_4498,N_3492,N_3226);
nand U4499 (N_4499,N_3384,N_3452);
nor U4500 (N_4500,N_3217,N_3413);
and U4501 (N_4501,N_3137,N_3942);
nor U4502 (N_4502,N_3607,N_3384);
or U4503 (N_4503,N_3581,N_3333);
nand U4504 (N_4504,N_3137,N_3876);
nor U4505 (N_4505,N_3429,N_3159);
nor U4506 (N_4506,N_3981,N_3100);
and U4507 (N_4507,N_3416,N_3644);
nor U4508 (N_4508,N_3607,N_3231);
nand U4509 (N_4509,N_3104,N_3954);
nand U4510 (N_4510,N_3563,N_3468);
nand U4511 (N_4511,N_3204,N_3917);
or U4512 (N_4512,N_3561,N_3920);
nor U4513 (N_4513,N_3074,N_3294);
and U4514 (N_4514,N_3621,N_3964);
nor U4515 (N_4515,N_3369,N_3728);
and U4516 (N_4516,N_3162,N_3247);
nand U4517 (N_4517,N_3792,N_3281);
and U4518 (N_4518,N_3472,N_3018);
nand U4519 (N_4519,N_3541,N_3918);
and U4520 (N_4520,N_3565,N_3725);
nand U4521 (N_4521,N_3363,N_3954);
or U4522 (N_4522,N_3841,N_3093);
or U4523 (N_4523,N_3305,N_3796);
nand U4524 (N_4524,N_3263,N_3672);
nor U4525 (N_4525,N_3381,N_3624);
xnor U4526 (N_4526,N_3073,N_3610);
or U4527 (N_4527,N_3045,N_3280);
nand U4528 (N_4528,N_3470,N_3977);
or U4529 (N_4529,N_3860,N_3385);
nor U4530 (N_4530,N_3587,N_3838);
nor U4531 (N_4531,N_3649,N_3282);
and U4532 (N_4532,N_3121,N_3380);
and U4533 (N_4533,N_3809,N_3119);
or U4534 (N_4534,N_3120,N_3594);
xor U4535 (N_4535,N_3791,N_3701);
or U4536 (N_4536,N_3575,N_3600);
or U4537 (N_4537,N_3885,N_3559);
nor U4538 (N_4538,N_3670,N_3039);
nand U4539 (N_4539,N_3226,N_3045);
and U4540 (N_4540,N_3567,N_3859);
nor U4541 (N_4541,N_3654,N_3225);
or U4542 (N_4542,N_3281,N_3224);
and U4543 (N_4543,N_3877,N_3731);
nor U4544 (N_4544,N_3943,N_3974);
nor U4545 (N_4545,N_3431,N_3467);
nor U4546 (N_4546,N_3910,N_3078);
or U4547 (N_4547,N_3967,N_3672);
xnor U4548 (N_4548,N_3721,N_3382);
nor U4549 (N_4549,N_3817,N_3418);
nor U4550 (N_4550,N_3832,N_3157);
and U4551 (N_4551,N_3995,N_3304);
nor U4552 (N_4552,N_3212,N_3544);
nor U4553 (N_4553,N_3781,N_3911);
nand U4554 (N_4554,N_3505,N_3436);
xnor U4555 (N_4555,N_3823,N_3072);
or U4556 (N_4556,N_3119,N_3868);
and U4557 (N_4557,N_3358,N_3309);
nor U4558 (N_4558,N_3695,N_3408);
or U4559 (N_4559,N_3704,N_3666);
and U4560 (N_4560,N_3032,N_3022);
or U4561 (N_4561,N_3060,N_3635);
nor U4562 (N_4562,N_3579,N_3301);
and U4563 (N_4563,N_3368,N_3122);
nor U4564 (N_4564,N_3348,N_3356);
or U4565 (N_4565,N_3278,N_3832);
nand U4566 (N_4566,N_3306,N_3752);
nor U4567 (N_4567,N_3608,N_3840);
nor U4568 (N_4568,N_3957,N_3250);
and U4569 (N_4569,N_3902,N_3846);
nand U4570 (N_4570,N_3287,N_3800);
nand U4571 (N_4571,N_3887,N_3219);
or U4572 (N_4572,N_3198,N_3384);
and U4573 (N_4573,N_3224,N_3237);
or U4574 (N_4574,N_3005,N_3255);
or U4575 (N_4575,N_3243,N_3794);
nand U4576 (N_4576,N_3876,N_3304);
nor U4577 (N_4577,N_3294,N_3379);
or U4578 (N_4578,N_3138,N_3066);
and U4579 (N_4579,N_3375,N_3121);
nor U4580 (N_4580,N_3324,N_3832);
nor U4581 (N_4581,N_3862,N_3464);
nor U4582 (N_4582,N_3474,N_3671);
nor U4583 (N_4583,N_3668,N_3366);
and U4584 (N_4584,N_3646,N_3064);
or U4585 (N_4585,N_3808,N_3419);
nor U4586 (N_4586,N_3988,N_3131);
and U4587 (N_4587,N_3028,N_3424);
and U4588 (N_4588,N_3502,N_3836);
or U4589 (N_4589,N_3510,N_3127);
nand U4590 (N_4590,N_3305,N_3533);
and U4591 (N_4591,N_3735,N_3596);
and U4592 (N_4592,N_3159,N_3166);
or U4593 (N_4593,N_3958,N_3647);
and U4594 (N_4594,N_3586,N_3698);
and U4595 (N_4595,N_3568,N_3130);
nor U4596 (N_4596,N_3850,N_3935);
and U4597 (N_4597,N_3955,N_3025);
nor U4598 (N_4598,N_3634,N_3338);
and U4599 (N_4599,N_3213,N_3904);
and U4600 (N_4600,N_3490,N_3081);
nand U4601 (N_4601,N_3992,N_3267);
or U4602 (N_4602,N_3749,N_3822);
nand U4603 (N_4603,N_3459,N_3615);
or U4604 (N_4604,N_3063,N_3199);
or U4605 (N_4605,N_3485,N_3665);
nand U4606 (N_4606,N_3575,N_3083);
nand U4607 (N_4607,N_3936,N_3914);
nor U4608 (N_4608,N_3224,N_3998);
and U4609 (N_4609,N_3654,N_3487);
and U4610 (N_4610,N_3790,N_3078);
nand U4611 (N_4611,N_3350,N_3326);
nand U4612 (N_4612,N_3462,N_3883);
or U4613 (N_4613,N_3258,N_3114);
nor U4614 (N_4614,N_3767,N_3029);
nor U4615 (N_4615,N_3855,N_3934);
nor U4616 (N_4616,N_3838,N_3238);
nor U4617 (N_4617,N_3877,N_3333);
and U4618 (N_4618,N_3226,N_3799);
and U4619 (N_4619,N_3790,N_3730);
nor U4620 (N_4620,N_3364,N_3108);
and U4621 (N_4621,N_3089,N_3281);
nor U4622 (N_4622,N_3025,N_3932);
or U4623 (N_4623,N_3131,N_3213);
and U4624 (N_4624,N_3976,N_3950);
and U4625 (N_4625,N_3406,N_3450);
or U4626 (N_4626,N_3882,N_3777);
nor U4627 (N_4627,N_3970,N_3317);
or U4628 (N_4628,N_3826,N_3856);
or U4629 (N_4629,N_3897,N_3055);
nor U4630 (N_4630,N_3865,N_3461);
or U4631 (N_4631,N_3270,N_3001);
and U4632 (N_4632,N_3946,N_3516);
or U4633 (N_4633,N_3430,N_3593);
and U4634 (N_4634,N_3514,N_3564);
or U4635 (N_4635,N_3201,N_3604);
nor U4636 (N_4636,N_3245,N_3950);
and U4637 (N_4637,N_3160,N_3493);
nand U4638 (N_4638,N_3280,N_3627);
and U4639 (N_4639,N_3434,N_3375);
or U4640 (N_4640,N_3857,N_3719);
nand U4641 (N_4641,N_3329,N_3745);
nand U4642 (N_4642,N_3883,N_3396);
nor U4643 (N_4643,N_3803,N_3290);
and U4644 (N_4644,N_3645,N_3267);
nor U4645 (N_4645,N_3800,N_3749);
nor U4646 (N_4646,N_3612,N_3873);
nand U4647 (N_4647,N_3026,N_3010);
nand U4648 (N_4648,N_3983,N_3561);
nor U4649 (N_4649,N_3338,N_3988);
nand U4650 (N_4650,N_3859,N_3468);
and U4651 (N_4651,N_3945,N_3621);
nand U4652 (N_4652,N_3819,N_3408);
or U4653 (N_4653,N_3638,N_3367);
nand U4654 (N_4654,N_3504,N_3516);
nor U4655 (N_4655,N_3554,N_3853);
nor U4656 (N_4656,N_3129,N_3915);
and U4657 (N_4657,N_3634,N_3104);
nand U4658 (N_4658,N_3634,N_3623);
nand U4659 (N_4659,N_3694,N_3959);
and U4660 (N_4660,N_3525,N_3471);
nand U4661 (N_4661,N_3226,N_3270);
and U4662 (N_4662,N_3521,N_3132);
and U4663 (N_4663,N_3099,N_3396);
nor U4664 (N_4664,N_3233,N_3827);
nand U4665 (N_4665,N_3178,N_3828);
and U4666 (N_4666,N_3678,N_3560);
or U4667 (N_4667,N_3459,N_3177);
or U4668 (N_4668,N_3161,N_3527);
or U4669 (N_4669,N_3370,N_3269);
or U4670 (N_4670,N_3189,N_3399);
nand U4671 (N_4671,N_3821,N_3691);
nor U4672 (N_4672,N_3133,N_3097);
and U4673 (N_4673,N_3915,N_3753);
or U4674 (N_4674,N_3430,N_3873);
or U4675 (N_4675,N_3389,N_3127);
nor U4676 (N_4676,N_3064,N_3011);
nor U4677 (N_4677,N_3492,N_3854);
and U4678 (N_4678,N_3089,N_3785);
xnor U4679 (N_4679,N_3210,N_3077);
nand U4680 (N_4680,N_3860,N_3851);
xor U4681 (N_4681,N_3143,N_3164);
nor U4682 (N_4682,N_3271,N_3714);
or U4683 (N_4683,N_3900,N_3203);
nand U4684 (N_4684,N_3352,N_3844);
nand U4685 (N_4685,N_3748,N_3443);
and U4686 (N_4686,N_3084,N_3270);
or U4687 (N_4687,N_3271,N_3690);
and U4688 (N_4688,N_3002,N_3600);
nand U4689 (N_4689,N_3783,N_3534);
or U4690 (N_4690,N_3169,N_3327);
nor U4691 (N_4691,N_3178,N_3219);
and U4692 (N_4692,N_3642,N_3077);
nor U4693 (N_4693,N_3793,N_3696);
or U4694 (N_4694,N_3714,N_3434);
or U4695 (N_4695,N_3737,N_3067);
nor U4696 (N_4696,N_3259,N_3621);
nand U4697 (N_4697,N_3732,N_3755);
xor U4698 (N_4698,N_3779,N_3499);
nand U4699 (N_4699,N_3639,N_3381);
and U4700 (N_4700,N_3045,N_3703);
and U4701 (N_4701,N_3517,N_3043);
nor U4702 (N_4702,N_3312,N_3113);
or U4703 (N_4703,N_3671,N_3995);
nand U4704 (N_4704,N_3142,N_3512);
nor U4705 (N_4705,N_3883,N_3933);
nor U4706 (N_4706,N_3239,N_3546);
and U4707 (N_4707,N_3612,N_3265);
or U4708 (N_4708,N_3366,N_3058);
or U4709 (N_4709,N_3298,N_3902);
or U4710 (N_4710,N_3346,N_3067);
and U4711 (N_4711,N_3311,N_3581);
and U4712 (N_4712,N_3364,N_3739);
nor U4713 (N_4713,N_3497,N_3977);
and U4714 (N_4714,N_3565,N_3509);
or U4715 (N_4715,N_3101,N_3235);
and U4716 (N_4716,N_3535,N_3385);
nand U4717 (N_4717,N_3388,N_3226);
or U4718 (N_4718,N_3507,N_3748);
nand U4719 (N_4719,N_3820,N_3838);
or U4720 (N_4720,N_3137,N_3221);
and U4721 (N_4721,N_3590,N_3247);
and U4722 (N_4722,N_3102,N_3000);
or U4723 (N_4723,N_3196,N_3058);
nand U4724 (N_4724,N_3203,N_3931);
nor U4725 (N_4725,N_3657,N_3422);
nor U4726 (N_4726,N_3984,N_3894);
and U4727 (N_4727,N_3045,N_3756);
and U4728 (N_4728,N_3567,N_3708);
nor U4729 (N_4729,N_3142,N_3147);
nand U4730 (N_4730,N_3832,N_3108);
nand U4731 (N_4731,N_3085,N_3290);
nor U4732 (N_4732,N_3609,N_3506);
and U4733 (N_4733,N_3426,N_3677);
nand U4734 (N_4734,N_3010,N_3533);
nor U4735 (N_4735,N_3334,N_3887);
or U4736 (N_4736,N_3513,N_3279);
nor U4737 (N_4737,N_3973,N_3240);
nand U4738 (N_4738,N_3769,N_3411);
nor U4739 (N_4739,N_3090,N_3732);
nand U4740 (N_4740,N_3861,N_3088);
and U4741 (N_4741,N_3885,N_3045);
nor U4742 (N_4742,N_3278,N_3261);
or U4743 (N_4743,N_3173,N_3531);
nor U4744 (N_4744,N_3484,N_3319);
nand U4745 (N_4745,N_3157,N_3433);
nand U4746 (N_4746,N_3573,N_3948);
nor U4747 (N_4747,N_3469,N_3767);
or U4748 (N_4748,N_3226,N_3499);
nand U4749 (N_4749,N_3595,N_3299);
and U4750 (N_4750,N_3479,N_3563);
nand U4751 (N_4751,N_3224,N_3483);
nor U4752 (N_4752,N_3664,N_3039);
or U4753 (N_4753,N_3875,N_3858);
nor U4754 (N_4754,N_3525,N_3869);
and U4755 (N_4755,N_3015,N_3255);
or U4756 (N_4756,N_3106,N_3689);
or U4757 (N_4757,N_3509,N_3908);
nand U4758 (N_4758,N_3750,N_3899);
and U4759 (N_4759,N_3678,N_3445);
or U4760 (N_4760,N_3717,N_3385);
and U4761 (N_4761,N_3198,N_3114);
nor U4762 (N_4762,N_3766,N_3824);
nand U4763 (N_4763,N_3111,N_3103);
nand U4764 (N_4764,N_3403,N_3110);
or U4765 (N_4765,N_3551,N_3372);
nor U4766 (N_4766,N_3989,N_3092);
nor U4767 (N_4767,N_3314,N_3034);
nor U4768 (N_4768,N_3227,N_3250);
or U4769 (N_4769,N_3610,N_3326);
or U4770 (N_4770,N_3371,N_3545);
and U4771 (N_4771,N_3446,N_3123);
and U4772 (N_4772,N_3097,N_3945);
nor U4773 (N_4773,N_3110,N_3756);
nor U4774 (N_4774,N_3286,N_3182);
nand U4775 (N_4775,N_3395,N_3336);
and U4776 (N_4776,N_3089,N_3710);
nand U4777 (N_4777,N_3688,N_3286);
nor U4778 (N_4778,N_3595,N_3622);
nor U4779 (N_4779,N_3409,N_3082);
nor U4780 (N_4780,N_3114,N_3619);
or U4781 (N_4781,N_3372,N_3487);
nand U4782 (N_4782,N_3939,N_3912);
nor U4783 (N_4783,N_3496,N_3616);
or U4784 (N_4784,N_3732,N_3619);
or U4785 (N_4785,N_3242,N_3171);
or U4786 (N_4786,N_3771,N_3380);
or U4787 (N_4787,N_3420,N_3599);
and U4788 (N_4788,N_3757,N_3484);
or U4789 (N_4789,N_3093,N_3715);
nand U4790 (N_4790,N_3106,N_3884);
or U4791 (N_4791,N_3090,N_3573);
nand U4792 (N_4792,N_3624,N_3329);
nand U4793 (N_4793,N_3498,N_3282);
nor U4794 (N_4794,N_3003,N_3735);
nor U4795 (N_4795,N_3914,N_3808);
nor U4796 (N_4796,N_3887,N_3489);
and U4797 (N_4797,N_3705,N_3695);
and U4798 (N_4798,N_3298,N_3944);
and U4799 (N_4799,N_3306,N_3271);
and U4800 (N_4800,N_3506,N_3777);
or U4801 (N_4801,N_3892,N_3010);
or U4802 (N_4802,N_3235,N_3038);
nand U4803 (N_4803,N_3951,N_3006);
and U4804 (N_4804,N_3713,N_3240);
and U4805 (N_4805,N_3714,N_3737);
and U4806 (N_4806,N_3743,N_3913);
or U4807 (N_4807,N_3797,N_3442);
and U4808 (N_4808,N_3498,N_3906);
or U4809 (N_4809,N_3120,N_3280);
nor U4810 (N_4810,N_3181,N_3731);
or U4811 (N_4811,N_3545,N_3395);
or U4812 (N_4812,N_3281,N_3801);
or U4813 (N_4813,N_3727,N_3739);
nor U4814 (N_4814,N_3198,N_3891);
and U4815 (N_4815,N_3343,N_3206);
nor U4816 (N_4816,N_3114,N_3369);
and U4817 (N_4817,N_3256,N_3972);
or U4818 (N_4818,N_3951,N_3746);
nor U4819 (N_4819,N_3756,N_3809);
nor U4820 (N_4820,N_3001,N_3595);
nor U4821 (N_4821,N_3323,N_3370);
nand U4822 (N_4822,N_3065,N_3449);
or U4823 (N_4823,N_3651,N_3244);
or U4824 (N_4824,N_3462,N_3383);
and U4825 (N_4825,N_3740,N_3561);
or U4826 (N_4826,N_3722,N_3770);
nor U4827 (N_4827,N_3693,N_3318);
nor U4828 (N_4828,N_3838,N_3781);
and U4829 (N_4829,N_3341,N_3852);
xnor U4830 (N_4830,N_3906,N_3678);
nand U4831 (N_4831,N_3655,N_3935);
nor U4832 (N_4832,N_3828,N_3418);
and U4833 (N_4833,N_3566,N_3890);
nand U4834 (N_4834,N_3905,N_3886);
or U4835 (N_4835,N_3331,N_3014);
nand U4836 (N_4836,N_3074,N_3609);
and U4837 (N_4837,N_3778,N_3481);
nor U4838 (N_4838,N_3636,N_3325);
and U4839 (N_4839,N_3828,N_3219);
nor U4840 (N_4840,N_3647,N_3020);
or U4841 (N_4841,N_3456,N_3854);
or U4842 (N_4842,N_3956,N_3129);
nor U4843 (N_4843,N_3820,N_3375);
or U4844 (N_4844,N_3417,N_3633);
nand U4845 (N_4845,N_3729,N_3236);
nand U4846 (N_4846,N_3123,N_3000);
nand U4847 (N_4847,N_3592,N_3252);
and U4848 (N_4848,N_3482,N_3223);
or U4849 (N_4849,N_3988,N_3801);
and U4850 (N_4850,N_3380,N_3622);
nand U4851 (N_4851,N_3338,N_3351);
and U4852 (N_4852,N_3684,N_3615);
or U4853 (N_4853,N_3143,N_3537);
nor U4854 (N_4854,N_3254,N_3062);
and U4855 (N_4855,N_3574,N_3822);
nor U4856 (N_4856,N_3455,N_3369);
or U4857 (N_4857,N_3794,N_3889);
and U4858 (N_4858,N_3949,N_3200);
and U4859 (N_4859,N_3636,N_3861);
and U4860 (N_4860,N_3271,N_3219);
nor U4861 (N_4861,N_3636,N_3878);
nand U4862 (N_4862,N_3472,N_3990);
nand U4863 (N_4863,N_3644,N_3898);
nand U4864 (N_4864,N_3896,N_3453);
nand U4865 (N_4865,N_3699,N_3212);
nor U4866 (N_4866,N_3447,N_3164);
or U4867 (N_4867,N_3744,N_3827);
nand U4868 (N_4868,N_3286,N_3488);
nand U4869 (N_4869,N_3183,N_3564);
nand U4870 (N_4870,N_3743,N_3574);
nand U4871 (N_4871,N_3928,N_3225);
and U4872 (N_4872,N_3794,N_3630);
and U4873 (N_4873,N_3463,N_3395);
nor U4874 (N_4874,N_3346,N_3641);
nor U4875 (N_4875,N_3065,N_3441);
and U4876 (N_4876,N_3158,N_3846);
nor U4877 (N_4877,N_3770,N_3039);
nor U4878 (N_4878,N_3378,N_3836);
nor U4879 (N_4879,N_3657,N_3477);
or U4880 (N_4880,N_3649,N_3541);
and U4881 (N_4881,N_3944,N_3681);
nor U4882 (N_4882,N_3145,N_3334);
or U4883 (N_4883,N_3185,N_3321);
and U4884 (N_4884,N_3704,N_3183);
or U4885 (N_4885,N_3009,N_3130);
and U4886 (N_4886,N_3867,N_3282);
and U4887 (N_4887,N_3611,N_3642);
and U4888 (N_4888,N_3745,N_3104);
nand U4889 (N_4889,N_3214,N_3012);
and U4890 (N_4890,N_3662,N_3421);
and U4891 (N_4891,N_3301,N_3733);
nand U4892 (N_4892,N_3573,N_3900);
or U4893 (N_4893,N_3644,N_3804);
or U4894 (N_4894,N_3191,N_3889);
nor U4895 (N_4895,N_3439,N_3713);
nand U4896 (N_4896,N_3638,N_3666);
nand U4897 (N_4897,N_3627,N_3699);
and U4898 (N_4898,N_3742,N_3428);
nor U4899 (N_4899,N_3226,N_3087);
or U4900 (N_4900,N_3927,N_3260);
or U4901 (N_4901,N_3546,N_3454);
or U4902 (N_4902,N_3035,N_3022);
nor U4903 (N_4903,N_3120,N_3276);
nor U4904 (N_4904,N_3816,N_3375);
nor U4905 (N_4905,N_3949,N_3371);
nand U4906 (N_4906,N_3349,N_3815);
nand U4907 (N_4907,N_3381,N_3912);
or U4908 (N_4908,N_3066,N_3610);
or U4909 (N_4909,N_3168,N_3275);
nor U4910 (N_4910,N_3820,N_3924);
and U4911 (N_4911,N_3253,N_3238);
nor U4912 (N_4912,N_3272,N_3695);
and U4913 (N_4913,N_3950,N_3944);
or U4914 (N_4914,N_3077,N_3097);
nand U4915 (N_4915,N_3487,N_3364);
or U4916 (N_4916,N_3580,N_3019);
nor U4917 (N_4917,N_3266,N_3213);
nor U4918 (N_4918,N_3612,N_3337);
nor U4919 (N_4919,N_3026,N_3322);
nor U4920 (N_4920,N_3041,N_3307);
nor U4921 (N_4921,N_3673,N_3216);
nand U4922 (N_4922,N_3752,N_3601);
or U4923 (N_4923,N_3343,N_3339);
or U4924 (N_4924,N_3306,N_3796);
or U4925 (N_4925,N_3680,N_3515);
or U4926 (N_4926,N_3758,N_3809);
and U4927 (N_4927,N_3494,N_3255);
nand U4928 (N_4928,N_3139,N_3622);
or U4929 (N_4929,N_3211,N_3221);
and U4930 (N_4930,N_3173,N_3421);
and U4931 (N_4931,N_3585,N_3145);
nor U4932 (N_4932,N_3534,N_3686);
nand U4933 (N_4933,N_3318,N_3087);
nand U4934 (N_4934,N_3800,N_3106);
or U4935 (N_4935,N_3066,N_3321);
nand U4936 (N_4936,N_3267,N_3638);
nand U4937 (N_4937,N_3812,N_3486);
xnor U4938 (N_4938,N_3219,N_3943);
and U4939 (N_4939,N_3977,N_3375);
nand U4940 (N_4940,N_3657,N_3117);
and U4941 (N_4941,N_3678,N_3838);
nor U4942 (N_4942,N_3714,N_3371);
nand U4943 (N_4943,N_3766,N_3307);
and U4944 (N_4944,N_3364,N_3983);
nand U4945 (N_4945,N_3227,N_3577);
nor U4946 (N_4946,N_3874,N_3038);
or U4947 (N_4947,N_3349,N_3819);
nor U4948 (N_4948,N_3343,N_3720);
or U4949 (N_4949,N_3466,N_3901);
or U4950 (N_4950,N_3046,N_3167);
and U4951 (N_4951,N_3593,N_3988);
or U4952 (N_4952,N_3923,N_3932);
nand U4953 (N_4953,N_3301,N_3732);
nand U4954 (N_4954,N_3697,N_3957);
or U4955 (N_4955,N_3903,N_3636);
and U4956 (N_4956,N_3068,N_3717);
and U4957 (N_4957,N_3336,N_3986);
nor U4958 (N_4958,N_3718,N_3560);
nand U4959 (N_4959,N_3971,N_3003);
nand U4960 (N_4960,N_3313,N_3783);
nand U4961 (N_4961,N_3754,N_3889);
nand U4962 (N_4962,N_3892,N_3819);
nand U4963 (N_4963,N_3621,N_3085);
nor U4964 (N_4964,N_3980,N_3454);
and U4965 (N_4965,N_3240,N_3083);
and U4966 (N_4966,N_3088,N_3218);
nor U4967 (N_4967,N_3749,N_3717);
and U4968 (N_4968,N_3486,N_3414);
and U4969 (N_4969,N_3015,N_3557);
nor U4970 (N_4970,N_3625,N_3649);
and U4971 (N_4971,N_3774,N_3557);
nand U4972 (N_4972,N_3873,N_3459);
nand U4973 (N_4973,N_3468,N_3630);
or U4974 (N_4974,N_3233,N_3042);
xnor U4975 (N_4975,N_3403,N_3585);
or U4976 (N_4976,N_3150,N_3008);
nor U4977 (N_4977,N_3645,N_3793);
and U4978 (N_4978,N_3696,N_3173);
and U4979 (N_4979,N_3985,N_3115);
or U4980 (N_4980,N_3636,N_3365);
nor U4981 (N_4981,N_3069,N_3951);
or U4982 (N_4982,N_3979,N_3621);
or U4983 (N_4983,N_3050,N_3792);
or U4984 (N_4984,N_3111,N_3186);
nand U4985 (N_4985,N_3529,N_3878);
nor U4986 (N_4986,N_3930,N_3006);
or U4987 (N_4987,N_3568,N_3942);
or U4988 (N_4988,N_3742,N_3599);
nor U4989 (N_4989,N_3946,N_3717);
nand U4990 (N_4990,N_3451,N_3819);
nand U4991 (N_4991,N_3627,N_3065);
or U4992 (N_4992,N_3816,N_3660);
and U4993 (N_4993,N_3755,N_3780);
nor U4994 (N_4994,N_3600,N_3261);
and U4995 (N_4995,N_3928,N_3683);
and U4996 (N_4996,N_3681,N_3828);
and U4997 (N_4997,N_3289,N_3799);
xor U4998 (N_4998,N_3533,N_3014);
nor U4999 (N_4999,N_3536,N_3660);
and UO_0 (O_0,N_4671,N_4713);
nor UO_1 (O_1,N_4210,N_4398);
nand UO_2 (O_2,N_4315,N_4628);
and UO_3 (O_3,N_4590,N_4108);
nor UO_4 (O_4,N_4490,N_4668);
nand UO_5 (O_5,N_4772,N_4260);
or UO_6 (O_6,N_4185,N_4664);
nand UO_7 (O_7,N_4451,N_4228);
or UO_8 (O_8,N_4280,N_4016);
nand UO_9 (O_9,N_4548,N_4096);
nor UO_10 (O_10,N_4598,N_4339);
xor UO_11 (O_11,N_4028,N_4361);
nand UO_12 (O_12,N_4699,N_4764);
nor UO_13 (O_13,N_4638,N_4927);
nor UO_14 (O_14,N_4393,N_4025);
nand UO_15 (O_15,N_4038,N_4765);
and UO_16 (O_16,N_4435,N_4661);
nand UO_17 (O_17,N_4005,N_4122);
nor UO_18 (O_18,N_4828,N_4763);
and UO_19 (O_19,N_4790,N_4984);
nor UO_20 (O_20,N_4876,N_4758);
or UO_21 (O_21,N_4870,N_4021);
nand UO_22 (O_22,N_4233,N_4417);
or UO_23 (O_23,N_4505,N_4866);
or UO_24 (O_24,N_4564,N_4766);
or UO_25 (O_25,N_4012,N_4113);
nand UO_26 (O_26,N_4329,N_4886);
nor UO_27 (O_27,N_4254,N_4566);
nand UO_28 (O_28,N_4854,N_4223);
nand UO_29 (O_29,N_4261,N_4582);
and UO_30 (O_30,N_4434,N_4229);
and UO_31 (O_31,N_4525,N_4808);
nor UO_32 (O_32,N_4104,N_4546);
or UO_33 (O_33,N_4344,N_4952);
and UO_34 (O_34,N_4889,N_4513);
nand UO_35 (O_35,N_4879,N_4636);
nand UO_36 (O_36,N_4819,N_4450);
or UO_37 (O_37,N_4703,N_4720);
nor UO_38 (O_38,N_4396,N_4920);
and UO_39 (O_39,N_4487,N_4863);
nand UO_40 (O_40,N_4418,N_4079);
nor UO_41 (O_41,N_4964,N_4144);
nor UO_42 (O_42,N_4107,N_4355);
or UO_43 (O_43,N_4284,N_4171);
or UO_44 (O_44,N_4717,N_4731);
nor UO_45 (O_45,N_4883,N_4724);
or UO_46 (O_46,N_4794,N_4508);
and UO_47 (O_47,N_4730,N_4756);
or UO_48 (O_48,N_4087,N_4799);
or UO_49 (O_49,N_4949,N_4608);
or UO_50 (O_50,N_4742,N_4409);
and UO_51 (O_51,N_4406,N_4175);
nor UO_52 (O_52,N_4888,N_4620);
and UO_53 (O_53,N_4629,N_4138);
nor UO_54 (O_54,N_4824,N_4156);
or UO_55 (O_55,N_4204,N_4959);
and UO_56 (O_56,N_4771,N_4786);
nand UO_57 (O_57,N_4504,N_4330);
nand UO_58 (O_58,N_4321,N_4390);
or UO_59 (O_59,N_4492,N_4547);
nand UO_60 (O_60,N_4923,N_4484);
nand UO_61 (O_61,N_4675,N_4813);
nand UO_62 (O_62,N_4779,N_4128);
nor UO_63 (O_63,N_4181,N_4563);
nand UO_64 (O_64,N_4930,N_4810);
nand UO_65 (O_65,N_4008,N_4585);
or UO_66 (O_66,N_4403,N_4896);
or UO_67 (O_67,N_4444,N_4732);
nor UO_68 (O_68,N_4076,N_4094);
and UO_69 (O_69,N_4066,N_4309);
nor UO_70 (O_70,N_4678,N_4437);
nand UO_71 (O_71,N_4855,N_4277);
or UO_72 (O_72,N_4022,N_4542);
and UO_73 (O_73,N_4902,N_4752);
and UO_74 (O_74,N_4065,N_4232);
nor UO_75 (O_75,N_4788,N_4818);
or UO_76 (O_76,N_4308,N_4827);
nor UO_77 (O_77,N_4226,N_4728);
nand UO_78 (O_78,N_4457,N_4432);
or UO_79 (O_79,N_4691,N_4734);
nor UO_80 (O_80,N_4419,N_4208);
nor UO_81 (O_81,N_4874,N_4967);
or UO_82 (O_82,N_4955,N_4755);
nor UO_83 (O_83,N_4074,N_4740);
or UO_84 (O_84,N_4999,N_4778);
nor UO_85 (O_85,N_4710,N_4535);
or UO_86 (O_86,N_4679,N_4759);
nand UO_87 (O_87,N_4520,N_4797);
nand UO_88 (O_88,N_4300,N_4946);
nand UO_89 (O_89,N_4338,N_4500);
and UO_90 (O_90,N_4268,N_4561);
nor UO_91 (O_91,N_4369,N_4873);
nand UO_92 (O_92,N_4847,N_4735);
or UO_93 (O_93,N_4626,N_4424);
or UO_94 (O_94,N_4426,N_4231);
and UO_95 (O_95,N_4793,N_4466);
nor UO_96 (O_96,N_4602,N_4979);
nand UO_97 (O_97,N_4910,N_4506);
nor UO_98 (O_98,N_4605,N_4032);
nand UO_99 (O_99,N_4106,N_4958);
nor UO_100 (O_100,N_4861,N_4634);
nor UO_101 (O_101,N_4407,N_4395);
xor UO_102 (O_102,N_4990,N_4892);
and UO_103 (O_103,N_4242,N_4502);
or UO_104 (O_104,N_4324,N_4286);
and UO_105 (O_105,N_4681,N_4622);
and UO_106 (O_106,N_4116,N_4310);
nand UO_107 (O_107,N_4187,N_4147);
nand UO_108 (O_108,N_4544,N_4439);
and UO_109 (O_109,N_4953,N_4741);
and UO_110 (O_110,N_4427,N_4648);
and UO_111 (O_111,N_4951,N_4976);
nor UO_112 (O_112,N_4317,N_4553);
nand UO_113 (O_113,N_4376,N_4467);
or UO_114 (O_114,N_4639,N_4482);
and UO_115 (O_115,N_4982,N_4379);
or UO_116 (O_116,N_4653,N_4770);
nand UO_117 (O_117,N_4158,N_4575);
or UO_118 (O_118,N_4545,N_4862);
nand UO_119 (O_119,N_4283,N_4265);
nand UO_120 (O_120,N_4531,N_4061);
and UO_121 (O_121,N_4216,N_4729);
nor UO_122 (O_122,N_4701,N_4841);
nand UO_123 (O_123,N_4491,N_4867);
nor UO_124 (O_124,N_4860,N_4781);
nor UO_125 (O_125,N_4987,N_4462);
nor UO_126 (O_126,N_4363,N_4213);
nand UO_127 (O_127,N_4239,N_4619);
nand UO_128 (O_128,N_4688,N_4472);
nor UO_129 (O_129,N_4095,N_4201);
and UO_130 (O_130,N_4932,N_4745);
nand UO_131 (O_131,N_4612,N_4938);
or UO_132 (O_132,N_4716,N_4336);
nor UO_133 (O_133,N_4000,N_4599);
nor UO_134 (O_134,N_4359,N_4807);
nor UO_135 (O_135,N_4684,N_4013);
or UO_136 (O_136,N_4798,N_4081);
nor UO_137 (O_137,N_4244,N_4843);
nand UO_138 (O_138,N_4045,N_4044);
nor UO_139 (O_139,N_4782,N_4658);
and UO_140 (O_140,N_4882,N_4551);
nor UO_141 (O_141,N_4459,N_4985);
nand UO_142 (O_142,N_4014,N_4596);
or UO_143 (O_143,N_4846,N_4934);
or UO_144 (O_144,N_4271,N_4868);
nor UO_145 (O_145,N_4978,N_4054);
and UO_146 (O_146,N_4230,N_4404);
nor UO_147 (O_147,N_4831,N_4067);
nor UO_148 (O_148,N_4263,N_4129);
or UO_149 (O_149,N_4683,N_4238);
nand UO_150 (O_150,N_4218,N_4307);
nor UO_151 (O_151,N_4665,N_4972);
xor UO_152 (O_152,N_4402,N_4919);
or UO_153 (O_153,N_4362,N_4420);
nand UO_154 (O_154,N_4891,N_4448);
nand UO_155 (O_155,N_4093,N_4311);
and UO_156 (O_156,N_4202,N_4225);
nor UO_157 (O_157,N_4182,N_4850);
or UO_158 (O_158,N_4885,N_4611);
or UO_159 (O_159,N_4627,N_4374);
nand UO_160 (O_160,N_4991,N_4249);
or UO_161 (O_161,N_4814,N_4774);
and UO_162 (O_162,N_4533,N_4989);
and UO_163 (O_163,N_4913,N_4852);
nand UO_164 (O_164,N_4077,N_4099);
nor UO_165 (O_165,N_4526,N_4801);
or UO_166 (O_166,N_4473,N_4948);
and UO_167 (O_167,N_4083,N_4800);
nand UO_168 (O_168,N_4997,N_4162);
and UO_169 (O_169,N_4121,N_4534);
nor UO_170 (O_170,N_4767,N_4647);
nand UO_171 (O_171,N_4371,N_4373);
nand UO_172 (O_172,N_4392,N_4893);
nor UO_173 (O_173,N_4170,N_4365);
nor UO_174 (O_174,N_4707,N_4836);
or UO_175 (O_175,N_4475,N_4273);
nand UO_176 (O_176,N_4141,N_4354);
nor UO_177 (O_177,N_4711,N_4441);
nand UO_178 (O_178,N_4837,N_4519);
nand UO_179 (O_179,N_4963,N_4222);
or UO_180 (O_180,N_4349,N_4199);
nand UO_181 (O_181,N_4118,N_4062);
nand UO_182 (O_182,N_4795,N_4574);
nor UO_183 (O_183,N_4060,N_4529);
and UO_184 (O_184,N_4188,N_4258);
and UO_185 (O_185,N_4649,N_4340);
and UO_186 (O_186,N_4486,N_4672);
or UO_187 (O_187,N_4298,N_4488);
or UO_188 (O_188,N_4055,N_4098);
and UO_189 (O_189,N_4119,N_4727);
and UO_190 (O_190,N_4718,N_4049);
nand UO_191 (O_191,N_4367,N_4697);
and UO_192 (O_192,N_4969,N_4498);
and UO_193 (O_193,N_4090,N_4089);
and UO_194 (O_194,N_4811,N_4133);
and UO_195 (O_195,N_4821,N_4645);
or UO_196 (O_196,N_4792,N_4986);
or UO_197 (O_197,N_4481,N_4802);
nor UO_198 (O_198,N_4072,N_4256);
nor UO_199 (O_199,N_4878,N_4624);
or UO_200 (O_200,N_4465,N_4235);
nor UO_201 (O_201,N_4370,N_4257);
and UO_202 (O_202,N_4043,N_4180);
nand UO_203 (O_203,N_4739,N_4521);
or UO_204 (O_204,N_4163,N_4197);
nand UO_205 (O_205,N_4956,N_4294);
nand UO_206 (O_206,N_4037,N_4001);
and UO_207 (O_207,N_4127,N_4944);
nor UO_208 (O_208,N_4646,N_4777);
nor UO_209 (O_209,N_4150,N_4306);
nor UO_210 (O_210,N_4686,N_4219);
and UO_211 (O_211,N_4161,N_4117);
nand UO_212 (O_212,N_4762,N_4183);
or UO_213 (O_213,N_4036,N_4805);
nor UO_214 (O_214,N_4319,N_4050);
nor UO_215 (O_215,N_4137,N_4559);
or UO_216 (O_216,N_4555,N_4543);
and UO_217 (O_217,N_4872,N_4041);
nand UO_218 (O_218,N_4082,N_4704);
or UO_219 (O_219,N_4125,N_4224);
nand UO_220 (O_220,N_4917,N_4884);
nand UO_221 (O_221,N_4829,N_4589);
and UO_222 (O_222,N_4215,N_4386);
and UO_223 (O_223,N_4943,N_4820);
nor UO_224 (O_224,N_4615,N_4754);
and UO_225 (O_225,N_4111,N_4293);
nand UO_226 (O_226,N_4924,N_4042);
or UO_227 (O_227,N_4676,N_4019);
nor UO_228 (O_228,N_4560,N_4549);
and UO_229 (O_229,N_4617,N_4415);
nor UO_230 (O_230,N_4904,N_4816);
nand UO_231 (O_231,N_4722,N_4532);
or UO_232 (O_232,N_4669,N_4911);
nand UO_233 (O_233,N_4130,N_4474);
and UO_234 (O_234,N_4101,N_4663);
nand UO_235 (O_235,N_4422,N_4579);
or UO_236 (O_236,N_4583,N_4894);
nand UO_237 (O_237,N_4656,N_4140);
nand UO_238 (O_238,N_4031,N_4453);
and UO_239 (O_239,N_4945,N_4973);
and UO_240 (O_240,N_4155,N_4842);
nand UO_241 (O_241,N_4591,N_4791);
nand UO_242 (O_242,N_4914,N_4918);
and UO_243 (O_243,N_4352,N_4761);
and UO_244 (O_244,N_4375,N_4580);
or UO_245 (O_245,N_4833,N_4205);
and UO_246 (O_246,N_4869,N_4017);
nand UO_247 (O_247,N_4296,N_4469);
nand UO_248 (O_248,N_4936,N_4974);
and UO_249 (O_249,N_4040,N_4123);
and UO_250 (O_250,N_4351,N_4614);
and UO_251 (O_251,N_4326,N_4423);
and UO_252 (O_252,N_4750,N_4994);
nand UO_253 (O_253,N_4259,N_4510);
and UO_254 (O_254,N_4499,N_4726);
nor UO_255 (O_255,N_4109,N_4922);
nand UO_256 (O_256,N_4558,N_4503);
nor UO_257 (O_257,N_4364,N_4288);
and UO_258 (O_258,N_4154,N_4901);
or UO_259 (O_259,N_4292,N_4737);
or UO_260 (O_260,N_4514,N_4931);
nor UO_261 (O_261,N_4241,N_4753);
nor UO_262 (O_262,N_4550,N_4557);
nand UO_263 (O_263,N_4832,N_4394);
nand UO_264 (O_264,N_4670,N_4020);
nor UO_265 (O_265,N_4975,N_4540);
nand UO_266 (O_266,N_4179,N_4586);
nand UO_267 (O_267,N_4442,N_4769);
and UO_268 (O_268,N_4815,N_4333);
or UO_269 (O_269,N_4530,N_4497);
and UO_270 (O_270,N_4220,N_4343);
nand UO_271 (O_271,N_4584,N_4186);
and UO_272 (O_272,N_4131,N_4518);
or UO_273 (O_273,N_4747,N_4399);
and UO_274 (O_274,N_4809,N_4695);
nor UO_275 (O_275,N_4160,N_4823);
nor UO_276 (O_276,N_4269,N_4071);
nor UO_277 (O_277,N_4966,N_4039);
and UO_278 (O_278,N_4954,N_4929);
and UO_279 (O_279,N_4248,N_4594);
nor UO_280 (O_280,N_4522,N_4251);
or UO_281 (O_281,N_4736,N_4942);
or UO_282 (O_282,N_4159,N_4102);
and UO_283 (O_283,N_4433,N_4124);
nor UO_284 (O_284,N_4282,N_4211);
nand UO_285 (O_285,N_4581,N_4988);
nor UO_286 (O_286,N_4011,N_4983);
nand UO_287 (O_287,N_4607,N_4312);
or UO_288 (O_288,N_4206,N_4709);
nor UO_289 (O_289,N_4112,N_4246);
nor UO_290 (O_290,N_4024,N_4511);
or UO_291 (O_291,N_4618,N_4412);
nor UO_292 (O_292,N_4088,N_4537);
nor UO_293 (O_293,N_4680,N_4026);
nor UO_294 (O_294,N_4323,N_4411);
xor UO_295 (O_295,N_4245,N_4184);
nor UO_296 (O_296,N_4278,N_4227);
or UO_297 (O_297,N_4992,N_4509);
nor UO_298 (O_298,N_4172,N_4078);
nor UO_299 (O_299,N_4881,N_4556);
nand UO_300 (O_300,N_4830,N_4413);
nor UO_301 (O_301,N_4712,N_4662);
nor UO_302 (O_302,N_4377,N_4673);
or UO_303 (O_303,N_4027,N_4776);
nor UO_304 (O_304,N_4057,N_4900);
or UO_305 (O_305,N_4950,N_4485);
nor UO_306 (O_306,N_4757,N_4252);
or UO_307 (O_307,N_4606,N_4470);
nand UO_308 (O_308,N_4652,N_4865);
and UO_309 (O_309,N_4597,N_4193);
nand UO_310 (O_310,N_4303,N_4857);
nand UO_311 (O_311,N_4493,N_4570);
nand UO_312 (O_312,N_4167,N_4237);
or UO_313 (O_313,N_4625,N_4700);
and UO_314 (O_314,N_4240,N_4477);
nor UO_315 (O_315,N_4084,N_4970);
nand UO_316 (O_316,N_4655,N_4743);
nand UO_317 (O_317,N_4203,N_4169);
and UO_318 (O_318,N_4682,N_4262);
nand UO_319 (O_319,N_4609,N_4177);
and UO_320 (O_320,N_4705,N_4642);
and UO_321 (O_321,N_4685,N_4314);
and UO_322 (O_322,N_4059,N_4796);
nor UO_323 (O_323,N_4838,N_4291);
nand UO_324 (O_324,N_4176,N_4780);
or UO_325 (O_325,N_4033,N_4301);
and UO_326 (O_326,N_4281,N_4304);
or UO_327 (O_327,N_4139,N_4483);
or UO_328 (O_328,N_4804,N_4004);
xnor UO_329 (O_329,N_4468,N_4864);
nand UO_330 (O_330,N_4906,N_4378);
and UO_331 (O_331,N_4603,N_4907);
nor UO_332 (O_332,N_4568,N_4103);
or UO_333 (O_333,N_4693,N_4368);
nand UO_334 (O_334,N_4178,N_4320);
or UO_335 (O_335,N_4601,N_4859);
and UO_336 (O_336,N_4476,N_4342);
nor UO_337 (O_337,N_4436,N_4714);
nor UO_338 (O_338,N_4051,N_4452);
or UO_339 (O_339,N_4998,N_4659);
nand UO_340 (O_340,N_4234,N_4496);
and UO_341 (O_341,N_4387,N_4926);
or UO_342 (O_342,N_4851,N_4209);
nor UO_343 (O_343,N_4858,N_4965);
xnor UO_344 (O_344,N_4775,N_4299);
and UO_345 (O_345,N_4723,N_4380);
and UO_346 (O_346,N_4035,N_4063);
or UO_347 (O_347,N_4751,N_4643);
nor UO_348 (O_348,N_4960,N_4135);
and UO_349 (O_349,N_4455,N_4637);
nand UO_350 (O_350,N_4787,N_4631);
nor UO_351 (O_351,N_4623,N_4070);
and UO_352 (O_352,N_4207,N_4822);
nand UO_353 (O_353,N_4198,N_4853);
and UO_354 (O_354,N_4725,N_4153);
nor UO_355 (O_355,N_4463,N_4405);
nor UO_356 (O_356,N_4385,N_4494);
and UO_357 (O_357,N_4047,N_4285);
or UO_358 (O_358,N_4632,N_4554);
nor UO_359 (O_359,N_4640,N_4048);
and UO_360 (O_360,N_4414,N_4318);
nor UO_361 (O_361,N_4266,N_4428);
nand UO_362 (O_362,N_4357,N_4250);
nor UO_363 (O_363,N_4267,N_4275);
or UO_364 (O_364,N_4692,N_4322);
and UO_365 (O_365,N_4947,N_4327);
nor UO_366 (O_366,N_4993,N_4844);
or UO_367 (O_367,N_4046,N_4243);
and UO_368 (O_368,N_4196,N_4236);
or UO_369 (O_369,N_4962,N_4290);
nor UO_370 (O_370,N_4995,N_4091);
and UO_371 (O_371,N_4080,N_4454);
nor UO_372 (O_372,N_4287,N_4408);
nand UO_373 (O_373,N_4097,N_4567);
and UO_374 (O_374,N_4075,N_4641);
nor UO_375 (O_375,N_4677,N_4507);
nand UO_376 (O_376,N_4773,N_4007);
and UO_377 (O_377,N_4501,N_4908);
nor UO_378 (O_378,N_4996,N_4935);
or UO_379 (O_379,N_4495,N_4136);
nor UO_380 (O_380,N_4621,N_4114);
and UO_381 (O_381,N_4410,N_4142);
nor UO_382 (O_382,N_4200,N_4400);
and UO_383 (O_383,N_4576,N_4023);
nor UO_384 (O_384,N_4980,N_4069);
nor UO_385 (O_385,N_4429,N_4536);
nand UO_386 (O_386,N_4616,N_4143);
xnor UO_387 (O_387,N_4157,N_4110);
nand UO_388 (O_388,N_4030,N_4887);
and UO_389 (O_389,N_4445,N_4562);
nand UO_390 (O_390,N_4721,N_4276);
or UO_391 (O_391,N_4191,N_4383);
nor UO_392 (O_392,N_4633,N_4430);
nor UO_393 (O_393,N_4458,N_4600);
or UO_394 (O_394,N_4971,N_4748);
or UO_395 (O_395,N_4541,N_4438);
nand UO_396 (O_396,N_4571,N_4347);
and UO_397 (O_397,N_4587,N_4145);
nor UO_398 (O_398,N_4528,N_4706);
nand UO_399 (O_399,N_4595,N_4981);
nand UO_400 (O_400,N_4003,N_4381);
nor UO_401 (O_401,N_4389,N_4746);
or UO_402 (O_402,N_4667,N_4825);
nor UO_403 (O_403,N_4134,N_4443);
nand UO_404 (O_404,N_4316,N_4527);
or UO_405 (O_405,N_4337,N_4190);
nand UO_406 (O_406,N_4391,N_4925);
nand UO_407 (O_407,N_4328,N_4877);
or UO_408 (O_408,N_4489,N_4895);
xor UO_409 (O_409,N_4092,N_4897);
and UO_410 (O_410,N_4875,N_4849);
and UO_411 (O_411,N_4073,N_4698);
nand UO_412 (O_412,N_4297,N_4382);
nor UO_413 (O_413,N_4690,N_4856);
nand UO_414 (O_414,N_4898,N_4064);
and UO_415 (O_415,N_4715,N_4916);
nor UO_416 (O_416,N_4397,N_4593);
or UO_417 (O_417,N_4940,N_4350);
or UO_418 (O_418,N_4151,N_4480);
nand UO_419 (O_419,N_4968,N_4921);
and UO_420 (O_420,N_4977,N_4416);
and UO_421 (O_421,N_4086,N_4660);
nand UO_422 (O_422,N_4744,N_4341);
nand UO_423 (O_423,N_4903,N_4784);
nor UO_424 (O_424,N_4345,N_4578);
nor UO_425 (O_425,N_4738,N_4305);
xnor UO_426 (O_426,N_4270,N_4961);
and UO_427 (O_427,N_4289,N_4512);
or UO_428 (O_428,N_4168,N_4253);
and UO_429 (O_429,N_4471,N_4933);
or UO_430 (O_430,N_4010,N_4654);
nor UO_431 (O_431,N_4517,N_4302);
nand UO_432 (O_432,N_4388,N_4915);
and UO_433 (O_433,N_4783,N_4569);
and UO_434 (O_434,N_4817,N_4194);
nor UO_435 (O_435,N_4789,N_4214);
nor UO_436 (O_436,N_4604,N_4702);
or UO_437 (O_437,N_4689,N_4313);
and UO_438 (O_438,N_4479,N_4425);
and UO_439 (O_439,N_4446,N_4733);
nor UO_440 (O_440,N_4018,N_4166);
nand UO_441 (O_441,N_4447,N_4666);
nor UO_442 (O_442,N_4034,N_4478);
nand UO_443 (O_443,N_4346,N_4939);
nor UO_444 (O_444,N_4674,N_4610);
and UO_445 (O_445,N_4812,N_4195);
or UO_446 (O_446,N_4053,N_4348);
and UO_447 (O_447,N_4356,N_4928);
nor UO_448 (O_448,N_4335,N_4785);
nand UO_449 (O_449,N_4331,N_4871);
nor UO_450 (O_450,N_4120,N_4464);
nor UO_451 (O_451,N_4440,N_4058);
and UO_452 (O_452,N_4840,N_4221);
nor UO_453 (O_453,N_4272,N_4449);
or UO_454 (O_454,N_4052,N_4015);
or UO_455 (O_455,N_4539,N_4899);
and UO_456 (O_456,N_4279,N_4749);
nor UO_457 (O_457,N_4152,N_4565);
and UO_458 (O_458,N_4126,N_4149);
and UO_459 (O_459,N_4100,N_4009);
or UO_460 (O_460,N_4880,N_4573);
nand UO_461 (O_461,N_4909,N_4760);
or UO_462 (O_462,N_4325,N_4431);
nor UO_463 (O_463,N_4132,N_4552);
nand UO_464 (O_464,N_4848,N_4115);
nor UO_465 (O_465,N_4687,N_4912);
nor UO_466 (O_466,N_4719,N_4274);
nand UO_467 (O_467,N_4173,N_4696);
nand UO_468 (O_468,N_4366,N_4264);
nand UO_469 (O_469,N_4372,N_4592);
and UO_470 (O_470,N_4635,N_4806);
and UO_471 (O_471,N_4353,N_4295);
and UO_472 (O_472,N_4644,N_4516);
xor UO_473 (O_473,N_4905,N_4577);
or UO_474 (O_474,N_4630,N_4523);
nand UO_475 (O_475,N_4708,N_4515);
and UO_476 (O_476,N_4358,N_4834);
or UO_477 (O_477,N_4651,N_4212);
nand UO_478 (O_478,N_4572,N_4456);
and UO_479 (O_479,N_4538,N_4146);
or UO_480 (O_480,N_4937,N_4192);
and UO_481 (O_481,N_4332,N_4189);
nand UO_482 (O_482,N_4839,N_4029);
and UO_483 (O_483,N_4957,N_4360);
nand UO_484 (O_484,N_4461,N_4334);
and UO_485 (O_485,N_4803,N_4835);
nor UO_486 (O_486,N_4164,N_4002);
and UO_487 (O_487,N_4401,N_4657);
or UO_488 (O_488,N_4460,N_4941);
nor UO_489 (O_489,N_4524,N_4588);
or UO_490 (O_490,N_4085,N_4384);
or UO_491 (O_491,N_4217,N_4613);
nor UO_492 (O_492,N_4845,N_4694);
and UO_493 (O_493,N_4650,N_4247);
and UO_494 (O_494,N_4826,N_4148);
nand UO_495 (O_495,N_4056,N_4105);
or UO_496 (O_496,N_4768,N_4255);
nand UO_497 (O_497,N_4006,N_4890);
or UO_498 (O_498,N_4421,N_4174);
nand UO_499 (O_499,N_4068,N_4165);
nand UO_500 (O_500,N_4862,N_4454);
nand UO_501 (O_501,N_4006,N_4138);
nor UO_502 (O_502,N_4089,N_4796);
and UO_503 (O_503,N_4238,N_4763);
or UO_504 (O_504,N_4851,N_4401);
nor UO_505 (O_505,N_4839,N_4542);
and UO_506 (O_506,N_4146,N_4390);
and UO_507 (O_507,N_4232,N_4195);
nand UO_508 (O_508,N_4152,N_4103);
nand UO_509 (O_509,N_4723,N_4776);
nor UO_510 (O_510,N_4784,N_4416);
or UO_511 (O_511,N_4832,N_4190);
nand UO_512 (O_512,N_4317,N_4613);
or UO_513 (O_513,N_4828,N_4659);
nor UO_514 (O_514,N_4939,N_4754);
and UO_515 (O_515,N_4246,N_4374);
nand UO_516 (O_516,N_4911,N_4888);
nor UO_517 (O_517,N_4392,N_4560);
nand UO_518 (O_518,N_4181,N_4941);
and UO_519 (O_519,N_4337,N_4531);
and UO_520 (O_520,N_4123,N_4318);
and UO_521 (O_521,N_4770,N_4756);
nor UO_522 (O_522,N_4903,N_4735);
nor UO_523 (O_523,N_4753,N_4934);
nand UO_524 (O_524,N_4706,N_4140);
nor UO_525 (O_525,N_4226,N_4088);
and UO_526 (O_526,N_4205,N_4989);
nand UO_527 (O_527,N_4987,N_4101);
nor UO_528 (O_528,N_4927,N_4970);
nor UO_529 (O_529,N_4145,N_4190);
and UO_530 (O_530,N_4415,N_4726);
and UO_531 (O_531,N_4733,N_4145);
and UO_532 (O_532,N_4915,N_4800);
and UO_533 (O_533,N_4887,N_4946);
nor UO_534 (O_534,N_4223,N_4157);
and UO_535 (O_535,N_4020,N_4721);
nor UO_536 (O_536,N_4187,N_4018);
or UO_537 (O_537,N_4375,N_4121);
nor UO_538 (O_538,N_4029,N_4261);
nand UO_539 (O_539,N_4285,N_4735);
nor UO_540 (O_540,N_4332,N_4464);
nor UO_541 (O_541,N_4014,N_4642);
or UO_542 (O_542,N_4055,N_4158);
nand UO_543 (O_543,N_4743,N_4015);
or UO_544 (O_544,N_4533,N_4484);
and UO_545 (O_545,N_4775,N_4612);
nor UO_546 (O_546,N_4345,N_4564);
nand UO_547 (O_547,N_4581,N_4138);
nor UO_548 (O_548,N_4629,N_4966);
and UO_549 (O_549,N_4452,N_4837);
and UO_550 (O_550,N_4180,N_4839);
or UO_551 (O_551,N_4485,N_4870);
nand UO_552 (O_552,N_4078,N_4955);
nor UO_553 (O_553,N_4774,N_4791);
nand UO_554 (O_554,N_4165,N_4573);
and UO_555 (O_555,N_4360,N_4168);
or UO_556 (O_556,N_4011,N_4835);
and UO_557 (O_557,N_4073,N_4129);
nand UO_558 (O_558,N_4916,N_4658);
nand UO_559 (O_559,N_4657,N_4176);
nand UO_560 (O_560,N_4888,N_4095);
or UO_561 (O_561,N_4815,N_4807);
or UO_562 (O_562,N_4603,N_4953);
nand UO_563 (O_563,N_4164,N_4023);
nor UO_564 (O_564,N_4843,N_4599);
and UO_565 (O_565,N_4121,N_4843);
or UO_566 (O_566,N_4983,N_4919);
or UO_567 (O_567,N_4469,N_4508);
and UO_568 (O_568,N_4461,N_4858);
nand UO_569 (O_569,N_4715,N_4910);
nand UO_570 (O_570,N_4488,N_4793);
or UO_571 (O_571,N_4478,N_4338);
nand UO_572 (O_572,N_4055,N_4111);
and UO_573 (O_573,N_4533,N_4414);
and UO_574 (O_574,N_4702,N_4363);
nand UO_575 (O_575,N_4245,N_4373);
nand UO_576 (O_576,N_4728,N_4796);
and UO_577 (O_577,N_4707,N_4576);
or UO_578 (O_578,N_4940,N_4734);
or UO_579 (O_579,N_4982,N_4124);
and UO_580 (O_580,N_4222,N_4308);
nor UO_581 (O_581,N_4126,N_4735);
or UO_582 (O_582,N_4456,N_4512);
or UO_583 (O_583,N_4605,N_4804);
nand UO_584 (O_584,N_4695,N_4108);
and UO_585 (O_585,N_4281,N_4105);
nand UO_586 (O_586,N_4274,N_4142);
or UO_587 (O_587,N_4729,N_4762);
and UO_588 (O_588,N_4020,N_4555);
or UO_589 (O_589,N_4457,N_4847);
and UO_590 (O_590,N_4010,N_4559);
nand UO_591 (O_591,N_4156,N_4195);
nand UO_592 (O_592,N_4886,N_4025);
nor UO_593 (O_593,N_4832,N_4012);
or UO_594 (O_594,N_4143,N_4868);
and UO_595 (O_595,N_4078,N_4261);
or UO_596 (O_596,N_4091,N_4280);
or UO_597 (O_597,N_4103,N_4995);
or UO_598 (O_598,N_4009,N_4595);
or UO_599 (O_599,N_4229,N_4617);
and UO_600 (O_600,N_4445,N_4127);
nor UO_601 (O_601,N_4597,N_4558);
nor UO_602 (O_602,N_4064,N_4458);
or UO_603 (O_603,N_4001,N_4231);
or UO_604 (O_604,N_4467,N_4893);
or UO_605 (O_605,N_4031,N_4177);
nand UO_606 (O_606,N_4837,N_4343);
and UO_607 (O_607,N_4209,N_4950);
or UO_608 (O_608,N_4222,N_4041);
and UO_609 (O_609,N_4252,N_4509);
nor UO_610 (O_610,N_4095,N_4001);
nand UO_611 (O_611,N_4770,N_4217);
nor UO_612 (O_612,N_4457,N_4697);
nor UO_613 (O_613,N_4141,N_4872);
nor UO_614 (O_614,N_4158,N_4964);
and UO_615 (O_615,N_4650,N_4691);
nand UO_616 (O_616,N_4715,N_4606);
and UO_617 (O_617,N_4420,N_4006);
nand UO_618 (O_618,N_4525,N_4879);
nand UO_619 (O_619,N_4868,N_4580);
nand UO_620 (O_620,N_4483,N_4178);
and UO_621 (O_621,N_4644,N_4988);
and UO_622 (O_622,N_4112,N_4641);
and UO_623 (O_623,N_4135,N_4832);
nand UO_624 (O_624,N_4121,N_4875);
nand UO_625 (O_625,N_4877,N_4699);
nand UO_626 (O_626,N_4131,N_4469);
or UO_627 (O_627,N_4027,N_4735);
nor UO_628 (O_628,N_4769,N_4725);
nand UO_629 (O_629,N_4386,N_4980);
xnor UO_630 (O_630,N_4487,N_4361);
or UO_631 (O_631,N_4499,N_4225);
or UO_632 (O_632,N_4886,N_4949);
and UO_633 (O_633,N_4819,N_4409);
nor UO_634 (O_634,N_4847,N_4866);
nor UO_635 (O_635,N_4040,N_4522);
or UO_636 (O_636,N_4776,N_4913);
and UO_637 (O_637,N_4313,N_4475);
or UO_638 (O_638,N_4442,N_4975);
and UO_639 (O_639,N_4745,N_4993);
xnor UO_640 (O_640,N_4105,N_4253);
and UO_641 (O_641,N_4080,N_4582);
and UO_642 (O_642,N_4226,N_4235);
or UO_643 (O_643,N_4672,N_4122);
and UO_644 (O_644,N_4254,N_4992);
or UO_645 (O_645,N_4961,N_4403);
nor UO_646 (O_646,N_4761,N_4181);
nor UO_647 (O_647,N_4697,N_4393);
or UO_648 (O_648,N_4215,N_4796);
nand UO_649 (O_649,N_4938,N_4948);
and UO_650 (O_650,N_4976,N_4751);
or UO_651 (O_651,N_4021,N_4742);
or UO_652 (O_652,N_4020,N_4991);
nand UO_653 (O_653,N_4654,N_4623);
nand UO_654 (O_654,N_4833,N_4159);
and UO_655 (O_655,N_4010,N_4981);
nor UO_656 (O_656,N_4004,N_4230);
and UO_657 (O_657,N_4816,N_4377);
nor UO_658 (O_658,N_4708,N_4946);
nand UO_659 (O_659,N_4685,N_4000);
or UO_660 (O_660,N_4514,N_4868);
or UO_661 (O_661,N_4819,N_4909);
nand UO_662 (O_662,N_4511,N_4095);
and UO_663 (O_663,N_4546,N_4896);
nand UO_664 (O_664,N_4542,N_4715);
or UO_665 (O_665,N_4198,N_4580);
nor UO_666 (O_666,N_4133,N_4250);
nand UO_667 (O_667,N_4070,N_4594);
nor UO_668 (O_668,N_4557,N_4620);
and UO_669 (O_669,N_4408,N_4038);
and UO_670 (O_670,N_4538,N_4156);
nand UO_671 (O_671,N_4202,N_4540);
nand UO_672 (O_672,N_4066,N_4102);
nand UO_673 (O_673,N_4684,N_4398);
and UO_674 (O_674,N_4986,N_4595);
nor UO_675 (O_675,N_4551,N_4462);
and UO_676 (O_676,N_4583,N_4334);
nand UO_677 (O_677,N_4470,N_4999);
nand UO_678 (O_678,N_4017,N_4671);
nor UO_679 (O_679,N_4207,N_4453);
and UO_680 (O_680,N_4057,N_4697);
or UO_681 (O_681,N_4169,N_4483);
or UO_682 (O_682,N_4325,N_4856);
nand UO_683 (O_683,N_4752,N_4854);
nand UO_684 (O_684,N_4858,N_4293);
or UO_685 (O_685,N_4634,N_4640);
and UO_686 (O_686,N_4668,N_4406);
and UO_687 (O_687,N_4223,N_4983);
nor UO_688 (O_688,N_4997,N_4388);
and UO_689 (O_689,N_4456,N_4752);
and UO_690 (O_690,N_4852,N_4373);
nor UO_691 (O_691,N_4735,N_4634);
nor UO_692 (O_692,N_4997,N_4419);
and UO_693 (O_693,N_4100,N_4704);
and UO_694 (O_694,N_4076,N_4720);
nand UO_695 (O_695,N_4829,N_4471);
xnor UO_696 (O_696,N_4237,N_4069);
nand UO_697 (O_697,N_4556,N_4378);
and UO_698 (O_698,N_4455,N_4118);
xor UO_699 (O_699,N_4893,N_4412);
nor UO_700 (O_700,N_4465,N_4969);
or UO_701 (O_701,N_4144,N_4913);
or UO_702 (O_702,N_4765,N_4683);
or UO_703 (O_703,N_4552,N_4577);
or UO_704 (O_704,N_4916,N_4706);
and UO_705 (O_705,N_4259,N_4158);
or UO_706 (O_706,N_4980,N_4221);
or UO_707 (O_707,N_4166,N_4148);
nor UO_708 (O_708,N_4116,N_4128);
or UO_709 (O_709,N_4581,N_4427);
nor UO_710 (O_710,N_4331,N_4003);
or UO_711 (O_711,N_4030,N_4368);
nand UO_712 (O_712,N_4261,N_4796);
and UO_713 (O_713,N_4180,N_4726);
and UO_714 (O_714,N_4109,N_4856);
and UO_715 (O_715,N_4919,N_4748);
or UO_716 (O_716,N_4571,N_4123);
nand UO_717 (O_717,N_4277,N_4316);
xor UO_718 (O_718,N_4973,N_4020);
or UO_719 (O_719,N_4213,N_4339);
and UO_720 (O_720,N_4088,N_4364);
nand UO_721 (O_721,N_4610,N_4785);
or UO_722 (O_722,N_4072,N_4764);
or UO_723 (O_723,N_4899,N_4511);
or UO_724 (O_724,N_4254,N_4040);
or UO_725 (O_725,N_4354,N_4372);
nor UO_726 (O_726,N_4750,N_4068);
nand UO_727 (O_727,N_4034,N_4473);
and UO_728 (O_728,N_4476,N_4487);
or UO_729 (O_729,N_4185,N_4047);
nor UO_730 (O_730,N_4459,N_4946);
nand UO_731 (O_731,N_4817,N_4522);
nor UO_732 (O_732,N_4450,N_4802);
or UO_733 (O_733,N_4931,N_4821);
or UO_734 (O_734,N_4562,N_4985);
or UO_735 (O_735,N_4848,N_4546);
or UO_736 (O_736,N_4733,N_4036);
and UO_737 (O_737,N_4569,N_4804);
and UO_738 (O_738,N_4517,N_4415);
nand UO_739 (O_739,N_4778,N_4956);
nand UO_740 (O_740,N_4689,N_4020);
or UO_741 (O_741,N_4729,N_4933);
nor UO_742 (O_742,N_4561,N_4058);
or UO_743 (O_743,N_4650,N_4601);
nand UO_744 (O_744,N_4284,N_4580);
or UO_745 (O_745,N_4771,N_4660);
and UO_746 (O_746,N_4632,N_4336);
nand UO_747 (O_747,N_4701,N_4262);
or UO_748 (O_748,N_4943,N_4560);
or UO_749 (O_749,N_4061,N_4877);
or UO_750 (O_750,N_4013,N_4142);
nand UO_751 (O_751,N_4728,N_4361);
nor UO_752 (O_752,N_4100,N_4515);
nor UO_753 (O_753,N_4936,N_4947);
nand UO_754 (O_754,N_4345,N_4384);
and UO_755 (O_755,N_4623,N_4179);
or UO_756 (O_756,N_4271,N_4060);
nor UO_757 (O_757,N_4872,N_4556);
nor UO_758 (O_758,N_4118,N_4525);
nor UO_759 (O_759,N_4283,N_4447);
nand UO_760 (O_760,N_4214,N_4727);
or UO_761 (O_761,N_4995,N_4911);
nor UO_762 (O_762,N_4785,N_4476);
and UO_763 (O_763,N_4722,N_4745);
nand UO_764 (O_764,N_4671,N_4220);
nand UO_765 (O_765,N_4679,N_4967);
nor UO_766 (O_766,N_4305,N_4216);
and UO_767 (O_767,N_4520,N_4256);
nor UO_768 (O_768,N_4601,N_4858);
nand UO_769 (O_769,N_4934,N_4434);
nand UO_770 (O_770,N_4489,N_4103);
nor UO_771 (O_771,N_4779,N_4815);
and UO_772 (O_772,N_4128,N_4523);
nand UO_773 (O_773,N_4898,N_4184);
nor UO_774 (O_774,N_4997,N_4735);
or UO_775 (O_775,N_4114,N_4314);
nor UO_776 (O_776,N_4880,N_4168);
nand UO_777 (O_777,N_4203,N_4451);
nor UO_778 (O_778,N_4850,N_4708);
nand UO_779 (O_779,N_4734,N_4362);
nand UO_780 (O_780,N_4648,N_4819);
and UO_781 (O_781,N_4655,N_4756);
nand UO_782 (O_782,N_4397,N_4018);
nand UO_783 (O_783,N_4847,N_4738);
or UO_784 (O_784,N_4915,N_4106);
nor UO_785 (O_785,N_4460,N_4123);
or UO_786 (O_786,N_4274,N_4403);
nor UO_787 (O_787,N_4528,N_4458);
and UO_788 (O_788,N_4927,N_4809);
nor UO_789 (O_789,N_4333,N_4335);
and UO_790 (O_790,N_4996,N_4481);
or UO_791 (O_791,N_4531,N_4911);
nand UO_792 (O_792,N_4753,N_4794);
and UO_793 (O_793,N_4996,N_4887);
nand UO_794 (O_794,N_4059,N_4149);
nor UO_795 (O_795,N_4806,N_4326);
and UO_796 (O_796,N_4069,N_4473);
and UO_797 (O_797,N_4497,N_4800);
and UO_798 (O_798,N_4735,N_4509);
nand UO_799 (O_799,N_4364,N_4846);
nor UO_800 (O_800,N_4868,N_4133);
or UO_801 (O_801,N_4565,N_4506);
nand UO_802 (O_802,N_4604,N_4795);
or UO_803 (O_803,N_4208,N_4267);
or UO_804 (O_804,N_4673,N_4505);
and UO_805 (O_805,N_4380,N_4534);
nor UO_806 (O_806,N_4756,N_4554);
and UO_807 (O_807,N_4143,N_4167);
or UO_808 (O_808,N_4978,N_4572);
and UO_809 (O_809,N_4531,N_4891);
nand UO_810 (O_810,N_4211,N_4608);
and UO_811 (O_811,N_4594,N_4711);
and UO_812 (O_812,N_4312,N_4174);
or UO_813 (O_813,N_4034,N_4746);
nand UO_814 (O_814,N_4990,N_4828);
and UO_815 (O_815,N_4467,N_4398);
or UO_816 (O_816,N_4628,N_4073);
and UO_817 (O_817,N_4070,N_4888);
and UO_818 (O_818,N_4825,N_4774);
xnor UO_819 (O_819,N_4603,N_4214);
nor UO_820 (O_820,N_4728,N_4916);
nand UO_821 (O_821,N_4629,N_4769);
or UO_822 (O_822,N_4996,N_4817);
nand UO_823 (O_823,N_4855,N_4127);
nor UO_824 (O_824,N_4939,N_4865);
nand UO_825 (O_825,N_4509,N_4774);
or UO_826 (O_826,N_4560,N_4675);
and UO_827 (O_827,N_4967,N_4196);
nor UO_828 (O_828,N_4738,N_4072);
and UO_829 (O_829,N_4127,N_4999);
nor UO_830 (O_830,N_4005,N_4716);
and UO_831 (O_831,N_4616,N_4693);
nand UO_832 (O_832,N_4731,N_4333);
or UO_833 (O_833,N_4201,N_4804);
or UO_834 (O_834,N_4938,N_4015);
or UO_835 (O_835,N_4028,N_4428);
or UO_836 (O_836,N_4848,N_4802);
or UO_837 (O_837,N_4927,N_4923);
or UO_838 (O_838,N_4895,N_4061);
or UO_839 (O_839,N_4683,N_4123);
nand UO_840 (O_840,N_4810,N_4315);
nand UO_841 (O_841,N_4940,N_4652);
and UO_842 (O_842,N_4908,N_4449);
and UO_843 (O_843,N_4540,N_4084);
and UO_844 (O_844,N_4597,N_4194);
nand UO_845 (O_845,N_4705,N_4939);
or UO_846 (O_846,N_4335,N_4791);
nor UO_847 (O_847,N_4070,N_4266);
or UO_848 (O_848,N_4928,N_4088);
or UO_849 (O_849,N_4674,N_4758);
nand UO_850 (O_850,N_4653,N_4509);
or UO_851 (O_851,N_4882,N_4581);
nor UO_852 (O_852,N_4776,N_4879);
and UO_853 (O_853,N_4987,N_4300);
nand UO_854 (O_854,N_4286,N_4114);
nand UO_855 (O_855,N_4906,N_4519);
nor UO_856 (O_856,N_4454,N_4293);
nor UO_857 (O_857,N_4695,N_4749);
or UO_858 (O_858,N_4296,N_4498);
nand UO_859 (O_859,N_4037,N_4647);
and UO_860 (O_860,N_4001,N_4834);
or UO_861 (O_861,N_4937,N_4694);
or UO_862 (O_862,N_4722,N_4694);
nand UO_863 (O_863,N_4734,N_4688);
or UO_864 (O_864,N_4837,N_4115);
and UO_865 (O_865,N_4673,N_4264);
or UO_866 (O_866,N_4452,N_4264);
and UO_867 (O_867,N_4026,N_4740);
nand UO_868 (O_868,N_4916,N_4018);
and UO_869 (O_869,N_4653,N_4524);
nor UO_870 (O_870,N_4395,N_4628);
or UO_871 (O_871,N_4321,N_4064);
nor UO_872 (O_872,N_4503,N_4856);
or UO_873 (O_873,N_4414,N_4469);
and UO_874 (O_874,N_4257,N_4099);
or UO_875 (O_875,N_4253,N_4838);
or UO_876 (O_876,N_4961,N_4243);
nand UO_877 (O_877,N_4788,N_4559);
and UO_878 (O_878,N_4941,N_4463);
or UO_879 (O_879,N_4341,N_4353);
and UO_880 (O_880,N_4079,N_4792);
and UO_881 (O_881,N_4088,N_4215);
nor UO_882 (O_882,N_4347,N_4359);
and UO_883 (O_883,N_4755,N_4628);
or UO_884 (O_884,N_4016,N_4588);
and UO_885 (O_885,N_4301,N_4923);
and UO_886 (O_886,N_4577,N_4470);
nor UO_887 (O_887,N_4861,N_4237);
and UO_888 (O_888,N_4253,N_4757);
or UO_889 (O_889,N_4617,N_4427);
nor UO_890 (O_890,N_4114,N_4974);
nor UO_891 (O_891,N_4427,N_4544);
nand UO_892 (O_892,N_4871,N_4921);
nor UO_893 (O_893,N_4696,N_4910);
or UO_894 (O_894,N_4074,N_4984);
nand UO_895 (O_895,N_4836,N_4478);
nor UO_896 (O_896,N_4138,N_4941);
and UO_897 (O_897,N_4778,N_4693);
nor UO_898 (O_898,N_4815,N_4824);
nand UO_899 (O_899,N_4751,N_4204);
nand UO_900 (O_900,N_4908,N_4822);
and UO_901 (O_901,N_4867,N_4064);
nor UO_902 (O_902,N_4853,N_4558);
nand UO_903 (O_903,N_4572,N_4687);
nor UO_904 (O_904,N_4588,N_4736);
and UO_905 (O_905,N_4023,N_4803);
nor UO_906 (O_906,N_4378,N_4160);
nand UO_907 (O_907,N_4094,N_4034);
nor UO_908 (O_908,N_4186,N_4951);
and UO_909 (O_909,N_4079,N_4276);
or UO_910 (O_910,N_4987,N_4647);
and UO_911 (O_911,N_4320,N_4493);
and UO_912 (O_912,N_4646,N_4359);
and UO_913 (O_913,N_4840,N_4342);
or UO_914 (O_914,N_4401,N_4382);
or UO_915 (O_915,N_4083,N_4472);
or UO_916 (O_916,N_4332,N_4482);
and UO_917 (O_917,N_4351,N_4280);
and UO_918 (O_918,N_4010,N_4107);
or UO_919 (O_919,N_4143,N_4884);
or UO_920 (O_920,N_4085,N_4563);
nor UO_921 (O_921,N_4321,N_4929);
or UO_922 (O_922,N_4736,N_4287);
nand UO_923 (O_923,N_4736,N_4122);
nor UO_924 (O_924,N_4920,N_4784);
nor UO_925 (O_925,N_4953,N_4443);
and UO_926 (O_926,N_4573,N_4843);
or UO_927 (O_927,N_4472,N_4412);
and UO_928 (O_928,N_4030,N_4429);
or UO_929 (O_929,N_4213,N_4045);
nor UO_930 (O_930,N_4033,N_4840);
nor UO_931 (O_931,N_4512,N_4396);
nor UO_932 (O_932,N_4128,N_4557);
or UO_933 (O_933,N_4093,N_4296);
nand UO_934 (O_934,N_4286,N_4283);
or UO_935 (O_935,N_4641,N_4217);
and UO_936 (O_936,N_4115,N_4886);
and UO_937 (O_937,N_4718,N_4905);
nand UO_938 (O_938,N_4631,N_4707);
nand UO_939 (O_939,N_4648,N_4702);
nand UO_940 (O_940,N_4410,N_4765);
and UO_941 (O_941,N_4786,N_4009);
nand UO_942 (O_942,N_4413,N_4911);
or UO_943 (O_943,N_4061,N_4702);
nor UO_944 (O_944,N_4251,N_4468);
nand UO_945 (O_945,N_4251,N_4619);
and UO_946 (O_946,N_4960,N_4941);
or UO_947 (O_947,N_4204,N_4660);
nor UO_948 (O_948,N_4511,N_4957);
nand UO_949 (O_949,N_4530,N_4631);
nand UO_950 (O_950,N_4616,N_4937);
nor UO_951 (O_951,N_4860,N_4415);
and UO_952 (O_952,N_4394,N_4549);
or UO_953 (O_953,N_4937,N_4688);
nand UO_954 (O_954,N_4611,N_4536);
nor UO_955 (O_955,N_4911,N_4720);
nor UO_956 (O_956,N_4906,N_4872);
or UO_957 (O_957,N_4528,N_4213);
nor UO_958 (O_958,N_4709,N_4531);
nor UO_959 (O_959,N_4297,N_4084);
or UO_960 (O_960,N_4249,N_4177);
nand UO_961 (O_961,N_4145,N_4029);
nor UO_962 (O_962,N_4569,N_4875);
nor UO_963 (O_963,N_4154,N_4804);
or UO_964 (O_964,N_4384,N_4180);
and UO_965 (O_965,N_4457,N_4075);
or UO_966 (O_966,N_4926,N_4468);
nor UO_967 (O_967,N_4153,N_4998);
and UO_968 (O_968,N_4106,N_4022);
or UO_969 (O_969,N_4720,N_4187);
and UO_970 (O_970,N_4476,N_4656);
nor UO_971 (O_971,N_4258,N_4330);
nand UO_972 (O_972,N_4821,N_4372);
or UO_973 (O_973,N_4238,N_4627);
nor UO_974 (O_974,N_4205,N_4128);
and UO_975 (O_975,N_4823,N_4080);
nand UO_976 (O_976,N_4095,N_4469);
nand UO_977 (O_977,N_4965,N_4776);
or UO_978 (O_978,N_4535,N_4212);
or UO_979 (O_979,N_4371,N_4249);
and UO_980 (O_980,N_4079,N_4500);
nor UO_981 (O_981,N_4470,N_4413);
nor UO_982 (O_982,N_4581,N_4003);
and UO_983 (O_983,N_4490,N_4589);
or UO_984 (O_984,N_4773,N_4452);
nor UO_985 (O_985,N_4001,N_4662);
nor UO_986 (O_986,N_4684,N_4923);
and UO_987 (O_987,N_4825,N_4350);
nand UO_988 (O_988,N_4731,N_4986);
and UO_989 (O_989,N_4351,N_4982);
or UO_990 (O_990,N_4013,N_4441);
nor UO_991 (O_991,N_4132,N_4462);
nand UO_992 (O_992,N_4830,N_4727);
nor UO_993 (O_993,N_4996,N_4435);
or UO_994 (O_994,N_4184,N_4138);
nand UO_995 (O_995,N_4993,N_4079);
nor UO_996 (O_996,N_4777,N_4781);
nand UO_997 (O_997,N_4668,N_4545);
nand UO_998 (O_998,N_4289,N_4526);
and UO_999 (O_999,N_4255,N_4994);
endmodule