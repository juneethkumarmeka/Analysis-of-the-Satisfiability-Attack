module basic_1500_15000_2000_60_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_855,In_573);
nor U1 (N_1,In_338,In_1042);
xnor U2 (N_2,In_1273,In_1163);
or U3 (N_3,In_930,In_4);
or U4 (N_4,In_702,In_538);
or U5 (N_5,In_1387,In_931);
xnor U6 (N_6,In_360,In_1095);
nand U7 (N_7,In_946,In_762);
nand U8 (N_8,In_269,In_1074);
and U9 (N_9,In_381,In_178);
nand U10 (N_10,In_1106,In_172);
nand U11 (N_11,In_1253,In_694);
or U12 (N_12,In_242,In_1043);
and U13 (N_13,In_158,In_1378);
xor U14 (N_14,In_1499,In_549);
or U15 (N_15,In_1394,In_998);
nand U16 (N_16,In_0,In_728);
xnor U17 (N_17,In_128,In_143);
and U18 (N_18,In_30,In_847);
and U19 (N_19,In_357,In_1237);
nor U20 (N_20,In_699,In_590);
or U21 (N_21,In_1132,In_845);
and U22 (N_22,In_817,In_173);
nand U23 (N_23,In_480,In_92);
xnor U24 (N_24,In_1377,In_760);
and U25 (N_25,In_994,In_1017);
and U26 (N_26,In_1191,In_1137);
nand U27 (N_27,In_1103,In_955);
or U28 (N_28,In_595,In_1285);
and U29 (N_29,In_1458,In_33);
and U30 (N_30,In_616,In_96);
and U31 (N_31,In_28,In_1337);
nand U32 (N_32,In_112,In_816);
nand U33 (N_33,In_981,In_24);
or U34 (N_34,In_336,In_634);
or U35 (N_35,In_442,In_1482);
nand U36 (N_36,In_376,In_365);
nor U37 (N_37,In_505,In_471);
nand U38 (N_38,In_351,In_1466);
nand U39 (N_39,In_137,In_940);
and U40 (N_40,In_1369,In_753);
and U41 (N_41,In_1047,In_303);
nand U42 (N_42,In_77,In_1179);
xor U43 (N_43,In_990,In_222);
or U44 (N_44,In_316,In_240);
and U45 (N_45,In_718,In_514);
nor U46 (N_46,In_1399,In_36);
nand U47 (N_47,In_1052,In_1129);
or U48 (N_48,In_314,In_1321);
or U49 (N_49,In_1423,In_440);
xor U50 (N_50,In_770,In_65);
nand U51 (N_51,In_244,In_191);
nand U52 (N_52,In_315,In_127);
nor U53 (N_53,In_1157,In_181);
nand U54 (N_54,In_572,In_1371);
nand U55 (N_55,In_1242,In_1492);
or U56 (N_56,In_1488,In_182);
xnor U57 (N_57,In_796,In_900);
nand U58 (N_58,In_1214,In_526);
nor U59 (N_59,In_122,In_427);
nand U60 (N_60,In_783,In_246);
or U61 (N_61,In_1056,In_1083);
xnor U62 (N_62,In_742,In_767);
nand U63 (N_63,In_39,In_682);
nand U64 (N_64,In_1138,In_279);
nand U65 (N_65,In_424,In_152);
nor U66 (N_66,In_986,In_686);
nor U67 (N_67,In_693,In_1364);
and U68 (N_68,In_923,In_370);
or U69 (N_69,In_681,In_1353);
nand U70 (N_70,In_1155,In_287);
xnor U71 (N_71,In_993,In_547);
nor U72 (N_72,In_881,In_611);
xnor U73 (N_73,In_700,In_142);
xnor U74 (N_74,In_1101,In_899);
nor U75 (N_75,In_621,In_1235);
or U76 (N_76,In_1259,In_619);
and U77 (N_77,In_1325,In_679);
nand U78 (N_78,In_6,In_73);
and U79 (N_79,In_1421,In_1429);
and U80 (N_80,In_964,In_866);
and U81 (N_81,In_1339,In_1107);
xnor U82 (N_82,In_492,In_493);
and U83 (N_83,In_1049,In_443);
xor U84 (N_84,In_1055,In_667);
or U85 (N_85,In_1396,In_922);
nand U86 (N_86,In_130,In_482);
nor U87 (N_87,In_528,In_1301);
xor U88 (N_88,In_836,In_448);
and U89 (N_89,In_1463,In_1199);
nor U90 (N_90,In_620,In_1001);
or U91 (N_91,In_1197,In_456);
or U92 (N_92,In_985,In_1408);
nor U93 (N_93,In_614,In_1252);
xor U94 (N_94,In_1100,In_598);
nor U95 (N_95,In_856,In_459);
or U96 (N_96,In_221,In_974);
xnor U97 (N_97,In_632,In_730);
nor U98 (N_98,In_194,In_190);
and U99 (N_99,In_743,In_1334);
and U100 (N_100,In_1069,In_195);
xor U101 (N_101,In_1133,In_329);
nand U102 (N_102,In_685,In_476);
or U103 (N_103,In_1119,In_1355);
and U104 (N_104,In_59,In_1067);
nor U105 (N_105,In_826,In_987);
nand U106 (N_106,In_466,In_1306);
xnor U107 (N_107,In_290,In_537);
nor U108 (N_108,In_1267,In_789);
or U109 (N_109,In_1478,In_819);
xnor U110 (N_110,In_921,In_54);
nand U111 (N_111,In_624,In_601);
nor U112 (N_112,In_835,In_1118);
nor U113 (N_113,In_1323,In_1114);
or U114 (N_114,In_1102,In_709);
and U115 (N_115,In_1205,In_43);
nand U116 (N_116,In_989,In_733);
nand U117 (N_117,In_727,In_45);
and U118 (N_118,In_636,In_1181);
or U119 (N_119,In_458,In_646);
nor U120 (N_120,In_121,In_648);
nand U121 (N_121,In_1344,In_1449);
or U122 (N_122,In_1204,In_698);
nor U123 (N_123,In_1094,In_656);
nor U124 (N_124,In_979,In_348);
nand U125 (N_125,In_486,In_1281);
nor U126 (N_126,In_429,In_89);
xor U127 (N_127,In_655,In_695);
nor U128 (N_128,In_1195,In_405);
and U129 (N_129,In_754,In_903);
or U130 (N_130,In_227,In_477);
or U131 (N_131,In_109,In_1156);
nand U132 (N_132,In_734,In_829);
or U133 (N_133,In_1041,In_93);
nor U134 (N_134,In_706,In_561);
nor U135 (N_135,In_475,In_208);
xor U136 (N_136,In_48,In_1333);
nand U137 (N_137,In_1006,In_201);
nand U138 (N_138,In_1079,In_1122);
xor U139 (N_139,In_44,In_740);
nor U140 (N_140,In_557,In_520);
or U141 (N_141,In_649,In_125);
xor U142 (N_142,In_696,In_1424);
nand U143 (N_143,In_1342,In_1021);
nor U144 (N_144,In_997,In_422);
xor U145 (N_145,In_284,In_1228);
nand U146 (N_146,In_20,In_961);
nor U147 (N_147,In_29,In_364);
and U148 (N_148,In_32,In_7);
and U149 (N_149,In_46,In_209);
or U150 (N_150,In_5,In_1431);
nor U151 (N_151,In_183,In_896);
nand U152 (N_152,In_331,In_971);
nor U153 (N_153,In_230,In_34);
nor U154 (N_154,In_1341,In_1283);
and U155 (N_155,In_23,In_1479);
nor U156 (N_156,In_1254,In_155);
xor U157 (N_157,In_319,In_1028);
nor U158 (N_158,In_210,In_1091);
xor U159 (N_159,In_1140,In_363);
nand U160 (N_160,In_1326,In_504);
and U161 (N_161,In_1291,In_1023);
nor U162 (N_162,In_1409,In_941);
xnor U163 (N_163,In_1264,In_1470);
nor U164 (N_164,In_1246,In_219);
nand U165 (N_165,In_562,In_943);
and U166 (N_166,In_463,In_280);
and U167 (N_167,In_568,In_1000);
nand U168 (N_168,In_759,In_428);
or U169 (N_169,In_1165,In_318);
nand U170 (N_170,In_633,In_776);
nand U171 (N_171,In_723,In_737);
nand U172 (N_172,In_1381,In_168);
or U173 (N_173,In_772,In_116);
nor U174 (N_174,In_1483,In_15);
and U175 (N_175,In_1328,In_973);
or U176 (N_176,In_1416,In_1367);
nand U177 (N_177,In_1024,In_1033);
or U178 (N_178,In_1365,In_170);
nand U179 (N_179,In_1230,In_811);
nand U180 (N_180,In_485,In_642);
or U181 (N_181,In_1271,In_1293);
nand U182 (N_182,In_410,In_1497);
and U183 (N_183,In_758,In_132);
nor U184 (N_184,In_293,In_1314);
xor U185 (N_185,In_798,In_272);
nand U186 (N_186,In_1274,In_115);
nand U187 (N_187,In_784,In_1109);
and U188 (N_188,In_204,In_1151);
or U189 (N_189,In_390,In_512);
nor U190 (N_190,In_1180,In_749);
and U191 (N_191,In_1417,In_1234);
and U192 (N_192,In_175,In_999);
or U193 (N_193,In_53,In_814);
nor U194 (N_194,In_304,In_1422);
nor U195 (N_195,In_1112,In_1393);
or U196 (N_196,In_3,In_498);
nand U197 (N_197,In_1414,In_892);
xor U198 (N_198,In_355,In_484);
or U199 (N_199,In_263,In_1121);
nand U200 (N_200,In_791,In_213);
nand U201 (N_201,In_757,In_1038);
or U202 (N_202,In_321,In_445);
xnor U203 (N_203,In_1395,In_1372);
or U204 (N_204,In_37,In_1298);
nand U205 (N_205,In_703,In_327);
nand U206 (N_206,In_761,In_305);
and U207 (N_207,In_799,In_345);
nand U208 (N_208,In_266,In_1468);
nor U209 (N_209,In_932,In_285);
xnor U210 (N_210,In_42,In_548);
or U211 (N_211,In_1051,In_1073);
xnor U212 (N_212,In_877,In_1498);
and U213 (N_213,In_206,In_1012);
or U214 (N_214,In_1437,In_968);
nand U215 (N_215,In_380,In_105);
and U216 (N_216,In_567,In_854);
and U217 (N_217,In_984,In_1441);
xnor U218 (N_218,In_1359,In_744);
nand U219 (N_219,In_1169,In_953);
xor U220 (N_220,In_420,In_1116);
and U221 (N_221,In_1225,In_1436);
and U222 (N_222,In_827,In_1215);
nor U223 (N_223,In_1087,In_57);
nor U224 (N_224,In_1402,In_797);
nor U225 (N_225,In_507,In_1320);
nor U226 (N_226,In_1315,In_1340);
and U227 (N_227,In_625,In_450);
xor U228 (N_228,In_1131,In_430);
nor U229 (N_229,In_1316,In_676);
nand U230 (N_230,In_1226,In_1211);
nand U231 (N_231,In_1307,In_464);
and U232 (N_232,In_368,In_782);
and U233 (N_233,In_637,In_947);
nand U234 (N_234,In_78,In_479);
and U235 (N_235,In_1335,In_1212);
nor U236 (N_236,In_1311,In_497);
nor U237 (N_237,In_914,In_608);
or U238 (N_238,In_556,In_359);
nand U239 (N_239,In_1308,In_212);
nand U240 (N_240,In_666,In_1456);
xor U241 (N_241,In_436,In_593);
or U242 (N_242,In_902,In_735);
xnor U243 (N_243,In_169,In_553);
nor U244 (N_244,In_1086,In_1282);
or U245 (N_245,In_818,In_848);
or U246 (N_246,In_22,In_780);
xnor U247 (N_247,In_1113,In_645);
or U248 (N_248,In_1257,In_1238);
xnor U249 (N_249,In_1389,In_111);
and U250 (N_250,In_613,In_1039);
nor U251 (N_251,In_391,In_374);
or U252 (N_252,In_320,In_785);
xor U253 (N_253,In_1174,N_111);
nor U254 (N_254,In_518,In_741);
and U255 (N_255,In_1480,In_612);
nor U256 (N_256,In_1440,In_875);
and U257 (N_257,N_29,N_86);
or U258 (N_258,In_867,In_635);
nor U259 (N_259,In_1018,In_133);
nand U260 (N_260,In_1373,N_170);
nand U261 (N_261,In_969,In_707);
or U262 (N_262,N_167,N_183);
nor U263 (N_263,In_64,In_630);
and U264 (N_264,In_461,In_1142);
nand U265 (N_265,In_404,In_1419);
and U266 (N_266,In_180,N_32);
xnor U267 (N_267,In_1430,N_133);
or U268 (N_268,In_1198,In_135);
xor U269 (N_269,In_1462,In_623);
and U270 (N_270,N_7,In_198);
nand U271 (N_271,In_738,N_48);
and U272 (N_272,N_168,In_226);
nand U273 (N_273,In_853,In_432);
and U274 (N_274,N_10,In_844);
nand U275 (N_275,N_22,In_926);
nand U276 (N_276,In_1454,In_535);
nor U277 (N_277,In_851,In_369);
xor U278 (N_278,In_673,In_274);
xnor U279 (N_279,In_1015,N_40);
and U280 (N_280,In_1432,N_56);
and U281 (N_281,In_438,In_1294);
or U282 (N_282,In_211,In_675);
nand U283 (N_283,In_1412,In_249);
xnor U284 (N_284,In_153,In_1136);
xnor U285 (N_285,In_1425,In_378);
or U286 (N_286,In_591,N_128);
nand U287 (N_287,In_869,In_1413);
nand U288 (N_288,In_187,In_887);
nor U289 (N_289,In_40,In_86);
and U290 (N_290,N_247,In_995);
nand U291 (N_291,N_245,N_117);
xor U292 (N_292,In_1193,In_61);
xnor U293 (N_293,In_585,In_1089);
nor U294 (N_294,In_752,In_238);
or U295 (N_295,In_56,In_581);
or U296 (N_296,In_254,In_747);
or U297 (N_297,N_220,In_1460);
and U298 (N_298,In_384,N_33);
nand U299 (N_299,In_725,In_102);
xor U300 (N_300,In_500,N_190);
or U301 (N_301,N_166,In_1096);
nand U302 (N_302,In_273,In_936);
xnor U303 (N_303,In_330,In_513);
nor U304 (N_304,In_1491,In_1097);
or U305 (N_305,In_1471,N_36);
xnor U306 (N_306,In_1494,In_1442);
nand U307 (N_307,In_607,In_1161);
or U308 (N_308,In_909,In_672);
nor U309 (N_309,In_988,In_403);
or U310 (N_310,In_840,N_218);
nand U311 (N_311,In_1054,In_1034);
and U312 (N_312,In_298,In_924);
or U313 (N_313,N_171,In_523);
nand U314 (N_314,In_710,N_211);
and U315 (N_315,In_367,In_481);
or U316 (N_316,In_868,In_70);
xnor U317 (N_317,N_107,In_312);
or U318 (N_318,In_543,In_774);
xnor U319 (N_319,In_241,In_722);
nor U320 (N_320,In_262,In_1477);
nand U321 (N_321,In_717,N_24);
or U322 (N_322,In_229,In_662);
and U323 (N_323,In_1376,In_842);
nor U324 (N_324,N_77,In_1217);
and U325 (N_325,In_1160,N_85);
nor U326 (N_326,In_1146,In_1266);
nand U327 (N_327,In_1380,In_1166);
and U328 (N_328,In_582,In_455);
xnor U329 (N_329,In_944,In_1233);
nand U330 (N_330,In_503,In_889);
and U331 (N_331,In_394,In_641);
xnor U332 (N_332,In_713,In_1105);
xnor U333 (N_333,In_1493,In_408);
xnor U334 (N_334,N_246,In_843);
and U335 (N_335,In_460,In_18);
nand U336 (N_336,In_962,In_289);
nor U337 (N_337,N_201,In_775);
or U338 (N_338,In_506,In_1231);
nor U339 (N_339,In_898,In_192);
or U340 (N_340,In_1304,In_1249);
nand U341 (N_341,In_147,N_199);
xnor U342 (N_342,In_277,N_169);
xnor U343 (N_343,In_1148,In_1187);
xnor U344 (N_344,In_1026,In_239);
nand U345 (N_345,N_228,In_1078);
and U346 (N_346,In_669,In_559);
xnor U347 (N_347,In_639,In_265);
and U348 (N_348,In_546,In_76);
xnor U349 (N_349,In_1275,In_1329);
nor U350 (N_350,In_963,In_176);
nor U351 (N_351,In_833,In_161);
xnor U352 (N_352,N_155,In_704);
nor U353 (N_353,In_1481,N_102);
xnor U354 (N_354,In_301,In_496);
xor U355 (N_355,N_187,In_715);
and U356 (N_356,In_522,In_1125);
xor U357 (N_357,In_317,In_532);
nand U358 (N_358,In_282,N_126);
nor U359 (N_359,In_1115,In_604);
nor U360 (N_360,N_226,N_206);
nand U361 (N_361,In_323,In_970);
or U362 (N_362,In_587,In_1189);
nand U363 (N_363,N_221,In_1072);
nand U364 (N_364,In_488,In_787);
nand U365 (N_365,N_197,N_83);
or U366 (N_366,In_720,In_688);
nor U367 (N_367,N_21,In_200);
or U368 (N_368,In_982,In_361);
or U369 (N_369,N_136,In_751);
and U370 (N_370,In_769,In_167);
nand U371 (N_371,In_1490,N_146);
xnor U372 (N_372,In_409,In_1168);
or U373 (N_373,In_540,In_830);
nor U374 (N_374,In_1209,In_346);
xor U375 (N_375,N_160,N_159);
xnor U376 (N_376,In_765,In_805);
and U377 (N_377,In_193,In_939);
and U378 (N_378,In_945,In_1066);
and U379 (N_379,In_237,In_1227);
and U380 (N_380,In_925,In_297);
and U381 (N_381,In_1050,In_156);
nand U382 (N_382,N_113,In_1172);
nor U383 (N_383,N_79,In_426);
and U384 (N_384,N_89,N_9);
nor U385 (N_385,In_580,In_157);
and U386 (N_386,N_200,N_2);
nor U387 (N_387,In_474,In_516);
or U388 (N_388,In_60,In_628);
nor U389 (N_389,In_647,N_178);
nand U390 (N_390,In_1330,In_184);
or U391 (N_391,In_991,N_11);
and U392 (N_392,In_1473,In_1263);
xor U393 (N_393,In_1076,In_605);
and U394 (N_394,In_1345,In_421);
xor U395 (N_395,In_140,In_275);
nand U396 (N_396,In_90,In_478);
and U397 (N_397,N_238,In_1452);
nand U398 (N_398,In_732,In_721);
and U399 (N_399,N_176,In_214);
xor U400 (N_400,N_204,In_951);
and U401 (N_401,In_1185,N_34);
and U402 (N_402,In_822,N_38);
or U403 (N_403,In_389,In_729);
xnor U404 (N_404,In_948,In_1104);
xor U405 (N_405,In_80,In_356);
nand U406 (N_406,In_1453,N_99);
and U407 (N_407,In_1057,N_17);
nor U408 (N_408,In_956,In_1154);
and U409 (N_409,In_382,N_164);
and U410 (N_410,In_228,In_542);
or U411 (N_411,In_1232,In_472);
or U412 (N_412,In_1020,In_41);
and U413 (N_413,In_793,In_82);
xor U414 (N_414,In_849,N_149);
nand U415 (N_415,In_55,In_1260);
and U416 (N_416,In_113,In_992);
nand U417 (N_417,In_103,N_0);
or U418 (N_418,In_651,In_788);
nand U419 (N_419,N_196,In_417);
nand U420 (N_420,In_1070,N_154);
or U421 (N_421,In_1110,N_91);
or U422 (N_422,In_1196,In_313);
nor U423 (N_423,In_38,In_841);
xor U424 (N_424,In_1270,In_1310);
nor U425 (N_425,In_12,In_719);
nor U426 (N_426,In_234,In_544);
xnor U427 (N_427,In_1400,In_912);
nor U428 (N_428,In_726,In_1240);
nand U429 (N_429,In_653,In_859);
or U430 (N_430,In_1446,In_177);
and U431 (N_431,In_654,N_28);
nor U432 (N_432,In_1220,In_1391);
or U433 (N_433,In_1461,In_777);
or U434 (N_434,In_1450,N_202);
nor U435 (N_435,N_181,In_831);
nor U436 (N_436,N_60,In_1124);
and U437 (N_437,In_126,In_260);
nor U438 (N_438,N_207,In_1243);
xnor U439 (N_439,In_8,In_705);
nor U440 (N_440,In_162,In_97);
xor U441 (N_441,In_803,In_129);
or U442 (N_442,N_119,In_617);
xnor U443 (N_443,N_90,In_1455);
and U444 (N_444,In_95,In_884);
nand U445 (N_445,In_745,In_1016);
or U446 (N_446,N_231,In_407);
or U447 (N_447,In_337,In_1222);
nand U448 (N_448,In_1139,In_267);
or U449 (N_449,N_39,In_1037);
nand U450 (N_450,N_135,In_258);
or U451 (N_451,In_687,N_25);
xor U452 (N_452,N_4,In_1141);
nand U453 (N_453,N_223,In_1201);
or U454 (N_454,In_91,In_660);
xor U455 (N_455,In_1123,N_131);
nand U456 (N_456,In_159,In_610);
or U457 (N_457,In_85,In_652);
or U458 (N_458,N_18,N_87);
nor U459 (N_459,In_558,In_163);
nand U460 (N_460,In_966,In_491);
xnor U461 (N_461,In_570,In_470);
nor U462 (N_462,In_857,N_57);
nand U463 (N_463,In_1022,In_413);
and U464 (N_464,In_1464,N_139);
and U465 (N_465,In_1013,N_212);
xnor U466 (N_466,In_766,In_906);
nor U467 (N_467,In_1467,In_813);
xor U468 (N_468,In_756,In_684);
nand U469 (N_469,N_180,In_960);
or U470 (N_470,In_586,In_310);
nor U471 (N_471,In_67,In_731);
nor U472 (N_472,N_97,In_1153);
or U473 (N_473,In_1130,In_124);
or U474 (N_474,In_919,In_1265);
and U475 (N_475,In_1063,In_216);
nand U476 (N_476,In_680,In_81);
or U477 (N_477,In_957,In_94);
nand U478 (N_478,In_911,In_1010);
or U479 (N_479,N_140,N_45);
nor U480 (N_480,In_328,In_1258);
or U481 (N_481,In_1245,N_142);
and U482 (N_482,In_781,In_755);
nand U483 (N_483,In_288,In_100);
nor U484 (N_484,In_202,In_517);
nor U485 (N_485,In_530,In_1299);
and U486 (N_486,In_629,In_1071);
nor U487 (N_487,In_1150,In_708);
nand U488 (N_488,In_307,In_58);
nor U489 (N_489,In_1476,In_1351);
and U490 (N_490,In_644,N_125);
nor U491 (N_491,N_5,In_1241);
nor U492 (N_492,In_1178,In_247);
or U493 (N_493,In_188,N_69);
nand U494 (N_494,In_1058,In_907);
nand U495 (N_495,In_231,In_671);
xor U496 (N_496,In_1170,In_1223);
or U497 (N_497,In_145,In_839);
nand U498 (N_498,In_937,In_560);
or U499 (N_499,N_239,In_270);
or U500 (N_500,N_301,N_255);
or U501 (N_501,N_334,N_391);
nand U502 (N_502,N_279,In_379);
or U503 (N_503,N_478,In_339);
and U504 (N_504,In_467,In_712);
nor U505 (N_505,N_104,N_233);
or U506 (N_506,N_489,N_344);
and U507 (N_507,N_59,N_241);
and U508 (N_508,N_303,N_364);
nor U509 (N_509,In_411,N_324);
and U510 (N_510,In_763,In_386);
or U511 (N_511,N_161,In_1075);
nand U512 (N_512,N_323,N_100);
nor U513 (N_513,In_120,In_511);
and U514 (N_514,In_283,In_333);
nand U515 (N_515,N_82,N_253);
xor U516 (N_516,In_935,N_397);
nand U517 (N_517,N_384,In_490);
xor U518 (N_518,N_358,In_812);
xnor U519 (N_519,N_35,N_390);
xnor U520 (N_520,N_298,In_396);
nand U521 (N_521,In_1027,N_402);
or U522 (N_522,In_31,N_274);
or U523 (N_523,In_495,In_897);
and U524 (N_524,In_160,N_428);
nand U525 (N_525,In_1218,In_565);
and U526 (N_526,In_502,In_1305);
nor U527 (N_527,N_349,N_115);
and U528 (N_528,In_309,In_1302);
nand U529 (N_529,N_430,N_216);
xor U530 (N_530,In_977,In_84);
xnor U531 (N_531,N_265,In_908);
or U532 (N_532,In_358,N_123);
nand U533 (N_533,In_1363,In_406);
xor U534 (N_534,In_815,N_389);
nor U535 (N_535,In_1295,In_1420);
nor U536 (N_536,N_361,In_697);
xor U537 (N_537,N_251,In_1008);
nand U538 (N_538,In_372,N_152);
xnor U539 (N_539,In_392,In_594);
nor U540 (N_540,N_424,In_916);
xnor U541 (N_541,In_1434,In_207);
nand U542 (N_542,In_596,In_527);
and U543 (N_543,In_683,N_73);
nor U544 (N_544,In_1065,In_1);
nor U545 (N_545,N_385,N_452);
or U546 (N_546,In_1134,In_800);
nand U547 (N_547,In_377,N_337);
or U548 (N_548,In_395,N_352);
nand U549 (N_549,In_469,In_281);
nand U550 (N_550,N_134,In_243);
and U551 (N_551,N_434,In_934);
and U552 (N_552,In_179,In_1366);
nand U553 (N_553,N_203,N_145);
nand U554 (N_554,In_107,N_493);
xnor U555 (N_555,In_668,In_905);
nor U556 (N_556,N_431,In_885);
or U557 (N_557,N_208,In_1117);
nand U558 (N_558,N_8,N_497);
nand U559 (N_559,In_980,In_98);
or U560 (N_560,In_615,N_43);
xor U561 (N_561,N_116,N_436);
or U562 (N_562,In_1346,In_1297);
xor U563 (N_563,N_230,N_213);
or U564 (N_564,N_355,In_203);
nand U565 (N_565,In_978,N_401);
and U566 (N_566,N_98,In_362);
xnor U567 (N_567,N_420,In_1404);
or U568 (N_568,In_790,In_1489);
nand U569 (N_569,N_275,In_1188);
xor U570 (N_570,In_1210,N_264);
xnor U571 (N_571,In_118,In_534);
or U572 (N_572,N_414,N_396);
nand U573 (N_573,In_171,In_1192);
or U574 (N_574,In_149,In_1152);
xor U575 (N_575,N_468,N_318);
nor U576 (N_576,N_289,In_1327);
or U577 (N_577,In_701,N_367);
nand U578 (N_578,In_452,In_248);
and U579 (N_579,In_950,In_311);
or U580 (N_580,In_88,In_1447);
and U581 (N_581,In_638,N_103);
nor U582 (N_582,In_1338,In_519);
nand U583 (N_583,In_714,N_37);
nand U584 (N_584,In_860,In_1374);
or U585 (N_585,In_106,In_794);
nor U586 (N_586,In_1401,In_870);
and U587 (N_587,In_1358,In_821);
and U588 (N_588,N_466,N_165);
nor U589 (N_589,In_965,In_236);
xnor U590 (N_590,N_331,In_1405);
xnor U591 (N_591,In_286,In_108);
and U592 (N_592,N_269,In_1031);
xnor U593 (N_593,In_468,In_1044);
or U594 (N_594,N_365,In_489);
or U595 (N_595,In_1496,N_44);
nand U596 (N_596,In_1361,In_554);
xor U597 (N_597,N_380,In_692);
and U598 (N_598,In_1045,In_878);
nand U599 (N_599,In_189,N_471);
and U600 (N_600,N_339,In_174);
xnor U601 (N_601,N_437,In_1487);
or U602 (N_602,In_716,In_1036);
and U603 (N_603,In_342,In_259);
nor U604 (N_604,In_205,N_217);
nand U605 (N_605,In_972,In_1255);
nor U606 (N_606,In_1093,N_137);
or U607 (N_607,In_449,In_1060);
and U608 (N_608,In_810,N_378);
nand U609 (N_609,N_382,In_1287);
and U610 (N_610,N_476,N_374);
xnor U611 (N_611,In_1173,N_74);
or U612 (N_612,N_320,N_329);
xnor U613 (N_613,N_129,N_42);
nor U614 (N_614,In_1397,In_958);
nor U615 (N_615,N_295,In_1336);
and U616 (N_616,N_54,N_225);
and U617 (N_617,In_110,In_746);
nor U618 (N_618,N_81,In_1332);
and U619 (N_619,In_499,N_381);
or U620 (N_620,In_1088,N_242);
nor U621 (N_621,N_398,N_456);
or U622 (N_622,In_50,In_1224);
and U623 (N_623,In_451,In_47);
or U624 (N_624,In_1176,In_1356);
and U625 (N_625,N_496,In_268);
xnor U626 (N_626,In_650,N_156);
nor U627 (N_627,N_294,N_438);
nor U628 (N_628,N_432,In_1384);
nor U629 (N_629,In_416,In_1048);
nor U630 (N_630,In_1025,N_499);
nor U631 (N_631,In_1061,In_563);
or U632 (N_632,In_235,In_412);
nor U633 (N_633,In_1443,N_464);
xnor U634 (N_634,In_264,In_938);
and U635 (N_635,In_439,In_809);
and U636 (N_636,In_295,In_255);
and U637 (N_637,In_1360,N_427);
nand U638 (N_638,In_724,N_30);
nor U639 (N_639,In_462,In_873);
nor U640 (N_640,N_3,N_342);
nor U641 (N_641,N_271,In_1284);
or U642 (N_642,N_198,In_894);
nand U643 (N_643,N_457,N_421);
nor U644 (N_644,In_278,In_233);
and U645 (N_645,In_1175,N_327);
or U646 (N_646,In_1126,In_664);
nand U647 (N_647,In_131,N_153);
or U648 (N_648,In_825,In_473);
xor U649 (N_649,N_23,In_341);
nand U650 (N_650,N_407,In_1120);
nand U651 (N_651,In_299,In_292);
nand U652 (N_652,N_95,N_447);
or U653 (N_653,In_322,N_388);
or U654 (N_654,In_1159,N_188);
and U655 (N_655,In_1382,N_16);
nor U656 (N_656,In_711,N_399);
or U657 (N_657,In_10,In_1312);
or U658 (N_658,In_584,In_2);
and U659 (N_659,N_338,In_1216);
and U660 (N_660,N_244,In_659);
or U661 (N_661,In_388,N_141);
xnor U662 (N_662,N_173,In_1427);
xor U663 (N_663,N_259,N_78);
or U664 (N_664,In_164,In_773);
xnor U665 (N_665,N_297,In_257);
nand U666 (N_666,In_626,In_515);
nand U667 (N_667,In_138,In_508);
or U668 (N_668,In_1247,N_191);
or U669 (N_669,N_106,N_405);
or U670 (N_670,In_483,N_240);
or U671 (N_671,In_1457,In_609);
xnor U672 (N_672,N_483,In_691);
nor U673 (N_673,N_234,N_118);
nand U674 (N_674,In_435,N_75);
xor U675 (N_675,N_27,In_75);
nor U676 (N_676,In_1438,In_529);
nand U677 (N_677,In_253,In_393);
or U678 (N_678,N_280,N_88);
nor U679 (N_679,In_678,In_215);
and U680 (N_680,In_1221,In_893);
nor U681 (N_681,N_371,In_1030);
or U682 (N_682,N_314,In_1495);
nor U683 (N_683,In_1135,In_1177);
or U684 (N_684,In_913,N_120);
or U685 (N_685,N_312,In_340);
nor U686 (N_686,N_495,In_879);
or U687 (N_687,In_1171,N_132);
xor U688 (N_688,In_996,N_292);
nand U689 (N_689,In_1014,In_300);
or U690 (N_690,In_308,In_764);
and U691 (N_691,N_450,N_469);
and U692 (N_692,In_915,N_209);
and U693 (N_693,N_127,In_296);
xor U694 (N_694,N_400,In_1410);
nor U695 (N_695,N_317,In_250);
or U696 (N_696,In_657,N_144);
or U697 (N_697,N_55,N_412);
and U698 (N_698,In_35,N_326);
nor U699 (N_699,In_927,In_882);
and U700 (N_700,In_1331,N_488);
xnor U701 (N_701,N_467,In_658);
and U702 (N_702,In_27,In_256);
nand U703 (N_703,N_237,N_316);
or U704 (N_704,In_148,In_1388);
and U705 (N_705,In_750,N_76);
nand U706 (N_706,N_235,In_1278);
or U707 (N_707,N_287,In_1357);
and U708 (N_708,N_157,In_326);
and U709 (N_709,In_1261,N_386);
xor U710 (N_710,In_1317,N_440);
nand U711 (N_711,N_49,In_861);
and U712 (N_712,In_574,In_1236);
nor U713 (N_713,N_366,In_245);
xnor U714 (N_714,In_419,In_1390);
xor U715 (N_715,N_473,N_392);
xor U716 (N_716,In_588,In_795);
and U717 (N_717,N_138,In_771);
xnor U718 (N_718,In_975,N_480);
and U719 (N_719,In_1347,In_1029);
nor U720 (N_720,In_1469,In_252);
nor U721 (N_721,In_592,In_324);
nor U722 (N_722,N_321,N_177);
nand U723 (N_723,In_670,In_862);
xor U724 (N_724,N_299,N_50);
nand U725 (N_725,N_272,N_257);
nor U726 (N_726,In_1418,N_330);
nand U727 (N_727,In_101,In_13);
and U728 (N_728,In_1368,In_1486);
xor U729 (N_729,N_350,N_266);
or U730 (N_730,In_920,In_627);
or U731 (N_731,N_347,In_501);
xnor U732 (N_732,In_566,In_863);
nand U733 (N_733,In_689,In_792);
nor U734 (N_734,N_340,N_461);
and U735 (N_735,N_193,In_1145);
nand U736 (N_736,N_311,N_232);
nand U737 (N_737,In_1084,In_123);
xor U738 (N_738,In_663,N_41);
or U739 (N_739,In_397,In_864);
nor U740 (N_740,In_1162,N_319);
xnor U741 (N_741,In_1459,N_328);
and U742 (N_742,N_112,N_494);
or U743 (N_743,N_395,In_804);
or U744 (N_744,In_536,N_243);
nand U745 (N_745,In_21,In_1343);
nor U746 (N_746,N_387,N_403);
nor U747 (N_747,In_444,In_465);
nor U748 (N_748,In_232,In_1035);
nand U749 (N_749,In_1229,In_917);
and U750 (N_750,N_179,N_276);
nand U751 (N_751,N_612,In_196);
nor U752 (N_752,N_410,In_134);
nor U753 (N_753,N_446,N_519);
nand U754 (N_754,In_779,N_250);
xor U755 (N_755,In_910,In_454);
nor U756 (N_756,N_746,In_431);
or U757 (N_757,In_117,N_459);
nor U758 (N_758,N_31,In_335);
or U759 (N_759,N_570,N_394);
or U760 (N_760,N_543,N_554);
nand U761 (N_761,N_727,N_610);
xor U762 (N_762,N_463,In_1444);
or U763 (N_763,In_876,In_739);
xor U764 (N_764,N_93,N_707);
and U765 (N_765,N_418,N_582);
xnor U766 (N_766,In_49,In_1248);
nand U767 (N_767,N_693,N_256);
or U768 (N_768,In_433,In_399);
and U769 (N_769,In_68,N_625);
or U770 (N_770,In_1158,N_510);
nor U771 (N_771,In_1046,In_74);
nor U772 (N_772,N_46,N_718);
nor U773 (N_773,In_1040,N_65);
xnor U774 (N_774,N_692,In_294);
nand U775 (N_775,N_372,N_677);
nand U776 (N_776,In_291,N_647);
and U777 (N_777,In_904,In_1433);
xor U778 (N_778,N_583,In_1167);
xnor U779 (N_779,N_511,N_520);
or U780 (N_780,N_296,N_66);
or U781 (N_781,N_720,In_185);
nor U782 (N_782,In_1203,N_531);
nand U783 (N_783,N_278,N_182);
nand U784 (N_784,In_1288,N_565);
xnor U785 (N_785,N_268,N_571);
nor U786 (N_786,In_402,N_479);
nor U787 (N_787,N_533,In_1092);
or U788 (N_788,N_705,N_62);
xor U789 (N_789,N_624,N_96);
and U790 (N_790,N_703,N_581);
nor U791 (N_791,In_952,In_418);
and U792 (N_792,N_194,In_888);
and U793 (N_793,N_490,In_9);
or U794 (N_794,N_724,In_824);
xnor U795 (N_795,N_662,In_871);
or U796 (N_796,In_578,N_283);
xor U797 (N_797,In_865,N_538);
nand U798 (N_798,In_886,In_1439);
nor U799 (N_799,N_393,N_375);
nand U800 (N_800,In_575,In_1465);
and U801 (N_801,N_84,In_306);
xor U802 (N_802,N_47,N_563);
nor U803 (N_803,N_557,In_11);
xor U804 (N_804,In_1362,N_512);
nor U805 (N_805,In_550,N_649);
or U806 (N_806,N_290,In_139);
nor U807 (N_807,N_738,N_20);
or U808 (N_808,N_492,In_1059);
xnor U809 (N_809,N_453,In_949);
xnor U810 (N_810,In_1213,N_648);
nand U811 (N_811,In_690,N_732);
and U812 (N_812,In_1303,N_186);
xor U813 (N_813,In_398,N_733);
and U814 (N_814,In_564,N_712);
nor U815 (N_815,N_518,In_401);
nand U816 (N_816,In_539,In_353);
xnor U817 (N_817,In_1090,In_1319);
or U818 (N_818,In_1064,In_933);
nand U819 (N_819,N_689,In_1269);
nor U820 (N_820,In_880,In_606);
or U821 (N_821,N_475,In_1202);
xor U822 (N_822,N_195,N_150);
xor U823 (N_823,N_719,N_659);
or U824 (N_824,N_723,N_377);
nor U825 (N_825,In_261,N_6);
or U826 (N_826,N_660,N_481);
xnor U827 (N_827,In_748,N_151);
or U828 (N_828,In_375,In_579);
and U829 (N_829,N_504,In_850);
xnor U830 (N_830,N_376,In_25);
or U831 (N_831,N_672,In_1289);
or U832 (N_832,In_400,In_928);
nand U833 (N_833,In_1268,N_686);
nor U834 (N_834,N_335,N_449);
or U835 (N_835,N_460,N_508);
nor U836 (N_836,N_262,In_347);
or U837 (N_837,In_832,In_768);
nand U838 (N_838,In_494,N_621);
or U839 (N_839,In_385,N_522);
or U840 (N_840,In_1144,N_650);
and U841 (N_841,In_808,In_1403);
and U842 (N_842,In_806,N_729);
nand U843 (N_843,In_802,N_501);
nor U844 (N_844,N_706,N_286);
xor U845 (N_845,N_516,N_559);
nand U846 (N_846,In_271,In_1250);
nand U847 (N_847,N_51,N_163);
nor U848 (N_848,N_584,In_890);
xor U849 (N_849,N_332,In_583);
nand U850 (N_850,In_441,N_210);
xnor U851 (N_851,In_276,N_71);
or U852 (N_852,N_529,N_606);
and U853 (N_853,N_362,N_683);
xor U854 (N_854,N_644,N_657);
nand U855 (N_855,In_531,In_1428);
or U856 (N_856,In_51,N_61);
xor U857 (N_857,In_447,In_1108);
or U858 (N_858,N_640,N_484);
nand U859 (N_859,N_575,N_740);
nand U860 (N_860,N_19,In_83);
xnor U861 (N_861,N_185,In_366);
xor U862 (N_862,In_119,N_354);
nand U863 (N_863,In_104,N_451);
and U864 (N_864,In_891,In_918);
xor U865 (N_865,N_711,N_348);
xnor U866 (N_866,N_58,N_696);
xnor U867 (N_867,N_260,N_307);
xor U868 (N_868,In_1406,N_470);
xor U869 (N_869,In_823,N_551);
or U870 (N_870,In_344,In_1292);
or U871 (N_871,In_220,N_564);
nor U872 (N_872,In_643,N_637);
and U873 (N_873,In_1183,In_251);
or U874 (N_874,In_1448,N_679);
nor U875 (N_875,In_1164,In_1280);
xnor U876 (N_876,In_1277,N_617);
or U877 (N_877,N_602,In_1415);
xor U878 (N_878,N_555,N_285);
and U879 (N_879,N_748,N_454);
xor U880 (N_880,In_1276,N_726);
nand U881 (N_881,N_631,N_669);
nand U882 (N_882,N_687,In_144);
xnor U883 (N_883,N_448,N_80);
or U884 (N_884,In_434,N_304);
xor U885 (N_885,N_506,N_485);
nand U886 (N_886,In_350,In_387);
or U887 (N_887,In_828,N_735);
and U888 (N_888,N_676,In_1062);
or U889 (N_889,N_404,In_600);
and U890 (N_890,In_846,N_576);
or U891 (N_891,N_668,In_217);
and U892 (N_892,N_442,In_218);
or U893 (N_893,N_562,N_714);
and U894 (N_894,In_901,N_205);
or U895 (N_895,In_453,N_544);
or U896 (N_896,N_629,In_895);
xor U897 (N_897,N_725,N_63);
nor U898 (N_898,N_505,N_64);
nor U899 (N_899,In_525,N_313);
nand U900 (N_900,In_1290,In_1398);
nor U901 (N_901,In_151,N_513);
xnor U902 (N_902,In_801,In_533);
or U903 (N_903,N_553,In_1082);
xor U904 (N_904,In_1348,N_148);
or U905 (N_905,In_545,N_567);
xnor U906 (N_906,N_472,N_569);
or U907 (N_907,N_507,In_1407);
xnor U908 (N_908,In_1194,In_325);
xnor U909 (N_909,In_1003,N_666);
nor U910 (N_910,In_942,In_1352);
nor U911 (N_911,N_675,In_1354);
and U912 (N_912,In_154,N_67);
and U913 (N_913,N_709,N_353);
nand U914 (N_914,N_270,In_1184);
xor U915 (N_915,In_661,N_370);
nor U916 (N_916,N_585,N_639);
or U917 (N_917,In_19,N_68);
nand U918 (N_918,In_736,N_310);
nor U919 (N_919,In_79,N_745);
or U920 (N_920,In_1383,N_739);
or U921 (N_921,N_13,N_598);
nor U922 (N_922,In_858,In_354);
and U923 (N_923,N_411,In_603);
nand U924 (N_924,N_577,N_517);
or U925 (N_925,N_425,In_371);
xor U926 (N_926,N_114,N_592);
nor U927 (N_927,In_1219,N_474);
or U928 (N_928,In_197,In_837);
nor U929 (N_929,N_593,In_1313);
or U930 (N_930,In_1350,In_1349);
and U931 (N_931,N_130,In_983);
xnor U932 (N_932,N_281,N_590);
or U933 (N_933,N_343,N_458);
nor U934 (N_934,N_737,N_604);
nor U935 (N_935,N_635,N_101);
xor U936 (N_936,In_1239,N_122);
and U937 (N_937,In_1149,In_541);
nand U938 (N_938,In_551,N_716);
nor U939 (N_939,In_352,N_525);
nor U940 (N_940,N_14,In_1324);
nand U941 (N_941,N_700,In_872);
or U942 (N_942,N_704,N_652);
nand U943 (N_943,N_678,N_445);
nand U944 (N_944,N_282,In_26);
and U945 (N_945,In_17,N_741);
or U946 (N_946,In_150,In_199);
and U947 (N_947,N_702,In_1081);
and U948 (N_948,N_124,N_305);
nor U949 (N_949,N_736,N_552);
nor U950 (N_950,N_110,N_655);
xnor U951 (N_951,In_52,N_174);
and U952 (N_952,N_53,N_742);
or U953 (N_953,In_1485,N_379);
nor U954 (N_954,In_834,N_614);
nor U955 (N_955,In_1322,In_640);
and U956 (N_956,N_651,In_87);
nor U957 (N_957,In_820,N_607);
or U958 (N_958,N_708,N_667);
or U959 (N_959,N_540,In_66);
nand U960 (N_960,N_263,In_521);
and U961 (N_961,N_561,N_597);
xor U962 (N_962,N_308,N_599);
nand U963 (N_963,N_26,N_415);
nor U964 (N_964,N_623,N_356);
nand U965 (N_965,In_1068,N_615);
or U966 (N_966,In_674,N_697);
nor U967 (N_967,In_967,N_514);
or U968 (N_968,In_1445,In_1186);
and U969 (N_969,In_577,In_1386);
nor U970 (N_970,N_94,N_258);
or U971 (N_971,N_92,N_680);
or U972 (N_972,In_457,N_433);
and U973 (N_973,N_121,N_503);
nor U974 (N_974,In_166,N_184);
and U975 (N_975,N_158,N_611);
nor U976 (N_976,N_523,N_408);
and U977 (N_977,In_1484,N_322);
and U978 (N_978,N_482,In_509);
xor U979 (N_979,N_108,N_52);
and U980 (N_980,N_586,N_351);
nor U981 (N_981,N_641,In_343);
xor U982 (N_982,N_550,N_413);
nor U983 (N_983,N_674,N_534);
nand U984 (N_984,N_628,N_658);
or U985 (N_985,N_579,In_332);
xor U986 (N_986,N_694,In_1256);
or U987 (N_987,N_645,In_302);
or U988 (N_988,N_346,In_807);
nor U989 (N_989,In_929,In_1005);
or U990 (N_990,In_373,N_698);
xor U991 (N_991,N_730,In_1379);
xnor U992 (N_992,In_510,In_1004);
nand U993 (N_993,N_300,N_336);
xnor U994 (N_994,N_306,In_146);
or U995 (N_995,N_613,In_165);
xor U996 (N_996,N_728,N_528);
nand U997 (N_997,N_671,N_556);
and U998 (N_998,N_288,N_633);
nand U999 (N_999,N_369,N_465);
nor U1000 (N_1000,N_770,N_249);
nand U1001 (N_1001,N_785,N_842);
and U1002 (N_1002,N_950,N_638);
xor U1003 (N_1003,In_1318,In_1143);
and U1004 (N_1004,N_572,N_940);
or U1005 (N_1005,N_359,N_846);
and U1006 (N_1006,N_532,In_874);
xnor U1007 (N_1007,N_261,In_1077);
or U1008 (N_1008,N_769,N_619);
or U1009 (N_1009,N_912,N_911);
nor U1010 (N_1010,N_844,N_747);
nand U1011 (N_1011,N_636,In_1426);
nor U1012 (N_1012,N_861,N_515);
and U1013 (N_1013,N_920,N_802);
nand U1014 (N_1014,N_357,N_690);
nand U1015 (N_1015,In_1011,N_901);
xnor U1016 (N_1016,N_373,In_69);
xnor U1017 (N_1017,N_763,N_836);
xnor U1018 (N_1018,N_977,N_462);
and U1019 (N_1019,N_363,N_673);
nand U1020 (N_1020,N_992,N_841);
xnor U1021 (N_1021,N_277,N_682);
xnor U1022 (N_1022,N_656,N_856);
or U1023 (N_1023,N_761,N_818);
and U1024 (N_1024,N_603,In_1127);
and U1025 (N_1025,N_819,N_788);
or U1026 (N_1026,N_416,N_937);
or U1027 (N_1027,N_948,In_334);
xnor U1028 (N_1028,In_425,N_882);
xnor U1029 (N_1029,N_809,In_1251);
or U1030 (N_1030,N_254,N_601);
nor U1031 (N_1031,In_1411,N_835);
nor U1032 (N_1032,N_975,N_953);
and U1033 (N_1033,In_524,N_828);
and U1034 (N_1034,N_773,N_814);
nand U1035 (N_1035,N_993,N_851);
nor U1036 (N_1036,N_891,N_839);
nor U1037 (N_1037,N_608,N_248);
and U1038 (N_1038,N_587,N_796);
xor U1039 (N_1039,In_552,N_1);
nor U1040 (N_1040,N_634,In_1009);
or U1041 (N_1041,In_1206,N_143);
nor U1042 (N_1042,N_947,N_877);
nand U1043 (N_1043,N_643,N_605);
xnor U1044 (N_1044,N_779,N_906);
nand U1045 (N_1045,N_996,N_383);
nand U1046 (N_1046,N_869,In_954);
or U1047 (N_1047,In_446,N_595);
nand U1048 (N_1048,N_749,In_677);
and U1049 (N_1049,In_62,N_966);
nor U1050 (N_1050,N_406,N_630);
and U1051 (N_1051,N_898,N_423);
xnor U1052 (N_1052,In_225,In_622);
xor U1053 (N_1053,N_713,N_717);
nand U1054 (N_1054,N_439,In_1300);
or U1055 (N_1055,N_684,N_710);
nor U1056 (N_1056,N_959,N_616);
and U1057 (N_1057,N_172,N_908);
nor U1058 (N_1058,N_15,N_867);
and U1059 (N_1059,N_870,In_414);
nor U1060 (N_1060,N_957,N_822);
xnor U1061 (N_1061,N_566,N_798);
and U1062 (N_1062,N_175,N_368);
nor U1063 (N_1063,In_415,N_881);
or U1064 (N_1064,N_873,N_897);
nor U1065 (N_1065,N_626,N_293);
nor U1066 (N_1066,N_800,N_509);
and U1067 (N_1067,In_136,N_958);
nand U1068 (N_1068,N_917,N_803);
and U1069 (N_1069,In_1111,N_827);
xnor U1070 (N_1070,N_878,N_964);
nand U1071 (N_1071,N_843,N_189);
nand U1072 (N_1072,N_653,N_12);
nor U1073 (N_1073,N_219,N_789);
nand U1074 (N_1074,In_1002,N_539);
or U1075 (N_1075,N_548,In_1262);
xor U1076 (N_1076,N_663,N_793);
nor U1077 (N_1077,N_960,N_916);
nor U1078 (N_1078,N_962,N_990);
nor U1079 (N_1079,In_99,N_840);
and U1080 (N_1080,N_781,In_1182);
nor U1081 (N_1081,N_942,N_721);
xor U1082 (N_1082,N_933,N_857);
and U1083 (N_1083,N_875,N_521);
xnor U1084 (N_1084,In_569,N_227);
nand U1085 (N_1085,N_808,N_455);
xnor U1086 (N_1086,N_874,N_771);
and U1087 (N_1087,N_986,N_815);
or U1088 (N_1088,In_1385,N_995);
or U1089 (N_1089,N_907,N_762);
or U1090 (N_1090,N_527,In_1392);
or U1091 (N_1091,N_983,In_631);
xnor U1092 (N_1092,In_114,N_801);
xor U1093 (N_1093,N_994,In_959);
and U1094 (N_1094,N_941,N_894);
nor U1095 (N_1095,N_502,In_1200);
and U1096 (N_1096,N_755,N_830);
or U1097 (N_1097,N_943,N_309);
or U1098 (N_1098,N_409,N_775);
or U1099 (N_1099,N_743,N_871);
nor U1100 (N_1100,N_921,In_141);
nand U1101 (N_1101,N_949,N_931);
nor U1102 (N_1102,N_753,N_498);
and U1103 (N_1103,N_443,In_1286);
xor U1104 (N_1104,N_778,N_273);
xnor U1105 (N_1105,N_722,N_701);
and U1106 (N_1106,N_930,N_845);
nor U1107 (N_1107,N_919,N_969);
or U1108 (N_1108,In_437,N_890);
xnor U1109 (N_1109,N_782,In_1375);
and U1110 (N_1110,N_596,In_786);
or U1111 (N_1111,N_487,N_715);
nor U1112 (N_1112,N_620,In_1207);
nor U1113 (N_1113,In_1272,N_945);
xor U1114 (N_1114,N_859,N_224);
or U1115 (N_1115,N_812,N_105);
and U1116 (N_1116,In_1190,N_345);
nor U1117 (N_1117,N_847,N_665);
or U1118 (N_1118,N_214,N_766);
nor U1119 (N_1119,In_1128,N_888);
or U1120 (N_1120,N_622,In_1080);
or U1121 (N_1121,N_685,N_560);
nand U1122 (N_1122,N_558,N_491);
or U1123 (N_1123,N_886,N_862);
nor U1124 (N_1124,N_925,In_1435);
xor U1125 (N_1125,N_849,N_853);
and U1126 (N_1126,In_1474,N_952);
or U1127 (N_1127,N_600,N_795);
and U1128 (N_1128,N_999,N_790);
xnor U1129 (N_1129,N_588,N_222);
xor U1130 (N_1130,N_765,N_981);
or U1131 (N_1131,In_1296,N_985);
xnor U1132 (N_1132,In_1147,N_825);
nand U1133 (N_1133,N_922,N_632);
and U1134 (N_1134,N_341,N_924);
xnor U1135 (N_1135,N_967,N_971);
nor U1136 (N_1136,N_792,N_302);
and U1137 (N_1137,N_932,N_426);
xor U1138 (N_1138,N_887,N_885);
or U1139 (N_1139,N_903,In_555);
nand U1140 (N_1140,N_978,N_252);
nand U1141 (N_1141,N_444,N_435);
or U1142 (N_1142,N_192,N_759);
nor U1143 (N_1143,N_546,N_935);
nor U1144 (N_1144,N_688,N_872);
xor U1145 (N_1145,In_1007,N_791);
nand U1146 (N_1146,N_864,N_654);
and U1147 (N_1147,In_589,N_889);
and U1148 (N_1148,N_758,N_936);
nand U1149 (N_1149,N_545,N_883);
or U1150 (N_1150,N_750,N_530);
nor U1151 (N_1151,N_961,N_589);
nand U1152 (N_1152,N_834,N_973);
nor U1153 (N_1153,N_909,In_71);
xnor U1154 (N_1154,N_824,N_70);
or U1155 (N_1155,N_642,N_787);
and U1156 (N_1156,N_768,N_291);
xnor U1157 (N_1157,N_972,N_879);
xor U1158 (N_1158,N_756,In_63);
xor U1159 (N_1159,N_315,N_979);
and U1160 (N_1160,N_681,N_754);
nor U1161 (N_1161,N_831,N_422);
or U1162 (N_1162,N_915,N_578);
or U1163 (N_1163,In_1085,In_1099);
nor U1164 (N_1164,In_223,N_982);
or U1165 (N_1165,N_811,N_580);
and U1166 (N_1166,N_757,N_866);
or U1167 (N_1167,In_423,N_852);
xor U1168 (N_1168,N_441,N_826);
and U1169 (N_1169,N_776,N_236);
nor U1170 (N_1170,N_837,N_661);
and U1171 (N_1171,In_1309,N_850);
nor U1172 (N_1172,N_910,In_883);
and U1173 (N_1173,N_980,In_186);
nand U1174 (N_1174,N_860,N_829);
xnor U1175 (N_1175,N_751,N_833);
and U1176 (N_1176,N_938,N_486);
xor U1177 (N_1177,N_820,In_976);
and U1178 (N_1178,N_880,N_900);
xnor U1179 (N_1179,N_956,In_1370);
xnor U1180 (N_1180,N_951,N_895);
and U1181 (N_1181,In_383,In_72);
or U1182 (N_1182,N_537,N_863);
xnor U1183 (N_1183,In_1053,N_524);
and U1184 (N_1184,N_892,N_429);
or U1185 (N_1185,N_904,N_902);
nor U1186 (N_1186,N_823,N_731);
or U1187 (N_1187,N_695,N_968);
xor U1188 (N_1188,N_627,N_913);
nor U1189 (N_1189,N_477,N_419);
and U1190 (N_1190,N_784,N_215);
or U1191 (N_1191,N_760,N_868);
and U1192 (N_1192,In_1475,N_772);
nand U1193 (N_1193,In_1032,N_670);
xor U1194 (N_1194,N_535,In_1279);
or U1195 (N_1195,In_1451,N_574);
or U1196 (N_1196,N_816,N_767);
nand U1197 (N_1197,N_926,In_602);
or U1198 (N_1198,N_699,N_618);
xor U1199 (N_1199,N_284,N_984);
xor U1200 (N_1200,In_838,N_832);
or U1201 (N_1201,In_487,N_536);
nor U1202 (N_1202,N_325,N_547);
nor U1203 (N_1203,N_591,N_594);
nor U1204 (N_1204,N_780,In_597);
nor U1205 (N_1205,N_774,N_970);
and U1206 (N_1206,N_848,In_599);
nand U1207 (N_1207,N_807,In_1208);
and U1208 (N_1208,N_854,N_965);
xor U1209 (N_1209,In_1019,N_646);
xor U1210 (N_1210,N_899,In_852);
nand U1211 (N_1211,N_923,In_1244);
nor U1212 (N_1212,N_954,In_1472);
or U1213 (N_1213,N_963,In_665);
nand U1214 (N_1214,N_821,In_576);
nor U1215 (N_1215,N_147,N_927);
and U1216 (N_1216,N_928,N_542);
nand U1217 (N_1217,N_944,N_799);
or U1218 (N_1218,N_797,N_865);
and U1219 (N_1219,N_72,N_805);
nand U1220 (N_1220,N_804,N_162);
nand U1221 (N_1221,N_893,N_855);
or U1222 (N_1222,N_810,N_997);
nor U1223 (N_1223,N_929,N_783);
xor U1224 (N_1224,N_794,N_664);
xor U1225 (N_1225,N_918,N_333);
nor U1226 (N_1226,N_691,N_934);
and U1227 (N_1227,N_974,N_777);
nor U1228 (N_1228,In_571,In_14);
nor U1229 (N_1229,N_998,N_752);
nor U1230 (N_1230,N_905,In_1098);
xor U1231 (N_1231,In_349,N_360);
nand U1232 (N_1232,N_988,N_764);
nand U1233 (N_1233,N_786,N_549);
and U1234 (N_1234,N_417,N_991);
nand U1235 (N_1235,N_989,N_876);
and U1236 (N_1236,N_813,N_914);
or U1237 (N_1237,N_858,N_744);
nand U1238 (N_1238,In_778,N_939);
nor U1239 (N_1239,N_267,N_955);
and U1240 (N_1240,N_573,N_568);
nand U1241 (N_1241,N_817,N_946);
nor U1242 (N_1242,N_884,N_734);
or U1243 (N_1243,N_987,N_541);
and U1244 (N_1244,N_976,N_500);
nor U1245 (N_1245,N_526,In_618);
xor U1246 (N_1246,In_16,N_838);
and U1247 (N_1247,N_609,N_806);
nand U1248 (N_1248,N_896,N_109);
nand U1249 (N_1249,In_224,N_229);
nor U1250 (N_1250,N_1133,N_1162);
nor U1251 (N_1251,N_1059,N_1093);
nor U1252 (N_1252,N_1129,N_1236);
or U1253 (N_1253,N_1148,N_1001);
or U1254 (N_1254,N_1054,N_1003);
xor U1255 (N_1255,N_1026,N_1194);
xnor U1256 (N_1256,N_1110,N_1069);
nand U1257 (N_1257,N_1083,N_1157);
and U1258 (N_1258,N_1113,N_1219);
xnor U1259 (N_1259,N_1057,N_1099);
and U1260 (N_1260,N_1237,N_1096);
xor U1261 (N_1261,N_1240,N_1078);
nor U1262 (N_1262,N_1092,N_1227);
and U1263 (N_1263,N_1156,N_1060);
nand U1264 (N_1264,N_1152,N_1126);
or U1265 (N_1265,N_1010,N_1134);
or U1266 (N_1266,N_1241,N_1072);
nand U1267 (N_1267,N_1013,N_1064);
or U1268 (N_1268,N_1051,N_1031);
xnor U1269 (N_1269,N_1104,N_1128);
or U1270 (N_1270,N_1008,N_1208);
and U1271 (N_1271,N_1205,N_1226);
xor U1272 (N_1272,N_1118,N_1087);
nand U1273 (N_1273,N_1039,N_1005);
or U1274 (N_1274,N_1027,N_1169);
nand U1275 (N_1275,N_1167,N_1102);
and U1276 (N_1276,N_1040,N_1207);
or U1277 (N_1277,N_1066,N_1018);
and U1278 (N_1278,N_1090,N_1037);
nor U1279 (N_1279,N_1124,N_1084);
or U1280 (N_1280,N_1015,N_1123);
xnor U1281 (N_1281,N_1197,N_1000);
nand U1282 (N_1282,N_1075,N_1222);
nand U1283 (N_1283,N_1245,N_1213);
nor U1284 (N_1284,N_1056,N_1105);
nand U1285 (N_1285,N_1136,N_1085);
nand U1286 (N_1286,N_1188,N_1025);
xnor U1287 (N_1287,N_1074,N_1073);
xor U1288 (N_1288,N_1142,N_1199);
nand U1289 (N_1289,N_1247,N_1082);
xnor U1290 (N_1290,N_1233,N_1146);
xor U1291 (N_1291,N_1230,N_1112);
nand U1292 (N_1292,N_1007,N_1243);
nand U1293 (N_1293,N_1165,N_1049);
xnor U1294 (N_1294,N_1019,N_1016);
nor U1295 (N_1295,N_1065,N_1140);
and U1296 (N_1296,N_1130,N_1176);
or U1297 (N_1297,N_1042,N_1097);
nor U1298 (N_1298,N_1221,N_1212);
xnor U1299 (N_1299,N_1145,N_1101);
nand U1300 (N_1300,N_1232,N_1137);
nand U1301 (N_1301,N_1242,N_1190);
or U1302 (N_1302,N_1038,N_1191);
xnor U1303 (N_1303,N_1211,N_1131);
nor U1304 (N_1304,N_1114,N_1006);
nor U1305 (N_1305,N_1185,N_1067);
nand U1306 (N_1306,N_1091,N_1011);
and U1307 (N_1307,N_1249,N_1076);
nor U1308 (N_1308,N_1228,N_1106);
and U1309 (N_1309,N_1047,N_1141);
nor U1310 (N_1310,N_1021,N_1044);
or U1311 (N_1311,N_1159,N_1171);
xor U1312 (N_1312,N_1043,N_1132);
nand U1313 (N_1313,N_1210,N_1238);
or U1314 (N_1314,N_1052,N_1229);
and U1315 (N_1315,N_1111,N_1070);
nor U1316 (N_1316,N_1138,N_1095);
or U1317 (N_1317,N_1173,N_1028);
xor U1318 (N_1318,N_1217,N_1023);
nand U1319 (N_1319,N_1081,N_1122);
and U1320 (N_1320,N_1154,N_1223);
xnor U1321 (N_1321,N_1046,N_1135);
or U1322 (N_1322,N_1048,N_1115);
nor U1323 (N_1323,N_1149,N_1094);
nor U1324 (N_1324,N_1166,N_1235);
or U1325 (N_1325,N_1024,N_1062);
and U1326 (N_1326,N_1035,N_1218);
xor U1327 (N_1327,N_1186,N_1151);
nand U1328 (N_1328,N_1161,N_1068);
nand U1329 (N_1329,N_1220,N_1170);
or U1330 (N_1330,N_1187,N_1120);
and U1331 (N_1331,N_1125,N_1127);
xnor U1332 (N_1332,N_1203,N_1164);
or U1333 (N_1333,N_1189,N_1178);
nor U1334 (N_1334,N_1050,N_1200);
and U1335 (N_1335,N_1030,N_1244);
or U1336 (N_1336,N_1175,N_1103);
nor U1337 (N_1337,N_1063,N_1079);
and U1338 (N_1338,N_1174,N_1179);
nor U1339 (N_1339,N_1248,N_1182);
or U1340 (N_1340,N_1116,N_1180);
xor U1341 (N_1341,N_1163,N_1139);
and U1342 (N_1342,N_1196,N_1225);
or U1343 (N_1343,N_1246,N_1193);
and U1344 (N_1344,N_1158,N_1109);
xnor U1345 (N_1345,N_1041,N_1231);
nand U1346 (N_1346,N_1058,N_1086);
or U1347 (N_1347,N_1029,N_1121);
xor U1348 (N_1348,N_1032,N_1034);
nand U1349 (N_1349,N_1215,N_1239);
nand U1350 (N_1350,N_1234,N_1160);
nor U1351 (N_1351,N_1061,N_1033);
xor U1352 (N_1352,N_1004,N_1045);
or U1353 (N_1353,N_1192,N_1009);
or U1354 (N_1354,N_1053,N_1071);
nor U1355 (N_1355,N_1107,N_1144);
nand U1356 (N_1356,N_1036,N_1181);
nor U1357 (N_1357,N_1055,N_1150);
xnor U1358 (N_1358,N_1201,N_1143);
nor U1359 (N_1359,N_1119,N_1172);
nand U1360 (N_1360,N_1177,N_1002);
nor U1361 (N_1361,N_1216,N_1184);
and U1362 (N_1362,N_1088,N_1077);
or U1363 (N_1363,N_1195,N_1108);
nor U1364 (N_1364,N_1224,N_1098);
or U1365 (N_1365,N_1100,N_1020);
xor U1366 (N_1366,N_1089,N_1147);
nand U1367 (N_1367,N_1117,N_1206);
or U1368 (N_1368,N_1209,N_1022);
nand U1369 (N_1369,N_1198,N_1153);
nand U1370 (N_1370,N_1202,N_1183);
and U1371 (N_1371,N_1214,N_1080);
nand U1372 (N_1372,N_1155,N_1204);
nor U1373 (N_1373,N_1014,N_1168);
and U1374 (N_1374,N_1012,N_1017);
and U1375 (N_1375,N_1111,N_1021);
and U1376 (N_1376,N_1092,N_1047);
or U1377 (N_1377,N_1209,N_1072);
or U1378 (N_1378,N_1008,N_1207);
and U1379 (N_1379,N_1189,N_1046);
nor U1380 (N_1380,N_1075,N_1161);
nor U1381 (N_1381,N_1233,N_1023);
nor U1382 (N_1382,N_1079,N_1130);
or U1383 (N_1383,N_1149,N_1117);
xor U1384 (N_1384,N_1087,N_1034);
nand U1385 (N_1385,N_1136,N_1113);
nand U1386 (N_1386,N_1050,N_1210);
nand U1387 (N_1387,N_1184,N_1031);
or U1388 (N_1388,N_1049,N_1080);
and U1389 (N_1389,N_1245,N_1065);
nand U1390 (N_1390,N_1244,N_1000);
nor U1391 (N_1391,N_1245,N_1001);
xor U1392 (N_1392,N_1239,N_1207);
and U1393 (N_1393,N_1076,N_1170);
and U1394 (N_1394,N_1166,N_1203);
nor U1395 (N_1395,N_1060,N_1193);
and U1396 (N_1396,N_1009,N_1227);
nor U1397 (N_1397,N_1197,N_1048);
nor U1398 (N_1398,N_1185,N_1133);
and U1399 (N_1399,N_1173,N_1074);
and U1400 (N_1400,N_1067,N_1124);
and U1401 (N_1401,N_1023,N_1076);
or U1402 (N_1402,N_1121,N_1027);
nand U1403 (N_1403,N_1020,N_1217);
and U1404 (N_1404,N_1225,N_1234);
xor U1405 (N_1405,N_1036,N_1247);
xor U1406 (N_1406,N_1209,N_1141);
and U1407 (N_1407,N_1118,N_1156);
nor U1408 (N_1408,N_1166,N_1165);
nand U1409 (N_1409,N_1045,N_1237);
xor U1410 (N_1410,N_1096,N_1094);
nor U1411 (N_1411,N_1241,N_1178);
nand U1412 (N_1412,N_1080,N_1040);
xor U1413 (N_1413,N_1225,N_1022);
or U1414 (N_1414,N_1142,N_1195);
or U1415 (N_1415,N_1043,N_1068);
or U1416 (N_1416,N_1075,N_1062);
and U1417 (N_1417,N_1230,N_1099);
xor U1418 (N_1418,N_1219,N_1117);
nand U1419 (N_1419,N_1176,N_1249);
and U1420 (N_1420,N_1128,N_1132);
nor U1421 (N_1421,N_1119,N_1156);
nor U1422 (N_1422,N_1033,N_1180);
nand U1423 (N_1423,N_1079,N_1018);
and U1424 (N_1424,N_1000,N_1232);
and U1425 (N_1425,N_1033,N_1073);
or U1426 (N_1426,N_1100,N_1128);
nor U1427 (N_1427,N_1055,N_1193);
or U1428 (N_1428,N_1239,N_1143);
xor U1429 (N_1429,N_1015,N_1057);
and U1430 (N_1430,N_1133,N_1184);
nand U1431 (N_1431,N_1085,N_1017);
nor U1432 (N_1432,N_1181,N_1236);
nand U1433 (N_1433,N_1197,N_1002);
xor U1434 (N_1434,N_1168,N_1050);
nand U1435 (N_1435,N_1244,N_1174);
nor U1436 (N_1436,N_1244,N_1241);
nor U1437 (N_1437,N_1133,N_1030);
nor U1438 (N_1438,N_1043,N_1202);
and U1439 (N_1439,N_1025,N_1153);
nand U1440 (N_1440,N_1152,N_1213);
nand U1441 (N_1441,N_1159,N_1222);
nand U1442 (N_1442,N_1225,N_1190);
nor U1443 (N_1443,N_1046,N_1058);
or U1444 (N_1444,N_1051,N_1192);
nor U1445 (N_1445,N_1020,N_1058);
or U1446 (N_1446,N_1009,N_1099);
nor U1447 (N_1447,N_1211,N_1224);
or U1448 (N_1448,N_1115,N_1021);
and U1449 (N_1449,N_1065,N_1097);
xor U1450 (N_1450,N_1064,N_1247);
nand U1451 (N_1451,N_1247,N_1060);
nor U1452 (N_1452,N_1057,N_1026);
nor U1453 (N_1453,N_1202,N_1052);
nand U1454 (N_1454,N_1015,N_1061);
xnor U1455 (N_1455,N_1064,N_1021);
nand U1456 (N_1456,N_1052,N_1075);
xor U1457 (N_1457,N_1062,N_1219);
xnor U1458 (N_1458,N_1100,N_1190);
nand U1459 (N_1459,N_1185,N_1005);
and U1460 (N_1460,N_1010,N_1192);
nand U1461 (N_1461,N_1063,N_1194);
or U1462 (N_1462,N_1156,N_1226);
or U1463 (N_1463,N_1084,N_1249);
and U1464 (N_1464,N_1226,N_1039);
nand U1465 (N_1465,N_1240,N_1179);
nor U1466 (N_1466,N_1220,N_1134);
nand U1467 (N_1467,N_1223,N_1029);
and U1468 (N_1468,N_1217,N_1153);
and U1469 (N_1469,N_1153,N_1105);
nand U1470 (N_1470,N_1010,N_1208);
and U1471 (N_1471,N_1014,N_1141);
and U1472 (N_1472,N_1214,N_1188);
nand U1473 (N_1473,N_1032,N_1026);
xor U1474 (N_1474,N_1166,N_1190);
and U1475 (N_1475,N_1149,N_1200);
or U1476 (N_1476,N_1180,N_1058);
or U1477 (N_1477,N_1049,N_1024);
xor U1478 (N_1478,N_1166,N_1216);
xor U1479 (N_1479,N_1046,N_1174);
or U1480 (N_1480,N_1061,N_1055);
nand U1481 (N_1481,N_1182,N_1030);
nand U1482 (N_1482,N_1101,N_1208);
nor U1483 (N_1483,N_1089,N_1006);
or U1484 (N_1484,N_1024,N_1164);
nand U1485 (N_1485,N_1220,N_1146);
and U1486 (N_1486,N_1011,N_1242);
or U1487 (N_1487,N_1109,N_1053);
or U1488 (N_1488,N_1199,N_1130);
or U1489 (N_1489,N_1051,N_1058);
and U1490 (N_1490,N_1088,N_1214);
and U1491 (N_1491,N_1224,N_1050);
and U1492 (N_1492,N_1108,N_1096);
nand U1493 (N_1493,N_1240,N_1234);
xor U1494 (N_1494,N_1071,N_1136);
nor U1495 (N_1495,N_1038,N_1036);
xor U1496 (N_1496,N_1240,N_1061);
and U1497 (N_1497,N_1215,N_1123);
nor U1498 (N_1498,N_1017,N_1052);
nor U1499 (N_1499,N_1101,N_1173);
xor U1500 (N_1500,N_1350,N_1344);
xnor U1501 (N_1501,N_1487,N_1271);
nand U1502 (N_1502,N_1282,N_1431);
xor U1503 (N_1503,N_1278,N_1415);
xor U1504 (N_1504,N_1286,N_1291);
nor U1505 (N_1505,N_1296,N_1311);
and U1506 (N_1506,N_1378,N_1470);
nor U1507 (N_1507,N_1460,N_1448);
or U1508 (N_1508,N_1413,N_1375);
nor U1509 (N_1509,N_1301,N_1492);
nor U1510 (N_1510,N_1373,N_1370);
xor U1511 (N_1511,N_1351,N_1359);
nand U1512 (N_1512,N_1357,N_1442);
nor U1513 (N_1513,N_1485,N_1428);
or U1514 (N_1514,N_1489,N_1406);
or U1515 (N_1515,N_1443,N_1257);
and U1516 (N_1516,N_1481,N_1410);
or U1517 (N_1517,N_1387,N_1440);
or U1518 (N_1518,N_1273,N_1491);
nand U1519 (N_1519,N_1379,N_1260);
nor U1520 (N_1520,N_1386,N_1272);
and U1521 (N_1521,N_1416,N_1496);
nor U1522 (N_1522,N_1333,N_1303);
nand U1523 (N_1523,N_1289,N_1306);
or U1524 (N_1524,N_1288,N_1399);
and U1525 (N_1525,N_1336,N_1316);
xnor U1526 (N_1526,N_1456,N_1477);
nor U1527 (N_1527,N_1328,N_1281);
nor U1528 (N_1528,N_1352,N_1262);
or U1529 (N_1529,N_1374,N_1309);
and U1530 (N_1530,N_1381,N_1455);
nor U1531 (N_1531,N_1433,N_1444);
xor U1532 (N_1532,N_1466,N_1339);
and U1533 (N_1533,N_1364,N_1493);
nor U1534 (N_1534,N_1422,N_1361);
and U1535 (N_1535,N_1312,N_1467);
nor U1536 (N_1536,N_1363,N_1330);
nand U1537 (N_1537,N_1277,N_1497);
nand U1538 (N_1538,N_1382,N_1356);
nor U1539 (N_1539,N_1384,N_1326);
or U1540 (N_1540,N_1294,N_1459);
or U1541 (N_1541,N_1426,N_1342);
nand U1542 (N_1542,N_1494,N_1395);
or U1543 (N_1543,N_1343,N_1365);
nor U1544 (N_1544,N_1321,N_1441);
and U1545 (N_1545,N_1334,N_1264);
and U1546 (N_1546,N_1376,N_1347);
nand U1547 (N_1547,N_1469,N_1451);
or U1548 (N_1548,N_1325,N_1421);
or U1549 (N_1549,N_1367,N_1394);
xnor U1550 (N_1550,N_1340,N_1423);
and U1551 (N_1551,N_1420,N_1358);
nand U1552 (N_1552,N_1298,N_1317);
nand U1553 (N_1553,N_1323,N_1471);
xor U1554 (N_1554,N_1267,N_1414);
xor U1555 (N_1555,N_1337,N_1253);
nor U1556 (N_1556,N_1424,N_1419);
nor U1557 (N_1557,N_1427,N_1432);
nor U1558 (N_1558,N_1322,N_1452);
and U1559 (N_1559,N_1258,N_1266);
nor U1560 (N_1560,N_1393,N_1256);
nor U1561 (N_1561,N_1478,N_1255);
and U1562 (N_1562,N_1369,N_1283);
xnor U1563 (N_1563,N_1429,N_1486);
nor U1564 (N_1564,N_1483,N_1315);
nor U1565 (N_1565,N_1263,N_1476);
or U1566 (N_1566,N_1304,N_1310);
or U1567 (N_1567,N_1360,N_1465);
and U1568 (N_1568,N_1252,N_1391);
and U1569 (N_1569,N_1468,N_1474);
or U1570 (N_1570,N_1464,N_1450);
nand U1571 (N_1571,N_1409,N_1348);
xor U1572 (N_1572,N_1318,N_1280);
nor U1573 (N_1573,N_1307,N_1453);
nand U1574 (N_1574,N_1411,N_1439);
and U1575 (N_1575,N_1377,N_1498);
nor U1576 (N_1576,N_1259,N_1276);
or U1577 (N_1577,N_1355,N_1462);
and U1578 (N_1578,N_1314,N_1473);
and U1579 (N_1579,N_1366,N_1446);
and U1580 (N_1580,N_1401,N_1482);
nor U1581 (N_1581,N_1324,N_1472);
nor U1582 (N_1582,N_1418,N_1402);
nand U1583 (N_1583,N_1495,N_1284);
nand U1584 (N_1584,N_1463,N_1308);
nor U1585 (N_1585,N_1269,N_1396);
or U1586 (N_1586,N_1438,N_1372);
nor U1587 (N_1587,N_1254,N_1454);
nand U1588 (N_1588,N_1354,N_1265);
nand U1589 (N_1589,N_1405,N_1346);
and U1590 (N_1590,N_1435,N_1295);
nor U1591 (N_1591,N_1449,N_1397);
nor U1592 (N_1592,N_1484,N_1480);
nand U1593 (N_1593,N_1488,N_1457);
nor U1594 (N_1594,N_1251,N_1368);
and U1595 (N_1595,N_1403,N_1292);
or U1596 (N_1596,N_1274,N_1293);
or U1597 (N_1597,N_1353,N_1341);
or U1598 (N_1598,N_1407,N_1299);
xor U1599 (N_1599,N_1445,N_1327);
or U1600 (N_1600,N_1279,N_1331);
nand U1601 (N_1601,N_1285,N_1250);
nor U1602 (N_1602,N_1287,N_1261);
nor U1603 (N_1603,N_1398,N_1362);
or U1604 (N_1604,N_1447,N_1412);
or U1605 (N_1605,N_1268,N_1389);
nor U1606 (N_1606,N_1479,N_1388);
nand U1607 (N_1607,N_1297,N_1408);
or U1608 (N_1608,N_1475,N_1320);
nand U1609 (N_1609,N_1392,N_1319);
xnor U1610 (N_1610,N_1302,N_1461);
xnor U1611 (N_1611,N_1425,N_1371);
xor U1612 (N_1612,N_1390,N_1436);
nor U1613 (N_1613,N_1275,N_1329);
xor U1614 (N_1614,N_1499,N_1434);
or U1615 (N_1615,N_1437,N_1305);
nand U1616 (N_1616,N_1349,N_1490);
or U1617 (N_1617,N_1380,N_1430);
and U1618 (N_1618,N_1270,N_1338);
nor U1619 (N_1619,N_1385,N_1417);
nand U1620 (N_1620,N_1345,N_1332);
and U1621 (N_1621,N_1313,N_1458);
or U1622 (N_1622,N_1400,N_1290);
nand U1623 (N_1623,N_1404,N_1335);
nand U1624 (N_1624,N_1300,N_1383);
and U1625 (N_1625,N_1308,N_1315);
and U1626 (N_1626,N_1406,N_1355);
xor U1627 (N_1627,N_1251,N_1258);
xor U1628 (N_1628,N_1256,N_1342);
nand U1629 (N_1629,N_1475,N_1409);
nor U1630 (N_1630,N_1273,N_1348);
nor U1631 (N_1631,N_1361,N_1485);
xnor U1632 (N_1632,N_1346,N_1381);
or U1633 (N_1633,N_1342,N_1347);
nor U1634 (N_1634,N_1429,N_1353);
nand U1635 (N_1635,N_1272,N_1287);
nand U1636 (N_1636,N_1298,N_1353);
nor U1637 (N_1637,N_1319,N_1291);
nand U1638 (N_1638,N_1358,N_1439);
or U1639 (N_1639,N_1290,N_1272);
nor U1640 (N_1640,N_1354,N_1303);
xnor U1641 (N_1641,N_1319,N_1473);
and U1642 (N_1642,N_1389,N_1291);
nand U1643 (N_1643,N_1466,N_1415);
xnor U1644 (N_1644,N_1370,N_1266);
or U1645 (N_1645,N_1324,N_1366);
nand U1646 (N_1646,N_1393,N_1441);
nand U1647 (N_1647,N_1385,N_1445);
and U1648 (N_1648,N_1390,N_1375);
and U1649 (N_1649,N_1316,N_1268);
nor U1650 (N_1650,N_1431,N_1422);
nor U1651 (N_1651,N_1347,N_1462);
nor U1652 (N_1652,N_1365,N_1342);
or U1653 (N_1653,N_1489,N_1417);
or U1654 (N_1654,N_1468,N_1459);
and U1655 (N_1655,N_1431,N_1462);
nand U1656 (N_1656,N_1301,N_1408);
nand U1657 (N_1657,N_1457,N_1406);
nor U1658 (N_1658,N_1400,N_1476);
nor U1659 (N_1659,N_1444,N_1282);
nor U1660 (N_1660,N_1295,N_1459);
nor U1661 (N_1661,N_1401,N_1442);
xnor U1662 (N_1662,N_1412,N_1432);
nand U1663 (N_1663,N_1329,N_1305);
xnor U1664 (N_1664,N_1255,N_1351);
or U1665 (N_1665,N_1384,N_1358);
and U1666 (N_1666,N_1497,N_1462);
nand U1667 (N_1667,N_1263,N_1481);
and U1668 (N_1668,N_1277,N_1348);
and U1669 (N_1669,N_1314,N_1290);
or U1670 (N_1670,N_1307,N_1451);
xor U1671 (N_1671,N_1399,N_1385);
and U1672 (N_1672,N_1321,N_1481);
xnor U1673 (N_1673,N_1358,N_1457);
xor U1674 (N_1674,N_1331,N_1306);
nand U1675 (N_1675,N_1384,N_1396);
xor U1676 (N_1676,N_1353,N_1287);
or U1677 (N_1677,N_1454,N_1429);
nand U1678 (N_1678,N_1347,N_1323);
nand U1679 (N_1679,N_1333,N_1481);
and U1680 (N_1680,N_1390,N_1362);
nor U1681 (N_1681,N_1280,N_1297);
xnor U1682 (N_1682,N_1498,N_1296);
and U1683 (N_1683,N_1423,N_1386);
xnor U1684 (N_1684,N_1259,N_1288);
or U1685 (N_1685,N_1454,N_1491);
nand U1686 (N_1686,N_1475,N_1335);
or U1687 (N_1687,N_1410,N_1478);
nor U1688 (N_1688,N_1274,N_1256);
nand U1689 (N_1689,N_1490,N_1411);
or U1690 (N_1690,N_1470,N_1483);
nand U1691 (N_1691,N_1390,N_1328);
and U1692 (N_1692,N_1479,N_1266);
xnor U1693 (N_1693,N_1464,N_1299);
and U1694 (N_1694,N_1392,N_1415);
nor U1695 (N_1695,N_1469,N_1372);
xor U1696 (N_1696,N_1283,N_1484);
or U1697 (N_1697,N_1428,N_1440);
and U1698 (N_1698,N_1381,N_1413);
or U1699 (N_1699,N_1363,N_1325);
xor U1700 (N_1700,N_1266,N_1476);
or U1701 (N_1701,N_1390,N_1447);
nand U1702 (N_1702,N_1291,N_1498);
or U1703 (N_1703,N_1311,N_1413);
and U1704 (N_1704,N_1326,N_1424);
and U1705 (N_1705,N_1264,N_1365);
and U1706 (N_1706,N_1423,N_1338);
or U1707 (N_1707,N_1495,N_1424);
and U1708 (N_1708,N_1298,N_1327);
and U1709 (N_1709,N_1437,N_1489);
or U1710 (N_1710,N_1394,N_1441);
nor U1711 (N_1711,N_1483,N_1285);
or U1712 (N_1712,N_1347,N_1365);
and U1713 (N_1713,N_1322,N_1371);
xnor U1714 (N_1714,N_1393,N_1286);
xor U1715 (N_1715,N_1464,N_1413);
and U1716 (N_1716,N_1411,N_1341);
nor U1717 (N_1717,N_1434,N_1483);
nand U1718 (N_1718,N_1381,N_1285);
nand U1719 (N_1719,N_1350,N_1317);
or U1720 (N_1720,N_1480,N_1492);
xor U1721 (N_1721,N_1256,N_1329);
nand U1722 (N_1722,N_1351,N_1267);
nand U1723 (N_1723,N_1312,N_1426);
and U1724 (N_1724,N_1339,N_1289);
nor U1725 (N_1725,N_1366,N_1265);
or U1726 (N_1726,N_1390,N_1469);
nor U1727 (N_1727,N_1399,N_1383);
xor U1728 (N_1728,N_1467,N_1396);
or U1729 (N_1729,N_1398,N_1469);
xnor U1730 (N_1730,N_1386,N_1261);
xor U1731 (N_1731,N_1320,N_1404);
nand U1732 (N_1732,N_1463,N_1277);
nand U1733 (N_1733,N_1313,N_1302);
and U1734 (N_1734,N_1460,N_1404);
or U1735 (N_1735,N_1423,N_1404);
nand U1736 (N_1736,N_1390,N_1254);
xor U1737 (N_1737,N_1285,N_1480);
nor U1738 (N_1738,N_1390,N_1291);
and U1739 (N_1739,N_1347,N_1473);
or U1740 (N_1740,N_1376,N_1470);
nor U1741 (N_1741,N_1472,N_1340);
or U1742 (N_1742,N_1417,N_1391);
nand U1743 (N_1743,N_1324,N_1288);
or U1744 (N_1744,N_1300,N_1387);
or U1745 (N_1745,N_1498,N_1333);
nor U1746 (N_1746,N_1434,N_1390);
or U1747 (N_1747,N_1449,N_1351);
nor U1748 (N_1748,N_1470,N_1457);
and U1749 (N_1749,N_1413,N_1405);
nor U1750 (N_1750,N_1540,N_1663);
nor U1751 (N_1751,N_1612,N_1658);
and U1752 (N_1752,N_1742,N_1592);
and U1753 (N_1753,N_1546,N_1523);
nor U1754 (N_1754,N_1641,N_1739);
or U1755 (N_1755,N_1508,N_1733);
and U1756 (N_1756,N_1529,N_1655);
nand U1757 (N_1757,N_1677,N_1621);
or U1758 (N_1758,N_1571,N_1543);
and U1759 (N_1759,N_1578,N_1706);
xor U1760 (N_1760,N_1633,N_1747);
or U1761 (N_1761,N_1598,N_1712);
xor U1762 (N_1762,N_1718,N_1600);
or U1763 (N_1763,N_1613,N_1521);
and U1764 (N_1764,N_1535,N_1639);
nor U1765 (N_1765,N_1628,N_1515);
xor U1766 (N_1766,N_1642,N_1679);
and U1767 (N_1767,N_1653,N_1561);
and U1768 (N_1768,N_1737,N_1720);
xnor U1769 (N_1769,N_1630,N_1565);
nand U1770 (N_1770,N_1619,N_1601);
nor U1771 (N_1771,N_1549,N_1519);
nor U1772 (N_1772,N_1525,N_1729);
and U1773 (N_1773,N_1513,N_1645);
nor U1774 (N_1774,N_1577,N_1553);
or U1775 (N_1775,N_1596,N_1556);
or U1776 (N_1776,N_1744,N_1638);
or U1777 (N_1777,N_1656,N_1657);
and U1778 (N_1778,N_1659,N_1674);
nor U1779 (N_1779,N_1646,N_1579);
nor U1780 (N_1780,N_1688,N_1709);
or U1781 (N_1781,N_1607,N_1622);
nand U1782 (N_1782,N_1698,N_1667);
or U1783 (N_1783,N_1618,N_1554);
nand U1784 (N_1784,N_1584,N_1678);
and U1785 (N_1785,N_1572,N_1748);
or U1786 (N_1786,N_1620,N_1588);
and U1787 (N_1787,N_1662,N_1727);
xor U1788 (N_1788,N_1710,N_1551);
or U1789 (N_1789,N_1697,N_1568);
nand U1790 (N_1790,N_1722,N_1714);
or U1791 (N_1791,N_1696,N_1539);
nand U1792 (N_1792,N_1564,N_1616);
nor U1793 (N_1793,N_1567,N_1548);
xor U1794 (N_1794,N_1725,N_1627);
nand U1795 (N_1795,N_1651,N_1583);
nand U1796 (N_1796,N_1511,N_1603);
nand U1797 (N_1797,N_1581,N_1644);
xnor U1798 (N_1798,N_1575,N_1626);
and U1799 (N_1799,N_1558,N_1676);
and U1800 (N_1800,N_1640,N_1649);
and U1801 (N_1801,N_1695,N_1717);
nor U1802 (N_1802,N_1566,N_1602);
nor U1803 (N_1803,N_1623,N_1668);
nor U1804 (N_1804,N_1506,N_1501);
or U1805 (N_1805,N_1563,N_1636);
or U1806 (N_1806,N_1547,N_1541);
nor U1807 (N_1807,N_1586,N_1593);
and U1808 (N_1808,N_1504,N_1537);
or U1809 (N_1809,N_1634,N_1719);
nand U1810 (N_1810,N_1685,N_1605);
nand U1811 (N_1811,N_1721,N_1609);
nand U1812 (N_1812,N_1632,N_1587);
and U1813 (N_1813,N_1522,N_1694);
nor U1814 (N_1814,N_1716,N_1687);
nand U1815 (N_1815,N_1544,N_1517);
nand U1816 (N_1816,N_1562,N_1532);
and U1817 (N_1817,N_1680,N_1699);
xnor U1818 (N_1818,N_1538,N_1557);
xor U1819 (N_1819,N_1560,N_1713);
nand U1820 (N_1820,N_1731,N_1555);
nand U1821 (N_1821,N_1503,N_1617);
nand U1822 (N_1822,N_1711,N_1610);
or U1823 (N_1823,N_1732,N_1570);
or U1824 (N_1824,N_1512,N_1614);
and U1825 (N_1825,N_1684,N_1629);
and U1826 (N_1826,N_1664,N_1533);
xor U1827 (N_1827,N_1745,N_1700);
xor U1828 (N_1828,N_1736,N_1502);
xor U1829 (N_1829,N_1585,N_1580);
or U1830 (N_1830,N_1527,N_1734);
nand U1831 (N_1831,N_1749,N_1635);
xnor U1832 (N_1832,N_1589,N_1730);
nand U1833 (N_1833,N_1599,N_1665);
or U1834 (N_1834,N_1693,N_1650);
or U1835 (N_1835,N_1576,N_1595);
nand U1836 (N_1836,N_1643,N_1654);
and U1837 (N_1837,N_1735,N_1507);
and U1838 (N_1838,N_1704,N_1746);
and U1839 (N_1839,N_1569,N_1701);
nand U1840 (N_1840,N_1524,N_1724);
and U1841 (N_1841,N_1573,N_1670);
or U1842 (N_1842,N_1545,N_1590);
nor U1843 (N_1843,N_1597,N_1647);
nor U1844 (N_1844,N_1514,N_1715);
nor U1845 (N_1845,N_1669,N_1682);
and U1846 (N_1846,N_1606,N_1530);
xor U1847 (N_1847,N_1559,N_1690);
nand U1848 (N_1848,N_1666,N_1552);
or U1849 (N_1849,N_1691,N_1686);
xnor U1850 (N_1850,N_1681,N_1615);
xnor U1851 (N_1851,N_1526,N_1692);
xnor U1852 (N_1852,N_1741,N_1631);
and U1853 (N_1853,N_1708,N_1624);
nand U1854 (N_1854,N_1516,N_1509);
xor U1855 (N_1855,N_1550,N_1726);
and U1856 (N_1856,N_1625,N_1594);
xnor U1857 (N_1857,N_1518,N_1611);
nand U1858 (N_1858,N_1672,N_1528);
or U1859 (N_1859,N_1574,N_1520);
nor U1860 (N_1860,N_1705,N_1591);
or U1861 (N_1861,N_1689,N_1510);
nand U1862 (N_1862,N_1707,N_1648);
or U1863 (N_1863,N_1652,N_1740);
nor U1864 (N_1864,N_1608,N_1660);
xor U1865 (N_1865,N_1542,N_1500);
nand U1866 (N_1866,N_1536,N_1738);
or U1867 (N_1867,N_1728,N_1604);
and U1868 (N_1868,N_1673,N_1671);
xor U1869 (N_1869,N_1582,N_1703);
or U1870 (N_1870,N_1683,N_1531);
nor U1871 (N_1871,N_1702,N_1505);
nor U1872 (N_1872,N_1534,N_1637);
nand U1873 (N_1873,N_1723,N_1675);
nand U1874 (N_1874,N_1743,N_1661);
nor U1875 (N_1875,N_1550,N_1555);
or U1876 (N_1876,N_1535,N_1635);
and U1877 (N_1877,N_1651,N_1532);
xnor U1878 (N_1878,N_1725,N_1672);
or U1879 (N_1879,N_1714,N_1735);
nand U1880 (N_1880,N_1702,N_1606);
nand U1881 (N_1881,N_1577,N_1683);
nand U1882 (N_1882,N_1583,N_1627);
and U1883 (N_1883,N_1604,N_1503);
xnor U1884 (N_1884,N_1624,N_1706);
or U1885 (N_1885,N_1691,N_1664);
or U1886 (N_1886,N_1571,N_1615);
and U1887 (N_1887,N_1608,N_1726);
nor U1888 (N_1888,N_1592,N_1536);
xor U1889 (N_1889,N_1588,N_1662);
xnor U1890 (N_1890,N_1638,N_1719);
and U1891 (N_1891,N_1716,N_1651);
xor U1892 (N_1892,N_1633,N_1707);
nor U1893 (N_1893,N_1727,N_1503);
xor U1894 (N_1894,N_1740,N_1545);
xnor U1895 (N_1895,N_1623,N_1718);
and U1896 (N_1896,N_1580,N_1604);
or U1897 (N_1897,N_1504,N_1640);
and U1898 (N_1898,N_1525,N_1533);
nor U1899 (N_1899,N_1676,N_1747);
or U1900 (N_1900,N_1541,N_1688);
nand U1901 (N_1901,N_1605,N_1625);
or U1902 (N_1902,N_1506,N_1558);
nor U1903 (N_1903,N_1630,N_1568);
xnor U1904 (N_1904,N_1569,N_1607);
nand U1905 (N_1905,N_1588,N_1517);
nand U1906 (N_1906,N_1719,N_1746);
xnor U1907 (N_1907,N_1533,N_1587);
or U1908 (N_1908,N_1601,N_1722);
nor U1909 (N_1909,N_1625,N_1555);
nor U1910 (N_1910,N_1590,N_1663);
nand U1911 (N_1911,N_1662,N_1642);
and U1912 (N_1912,N_1740,N_1707);
nand U1913 (N_1913,N_1534,N_1669);
nor U1914 (N_1914,N_1617,N_1535);
nand U1915 (N_1915,N_1735,N_1531);
nor U1916 (N_1916,N_1534,N_1544);
nor U1917 (N_1917,N_1635,N_1703);
xnor U1918 (N_1918,N_1654,N_1547);
or U1919 (N_1919,N_1642,N_1547);
nand U1920 (N_1920,N_1506,N_1668);
nand U1921 (N_1921,N_1640,N_1611);
nand U1922 (N_1922,N_1583,N_1589);
nand U1923 (N_1923,N_1641,N_1691);
nor U1924 (N_1924,N_1736,N_1662);
nor U1925 (N_1925,N_1696,N_1687);
nand U1926 (N_1926,N_1730,N_1697);
nor U1927 (N_1927,N_1625,N_1745);
xnor U1928 (N_1928,N_1606,N_1734);
nand U1929 (N_1929,N_1632,N_1537);
nand U1930 (N_1930,N_1675,N_1607);
xor U1931 (N_1931,N_1702,N_1615);
xor U1932 (N_1932,N_1634,N_1607);
and U1933 (N_1933,N_1676,N_1728);
or U1934 (N_1934,N_1652,N_1660);
or U1935 (N_1935,N_1740,N_1605);
and U1936 (N_1936,N_1616,N_1570);
xnor U1937 (N_1937,N_1686,N_1575);
and U1938 (N_1938,N_1686,N_1717);
nand U1939 (N_1939,N_1733,N_1693);
nor U1940 (N_1940,N_1695,N_1577);
xor U1941 (N_1941,N_1589,N_1509);
or U1942 (N_1942,N_1635,N_1605);
nor U1943 (N_1943,N_1692,N_1530);
nor U1944 (N_1944,N_1540,N_1645);
xor U1945 (N_1945,N_1743,N_1600);
or U1946 (N_1946,N_1714,N_1556);
xnor U1947 (N_1947,N_1547,N_1687);
xnor U1948 (N_1948,N_1650,N_1554);
nand U1949 (N_1949,N_1627,N_1727);
and U1950 (N_1950,N_1667,N_1527);
nand U1951 (N_1951,N_1633,N_1713);
xor U1952 (N_1952,N_1666,N_1668);
nor U1953 (N_1953,N_1564,N_1667);
xnor U1954 (N_1954,N_1743,N_1539);
xnor U1955 (N_1955,N_1617,N_1674);
nor U1956 (N_1956,N_1691,N_1698);
and U1957 (N_1957,N_1709,N_1733);
nor U1958 (N_1958,N_1693,N_1520);
nand U1959 (N_1959,N_1729,N_1668);
nand U1960 (N_1960,N_1647,N_1551);
nand U1961 (N_1961,N_1679,N_1586);
nor U1962 (N_1962,N_1607,N_1576);
nand U1963 (N_1963,N_1550,N_1611);
nor U1964 (N_1964,N_1570,N_1608);
xor U1965 (N_1965,N_1678,N_1527);
xnor U1966 (N_1966,N_1577,N_1631);
or U1967 (N_1967,N_1525,N_1673);
nand U1968 (N_1968,N_1526,N_1704);
nand U1969 (N_1969,N_1625,N_1548);
or U1970 (N_1970,N_1638,N_1712);
or U1971 (N_1971,N_1529,N_1653);
nand U1972 (N_1972,N_1530,N_1596);
or U1973 (N_1973,N_1721,N_1560);
xor U1974 (N_1974,N_1530,N_1502);
or U1975 (N_1975,N_1642,N_1747);
nand U1976 (N_1976,N_1696,N_1544);
and U1977 (N_1977,N_1723,N_1612);
and U1978 (N_1978,N_1649,N_1609);
and U1979 (N_1979,N_1734,N_1624);
nand U1980 (N_1980,N_1664,N_1575);
xnor U1981 (N_1981,N_1523,N_1728);
and U1982 (N_1982,N_1581,N_1511);
nor U1983 (N_1983,N_1553,N_1651);
and U1984 (N_1984,N_1553,N_1534);
nand U1985 (N_1985,N_1640,N_1741);
and U1986 (N_1986,N_1510,N_1610);
and U1987 (N_1987,N_1509,N_1576);
or U1988 (N_1988,N_1531,N_1639);
xor U1989 (N_1989,N_1632,N_1713);
nor U1990 (N_1990,N_1644,N_1678);
or U1991 (N_1991,N_1543,N_1628);
xor U1992 (N_1992,N_1519,N_1594);
nand U1993 (N_1993,N_1735,N_1509);
xor U1994 (N_1994,N_1670,N_1624);
or U1995 (N_1995,N_1730,N_1602);
xor U1996 (N_1996,N_1698,N_1732);
or U1997 (N_1997,N_1735,N_1629);
and U1998 (N_1998,N_1672,N_1628);
xnor U1999 (N_1999,N_1597,N_1737);
and U2000 (N_2000,N_1904,N_1828);
nand U2001 (N_2001,N_1906,N_1805);
or U2002 (N_2002,N_1974,N_1775);
nor U2003 (N_2003,N_1884,N_1953);
nor U2004 (N_2004,N_1773,N_1881);
and U2005 (N_2005,N_1858,N_1809);
nor U2006 (N_2006,N_1945,N_1813);
or U2007 (N_2007,N_1819,N_1928);
xor U2008 (N_2008,N_1804,N_1783);
xnor U2009 (N_2009,N_1888,N_1873);
nand U2010 (N_2010,N_1855,N_1808);
or U2011 (N_2011,N_1810,N_1815);
nor U2012 (N_2012,N_1817,N_1982);
nor U2013 (N_2013,N_1753,N_1867);
xor U2014 (N_2014,N_1957,N_1921);
nor U2015 (N_2015,N_1859,N_1849);
and U2016 (N_2016,N_1781,N_1825);
and U2017 (N_2017,N_1779,N_1983);
or U2018 (N_2018,N_1768,N_1896);
or U2019 (N_2019,N_1919,N_1901);
nand U2020 (N_2020,N_1834,N_1790);
nand U2021 (N_2021,N_1822,N_1940);
nand U2022 (N_2022,N_1878,N_1898);
or U2023 (N_2023,N_1777,N_1767);
and U2024 (N_2024,N_1992,N_1948);
nand U2025 (N_2025,N_1946,N_1934);
xnor U2026 (N_2026,N_1869,N_1877);
nor U2027 (N_2027,N_1915,N_1831);
nor U2028 (N_2028,N_1792,N_1991);
xnor U2029 (N_2029,N_1923,N_1968);
nand U2030 (N_2030,N_1864,N_1903);
or U2031 (N_2031,N_1848,N_1750);
or U2032 (N_2032,N_1821,N_1835);
and U2033 (N_2033,N_1861,N_1761);
or U2034 (N_2034,N_1943,N_1846);
nand U2035 (N_2035,N_1944,N_1863);
nand U2036 (N_2036,N_1889,N_1971);
and U2037 (N_2037,N_1987,N_1988);
or U2038 (N_2038,N_1841,N_1771);
xor U2039 (N_2039,N_1796,N_1969);
xor U2040 (N_2040,N_1832,N_1905);
or U2041 (N_2041,N_1812,N_1997);
or U2042 (N_2042,N_1998,N_1980);
nor U2043 (N_2043,N_1801,N_1978);
xnor U2044 (N_2044,N_1788,N_1836);
nand U2045 (N_2045,N_1875,N_1897);
nand U2046 (N_2046,N_1938,N_1840);
and U2047 (N_2047,N_1927,N_1918);
and U2048 (N_2048,N_1929,N_1935);
nand U2049 (N_2049,N_1757,N_1981);
nand U2050 (N_2050,N_1937,N_1760);
nand U2051 (N_2051,N_1764,N_1965);
xnor U2052 (N_2052,N_1860,N_1885);
or U2053 (N_2053,N_1914,N_1870);
nor U2054 (N_2054,N_1778,N_1823);
or U2055 (N_2055,N_1887,N_1789);
or U2056 (N_2056,N_1772,N_1993);
nand U2057 (N_2057,N_1916,N_1833);
nand U2058 (N_2058,N_1871,N_1984);
nor U2059 (N_2059,N_1883,N_1795);
or U2060 (N_2060,N_1932,N_1924);
nand U2061 (N_2061,N_1895,N_1824);
nor U2062 (N_2062,N_1798,N_1926);
or U2063 (N_2063,N_1985,N_1942);
or U2064 (N_2064,N_1791,N_1838);
or U2065 (N_2065,N_1959,N_1892);
xnor U2066 (N_2066,N_1752,N_1842);
nor U2067 (N_2067,N_1759,N_1862);
and U2068 (N_2068,N_1852,N_1908);
or U2069 (N_2069,N_1879,N_1837);
xor U2070 (N_2070,N_1939,N_1976);
xor U2071 (N_2071,N_1853,N_1977);
nand U2072 (N_2072,N_1956,N_1784);
and U2073 (N_2073,N_1845,N_1811);
and U2074 (N_2074,N_1814,N_1962);
nand U2075 (N_2075,N_1787,N_1893);
or U2076 (N_2076,N_1806,N_1900);
xnor U2077 (N_2077,N_1803,N_1961);
nand U2078 (N_2078,N_1886,N_1816);
and U2079 (N_2079,N_1949,N_1912);
xnor U2080 (N_2080,N_1996,N_1973);
xnor U2081 (N_2081,N_1882,N_1909);
xor U2082 (N_2082,N_1979,N_1989);
or U2083 (N_2083,N_1910,N_1990);
nor U2084 (N_2084,N_1765,N_1960);
xor U2085 (N_2085,N_1865,N_1899);
nor U2086 (N_2086,N_1933,N_1820);
nor U2087 (N_2087,N_1890,N_1955);
xnor U2088 (N_2088,N_1894,N_1913);
nand U2089 (N_2089,N_1970,N_1839);
nand U2090 (N_2090,N_1756,N_1950);
and U2091 (N_2091,N_1876,N_1826);
and U2092 (N_2092,N_1850,N_1774);
or U2093 (N_2093,N_1800,N_1770);
xnor U2094 (N_2094,N_1818,N_1995);
and U2095 (N_2095,N_1902,N_1958);
xnor U2096 (N_2096,N_1755,N_1751);
and U2097 (N_2097,N_1793,N_1936);
nor U2098 (N_2098,N_1964,N_1930);
and U2099 (N_2099,N_1941,N_1925);
nand U2100 (N_2100,N_1857,N_1769);
nor U2101 (N_2101,N_1843,N_1847);
and U2102 (N_2102,N_1766,N_1854);
or U2103 (N_2103,N_1880,N_1844);
xnor U2104 (N_2104,N_1797,N_1907);
xor U2105 (N_2105,N_1782,N_1799);
and U2106 (N_2106,N_1866,N_1872);
xor U2107 (N_2107,N_1952,N_1966);
xor U2108 (N_2108,N_1830,N_1911);
nor U2109 (N_2109,N_1776,N_1999);
nor U2110 (N_2110,N_1786,N_1917);
or U2111 (N_2111,N_1754,N_1972);
nor U2112 (N_2112,N_1975,N_1931);
and U2113 (N_2113,N_1851,N_1794);
nand U2114 (N_2114,N_1802,N_1986);
and U2115 (N_2115,N_1829,N_1954);
or U2116 (N_2116,N_1994,N_1758);
or U2117 (N_2117,N_1920,N_1947);
xnor U2118 (N_2118,N_1780,N_1763);
and U2119 (N_2119,N_1785,N_1762);
xnor U2120 (N_2120,N_1868,N_1891);
nor U2121 (N_2121,N_1827,N_1807);
nand U2122 (N_2122,N_1874,N_1951);
nand U2123 (N_2123,N_1967,N_1922);
xor U2124 (N_2124,N_1963,N_1856);
nand U2125 (N_2125,N_1853,N_1979);
and U2126 (N_2126,N_1988,N_1985);
nor U2127 (N_2127,N_1932,N_1972);
nand U2128 (N_2128,N_1997,N_1898);
nand U2129 (N_2129,N_1931,N_1835);
nand U2130 (N_2130,N_1948,N_1894);
xor U2131 (N_2131,N_1986,N_1967);
nor U2132 (N_2132,N_1970,N_1855);
nand U2133 (N_2133,N_1946,N_1906);
nand U2134 (N_2134,N_1910,N_1950);
nand U2135 (N_2135,N_1752,N_1844);
nor U2136 (N_2136,N_1996,N_1759);
and U2137 (N_2137,N_1877,N_1898);
or U2138 (N_2138,N_1779,N_1881);
or U2139 (N_2139,N_1860,N_1876);
nor U2140 (N_2140,N_1995,N_1783);
or U2141 (N_2141,N_1959,N_1870);
nand U2142 (N_2142,N_1755,N_1924);
xnor U2143 (N_2143,N_1810,N_1788);
or U2144 (N_2144,N_1860,N_1803);
nand U2145 (N_2145,N_1841,N_1899);
nand U2146 (N_2146,N_1894,N_1781);
xor U2147 (N_2147,N_1810,N_1806);
or U2148 (N_2148,N_1808,N_1834);
nor U2149 (N_2149,N_1892,N_1868);
xor U2150 (N_2150,N_1823,N_1905);
nor U2151 (N_2151,N_1866,N_1877);
nor U2152 (N_2152,N_1942,N_1951);
nor U2153 (N_2153,N_1915,N_1951);
or U2154 (N_2154,N_1945,N_1834);
xor U2155 (N_2155,N_1881,N_1989);
xnor U2156 (N_2156,N_1795,N_1838);
nand U2157 (N_2157,N_1892,N_1831);
or U2158 (N_2158,N_1831,N_1821);
xnor U2159 (N_2159,N_1833,N_1872);
nand U2160 (N_2160,N_1962,N_1825);
and U2161 (N_2161,N_1772,N_1868);
or U2162 (N_2162,N_1993,N_1805);
or U2163 (N_2163,N_1750,N_1898);
nor U2164 (N_2164,N_1831,N_1779);
nand U2165 (N_2165,N_1809,N_1844);
and U2166 (N_2166,N_1896,N_1991);
nor U2167 (N_2167,N_1811,N_1899);
and U2168 (N_2168,N_1932,N_1896);
nand U2169 (N_2169,N_1804,N_1779);
or U2170 (N_2170,N_1799,N_1981);
and U2171 (N_2171,N_1955,N_1848);
and U2172 (N_2172,N_1935,N_1820);
and U2173 (N_2173,N_1959,N_1797);
xnor U2174 (N_2174,N_1940,N_1800);
xor U2175 (N_2175,N_1924,N_1818);
nand U2176 (N_2176,N_1889,N_1750);
nor U2177 (N_2177,N_1977,N_1952);
nand U2178 (N_2178,N_1861,N_1752);
nand U2179 (N_2179,N_1983,N_1956);
and U2180 (N_2180,N_1781,N_1990);
nand U2181 (N_2181,N_1952,N_1793);
xnor U2182 (N_2182,N_1860,N_1957);
or U2183 (N_2183,N_1811,N_1937);
nor U2184 (N_2184,N_1965,N_1928);
xnor U2185 (N_2185,N_1935,N_1960);
nor U2186 (N_2186,N_1846,N_1783);
nand U2187 (N_2187,N_1788,N_1960);
nor U2188 (N_2188,N_1940,N_1876);
xnor U2189 (N_2189,N_1883,N_1910);
or U2190 (N_2190,N_1803,N_1989);
or U2191 (N_2191,N_1977,N_1901);
xnor U2192 (N_2192,N_1825,N_1815);
nor U2193 (N_2193,N_1917,N_1880);
nor U2194 (N_2194,N_1753,N_1824);
nand U2195 (N_2195,N_1825,N_1793);
nor U2196 (N_2196,N_1802,N_1998);
and U2197 (N_2197,N_1966,N_1933);
nand U2198 (N_2198,N_1819,N_1846);
xnor U2199 (N_2199,N_1775,N_1902);
xnor U2200 (N_2200,N_1810,N_1960);
nor U2201 (N_2201,N_1914,N_1920);
or U2202 (N_2202,N_1967,N_1993);
nand U2203 (N_2203,N_1822,N_1807);
nand U2204 (N_2204,N_1895,N_1922);
nand U2205 (N_2205,N_1754,N_1996);
or U2206 (N_2206,N_1991,N_1941);
and U2207 (N_2207,N_1895,N_1764);
and U2208 (N_2208,N_1805,N_1784);
and U2209 (N_2209,N_1888,N_1778);
nand U2210 (N_2210,N_1904,N_1846);
nand U2211 (N_2211,N_1942,N_1967);
or U2212 (N_2212,N_1978,N_1974);
xor U2213 (N_2213,N_1918,N_1834);
and U2214 (N_2214,N_1834,N_1890);
xnor U2215 (N_2215,N_1948,N_1752);
and U2216 (N_2216,N_1950,N_1996);
nor U2217 (N_2217,N_1956,N_1962);
or U2218 (N_2218,N_1795,N_1907);
nor U2219 (N_2219,N_1987,N_1873);
xnor U2220 (N_2220,N_1978,N_1921);
and U2221 (N_2221,N_1795,N_1915);
nor U2222 (N_2222,N_1938,N_1829);
nand U2223 (N_2223,N_1975,N_1771);
and U2224 (N_2224,N_1847,N_1842);
xnor U2225 (N_2225,N_1754,N_1898);
xor U2226 (N_2226,N_1832,N_1975);
nor U2227 (N_2227,N_1937,N_1775);
or U2228 (N_2228,N_1978,N_1920);
xor U2229 (N_2229,N_1893,N_1979);
xnor U2230 (N_2230,N_1757,N_1884);
nor U2231 (N_2231,N_1985,N_1838);
and U2232 (N_2232,N_1779,N_1815);
or U2233 (N_2233,N_1957,N_1996);
and U2234 (N_2234,N_1949,N_1930);
nand U2235 (N_2235,N_1777,N_1917);
nand U2236 (N_2236,N_1943,N_1955);
or U2237 (N_2237,N_1988,N_1813);
xnor U2238 (N_2238,N_1965,N_1840);
or U2239 (N_2239,N_1808,N_1967);
or U2240 (N_2240,N_1766,N_1934);
and U2241 (N_2241,N_1831,N_1903);
nand U2242 (N_2242,N_1982,N_1828);
nor U2243 (N_2243,N_1893,N_1938);
or U2244 (N_2244,N_1829,N_1909);
or U2245 (N_2245,N_1792,N_1757);
xor U2246 (N_2246,N_1789,N_1938);
or U2247 (N_2247,N_1893,N_1983);
or U2248 (N_2248,N_1764,N_1802);
and U2249 (N_2249,N_1947,N_1834);
xor U2250 (N_2250,N_2248,N_2062);
nand U2251 (N_2251,N_2149,N_2217);
and U2252 (N_2252,N_2061,N_2159);
or U2253 (N_2253,N_2028,N_2016);
and U2254 (N_2254,N_2026,N_2229);
nor U2255 (N_2255,N_2010,N_2204);
nand U2256 (N_2256,N_2102,N_2019);
xnor U2257 (N_2257,N_2111,N_2041);
nor U2258 (N_2258,N_2169,N_2063);
nor U2259 (N_2259,N_2209,N_2178);
and U2260 (N_2260,N_2237,N_2116);
and U2261 (N_2261,N_2068,N_2048);
and U2262 (N_2262,N_2230,N_2094);
nand U2263 (N_2263,N_2153,N_2191);
nor U2264 (N_2264,N_2206,N_2152);
nand U2265 (N_2265,N_2140,N_2012);
xnor U2266 (N_2266,N_2138,N_2042);
xnor U2267 (N_2267,N_2188,N_2080);
nor U2268 (N_2268,N_2056,N_2037);
xnor U2269 (N_2269,N_2090,N_2238);
nor U2270 (N_2270,N_2077,N_2194);
and U2271 (N_2271,N_2113,N_2122);
and U2272 (N_2272,N_2129,N_2211);
xnor U2273 (N_2273,N_2239,N_2166);
xnor U2274 (N_2274,N_2224,N_2155);
xor U2275 (N_2275,N_2084,N_2137);
or U2276 (N_2276,N_2228,N_2045);
and U2277 (N_2277,N_2064,N_2024);
nand U2278 (N_2278,N_2076,N_2114);
or U2279 (N_2279,N_2190,N_2157);
or U2280 (N_2280,N_2241,N_2003);
and U2281 (N_2281,N_2220,N_2074);
or U2282 (N_2282,N_2099,N_2156);
nor U2283 (N_2283,N_2004,N_2146);
nor U2284 (N_2284,N_2070,N_2179);
nor U2285 (N_2285,N_2069,N_2222);
nand U2286 (N_2286,N_2075,N_2040);
xor U2287 (N_2287,N_2225,N_2135);
and U2288 (N_2288,N_2242,N_2203);
xnor U2289 (N_2289,N_2072,N_2215);
nor U2290 (N_2290,N_2196,N_2112);
nand U2291 (N_2291,N_2066,N_2086);
xnor U2292 (N_2292,N_2134,N_2243);
xor U2293 (N_2293,N_2036,N_2044);
nor U2294 (N_2294,N_2001,N_2124);
or U2295 (N_2295,N_2088,N_2136);
or U2296 (N_2296,N_2052,N_2235);
nor U2297 (N_2297,N_2150,N_2067);
or U2298 (N_2298,N_2121,N_2180);
nor U2299 (N_2299,N_2207,N_2192);
nand U2300 (N_2300,N_2198,N_2148);
nand U2301 (N_2301,N_2014,N_2210);
and U2302 (N_2302,N_2038,N_2212);
and U2303 (N_2303,N_2171,N_2170);
and U2304 (N_2304,N_2175,N_2050);
nor U2305 (N_2305,N_2234,N_2176);
nand U2306 (N_2306,N_2087,N_2115);
xor U2307 (N_2307,N_2034,N_2128);
nor U2308 (N_2308,N_2089,N_2177);
or U2309 (N_2309,N_2083,N_2033);
or U2310 (N_2310,N_2218,N_2123);
xnor U2311 (N_2311,N_2002,N_2055);
and U2312 (N_2312,N_2018,N_2201);
nand U2313 (N_2313,N_2199,N_2236);
xor U2314 (N_2314,N_2017,N_2223);
nor U2315 (N_2315,N_2232,N_2096);
nand U2316 (N_2316,N_2189,N_2151);
and U2317 (N_2317,N_2058,N_2132);
nand U2318 (N_2318,N_2130,N_2008);
nor U2319 (N_2319,N_2214,N_2163);
or U2320 (N_2320,N_2082,N_2208);
nand U2321 (N_2321,N_2244,N_2143);
nand U2322 (N_2322,N_2039,N_2221);
xnor U2323 (N_2323,N_2073,N_2095);
and U2324 (N_2324,N_2186,N_2158);
and U2325 (N_2325,N_2059,N_2162);
or U2326 (N_2326,N_2043,N_2168);
nand U2327 (N_2327,N_2184,N_2197);
nor U2328 (N_2328,N_2110,N_2107);
xnor U2329 (N_2329,N_2200,N_2249);
or U2330 (N_2330,N_2023,N_2022);
nand U2331 (N_2331,N_2020,N_2097);
and U2332 (N_2332,N_2098,N_2185);
or U2333 (N_2333,N_2009,N_2007);
or U2334 (N_2334,N_2051,N_2182);
or U2335 (N_2335,N_2144,N_2226);
nand U2336 (N_2336,N_2120,N_2101);
and U2337 (N_2337,N_2131,N_2142);
or U2338 (N_2338,N_2127,N_2047);
nor U2339 (N_2339,N_2032,N_2118);
nand U2340 (N_2340,N_2161,N_2181);
or U2341 (N_2341,N_2029,N_2005);
nor U2342 (N_2342,N_2233,N_2213);
xnor U2343 (N_2343,N_2015,N_2100);
nor U2344 (N_2344,N_2108,N_2006);
or U2345 (N_2345,N_2035,N_2054);
or U2346 (N_2346,N_2000,N_2147);
nor U2347 (N_2347,N_2245,N_2046);
xor U2348 (N_2348,N_2104,N_2173);
nand U2349 (N_2349,N_2172,N_2078);
or U2350 (N_2350,N_2011,N_2091);
or U2351 (N_2351,N_2139,N_2030);
or U2352 (N_2352,N_2227,N_2085);
nor U2353 (N_2353,N_2246,N_2065);
or U2354 (N_2354,N_2092,N_2216);
xnor U2355 (N_2355,N_2202,N_2125);
and U2356 (N_2356,N_2071,N_2013);
or U2357 (N_2357,N_2154,N_2079);
or U2358 (N_2358,N_2145,N_2081);
or U2359 (N_2359,N_2106,N_2053);
and U2360 (N_2360,N_2193,N_2183);
nor U2361 (N_2361,N_2049,N_2025);
or U2362 (N_2362,N_2105,N_2195);
or U2363 (N_2363,N_2117,N_2093);
nand U2364 (N_2364,N_2021,N_2060);
and U2365 (N_2365,N_2126,N_2247);
nor U2366 (N_2366,N_2219,N_2164);
xnor U2367 (N_2367,N_2231,N_2109);
or U2368 (N_2368,N_2174,N_2057);
xnor U2369 (N_2369,N_2167,N_2160);
nor U2370 (N_2370,N_2165,N_2133);
nor U2371 (N_2371,N_2240,N_2031);
xnor U2372 (N_2372,N_2119,N_2187);
nor U2373 (N_2373,N_2103,N_2141);
nand U2374 (N_2374,N_2205,N_2027);
nand U2375 (N_2375,N_2138,N_2202);
and U2376 (N_2376,N_2088,N_2214);
nor U2377 (N_2377,N_2029,N_2089);
xnor U2378 (N_2378,N_2077,N_2146);
nand U2379 (N_2379,N_2092,N_2066);
or U2380 (N_2380,N_2042,N_2227);
nor U2381 (N_2381,N_2212,N_2166);
or U2382 (N_2382,N_2056,N_2101);
or U2383 (N_2383,N_2205,N_2076);
and U2384 (N_2384,N_2215,N_2071);
nand U2385 (N_2385,N_2039,N_2085);
and U2386 (N_2386,N_2205,N_2125);
nor U2387 (N_2387,N_2225,N_2037);
nor U2388 (N_2388,N_2234,N_2160);
and U2389 (N_2389,N_2093,N_2208);
xnor U2390 (N_2390,N_2001,N_2156);
and U2391 (N_2391,N_2094,N_2163);
and U2392 (N_2392,N_2143,N_2198);
nand U2393 (N_2393,N_2164,N_2109);
nor U2394 (N_2394,N_2228,N_2150);
xnor U2395 (N_2395,N_2161,N_2091);
xnor U2396 (N_2396,N_2085,N_2199);
and U2397 (N_2397,N_2236,N_2066);
xnor U2398 (N_2398,N_2113,N_2001);
nor U2399 (N_2399,N_2091,N_2215);
nand U2400 (N_2400,N_2105,N_2139);
or U2401 (N_2401,N_2142,N_2079);
nand U2402 (N_2402,N_2164,N_2007);
and U2403 (N_2403,N_2022,N_2052);
or U2404 (N_2404,N_2137,N_2224);
and U2405 (N_2405,N_2169,N_2030);
and U2406 (N_2406,N_2151,N_2081);
and U2407 (N_2407,N_2092,N_2005);
nor U2408 (N_2408,N_2159,N_2202);
and U2409 (N_2409,N_2226,N_2036);
nor U2410 (N_2410,N_2192,N_2170);
nor U2411 (N_2411,N_2109,N_2206);
nor U2412 (N_2412,N_2167,N_2202);
or U2413 (N_2413,N_2229,N_2089);
xnor U2414 (N_2414,N_2237,N_2000);
nor U2415 (N_2415,N_2150,N_2024);
and U2416 (N_2416,N_2191,N_2209);
or U2417 (N_2417,N_2003,N_2246);
xnor U2418 (N_2418,N_2090,N_2172);
nor U2419 (N_2419,N_2082,N_2004);
xnor U2420 (N_2420,N_2004,N_2236);
nor U2421 (N_2421,N_2081,N_2057);
nor U2422 (N_2422,N_2196,N_2055);
nor U2423 (N_2423,N_2214,N_2239);
nand U2424 (N_2424,N_2088,N_2055);
and U2425 (N_2425,N_2225,N_2053);
nor U2426 (N_2426,N_2199,N_2164);
xor U2427 (N_2427,N_2214,N_2153);
xor U2428 (N_2428,N_2037,N_2189);
nor U2429 (N_2429,N_2230,N_2105);
nor U2430 (N_2430,N_2178,N_2084);
and U2431 (N_2431,N_2039,N_2016);
nor U2432 (N_2432,N_2039,N_2044);
and U2433 (N_2433,N_2191,N_2212);
nor U2434 (N_2434,N_2175,N_2173);
nand U2435 (N_2435,N_2067,N_2176);
nand U2436 (N_2436,N_2004,N_2140);
nand U2437 (N_2437,N_2097,N_2092);
nand U2438 (N_2438,N_2160,N_2060);
or U2439 (N_2439,N_2177,N_2094);
xor U2440 (N_2440,N_2209,N_2005);
xnor U2441 (N_2441,N_2014,N_2013);
or U2442 (N_2442,N_2016,N_2122);
xor U2443 (N_2443,N_2152,N_2243);
or U2444 (N_2444,N_2229,N_2186);
nand U2445 (N_2445,N_2081,N_2193);
nand U2446 (N_2446,N_2158,N_2066);
or U2447 (N_2447,N_2038,N_2006);
xor U2448 (N_2448,N_2147,N_2191);
xor U2449 (N_2449,N_2053,N_2056);
nor U2450 (N_2450,N_2151,N_2197);
xnor U2451 (N_2451,N_2047,N_2066);
or U2452 (N_2452,N_2202,N_2086);
xnor U2453 (N_2453,N_2133,N_2036);
nand U2454 (N_2454,N_2002,N_2147);
or U2455 (N_2455,N_2130,N_2114);
or U2456 (N_2456,N_2011,N_2049);
xor U2457 (N_2457,N_2086,N_2112);
or U2458 (N_2458,N_2200,N_2120);
and U2459 (N_2459,N_2005,N_2246);
nand U2460 (N_2460,N_2163,N_2111);
and U2461 (N_2461,N_2000,N_2001);
xor U2462 (N_2462,N_2088,N_2020);
nor U2463 (N_2463,N_2237,N_2103);
nand U2464 (N_2464,N_2021,N_2141);
nor U2465 (N_2465,N_2007,N_2117);
and U2466 (N_2466,N_2229,N_2014);
or U2467 (N_2467,N_2108,N_2078);
nand U2468 (N_2468,N_2190,N_2230);
or U2469 (N_2469,N_2183,N_2097);
nor U2470 (N_2470,N_2249,N_2130);
nor U2471 (N_2471,N_2096,N_2073);
or U2472 (N_2472,N_2143,N_2025);
xor U2473 (N_2473,N_2027,N_2066);
nor U2474 (N_2474,N_2157,N_2033);
and U2475 (N_2475,N_2093,N_2231);
nor U2476 (N_2476,N_2077,N_2094);
nor U2477 (N_2477,N_2239,N_2085);
xor U2478 (N_2478,N_2154,N_2205);
nand U2479 (N_2479,N_2215,N_2010);
nand U2480 (N_2480,N_2228,N_2018);
nor U2481 (N_2481,N_2249,N_2067);
or U2482 (N_2482,N_2190,N_2160);
nand U2483 (N_2483,N_2076,N_2236);
xor U2484 (N_2484,N_2191,N_2077);
or U2485 (N_2485,N_2214,N_2137);
nand U2486 (N_2486,N_2078,N_2161);
nor U2487 (N_2487,N_2140,N_2022);
nand U2488 (N_2488,N_2179,N_2196);
and U2489 (N_2489,N_2234,N_2142);
and U2490 (N_2490,N_2049,N_2143);
or U2491 (N_2491,N_2246,N_2205);
and U2492 (N_2492,N_2208,N_2142);
xor U2493 (N_2493,N_2005,N_2098);
xor U2494 (N_2494,N_2059,N_2008);
nand U2495 (N_2495,N_2106,N_2060);
nand U2496 (N_2496,N_2182,N_2054);
or U2497 (N_2497,N_2106,N_2006);
and U2498 (N_2498,N_2058,N_2144);
nor U2499 (N_2499,N_2189,N_2095);
nor U2500 (N_2500,N_2428,N_2433);
and U2501 (N_2501,N_2486,N_2467);
or U2502 (N_2502,N_2445,N_2479);
nor U2503 (N_2503,N_2458,N_2348);
nor U2504 (N_2504,N_2455,N_2372);
nand U2505 (N_2505,N_2318,N_2463);
and U2506 (N_2506,N_2459,N_2304);
nor U2507 (N_2507,N_2332,N_2277);
and U2508 (N_2508,N_2404,N_2361);
or U2509 (N_2509,N_2424,N_2383);
and U2510 (N_2510,N_2268,N_2476);
nor U2511 (N_2511,N_2466,N_2346);
and U2512 (N_2512,N_2315,N_2490);
nor U2513 (N_2513,N_2289,N_2425);
nor U2514 (N_2514,N_2392,N_2331);
xor U2515 (N_2515,N_2473,N_2498);
xor U2516 (N_2516,N_2307,N_2482);
nand U2517 (N_2517,N_2415,N_2265);
nand U2518 (N_2518,N_2366,N_2300);
nand U2519 (N_2519,N_2485,N_2396);
or U2520 (N_2520,N_2439,N_2382);
or U2521 (N_2521,N_2395,N_2481);
xor U2522 (N_2522,N_2368,N_2355);
xnor U2523 (N_2523,N_2278,N_2305);
nor U2524 (N_2524,N_2369,N_2436);
nor U2525 (N_2525,N_2281,N_2334);
xnor U2526 (N_2526,N_2344,N_2312);
and U2527 (N_2527,N_2260,N_2356);
or U2528 (N_2528,N_2343,N_2388);
nor U2529 (N_2529,N_2474,N_2447);
xor U2530 (N_2530,N_2352,N_2462);
nand U2531 (N_2531,N_2386,N_2333);
or U2532 (N_2532,N_2391,N_2350);
xor U2533 (N_2533,N_2370,N_2435);
nand U2534 (N_2534,N_2470,N_2446);
or U2535 (N_2535,N_2469,N_2314);
and U2536 (N_2536,N_2283,N_2279);
or U2537 (N_2537,N_2253,N_2472);
nand U2538 (N_2538,N_2270,N_2359);
nand U2539 (N_2539,N_2398,N_2257);
and U2540 (N_2540,N_2256,N_2387);
nor U2541 (N_2541,N_2339,N_2464);
and U2542 (N_2542,N_2454,N_2293);
nand U2543 (N_2543,N_2258,N_2407);
nor U2544 (N_2544,N_2456,N_2313);
nand U2545 (N_2545,N_2403,N_2401);
nand U2546 (N_2546,N_2326,N_2471);
nor U2547 (N_2547,N_2271,N_2274);
xnor U2548 (N_2548,N_2477,N_2457);
and U2549 (N_2549,N_2319,N_2328);
nand U2550 (N_2550,N_2438,N_2309);
xnor U2551 (N_2551,N_2374,N_2418);
nor U2552 (N_2552,N_2347,N_2285);
nand U2553 (N_2553,N_2384,N_2295);
xor U2554 (N_2554,N_2365,N_2272);
nor U2555 (N_2555,N_2488,N_2349);
nand U2556 (N_2556,N_2302,N_2414);
xor U2557 (N_2557,N_2310,N_2335);
or U2558 (N_2558,N_2451,N_2341);
and U2559 (N_2559,N_2294,N_2354);
nor U2560 (N_2560,N_2440,N_2437);
or U2561 (N_2561,N_2377,N_2389);
nand U2562 (N_2562,N_2376,N_2429);
xor U2563 (N_2563,N_2252,N_2322);
nor U2564 (N_2564,N_2373,N_2410);
or U2565 (N_2565,N_2450,N_2323);
or U2566 (N_2566,N_2416,N_2351);
nand U2567 (N_2567,N_2284,N_2460);
nor U2568 (N_2568,N_2495,N_2259);
nor U2569 (N_2569,N_2282,N_2303);
xnor U2570 (N_2570,N_2321,N_2385);
or U2571 (N_2571,N_2492,N_2381);
nand U2572 (N_2572,N_2299,N_2306);
nor U2573 (N_2573,N_2426,N_2399);
or U2574 (N_2574,N_2327,N_2308);
or U2575 (N_2575,N_2262,N_2276);
or U2576 (N_2576,N_2380,N_2263);
xor U2577 (N_2577,N_2417,N_2291);
nor U2578 (N_2578,N_2441,N_2296);
nand U2579 (N_2579,N_2421,N_2367);
xor U2580 (N_2580,N_2340,N_2409);
and U2581 (N_2581,N_2408,N_2342);
xnor U2582 (N_2582,N_2432,N_2362);
nor U2583 (N_2583,N_2280,N_2419);
xor U2584 (N_2584,N_2267,N_2336);
nor U2585 (N_2585,N_2444,N_2468);
or U2586 (N_2586,N_2375,N_2483);
and U2587 (N_2587,N_2412,N_2378);
nand U2588 (N_2588,N_2329,N_2431);
nand U2589 (N_2589,N_2478,N_2453);
and U2590 (N_2590,N_2255,N_2434);
or U2591 (N_2591,N_2449,N_2484);
nand U2592 (N_2592,N_2406,N_2400);
nor U2593 (N_2593,N_2371,N_2496);
xnor U2594 (N_2594,N_2250,N_2413);
xnor U2595 (N_2595,N_2266,N_2423);
nand U2596 (N_2596,N_2487,N_2287);
xor U2597 (N_2597,N_2442,N_2489);
and U2598 (N_2598,N_2325,N_2324);
and U2599 (N_2599,N_2288,N_2499);
xnor U2600 (N_2600,N_2298,N_2364);
nand U2601 (N_2601,N_2358,N_2452);
and U2602 (N_2602,N_2269,N_2337);
and U2603 (N_2603,N_2390,N_2493);
and U2604 (N_2604,N_2254,N_2402);
or U2605 (N_2605,N_2461,N_2311);
xor U2606 (N_2606,N_2301,N_2363);
nand U2607 (N_2607,N_2420,N_2397);
nand U2608 (N_2608,N_2465,N_2345);
nor U2609 (N_2609,N_2394,N_2261);
nor U2610 (N_2610,N_2443,N_2491);
and U2611 (N_2611,N_2338,N_2422);
nand U2612 (N_2612,N_2427,N_2497);
xnor U2613 (N_2613,N_2448,N_2251);
or U2614 (N_2614,N_2273,N_2292);
xor U2615 (N_2615,N_2480,N_2393);
or U2616 (N_2616,N_2286,N_2475);
xor U2617 (N_2617,N_2330,N_2317);
or U2618 (N_2618,N_2494,N_2357);
nand U2619 (N_2619,N_2264,N_2320);
or U2620 (N_2620,N_2379,N_2275);
and U2621 (N_2621,N_2353,N_2360);
or U2622 (N_2622,N_2316,N_2297);
and U2623 (N_2623,N_2411,N_2430);
or U2624 (N_2624,N_2405,N_2290);
nor U2625 (N_2625,N_2479,N_2293);
and U2626 (N_2626,N_2300,N_2385);
xnor U2627 (N_2627,N_2280,N_2349);
and U2628 (N_2628,N_2305,N_2395);
nor U2629 (N_2629,N_2273,N_2441);
or U2630 (N_2630,N_2353,N_2419);
nor U2631 (N_2631,N_2268,N_2260);
nand U2632 (N_2632,N_2278,N_2259);
nor U2633 (N_2633,N_2406,N_2426);
xnor U2634 (N_2634,N_2471,N_2372);
or U2635 (N_2635,N_2423,N_2289);
or U2636 (N_2636,N_2407,N_2490);
xnor U2637 (N_2637,N_2439,N_2498);
or U2638 (N_2638,N_2380,N_2428);
nor U2639 (N_2639,N_2350,N_2463);
nand U2640 (N_2640,N_2462,N_2399);
or U2641 (N_2641,N_2469,N_2308);
xnor U2642 (N_2642,N_2366,N_2364);
nor U2643 (N_2643,N_2307,N_2356);
xor U2644 (N_2644,N_2364,N_2490);
or U2645 (N_2645,N_2455,N_2405);
nor U2646 (N_2646,N_2426,N_2268);
and U2647 (N_2647,N_2257,N_2297);
or U2648 (N_2648,N_2417,N_2309);
or U2649 (N_2649,N_2492,N_2379);
nor U2650 (N_2650,N_2333,N_2318);
nand U2651 (N_2651,N_2421,N_2416);
or U2652 (N_2652,N_2419,N_2442);
or U2653 (N_2653,N_2459,N_2398);
or U2654 (N_2654,N_2299,N_2419);
nand U2655 (N_2655,N_2278,N_2280);
and U2656 (N_2656,N_2400,N_2349);
nor U2657 (N_2657,N_2463,N_2488);
nand U2658 (N_2658,N_2288,N_2387);
nand U2659 (N_2659,N_2336,N_2390);
nand U2660 (N_2660,N_2357,N_2485);
nand U2661 (N_2661,N_2318,N_2422);
nand U2662 (N_2662,N_2467,N_2374);
and U2663 (N_2663,N_2387,N_2409);
nor U2664 (N_2664,N_2327,N_2395);
and U2665 (N_2665,N_2466,N_2322);
and U2666 (N_2666,N_2494,N_2258);
nand U2667 (N_2667,N_2365,N_2311);
and U2668 (N_2668,N_2424,N_2266);
or U2669 (N_2669,N_2288,N_2307);
nand U2670 (N_2670,N_2433,N_2328);
and U2671 (N_2671,N_2483,N_2260);
xor U2672 (N_2672,N_2457,N_2433);
nand U2673 (N_2673,N_2350,N_2289);
nand U2674 (N_2674,N_2409,N_2320);
and U2675 (N_2675,N_2275,N_2301);
nor U2676 (N_2676,N_2491,N_2377);
or U2677 (N_2677,N_2402,N_2480);
or U2678 (N_2678,N_2449,N_2379);
nor U2679 (N_2679,N_2437,N_2398);
nor U2680 (N_2680,N_2252,N_2402);
and U2681 (N_2681,N_2362,N_2372);
nor U2682 (N_2682,N_2481,N_2433);
or U2683 (N_2683,N_2356,N_2445);
or U2684 (N_2684,N_2444,N_2361);
and U2685 (N_2685,N_2372,N_2485);
xnor U2686 (N_2686,N_2289,N_2458);
xnor U2687 (N_2687,N_2480,N_2326);
nand U2688 (N_2688,N_2281,N_2284);
or U2689 (N_2689,N_2300,N_2415);
nand U2690 (N_2690,N_2472,N_2250);
xor U2691 (N_2691,N_2283,N_2250);
nand U2692 (N_2692,N_2261,N_2415);
nand U2693 (N_2693,N_2271,N_2269);
nand U2694 (N_2694,N_2383,N_2470);
or U2695 (N_2695,N_2291,N_2338);
nor U2696 (N_2696,N_2488,N_2285);
and U2697 (N_2697,N_2452,N_2478);
nor U2698 (N_2698,N_2285,N_2437);
and U2699 (N_2699,N_2370,N_2283);
xor U2700 (N_2700,N_2396,N_2262);
and U2701 (N_2701,N_2272,N_2271);
or U2702 (N_2702,N_2300,N_2463);
xor U2703 (N_2703,N_2388,N_2446);
nor U2704 (N_2704,N_2265,N_2262);
nand U2705 (N_2705,N_2449,N_2264);
xnor U2706 (N_2706,N_2394,N_2287);
and U2707 (N_2707,N_2306,N_2494);
nand U2708 (N_2708,N_2342,N_2461);
nor U2709 (N_2709,N_2392,N_2467);
or U2710 (N_2710,N_2430,N_2478);
nor U2711 (N_2711,N_2347,N_2292);
nand U2712 (N_2712,N_2326,N_2476);
nor U2713 (N_2713,N_2250,N_2350);
or U2714 (N_2714,N_2350,N_2298);
nor U2715 (N_2715,N_2454,N_2484);
nor U2716 (N_2716,N_2333,N_2370);
nand U2717 (N_2717,N_2384,N_2436);
nand U2718 (N_2718,N_2429,N_2309);
nor U2719 (N_2719,N_2456,N_2362);
or U2720 (N_2720,N_2333,N_2255);
xnor U2721 (N_2721,N_2484,N_2440);
nor U2722 (N_2722,N_2430,N_2354);
and U2723 (N_2723,N_2478,N_2290);
nor U2724 (N_2724,N_2427,N_2357);
or U2725 (N_2725,N_2494,N_2339);
or U2726 (N_2726,N_2347,N_2356);
xnor U2727 (N_2727,N_2320,N_2383);
xnor U2728 (N_2728,N_2440,N_2361);
xnor U2729 (N_2729,N_2427,N_2480);
and U2730 (N_2730,N_2290,N_2267);
nor U2731 (N_2731,N_2411,N_2422);
nand U2732 (N_2732,N_2378,N_2476);
xnor U2733 (N_2733,N_2352,N_2351);
and U2734 (N_2734,N_2410,N_2422);
xnor U2735 (N_2735,N_2431,N_2417);
and U2736 (N_2736,N_2472,N_2444);
xnor U2737 (N_2737,N_2394,N_2457);
and U2738 (N_2738,N_2254,N_2382);
and U2739 (N_2739,N_2499,N_2401);
nand U2740 (N_2740,N_2413,N_2381);
or U2741 (N_2741,N_2353,N_2451);
nand U2742 (N_2742,N_2317,N_2347);
and U2743 (N_2743,N_2444,N_2299);
nor U2744 (N_2744,N_2480,N_2449);
nor U2745 (N_2745,N_2335,N_2386);
xnor U2746 (N_2746,N_2412,N_2381);
and U2747 (N_2747,N_2356,N_2432);
or U2748 (N_2748,N_2426,N_2296);
xnor U2749 (N_2749,N_2440,N_2317);
and U2750 (N_2750,N_2556,N_2701);
or U2751 (N_2751,N_2531,N_2640);
or U2752 (N_2752,N_2634,N_2706);
nand U2753 (N_2753,N_2560,N_2532);
nand U2754 (N_2754,N_2605,N_2519);
xnor U2755 (N_2755,N_2696,N_2530);
nand U2756 (N_2756,N_2685,N_2680);
and U2757 (N_2757,N_2727,N_2650);
nand U2758 (N_2758,N_2636,N_2665);
nor U2759 (N_2759,N_2736,N_2645);
xnor U2760 (N_2760,N_2508,N_2611);
or U2761 (N_2761,N_2525,N_2565);
xnor U2762 (N_2762,N_2714,N_2666);
nand U2763 (N_2763,N_2596,N_2509);
and U2764 (N_2764,N_2593,N_2534);
xor U2765 (N_2765,N_2647,N_2687);
xor U2766 (N_2766,N_2747,N_2661);
and U2767 (N_2767,N_2579,N_2697);
or U2768 (N_2768,N_2651,N_2566);
or U2769 (N_2769,N_2553,N_2575);
xor U2770 (N_2770,N_2628,N_2742);
nor U2771 (N_2771,N_2540,N_2598);
and U2772 (N_2772,N_2613,N_2501);
nor U2773 (N_2773,N_2554,N_2510);
or U2774 (N_2774,N_2662,N_2577);
nand U2775 (N_2775,N_2582,N_2737);
xor U2776 (N_2776,N_2623,N_2709);
or U2777 (N_2777,N_2604,N_2734);
nor U2778 (N_2778,N_2619,N_2620);
or U2779 (N_2779,N_2589,N_2561);
nand U2780 (N_2780,N_2723,N_2739);
and U2781 (N_2781,N_2590,N_2683);
nor U2782 (N_2782,N_2621,N_2667);
xnor U2783 (N_2783,N_2542,N_2688);
xnor U2784 (N_2784,N_2733,N_2545);
nand U2785 (N_2785,N_2588,N_2555);
xor U2786 (N_2786,N_2644,N_2731);
xnor U2787 (N_2787,N_2691,N_2618);
or U2788 (N_2788,N_2559,N_2592);
nand U2789 (N_2789,N_2516,N_2726);
nor U2790 (N_2790,N_2669,N_2586);
nand U2791 (N_2791,N_2728,N_2622);
or U2792 (N_2792,N_2576,N_2643);
and U2793 (N_2793,N_2500,N_2513);
nor U2794 (N_2794,N_2672,N_2537);
or U2795 (N_2795,N_2626,N_2692);
nand U2796 (N_2796,N_2673,N_2646);
xor U2797 (N_2797,N_2695,N_2741);
and U2798 (N_2798,N_2625,N_2567);
and U2799 (N_2799,N_2738,N_2558);
xnor U2800 (N_2800,N_2583,N_2682);
or U2801 (N_2801,N_2631,N_2681);
nor U2802 (N_2802,N_2549,N_2551);
or U2803 (N_2803,N_2670,N_2599);
and U2804 (N_2804,N_2703,N_2719);
nor U2805 (N_2805,N_2656,N_2690);
and U2806 (N_2806,N_2711,N_2720);
or U2807 (N_2807,N_2538,N_2633);
or U2808 (N_2808,N_2704,N_2657);
and U2809 (N_2809,N_2686,N_2529);
or U2810 (N_2810,N_2684,N_2648);
and U2811 (N_2811,N_2595,N_2649);
or U2812 (N_2812,N_2608,N_2572);
xnor U2813 (N_2813,N_2746,N_2743);
nand U2814 (N_2814,N_2663,N_2518);
xor U2815 (N_2815,N_2600,N_2677);
nor U2816 (N_2816,N_2503,N_2713);
nand U2817 (N_2817,N_2652,N_2718);
nor U2818 (N_2818,N_2678,N_2543);
or U2819 (N_2819,N_2632,N_2710);
nor U2820 (N_2820,N_2616,N_2587);
and U2821 (N_2821,N_2522,N_2612);
and U2822 (N_2822,N_2527,N_2707);
nand U2823 (N_2823,N_2735,N_2674);
nand U2824 (N_2824,N_2536,N_2721);
xnor U2825 (N_2825,N_2610,N_2578);
and U2826 (N_2826,N_2574,N_2528);
nand U2827 (N_2827,N_2526,N_2629);
or U2828 (N_2828,N_2539,N_2664);
nor U2829 (N_2829,N_2521,N_2745);
and U2830 (N_2830,N_2635,N_2725);
nand U2831 (N_2831,N_2642,N_2506);
and U2832 (N_2832,N_2507,N_2627);
or U2833 (N_2833,N_2563,N_2698);
or U2834 (N_2834,N_2580,N_2729);
xnor U2835 (N_2835,N_2594,N_2571);
xnor U2836 (N_2836,N_2607,N_2693);
xor U2837 (N_2837,N_2675,N_2603);
nor U2838 (N_2838,N_2740,N_2689);
nand U2839 (N_2839,N_2562,N_2548);
nand U2840 (N_2840,N_2638,N_2544);
xor U2841 (N_2841,N_2515,N_2564);
xnor U2842 (N_2842,N_2505,N_2585);
xor U2843 (N_2843,N_2705,N_2514);
or U2844 (N_2844,N_2601,N_2557);
and U2845 (N_2845,N_2581,N_2732);
or U2846 (N_2846,N_2524,N_2748);
or U2847 (N_2847,N_2717,N_2584);
nor U2848 (N_2848,N_2653,N_2569);
or U2849 (N_2849,N_2517,N_2749);
or U2850 (N_2850,N_2523,N_2655);
nor U2851 (N_2851,N_2671,N_2654);
or U2852 (N_2852,N_2668,N_2679);
nor U2853 (N_2853,N_2617,N_2744);
or U2854 (N_2854,N_2541,N_2614);
or U2855 (N_2855,N_2512,N_2552);
or U2856 (N_2856,N_2658,N_2659);
xnor U2857 (N_2857,N_2702,N_2724);
xnor U2858 (N_2858,N_2730,N_2639);
or U2859 (N_2859,N_2624,N_2641);
nor U2860 (N_2860,N_2676,N_2716);
xnor U2861 (N_2861,N_2550,N_2694);
nand U2862 (N_2862,N_2606,N_2511);
nor U2863 (N_2863,N_2722,N_2699);
and U2864 (N_2864,N_2547,N_2535);
and U2865 (N_2865,N_2615,N_2609);
or U2866 (N_2866,N_2597,N_2502);
nand U2867 (N_2867,N_2637,N_2573);
nor U2868 (N_2868,N_2570,N_2660);
and U2869 (N_2869,N_2591,N_2546);
nor U2870 (N_2870,N_2520,N_2630);
nor U2871 (N_2871,N_2504,N_2700);
xor U2872 (N_2872,N_2708,N_2602);
or U2873 (N_2873,N_2533,N_2568);
and U2874 (N_2874,N_2712,N_2715);
xnor U2875 (N_2875,N_2629,N_2617);
or U2876 (N_2876,N_2543,N_2679);
xor U2877 (N_2877,N_2714,N_2702);
xor U2878 (N_2878,N_2569,N_2607);
nand U2879 (N_2879,N_2580,N_2515);
nor U2880 (N_2880,N_2530,N_2579);
and U2881 (N_2881,N_2642,N_2651);
nand U2882 (N_2882,N_2554,N_2626);
xnor U2883 (N_2883,N_2639,N_2711);
nor U2884 (N_2884,N_2725,N_2647);
or U2885 (N_2885,N_2566,N_2617);
nand U2886 (N_2886,N_2622,N_2556);
or U2887 (N_2887,N_2591,N_2604);
xor U2888 (N_2888,N_2644,N_2582);
xor U2889 (N_2889,N_2550,N_2723);
or U2890 (N_2890,N_2572,N_2748);
and U2891 (N_2891,N_2735,N_2687);
or U2892 (N_2892,N_2742,N_2727);
or U2893 (N_2893,N_2643,N_2742);
or U2894 (N_2894,N_2552,N_2612);
xnor U2895 (N_2895,N_2735,N_2737);
nor U2896 (N_2896,N_2582,N_2656);
or U2897 (N_2897,N_2682,N_2684);
xor U2898 (N_2898,N_2569,N_2501);
nor U2899 (N_2899,N_2621,N_2514);
and U2900 (N_2900,N_2655,N_2730);
and U2901 (N_2901,N_2606,N_2662);
or U2902 (N_2902,N_2516,N_2577);
xor U2903 (N_2903,N_2523,N_2570);
nand U2904 (N_2904,N_2681,N_2628);
or U2905 (N_2905,N_2731,N_2554);
nand U2906 (N_2906,N_2565,N_2524);
or U2907 (N_2907,N_2569,N_2636);
xor U2908 (N_2908,N_2513,N_2743);
xnor U2909 (N_2909,N_2516,N_2529);
and U2910 (N_2910,N_2667,N_2549);
nor U2911 (N_2911,N_2658,N_2689);
nand U2912 (N_2912,N_2601,N_2687);
xor U2913 (N_2913,N_2599,N_2595);
and U2914 (N_2914,N_2618,N_2653);
or U2915 (N_2915,N_2531,N_2593);
xor U2916 (N_2916,N_2704,N_2506);
and U2917 (N_2917,N_2742,N_2717);
nand U2918 (N_2918,N_2665,N_2528);
and U2919 (N_2919,N_2549,N_2557);
nand U2920 (N_2920,N_2649,N_2527);
nand U2921 (N_2921,N_2559,N_2729);
xor U2922 (N_2922,N_2668,N_2525);
or U2923 (N_2923,N_2696,N_2545);
and U2924 (N_2924,N_2723,N_2655);
nor U2925 (N_2925,N_2532,N_2686);
or U2926 (N_2926,N_2723,N_2717);
nand U2927 (N_2927,N_2671,N_2720);
and U2928 (N_2928,N_2684,N_2655);
and U2929 (N_2929,N_2512,N_2568);
or U2930 (N_2930,N_2590,N_2546);
and U2931 (N_2931,N_2650,N_2526);
and U2932 (N_2932,N_2541,N_2699);
xnor U2933 (N_2933,N_2549,N_2686);
nor U2934 (N_2934,N_2534,N_2662);
nand U2935 (N_2935,N_2717,N_2577);
nor U2936 (N_2936,N_2540,N_2698);
nand U2937 (N_2937,N_2682,N_2563);
or U2938 (N_2938,N_2636,N_2683);
xnor U2939 (N_2939,N_2689,N_2621);
xnor U2940 (N_2940,N_2690,N_2640);
nand U2941 (N_2941,N_2573,N_2681);
and U2942 (N_2942,N_2553,N_2681);
nand U2943 (N_2943,N_2511,N_2637);
or U2944 (N_2944,N_2554,N_2550);
nor U2945 (N_2945,N_2684,N_2546);
or U2946 (N_2946,N_2681,N_2638);
and U2947 (N_2947,N_2557,N_2509);
nor U2948 (N_2948,N_2544,N_2685);
and U2949 (N_2949,N_2738,N_2506);
xnor U2950 (N_2950,N_2575,N_2520);
and U2951 (N_2951,N_2742,N_2514);
and U2952 (N_2952,N_2634,N_2742);
nor U2953 (N_2953,N_2690,N_2688);
and U2954 (N_2954,N_2678,N_2654);
nand U2955 (N_2955,N_2541,N_2567);
nand U2956 (N_2956,N_2672,N_2556);
and U2957 (N_2957,N_2661,N_2609);
and U2958 (N_2958,N_2653,N_2544);
and U2959 (N_2959,N_2610,N_2539);
nor U2960 (N_2960,N_2717,N_2598);
nor U2961 (N_2961,N_2745,N_2623);
nand U2962 (N_2962,N_2712,N_2535);
nor U2963 (N_2963,N_2569,N_2552);
nand U2964 (N_2964,N_2634,N_2725);
nor U2965 (N_2965,N_2725,N_2713);
nand U2966 (N_2966,N_2540,N_2565);
xnor U2967 (N_2967,N_2549,N_2579);
and U2968 (N_2968,N_2714,N_2732);
nand U2969 (N_2969,N_2631,N_2527);
nor U2970 (N_2970,N_2577,N_2532);
nor U2971 (N_2971,N_2739,N_2505);
nor U2972 (N_2972,N_2712,N_2702);
nand U2973 (N_2973,N_2695,N_2716);
or U2974 (N_2974,N_2608,N_2713);
nor U2975 (N_2975,N_2546,N_2508);
nor U2976 (N_2976,N_2661,N_2745);
or U2977 (N_2977,N_2691,N_2702);
nand U2978 (N_2978,N_2669,N_2707);
nor U2979 (N_2979,N_2659,N_2535);
xnor U2980 (N_2980,N_2508,N_2501);
nand U2981 (N_2981,N_2514,N_2545);
nor U2982 (N_2982,N_2521,N_2632);
and U2983 (N_2983,N_2509,N_2563);
or U2984 (N_2984,N_2666,N_2648);
or U2985 (N_2985,N_2735,N_2749);
and U2986 (N_2986,N_2704,N_2547);
nand U2987 (N_2987,N_2725,N_2594);
nand U2988 (N_2988,N_2564,N_2581);
or U2989 (N_2989,N_2659,N_2716);
or U2990 (N_2990,N_2621,N_2699);
xnor U2991 (N_2991,N_2587,N_2605);
xnor U2992 (N_2992,N_2669,N_2559);
nand U2993 (N_2993,N_2573,N_2564);
and U2994 (N_2994,N_2610,N_2522);
nor U2995 (N_2995,N_2595,N_2622);
or U2996 (N_2996,N_2537,N_2651);
nor U2997 (N_2997,N_2744,N_2721);
nor U2998 (N_2998,N_2630,N_2536);
nor U2999 (N_2999,N_2723,N_2573);
xor U3000 (N_3000,N_2897,N_2880);
xnor U3001 (N_3001,N_2774,N_2885);
nand U3002 (N_3002,N_2988,N_2982);
and U3003 (N_3003,N_2758,N_2782);
xor U3004 (N_3004,N_2808,N_2812);
nor U3005 (N_3005,N_2950,N_2766);
nand U3006 (N_3006,N_2815,N_2964);
and U3007 (N_3007,N_2989,N_2901);
nor U3008 (N_3008,N_2846,N_2961);
nor U3009 (N_3009,N_2835,N_2765);
nand U3010 (N_3010,N_2759,N_2763);
nor U3011 (N_3011,N_2966,N_2911);
nand U3012 (N_3012,N_2868,N_2916);
or U3013 (N_3013,N_2893,N_2894);
xnor U3014 (N_3014,N_2956,N_2833);
xor U3015 (N_3015,N_2998,N_2898);
or U3016 (N_3016,N_2960,N_2990);
nor U3017 (N_3017,N_2972,N_2802);
nand U3018 (N_3018,N_2952,N_2849);
nor U3019 (N_3019,N_2983,N_2896);
nand U3020 (N_3020,N_2805,N_2884);
or U3021 (N_3021,N_2903,N_2752);
xnor U3022 (N_3022,N_2797,N_2912);
xor U3023 (N_3023,N_2855,N_2779);
or U3024 (N_3024,N_2858,N_2900);
nor U3025 (N_3025,N_2778,N_2847);
or U3026 (N_3026,N_2892,N_2940);
and U3027 (N_3027,N_2877,N_2790);
and U3028 (N_3028,N_2804,N_2936);
and U3029 (N_3029,N_2922,N_2965);
xor U3030 (N_3030,N_2913,N_2992);
and U3031 (N_3031,N_2934,N_2861);
nor U3032 (N_3032,N_2881,N_2906);
or U3033 (N_3033,N_2838,N_2895);
or U3034 (N_3034,N_2957,N_2785);
nor U3035 (N_3035,N_2879,N_2996);
nor U3036 (N_3036,N_2828,N_2902);
xnor U3037 (N_3037,N_2919,N_2968);
or U3038 (N_3038,N_2811,N_2888);
nor U3039 (N_3039,N_2920,N_2824);
xnor U3040 (N_3040,N_2818,N_2832);
or U3041 (N_3041,N_2869,N_2974);
nand U3042 (N_3042,N_2971,N_2946);
nand U3043 (N_3043,N_2866,N_2945);
nor U3044 (N_3044,N_2925,N_2874);
or U3045 (N_3045,N_2768,N_2784);
nand U3046 (N_3046,N_2969,N_2769);
xnor U3047 (N_3047,N_2840,N_2928);
nand U3048 (N_3048,N_2949,N_2848);
and U3049 (N_3049,N_2942,N_2841);
nand U3050 (N_3050,N_2886,N_2986);
and U3051 (N_3051,N_2856,N_2844);
or U3052 (N_3052,N_2924,N_2978);
xor U3053 (N_3053,N_2780,N_2870);
nand U3054 (N_3054,N_2979,N_2943);
nand U3055 (N_3055,N_2822,N_2984);
or U3056 (N_3056,N_2851,N_2944);
nand U3057 (N_3057,N_2921,N_2850);
nand U3058 (N_3058,N_2951,N_2939);
nand U3059 (N_3059,N_2825,N_2975);
and U3060 (N_3060,N_2904,N_2771);
xor U3061 (N_3061,N_2770,N_2862);
xnor U3062 (N_3062,N_2823,N_2923);
nor U3063 (N_3063,N_2908,N_2753);
xor U3064 (N_3064,N_2887,N_2754);
nand U3065 (N_3065,N_2757,N_2958);
nand U3066 (N_3066,N_2926,N_2854);
nor U3067 (N_3067,N_2830,N_2793);
nor U3068 (N_3068,N_2860,N_2963);
nand U3069 (N_3069,N_2997,N_2821);
and U3070 (N_3070,N_2935,N_2930);
nor U3071 (N_3071,N_2773,N_2801);
xnor U3072 (N_3072,N_2864,N_2937);
nand U3073 (N_3073,N_2967,N_2814);
or U3074 (N_3074,N_2867,N_2777);
nand U3075 (N_3075,N_2813,N_2786);
and U3076 (N_3076,N_2985,N_2816);
xnor U3077 (N_3077,N_2829,N_2762);
nand U3078 (N_3078,N_2938,N_2819);
or U3079 (N_3079,N_2918,N_2755);
or U3080 (N_3080,N_2800,N_2826);
nor U3081 (N_3081,N_2852,N_2932);
nand U3082 (N_3082,N_2905,N_2781);
nand U3083 (N_3083,N_2889,N_2863);
nor U3084 (N_3084,N_2875,N_2817);
xor U3085 (N_3085,N_2839,N_2917);
nand U3086 (N_3086,N_2791,N_2959);
and U3087 (N_3087,N_2994,N_2809);
nor U3088 (N_3088,N_2837,N_2842);
nand U3089 (N_3089,N_2853,N_2970);
nand U3090 (N_3090,N_2955,N_2987);
or U3091 (N_3091,N_2806,N_2798);
or U3092 (N_3092,N_2783,N_2991);
or U3093 (N_3093,N_2789,N_2976);
nor U3094 (N_3094,N_2764,N_2776);
nor U3095 (N_3095,N_2799,N_2907);
nor U3096 (N_3096,N_2767,N_2931);
nand U3097 (N_3097,N_2910,N_2792);
nor U3098 (N_3098,N_2756,N_2788);
or U3099 (N_3099,N_2795,N_2891);
or U3100 (N_3100,N_2873,N_2980);
and U3101 (N_3101,N_2948,N_2794);
xnor U3102 (N_3102,N_2834,N_2941);
nand U3103 (N_3103,N_2977,N_2876);
nor U3104 (N_3104,N_2843,N_2890);
nor U3105 (N_3105,N_2962,N_2807);
nand U3106 (N_3106,N_2927,N_2772);
xnor U3107 (N_3107,N_2953,N_2993);
and U3108 (N_3108,N_2796,N_2803);
and U3109 (N_3109,N_2883,N_2947);
nand U3110 (N_3110,N_2761,N_2914);
xor U3111 (N_3111,N_2981,N_2878);
nor U3112 (N_3112,N_2827,N_2831);
nor U3113 (N_3113,N_2999,N_2995);
or U3114 (N_3114,N_2909,N_2760);
or U3115 (N_3115,N_2871,N_2775);
nor U3116 (N_3116,N_2915,N_2954);
and U3117 (N_3117,N_2865,N_2845);
nand U3118 (N_3118,N_2929,N_2859);
or U3119 (N_3119,N_2820,N_2857);
and U3120 (N_3120,N_2899,N_2872);
or U3121 (N_3121,N_2787,N_2750);
and U3122 (N_3122,N_2882,N_2933);
xor U3123 (N_3123,N_2836,N_2973);
nor U3124 (N_3124,N_2751,N_2810);
xnor U3125 (N_3125,N_2899,N_2955);
nand U3126 (N_3126,N_2856,N_2993);
or U3127 (N_3127,N_2814,N_2833);
xor U3128 (N_3128,N_2760,N_2960);
nor U3129 (N_3129,N_2831,N_2962);
or U3130 (N_3130,N_2769,N_2866);
xnor U3131 (N_3131,N_2782,N_2783);
nor U3132 (N_3132,N_2803,N_2778);
or U3133 (N_3133,N_2988,N_2822);
nor U3134 (N_3134,N_2758,N_2885);
nand U3135 (N_3135,N_2879,N_2882);
or U3136 (N_3136,N_2821,N_2795);
nor U3137 (N_3137,N_2992,N_2975);
and U3138 (N_3138,N_2754,N_2874);
nand U3139 (N_3139,N_2944,N_2865);
nand U3140 (N_3140,N_2869,N_2887);
or U3141 (N_3141,N_2804,N_2798);
and U3142 (N_3142,N_2879,N_2784);
and U3143 (N_3143,N_2839,N_2993);
and U3144 (N_3144,N_2995,N_2869);
nor U3145 (N_3145,N_2841,N_2816);
and U3146 (N_3146,N_2946,N_2889);
nor U3147 (N_3147,N_2889,N_2994);
or U3148 (N_3148,N_2936,N_2872);
and U3149 (N_3149,N_2817,N_2871);
nand U3150 (N_3150,N_2983,N_2798);
nor U3151 (N_3151,N_2796,N_2887);
and U3152 (N_3152,N_2919,N_2901);
nand U3153 (N_3153,N_2891,N_2850);
and U3154 (N_3154,N_2878,N_2818);
or U3155 (N_3155,N_2983,N_2863);
nor U3156 (N_3156,N_2973,N_2982);
and U3157 (N_3157,N_2788,N_2823);
or U3158 (N_3158,N_2915,N_2918);
or U3159 (N_3159,N_2922,N_2913);
xor U3160 (N_3160,N_2966,N_2922);
nor U3161 (N_3161,N_2837,N_2761);
nand U3162 (N_3162,N_2757,N_2807);
or U3163 (N_3163,N_2920,N_2949);
nor U3164 (N_3164,N_2928,N_2894);
or U3165 (N_3165,N_2761,N_2826);
nor U3166 (N_3166,N_2982,N_2938);
nor U3167 (N_3167,N_2893,N_2805);
nand U3168 (N_3168,N_2782,N_2837);
or U3169 (N_3169,N_2892,N_2882);
or U3170 (N_3170,N_2792,N_2794);
or U3171 (N_3171,N_2803,N_2932);
or U3172 (N_3172,N_2786,N_2985);
and U3173 (N_3173,N_2901,N_2910);
xor U3174 (N_3174,N_2819,N_2906);
xnor U3175 (N_3175,N_2800,N_2788);
nor U3176 (N_3176,N_2979,N_2811);
or U3177 (N_3177,N_2830,N_2948);
xor U3178 (N_3178,N_2989,N_2842);
xnor U3179 (N_3179,N_2776,N_2757);
or U3180 (N_3180,N_2867,N_2853);
xnor U3181 (N_3181,N_2898,N_2788);
xnor U3182 (N_3182,N_2836,N_2782);
nand U3183 (N_3183,N_2983,N_2772);
nor U3184 (N_3184,N_2896,N_2825);
nor U3185 (N_3185,N_2977,N_2781);
xnor U3186 (N_3186,N_2811,N_2960);
or U3187 (N_3187,N_2773,N_2953);
nor U3188 (N_3188,N_2880,N_2967);
nor U3189 (N_3189,N_2885,N_2872);
nand U3190 (N_3190,N_2750,N_2964);
xor U3191 (N_3191,N_2964,N_2838);
or U3192 (N_3192,N_2780,N_2860);
nor U3193 (N_3193,N_2902,N_2888);
or U3194 (N_3194,N_2976,N_2906);
xnor U3195 (N_3195,N_2929,N_2953);
nor U3196 (N_3196,N_2875,N_2800);
nand U3197 (N_3197,N_2964,N_2907);
nor U3198 (N_3198,N_2970,N_2914);
nand U3199 (N_3199,N_2918,N_2848);
and U3200 (N_3200,N_2776,N_2937);
and U3201 (N_3201,N_2995,N_2905);
xor U3202 (N_3202,N_2944,N_2825);
nand U3203 (N_3203,N_2793,N_2858);
nor U3204 (N_3204,N_2883,N_2980);
or U3205 (N_3205,N_2988,N_2959);
or U3206 (N_3206,N_2750,N_2934);
or U3207 (N_3207,N_2952,N_2992);
nand U3208 (N_3208,N_2888,N_2796);
and U3209 (N_3209,N_2991,N_2896);
nand U3210 (N_3210,N_2948,N_2935);
xor U3211 (N_3211,N_2758,N_2993);
nand U3212 (N_3212,N_2810,N_2923);
and U3213 (N_3213,N_2896,N_2997);
or U3214 (N_3214,N_2932,N_2873);
or U3215 (N_3215,N_2773,N_2758);
nand U3216 (N_3216,N_2757,N_2915);
and U3217 (N_3217,N_2995,N_2825);
nor U3218 (N_3218,N_2872,N_2998);
xnor U3219 (N_3219,N_2835,N_2864);
xnor U3220 (N_3220,N_2977,N_2871);
and U3221 (N_3221,N_2750,N_2956);
and U3222 (N_3222,N_2963,N_2957);
and U3223 (N_3223,N_2961,N_2813);
and U3224 (N_3224,N_2829,N_2904);
or U3225 (N_3225,N_2894,N_2959);
nor U3226 (N_3226,N_2771,N_2912);
nor U3227 (N_3227,N_2972,N_2940);
or U3228 (N_3228,N_2884,N_2814);
xnor U3229 (N_3229,N_2961,N_2819);
xor U3230 (N_3230,N_2784,N_2782);
nand U3231 (N_3231,N_2764,N_2978);
nor U3232 (N_3232,N_2772,N_2996);
xor U3233 (N_3233,N_2981,N_2862);
and U3234 (N_3234,N_2955,N_2872);
or U3235 (N_3235,N_2911,N_2902);
or U3236 (N_3236,N_2957,N_2864);
nor U3237 (N_3237,N_2881,N_2819);
nand U3238 (N_3238,N_2893,N_2752);
nand U3239 (N_3239,N_2822,N_2833);
nand U3240 (N_3240,N_2791,N_2946);
and U3241 (N_3241,N_2894,N_2881);
and U3242 (N_3242,N_2801,N_2855);
xnor U3243 (N_3243,N_2987,N_2767);
nor U3244 (N_3244,N_2750,N_2751);
or U3245 (N_3245,N_2785,N_2962);
or U3246 (N_3246,N_2937,N_2917);
nor U3247 (N_3247,N_2796,N_2848);
nand U3248 (N_3248,N_2876,N_2948);
and U3249 (N_3249,N_2934,N_2778);
nor U3250 (N_3250,N_3019,N_3034);
or U3251 (N_3251,N_3047,N_3129);
nor U3252 (N_3252,N_3070,N_3012);
xnor U3253 (N_3253,N_3192,N_3037);
and U3254 (N_3254,N_3228,N_3089);
and U3255 (N_3255,N_3081,N_3184);
and U3256 (N_3256,N_3156,N_3105);
or U3257 (N_3257,N_3182,N_3014);
and U3258 (N_3258,N_3073,N_3246);
nand U3259 (N_3259,N_3234,N_3003);
xor U3260 (N_3260,N_3131,N_3122);
nand U3261 (N_3261,N_3226,N_3168);
and U3262 (N_3262,N_3169,N_3062);
nand U3263 (N_3263,N_3078,N_3083);
and U3264 (N_3264,N_3093,N_3204);
xnor U3265 (N_3265,N_3024,N_3229);
nor U3266 (N_3266,N_3187,N_3152);
nand U3267 (N_3267,N_3106,N_3243);
and U3268 (N_3268,N_3032,N_3209);
nand U3269 (N_3269,N_3038,N_3185);
nand U3270 (N_3270,N_3137,N_3202);
or U3271 (N_3271,N_3061,N_3028);
xnor U3272 (N_3272,N_3171,N_3084);
nand U3273 (N_3273,N_3102,N_3245);
xnor U3274 (N_3274,N_3099,N_3203);
nand U3275 (N_3275,N_3205,N_3180);
nor U3276 (N_3276,N_3159,N_3026);
or U3277 (N_3277,N_3216,N_3142);
xnor U3278 (N_3278,N_3086,N_3068);
or U3279 (N_3279,N_3053,N_3238);
nor U3280 (N_3280,N_3018,N_3095);
and U3281 (N_3281,N_3115,N_3045);
or U3282 (N_3282,N_3029,N_3139);
or U3283 (N_3283,N_3031,N_3186);
xor U3284 (N_3284,N_3021,N_3085);
xnor U3285 (N_3285,N_3001,N_3048);
and U3286 (N_3286,N_3136,N_3017);
nor U3287 (N_3287,N_3199,N_3221);
nand U3288 (N_3288,N_3235,N_3239);
and U3289 (N_3289,N_3125,N_3094);
or U3290 (N_3290,N_3213,N_3218);
nand U3291 (N_3291,N_3044,N_3002);
or U3292 (N_3292,N_3176,N_3097);
and U3293 (N_3293,N_3051,N_3178);
xnor U3294 (N_3294,N_3046,N_3076);
or U3295 (N_3295,N_3163,N_3007);
xor U3296 (N_3296,N_3058,N_3100);
xor U3297 (N_3297,N_3116,N_3030);
and U3298 (N_3298,N_3150,N_3191);
nand U3299 (N_3299,N_3049,N_3114);
and U3300 (N_3300,N_3013,N_3000);
nor U3301 (N_3301,N_3120,N_3067);
nor U3302 (N_3302,N_3040,N_3090);
nand U3303 (N_3303,N_3057,N_3056);
or U3304 (N_3304,N_3208,N_3195);
or U3305 (N_3305,N_3183,N_3157);
and U3306 (N_3306,N_3103,N_3211);
nor U3307 (N_3307,N_3091,N_3121);
and U3308 (N_3308,N_3127,N_3008);
nand U3309 (N_3309,N_3124,N_3227);
and U3310 (N_3310,N_3119,N_3217);
or U3311 (N_3311,N_3172,N_3009);
xnor U3312 (N_3312,N_3054,N_3098);
and U3313 (N_3313,N_3161,N_3027);
or U3314 (N_3314,N_3200,N_3166);
nand U3315 (N_3315,N_3167,N_3066);
nand U3316 (N_3316,N_3074,N_3079);
or U3317 (N_3317,N_3140,N_3052);
or U3318 (N_3318,N_3011,N_3237);
or U3319 (N_3319,N_3212,N_3110);
nor U3320 (N_3320,N_3035,N_3194);
nand U3321 (N_3321,N_3232,N_3214);
nor U3322 (N_3322,N_3155,N_3225);
and U3323 (N_3323,N_3112,N_3145);
xnor U3324 (N_3324,N_3181,N_3196);
or U3325 (N_3325,N_3077,N_3158);
or U3326 (N_3326,N_3064,N_3113);
xnor U3327 (N_3327,N_3177,N_3224);
or U3328 (N_3328,N_3022,N_3207);
xnor U3329 (N_3329,N_3015,N_3240);
or U3330 (N_3330,N_3020,N_3248);
nor U3331 (N_3331,N_3123,N_3118);
nor U3332 (N_3332,N_3060,N_3174);
and U3333 (N_3333,N_3088,N_3010);
xnor U3334 (N_3334,N_3175,N_3222);
and U3335 (N_3335,N_3126,N_3059);
xor U3336 (N_3336,N_3162,N_3165);
and U3337 (N_3337,N_3197,N_3242);
and U3338 (N_3338,N_3117,N_3146);
nor U3339 (N_3339,N_3154,N_3039);
xnor U3340 (N_3340,N_3033,N_3219);
nor U3341 (N_3341,N_3190,N_3188);
and U3342 (N_3342,N_3096,N_3087);
nor U3343 (N_3343,N_3050,N_3173);
xor U3344 (N_3344,N_3041,N_3233);
xnor U3345 (N_3345,N_3230,N_3107);
xnor U3346 (N_3346,N_3036,N_3042);
nand U3347 (N_3347,N_3104,N_3241);
or U3348 (N_3348,N_3170,N_3108);
nor U3349 (N_3349,N_3147,N_3135);
or U3350 (N_3350,N_3198,N_3016);
and U3351 (N_3351,N_3244,N_3130);
nand U3352 (N_3352,N_3111,N_3236);
xor U3353 (N_3353,N_3092,N_3249);
nand U3354 (N_3354,N_3071,N_3075);
or U3355 (N_3355,N_3148,N_3134);
or U3356 (N_3356,N_3138,N_3189);
nor U3357 (N_3357,N_3201,N_3069);
nor U3358 (N_3358,N_3080,N_3072);
nand U3359 (N_3359,N_3206,N_3160);
and U3360 (N_3360,N_3005,N_3164);
and U3361 (N_3361,N_3109,N_3004);
or U3362 (N_3362,N_3151,N_3055);
nand U3363 (N_3363,N_3043,N_3141);
nand U3364 (N_3364,N_3063,N_3082);
nor U3365 (N_3365,N_3144,N_3025);
or U3366 (N_3366,N_3128,N_3193);
nand U3367 (N_3367,N_3133,N_3247);
nand U3368 (N_3368,N_3132,N_3143);
and U3369 (N_3369,N_3220,N_3149);
xor U3370 (N_3370,N_3101,N_3210);
nor U3371 (N_3371,N_3006,N_3153);
nand U3372 (N_3372,N_3215,N_3223);
nand U3373 (N_3373,N_3231,N_3023);
and U3374 (N_3374,N_3179,N_3065);
xor U3375 (N_3375,N_3244,N_3062);
or U3376 (N_3376,N_3091,N_3134);
nor U3377 (N_3377,N_3076,N_3078);
xnor U3378 (N_3378,N_3106,N_3211);
or U3379 (N_3379,N_3169,N_3149);
nor U3380 (N_3380,N_3133,N_3175);
xor U3381 (N_3381,N_3226,N_3127);
nand U3382 (N_3382,N_3126,N_3061);
xnor U3383 (N_3383,N_3150,N_3111);
xor U3384 (N_3384,N_3077,N_3069);
nand U3385 (N_3385,N_3013,N_3249);
nand U3386 (N_3386,N_3023,N_3210);
or U3387 (N_3387,N_3056,N_3230);
or U3388 (N_3388,N_3244,N_3219);
nand U3389 (N_3389,N_3073,N_3186);
nor U3390 (N_3390,N_3170,N_3239);
or U3391 (N_3391,N_3072,N_3123);
xor U3392 (N_3392,N_3040,N_3119);
or U3393 (N_3393,N_3089,N_3051);
nand U3394 (N_3394,N_3082,N_3102);
nor U3395 (N_3395,N_3197,N_3231);
and U3396 (N_3396,N_3231,N_3188);
and U3397 (N_3397,N_3192,N_3242);
nand U3398 (N_3398,N_3221,N_3033);
xor U3399 (N_3399,N_3010,N_3026);
and U3400 (N_3400,N_3016,N_3082);
xnor U3401 (N_3401,N_3106,N_3060);
and U3402 (N_3402,N_3147,N_3029);
nor U3403 (N_3403,N_3103,N_3106);
nand U3404 (N_3404,N_3128,N_3039);
or U3405 (N_3405,N_3175,N_3079);
or U3406 (N_3406,N_3231,N_3204);
nor U3407 (N_3407,N_3245,N_3107);
nor U3408 (N_3408,N_3187,N_3064);
nand U3409 (N_3409,N_3048,N_3122);
xnor U3410 (N_3410,N_3184,N_3150);
nand U3411 (N_3411,N_3037,N_3146);
or U3412 (N_3412,N_3027,N_3007);
and U3413 (N_3413,N_3012,N_3159);
nor U3414 (N_3414,N_3026,N_3054);
xnor U3415 (N_3415,N_3025,N_3100);
nor U3416 (N_3416,N_3153,N_3050);
or U3417 (N_3417,N_3156,N_3040);
xor U3418 (N_3418,N_3210,N_3135);
or U3419 (N_3419,N_3084,N_3242);
nand U3420 (N_3420,N_3114,N_3061);
nand U3421 (N_3421,N_3075,N_3161);
nor U3422 (N_3422,N_3064,N_3137);
or U3423 (N_3423,N_3135,N_3189);
nand U3424 (N_3424,N_3049,N_3173);
and U3425 (N_3425,N_3059,N_3058);
and U3426 (N_3426,N_3179,N_3064);
and U3427 (N_3427,N_3166,N_3013);
nor U3428 (N_3428,N_3161,N_3219);
xor U3429 (N_3429,N_3052,N_3059);
nand U3430 (N_3430,N_3165,N_3231);
xor U3431 (N_3431,N_3092,N_3013);
nand U3432 (N_3432,N_3046,N_3230);
and U3433 (N_3433,N_3028,N_3204);
nand U3434 (N_3434,N_3013,N_3174);
or U3435 (N_3435,N_3178,N_3139);
xor U3436 (N_3436,N_3184,N_3218);
xor U3437 (N_3437,N_3201,N_3037);
nand U3438 (N_3438,N_3029,N_3143);
or U3439 (N_3439,N_3068,N_3089);
nand U3440 (N_3440,N_3013,N_3167);
or U3441 (N_3441,N_3209,N_3138);
nor U3442 (N_3442,N_3216,N_3010);
xnor U3443 (N_3443,N_3225,N_3041);
and U3444 (N_3444,N_3123,N_3179);
or U3445 (N_3445,N_3219,N_3153);
xnor U3446 (N_3446,N_3203,N_3082);
and U3447 (N_3447,N_3081,N_3033);
nand U3448 (N_3448,N_3244,N_3030);
xor U3449 (N_3449,N_3061,N_3091);
xor U3450 (N_3450,N_3228,N_3248);
nor U3451 (N_3451,N_3023,N_3174);
xnor U3452 (N_3452,N_3167,N_3130);
xnor U3453 (N_3453,N_3155,N_3217);
or U3454 (N_3454,N_3143,N_3194);
xor U3455 (N_3455,N_3067,N_3225);
xor U3456 (N_3456,N_3237,N_3183);
or U3457 (N_3457,N_3239,N_3151);
nand U3458 (N_3458,N_3022,N_3112);
xnor U3459 (N_3459,N_3067,N_3105);
nand U3460 (N_3460,N_3177,N_3157);
xor U3461 (N_3461,N_3021,N_3095);
xor U3462 (N_3462,N_3203,N_3205);
or U3463 (N_3463,N_3020,N_3107);
xor U3464 (N_3464,N_3154,N_3090);
xnor U3465 (N_3465,N_3138,N_3131);
and U3466 (N_3466,N_3137,N_3194);
or U3467 (N_3467,N_3170,N_3101);
nor U3468 (N_3468,N_3203,N_3238);
and U3469 (N_3469,N_3139,N_3148);
or U3470 (N_3470,N_3086,N_3158);
xor U3471 (N_3471,N_3244,N_3140);
nor U3472 (N_3472,N_3033,N_3247);
nand U3473 (N_3473,N_3091,N_3176);
nor U3474 (N_3474,N_3213,N_3207);
xnor U3475 (N_3475,N_3209,N_3141);
xnor U3476 (N_3476,N_3202,N_3047);
and U3477 (N_3477,N_3061,N_3145);
nand U3478 (N_3478,N_3064,N_3046);
nor U3479 (N_3479,N_3091,N_3219);
or U3480 (N_3480,N_3013,N_3016);
nor U3481 (N_3481,N_3180,N_3026);
or U3482 (N_3482,N_3082,N_3012);
nand U3483 (N_3483,N_3245,N_3010);
xor U3484 (N_3484,N_3087,N_3249);
xor U3485 (N_3485,N_3093,N_3176);
xor U3486 (N_3486,N_3165,N_3230);
or U3487 (N_3487,N_3128,N_3194);
and U3488 (N_3488,N_3184,N_3110);
xor U3489 (N_3489,N_3187,N_3185);
nor U3490 (N_3490,N_3196,N_3065);
xor U3491 (N_3491,N_3141,N_3246);
or U3492 (N_3492,N_3051,N_3113);
or U3493 (N_3493,N_3046,N_3075);
or U3494 (N_3494,N_3100,N_3134);
nor U3495 (N_3495,N_3159,N_3059);
or U3496 (N_3496,N_3016,N_3025);
and U3497 (N_3497,N_3201,N_3080);
nor U3498 (N_3498,N_3236,N_3036);
nor U3499 (N_3499,N_3198,N_3218);
nand U3500 (N_3500,N_3275,N_3333);
or U3501 (N_3501,N_3498,N_3475);
xor U3502 (N_3502,N_3369,N_3420);
and U3503 (N_3503,N_3331,N_3439);
nand U3504 (N_3504,N_3457,N_3378);
or U3505 (N_3505,N_3251,N_3325);
and U3506 (N_3506,N_3414,N_3407);
nand U3507 (N_3507,N_3412,N_3484);
or U3508 (N_3508,N_3421,N_3317);
or U3509 (N_3509,N_3358,N_3494);
xnor U3510 (N_3510,N_3393,N_3499);
or U3511 (N_3511,N_3367,N_3336);
and U3512 (N_3512,N_3303,N_3487);
xnor U3513 (N_3513,N_3370,N_3423);
nor U3514 (N_3514,N_3282,N_3448);
nand U3515 (N_3515,N_3474,N_3352);
nor U3516 (N_3516,N_3426,N_3322);
or U3517 (N_3517,N_3374,N_3492);
xnor U3518 (N_3518,N_3360,N_3302);
and U3519 (N_3519,N_3337,N_3372);
or U3520 (N_3520,N_3306,N_3481);
and U3521 (N_3521,N_3383,N_3379);
and U3522 (N_3522,N_3279,N_3418);
nor U3523 (N_3523,N_3410,N_3459);
nand U3524 (N_3524,N_3416,N_3485);
nor U3525 (N_3525,N_3315,N_3253);
nand U3526 (N_3526,N_3375,N_3347);
nor U3527 (N_3527,N_3404,N_3344);
xnor U3528 (N_3528,N_3376,N_3364);
xnor U3529 (N_3529,N_3283,N_3377);
nand U3530 (N_3530,N_3497,N_3434);
nor U3531 (N_3531,N_3483,N_3281);
nor U3532 (N_3532,N_3478,N_3396);
xnor U3533 (N_3533,N_3428,N_3442);
xor U3534 (N_3534,N_3384,N_3400);
or U3535 (N_3535,N_3305,N_3272);
nor U3536 (N_3536,N_3339,N_3263);
xor U3537 (N_3537,N_3346,N_3465);
xnor U3538 (N_3538,N_3461,N_3496);
xnor U3539 (N_3539,N_3311,N_3354);
or U3540 (N_3540,N_3493,N_3271);
nor U3541 (N_3541,N_3313,N_3309);
and U3542 (N_3542,N_3291,N_3334);
and U3543 (N_3543,N_3362,N_3489);
and U3544 (N_3544,N_3264,N_3326);
nand U3545 (N_3545,N_3385,N_3327);
nand U3546 (N_3546,N_3301,N_3390);
and U3547 (N_3547,N_3386,N_3340);
and U3548 (N_3548,N_3366,N_3401);
nand U3549 (N_3549,N_3330,N_3402);
nand U3550 (N_3550,N_3391,N_3329);
nor U3551 (N_3551,N_3293,N_3389);
and U3552 (N_3552,N_3350,N_3357);
nor U3553 (N_3553,N_3268,N_3314);
or U3554 (N_3554,N_3463,N_3419);
nand U3555 (N_3555,N_3411,N_3335);
or U3556 (N_3556,N_3368,N_3365);
nor U3557 (N_3557,N_3491,N_3287);
nor U3558 (N_3558,N_3332,N_3417);
and U3559 (N_3559,N_3468,N_3394);
nand U3560 (N_3560,N_3467,N_3424);
xor U3561 (N_3561,N_3297,N_3342);
xor U3562 (N_3562,N_3257,N_3443);
or U3563 (N_3563,N_3278,N_3361);
or U3564 (N_3564,N_3298,N_3296);
or U3565 (N_3565,N_3260,N_3318);
and U3566 (N_3566,N_3415,N_3324);
or U3567 (N_3567,N_3250,N_3464);
or U3568 (N_3568,N_3274,N_3422);
nand U3569 (N_3569,N_3295,N_3458);
and U3570 (N_3570,N_3425,N_3265);
or U3571 (N_3571,N_3310,N_3321);
and U3572 (N_3572,N_3280,N_3399);
nand U3573 (N_3573,N_3363,N_3398);
or U3574 (N_3574,N_3288,N_3254);
and U3575 (N_3575,N_3433,N_3444);
nand U3576 (N_3576,N_3447,N_3453);
xnor U3577 (N_3577,N_3482,N_3446);
nor U3578 (N_3578,N_3450,N_3276);
nand U3579 (N_3579,N_3353,N_3452);
and U3580 (N_3580,N_3256,N_3359);
and U3581 (N_3581,N_3307,N_3395);
nor U3582 (N_3582,N_3472,N_3351);
and U3583 (N_3583,N_3266,N_3308);
nand U3584 (N_3584,N_3338,N_3408);
and U3585 (N_3585,N_3294,N_3381);
or U3586 (N_3586,N_3462,N_3388);
nor U3587 (N_3587,N_3409,N_3285);
nor U3588 (N_3588,N_3460,N_3471);
nand U3589 (N_3589,N_3392,N_3341);
nor U3590 (N_3590,N_3455,N_3441);
xor U3591 (N_3591,N_3427,N_3328);
or U3592 (N_3592,N_3255,N_3429);
nor U3593 (N_3593,N_3270,N_3316);
and U3594 (N_3594,N_3300,N_3406);
xnor U3595 (N_3595,N_3284,N_3349);
or U3596 (N_3596,N_3435,N_3345);
and U3597 (N_3597,N_3486,N_3405);
and U3598 (N_3598,N_3262,N_3430);
nand U3599 (N_3599,N_3371,N_3437);
nand U3600 (N_3600,N_3312,N_3380);
nor U3601 (N_3601,N_3403,N_3319);
or U3602 (N_3602,N_3292,N_3320);
nor U3603 (N_3603,N_3436,N_3290);
or U3604 (N_3604,N_3299,N_3466);
nand U3605 (N_3605,N_3480,N_3289);
xor U3606 (N_3606,N_3304,N_3473);
or U3607 (N_3607,N_3470,N_3490);
and U3608 (N_3608,N_3495,N_3356);
and U3609 (N_3609,N_3343,N_3323);
and U3610 (N_3610,N_3252,N_3477);
xor U3611 (N_3611,N_3382,N_3397);
nand U3612 (N_3612,N_3348,N_3476);
nand U3613 (N_3613,N_3440,N_3469);
nand U3614 (N_3614,N_3269,N_3373);
or U3615 (N_3615,N_3277,N_3259);
and U3616 (N_3616,N_3456,N_3479);
nand U3617 (N_3617,N_3432,N_3438);
or U3618 (N_3618,N_3261,N_3387);
nand U3619 (N_3619,N_3451,N_3355);
nand U3620 (N_3620,N_3413,N_3445);
nor U3621 (N_3621,N_3273,N_3431);
or U3622 (N_3622,N_3258,N_3267);
xor U3623 (N_3623,N_3454,N_3286);
or U3624 (N_3624,N_3449,N_3488);
xnor U3625 (N_3625,N_3266,N_3315);
nand U3626 (N_3626,N_3427,N_3456);
nand U3627 (N_3627,N_3309,N_3291);
xor U3628 (N_3628,N_3295,N_3293);
nor U3629 (N_3629,N_3263,N_3269);
nor U3630 (N_3630,N_3415,N_3256);
xnor U3631 (N_3631,N_3403,N_3271);
and U3632 (N_3632,N_3490,N_3292);
xnor U3633 (N_3633,N_3323,N_3304);
xor U3634 (N_3634,N_3395,N_3476);
nand U3635 (N_3635,N_3278,N_3305);
nand U3636 (N_3636,N_3304,N_3458);
nand U3637 (N_3637,N_3386,N_3317);
nand U3638 (N_3638,N_3373,N_3343);
xor U3639 (N_3639,N_3284,N_3338);
and U3640 (N_3640,N_3370,N_3481);
nand U3641 (N_3641,N_3418,N_3455);
and U3642 (N_3642,N_3339,N_3422);
nand U3643 (N_3643,N_3488,N_3398);
or U3644 (N_3644,N_3318,N_3271);
nor U3645 (N_3645,N_3278,N_3337);
nand U3646 (N_3646,N_3419,N_3455);
nand U3647 (N_3647,N_3299,N_3314);
or U3648 (N_3648,N_3467,N_3488);
nand U3649 (N_3649,N_3362,N_3334);
nor U3650 (N_3650,N_3302,N_3365);
and U3651 (N_3651,N_3336,N_3310);
nand U3652 (N_3652,N_3443,N_3299);
nand U3653 (N_3653,N_3322,N_3314);
nor U3654 (N_3654,N_3326,N_3332);
xor U3655 (N_3655,N_3300,N_3293);
nand U3656 (N_3656,N_3309,N_3499);
xor U3657 (N_3657,N_3266,N_3314);
and U3658 (N_3658,N_3489,N_3408);
nand U3659 (N_3659,N_3446,N_3357);
nor U3660 (N_3660,N_3400,N_3448);
and U3661 (N_3661,N_3331,N_3475);
nor U3662 (N_3662,N_3383,N_3407);
nor U3663 (N_3663,N_3321,N_3377);
or U3664 (N_3664,N_3419,N_3347);
and U3665 (N_3665,N_3499,N_3278);
nand U3666 (N_3666,N_3478,N_3375);
xnor U3667 (N_3667,N_3341,N_3390);
and U3668 (N_3668,N_3439,N_3328);
or U3669 (N_3669,N_3454,N_3362);
xnor U3670 (N_3670,N_3294,N_3275);
nand U3671 (N_3671,N_3284,N_3431);
nor U3672 (N_3672,N_3288,N_3490);
xnor U3673 (N_3673,N_3311,N_3407);
nand U3674 (N_3674,N_3310,N_3279);
and U3675 (N_3675,N_3427,N_3385);
xor U3676 (N_3676,N_3467,N_3316);
nor U3677 (N_3677,N_3439,N_3305);
and U3678 (N_3678,N_3458,N_3253);
or U3679 (N_3679,N_3384,N_3423);
xor U3680 (N_3680,N_3260,N_3288);
nor U3681 (N_3681,N_3468,N_3312);
nor U3682 (N_3682,N_3423,N_3371);
xnor U3683 (N_3683,N_3410,N_3250);
nand U3684 (N_3684,N_3467,N_3416);
nor U3685 (N_3685,N_3400,N_3254);
nor U3686 (N_3686,N_3475,N_3393);
and U3687 (N_3687,N_3414,N_3442);
nand U3688 (N_3688,N_3450,N_3323);
nand U3689 (N_3689,N_3370,N_3425);
and U3690 (N_3690,N_3367,N_3383);
or U3691 (N_3691,N_3277,N_3490);
xor U3692 (N_3692,N_3444,N_3312);
nand U3693 (N_3693,N_3333,N_3331);
xnor U3694 (N_3694,N_3405,N_3423);
xnor U3695 (N_3695,N_3378,N_3422);
nor U3696 (N_3696,N_3430,N_3389);
nor U3697 (N_3697,N_3252,N_3387);
and U3698 (N_3698,N_3385,N_3309);
nand U3699 (N_3699,N_3342,N_3371);
and U3700 (N_3700,N_3378,N_3292);
nand U3701 (N_3701,N_3441,N_3325);
xor U3702 (N_3702,N_3383,N_3276);
nand U3703 (N_3703,N_3285,N_3268);
xnor U3704 (N_3704,N_3472,N_3311);
and U3705 (N_3705,N_3364,N_3316);
nor U3706 (N_3706,N_3348,N_3435);
or U3707 (N_3707,N_3481,N_3479);
or U3708 (N_3708,N_3395,N_3440);
xor U3709 (N_3709,N_3419,N_3344);
nand U3710 (N_3710,N_3329,N_3251);
xnor U3711 (N_3711,N_3437,N_3481);
xor U3712 (N_3712,N_3264,N_3484);
nor U3713 (N_3713,N_3318,N_3335);
nor U3714 (N_3714,N_3333,N_3416);
nor U3715 (N_3715,N_3396,N_3470);
xor U3716 (N_3716,N_3336,N_3254);
nor U3717 (N_3717,N_3310,N_3445);
or U3718 (N_3718,N_3390,N_3404);
and U3719 (N_3719,N_3329,N_3272);
and U3720 (N_3720,N_3420,N_3258);
nand U3721 (N_3721,N_3397,N_3319);
and U3722 (N_3722,N_3439,N_3267);
and U3723 (N_3723,N_3286,N_3443);
nor U3724 (N_3724,N_3260,N_3353);
nor U3725 (N_3725,N_3402,N_3380);
xnor U3726 (N_3726,N_3455,N_3499);
or U3727 (N_3727,N_3353,N_3444);
xnor U3728 (N_3728,N_3312,N_3443);
and U3729 (N_3729,N_3378,N_3303);
nand U3730 (N_3730,N_3386,N_3414);
xnor U3731 (N_3731,N_3469,N_3291);
xor U3732 (N_3732,N_3417,N_3457);
or U3733 (N_3733,N_3394,N_3330);
xnor U3734 (N_3734,N_3487,N_3276);
or U3735 (N_3735,N_3256,N_3342);
or U3736 (N_3736,N_3479,N_3348);
and U3737 (N_3737,N_3430,N_3483);
nor U3738 (N_3738,N_3422,N_3273);
or U3739 (N_3739,N_3342,N_3438);
xnor U3740 (N_3740,N_3318,N_3497);
xor U3741 (N_3741,N_3336,N_3284);
nand U3742 (N_3742,N_3342,N_3449);
and U3743 (N_3743,N_3305,N_3386);
nor U3744 (N_3744,N_3401,N_3298);
xnor U3745 (N_3745,N_3464,N_3337);
xnor U3746 (N_3746,N_3368,N_3481);
nor U3747 (N_3747,N_3397,N_3473);
xnor U3748 (N_3748,N_3291,N_3297);
or U3749 (N_3749,N_3396,N_3253);
and U3750 (N_3750,N_3690,N_3597);
nand U3751 (N_3751,N_3577,N_3562);
nor U3752 (N_3752,N_3634,N_3726);
and U3753 (N_3753,N_3607,N_3600);
and U3754 (N_3754,N_3630,N_3549);
nor U3755 (N_3755,N_3535,N_3512);
nor U3756 (N_3756,N_3553,N_3640);
nand U3757 (N_3757,N_3674,N_3656);
xor U3758 (N_3758,N_3560,N_3647);
nor U3759 (N_3759,N_3529,N_3532);
xnor U3760 (N_3760,N_3705,N_3525);
nor U3761 (N_3761,N_3661,N_3644);
nor U3762 (N_3762,N_3722,N_3591);
and U3763 (N_3763,N_3626,N_3513);
and U3764 (N_3764,N_3703,N_3531);
nor U3765 (N_3765,N_3565,N_3524);
nor U3766 (N_3766,N_3730,N_3545);
xnor U3767 (N_3767,N_3625,N_3541);
and U3768 (N_3768,N_3677,N_3701);
nor U3769 (N_3769,N_3696,N_3624);
nor U3770 (N_3770,N_3686,N_3694);
nor U3771 (N_3771,N_3539,N_3592);
nor U3772 (N_3772,N_3594,N_3520);
nand U3773 (N_3773,N_3516,N_3582);
and U3774 (N_3774,N_3645,N_3676);
or U3775 (N_3775,N_3663,N_3551);
nor U3776 (N_3776,N_3585,N_3540);
or U3777 (N_3777,N_3604,N_3507);
or U3778 (N_3778,N_3695,N_3687);
xnor U3779 (N_3779,N_3713,N_3558);
nand U3780 (N_3780,N_3720,N_3574);
nand U3781 (N_3781,N_3724,N_3590);
and U3782 (N_3782,N_3537,N_3559);
or U3783 (N_3783,N_3614,N_3605);
nor U3784 (N_3784,N_3621,N_3567);
xor U3785 (N_3785,N_3685,N_3650);
or U3786 (N_3786,N_3627,N_3564);
and U3787 (N_3787,N_3514,N_3623);
nand U3788 (N_3788,N_3629,N_3569);
and U3789 (N_3789,N_3671,N_3509);
xor U3790 (N_3790,N_3723,N_3683);
nor U3791 (N_3791,N_3547,N_3662);
nand U3792 (N_3792,N_3572,N_3533);
or U3793 (N_3793,N_3588,N_3746);
xor U3794 (N_3794,N_3620,N_3680);
and U3795 (N_3795,N_3631,N_3527);
and U3796 (N_3796,N_3733,N_3519);
and U3797 (N_3797,N_3670,N_3700);
and U3798 (N_3798,N_3616,N_3609);
xor U3799 (N_3799,N_3727,N_3708);
or U3800 (N_3800,N_3579,N_3688);
or U3801 (N_3801,N_3575,N_3717);
nor U3802 (N_3802,N_3595,N_3578);
and U3803 (N_3803,N_3593,N_3521);
nand U3804 (N_3804,N_3666,N_3504);
or U3805 (N_3805,N_3704,N_3611);
or U3806 (N_3806,N_3500,N_3745);
and U3807 (N_3807,N_3603,N_3652);
or U3808 (N_3808,N_3530,N_3546);
nor U3809 (N_3809,N_3502,N_3550);
and U3810 (N_3810,N_3668,N_3568);
or U3811 (N_3811,N_3736,N_3684);
and U3812 (N_3812,N_3654,N_3747);
xor U3813 (N_3813,N_3526,N_3664);
nor U3814 (N_3814,N_3602,N_3682);
and U3815 (N_3815,N_3693,N_3731);
nand U3816 (N_3816,N_3710,N_3675);
xor U3817 (N_3817,N_3641,N_3544);
nor U3818 (N_3818,N_3698,N_3584);
or U3819 (N_3819,N_3732,N_3503);
xor U3820 (N_3820,N_3718,N_3543);
xnor U3821 (N_3821,N_3639,N_3598);
nand U3822 (N_3822,N_3534,N_3749);
nor U3823 (N_3823,N_3721,N_3658);
or U3824 (N_3824,N_3643,N_3744);
xor U3825 (N_3825,N_3743,N_3505);
and U3826 (N_3826,N_3587,N_3714);
or U3827 (N_3827,N_3649,N_3612);
or U3828 (N_3828,N_3515,N_3608);
nand U3829 (N_3829,N_3518,N_3511);
nor U3830 (N_3830,N_3699,N_3660);
nand U3831 (N_3831,N_3622,N_3536);
nand U3832 (N_3832,N_3542,N_3729);
xnor U3833 (N_3833,N_3734,N_3655);
nor U3834 (N_3834,N_3702,N_3646);
nand U3835 (N_3835,N_3555,N_3738);
nor U3836 (N_3836,N_3617,N_3667);
and U3837 (N_3837,N_3566,N_3659);
nor U3838 (N_3838,N_3712,N_3508);
nor U3839 (N_3839,N_3692,N_3635);
nor U3840 (N_3840,N_3711,N_3678);
nand U3841 (N_3841,N_3632,N_3707);
nor U3842 (N_3842,N_3725,N_3552);
nor U3843 (N_3843,N_3601,N_3580);
and U3844 (N_3844,N_3596,N_3653);
and U3845 (N_3845,N_3571,N_3583);
nor U3846 (N_3846,N_3672,N_3741);
or U3847 (N_3847,N_3665,N_3735);
nand U3848 (N_3848,N_3556,N_3673);
nor U3849 (N_3849,N_3610,N_3669);
or U3850 (N_3850,N_3538,N_3510);
or U3851 (N_3851,N_3522,N_3563);
or U3852 (N_3852,N_3691,N_3618);
nand U3853 (N_3853,N_3581,N_3528);
nand U3854 (N_3854,N_3648,N_3606);
xnor U3855 (N_3855,N_3554,N_3709);
xnor U3856 (N_3856,N_3679,N_3576);
or U3857 (N_3857,N_3615,N_3657);
or U3858 (N_3858,N_3506,N_3613);
xnor U3859 (N_3859,N_3651,N_3728);
or U3860 (N_3860,N_3517,N_3742);
or U3861 (N_3861,N_3748,N_3548);
xnor U3862 (N_3862,N_3681,N_3633);
nor U3863 (N_3863,N_3740,N_3619);
xnor U3864 (N_3864,N_3636,N_3570);
or U3865 (N_3865,N_3523,N_3637);
nand U3866 (N_3866,N_3719,N_3586);
nand U3867 (N_3867,N_3706,N_3557);
xnor U3868 (N_3868,N_3501,N_3642);
xnor U3869 (N_3869,N_3689,N_3697);
xor U3870 (N_3870,N_3739,N_3589);
or U3871 (N_3871,N_3628,N_3573);
nor U3872 (N_3872,N_3561,N_3716);
and U3873 (N_3873,N_3599,N_3737);
nor U3874 (N_3874,N_3638,N_3715);
nand U3875 (N_3875,N_3515,N_3618);
or U3876 (N_3876,N_3588,N_3711);
nand U3877 (N_3877,N_3522,N_3693);
nor U3878 (N_3878,N_3745,N_3607);
or U3879 (N_3879,N_3701,N_3540);
nand U3880 (N_3880,N_3742,N_3577);
nand U3881 (N_3881,N_3695,N_3534);
xnor U3882 (N_3882,N_3532,N_3591);
nor U3883 (N_3883,N_3598,N_3698);
and U3884 (N_3884,N_3531,N_3539);
or U3885 (N_3885,N_3627,N_3710);
nor U3886 (N_3886,N_3546,N_3517);
or U3887 (N_3887,N_3723,N_3520);
nor U3888 (N_3888,N_3606,N_3730);
nor U3889 (N_3889,N_3727,N_3554);
nor U3890 (N_3890,N_3699,N_3506);
xnor U3891 (N_3891,N_3657,N_3649);
nand U3892 (N_3892,N_3557,N_3632);
or U3893 (N_3893,N_3685,N_3726);
nor U3894 (N_3894,N_3537,N_3638);
nor U3895 (N_3895,N_3649,N_3712);
nand U3896 (N_3896,N_3596,N_3524);
or U3897 (N_3897,N_3658,N_3741);
nand U3898 (N_3898,N_3644,N_3574);
xnor U3899 (N_3899,N_3693,N_3549);
or U3900 (N_3900,N_3521,N_3708);
and U3901 (N_3901,N_3548,N_3504);
and U3902 (N_3902,N_3649,N_3717);
xor U3903 (N_3903,N_3574,N_3704);
or U3904 (N_3904,N_3653,N_3520);
nand U3905 (N_3905,N_3567,N_3719);
nor U3906 (N_3906,N_3659,N_3519);
xnor U3907 (N_3907,N_3598,N_3610);
nor U3908 (N_3908,N_3740,N_3539);
or U3909 (N_3909,N_3580,N_3674);
nand U3910 (N_3910,N_3720,N_3597);
or U3911 (N_3911,N_3640,N_3670);
and U3912 (N_3912,N_3519,N_3674);
nand U3913 (N_3913,N_3741,N_3566);
xor U3914 (N_3914,N_3744,N_3707);
nand U3915 (N_3915,N_3546,N_3739);
xnor U3916 (N_3916,N_3637,N_3593);
and U3917 (N_3917,N_3604,N_3513);
or U3918 (N_3918,N_3656,N_3536);
nor U3919 (N_3919,N_3730,N_3533);
or U3920 (N_3920,N_3671,N_3654);
xnor U3921 (N_3921,N_3514,N_3693);
or U3922 (N_3922,N_3606,N_3673);
xnor U3923 (N_3923,N_3604,N_3629);
nor U3924 (N_3924,N_3546,N_3741);
or U3925 (N_3925,N_3595,N_3710);
and U3926 (N_3926,N_3693,N_3661);
and U3927 (N_3927,N_3661,N_3627);
nand U3928 (N_3928,N_3613,N_3524);
nor U3929 (N_3929,N_3742,N_3507);
xor U3930 (N_3930,N_3601,N_3708);
nand U3931 (N_3931,N_3579,N_3720);
xnor U3932 (N_3932,N_3529,N_3712);
or U3933 (N_3933,N_3655,N_3640);
nor U3934 (N_3934,N_3505,N_3726);
xnor U3935 (N_3935,N_3606,N_3559);
nor U3936 (N_3936,N_3563,N_3604);
or U3937 (N_3937,N_3683,N_3692);
nand U3938 (N_3938,N_3695,N_3513);
nand U3939 (N_3939,N_3675,N_3731);
or U3940 (N_3940,N_3654,N_3634);
nand U3941 (N_3941,N_3575,N_3646);
xnor U3942 (N_3942,N_3632,N_3618);
or U3943 (N_3943,N_3645,N_3614);
nand U3944 (N_3944,N_3611,N_3528);
and U3945 (N_3945,N_3726,N_3733);
nor U3946 (N_3946,N_3741,N_3749);
nor U3947 (N_3947,N_3570,N_3550);
nor U3948 (N_3948,N_3721,N_3504);
xnor U3949 (N_3949,N_3643,N_3594);
xnor U3950 (N_3950,N_3590,N_3654);
nor U3951 (N_3951,N_3677,N_3579);
nor U3952 (N_3952,N_3591,N_3746);
or U3953 (N_3953,N_3733,N_3657);
nand U3954 (N_3954,N_3554,N_3632);
nor U3955 (N_3955,N_3642,N_3700);
xnor U3956 (N_3956,N_3705,N_3507);
nand U3957 (N_3957,N_3650,N_3609);
or U3958 (N_3958,N_3738,N_3642);
and U3959 (N_3959,N_3559,N_3637);
xnor U3960 (N_3960,N_3583,N_3536);
nor U3961 (N_3961,N_3550,N_3519);
or U3962 (N_3962,N_3606,N_3701);
nor U3963 (N_3963,N_3748,N_3582);
nand U3964 (N_3964,N_3526,N_3582);
xor U3965 (N_3965,N_3694,N_3743);
nor U3966 (N_3966,N_3560,N_3614);
nand U3967 (N_3967,N_3554,N_3597);
nand U3968 (N_3968,N_3656,N_3525);
xnor U3969 (N_3969,N_3584,N_3592);
nand U3970 (N_3970,N_3547,N_3608);
or U3971 (N_3971,N_3625,N_3691);
and U3972 (N_3972,N_3704,N_3543);
nand U3973 (N_3973,N_3640,N_3709);
and U3974 (N_3974,N_3500,N_3677);
nand U3975 (N_3975,N_3533,N_3642);
nand U3976 (N_3976,N_3503,N_3507);
or U3977 (N_3977,N_3608,N_3611);
nand U3978 (N_3978,N_3643,N_3690);
or U3979 (N_3979,N_3696,N_3597);
nand U3980 (N_3980,N_3585,N_3599);
nor U3981 (N_3981,N_3705,N_3720);
nor U3982 (N_3982,N_3621,N_3652);
nor U3983 (N_3983,N_3518,N_3596);
or U3984 (N_3984,N_3592,N_3747);
or U3985 (N_3985,N_3728,N_3618);
xnor U3986 (N_3986,N_3637,N_3609);
or U3987 (N_3987,N_3581,N_3610);
xor U3988 (N_3988,N_3594,N_3613);
xor U3989 (N_3989,N_3553,N_3718);
xor U3990 (N_3990,N_3613,N_3612);
nor U3991 (N_3991,N_3605,N_3578);
nand U3992 (N_3992,N_3546,N_3676);
xnor U3993 (N_3993,N_3660,N_3564);
or U3994 (N_3994,N_3569,N_3632);
nand U3995 (N_3995,N_3614,N_3622);
nand U3996 (N_3996,N_3595,N_3736);
or U3997 (N_3997,N_3567,N_3677);
nor U3998 (N_3998,N_3508,N_3536);
nand U3999 (N_3999,N_3511,N_3532);
xnor U4000 (N_4000,N_3854,N_3797);
xor U4001 (N_4001,N_3991,N_3790);
or U4002 (N_4002,N_3807,N_3921);
nand U4003 (N_4003,N_3976,N_3970);
nand U4004 (N_4004,N_3752,N_3924);
nor U4005 (N_4005,N_3905,N_3755);
nor U4006 (N_4006,N_3802,N_3965);
nor U4007 (N_4007,N_3899,N_3968);
nand U4008 (N_4008,N_3986,N_3978);
or U4009 (N_4009,N_3888,N_3915);
nand U4010 (N_4010,N_3935,N_3959);
nand U4011 (N_4011,N_3760,N_3946);
and U4012 (N_4012,N_3814,N_3887);
and U4013 (N_4013,N_3889,N_3766);
and U4014 (N_4014,N_3923,N_3855);
xnor U4015 (N_4015,N_3901,N_3910);
xor U4016 (N_4016,N_3800,N_3780);
or U4017 (N_4017,N_3831,N_3828);
nor U4018 (N_4018,N_3811,N_3999);
or U4019 (N_4019,N_3801,N_3840);
nor U4020 (N_4020,N_3871,N_3988);
nand U4021 (N_4021,N_3989,N_3825);
nand U4022 (N_4022,N_3868,N_3764);
xnor U4023 (N_4023,N_3847,N_3784);
nand U4024 (N_4024,N_3805,N_3884);
nand U4025 (N_4025,N_3974,N_3830);
nor U4026 (N_4026,N_3956,N_3955);
and U4027 (N_4027,N_3757,N_3776);
and U4028 (N_4028,N_3864,N_3866);
or U4029 (N_4029,N_3973,N_3950);
and U4030 (N_4030,N_3917,N_3879);
and U4031 (N_4031,N_3856,N_3853);
and U4032 (N_4032,N_3961,N_3778);
nor U4033 (N_4033,N_3874,N_3931);
nand U4034 (N_4034,N_3803,N_3812);
nor U4035 (N_4035,N_3971,N_3983);
nand U4036 (N_4036,N_3926,N_3966);
nand U4037 (N_4037,N_3779,N_3810);
xnor U4038 (N_4038,N_3785,N_3838);
xor U4039 (N_4039,N_3791,N_3839);
nand U4040 (N_4040,N_3756,N_3827);
or U4041 (N_4041,N_3944,N_3804);
nor U4042 (N_4042,N_3750,N_3891);
xnor U4043 (N_4043,N_3953,N_3775);
xor U4044 (N_4044,N_3957,N_3951);
and U4045 (N_4045,N_3809,N_3904);
nor U4046 (N_4046,N_3943,N_3898);
or U4047 (N_4047,N_3788,N_3796);
nor U4048 (N_4048,N_3967,N_3930);
nor U4049 (N_4049,N_3751,N_3833);
and U4050 (N_4050,N_3857,N_3952);
and U4051 (N_4051,N_3993,N_3977);
or U4052 (N_4052,N_3895,N_3861);
or U4053 (N_4053,N_3858,N_3820);
xor U4054 (N_4054,N_3964,N_3920);
nand U4055 (N_4055,N_3906,N_3997);
or U4056 (N_4056,N_3947,N_3850);
or U4057 (N_4057,N_3945,N_3972);
nor U4058 (N_4058,N_3893,N_3892);
nor U4059 (N_4059,N_3940,N_3794);
nand U4060 (N_4060,N_3815,N_3882);
xnor U4061 (N_4061,N_3938,N_3897);
nand U4062 (N_4062,N_3900,N_3909);
and U4063 (N_4063,N_3948,N_3767);
nor U4064 (N_4064,N_3979,N_3792);
and U4065 (N_4065,N_3937,N_3754);
and U4066 (N_4066,N_3761,N_3782);
or U4067 (N_4067,N_3862,N_3759);
or U4068 (N_4068,N_3992,N_3949);
nor U4069 (N_4069,N_3823,N_3772);
nand U4070 (N_4070,N_3934,N_3995);
or U4071 (N_4071,N_3942,N_3786);
and U4072 (N_4072,N_3819,N_3837);
nor U4073 (N_4073,N_3834,N_3962);
xor U4074 (N_4074,N_3798,N_3762);
and U4075 (N_4075,N_3829,N_3911);
nand U4076 (N_4076,N_3870,N_3922);
nand U4077 (N_4077,N_3984,N_3821);
and U4078 (N_4078,N_3876,N_3769);
or U4079 (N_4079,N_3980,N_3960);
nand U4080 (N_4080,N_3774,N_3771);
and U4081 (N_4081,N_3860,N_3890);
nor U4082 (N_4082,N_3824,N_3982);
nand U4083 (N_4083,N_3913,N_3845);
or U4084 (N_4084,N_3896,N_3996);
nand U4085 (N_4085,N_3975,N_3933);
nor U4086 (N_4086,N_3813,N_3902);
or U4087 (N_4087,N_3885,N_3981);
or U4088 (N_4088,N_3768,N_3765);
nor U4089 (N_4089,N_3877,N_3806);
xor U4090 (N_4090,N_3941,N_3936);
xnor U4091 (N_4091,N_3883,N_3846);
and U4092 (N_4092,N_3954,N_3963);
nand U4093 (N_4093,N_3835,N_3826);
and U4094 (N_4094,N_3886,N_3929);
nand U4095 (N_4095,N_3863,N_3998);
nand U4096 (N_4096,N_3969,N_3851);
xor U4097 (N_4097,N_3808,N_3867);
xor U4098 (N_4098,N_3880,N_3990);
or U4099 (N_4099,N_3770,N_3859);
nand U4100 (N_4100,N_3916,N_3939);
or U4101 (N_4101,N_3908,N_3789);
xnor U4102 (N_4102,N_3894,N_3849);
or U4103 (N_4103,N_3842,N_3918);
xor U4104 (N_4104,N_3994,N_3925);
nor U4105 (N_4105,N_3881,N_3836);
xor U4106 (N_4106,N_3928,N_3832);
xnor U4107 (N_4107,N_3958,N_3841);
or U4108 (N_4108,N_3818,N_3927);
nor U4109 (N_4109,N_3817,N_3793);
nor U4110 (N_4110,N_3843,N_3985);
xnor U4111 (N_4111,N_3987,N_3869);
xor U4112 (N_4112,N_3758,N_3919);
and U4113 (N_4113,N_3903,N_3875);
nor U4114 (N_4114,N_3816,N_3932);
nor U4115 (N_4115,N_3878,N_3763);
or U4116 (N_4116,N_3848,N_3795);
and U4117 (N_4117,N_3781,N_3777);
nor U4118 (N_4118,N_3783,N_3753);
or U4119 (N_4119,N_3822,N_3872);
nand U4120 (N_4120,N_3873,N_3914);
and U4121 (N_4121,N_3907,N_3844);
nor U4122 (N_4122,N_3773,N_3799);
nand U4123 (N_4123,N_3787,N_3865);
nor U4124 (N_4124,N_3852,N_3912);
nor U4125 (N_4125,N_3758,N_3801);
nor U4126 (N_4126,N_3964,N_3941);
or U4127 (N_4127,N_3866,N_3968);
xor U4128 (N_4128,N_3913,N_3839);
xnor U4129 (N_4129,N_3930,N_3984);
or U4130 (N_4130,N_3904,N_3865);
xnor U4131 (N_4131,N_3934,N_3917);
nor U4132 (N_4132,N_3945,N_3790);
nand U4133 (N_4133,N_3894,N_3801);
or U4134 (N_4134,N_3819,N_3857);
and U4135 (N_4135,N_3832,N_3870);
and U4136 (N_4136,N_3930,N_3924);
nor U4137 (N_4137,N_3918,N_3879);
and U4138 (N_4138,N_3868,N_3852);
or U4139 (N_4139,N_3769,N_3998);
xnor U4140 (N_4140,N_3855,N_3762);
or U4141 (N_4141,N_3801,N_3939);
nand U4142 (N_4142,N_3959,N_3963);
xnor U4143 (N_4143,N_3941,N_3846);
nor U4144 (N_4144,N_3903,N_3848);
and U4145 (N_4145,N_3935,N_3879);
or U4146 (N_4146,N_3878,N_3785);
nand U4147 (N_4147,N_3950,N_3884);
nand U4148 (N_4148,N_3777,N_3838);
xnor U4149 (N_4149,N_3885,N_3970);
nand U4150 (N_4150,N_3803,N_3937);
and U4151 (N_4151,N_3931,N_3750);
xnor U4152 (N_4152,N_3825,N_3979);
nor U4153 (N_4153,N_3819,N_3975);
nor U4154 (N_4154,N_3853,N_3758);
and U4155 (N_4155,N_3997,N_3898);
nor U4156 (N_4156,N_3872,N_3784);
nand U4157 (N_4157,N_3776,N_3966);
xor U4158 (N_4158,N_3964,N_3848);
xnor U4159 (N_4159,N_3824,N_3986);
nor U4160 (N_4160,N_3874,N_3891);
nand U4161 (N_4161,N_3758,N_3924);
and U4162 (N_4162,N_3977,N_3800);
or U4163 (N_4163,N_3918,N_3954);
or U4164 (N_4164,N_3975,N_3912);
or U4165 (N_4165,N_3759,N_3975);
xor U4166 (N_4166,N_3927,N_3780);
xor U4167 (N_4167,N_3934,N_3782);
or U4168 (N_4168,N_3803,N_3875);
nor U4169 (N_4169,N_3811,N_3843);
or U4170 (N_4170,N_3950,N_3954);
nand U4171 (N_4171,N_3944,N_3942);
nand U4172 (N_4172,N_3961,N_3879);
nor U4173 (N_4173,N_3799,N_3921);
nor U4174 (N_4174,N_3851,N_3928);
nand U4175 (N_4175,N_3902,N_3878);
and U4176 (N_4176,N_3847,N_3830);
or U4177 (N_4177,N_3860,N_3799);
xor U4178 (N_4178,N_3943,N_3910);
xnor U4179 (N_4179,N_3856,N_3930);
and U4180 (N_4180,N_3786,N_3799);
nand U4181 (N_4181,N_3982,N_3990);
nor U4182 (N_4182,N_3878,N_3895);
or U4183 (N_4183,N_3780,N_3847);
nand U4184 (N_4184,N_3910,N_3968);
or U4185 (N_4185,N_3988,N_3903);
xor U4186 (N_4186,N_3849,N_3951);
or U4187 (N_4187,N_3855,N_3816);
nand U4188 (N_4188,N_3979,N_3894);
nand U4189 (N_4189,N_3898,N_3924);
and U4190 (N_4190,N_3764,N_3949);
or U4191 (N_4191,N_3932,N_3778);
nand U4192 (N_4192,N_3901,N_3955);
nor U4193 (N_4193,N_3906,N_3752);
nor U4194 (N_4194,N_3873,N_3990);
nand U4195 (N_4195,N_3919,N_3885);
xnor U4196 (N_4196,N_3823,N_3952);
xnor U4197 (N_4197,N_3941,N_3811);
xnor U4198 (N_4198,N_3924,N_3969);
or U4199 (N_4199,N_3818,N_3935);
xnor U4200 (N_4200,N_3977,N_3906);
and U4201 (N_4201,N_3761,N_3969);
nand U4202 (N_4202,N_3878,N_3865);
and U4203 (N_4203,N_3980,N_3871);
xor U4204 (N_4204,N_3803,N_3850);
and U4205 (N_4205,N_3784,N_3985);
nand U4206 (N_4206,N_3802,N_3900);
xnor U4207 (N_4207,N_3898,N_3804);
xor U4208 (N_4208,N_3952,N_3759);
xnor U4209 (N_4209,N_3764,N_3769);
xnor U4210 (N_4210,N_3805,N_3842);
and U4211 (N_4211,N_3986,N_3911);
xnor U4212 (N_4212,N_3886,N_3854);
nand U4213 (N_4213,N_3970,N_3926);
xnor U4214 (N_4214,N_3943,N_3893);
or U4215 (N_4215,N_3900,N_3758);
or U4216 (N_4216,N_3961,N_3817);
or U4217 (N_4217,N_3870,N_3836);
and U4218 (N_4218,N_3836,N_3869);
nand U4219 (N_4219,N_3976,N_3826);
or U4220 (N_4220,N_3832,N_3853);
and U4221 (N_4221,N_3950,N_3960);
nand U4222 (N_4222,N_3928,N_3829);
or U4223 (N_4223,N_3769,N_3782);
nor U4224 (N_4224,N_3787,N_3791);
nand U4225 (N_4225,N_3829,N_3852);
xnor U4226 (N_4226,N_3834,N_3873);
nand U4227 (N_4227,N_3839,N_3902);
and U4228 (N_4228,N_3871,N_3984);
and U4229 (N_4229,N_3818,N_3750);
and U4230 (N_4230,N_3826,N_3993);
or U4231 (N_4231,N_3895,N_3885);
nor U4232 (N_4232,N_3771,N_3960);
nand U4233 (N_4233,N_3937,N_3802);
xor U4234 (N_4234,N_3844,N_3764);
or U4235 (N_4235,N_3897,N_3833);
or U4236 (N_4236,N_3913,N_3855);
and U4237 (N_4237,N_3995,N_3868);
nand U4238 (N_4238,N_3906,N_3816);
nand U4239 (N_4239,N_3942,N_3933);
and U4240 (N_4240,N_3942,N_3831);
xor U4241 (N_4241,N_3791,N_3831);
nor U4242 (N_4242,N_3913,N_3831);
or U4243 (N_4243,N_3763,N_3780);
xnor U4244 (N_4244,N_3952,N_3967);
and U4245 (N_4245,N_3847,N_3960);
xnor U4246 (N_4246,N_3929,N_3902);
or U4247 (N_4247,N_3761,N_3786);
nor U4248 (N_4248,N_3757,N_3941);
nor U4249 (N_4249,N_3962,N_3994);
or U4250 (N_4250,N_4035,N_4235);
nor U4251 (N_4251,N_4174,N_4110);
or U4252 (N_4252,N_4147,N_4062);
nand U4253 (N_4253,N_4156,N_4045);
xor U4254 (N_4254,N_4184,N_4221);
or U4255 (N_4255,N_4140,N_4016);
nor U4256 (N_4256,N_4182,N_4172);
or U4257 (N_4257,N_4117,N_4162);
or U4258 (N_4258,N_4055,N_4018);
xnor U4259 (N_4259,N_4158,N_4098);
and U4260 (N_4260,N_4243,N_4080);
or U4261 (N_4261,N_4200,N_4166);
xor U4262 (N_4262,N_4227,N_4027);
or U4263 (N_4263,N_4069,N_4122);
nand U4264 (N_4264,N_4044,N_4099);
nor U4265 (N_4265,N_4116,N_4124);
and U4266 (N_4266,N_4230,N_4036);
nor U4267 (N_4267,N_4161,N_4146);
and U4268 (N_4268,N_4056,N_4176);
xor U4269 (N_4269,N_4127,N_4189);
nand U4270 (N_4270,N_4128,N_4096);
or U4271 (N_4271,N_4178,N_4171);
nand U4272 (N_4272,N_4020,N_4143);
and U4273 (N_4273,N_4012,N_4148);
nand U4274 (N_4274,N_4058,N_4231);
or U4275 (N_4275,N_4113,N_4205);
nor U4276 (N_4276,N_4002,N_4085);
nor U4277 (N_4277,N_4167,N_4152);
or U4278 (N_4278,N_4194,N_4144);
xor U4279 (N_4279,N_4028,N_4212);
and U4280 (N_4280,N_4179,N_4213);
nand U4281 (N_4281,N_4047,N_4219);
xnor U4282 (N_4282,N_4180,N_4188);
or U4283 (N_4283,N_4087,N_4203);
xor U4284 (N_4284,N_4217,N_4070);
nor U4285 (N_4285,N_4092,N_4159);
and U4286 (N_4286,N_4126,N_4223);
xor U4287 (N_4287,N_4014,N_4032);
or U4288 (N_4288,N_4043,N_4195);
nand U4289 (N_4289,N_4086,N_4061);
nor U4290 (N_4290,N_4076,N_4067);
xnor U4291 (N_4291,N_4102,N_4054);
and U4292 (N_4292,N_4063,N_4077);
or U4293 (N_4293,N_4083,N_4071);
nand U4294 (N_4294,N_4081,N_4187);
or U4295 (N_4295,N_4015,N_4109);
nand U4296 (N_4296,N_4193,N_4153);
nand U4297 (N_4297,N_4030,N_4094);
nand U4298 (N_4298,N_4136,N_4238);
or U4299 (N_4299,N_4120,N_4064);
or U4300 (N_4300,N_4079,N_4066);
and U4301 (N_4301,N_4199,N_4100);
and U4302 (N_4302,N_4220,N_4041);
and U4303 (N_4303,N_4134,N_4129);
nor U4304 (N_4304,N_4190,N_4137);
and U4305 (N_4305,N_4068,N_4225);
xnor U4306 (N_4306,N_4097,N_4165);
nand U4307 (N_4307,N_4115,N_4034);
nand U4308 (N_4308,N_4095,N_4224);
xnor U4309 (N_4309,N_4154,N_4057);
nor U4310 (N_4310,N_4025,N_4233);
nand U4311 (N_4311,N_4145,N_4059);
and U4312 (N_4312,N_4218,N_4151);
nand U4313 (N_4313,N_4138,N_4135);
and U4314 (N_4314,N_4021,N_4022);
nor U4315 (N_4315,N_4112,N_4000);
and U4316 (N_4316,N_4239,N_4222);
nor U4317 (N_4317,N_4101,N_4038);
xnor U4318 (N_4318,N_4150,N_4160);
or U4319 (N_4319,N_4084,N_4093);
and U4320 (N_4320,N_4065,N_4164);
or U4321 (N_4321,N_4073,N_4175);
or U4322 (N_4322,N_4111,N_4236);
xnor U4323 (N_4323,N_4001,N_4037);
xnor U4324 (N_4324,N_4209,N_4040);
nor U4325 (N_4325,N_4107,N_4139);
or U4326 (N_4326,N_4060,N_4181);
xnor U4327 (N_4327,N_4170,N_4186);
xnor U4328 (N_4328,N_4123,N_4132);
nor U4329 (N_4329,N_4042,N_4046);
nor U4330 (N_4330,N_4005,N_4078);
nand U4331 (N_4331,N_4248,N_4197);
nand U4332 (N_4332,N_4074,N_4108);
nand U4333 (N_4333,N_4245,N_4052);
and U4334 (N_4334,N_4121,N_4019);
and U4335 (N_4335,N_4249,N_4214);
nand U4336 (N_4336,N_4177,N_4229);
xor U4337 (N_4337,N_4050,N_4119);
nor U4338 (N_4338,N_4017,N_4244);
nor U4339 (N_4339,N_4039,N_4207);
nand U4340 (N_4340,N_4149,N_4211);
nand U4341 (N_4341,N_4168,N_4141);
xnor U4342 (N_4342,N_4206,N_4169);
nand U4343 (N_4343,N_4026,N_4029);
or U4344 (N_4344,N_4088,N_4006);
or U4345 (N_4345,N_4185,N_4163);
nor U4346 (N_4346,N_4173,N_4242);
nand U4347 (N_4347,N_4183,N_4202);
nor U4348 (N_4348,N_4191,N_4226);
or U4349 (N_4349,N_4106,N_4246);
and U4350 (N_4350,N_4023,N_4008);
nor U4351 (N_4351,N_4051,N_4011);
nand U4352 (N_4352,N_4198,N_4192);
xor U4353 (N_4353,N_4247,N_4204);
xnor U4354 (N_4354,N_4082,N_4114);
nor U4355 (N_4355,N_4010,N_4157);
nor U4356 (N_4356,N_4142,N_4075);
and U4357 (N_4357,N_4232,N_4024);
and U4358 (N_4358,N_4234,N_4237);
and U4359 (N_4359,N_4013,N_4240);
nand U4360 (N_4360,N_4155,N_4033);
or U4361 (N_4361,N_4241,N_4049);
or U4362 (N_4362,N_4104,N_4048);
xnor U4363 (N_4363,N_4103,N_4004);
nand U4364 (N_4364,N_4208,N_4133);
nor U4365 (N_4365,N_4118,N_4031);
xor U4366 (N_4366,N_4215,N_4131);
nand U4367 (N_4367,N_4196,N_4210);
or U4368 (N_4368,N_4007,N_4091);
nand U4369 (N_4369,N_4090,N_4053);
nand U4370 (N_4370,N_4009,N_4130);
or U4371 (N_4371,N_4201,N_4072);
nor U4372 (N_4372,N_4228,N_4089);
or U4373 (N_4373,N_4216,N_4003);
nor U4374 (N_4374,N_4105,N_4125);
or U4375 (N_4375,N_4136,N_4222);
and U4376 (N_4376,N_4019,N_4033);
nand U4377 (N_4377,N_4117,N_4243);
nor U4378 (N_4378,N_4092,N_4090);
and U4379 (N_4379,N_4094,N_4027);
xnor U4380 (N_4380,N_4054,N_4161);
xor U4381 (N_4381,N_4083,N_4066);
nand U4382 (N_4382,N_4174,N_4152);
nor U4383 (N_4383,N_4234,N_4112);
nor U4384 (N_4384,N_4107,N_4035);
xnor U4385 (N_4385,N_4045,N_4134);
and U4386 (N_4386,N_4230,N_4203);
nand U4387 (N_4387,N_4217,N_4203);
xnor U4388 (N_4388,N_4086,N_4194);
or U4389 (N_4389,N_4094,N_4111);
xnor U4390 (N_4390,N_4235,N_4058);
and U4391 (N_4391,N_4037,N_4107);
xor U4392 (N_4392,N_4046,N_4247);
xor U4393 (N_4393,N_4157,N_4031);
or U4394 (N_4394,N_4030,N_4217);
nor U4395 (N_4395,N_4101,N_4131);
xor U4396 (N_4396,N_4137,N_4234);
nand U4397 (N_4397,N_4205,N_4005);
nor U4398 (N_4398,N_4049,N_4076);
or U4399 (N_4399,N_4034,N_4219);
xnor U4400 (N_4400,N_4148,N_4226);
nand U4401 (N_4401,N_4017,N_4064);
nor U4402 (N_4402,N_4028,N_4190);
xnor U4403 (N_4403,N_4060,N_4236);
xnor U4404 (N_4404,N_4002,N_4245);
xor U4405 (N_4405,N_4130,N_4087);
and U4406 (N_4406,N_4158,N_4002);
or U4407 (N_4407,N_4126,N_4201);
xnor U4408 (N_4408,N_4162,N_4105);
nor U4409 (N_4409,N_4008,N_4161);
or U4410 (N_4410,N_4089,N_4196);
or U4411 (N_4411,N_4039,N_4231);
nor U4412 (N_4412,N_4139,N_4193);
nand U4413 (N_4413,N_4088,N_4049);
and U4414 (N_4414,N_4063,N_4003);
nor U4415 (N_4415,N_4201,N_4125);
and U4416 (N_4416,N_4047,N_4235);
or U4417 (N_4417,N_4234,N_4139);
or U4418 (N_4418,N_4172,N_4037);
and U4419 (N_4419,N_4220,N_4179);
or U4420 (N_4420,N_4048,N_4151);
nand U4421 (N_4421,N_4038,N_4124);
nand U4422 (N_4422,N_4148,N_4057);
xnor U4423 (N_4423,N_4134,N_4128);
and U4424 (N_4424,N_4223,N_4075);
nor U4425 (N_4425,N_4242,N_4054);
xor U4426 (N_4426,N_4181,N_4090);
or U4427 (N_4427,N_4188,N_4247);
or U4428 (N_4428,N_4094,N_4009);
nand U4429 (N_4429,N_4235,N_4138);
and U4430 (N_4430,N_4170,N_4192);
nand U4431 (N_4431,N_4216,N_4225);
or U4432 (N_4432,N_4045,N_4033);
or U4433 (N_4433,N_4083,N_4139);
nand U4434 (N_4434,N_4200,N_4089);
or U4435 (N_4435,N_4028,N_4128);
nand U4436 (N_4436,N_4057,N_4236);
nor U4437 (N_4437,N_4071,N_4202);
nor U4438 (N_4438,N_4177,N_4086);
xnor U4439 (N_4439,N_4032,N_4116);
and U4440 (N_4440,N_4201,N_4016);
xnor U4441 (N_4441,N_4125,N_4129);
and U4442 (N_4442,N_4214,N_4000);
nor U4443 (N_4443,N_4230,N_4052);
and U4444 (N_4444,N_4031,N_4104);
and U4445 (N_4445,N_4033,N_4000);
xnor U4446 (N_4446,N_4194,N_4042);
nand U4447 (N_4447,N_4064,N_4059);
nand U4448 (N_4448,N_4042,N_4142);
xnor U4449 (N_4449,N_4156,N_4205);
and U4450 (N_4450,N_4087,N_4166);
nand U4451 (N_4451,N_4233,N_4229);
or U4452 (N_4452,N_4103,N_4190);
xor U4453 (N_4453,N_4119,N_4128);
or U4454 (N_4454,N_4202,N_4142);
nand U4455 (N_4455,N_4147,N_4080);
nand U4456 (N_4456,N_4227,N_4176);
nor U4457 (N_4457,N_4235,N_4076);
and U4458 (N_4458,N_4212,N_4015);
and U4459 (N_4459,N_4166,N_4142);
nor U4460 (N_4460,N_4089,N_4204);
xnor U4461 (N_4461,N_4159,N_4207);
or U4462 (N_4462,N_4216,N_4184);
nand U4463 (N_4463,N_4004,N_4210);
or U4464 (N_4464,N_4191,N_4160);
or U4465 (N_4465,N_4156,N_4087);
xor U4466 (N_4466,N_4076,N_4020);
nand U4467 (N_4467,N_4247,N_4027);
and U4468 (N_4468,N_4184,N_4191);
and U4469 (N_4469,N_4013,N_4067);
xor U4470 (N_4470,N_4047,N_4092);
xor U4471 (N_4471,N_4013,N_4206);
xor U4472 (N_4472,N_4248,N_4171);
xor U4473 (N_4473,N_4190,N_4116);
or U4474 (N_4474,N_4110,N_4216);
or U4475 (N_4475,N_4154,N_4130);
xor U4476 (N_4476,N_4092,N_4158);
or U4477 (N_4477,N_4029,N_4129);
nand U4478 (N_4478,N_4104,N_4123);
nand U4479 (N_4479,N_4079,N_4030);
xnor U4480 (N_4480,N_4011,N_4239);
and U4481 (N_4481,N_4134,N_4048);
nor U4482 (N_4482,N_4087,N_4190);
and U4483 (N_4483,N_4034,N_4164);
nand U4484 (N_4484,N_4248,N_4145);
or U4485 (N_4485,N_4017,N_4055);
or U4486 (N_4486,N_4098,N_4205);
and U4487 (N_4487,N_4030,N_4199);
nand U4488 (N_4488,N_4040,N_4242);
and U4489 (N_4489,N_4126,N_4208);
nand U4490 (N_4490,N_4147,N_4246);
xnor U4491 (N_4491,N_4140,N_4170);
or U4492 (N_4492,N_4184,N_4104);
or U4493 (N_4493,N_4076,N_4220);
xor U4494 (N_4494,N_4087,N_4207);
nand U4495 (N_4495,N_4110,N_4155);
nor U4496 (N_4496,N_4066,N_4091);
or U4497 (N_4497,N_4046,N_4179);
xnor U4498 (N_4498,N_4059,N_4219);
nand U4499 (N_4499,N_4153,N_4059);
xor U4500 (N_4500,N_4457,N_4441);
nand U4501 (N_4501,N_4292,N_4384);
nor U4502 (N_4502,N_4493,N_4321);
nand U4503 (N_4503,N_4456,N_4461);
xor U4504 (N_4504,N_4278,N_4403);
nand U4505 (N_4505,N_4322,N_4317);
xnor U4506 (N_4506,N_4395,N_4458);
xor U4507 (N_4507,N_4365,N_4432);
nor U4508 (N_4508,N_4446,N_4258);
xnor U4509 (N_4509,N_4295,N_4468);
and U4510 (N_4510,N_4499,N_4439);
nand U4511 (N_4511,N_4283,N_4455);
nor U4512 (N_4512,N_4336,N_4299);
and U4513 (N_4513,N_4472,N_4352);
nor U4514 (N_4514,N_4325,N_4318);
or U4515 (N_4515,N_4451,N_4261);
nor U4516 (N_4516,N_4427,N_4443);
xor U4517 (N_4517,N_4313,N_4356);
and U4518 (N_4518,N_4492,N_4447);
nor U4519 (N_4519,N_4320,N_4355);
nand U4520 (N_4520,N_4288,N_4474);
and U4521 (N_4521,N_4297,N_4342);
xnor U4522 (N_4522,N_4467,N_4453);
xnor U4523 (N_4523,N_4268,N_4480);
or U4524 (N_4524,N_4280,N_4300);
nand U4525 (N_4525,N_4359,N_4285);
or U4526 (N_4526,N_4481,N_4330);
nor U4527 (N_4527,N_4296,N_4362);
nand U4528 (N_4528,N_4364,N_4314);
nor U4529 (N_4529,N_4389,N_4390);
and U4530 (N_4530,N_4411,N_4361);
and U4531 (N_4531,N_4282,N_4404);
xnor U4532 (N_4532,N_4399,N_4331);
or U4533 (N_4533,N_4406,N_4375);
and U4534 (N_4534,N_4351,N_4421);
xor U4535 (N_4535,N_4339,N_4327);
nor U4536 (N_4536,N_4440,N_4435);
nand U4537 (N_4537,N_4332,N_4425);
and U4538 (N_4538,N_4279,N_4289);
and U4539 (N_4539,N_4445,N_4433);
or U4540 (N_4540,N_4496,N_4312);
or U4541 (N_4541,N_4298,N_4482);
or U4542 (N_4542,N_4415,N_4388);
nand U4543 (N_4543,N_4442,N_4418);
and U4544 (N_4544,N_4497,N_4437);
or U4545 (N_4545,N_4402,N_4464);
or U4546 (N_4546,N_4469,N_4477);
xor U4547 (N_4547,N_4274,N_4329);
or U4548 (N_4548,N_4428,N_4422);
nor U4549 (N_4549,N_4408,N_4378);
or U4550 (N_4550,N_4264,N_4387);
xnor U4551 (N_4551,N_4392,N_4346);
and U4552 (N_4552,N_4273,N_4368);
nor U4553 (N_4553,N_4462,N_4251);
or U4554 (N_4554,N_4423,N_4444);
nand U4555 (N_4555,N_4271,N_4385);
nand U4556 (N_4556,N_4483,N_4269);
or U4557 (N_4557,N_4380,N_4347);
xnor U4558 (N_4558,N_4250,N_4405);
nand U4559 (N_4559,N_4372,N_4391);
nor U4560 (N_4560,N_4484,N_4479);
xor U4561 (N_4561,N_4256,N_4454);
nor U4562 (N_4562,N_4284,N_4383);
xor U4563 (N_4563,N_4373,N_4489);
and U4564 (N_4564,N_4315,N_4307);
nand U4565 (N_4565,N_4323,N_4379);
xor U4566 (N_4566,N_4255,N_4253);
or U4567 (N_4567,N_4302,N_4294);
and U4568 (N_4568,N_4449,N_4358);
nor U4569 (N_4569,N_4293,N_4376);
or U4570 (N_4570,N_4267,N_4337);
or U4571 (N_4571,N_4400,N_4326);
or U4572 (N_4572,N_4491,N_4354);
xnor U4573 (N_4573,N_4290,N_4448);
and U4574 (N_4574,N_4487,N_4270);
or U4575 (N_4575,N_4398,N_4420);
nor U4576 (N_4576,N_4377,N_4305);
and U4577 (N_4577,N_4475,N_4452);
nor U4578 (N_4578,N_4419,N_4338);
nor U4579 (N_4579,N_4360,N_4429);
nand U4580 (N_4580,N_4396,N_4438);
and U4581 (N_4581,N_4486,N_4465);
xor U4582 (N_4582,N_4343,N_4345);
nand U4583 (N_4583,N_4357,N_4324);
and U4584 (N_4584,N_4369,N_4450);
nor U4585 (N_4585,N_4281,N_4308);
nand U4586 (N_4586,N_4431,N_4416);
or U4587 (N_4587,N_4350,N_4485);
nor U4588 (N_4588,N_4311,N_4410);
nor U4589 (N_4589,N_4263,N_4303);
nor U4590 (N_4590,N_4490,N_4494);
or U4591 (N_4591,N_4426,N_4488);
or U4592 (N_4592,N_4382,N_4417);
or U4593 (N_4593,N_4353,N_4463);
or U4594 (N_4594,N_4401,N_4265);
nor U4595 (N_4595,N_4252,N_4367);
and U4596 (N_4596,N_4257,N_4319);
xnor U4597 (N_4597,N_4309,N_4287);
xnor U4598 (N_4598,N_4407,N_4371);
nand U4599 (N_4599,N_4478,N_4344);
or U4600 (N_4600,N_4272,N_4413);
and U4601 (N_4601,N_4473,N_4276);
xnor U4602 (N_4602,N_4277,N_4460);
and U4603 (N_4603,N_4260,N_4341);
nor U4604 (N_4604,N_4306,N_4381);
nand U4605 (N_4605,N_4335,N_4495);
xor U4606 (N_4606,N_4340,N_4412);
nand U4607 (N_4607,N_4316,N_4397);
and U4608 (N_4608,N_4262,N_4363);
nor U4609 (N_4609,N_4291,N_4259);
xnor U4610 (N_4610,N_4334,N_4430);
and U4611 (N_4611,N_4498,N_4301);
nor U4612 (N_4612,N_4436,N_4349);
and U4613 (N_4613,N_4366,N_4275);
nand U4614 (N_4614,N_4254,N_4459);
nand U4615 (N_4615,N_4348,N_4470);
and U4616 (N_4616,N_4374,N_4328);
nand U4617 (N_4617,N_4266,N_4386);
xnor U4618 (N_4618,N_4333,N_4476);
nor U4619 (N_4619,N_4394,N_4466);
and U4620 (N_4620,N_4409,N_4310);
nand U4621 (N_4621,N_4286,N_4414);
xor U4622 (N_4622,N_4304,N_4393);
xnor U4623 (N_4623,N_4471,N_4434);
nand U4624 (N_4624,N_4370,N_4424);
and U4625 (N_4625,N_4382,N_4487);
nor U4626 (N_4626,N_4420,N_4299);
xor U4627 (N_4627,N_4288,N_4307);
and U4628 (N_4628,N_4327,N_4477);
nor U4629 (N_4629,N_4313,N_4469);
or U4630 (N_4630,N_4317,N_4461);
xor U4631 (N_4631,N_4313,N_4316);
and U4632 (N_4632,N_4279,N_4472);
and U4633 (N_4633,N_4288,N_4436);
nor U4634 (N_4634,N_4377,N_4463);
or U4635 (N_4635,N_4398,N_4426);
nor U4636 (N_4636,N_4326,N_4375);
xor U4637 (N_4637,N_4429,N_4286);
or U4638 (N_4638,N_4327,N_4475);
or U4639 (N_4639,N_4285,N_4283);
or U4640 (N_4640,N_4378,N_4477);
or U4641 (N_4641,N_4473,N_4336);
nand U4642 (N_4642,N_4414,N_4441);
or U4643 (N_4643,N_4314,N_4310);
and U4644 (N_4644,N_4384,N_4251);
nor U4645 (N_4645,N_4336,N_4396);
and U4646 (N_4646,N_4305,N_4468);
xor U4647 (N_4647,N_4379,N_4461);
xnor U4648 (N_4648,N_4286,N_4263);
nand U4649 (N_4649,N_4463,N_4369);
or U4650 (N_4650,N_4304,N_4433);
xnor U4651 (N_4651,N_4403,N_4498);
xnor U4652 (N_4652,N_4395,N_4320);
nand U4653 (N_4653,N_4256,N_4339);
and U4654 (N_4654,N_4494,N_4375);
nand U4655 (N_4655,N_4370,N_4290);
and U4656 (N_4656,N_4496,N_4317);
or U4657 (N_4657,N_4322,N_4395);
and U4658 (N_4658,N_4420,N_4268);
or U4659 (N_4659,N_4353,N_4286);
nor U4660 (N_4660,N_4355,N_4455);
or U4661 (N_4661,N_4401,N_4296);
nor U4662 (N_4662,N_4332,N_4393);
xnor U4663 (N_4663,N_4256,N_4497);
xnor U4664 (N_4664,N_4407,N_4355);
nand U4665 (N_4665,N_4250,N_4263);
nor U4666 (N_4666,N_4476,N_4277);
or U4667 (N_4667,N_4434,N_4435);
or U4668 (N_4668,N_4358,N_4375);
nand U4669 (N_4669,N_4337,N_4283);
xor U4670 (N_4670,N_4362,N_4423);
nand U4671 (N_4671,N_4458,N_4280);
nand U4672 (N_4672,N_4391,N_4263);
nor U4673 (N_4673,N_4330,N_4332);
nand U4674 (N_4674,N_4365,N_4320);
nor U4675 (N_4675,N_4291,N_4280);
and U4676 (N_4676,N_4408,N_4488);
or U4677 (N_4677,N_4253,N_4367);
and U4678 (N_4678,N_4452,N_4370);
nand U4679 (N_4679,N_4468,N_4335);
nor U4680 (N_4680,N_4349,N_4285);
xor U4681 (N_4681,N_4462,N_4467);
or U4682 (N_4682,N_4470,N_4463);
and U4683 (N_4683,N_4404,N_4350);
and U4684 (N_4684,N_4382,N_4437);
and U4685 (N_4685,N_4267,N_4334);
nor U4686 (N_4686,N_4303,N_4432);
and U4687 (N_4687,N_4412,N_4327);
or U4688 (N_4688,N_4286,N_4296);
or U4689 (N_4689,N_4489,N_4466);
nand U4690 (N_4690,N_4493,N_4469);
nand U4691 (N_4691,N_4395,N_4266);
xnor U4692 (N_4692,N_4306,N_4307);
or U4693 (N_4693,N_4386,N_4337);
nand U4694 (N_4694,N_4258,N_4443);
or U4695 (N_4695,N_4350,N_4300);
nor U4696 (N_4696,N_4487,N_4459);
and U4697 (N_4697,N_4366,N_4445);
nand U4698 (N_4698,N_4359,N_4380);
and U4699 (N_4699,N_4463,N_4324);
and U4700 (N_4700,N_4283,N_4326);
or U4701 (N_4701,N_4435,N_4416);
nor U4702 (N_4702,N_4301,N_4475);
nand U4703 (N_4703,N_4321,N_4426);
and U4704 (N_4704,N_4299,N_4267);
nand U4705 (N_4705,N_4275,N_4314);
xor U4706 (N_4706,N_4320,N_4324);
xnor U4707 (N_4707,N_4497,N_4349);
nand U4708 (N_4708,N_4396,N_4472);
xor U4709 (N_4709,N_4408,N_4384);
and U4710 (N_4710,N_4412,N_4428);
nand U4711 (N_4711,N_4450,N_4458);
nor U4712 (N_4712,N_4277,N_4470);
and U4713 (N_4713,N_4383,N_4312);
nor U4714 (N_4714,N_4470,N_4421);
xor U4715 (N_4715,N_4426,N_4250);
nand U4716 (N_4716,N_4333,N_4337);
xor U4717 (N_4717,N_4377,N_4362);
or U4718 (N_4718,N_4476,N_4456);
and U4719 (N_4719,N_4331,N_4318);
or U4720 (N_4720,N_4332,N_4460);
and U4721 (N_4721,N_4413,N_4456);
nor U4722 (N_4722,N_4465,N_4440);
or U4723 (N_4723,N_4485,N_4340);
and U4724 (N_4724,N_4491,N_4302);
or U4725 (N_4725,N_4391,N_4428);
nand U4726 (N_4726,N_4437,N_4361);
nand U4727 (N_4727,N_4253,N_4458);
xor U4728 (N_4728,N_4455,N_4486);
nand U4729 (N_4729,N_4327,N_4250);
or U4730 (N_4730,N_4324,N_4312);
and U4731 (N_4731,N_4329,N_4256);
xnor U4732 (N_4732,N_4310,N_4357);
or U4733 (N_4733,N_4371,N_4457);
nor U4734 (N_4734,N_4481,N_4462);
nand U4735 (N_4735,N_4372,N_4427);
nand U4736 (N_4736,N_4416,N_4482);
nor U4737 (N_4737,N_4362,N_4486);
nand U4738 (N_4738,N_4322,N_4451);
and U4739 (N_4739,N_4317,N_4468);
and U4740 (N_4740,N_4399,N_4349);
nor U4741 (N_4741,N_4312,N_4428);
xor U4742 (N_4742,N_4386,N_4400);
xor U4743 (N_4743,N_4255,N_4432);
or U4744 (N_4744,N_4266,N_4415);
or U4745 (N_4745,N_4342,N_4395);
and U4746 (N_4746,N_4431,N_4326);
nand U4747 (N_4747,N_4417,N_4341);
nor U4748 (N_4748,N_4339,N_4402);
nand U4749 (N_4749,N_4436,N_4407);
nor U4750 (N_4750,N_4567,N_4616);
nand U4751 (N_4751,N_4623,N_4644);
and U4752 (N_4752,N_4716,N_4631);
nor U4753 (N_4753,N_4640,N_4678);
xor U4754 (N_4754,N_4513,N_4683);
or U4755 (N_4755,N_4564,N_4520);
nand U4756 (N_4756,N_4516,N_4674);
nand U4757 (N_4757,N_4703,N_4585);
or U4758 (N_4758,N_4609,N_4548);
and U4759 (N_4759,N_4613,N_4663);
xnor U4760 (N_4760,N_4688,N_4582);
and U4761 (N_4761,N_4610,N_4675);
nand U4762 (N_4762,N_4671,N_4638);
xnor U4763 (N_4763,N_4555,N_4518);
nand U4764 (N_4764,N_4619,N_4690);
or U4765 (N_4765,N_4509,N_4627);
nor U4766 (N_4766,N_4649,N_4536);
or U4767 (N_4767,N_4707,N_4723);
xor U4768 (N_4768,N_4679,N_4658);
xnor U4769 (N_4769,N_4684,N_4522);
or U4770 (N_4770,N_4738,N_4664);
or U4771 (N_4771,N_4657,N_4622);
or U4772 (N_4772,N_4546,N_4540);
xnor U4773 (N_4773,N_4572,N_4532);
nand U4774 (N_4774,N_4511,N_4550);
or U4775 (N_4775,N_4709,N_4704);
or U4776 (N_4776,N_4605,N_4660);
nor U4777 (N_4777,N_4632,N_4641);
and U4778 (N_4778,N_4521,N_4538);
xor U4779 (N_4779,N_4625,N_4662);
nand U4780 (N_4780,N_4599,N_4576);
and U4781 (N_4781,N_4570,N_4504);
or U4782 (N_4782,N_4621,N_4677);
or U4783 (N_4783,N_4587,N_4589);
and U4784 (N_4784,N_4584,N_4552);
xnor U4785 (N_4785,N_4526,N_4531);
and U4786 (N_4786,N_4730,N_4724);
nor U4787 (N_4787,N_4544,N_4598);
or U4788 (N_4788,N_4732,N_4728);
nor U4789 (N_4789,N_4642,N_4514);
and U4790 (N_4790,N_4545,N_4594);
nand U4791 (N_4791,N_4593,N_4527);
or U4792 (N_4792,N_4528,N_4517);
nor U4793 (N_4793,N_4530,N_4571);
or U4794 (N_4794,N_4557,N_4636);
xnor U4795 (N_4795,N_4726,N_4574);
and U4796 (N_4796,N_4681,N_4612);
or U4797 (N_4797,N_4601,N_4706);
xnor U4798 (N_4798,N_4596,N_4523);
xnor U4799 (N_4799,N_4718,N_4624);
or U4800 (N_4800,N_4680,N_4586);
and U4801 (N_4801,N_4692,N_4719);
nand U4802 (N_4802,N_4676,N_4534);
nor U4803 (N_4803,N_4553,N_4620);
nor U4804 (N_4804,N_4629,N_4592);
xnor U4805 (N_4805,N_4600,N_4727);
nand U4806 (N_4806,N_4578,N_4645);
and U4807 (N_4807,N_4700,N_4618);
or U4808 (N_4808,N_4687,N_4670);
nor U4809 (N_4809,N_4734,N_4502);
xor U4810 (N_4810,N_4506,N_4560);
xor U4811 (N_4811,N_4659,N_4669);
nor U4812 (N_4812,N_4542,N_4501);
nor U4813 (N_4813,N_4666,N_4746);
xor U4814 (N_4814,N_4741,N_4736);
and U4815 (N_4815,N_4614,N_4583);
or U4816 (N_4816,N_4568,N_4512);
nand U4817 (N_4817,N_4712,N_4708);
nor U4818 (N_4818,N_4533,N_4561);
nor U4819 (N_4819,N_4588,N_4591);
and U4820 (N_4820,N_4643,N_4569);
and U4821 (N_4821,N_4733,N_4604);
xnor U4822 (N_4822,N_4529,N_4731);
nand U4823 (N_4823,N_4737,N_4580);
nand U4824 (N_4824,N_4717,N_4720);
xnor U4825 (N_4825,N_4710,N_4699);
nand U4826 (N_4826,N_4559,N_4749);
nand U4827 (N_4827,N_4646,N_4668);
nor U4828 (N_4828,N_4654,N_4608);
or U4829 (N_4829,N_4606,N_4505);
or U4830 (N_4830,N_4515,N_4508);
or U4831 (N_4831,N_4639,N_4597);
xnor U4832 (N_4832,N_4551,N_4558);
nand U4833 (N_4833,N_4693,N_4661);
or U4834 (N_4834,N_4653,N_4740);
nand U4835 (N_4835,N_4696,N_4650);
nor U4836 (N_4836,N_4739,N_4607);
nand U4837 (N_4837,N_4682,N_4547);
or U4838 (N_4838,N_4519,N_4603);
xnor U4839 (N_4839,N_4535,N_4563);
nand U4840 (N_4840,N_4573,N_4510);
xnor U4841 (N_4841,N_4565,N_4626);
nand U4842 (N_4842,N_4617,N_4655);
xor U4843 (N_4843,N_4702,N_4637);
or U4844 (N_4844,N_4579,N_4748);
xnor U4845 (N_4845,N_4525,N_4694);
nor U4846 (N_4846,N_4500,N_4651);
or U4847 (N_4847,N_4652,N_4685);
nor U4848 (N_4848,N_4747,N_4566);
and U4849 (N_4849,N_4647,N_4581);
nand U4850 (N_4850,N_4722,N_4543);
xor U4851 (N_4851,N_4634,N_4729);
xor U4852 (N_4852,N_4672,N_4721);
nand U4853 (N_4853,N_4615,N_4745);
nor U4854 (N_4854,N_4667,N_4507);
or U4855 (N_4855,N_4630,N_4656);
nor U4856 (N_4856,N_4744,N_4673);
nand U4857 (N_4857,N_4698,N_4714);
and U4858 (N_4858,N_4695,N_4715);
nand U4859 (N_4859,N_4701,N_4602);
nand U4860 (N_4860,N_4713,N_4742);
nor U4861 (N_4861,N_4735,N_4562);
or U4862 (N_4862,N_4691,N_4590);
xnor U4863 (N_4863,N_4611,N_4633);
nand U4864 (N_4864,N_4628,N_4697);
nand U4865 (N_4865,N_4539,N_4689);
nor U4866 (N_4866,N_4554,N_4711);
or U4867 (N_4867,N_4541,N_4686);
xnor U4868 (N_4868,N_4665,N_4705);
and U4869 (N_4869,N_4577,N_4524);
or U4870 (N_4870,N_4549,N_4648);
nand U4871 (N_4871,N_4725,N_4537);
xor U4872 (N_4872,N_4635,N_4503);
nand U4873 (N_4873,N_4595,N_4743);
nor U4874 (N_4874,N_4575,N_4556);
or U4875 (N_4875,N_4676,N_4594);
or U4876 (N_4876,N_4722,N_4573);
nor U4877 (N_4877,N_4554,N_4697);
nand U4878 (N_4878,N_4557,N_4640);
or U4879 (N_4879,N_4554,N_4611);
nor U4880 (N_4880,N_4592,N_4624);
nor U4881 (N_4881,N_4637,N_4515);
nand U4882 (N_4882,N_4584,N_4721);
nor U4883 (N_4883,N_4543,N_4628);
xnor U4884 (N_4884,N_4732,N_4651);
and U4885 (N_4885,N_4683,N_4530);
and U4886 (N_4886,N_4653,N_4532);
nor U4887 (N_4887,N_4561,N_4682);
or U4888 (N_4888,N_4547,N_4691);
xnor U4889 (N_4889,N_4672,N_4649);
xor U4890 (N_4890,N_4590,N_4630);
xnor U4891 (N_4891,N_4545,N_4738);
nor U4892 (N_4892,N_4649,N_4682);
nor U4893 (N_4893,N_4729,N_4505);
or U4894 (N_4894,N_4710,N_4557);
xnor U4895 (N_4895,N_4528,N_4513);
and U4896 (N_4896,N_4528,N_4504);
nand U4897 (N_4897,N_4657,N_4523);
nand U4898 (N_4898,N_4649,N_4633);
nand U4899 (N_4899,N_4683,N_4535);
and U4900 (N_4900,N_4703,N_4619);
nand U4901 (N_4901,N_4565,N_4604);
xnor U4902 (N_4902,N_4526,N_4684);
nand U4903 (N_4903,N_4699,N_4662);
and U4904 (N_4904,N_4742,N_4511);
nand U4905 (N_4905,N_4664,N_4714);
xor U4906 (N_4906,N_4635,N_4740);
or U4907 (N_4907,N_4536,N_4660);
nor U4908 (N_4908,N_4735,N_4694);
nor U4909 (N_4909,N_4537,N_4649);
nand U4910 (N_4910,N_4539,N_4709);
xor U4911 (N_4911,N_4606,N_4642);
or U4912 (N_4912,N_4526,N_4650);
and U4913 (N_4913,N_4746,N_4710);
nand U4914 (N_4914,N_4670,N_4627);
or U4915 (N_4915,N_4740,N_4697);
xor U4916 (N_4916,N_4562,N_4548);
xnor U4917 (N_4917,N_4634,N_4509);
or U4918 (N_4918,N_4607,N_4738);
nor U4919 (N_4919,N_4507,N_4508);
and U4920 (N_4920,N_4546,N_4574);
nor U4921 (N_4921,N_4655,N_4593);
nand U4922 (N_4922,N_4748,N_4583);
or U4923 (N_4923,N_4604,N_4576);
nor U4924 (N_4924,N_4540,N_4634);
and U4925 (N_4925,N_4501,N_4584);
xor U4926 (N_4926,N_4693,N_4730);
nand U4927 (N_4927,N_4577,N_4738);
and U4928 (N_4928,N_4718,N_4725);
nand U4929 (N_4929,N_4652,N_4542);
or U4930 (N_4930,N_4512,N_4733);
xnor U4931 (N_4931,N_4505,N_4735);
or U4932 (N_4932,N_4691,N_4697);
nand U4933 (N_4933,N_4513,N_4638);
nand U4934 (N_4934,N_4745,N_4623);
or U4935 (N_4935,N_4519,N_4749);
or U4936 (N_4936,N_4723,N_4612);
xnor U4937 (N_4937,N_4612,N_4652);
nand U4938 (N_4938,N_4529,N_4577);
nand U4939 (N_4939,N_4578,N_4547);
or U4940 (N_4940,N_4641,N_4569);
nand U4941 (N_4941,N_4728,N_4537);
xnor U4942 (N_4942,N_4518,N_4587);
xnor U4943 (N_4943,N_4608,N_4596);
and U4944 (N_4944,N_4580,N_4577);
nor U4945 (N_4945,N_4643,N_4616);
and U4946 (N_4946,N_4654,N_4602);
and U4947 (N_4947,N_4620,N_4509);
xnor U4948 (N_4948,N_4711,N_4532);
nand U4949 (N_4949,N_4660,N_4570);
nor U4950 (N_4950,N_4511,N_4725);
nand U4951 (N_4951,N_4667,N_4690);
nand U4952 (N_4952,N_4570,N_4723);
xnor U4953 (N_4953,N_4551,N_4554);
nand U4954 (N_4954,N_4654,N_4626);
or U4955 (N_4955,N_4664,N_4571);
and U4956 (N_4956,N_4552,N_4697);
nor U4957 (N_4957,N_4518,N_4502);
nand U4958 (N_4958,N_4704,N_4660);
nor U4959 (N_4959,N_4667,N_4609);
or U4960 (N_4960,N_4536,N_4626);
or U4961 (N_4961,N_4727,N_4591);
or U4962 (N_4962,N_4548,N_4661);
or U4963 (N_4963,N_4552,N_4587);
and U4964 (N_4964,N_4602,N_4691);
nor U4965 (N_4965,N_4679,N_4564);
nor U4966 (N_4966,N_4722,N_4528);
nor U4967 (N_4967,N_4583,N_4659);
xnor U4968 (N_4968,N_4696,N_4691);
nor U4969 (N_4969,N_4564,N_4619);
xnor U4970 (N_4970,N_4574,N_4700);
nand U4971 (N_4971,N_4622,N_4539);
and U4972 (N_4972,N_4742,N_4613);
xor U4973 (N_4973,N_4621,N_4723);
nor U4974 (N_4974,N_4746,N_4717);
nand U4975 (N_4975,N_4510,N_4582);
nor U4976 (N_4976,N_4735,N_4507);
or U4977 (N_4977,N_4522,N_4625);
nand U4978 (N_4978,N_4561,N_4583);
nand U4979 (N_4979,N_4520,N_4673);
or U4980 (N_4980,N_4518,N_4651);
and U4981 (N_4981,N_4567,N_4593);
xnor U4982 (N_4982,N_4657,N_4733);
nand U4983 (N_4983,N_4695,N_4501);
nor U4984 (N_4984,N_4640,N_4505);
nand U4985 (N_4985,N_4580,N_4518);
nand U4986 (N_4986,N_4691,N_4597);
nand U4987 (N_4987,N_4637,N_4689);
or U4988 (N_4988,N_4576,N_4506);
and U4989 (N_4989,N_4507,N_4590);
xnor U4990 (N_4990,N_4731,N_4745);
and U4991 (N_4991,N_4566,N_4704);
and U4992 (N_4992,N_4553,N_4712);
nand U4993 (N_4993,N_4612,N_4702);
nor U4994 (N_4994,N_4690,N_4551);
and U4995 (N_4995,N_4592,N_4724);
or U4996 (N_4996,N_4630,N_4597);
and U4997 (N_4997,N_4634,N_4617);
nand U4998 (N_4998,N_4623,N_4702);
nor U4999 (N_4999,N_4581,N_4714);
nand U5000 (N_5000,N_4990,N_4777);
xnor U5001 (N_5001,N_4783,N_4976);
xor U5002 (N_5002,N_4839,N_4863);
nand U5003 (N_5003,N_4834,N_4803);
xnor U5004 (N_5004,N_4984,N_4903);
or U5005 (N_5005,N_4944,N_4751);
or U5006 (N_5006,N_4757,N_4991);
or U5007 (N_5007,N_4812,N_4847);
xor U5008 (N_5008,N_4924,N_4987);
nor U5009 (N_5009,N_4951,N_4770);
nor U5010 (N_5010,N_4888,N_4977);
and U5011 (N_5011,N_4880,N_4796);
or U5012 (N_5012,N_4811,N_4848);
xor U5013 (N_5013,N_4845,N_4877);
or U5014 (N_5014,N_4829,N_4993);
nand U5015 (N_5015,N_4822,N_4872);
xnor U5016 (N_5016,N_4780,N_4909);
nor U5017 (N_5017,N_4755,N_4809);
nand U5018 (N_5018,N_4907,N_4833);
or U5019 (N_5019,N_4900,N_4767);
xnor U5020 (N_5020,N_4801,N_4805);
nor U5021 (N_5021,N_4896,N_4831);
and U5022 (N_5022,N_4952,N_4938);
or U5023 (N_5023,N_4788,N_4855);
nor U5024 (N_5024,N_4943,N_4852);
nand U5025 (N_5025,N_4949,N_4979);
or U5026 (N_5026,N_4956,N_4857);
and U5027 (N_5027,N_4786,N_4925);
or U5028 (N_5028,N_4981,N_4864);
and U5029 (N_5029,N_4887,N_4935);
nor U5030 (N_5030,N_4772,N_4816);
and U5031 (N_5031,N_4970,N_4837);
and U5032 (N_5032,N_4911,N_4775);
nand U5033 (N_5033,N_4937,N_4761);
and U5034 (N_5034,N_4930,N_4893);
nor U5035 (N_5035,N_4769,N_4969);
nor U5036 (N_5036,N_4750,N_4844);
and U5037 (N_5037,N_4905,N_4760);
or U5038 (N_5038,N_4778,N_4955);
or U5039 (N_5039,N_4752,N_4840);
nand U5040 (N_5040,N_4994,N_4957);
and U5041 (N_5041,N_4912,N_4860);
and U5042 (N_5042,N_4842,N_4975);
and U5043 (N_5043,N_4895,N_4963);
and U5044 (N_5044,N_4997,N_4879);
nand U5045 (N_5045,N_4869,N_4826);
nor U5046 (N_5046,N_4794,N_4962);
and U5047 (N_5047,N_4933,N_4968);
xnor U5048 (N_5048,N_4914,N_4960);
and U5049 (N_5049,N_4898,N_4908);
nor U5050 (N_5050,N_4807,N_4862);
nor U5051 (N_5051,N_4858,N_4874);
or U5052 (N_5052,N_4978,N_4929);
or U5053 (N_5053,N_4791,N_4999);
xnor U5054 (N_5054,N_4759,N_4841);
and U5055 (N_5055,N_4823,N_4771);
nand U5056 (N_5056,N_4779,N_4815);
and U5057 (N_5057,N_4921,N_4890);
nand U5058 (N_5058,N_4817,N_4953);
nor U5059 (N_5059,N_4828,N_4787);
nor U5060 (N_5060,N_4868,N_4998);
nand U5061 (N_5061,N_4849,N_4884);
nor U5062 (N_5062,N_4942,N_4982);
and U5063 (N_5063,N_4753,N_4931);
or U5064 (N_5064,N_4902,N_4870);
nand U5065 (N_5065,N_4934,N_4913);
nor U5066 (N_5066,N_4756,N_4790);
xor U5067 (N_5067,N_4776,N_4859);
xnor U5068 (N_5068,N_4873,N_4850);
nor U5069 (N_5069,N_4785,N_4853);
nor U5070 (N_5070,N_4838,N_4765);
nand U5071 (N_5071,N_4806,N_4854);
and U5072 (N_5072,N_4797,N_4856);
or U5073 (N_5073,N_4886,N_4795);
xnor U5074 (N_5074,N_4892,N_4989);
xnor U5075 (N_5075,N_4971,N_4808);
nor U5076 (N_5076,N_4945,N_4950);
and U5077 (N_5077,N_4926,N_4940);
nand U5078 (N_5078,N_4941,N_4851);
and U5079 (N_5079,N_4782,N_4897);
nor U5080 (N_5080,N_4954,N_4766);
nor U5081 (N_5081,N_4784,N_4818);
or U5082 (N_5082,N_4899,N_4825);
and U5083 (N_5083,N_4959,N_4754);
and U5084 (N_5084,N_4804,N_4768);
and U5085 (N_5085,N_4821,N_4813);
nor U5086 (N_5086,N_4819,N_4973);
or U5087 (N_5087,N_4832,N_4820);
xor U5088 (N_5088,N_4827,N_4918);
xnor U5089 (N_5089,N_4781,N_4965);
nand U5090 (N_5090,N_4904,N_4974);
and U5091 (N_5091,N_4936,N_4865);
xnor U5092 (N_5092,N_4876,N_4814);
and U5093 (N_5093,N_4983,N_4881);
nand U5094 (N_5094,N_4802,N_4861);
and U5095 (N_5095,N_4995,N_4922);
or U5096 (N_5096,N_4835,N_4906);
and U5097 (N_5097,N_4910,N_4883);
or U5098 (N_5098,N_4836,N_4966);
xnor U5099 (N_5099,N_4867,N_4946);
or U5100 (N_5100,N_4866,N_4762);
or U5101 (N_5101,N_4875,N_4799);
nand U5102 (N_5102,N_4798,N_4885);
xor U5103 (N_5103,N_4789,N_4773);
nand U5104 (N_5104,N_4964,N_4996);
and U5105 (N_5105,N_4980,N_4967);
nand U5106 (N_5106,N_4793,N_4932);
xnor U5107 (N_5107,N_4891,N_4916);
xor U5108 (N_5108,N_4917,N_4923);
nor U5109 (N_5109,N_4986,N_4920);
nand U5110 (N_5110,N_4800,N_4939);
or U5111 (N_5111,N_4901,N_4792);
nand U5112 (N_5112,N_4758,N_4947);
and U5113 (N_5113,N_4774,N_4992);
nand U5114 (N_5114,N_4958,N_4915);
or U5115 (N_5115,N_4846,N_4830);
xor U5116 (N_5116,N_4961,N_4948);
xnor U5117 (N_5117,N_4882,N_4894);
nor U5118 (N_5118,N_4927,N_4985);
xnor U5119 (N_5119,N_4764,N_4824);
nor U5120 (N_5120,N_4928,N_4889);
xor U5121 (N_5121,N_4972,N_4843);
or U5122 (N_5122,N_4871,N_4919);
xor U5123 (N_5123,N_4810,N_4878);
or U5124 (N_5124,N_4763,N_4988);
nand U5125 (N_5125,N_4795,N_4910);
or U5126 (N_5126,N_4897,N_4788);
nand U5127 (N_5127,N_4960,N_4838);
nor U5128 (N_5128,N_4823,N_4958);
xnor U5129 (N_5129,N_4953,N_4907);
nand U5130 (N_5130,N_4786,N_4848);
or U5131 (N_5131,N_4791,N_4952);
and U5132 (N_5132,N_4873,N_4892);
and U5133 (N_5133,N_4990,N_4976);
xnor U5134 (N_5134,N_4788,N_4956);
nor U5135 (N_5135,N_4861,N_4890);
and U5136 (N_5136,N_4907,N_4922);
or U5137 (N_5137,N_4988,N_4888);
and U5138 (N_5138,N_4830,N_4825);
and U5139 (N_5139,N_4947,N_4974);
or U5140 (N_5140,N_4950,N_4892);
nor U5141 (N_5141,N_4852,N_4861);
xor U5142 (N_5142,N_4901,N_4997);
nand U5143 (N_5143,N_4783,N_4928);
or U5144 (N_5144,N_4916,N_4755);
xor U5145 (N_5145,N_4836,N_4835);
nor U5146 (N_5146,N_4996,N_4768);
nand U5147 (N_5147,N_4935,N_4997);
nand U5148 (N_5148,N_4837,N_4897);
nor U5149 (N_5149,N_4852,N_4871);
or U5150 (N_5150,N_4874,N_4772);
or U5151 (N_5151,N_4802,N_4948);
or U5152 (N_5152,N_4796,N_4835);
or U5153 (N_5153,N_4972,N_4757);
xnor U5154 (N_5154,N_4771,N_4966);
and U5155 (N_5155,N_4784,N_4856);
and U5156 (N_5156,N_4883,N_4862);
nand U5157 (N_5157,N_4894,N_4874);
nand U5158 (N_5158,N_4834,N_4754);
and U5159 (N_5159,N_4971,N_4807);
and U5160 (N_5160,N_4799,N_4956);
nand U5161 (N_5161,N_4984,N_4842);
xnor U5162 (N_5162,N_4825,N_4946);
and U5163 (N_5163,N_4896,N_4814);
xnor U5164 (N_5164,N_4884,N_4906);
xor U5165 (N_5165,N_4876,N_4779);
xor U5166 (N_5166,N_4775,N_4953);
nand U5167 (N_5167,N_4887,N_4886);
or U5168 (N_5168,N_4906,N_4977);
xnor U5169 (N_5169,N_4751,N_4917);
and U5170 (N_5170,N_4758,N_4962);
or U5171 (N_5171,N_4977,N_4841);
and U5172 (N_5172,N_4989,N_4905);
or U5173 (N_5173,N_4770,N_4981);
nand U5174 (N_5174,N_4915,N_4818);
or U5175 (N_5175,N_4946,N_4982);
nand U5176 (N_5176,N_4932,N_4841);
nand U5177 (N_5177,N_4944,N_4959);
and U5178 (N_5178,N_4817,N_4963);
xnor U5179 (N_5179,N_4953,N_4779);
xnor U5180 (N_5180,N_4764,N_4809);
and U5181 (N_5181,N_4788,N_4958);
xor U5182 (N_5182,N_4759,N_4885);
nand U5183 (N_5183,N_4952,N_4787);
or U5184 (N_5184,N_4968,N_4859);
nand U5185 (N_5185,N_4959,N_4808);
xor U5186 (N_5186,N_4941,N_4958);
nand U5187 (N_5187,N_4875,N_4848);
nor U5188 (N_5188,N_4900,N_4941);
nor U5189 (N_5189,N_4863,N_4912);
nor U5190 (N_5190,N_4915,N_4900);
nand U5191 (N_5191,N_4774,N_4966);
nand U5192 (N_5192,N_4897,N_4951);
xor U5193 (N_5193,N_4791,N_4783);
or U5194 (N_5194,N_4842,N_4930);
xnor U5195 (N_5195,N_4918,N_4992);
or U5196 (N_5196,N_4921,N_4896);
and U5197 (N_5197,N_4837,N_4822);
nand U5198 (N_5198,N_4995,N_4939);
or U5199 (N_5199,N_4816,N_4783);
or U5200 (N_5200,N_4920,N_4998);
xnor U5201 (N_5201,N_4893,N_4850);
xor U5202 (N_5202,N_4985,N_4801);
nand U5203 (N_5203,N_4789,N_4851);
nor U5204 (N_5204,N_4764,N_4859);
or U5205 (N_5205,N_4926,N_4762);
and U5206 (N_5206,N_4892,N_4939);
nand U5207 (N_5207,N_4872,N_4784);
nand U5208 (N_5208,N_4963,N_4844);
nand U5209 (N_5209,N_4987,N_4919);
nand U5210 (N_5210,N_4807,N_4759);
xor U5211 (N_5211,N_4895,N_4803);
or U5212 (N_5212,N_4825,N_4930);
or U5213 (N_5213,N_4907,N_4766);
xnor U5214 (N_5214,N_4957,N_4894);
nor U5215 (N_5215,N_4929,N_4786);
xnor U5216 (N_5216,N_4878,N_4929);
nor U5217 (N_5217,N_4755,N_4914);
and U5218 (N_5218,N_4796,N_4764);
nand U5219 (N_5219,N_4789,N_4783);
nand U5220 (N_5220,N_4951,N_4845);
and U5221 (N_5221,N_4837,N_4877);
xnor U5222 (N_5222,N_4932,N_4796);
nand U5223 (N_5223,N_4871,N_4794);
or U5224 (N_5224,N_4847,N_4820);
nor U5225 (N_5225,N_4853,N_4998);
or U5226 (N_5226,N_4782,N_4926);
nand U5227 (N_5227,N_4995,N_4759);
nand U5228 (N_5228,N_4794,N_4898);
and U5229 (N_5229,N_4796,N_4818);
xor U5230 (N_5230,N_4874,N_4950);
xor U5231 (N_5231,N_4984,N_4935);
xor U5232 (N_5232,N_4871,N_4780);
xor U5233 (N_5233,N_4966,N_4862);
or U5234 (N_5234,N_4784,N_4800);
nand U5235 (N_5235,N_4957,N_4992);
nand U5236 (N_5236,N_4806,N_4753);
nor U5237 (N_5237,N_4798,N_4750);
nor U5238 (N_5238,N_4874,N_4944);
and U5239 (N_5239,N_4896,N_4987);
xnor U5240 (N_5240,N_4963,N_4950);
nor U5241 (N_5241,N_4928,N_4861);
and U5242 (N_5242,N_4904,N_4875);
or U5243 (N_5243,N_4954,N_4968);
or U5244 (N_5244,N_4950,N_4930);
or U5245 (N_5245,N_4993,N_4942);
and U5246 (N_5246,N_4968,N_4850);
or U5247 (N_5247,N_4843,N_4905);
xor U5248 (N_5248,N_4915,N_4879);
or U5249 (N_5249,N_4960,N_4966);
nor U5250 (N_5250,N_5037,N_5110);
xnor U5251 (N_5251,N_5192,N_5011);
or U5252 (N_5252,N_5242,N_5022);
xnor U5253 (N_5253,N_5156,N_5069);
xor U5254 (N_5254,N_5160,N_5164);
xor U5255 (N_5255,N_5155,N_5120);
or U5256 (N_5256,N_5051,N_5142);
or U5257 (N_5257,N_5139,N_5029);
nand U5258 (N_5258,N_5071,N_5053);
nand U5259 (N_5259,N_5040,N_5092);
xnor U5260 (N_5260,N_5196,N_5100);
xor U5261 (N_5261,N_5209,N_5178);
nand U5262 (N_5262,N_5055,N_5072);
and U5263 (N_5263,N_5171,N_5119);
xnor U5264 (N_5264,N_5202,N_5104);
nand U5265 (N_5265,N_5033,N_5025);
or U5266 (N_5266,N_5206,N_5005);
and U5267 (N_5267,N_5225,N_5246);
nand U5268 (N_5268,N_5030,N_5048);
nand U5269 (N_5269,N_5159,N_5168);
or U5270 (N_5270,N_5123,N_5230);
nand U5271 (N_5271,N_5162,N_5075);
and U5272 (N_5272,N_5204,N_5219);
xor U5273 (N_5273,N_5006,N_5080);
nor U5274 (N_5274,N_5107,N_5115);
xor U5275 (N_5275,N_5101,N_5086);
or U5276 (N_5276,N_5041,N_5042);
and U5277 (N_5277,N_5098,N_5131);
nor U5278 (N_5278,N_5111,N_5036);
xor U5279 (N_5279,N_5044,N_5108);
and U5280 (N_5280,N_5191,N_5085);
nand U5281 (N_5281,N_5243,N_5097);
nor U5282 (N_5282,N_5231,N_5017);
nand U5283 (N_5283,N_5163,N_5114);
or U5284 (N_5284,N_5102,N_5129);
nand U5285 (N_5285,N_5158,N_5176);
nand U5286 (N_5286,N_5004,N_5140);
or U5287 (N_5287,N_5014,N_5154);
nor U5288 (N_5288,N_5000,N_5028);
and U5289 (N_5289,N_5238,N_5064);
nor U5290 (N_5290,N_5147,N_5223);
and U5291 (N_5291,N_5150,N_5197);
nand U5292 (N_5292,N_5229,N_5118);
nor U5293 (N_5293,N_5239,N_5074);
xor U5294 (N_5294,N_5247,N_5057);
and U5295 (N_5295,N_5018,N_5058);
nor U5296 (N_5296,N_5094,N_5207);
and U5297 (N_5297,N_5039,N_5237);
xor U5298 (N_5298,N_5235,N_5077);
or U5299 (N_5299,N_5249,N_5054);
xor U5300 (N_5300,N_5153,N_5190);
and U5301 (N_5301,N_5134,N_5173);
nor U5302 (N_5302,N_5045,N_5091);
or U5303 (N_5303,N_5095,N_5245);
and U5304 (N_5304,N_5188,N_5001);
xor U5305 (N_5305,N_5081,N_5185);
xnor U5306 (N_5306,N_5138,N_5015);
and U5307 (N_5307,N_5215,N_5109);
nand U5308 (N_5308,N_5236,N_5047);
nor U5309 (N_5309,N_5093,N_5078);
or U5310 (N_5310,N_5193,N_5221);
or U5311 (N_5311,N_5046,N_5021);
nor U5312 (N_5312,N_5026,N_5052);
nor U5313 (N_5313,N_5208,N_5116);
nand U5314 (N_5314,N_5061,N_5205);
xor U5315 (N_5315,N_5177,N_5027);
or U5316 (N_5316,N_5184,N_5083);
xor U5317 (N_5317,N_5082,N_5186);
nor U5318 (N_5318,N_5244,N_5012);
and U5319 (N_5319,N_5210,N_5010);
and U5320 (N_5320,N_5013,N_5200);
or U5321 (N_5321,N_5175,N_5189);
xnor U5322 (N_5322,N_5035,N_5161);
and U5323 (N_5323,N_5224,N_5216);
xnor U5324 (N_5324,N_5169,N_5183);
xnor U5325 (N_5325,N_5063,N_5062);
or U5326 (N_5326,N_5034,N_5144);
or U5327 (N_5327,N_5234,N_5128);
nor U5328 (N_5328,N_5222,N_5066);
and U5329 (N_5329,N_5220,N_5137);
nor U5330 (N_5330,N_5143,N_5038);
and U5331 (N_5331,N_5132,N_5122);
xor U5332 (N_5332,N_5031,N_5126);
nand U5333 (N_5333,N_5228,N_5009);
xnor U5334 (N_5334,N_5020,N_5167);
nor U5335 (N_5335,N_5157,N_5073);
nor U5336 (N_5336,N_5124,N_5136);
xor U5337 (N_5337,N_5099,N_5056);
xor U5338 (N_5338,N_5130,N_5002);
xor U5339 (N_5339,N_5213,N_5172);
nor U5340 (N_5340,N_5194,N_5016);
nand U5341 (N_5341,N_5089,N_5096);
xnor U5342 (N_5342,N_5112,N_5240);
and U5343 (N_5343,N_5067,N_5133);
and U5344 (N_5344,N_5105,N_5084);
and U5345 (N_5345,N_5090,N_5008);
xor U5346 (N_5346,N_5151,N_5059);
and U5347 (N_5347,N_5195,N_5182);
xor U5348 (N_5348,N_5032,N_5141);
or U5349 (N_5349,N_5043,N_5174);
xor U5350 (N_5350,N_5233,N_5023);
nand U5351 (N_5351,N_5007,N_5113);
xor U5352 (N_5352,N_5070,N_5060);
nor U5353 (N_5353,N_5227,N_5146);
nand U5354 (N_5354,N_5165,N_5003);
nand U5355 (N_5355,N_5019,N_5217);
nor U5356 (N_5356,N_5024,N_5127);
nand U5357 (N_5357,N_5170,N_5149);
and U5358 (N_5358,N_5214,N_5248);
xnor U5359 (N_5359,N_5199,N_5121);
or U5360 (N_5360,N_5232,N_5145);
nand U5361 (N_5361,N_5125,N_5241);
nand U5362 (N_5362,N_5103,N_5065);
nor U5363 (N_5363,N_5050,N_5201);
nor U5364 (N_5364,N_5198,N_5212);
xor U5365 (N_5365,N_5135,N_5049);
nor U5366 (N_5366,N_5211,N_5218);
or U5367 (N_5367,N_5079,N_5068);
and U5368 (N_5368,N_5088,N_5166);
and U5369 (N_5369,N_5179,N_5187);
nand U5370 (N_5370,N_5106,N_5181);
or U5371 (N_5371,N_5117,N_5226);
and U5372 (N_5372,N_5180,N_5148);
nand U5373 (N_5373,N_5152,N_5203);
nor U5374 (N_5374,N_5076,N_5087);
nand U5375 (N_5375,N_5228,N_5249);
or U5376 (N_5376,N_5052,N_5249);
and U5377 (N_5377,N_5225,N_5051);
or U5378 (N_5378,N_5237,N_5066);
and U5379 (N_5379,N_5040,N_5178);
nor U5380 (N_5380,N_5169,N_5146);
and U5381 (N_5381,N_5080,N_5171);
xnor U5382 (N_5382,N_5013,N_5148);
or U5383 (N_5383,N_5051,N_5152);
nor U5384 (N_5384,N_5179,N_5154);
xor U5385 (N_5385,N_5015,N_5211);
nor U5386 (N_5386,N_5009,N_5214);
xnor U5387 (N_5387,N_5140,N_5003);
and U5388 (N_5388,N_5048,N_5160);
nand U5389 (N_5389,N_5205,N_5157);
and U5390 (N_5390,N_5154,N_5120);
nand U5391 (N_5391,N_5138,N_5006);
nor U5392 (N_5392,N_5084,N_5043);
or U5393 (N_5393,N_5168,N_5123);
xor U5394 (N_5394,N_5065,N_5196);
nor U5395 (N_5395,N_5078,N_5070);
xor U5396 (N_5396,N_5105,N_5149);
and U5397 (N_5397,N_5079,N_5069);
and U5398 (N_5398,N_5062,N_5049);
nand U5399 (N_5399,N_5105,N_5235);
and U5400 (N_5400,N_5232,N_5221);
or U5401 (N_5401,N_5118,N_5156);
or U5402 (N_5402,N_5160,N_5039);
xnor U5403 (N_5403,N_5026,N_5220);
xnor U5404 (N_5404,N_5193,N_5054);
and U5405 (N_5405,N_5187,N_5246);
nand U5406 (N_5406,N_5040,N_5006);
xnor U5407 (N_5407,N_5035,N_5124);
or U5408 (N_5408,N_5010,N_5169);
nand U5409 (N_5409,N_5137,N_5130);
nand U5410 (N_5410,N_5182,N_5176);
nand U5411 (N_5411,N_5214,N_5099);
nand U5412 (N_5412,N_5165,N_5231);
or U5413 (N_5413,N_5053,N_5029);
or U5414 (N_5414,N_5012,N_5126);
nand U5415 (N_5415,N_5221,N_5086);
xnor U5416 (N_5416,N_5008,N_5120);
nand U5417 (N_5417,N_5013,N_5012);
xnor U5418 (N_5418,N_5040,N_5236);
xnor U5419 (N_5419,N_5008,N_5177);
and U5420 (N_5420,N_5079,N_5005);
or U5421 (N_5421,N_5045,N_5135);
or U5422 (N_5422,N_5016,N_5047);
or U5423 (N_5423,N_5041,N_5153);
xor U5424 (N_5424,N_5061,N_5032);
nand U5425 (N_5425,N_5097,N_5011);
nand U5426 (N_5426,N_5217,N_5132);
nor U5427 (N_5427,N_5074,N_5058);
and U5428 (N_5428,N_5086,N_5013);
xor U5429 (N_5429,N_5023,N_5035);
nor U5430 (N_5430,N_5135,N_5070);
and U5431 (N_5431,N_5187,N_5080);
xor U5432 (N_5432,N_5001,N_5090);
nor U5433 (N_5433,N_5016,N_5104);
nand U5434 (N_5434,N_5194,N_5115);
nor U5435 (N_5435,N_5224,N_5077);
nor U5436 (N_5436,N_5098,N_5217);
nor U5437 (N_5437,N_5211,N_5148);
and U5438 (N_5438,N_5021,N_5230);
or U5439 (N_5439,N_5218,N_5050);
and U5440 (N_5440,N_5176,N_5207);
or U5441 (N_5441,N_5198,N_5227);
and U5442 (N_5442,N_5005,N_5128);
nor U5443 (N_5443,N_5046,N_5133);
or U5444 (N_5444,N_5162,N_5115);
nor U5445 (N_5445,N_5006,N_5023);
and U5446 (N_5446,N_5146,N_5219);
and U5447 (N_5447,N_5216,N_5062);
and U5448 (N_5448,N_5063,N_5210);
xor U5449 (N_5449,N_5000,N_5065);
nor U5450 (N_5450,N_5018,N_5200);
nor U5451 (N_5451,N_5184,N_5120);
nor U5452 (N_5452,N_5171,N_5043);
and U5453 (N_5453,N_5037,N_5090);
nor U5454 (N_5454,N_5109,N_5130);
and U5455 (N_5455,N_5040,N_5191);
nand U5456 (N_5456,N_5221,N_5091);
nor U5457 (N_5457,N_5180,N_5156);
and U5458 (N_5458,N_5107,N_5083);
or U5459 (N_5459,N_5066,N_5159);
and U5460 (N_5460,N_5220,N_5224);
nor U5461 (N_5461,N_5217,N_5212);
xnor U5462 (N_5462,N_5230,N_5142);
or U5463 (N_5463,N_5105,N_5167);
or U5464 (N_5464,N_5119,N_5089);
nor U5465 (N_5465,N_5161,N_5138);
or U5466 (N_5466,N_5083,N_5023);
nand U5467 (N_5467,N_5122,N_5164);
nand U5468 (N_5468,N_5047,N_5192);
or U5469 (N_5469,N_5083,N_5177);
nor U5470 (N_5470,N_5248,N_5127);
or U5471 (N_5471,N_5162,N_5024);
and U5472 (N_5472,N_5166,N_5092);
or U5473 (N_5473,N_5106,N_5022);
or U5474 (N_5474,N_5099,N_5037);
nand U5475 (N_5475,N_5106,N_5075);
and U5476 (N_5476,N_5153,N_5012);
xnor U5477 (N_5477,N_5016,N_5219);
nor U5478 (N_5478,N_5151,N_5027);
xnor U5479 (N_5479,N_5104,N_5086);
or U5480 (N_5480,N_5032,N_5234);
and U5481 (N_5481,N_5141,N_5224);
nor U5482 (N_5482,N_5042,N_5185);
or U5483 (N_5483,N_5019,N_5040);
or U5484 (N_5484,N_5140,N_5158);
and U5485 (N_5485,N_5076,N_5042);
and U5486 (N_5486,N_5233,N_5220);
nand U5487 (N_5487,N_5075,N_5058);
and U5488 (N_5488,N_5093,N_5088);
and U5489 (N_5489,N_5209,N_5216);
and U5490 (N_5490,N_5097,N_5197);
and U5491 (N_5491,N_5150,N_5151);
nand U5492 (N_5492,N_5017,N_5071);
nor U5493 (N_5493,N_5237,N_5242);
nor U5494 (N_5494,N_5014,N_5199);
xor U5495 (N_5495,N_5011,N_5176);
and U5496 (N_5496,N_5212,N_5044);
and U5497 (N_5497,N_5032,N_5089);
xnor U5498 (N_5498,N_5200,N_5066);
nor U5499 (N_5499,N_5045,N_5049);
or U5500 (N_5500,N_5423,N_5468);
xor U5501 (N_5501,N_5394,N_5340);
nor U5502 (N_5502,N_5427,N_5321);
or U5503 (N_5503,N_5457,N_5403);
and U5504 (N_5504,N_5475,N_5426);
nor U5505 (N_5505,N_5498,N_5291);
nand U5506 (N_5506,N_5370,N_5329);
xor U5507 (N_5507,N_5355,N_5465);
nand U5508 (N_5508,N_5385,N_5470);
nand U5509 (N_5509,N_5398,N_5318);
xor U5510 (N_5510,N_5311,N_5358);
nand U5511 (N_5511,N_5369,N_5407);
xor U5512 (N_5512,N_5364,N_5401);
xor U5513 (N_5513,N_5327,N_5346);
nand U5514 (N_5514,N_5303,N_5301);
nand U5515 (N_5515,N_5411,N_5477);
nand U5516 (N_5516,N_5491,N_5404);
nor U5517 (N_5517,N_5371,N_5268);
xnor U5518 (N_5518,N_5424,N_5255);
xnor U5519 (N_5519,N_5387,N_5383);
and U5520 (N_5520,N_5489,N_5494);
nor U5521 (N_5521,N_5484,N_5474);
nor U5522 (N_5522,N_5325,N_5386);
and U5523 (N_5523,N_5390,N_5342);
nor U5524 (N_5524,N_5436,N_5320);
and U5525 (N_5525,N_5377,N_5450);
or U5526 (N_5526,N_5391,N_5286);
nand U5527 (N_5527,N_5351,N_5372);
and U5528 (N_5528,N_5280,N_5428);
nand U5529 (N_5529,N_5365,N_5413);
xnor U5530 (N_5530,N_5375,N_5353);
or U5531 (N_5531,N_5282,N_5270);
nor U5532 (N_5532,N_5460,N_5308);
xor U5533 (N_5533,N_5279,N_5297);
and U5534 (N_5534,N_5402,N_5352);
nor U5535 (N_5535,N_5345,N_5343);
and U5536 (N_5536,N_5462,N_5488);
nor U5537 (N_5537,N_5322,N_5256);
xnor U5538 (N_5538,N_5487,N_5338);
or U5539 (N_5539,N_5493,N_5356);
nor U5540 (N_5540,N_5298,N_5389);
and U5541 (N_5541,N_5400,N_5478);
or U5542 (N_5542,N_5393,N_5271);
xnor U5543 (N_5543,N_5482,N_5348);
nor U5544 (N_5544,N_5419,N_5388);
and U5545 (N_5545,N_5454,N_5467);
xnor U5546 (N_5546,N_5319,N_5337);
nand U5547 (N_5547,N_5328,N_5366);
or U5548 (N_5548,N_5359,N_5485);
xor U5549 (N_5549,N_5284,N_5473);
xnor U5550 (N_5550,N_5379,N_5444);
or U5551 (N_5551,N_5492,N_5350);
nor U5552 (N_5552,N_5336,N_5331);
and U5553 (N_5553,N_5262,N_5252);
nor U5554 (N_5554,N_5480,N_5455);
xor U5555 (N_5555,N_5447,N_5274);
and U5556 (N_5556,N_5332,N_5437);
nand U5557 (N_5557,N_5368,N_5433);
and U5558 (N_5558,N_5281,N_5299);
nand U5559 (N_5559,N_5438,N_5333);
xnor U5560 (N_5560,N_5263,N_5324);
nand U5561 (N_5561,N_5452,N_5395);
or U5562 (N_5562,N_5373,N_5309);
or U5563 (N_5563,N_5314,N_5417);
nand U5564 (N_5564,N_5323,N_5440);
or U5565 (N_5565,N_5292,N_5431);
and U5566 (N_5566,N_5296,N_5254);
nand U5567 (N_5567,N_5310,N_5344);
or U5568 (N_5568,N_5415,N_5459);
xnor U5569 (N_5569,N_5432,N_5250);
xor U5570 (N_5570,N_5277,N_5283);
or U5571 (N_5571,N_5442,N_5464);
xnor U5572 (N_5572,N_5312,N_5429);
nand U5573 (N_5573,N_5305,N_5430);
nand U5574 (N_5574,N_5490,N_5294);
or U5575 (N_5575,N_5374,N_5414);
and U5576 (N_5576,N_5275,N_5330);
xor U5577 (N_5577,N_5316,N_5264);
nand U5578 (N_5578,N_5290,N_5251);
and U5579 (N_5579,N_5421,N_5361);
xnor U5580 (N_5580,N_5363,N_5453);
nand U5581 (N_5581,N_5258,N_5495);
nor U5582 (N_5582,N_5266,N_5260);
nand U5583 (N_5583,N_5339,N_5289);
and U5584 (N_5584,N_5441,N_5412);
or U5585 (N_5585,N_5253,N_5326);
nand U5586 (N_5586,N_5425,N_5313);
nand U5587 (N_5587,N_5472,N_5418);
or U5588 (N_5588,N_5461,N_5306);
nand U5589 (N_5589,N_5341,N_5392);
and U5590 (N_5590,N_5479,N_5448);
nand U5591 (N_5591,N_5302,N_5378);
nor U5592 (N_5592,N_5466,N_5410);
nor U5593 (N_5593,N_5420,N_5334);
and U5594 (N_5594,N_5259,N_5376);
or U5595 (N_5595,N_5382,N_5445);
and U5596 (N_5596,N_5416,N_5304);
nor U5597 (N_5597,N_5278,N_5384);
or U5598 (N_5598,N_5357,N_5471);
or U5599 (N_5599,N_5347,N_5497);
xor U5600 (N_5600,N_5273,N_5496);
or U5601 (N_5601,N_5399,N_5397);
or U5602 (N_5602,N_5481,N_5408);
nor U5603 (N_5603,N_5354,N_5272);
xor U5604 (N_5604,N_5261,N_5499);
or U5605 (N_5605,N_5265,N_5406);
or U5606 (N_5606,N_5367,N_5469);
nand U5607 (N_5607,N_5335,N_5267);
xnor U5608 (N_5608,N_5458,N_5439);
and U5609 (N_5609,N_5446,N_5288);
or U5610 (N_5610,N_5435,N_5409);
xor U5611 (N_5611,N_5434,N_5295);
and U5612 (N_5612,N_5349,N_5443);
or U5613 (N_5613,N_5483,N_5287);
nor U5614 (N_5614,N_5315,N_5476);
nor U5615 (N_5615,N_5360,N_5456);
or U5616 (N_5616,N_5463,N_5276);
nand U5617 (N_5617,N_5449,N_5451);
nand U5618 (N_5618,N_5307,N_5285);
and U5619 (N_5619,N_5381,N_5422);
nor U5620 (N_5620,N_5300,N_5362);
nor U5621 (N_5621,N_5293,N_5396);
nand U5622 (N_5622,N_5317,N_5380);
or U5623 (N_5623,N_5405,N_5486);
nor U5624 (N_5624,N_5257,N_5269);
or U5625 (N_5625,N_5476,N_5417);
nand U5626 (N_5626,N_5472,N_5490);
or U5627 (N_5627,N_5449,N_5406);
and U5628 (N_5628,N_5380,N_5481);
nor U5629 (N_5629,N_5327,N_5468);
nand U5630 (N_5630,N_5281,N_5394);
and U5631 (N_5631,N_5368,N_5337);
nor U5632 (N_5632,N_5261,N_5401);
xnor U5633 (N_5633,N_5493,N_5460);
and U5634 (N_5634,N_5312,N_5385);
or U5635 (N_5635,N_5276,N_5428);
nand U5636 (N_5636,N_5440,N_5328);
nor U5637 (N_5637,N_5402,N_5457);
xor U5638 (N_5638,N_5266,N_5406);
nand U5639 (N_5639,N_5280,N_5339);
or U5640 (N_5640,N_5258,N_5408);
or U5641 (N_5641,N_5306,N_5273);
and U5642 (N_5642,N_5315,N_5342);
nor U5643 (N_5643,N_5299,N_5301);
nor U5644 (N_5644,N_5395,N_5411);
and U5645 (N_5645,N_5463,N_5316);
nor U5646 (N_5646,N_5404,N_5497);
and U5647 (N_5647,N_5462,N_5313);
or U5648 (N_5648,N_5392,N_5417);
or U5649 (N_5649,N_5257,N_5491);
or U5650 (N_5650,N_5464,N_5272);
nor U5651 (N_5651,N_5460,N_5257);
nand U5652 (N_5652,N_5446,N_5463);
and U5653 (N_5653,N_5342,N_5344);
or U5654 (N_5654,N_5439,N_5327);
xnor U5655 (N_5655,N_5256,N_5470);
or U5656 (N_5656,N_5466,N_5407);
nor U5657 (N_5657,N_5363,N_5273);
nor U5658 (N_5658,N_5301,N_5291);
or U5659 (N_5659,N_5329,N_5297);
xor U5660 (N_5660,N_5329,N_5429);
nor U5661 (N_5661,N_5455,N_5484);
and U5662 (N_5662,N_5297,N_5260);
nor U5663 (N_5663,N_5302,N_5415);
and U5664 (N_5664,N_5492,N_5400);
nand U5665 (N_5665,N_5422,N_5441);
and U5666 (N_5666,N_5351,N_5380);
or U5667 (N_5667,N_5257,N_5260);
or U5668 (N_5668,N_5352,N_5400);
and U5669 (N_5669,N_5326,N_5399);
nand U5670 (N_5670,N_5293,N_5279);
and U5671 (N_5671,N_5451,N_5448);
and U5672 (N_5672,N_5475,N_5290);
or U5673 (N_5673,N_5378,N_5257);
and U5674 (N_5674,N_5323,N_5359);
and U5675 (N_5675,N_5487,N_5256);
nand U5676 (N_5676,N_5491,N_5493);
xor U5677 (N_5677,N_5484,N_5476);
xnor U5678 (N_5678,N_5344,N_5480);
xor U5679 (N_5679,N_5332,N_5341);
or U5680 (N_5680,N_5398,N_5362);
nor U5681 (N_5681,N_5381,N_5469);
or U5682 (N_5682,N_5488,N_5382);
nor U5683 (N_5683,N_5353,N_5448);
or U5684 (N_5684,N_5335,N_5457);
nand U5685 (N_5685,N_5352,N_5398);
or U5686 (N_5686,N_5449,N_5265);
nand U5687 (N_5687,N_5430,N_5497);
nor U5688 (N_5688,N_5342,N_5372);
nand U5689 (N_5689,N_5422,N_5417);
nand U5690 (N_5690,N_5355,N_5328);
xor U5691 (N_5691,N_5298,N_5315);
xnor U5692 (N_5692,N_5480,N_5498);
or U5693 (N_5693,N_5376,N_5368);
nand U5694 (N_5694,N_5402,N_5265);
and U5695 (N_5695,N_5419,N_5409);
nor U5696 (N_5696,N_5438,N_5491);
xor U5697 (N_5697,N_5447,N_5364);
nand U5698 (N_5698,N_5408,N_5355);
nand U5699 (N_5699,N_5418,N_5272);
xor U5700 (N_5700,N_5403,N_5265);
or U5701 (N_5701,N_5383,N_5453);
or U5702 (N_5702,N_5374,N_5339);
or U5703 (N_5703,N_5407,N_5333);
or U5704 (N_5704,N_5430,N_5464);
or U5705 (N_5705,N_5294,N_5372);
and U5706 (N_5706,N_5336,N_5445);
and U5707 (N_5707,N_5351,N_5411);
nor U5708 (N_5708,N_5398,N_5407);
nor U5709 (N_5709,N_5446,N_5309);
and U5710 (N_5710,N_5496,N_5406);
nor U5711 (N_5711,N_5455,N_5373);
nand U5712 (N_5712,N_5309,N_5474);
and U5713 (N_5713,N_5467,N_5409);
and U5714 (N_5714,N_5313,N_5274);
nand U5715 (N_5715,N_5486,N_5335);
nand U5716 (N_5716,N_5298,N_5308);
or U5717 (N_5717,N_5319,N_5272);
nor U5718 (N_5718,N_5334,N_5306);
nor U5719 (N_5719,N_5318,N_5294);
nand U5720 (N_5720,N_5412,N_5485);
xnor U5721 (N_5721,N_5279,N_5371);
and U5722 (N_5722,N_5458,N_5360);
nand U5723 (N_5723,N_5469,N_5448);
xor U5724 (N_5724,N_5330,N_5298);
and U5725 (N_5725,N_5390,N_5397);
or U5726 (N_5726,N_5306,N_5305);
nor U5727 (N_5727,N_5304,N_5494);
or U5728 (N_5728,N_5470,N_5264);
nor U5729 (N_5729,N_5331,N_5347);
and U5730 (N_5730,N_5269,N_5449);
and U5731 (N_5731,N_5448,N_5302);
or U5732 (N_5732,N_5369,N_5261);
xnor U5733 (N_5733,N_5293,N_5399);
or U5734 (N_5734,N_5452,N_5471);
nor U5735 (N_5735,N_5468,N_5450);
nand U5736 (N_5736,N_5366,N_5385);
xnor U5737 (N_5737,N_5309,N_5457);
or U5738 (N_5738,N_5476,N_5420);
nor U5739 (N_5739,N_5258,N_5317);
nor U5740 (N_5740,N_5290,N_5331);
or U5741 (N_5741,N_5482,N_5377);
nand U5742 (N_5742,N_5480,N_5469);
nor U5743 (N_5743,N_5320,N_5432);
xnor U5744 (N_5744,N_5393,N_5443);
nand U5745 (N_5745,N_5345,N_5259);
and U5746 (N_5746,N_5389,N_5264);
nand U5747 (N_5747,N_5317,N_5363);
and U5748 (N_5748,N_5369,N_5450);
or U5749 (N_5749,N_5376,N_5281);
xnor U5750 (N_5750,N_5632,N_5667);
and U5751 (N_5751,N_5704,N_5672);
nor U5752 (N_5752,N_5602,N_5531);
nor U5753 (N_5753,N_5567,N_5721);
xnor U5754 (N_5754,N_5702,N_5501);
xnor U5755 (N_5755,N_5689,N_5521);
or U5756 (N_5756,N_5722,N_5591);
nand U5757 (N_5757,N_5708,N_5514);
xnor U5758 (N_5758,N_5579,N_5601);
xor U5759 (N_5759,N_5636,N_5696);
nand U5760 (N_5760,N_5699,N_5691);
or U5761 (N_5761,N_5678,N_5538);
and U5762 (N_5762,N_5626,N_5551);
nand U5763 (N_5763,N_5652,N_5515);
nor U5764 (N_5764,N_5554,N_5629);
nor U5765 (N_5765,N_5736,N_5717);
nand U5766 (N_5766,N_5562,N_5525);
nand U5767 (N_5767,N_5507,N_5649);
and U5768 (N_5768,N_5547,N_5565);
and U5769 (N_5769,N_5533,N_5572);
xnor U5770 (N_5770,N_5552,N_5576);
nor U5771 (N_5771,N_5680,N_5613);
nor U5772 (N_5772,N_5697,N_5563);
nand U5773 (N_5773,N_5651,N_5719);
nor U5774 (N_5774,N_5596,N_5623);
nor U5775 (N_5775,N_5610,N_5738);
xor U5776 (N_5776,N_5612,N_5506);
and U5777 (N_5777,N_5509,N_5640);
nor U5778 (N_5778,N_5585,N_5664);
nor U5779 (N_5779,N_5677,N_5553);
xnor U5780 (N_5780,N_5542,N_5654);
xnor U5781 (N_5781,N_5526,N_5598);
and U5782 (N_5782,N_5695,N_5605);
nand U5783 (N_5783,N_5633,N_5622);
and U5784 (N_5784,N_5546,N_5663);
or U5785 (N_5785,N_5729,N_5684);
nor U5786 (N_5786,N_5643,N_5715);
xnor U5787 (N_5787,N_5517,N_5639);
and U5788 (N_5788,N_5524,N_5616);
or U5789 (N_5789,N_5726,N_5665);
xor U5790 (N_5790,N_5625,N_5518);
or U5791 (N_5791,N_5519,N_5559);
nor U5792 (N_5792,N_5549,N_5561);
xor U5793 (N_5793,N_5588,N_5737);
xnor U5794 (N_5794,N_5617,N_5637);
nor U5795 (N_5795,N_5535,N_5638);
xor U5796 (N_5796,N_5630,N_5734);
nor U5797 (N_5797,N_5582,N_5711);
nor U5798 (N_5798,N_5540,N_5668);
nand U5799 (N_5799,N_5730,N_5511);
xor U5800 (N_5800,N_5669,N_5682);
nand U5801 (N_5801,N_5568,N_5688);
nor U5802 (N_5802,N_5676,N_5523);
xor U5803 (N_5803,N_5544,N_5698);
or U5804 (N_5804,N_5714,N_5670);
nor U5805 (N_5805,N_5650,N_5543);
xor U5806 (N_5806,N_5709,N_5566);
nor U5807 (N_5807,N_5583,N_5619);
nand U5808 (N_5808,N_5683,N_5536);
nand U5809 (N_5809,N_5510,N_5621);
or U5810 (N_5810,N_5575,N_5646);
nand U5811 (N_5811,N_5614,N_5690);
and U5812 (N_5812,N_5679,N_5745);
nand U5813 (N_5813,N_5603,N_5586);
or U5814 (N_5814,N_5513,N_5671);
nand U5815 (N_5815,N_5674,N_5700);
xnor U5816 (N_5816,N_5716,N_5590);
or U5817 (N_5817,N_5604,N_5500);
nor U5818 (N_5818,N_5743,N_5686);
or U5819 (N_5819,N_5658,N_5520);
or U5820 (N_5820,N_5581,N_5611);
and U5821 (N_5821,N_5728,N_5600);
nor U5822 (N_5822,N_5587,N_5558);
xnor U5823 (N_5823,N_5701,N_5548);
nor U5824 (N_5824,N_5528,N_5733);
or U5825 (N_5825,N_5693,N_5731);
or U5826 (N_5826,N_5556,N_5584);
nor U5827 (N_5827,N_5748,N_5534);
xnor U5828 (N_5828,N_5620,N_5564);
xor U5829 (N_5829,N_5573,N_5712);
and U5830 (N_5830,N_5735,N_5615);
nor U5831 (N_5831,N_5607,N_5609);
or U5832 (N_5832,N_5560,N_5685);
nand U5833 (N_5833,N_5527,N_5694);
xnor U5834 (N_5834,N_5706,N_5634);
xnor U5835 (N_5835,N_5642,N_5530);
or U5836 (N_5836,N_5570,N_5522);
xnor U5837 (N_5837,N_5631,N_5645);
nor U5838 (N_5838,N_5641,N_5541);
nand U5839 (N_5839,N_5681,N_5687);
xor U5840 (N_5840,N_5569,N_5732);
and U5841 (N_5841,N_5739,N_5574);
nor U5842 (N_5842,N_5742,N_5624);
and U5843 (N_5843,N_5661,N_5746);
nand U5844 (N_5844,N_5618,N_5504);
nand U5845 (N_5845,N_5727,N_5508);
or U5846 (N_5846,N_5744,N_5662);
nand U5847 (N_5847,N_5571,N_5512);
or U5848 (N_5848,N_5647,N_5648);
xor U5849 (N_5849,N_5529,N_5592);
or U5850 (N_5850,N_5557,N_5657);
nand U5851 (N_5851,N_5595,N_5589);
and U5852 (N_5852,N_5505,N_5741);
and U5853 (N_5853,N_5580,N_5539);
xor U5854 (N_5854,N_5655,N_5725);
or U5855 (N_5855,N_5550,N_5555);
xor U5856 (N_5856,N_5628,N_5593);
nand U5857 (N_5857,N_5707,N_5718);
nand U5858 (N_5858,N_5740,N_5644);
or U5859 (N_5859,N_5627,N_5666);
nor U5860 (N_5860,N_5656,N_5608);
nor U5861 (N_5861,N_5577,N_5578);
nand U5862 (N_5862,N_5545,N_5503);
nand U5863 (N_5863,N_5532,N_5673);
xor U5864 (N_5864,N_5720,N_5705);
and U5865 (N_5865,N_5723,N_5749);
or U5866 (N_5866,N_5660,N_5710);
nor U5867 (N_5867,N_5606,N_5502);
xor U5868 (N_5868,N_5724,N_5703);
xor U5869 (N_5869,N_5675,N_5653);
and U5870 (N_5870,N_5537,N_5692);
xnor U5871 (N_5871,N_5635,N_5516);
or U5872 (N_5872,N_5747,N_5597);
or U5873 (N_5873,N_5599,N_5659);
and U5874 (N_5874,N_5594,N_5713);
nand U5875 (N_5875,N_5726,N_5518);
xor U5876 (N_5876,N_5550,N_5617);
xnor U5877 (N_5877,N_5662,N_5605);
nor U5878 (N_5878,N_5655,N_5583);
nand U5879 (N_5879,N_5529,N_5607);
xnor U5880 (N_5880,N_5655,N_5545);
nand U5881 (N_5881,N_5600,N_5510);
nor U5882 (N_5882,N_5589,N_5739);
xnor U5883 (N_5883,N_5729,N_5745);
and U5884 (N_5884,N_5617,N_5596);
or U5885 (N_5885,N_5729,N_5511);
nor U5886 (N_5886,N_5659,N_5651);
or U5887 (N_5887,N_5566,N_5625);
and U5888 (N_5888,N_5683,N_5743);
nand U5889 (N_5889,N_5724,N_5581);
and U5890 (N_5890,N_5674,N_5527);
xnor U5891 (N_5891,N_5500,N_5591);
nor U5892 (N_5892,N_5708,N_5655);
or U5893 (N_5893,N_5663,N_5565);
nand U5894 (N_5894,N_5613,N_5596);
nand U5895 (N_5895,N_5538,N_5733);
or U5896 (N_5896,N_5552,N_5587);
or U5897 (N_5897,N_5694,N_5550);
nor U5898 (N_5898,N_5720,N_5563);
nand U5899 (N_5899,N_5747,N_5542);
xnor U5900 (N_5900,N_5599,N_5704);
xnor U5901 (N_5901,N_5631,N_5571);
or U5902 (N_5902,N_5583,N_5667);
xor U5903 (N_5903,N_5733,N_5552);
nor U5904 (N_5904,N_5600,N_5727);
nor U5905 (N_5905,N_5543,N_5514);
nand U5906 (N_5906,N_5633,N_5616);
xor U5907 (N_5907,N_5743,N_5592);
nand U5908 (N_5908,N_5511,N_5652);
xor U5909 (N_5909,N_5524,N_5603);
and U5910 (N_5910,N_5558,N_5550);
or U5911 (N_5911,N_5577,N_5529);
xor U5912 (N_5912,N_5530,N_5645);
nor U5913 (N_5913,N_5662,N_5593);
nor U5914 (N_5914,N_5745,N_5696);
xor U5915 (N_5915,N_5726,N_5575);
nand U5916 (N_5916,N_5604,N_5606);
nor U5917 (N_5917,N_5715,N_5597);
and U5918 (N_5918,N_5700,N_5728);
nor U5919 (N_5919,N_5644,N_5512);
nor U5920 (N_5920,N_5636,N_5745);
or U5921 (N_5921,N_5705,N_5640);
xor U5922 (N_5922,N_5642,N_5721);
nor U5923 (N_5923,N_5704,N_5571);
nor U5924 (N_5924,N_5739,N_5555);
xnor U5925 (N_5925,N_5745,N_5734);
nor U5926 (N_5926,N_5569,N_5669);
and U5927 (N_5927,N_5721,N_5533);
nand U5928 (N_5928,N_5705,N_5665);
nor U5929 (N_5929,N_5625,N_5659);
or U5930 (N_5930,N_5645,N_5592);
nor U5931 (N_5931,N_5595,N_5563);
nor U5932 (N_5932,N_5584,N_5661);
nand U5933 (N_5933,N_5550,N_5628);
or U5934 (N_5934,N_5677,N_5510);
and U5935 (N_5935,N_5545,N_5729);
xnor U5936 (N_5936,N_5508,N_5583);
xor U5937 (N_5937,N_5699,N_5546);
nand U5938 (N_5938,N_5664,N_5672);
or U5939 (N_5939,N_5533,N_5629);
xnor U5940 (N_5940,N_5699,N_5666);
nor U5941 (N_5941,N_5719,N_5741);
xor U5942 (N_5942,N_5719,N_5511);
or U5943 (N_5943,N_5662,N_5749);
or U5944 (N_5944,N_5686,N_5716);
nor U5945 (N_5945,N_5749,N_5572);
and U5946 (N_5946,N_5518,N_5691);
nor U5947 (N_5947,N_5652,N_5616);
nand U5948 (N_5948,N_5554,N_5718);
nor U5949 (N_5949,N_5529,N_5739);
nor U5950 (N_5950,N_5573,N_5665);
nand U5951 (N_5951,N_5529,N_5736);
and U5952 (N_5952,N_5574,N_5563);
and U5953 (N_5953,N_5654,N_5521);
and U5954 (N_5954,N_5717,N_5529);
or U5955 (N_5955,N_5716,N_5742);
nand U5956 (N_5956,N_5631,N_5709);
xnor U5957 (N_5957,N_5650,N_5608);
or U5958 (N_5958,N_5673,N_5742);
and U5959 (N_5959,N_5618,N_5662);
or U5960 (N_5960,N_5542,N_5534);
nor U5961 (N_5961,N_5675,N_5683);
nor U5962 (N_5962,N_5622,N_5659);
nor U5963 (N_5963,N_5608,N_5679);
nand U5964 (N_5964,N_5560,N_5743);
or U5965 (N_5965,N_5628,N_5656);
or U5966 (N_5966,N_5605,N_5557);
nand U5967 (N_5967,N_5509,N_5531);
nand U5968 (N_5968,N_5602,N_5637);
nor U5969 (N_5969,N_5715,N_5559);
and U5970 (N_5970,N_5520,N_5593);
nor U5971 (N_5971,N_5745,N_5507);
nor U5972 (N_5972,N_5517,N_5604);
xor U5973 (N_5973,N_5532,N_5564);
nor U5974 (N_5974,N_5718,N_5524);
nor U5975 (N_5975,N_5678,N_5603);
nand U5976 (N_5976,N_5687,N_5625);
nor U5977 (N_5977,N_5582,N_5674);
nand U5978 (N_5978,N_5544,N_5712);
or U5979 (N_5979,N_5692,N_5566);
and U5980 (N_5980,N_5746,N_5503);
and U5981 (N_5981,N_5610,N_5737);
nor U5982 (N_5982,N_5574,N_5524);
xnor U5983 (N_5983,N_5596,N_5665);
xor U5984 (N_5984,N_5606,N_5504);
nor U5985 (N_5985,N_5736,N_5592);
nand U5986 (N_5986,N_5691,N_5622);
and U5987 (N_5987,N_5719,N_5646);
nor U5988 (N_5988,N_5579,N_5744);
or U5989 (N_5989,N_5636,N_5506);
or U5990 (N_5990,N_5565,N_5654);
nor U5991 (N_5991,N_5509,N_5501);
nand U5992 (N_5992,N_5529,N_5680);
or U5993 (N_5993,N_5729,N_5503);
xnor U5994 (N_5994,N_5723,N_5552);
nand U5995 (N_5995,N_5631,N_5574);
or U5996 (N_5996,N_5585,N_5674);
and U5997 (N_5997,N_5501,N_5684);
xnor U5998 (N_5998,N_5716,N_5704);
nand U5999 (N_5999,N_5573,N_5583);
and U6000 (N_6000,N_5999,N_5835);
or U6001 (N_6001,N_5790,N_5750);
nand U6002 (N_6002,N_5856,N_5858);
and U6003 (N_6003,N_5843,N_5759);
xnor U6004 (N_6004,N_5776,N_5883);
nor U6005 (N_6005,N_5939,N_5992);
nor U6006 (N_6006,N_5836,N_5851);
nand U6007 (N_6007,N_5787,N_5822);
or U6008 (N_6008,N_5782,N_5783);
or U6009 (N_6009,N_5954,N_5918);
xnor U6010 (N_6010,N_5844,N_5828);
xnor U6011 (N_6011,N_5961,N_5896);
nand U6012 (N_6012,N_5880,N_5838);
and U6013 (N_6013,N_5767,N_5842);
xor U6014 (N_6014,N_5934,N_5866);
xnor U6015 (N_6015,N_5957,N_5882);
xor U6016 (N_6016,N_5997,N_5801);
nand U6017 (N_6017,N_5834,N_5993);
nor U6018 (N_6018,N_5769,N_5873);
xor U6019 (N_6019,N_5974,N_5886);
xnor U6020 (N_6020,N_5906,N_5959);
nor U6021 (N_6021,N_5962,N_5865);
xor U6022 (N_6022,N_5871,N_5786);
xor U6023 (N_6023,N_5824,N_5755);
nand U6024 (N_6024,N_5812,N_5860);
or U6025 (N_6025,N_5995,N_5986);
nand U6026 (N_6026,N_5927,N_5916);
xor U6027 (N_6027,N_5756,N_5946);
xor U6028 (N_6028,N_5876,N_5968);
or U6029 (N_6029,N_5989,N_5940);
and U6030 (N_6030,N_5763,N_5966);
nor U6031 (N_6031,N_5823,N_5907);
or U6032 (N_6032,N_5789,N_5972);
xor U6033 (N_6033,N_5980,N_5874);
nand U6034 (N_6034,N_5803,N_5799);
nor U6035 (N_6035,N_5942,N_5788);
nand U6036 (N_6036,N_5936,N_5815);
and U6037 (N_6037,N_5955,N_5904);
or U6038 (N_6038,N_5963,N_5773);
nand U6039 (N_6039,N_5850,N_5821);
and U6040 (N_6040,N_5839,N_5784);
or U6041 (N_6041,N_5932,N_5967);
or U6042 (N_6042,N_5928,N_5827);
nor U6043 (N_6043,N_5899,N_5979);
and U6044 (N_6044,N_5833,N_5998);
xnor U6045 (N_6045,N_5900,N_5868);
and U6046 (N_6046,N_5973,N_5751);
nor U6047 (N_6047,N_5938,N_5914);
or U6048 (N_6048,N_5964,N_5853);
or U6049 (N_6049,N_5766,N_5798);
xor U6050 (N_6050,N_5826,N_5778);
xor U6051 (N_6051,N_5857,N_5920);
or U6052 (N_6052,N_5917,N_5921);
xor U6053 (N_6053,N_5820,N_5806);
xor U6054 (N_6054,N_5792,N_5831);
or U6055 (N_6055,N_5987,N_5791);
or U6056 (N_6056,N_5796,N_5847);
nor U6057 (N_6057,N_5802,N_5881);
or U6058 (N_6058,N_5922,N_5891);
xor U6059 (N_6059,N_5757,N_5867);
xor U6060 (N_6060,N_5794,N_5991);
and U6061 (N_6061,N_5912,N_5777);
xnor U6062 (N_6062,N_5800,N_5807);
nand U6063 (N_6063,N_5770,N_5852);
xor U6064 (N_6064,N_5864,N_5923);
nor U6065 (N_6065,N_5971,N_5895);
and U6066 (N_6066,N_5808,N_5772);
and U6067 (N_6067,N_5988,N_5976);
or U6068 (N_6068,N_5897,N_5981);
nor U6069 (N_6069,N_5945,N_5911);
nand U6070 (N_6070,N_5837,N_5996);
nand U6071 (N_6071,N_5930,N_5941);
nand U6072 (N_6072,N_5825,N_5848);
and U6073 (N_6073,N_5924,N_5944);
nor U6074 (N_6074,N_5951,N_5816);
nand U6075 (N_6075,N_5771,N_5785);
and U6076 (N_6076,N_5818,N_5926);
and U6077 (N_6077,N_5781,N_5810);
or U6078 (N_6078,N_5819,N_5870);
and U6079 (N_6079,N_5862,N_5931);
xnor U6080 (N_6080,N_5762,N_5947);
and U6081 (N_6081,N_5793,N_5948);
or U6082 (N_6082,N_5994,N_5805);
and U6083 (N_6083,N_5982,N_5985);
nand U6084 (N_6084,N_5840,N_5879);
nor U6085 (N_6085,N_5780,N_5950);
nor U6086 (N_6086,N_5872,N_5978);
or U6087 (N_6087,N_5887,N_5774);
nand U6088 (N_6088,N_5929,N_5841);
and U6089 (N_6089,N_5854,N_5814);
nand U6090 (N_6090,N_5885,N_5768);
or U6091 (N_6091,N_5925,N_5861);
or U6092 (N_6092,N_5811,N_5760);
xnor U6093 (N_6093,N_5977,N_5875);
nand U6094 (N_6094,N_5913,N_5965);
nor U6095 (N_6095,N_5845,N_5804);
xor U6096 (N_6096,N_5797,N_5910);
nor U6097 (N_6097,N_5958,N_5990);
or U6098 (N_6098,N_5901,N_5752);
nand U6099 (N_6099,N_5878,N_5813);
and U6100 (N_6100,N_5943,N_5753);
nand U6101 (N_6101,N_5859,N_5902);
or U6102 (N_6102,N_5949,N_5884);
and U6103 (N_6103,N_5758,N_5956);
xor U6104 (N_6104,N_5898,N_5937);
and U6105 (N_6105,N_5779,N_5795);
nand U6106 (N_6106,N_5764,N_5983);
or U6107 (N_6107,N_5830,N_5849);
nor U6108 (N_6108,N_5832,N_5893);
nor U6109 (N_6109,N_5855,N_5877);
or U6110 (N_6110,N_5909,N_5829);
xnor U6111 (N_6111,N_5765,N_5775);
or U6112 (N_6112,N_5888,N_5953);
nand U6113 (N_6113,N_5754,N_5890);
and U6114 (N_6114,N_5863,N_5915);
and U6115 (N_6115,N_5894,N_5969);
xor U6116 (N_6116,N_5933,N_5952);
nand U6117 (N_6117,N_5960,N_5984);
or U6118 (N_6118,N_5809,N_5919);
xor U6119 (N_6119,N_5846,N_5889);
xnor U6120 (N_6120,N_5975,N_5903);
xnor U6121 (N_6121,N_5970,N_5908);
xnor U6122 (N_6122,N_5869,N_5817);
or U6123 (N_6123,N_5905,N_5935);
xor U6124 (N_6124,N_5761,N_5892);
or U6125 (N_6125,N_5775,N_5771);
xor U6126 (N_6126,N_5865,N_5992);
or U6127 (N_6127,N_5979,N_5984);
nand U6128 (N_6128,N_5800,N_5791);
xnor U6129 (N_6129,N_5960,N_5861);
nor U6130 (N_6130,N_5803,N_5979);
xnor U6131 (N_6131,N_5844,N_5837);
nor U6132 (N_6132,N_5887,N_5998);
or U6133 (N_6133,N_5914,N_5750);
nand U6134 (N_6134,N_5878,N_5857);
nor U6135 (N_6135,N_5790,N_5999);
xnor U6136 (N_6136,N_5868,N_5861);
nor U6137 (N_6137,N_5799,N_5970);
and U6138 (N_6138,N_5752,N_5827);
nand U6139 (N_6139,N_5948,N_5847);
nor U6140 (N_6140,N_5836,N_5905);
nand U6141 (N_6141,N_5847,N_5862);
and U6142 (N_6142,N_5952,N_5864);
or U6143 (N_6143,N_5895,N_5925);
xor U6144 (N_6144,N_5872,N_5873);
nor U6145 (N_6145,N_5957,N_5951);
or U6146 (N_6146,N_5750,N_5816);
and U6147 (N_6147,N_5942,N_5815);
or U6148 (N_6148,N_5953,N_5972);
nor U6149 (N_6149,N_5766,N_5922);
or U6150 (N_6150,N_5912,N_5758);
or U6151 (N_6151,N_5837,N_5908);
nand U6152 (N_6152,N_5987,N_5768);
and U6153 (N_6153,N_5935,N_5992);
and U6154 (N_6154,N_5763,N_5797);
nor U6155 (N_6155,N_5793,N_5908);
nand U6156 (N_6156,N_5853,N_5889);
nor U6157 (N_6157,N_5761,N_5764);
or U6158 (N_6158,N_5933,N_5906);
nor U6159 (N_6159,N_5793,N_5936);
xor U6160 (N_6160,N_5963,N_5904);
and U6161 (N_6161,N_5757,N_5802);
nand U6162 (N_6162,N_5875,N_5894);
nand U6163 (N_6163,N_5832,N_5775);
xnor U6164 (N_6164,N_5779,N_5916);
nor U6165 (N_6165,N_5856,N_5813);
or U6166 (N_6166,N_5809,N_5887);
or U6167 (N_6167,N_5803,N_5763);
or U6168 (N_6168,N_5939,N_5853);
or U6169 (N_6169,N_5851,N_5884);
or U6170 (N_6170,N_5917,N_5956);
and U6171 (N_6171,N_5908,N_5933);
nand U6172 (N_6172,N_5852,N_5855);
xor U6173 (N_6173,N_5986,N_5916);
xor U6174 (N_6174,N_5857,N_5936);
xnor U6175 (N_6175,N_5903,N_5985);
nor U6176 (N_6176,N_5987,N_5751);
nor U6177 (N_6177,N_5778,N_5895);
xor U6178 (N_6178,N_5952,N_5782);
nor U6179 (N_6179,N_5869,N_5800);
or U6180 (N_6180,N_5828,N_5939);
and U6181 (N_6181,N_5986,N_5983);
nor U6182 (N_6182,N_5832,N_5804);
nand U6183 (N_6183,N_5779,N_5761);
nand U6184 (N_6184,N_5839,N_5893);
or U6185 (N_6185,N_5952,N_5823);
xor U6186 (N_6186,N_5986,N_5797);
nor U6187 (N_6187,N_5822,N_5758);
xor U6188 (N_6188,N_5778,N_5852);
or U6189 (N_6189,N_5958,N_5859);
and U6190 (N_6190,N_5925,N_5886);
nor U6191 (N_6191,N_5765,N_5983);
nor U6192 (N_6192,N_5779,N_5849);
and U6193 (N_6193,N_5786,N_5837);
and U6194 (N_6194,N_5890,N_5912);
and U6195 (N_6195,N_5988,N_5904);
or U6196 (N_6196,N_5961,N_5797);
xnor U6197 (N_6197,N_5894,N_5798);
or U6198 (N_6198,N_5902,N_5842);
nand U6199 (N_6199,N_5860,N_5996);
nand U6200 (N_6200,N_5973,N_5970);
and U6201 (N_6201,N_5958,N_5922);
nand U6202 (N_6202,N_5751,N_5808);
and U6203 (N_6203,N_5757,N_5904);
and U6204 (N_6204,N_5773,N_5765);
and U6205 (N_6205,N_5824,N_5939);
nand U6206 (N_6206,N_5772,N_5806);
or U6207 (N_6207,N_5871,N_5828);
nand U6208 (N_6208,N_5969,N_5931);
and U6209 (N_6209,N_5914,N_5884);
and U6210 (N_6210,N_5927,N_5786);
and U6211 (N_6211,N_5982,N_5906);
and U6212 (N_6212,N_5819,N_5826);
nor U6213 (N_6213,N_5925,N_5957);
xnor U6214 (N_6214,N_5909,N_5803);
xnor U6215 (N_6215,N_5961,N_5770);
nand U6216 (N_6216,N_5782,N_5979);
xor U6217 (N_6217,N_5826,N_5799);
xnor U6218 (N_6218,N_5862,N_5789);
or U6219 (N_6219,N_5847,N_5992);
nor U6220 (N_6220,N_5992,N_5896);
and U6221 (N_6221,N_5969,N_5911);
and U6222 (N_6222,N_5928,N_5794);
nand U6223 (N_6223,N_5984,N_5754);
nor U6224 (N_6224,N_5993,N_5975);
or U6225 (N_6225,N_5971,N_5792);
nor U6226 (N_6226,N_5969,N_5990);
or U6227 (N_6227,N_5882,N_5962);
or U6228 (N_6228,N_5907,N_5775);
nand U6229 (N_6229,N_5913,N_5907);
or U6230 (N_6230,N_5801,N_5950);
nor U6231 (N_6231,N_5827,N_5774);
nor U6232 (N_6232,N_5900,N_5954);
xor U6233 (N_6233,N_5953,N_5904);
or U6234 (N_6234,N_5867,N_5897);
nand U6235 (N_6235,N_5841,N_5907);
nand U6236 (N_6236,N_5966,N_5803);
or U6237 (N_6237,N_5796,N_5948);
xor U6238 (N_6238,N_5873,N_5968);
or U6239 (N_6239,N_5773,N_5803);
nand U6240 (N_6240,N_5939,N_5878);
xor U6241 (N_6241,N_5835,N_5783);
or U6242 (N_6242,N_5919,N_5836);
nor U6243 (N_6243,N_5997,N_5886);
or U6244 (N_6244,N_5988,N_5892);
xor U6245 (N_6245,N_5845,N_5899);
nor U6246 (N_6246,N_5799,N_5868);
nand U6247 (N_6247,N_5877,N_5968);
or U6248 (N_6248,N_5947,N_5981);
nand U6249 (N_6249,N_5959,N_5799);
and U6250 (N_6250,N_6121,N_6179);
xnor U6251 (N_6251,N_6102,N_6150);
or U6252 (N_6252,N_6117,N_6108);
nand U6253 (N_6253,N_6123,N_6238);
or U6254 (N_6254,N_6007,N_6120);
xnor U6255 (N_6255,N_6068,N_6057);
nand U6256 (N_6256,N_6138,N_6118);
nand U6257 (N_6257,N_6004,N_6223);
and U6258 (N_6258,N_6245,N_6033);
or U6259 (N_6259,N_6105,N_6205);
nand U6260 (N_6260,N_6030,N_6053);
xnor U6261 (N_6261,N_6008,N_6215);
or U6262 (N_6262,N_6106,N_6246);
xor U6263 (N_6263,N_6201,N_6147);
nor U6264 (N_6264,N_6186,N_6024);
or U6265 (N_6265,N_6097,N_6203);
and U6266 (N_6266,N_6211,N_6066);
and U6267 (N_6267,N_6141,N_6162);
xnor U6268 (N_6268,N_6222,N_6058);
nor U6269 (N_6269,N_6041,N_6200);
and U6270 (N_6270,N_6021,N_6192);
xor U6271 (N_6271,N_6137,N_6181);
nand U6272 (N_6272,N_6084,N_6166);
and U6273 (N_6273,N_6173,N_6175);
and U6274 (N_6274,N_6077,N_6226);
or U6275 (N_6275,N_6127,N_6026);
nand U6276 (N_6276,N_6048,N_6208);
and U6277 (N_6277,N_6159,N_6104);
and U6278 (N_6278,N_6047,N_6027);
or U6279 (N_6279,N_6195,N_6028);
or U6280 (N_6280,N_6210,N_6098);
and U6281 (N_6281,N_6091,N_6016);
nor U6282 (N_6282,N_6080,N_6038);
and U6283 (N_6283,N_6189,N_6235);
and U6284 (N_6284,N_6029,N_6229);
and U6285 (N_6285,N_6013,N_6221);
xnor U6286 (N_6286,N_6194,N_6193);
nor U6287 (N_6287,N_6003,N_6093);
nand U6288 (N_6288,N_6088,N_6202);
xor U6289 (N_6289,N_6163,N_6031);
and U6290 (N_6290,N_6144,N_6133);
and U6291 (N_6291,N_6050,N_6099);
nor U6292 (N_6292,N_6188,N_6178);
xnor U6293 (N_6293,N_6085,N_6051);
xor U6294 (N_6294,N_6247,N_6184);
nor U6295 (N_6295,N_6151,N_6236);
nor U6296 (N_6296,N_6190,N_6071);
xor U6297 (N_6297,N_6140,N_6002);
or U6298 (N_6298,N_6143,N_6227);
xnor U6299 (N_6299,N_6243,N_6185);
and U6300 (N_6300,N_6119,N_6055);
and U6301 (N_6301,N_6010,N_6040);
or U6302 (N_6302,N_6182,N_6165);
or U6303 (N_6303,N_6061,N_6191);
nand U6304 (N_6304,N_6213,N_6131);
nor U6305 (N_6305,N_6198,N_6220);
or U6306 (N_6306,N_6019,N_6239);
and U6307 (N_6307,N_6148,N_6241);
and U6308 (N_6308,N_6035,N_6012);
and U6309 (N_6309,N_6045,N_6153);
or U6310 (N_6310,N_6116,N_6103);
nand U6311 (N_6311,N_6204,N_6197);
or U6312 (N_6312,N_6096,N_6212);
xor U6313 (N_6313,N_6234,N_6072);
and U6314 (N_6314,N_6063,N_6078);
nand U6315 (N_6315,N_6124,N_6032);
and U6316 (N_6316,N_6042,N_6130);
xor U6317 (N_6317,N_6109,N_6139);
xnor U6318 (N_6318,N_6240,N_6218);
or U6319 (N_6319,N_6196,N_6017);
nand U6320 (N_6320,N_6064,N_6169);
nor U6321 (N_6321,N_6248,N_6217);
xnor U6322 (N_6322,N_6115,N_6237);
and U6323 (N_6323,N_6219,N_6230);
xnor U6324 (N_6324,N_6070,N_6225);
and U6325 (N_6325,N_6172,N_6060);
and U6326 (N_6326,N_6049,N_6065);
or U6327 (N_6327,N_6134,N_6039);
xor U6328 (N_6328,N_6152,N_6168);
nor U6329 (N_6329,N_6101,N_6009);
and U6330 (N_6330,N_6129,N_6224);
nor U6331 (N_6331,N_6054,N_6142);
and U6332 (N_6332,N_6110,N_6074);
nand U6333 (N_6333,N_6075,N_6136);
nor U6334 (N_6334,N_6037,N_6170);
nand U6335 (N_6335,N_6001,N_6231);
nor U6336 (N_6336,N_6107,N_6062);
or U6337 (N_6337,N_6244,N_6044);
nor U6338 (N_6338,N_6114,N_6125);
or U6339 (N_6339,N_6082,N_6034);
xnor U6340 (N_6340,N_6149,N_6086);
and U6341 (N_6341,N_6233,N_6059);
nand U6342 (N_6342,N_6087,N_6176);
nand U6343 (N_6343,N_6036,N_6014);
xor U6344 (N_6344,N_6135,N_6052);
nor U6345 (N_6345,N_6025,N_6083);
and U6346 (N_6346,N_6095,N_6160);
xor U6347 (N_6347,N_6122,N_6167);
or U6348 (N_6348,N_6164,N_6157);
nand U6349 (N_6349,N_6209,N_6011);
and U6350 (N_6350,N_6146,N_6092);
or U6351 (N_6351,N_6023,N_6177);
nand U6352 (N_6352,N_6022,N_6228);
nand U6353 (N_6353,N_6128,N_6111);
xnor U6354 (N_6354,N_6089,N_6020);
and U6355 (N_6355,N_6081,N_6079);
nand U6356 (N_6356,N_6249,N_6158);
and U6357 (N_6357,N_6067,N_6126);
and U6358 (N_6358,N_6069,N_6174);
or U6359 (N_6359,N_6171,N_6056);
nand U6360 (N_6360,N_6073,N_6132);
nand U6361 (N_6361,N_6183,N_6232);
xor U6362 (N_6362,N_6206,N_6216);
nand U6363 (N_6363,N_6161,N_6090);
nand U6364 (N_6364,N_6046,N_6155);
and U6365 (N_6365,N_6199,N_6156);
and U6366 (N_6366,N_6242,N_6076);
or U6367 (N_6367,N_6154,N_6112);
and U6368 (N_6368,N_6043,N_6018);
xnor U6369 (N_6369,N_6113,N_6005);
or U6370 (N_6370,N_6100,N_6207);
nand U6371 (N_6371,N_6000,N_6180);
and U6372 (N_6372,N_6145,N_6214);
xor U6373 (N_6373,N_6187,N_6006);
xor U6374 (N_6374,N_6094,N_6015);
or U6375 (N_6375,N_6218,N_6216);
nor U6376 (N_6376,N_6054,N_6118);
or U6377 (N_6377,N_6241,N_6202);
xor U6378 (N_6378,N_6248,N_6104);
nor U6379 (N_6379,N_6067,N_6092);
nor U6380 (N_6380,N_6110,N_6019);
or U6381 (N_6381,N_6234,N_6059);
and U6382 (N_6382,N_6243,N_6150);
and U6383 (N_6383,N_6146,N_6035);
nand U6384 (N_6384,N_6226,N_6020);
nand U6385 (N_6385,N_6135,N_6216);
xor U6386 (N_6386,N_6209,N_6171);
nand U6387 (N_6387,N_6152,N_6028);
and U6388 (N_6388,N_6013,N_6053);
xnor U6389 (N_6389,N_6038,N_6117);
and U6390 (N_6390,N_6039,N_6010);
or U6391 (N_6391,N_6001,N_6205);
nand U6392 (N_6392,N_6038,N_6132);
xnor U6393 (N_6393,N_6238,N_6207);
xnor U6394 (N_6394,N_6231,N_6120);
nor U6395 (N_6395,N_6188,N_6056);
or U6396 (N_6396,N_6078,N_6012);
nor U6397 (N_6397,N_6105,N_6212);
and U6398 (N_6398,N_6124,N_6114);
or U6399 (N_6399,N_6162,N_6117);
xnor U6400 (N_6400,N_6007,N_6143);
xnor U6401 (N_6401,N_6120,N_6023);
xnor U6402 (N_6402,N_6059,N_6054);
nand U6403 (N_6403,N_6090,N_6022);
and U6404 (N_6404,N_6210,N_6167);
and U6405 (N_6405,N_6099,N_6103);
xnor U6406 (N_6406,N_6058,N_6210);
xnor U6407 (N_6407,N_6204,N_6202);
nor U6408 (N_6408,N_6034,N_6212);
xnor U6409 (N_6409,N_6089,N_6126);
xor U6410 (N_6410,N_6139,N_6249);
or U6411 (N_6411,N_6017,N_6249);
nor U6412 (N_6412,N_6124,N_6174);
or U6413 (N_6413,N_6204,N_6037);
nand U6414 (N_6414,N_6221,N_6122);
or U6415 (N_6415,N_6050,N_6156);
nand U6416 (N_6416,N_6074,N_6132);
nor U6417 (N_6417,N_6032,N_6093);
or U6418 (N_6418,N_6170,N_6081);
nor U6419 (N_6419,N_6168,N_6171);
xor U6420 (N_6420,N_6216,N_6217);
or U6421 (N_6421,N_6246,N_6078);
xnor U6422 (N_6422,N_6000,N_6038);
nor U6423 (N_6423,N_6165,N_6044);
nand U6424 (N_6424,N_6012,N_6172);
or U6425 (N_6425,N_6034,N_6036);
or U6426 (N_6426,N_6183,N_6101);
nor U6427 (N_6427,N_6228,N_6105);
nand U6428 (N_6428,N_6041,N_6017);
xnor U6429 (N_6429,N_6081,N_6194);
and U6430 (N_6430,N_6064,N_6230);
or U6431 (N_6431,N_6099,N_6209);
nand U6432 (N_6432,N_6147,N_6002);
xnor U6433 (N_6433,N_6244,N_6157);
or U6434 (N_6434,N_6048,N_6173);
nor U6435 (N_6435,N_6224,N_6190);
or U6436 (N_6436,N_6217,N_6132);
and U6437 (N_6437,N_6102,N_6172);
xnor U6438 (N_6438,N_6201,N_6236);
or U6439 (N_6439,N_6171,N_6038);
xor U6440 (N_6440,N_6172,N_6147);
nand U6441 (N_6441,N_6112,N_6146);
and U6442 (N_6442,N_6217,N_6120);
xor U6443 (N_6443,N_6057,N_6049);
or U6444 (N_6444,N_6125,N_6241);
and U6445 (N_6445,N_6059,N_6203);
xnor U6446 (N_6446,N_6122,N_6090);
nand U6447 (N_6447,N_6109,N_6177);
or U6448 (N_6448,N_6244,N_6209);
or U6449 (N_6449,N_6247,N_6002);
and U6450 (N_6450,N_6098,N_6186);
nor U6451 (N_6451,N_6102,N_6137);
xnor U6452 (N_6452,N_6071,N_6082);
xnor U6453 (N_6453,N_6078,N_6182);
and U6454 (N_6454,N_6080,N_6215);
xnor U6455 (N_6455,N_6126,N_6170);
nor U6456 (N_6456,N_6048,N_6113);
and U6457 (N_6457,N_6029,N_6171);
xor U6458 (N_6458,N_6055,N_6132);
xor U6459 (N_6459,N_6089,N_6109);
nor U6460 (N_6460,N_6128,N_6066);
nor U6461 (N_6461,N_6094,N_6060);
and U6462 (N_6462,N_6194,N_6203);
nor U6463 (N_6463,N_6236,N_6199);
and U6464 (N_6464,N_6243,N_6007);
or U6465 (N_6465,N_6084,N_6076);
xnor U6466 (N_6466,N_6171,N_6085);
nor U6467 (N_6467,N_6209,N_6117);
xnor U6468 (N_6468,N_6130,N_6243);
xor U6469 (N_6469,N_6056,N_6164);
xor U6470 (N_6470,N_6033,N_6181);
and U6471 (N_6471,N_6026,N_6232);
nand U6472 (N_6472,N_6083,N_6011);
or U6473 (N_6473,N_6205,N_6215);
xnor U6474 (N_6474,N_6052,N_6099);
nand U6475 (N_6475,N_6157,N_6216);
nand U6476 (N_6476,N_6014,N_6175);
nand U6477 (N_6477,N_6123,N_6142);
or U6478 (N_6478,N_6204,N_6161);
and U6479 (N_6479,N_6188,N_6071);
nor U6480 (N_6480,N_6245,N_6194);
nand U6481 (N_6481,N_6101,N_6157);
nand U6482 (N_6482,N_6219,N_6040);
nor U6483 (N_6483,N_6180,N_6005);
nand U6484 (N_6484,N_6152,N_6140);
and U6485 (N_6485,N_6198,N_6111);
nand U6486 (N_6486,N_6175,N_6171);
or U6487 (N_6487,N_6026,N_6054);
xor U6488 (N_6488,N_6002,N_6028);
and U6489 (N_6489,N_6044,N_6149);
nand U6490 (N_6490,N_6047,N_6223);
nor U6491 (N_6491,N_6245,N_6241);
and U6492 (N_6492,N_6191,N_6171);
and U6493 (N_6493,N_6209,N_6010);
nor U6494 (N_6494,N_6120,N_6094);
xnor U6495 (N_6495,N_6101,N_6150);
nor U6496 (N_6496,N_6230,N_6148);
xor U6497 (N_6497,N_6033,N_6218);
nand U6498 (N_6498,N_6199,N_6050);
nand U6499 (N_6499,N_6072,N_6160);
nand U6500 (N_6500,N_6350,N_6328);
nor U6501 (N_6501,N_6375,N_6489);
or U6502 (N_6502,N_6292,N_6392);
nand U6503 (N_6503,N_6430,N_6408);
nor U6504 (N_6504,N_6391,N_6437);
nor U6505 (N_6505,N_6344,N_6379);
xnor U6506 (N_6506,N_6419,N_6455);
xor U6507 (N_6507,N_6323,N_6334);
nor U6508 (N_6508,N_6352,N_6409);
and U6509 (N_6509,N_6451,N_6368);
nor U6510 (N_6510,N_6441,N_6476);
nor U6511 (N_6511,N_6313,N_6376);
xnor U6512 (N_6512,N_6425,N_6257);
xor U6513 (N_6513,N_6499,N_6422);
xor U6514 (N_6514,N_6387,N_6351);
nand U6515 (N_6515,N_6343,N_6265);
and U6516 (N_6516,N_6278,N_6415);
xor U6517 (N_6517,N_6491,N_6370);
nand U6518 (N_6518,N_6464,N_6369);
and U6519 (N_6519,N_6268,N_6348);
nand U6520 (N_6520,N_6423,N_6367);
xnor U6521 (N_6521,N_6300,N_6453);
xor U6522 (N_6522,N_6452,N_6287);
and U6523 (N_6523,N_6250,N_6354);
xnor U6524 (N_6524,N_6373,N_6414);
nor U6525 (N_6525,N_6340,N_6438);
nand U6526 (N_6526,N_6450,N_6479);
nand U6527 (N_6527,N_6433,N_6311);
nand U6528 (N_6528,N_6478,N_6471);
nor U6529 (N_6529,N_6325,N_6283);
xor U6530 (N_6530,N_6332,N_6322);
nor U6531 (N_6531,N_6493,N_6255);
nor U6532 (N_6532,N_6293,N_6444);
and U6533 (N_6533,N_6458,N_6259);
nor U6534 (N_6534,N_6460,N_6400);
xor U6535 (N_6535,N_6318,N_6298);
nor U6536 (N_6536,N_6312,N_6289);
nor U6537 (N_6537,N_6411,N_6406);
and U6538 (N_6538,N_6429,N_6449);
xor U6539 (N_6539,N_6314,N_6389);
and U6540 (N_6540,N_6260,N_6333);
xnor U6541 (N_6541,N_6306,N_6412);
xor U6542 (N_6542,N_6290,N_6469);
or U6543 (N_6543,N_6277,N_6490);
nor U6544 (N_6544,N_6349,N_6362);
nor U6545 (N_6545,N_6345,N_6381);
and U6546 (N_6546,N_6299,N_6428);
and U6547 (N_6547,N_6434,N_6384);
nand U6548 (N_6548,N_6254,N_6463);
or U6549 (N_6549,N_6324,N_6439);
nand U6550 (N_6550,N_6273,N_6487);
nand U6551 (N_6551,N_6372,N_6468);
xnor U6552 (N_6552,N_6356,N_6473);
nand U6553 (N_6553,N_6341,N_6447);
xnor U6554 (N_6554,N_6303,N_6276);
or U6555 (N_6555,N_6302,N_6374);
xor U6556 (N_6556,N_6371,N_6363);
or U6557 (N_6557,N_6410,N_6456);
or U6558 (N_6558,N_6261,N_6398);
or U6559 (N_6559,N_6494,N_6316);
or U6560 (N_6560,N_6337,N_6294);
and U6561 (N_6561,N_6413,N_6359);
nor U6562 (N_6562,N_6485,N_6436);
or U6563 (N_6563,N_6421,N_6377);
xor U6564 (N_6564,N_6386,N_6495);
or U6565 (N_6565,N_6279,N_6467);
nand U6566 (N_6566,N_6420,N_6459);
xnor U6567 (N_6567,N_6383,N_6431);
nor U6568 (N_6568,N_6267,N_6427);
xnor U6569 (N_6569,N_6353,N_6317);
nor U6570 (N_6570,N_6329,N_6274);
xor U6571 (N_6571,N_6256,N_6264);
nor U6572 (N_6572,N_6321,N_6330);
and U6573 (N_6573,N_6393,N_6470);
nor U6574 (N_6574,N_6295,N_6364);
nor U6575 (N_6575,N_6315,N_6326);
xor U6576 (N_6576,N_6483,N_6390);
and U6577 (N_6577,N_6498,N_6327);
or U6578 (N_6578,N_6445,N_6440);
nand U6579 (N_6579,N_6358,N_6474);
nor U6580 (N_6580,N_6366,N_6484);
xor U6581 (N_6581,N_6401,N_6280);
nor U6582 (N_6582,N_6285,N_6380);
nand U6583 (N_6583,N_6272,N_6291);
nand U6584 (N_6584,N_6394,N_6403);
nor U6585 (N_6585,N_6397,N_6357);
and U6586 (N_6586,N_6395,N_6378);
or U6587 (N_6587,N_6480,N_6304);
or U6588 (N_6588,N_6461,N_6339);
and U6589 (N_6589,N_6307,N_6426);
nand U6590 (N_6590,N_6263,N_6405);
nor U6591 (N_6591,N_6488,N_6454);
or U6592 (N_6592,N_6336,N_6482);
nor U6593 (N_6593,N_6271,N_6432);
or U6594 (N_6594,N_6331,N_6472);
nor U6595 (N_6595,N_6262,N_6416);
or U6596 (N_6596,N_6481,N_6275);
nand U6597 (N_6597,N_6308,N_6443);
and U6598 (N_6598,N_6270,N_6266);
nor U6599 (N_6599,N_6346,N_6385);
or U6600 (N_6600,N_6497,N_6269);
and U6601 (N_6601,N_6281,N_6342);
or U6602 (N_6602,N_6301,N_6396);
and U6603 (N_6603,N_6388,N_6492);
nor U6604 (N_6604,N_6465,N_6407);
nor U6605 (N_6605,N_6399,N_6296);
xor U6606 (N_6606,N_6442,N_6338);
xnor U6607 (N_6607,N_6310,N_6462);
and U6608 (N_6608,N_6404,N_6347);
nand U6609 (N_6609,N_6496,N_6286);
xor U6610 (N_6610,N_6417,N_6335);
or U6611 (N_6611,N_6402,N_6365);
nand U6612 (N_6612,N_6360,N_6486);
nand U6613 (N_6613,N_6309,N_6253);
xor U6614 (N_6614,N_6424,N_6252);
xnor U6615 (N_6615,N_6466,N_6446);
xnor U6616 (N_6616,N_6258,N_6457);
or U6617 (N_6617,N_6288,N_6355);
or U6618 (N_6618,N_6361,N_6320);
and U6619 (N_6619,N_6435,N_6305);
xor U6620 (N_6620,N_6251,N_6477);
nand U6621 (N_6621,N_6282,N_6475);
and U6622 (N_6622,N_6297,N_6448);
nand U6623 (N_6623,N_6418,N_6382);
and U6624 (N_6624,N_6319,N_6284);
and U6625 (N_6625,N_6495,N_6429);
xor U6626 (N_6626,N_6302,N_6494);
xor U6627 (N_6627,N_6358,N_6323);
nand U6628 (N_6628,N_6254,N_6480);
xnor U6629 (N_6629,N_6280,N_6480);
nand U6630 (N_6630,N_6256,N_6432);
or U6631 (N_6631,N_6431,N_6307);
or U6632 (N_6632,N_6318,N_6334);
nand U6633 (N_6633,N_6340,N_6341);
xor U6634 (N_6634,N_6392,N_6475);
and U6635 (N_6635,N_6258,N_6488);
and U6636 (N_6636,N_6289,N_6268);
nor U6637 (N_6637,N_6433,N_6495);
xor U6638 (N_6638,N_6433,N_6422);
xor U6639 (N_6639,N_6367,N_6495);
nor U6640 (N_6640,N_6274,N_6484);
nor U6641 (N_6641,N_6368,N_6347);
xor U6642 (N_6642,N_6290,N_6260);
and U6643 (N_6643,N_6397,N_6372);
or U6644 (N_6644,N_6339,N_6466);
nor U6645 (N_6645,N_6440,N_6402);
xnor U6646 (N_6646,N_6473,N_6274);
nor U6647 (N_6647,N_6391,N_6295);
xor U6648 (N_6648,N_6412,N_6439);
or U6649 (N_6649,N_6385,N_6457);
nand U6650 (N_6650,N_6470,N_6494);
nand U6651 (N_6651,N_6376,N_6494);
and U6652 (N_6652,N_6409,N_6454);
nor U6653 (N_6653,N_6469,N_6372);
xnor U6654 (N_6654,N_6363,N_6336);
xnor U6655 (N_6655,N_6349,N_6460);
nor U6656 (N_6656,N_6349,N_6344);
nor U6657 (N_6657,N_6426,N_6488);
nand U6658 (N_6658,N_6375,N_6469);
nor U6659 (N_6659,N_6469,N_6488);
nand U6660 (N_6660,N_6459,N_6391);
nand U6661 (N_6661,N_6392,N_6306);
or U6662 (N_6662,N_6476,N_6290);
nand U6663 (N_6663,N_6385,N_6393);
and U6664 (N_6664,N_6354,N_6334);
or U6665 (N_6665,N_6336,N_6346);
nor U6666 (N_6666,N_6358,N_6439);
or U6667 (N_6667,N_6386,N_6261);
xnor U6668 (N_6668,N_6350,N_6321);
nor U6669 (N_6669,N_6324,N_6274);
xor U6670 (N_6670,N_6362,N_6268);
xor U6671 (N_6671,N_6473,N_6457);
and U6672 (N_6672,N_6310,N_6444);
nor U6673 (N_6673,N_6477,N_6421);
nor U6674 (N_6674,N_6376,N_6446);
nand U6675 (N_6675,N_6392,N_6410);
xnor U6676 (N_6676,N_6439,N_6378);
and U6677 (N_6677,N_6311,N_6361);
and U6678 (N_6678,N_6460,N_6292);
nor U6679 (N_6679,N_6379,N_6403);
or U6680 (N_6680,N_6327,N_6358);
xor U6681 (N_6681,N_6498,N_6456);
and U6682 (N_6682,N_6374,N_6481);
xnor U6683 (N_6683,N_6371,N_6279);
and U6684 (N_6684,N_6379,N_6276);
xnor U6685 (N_6685,N_6286,N_6452);
xnor U6686 (N_6686,N_6396,N_6349);
or U6687 (N_6687,N_6403,N_6404);
or U6688 (N_6688,N_6330,N_6326);
and U6689 (N_6689,N_6498,N_6272);
xor U6690 (N_6690,N_6371,N_6393);
or U6691 (N_6691,N_6278,N_6478);
nand U6692 (N_6692,N_6273,N_6331);
nand U6693 (N_6693,N_6498,N_6440);
or U6694 (N_6694,N_6267,N_6426);
nor U6695 (N_6695,N_6379,N_6314);
and U6696 (N_6696,N_6447,N_6327);
xor U6697 (N_6697,N_6286,N_6413);
xor U6698 (N_6698,N_6295,N_6352);
or U6699 (N_6699,N_6328,N_6378);
xor U6700 (N_6700,N_6260,N_6451);
or U6701 (N_6701,N_6482,N_6274);
or U6702 (N_6702,N_6395,N_6252);
xnor U6703 (N_6703,N_6390,N_6284);
nand U6704 (N_6704,N_6480,N_6460);
or U6705 (N_6705,N_6328,N_6304);
or U6706 (N_6706,N_6431,N_6376);
or U6707 (N_6707,N_6383,N_6322);
xor U6708 (N_6708,N_6491,N_6440);
nand U6709 (N_6709,N_6434,N_6404);
and U6710 (N_6710,N_6407,N_6355);
xnor U6711 (N_6711,N_6336,N_6308);
or U6712 (N_6712,N_6481,N_6477);
nor U6713 (N_6713,N_6429,N_6374);
nor U6714 (N_6714,N_6323,N_6348);
nand U6715 (N_6715,N_6403,N_6464);
nand U6716 (N_6716,N_6451,N_6295);
nand U6717 (N_6717,N_6328,N_6479);
or U6718 (N_6718,N_6368,N_6399);
or U6719 (N_6719,N_6471,N_6464);
nor U6720 (N_6720,N_6284,N_6295);
nor U6721 (N_6721,N_6459,N_6318);
nand U6722 (N_6722,N_6277,N_6486);
nand U6723 (N_6723,N_6329,N_6499);
and U6724 (N_6724,N_6330,N_6294);
or U6725 (N_6725,N_6448,N_6362);
nand U6726 (N_6726,N_6315,N_6495);
nor U6727 (N_6727,N_6270,N_6355);
nor U6728 (N_6728,N_6401,N_6377);
xor U6729 (N_6729,N_6257,N_6390);
nand U6730 (N_6730,N_6288,N_6386);
nor U6731 (N_6731,N_6431,N_6461);
and U6732 (N_6732,N_6450,N_6349);
or U6733 (N_6733,N_6464,N_6270);
xnor U6734 (N_6734,N_6401,N_6477);
or U6735 (N_6735,N_6252,N_6488);
nor U6736 (N_6736,N_6313,N_6327);
nor U6737 (N_6737,N_6403,N_6300);
nand U6738 (N_6738,N_6400,N_6465);
nor U6739 (N_6739,N_6481,N_6394);
xor U6740 (N_6740,N_6268,N_6458);
xnor U6741 (N_6741,N_6338,N_6420);
xnor U6742 (N_6742,N_6377,N_6462);
nand U6743 (N_6743,N_6286,N_6260);
or U6744 (N_6744,N_6265,N_6422);
nor U6745 (N_6745,N_6319,N_6396);
and U6746 (N_6746,N_6480,N_6322);
nor U6747 (N_6747,N_6363,N_6400);
nand U6748 (N_6748,N_6269,N_6311);
or U6749 (N_6749,N_6471,N_6281);
xnor U6750 (N_6750,N_6525,N_6726);
nand U6751 (N_6751,N_6538,N_6563);
nand U6752 (N_6752,N_6744,N_6618);
and U6753 (N_6753,N_6747,N_6518);
or U6754 (N_6754,N_6580,N_6748);
nand U6755 (N_6755,N_6697,N_6643);
nand U6756 (N_6756,N_6520,N_6621);
nor U6757 (N_6757,N_6590,N_6646);
nor U6758 (N_6758,N_6729,N_6708);
xor U6759 (N_6759,N_6584,N_6619);
or U6760 (N_6760,N_6540,N_6698);
nor U6761 (N_6761,N_6572,N_6651);
nor U6762 (N_6762,N_6608,N_6661);
and U6763 (N_6763,N_6675,N_6672);
xor U6764 (N_6764,N_6735,N_6534);
nor U6765 (N_6765,N_6571,N_6719);
nor U6766 (N_6766,N_6533,N_6693);
and U6767 (N_6767,N_6705,N_6650);
nor U6768 (N_6768,N_6596,N_6712);
or U6769 (N_6769,N_6567,N_6669);
xor U6770 (N_6770,N_6718,N_6657);
or U6771 (N_6771,N_6600,N_6516);
xnor U6772 (N_6772,N_6691,N_6521);
nand U6773 (N_6773,N_6677,N_6599);
nor U6774 (N_6774,N_6615,N_6656);
nor U6775 (N_6775,N_6736,N_6545);
and U6776 (N_6776,N_6720,N_6676);
or U6777 (N_6777,N_6586,N_6562);
or U6778 (N_6778,N_6611,N_6550);
nor U6779 (N_6779,N_6523,N_6522);
nor U6780 (N_6780,N_6542,N_6555);
and U6781 (N_6781,N_6631,N_6713);
xor U6782 (N_6782,N_6589,N_6566);
and U6783 (N_6783,N_6653,N_6727);
or U6784 (N_6784,N_6606,N_6527);
nand U6785 (N_6785,N_6728,N_6695);
nand U6786 (N_6786,N_6696,N_6711);
nand U6787 (N_6787,N_6535,N_6641);
and U6788 (N_6788,N_6707,N_6612);
or U6789 (N_6789,N_6548,N_6616);
xor U6790 (N_6790,N_6579,N_6725);
and U6791 (N_6791,N_6620,N_6577);
nor U6792 (N_6792,N_6687,N_6724);
nand U6793 (N_6793,N_6660,N_6554);
nor U6794 (N_6794,N_6515,N_6674);
nor U6795 (N_6795,N_6528,N_6565);
xor U6796 (N_6796,N_6564,N_6664);
and U6797 (N_6797,N_6625,N_6742);
or U6798 (N_6798,N_6671,N_6624);
and U6799 (N_6799,N_6723,N_6578);
nor U6800 (N_6800,N_6541,N_6721);
nor U6801 (N_6801,N_6576,N_6630);
nand U6802 (N_6802,N_6716,N_6617);
nor U6803 (N_6803,N_6574,N_6610);
nor U6804 (N_6804,N_6613,N_6678);
nand U6805 (N_6805,N_6680,N_6501);
and U6806 (N_6806,N_6598,N_6570);
nor U6807 (N_6807,N_6614,N_6642);
or U6808 (N_6808,N_6588,N_6645);
nor U6809 (N_6809,N_6667,N_6526);
xnor U6810 (N_6810,N_6623,N_6591);
nand U6811 (N_6811,N_6536,N_6551);
nor U6812 (N_6812,N_6530,N_6595);
nand U6813 (N_6813,N_6573,N_6581);
xnor U6814 (N_6814,N_6670,N_6517);
or U6815 (N_6815,N_6634,N_6597);
and U6816 (N_6816,N_6635,N_6512);
xor U6817 (N_6817,N_6605,N_6604);
nor U6818 (N_6818,N_6734,N_6544);
or U6819 (N_6819,N_6741,N_6547);
and U6820 (N_6820,N_6640,N_6513);
nor U6821 (N_6821,N_6583,N_6668);
nor U6822 (N_6822,N_6694,N_6717);
nor U6823 (N_6823,N_6568,N_6737);
xor U6824 (N_6824,N_6706,N_6585);
xnor U6825 (N_6825,N_6684,N_6704);
xor U6826 (N_6826,N_6637,N_6593);
nor U6827 (N_6827,N_6638,N_6663);
and U6828 (N_6828,N_6560,N_6594);
xor U6829 (N_6829,N_6529,N_6685);
or U6830 (N_6830,N_6662,N_6519);
nor U6831 (N_6831,N_6587,N_6592);
or U6832 (N_6832,N_6602,N_6556);
and U6833 (N_6833,N_6561,N_6699);
xnor U6834 (N_6834,N_6689,N_6703);
nor U6835 (N_6835,N_6553,N_6649);
nand U6836 (N_6836,N_6733,N_6739);
nor U6837 (N_6837,N_6692,N_6731);
and U6838 (N_6838,N_6652,N_6537);
xor U6839 (N_6839,N_6681,N_6508);
and U6840 (N_6840,N_6557,N_6509);
nand U6841 (N_6841,N_6506,N_6607);
xor U6842 (N_6842,N_6507,N_6546);
and U6843 (N_6843,N_6552,N_6673);
or U6844 (N_6844,N_6732,N_6505);
or U6845 (N_6845,N_6730,N_6715);
or U6846 (N_6846,N_6683,N_6665);
or U6847 (N_6847,N_6743,N_6629);
or U6848 (N_6848,N_6666,N_6738);
and U6849 (N_6849,N_6647,N_6644);
nand U6850 (N_6850,N_6558,N_6510);
or U6851 (N_6851,N_6633,N_6745);
nor U6852 (N_6852,N_6682,N_6648);
nand U6853 (N_6853,N_6601,N_6688);
and U6854 (N_6854,N_6749,N_6569);
or U6855 (N_6855,N_6514,N_6655);
xor U6856 (N_6856,N_6549,N_6740);
and U6857 (N_6857,N_6502,N_6659);
or U6858 (N_6858,N_6622,N_6679);
nor U6859 (N_6859,N_6700,N_6582);
nor U6860 (N_6860,N_6511,N_6543);
xor U6861 (N_6861,N_6654,N_6559);
nand U6862 (N_6862,N_6627,N_6746);
and U6863 (N_6863,N_6709,N_6710);
and U6864 (N_6864,N_6609,N_6722);
xor U6865 (N_6865,N_6690,N_6714);
nand U6866 (N_6866,N_6701,N_6500);
nor U6867 (N_6867,N_6504,N_6632);
xnor U6868 (N_6868,N_6636,N_6626);
nor U6869 (N_6869,N_6639,N_6658);
xor U6870 (N_6870,N_6524,N_6686);
and U6871 (N_6871,N_6532,N_6575);
nor U6872 (N_6872,N_6603,N_6628);
and U6873 (N_6873,N_6702,N_6539);
and U6874 (N_6874,N_6503,N_6531);
nand U6875 (N_6875,N_6652,N_6686);
or U6876 (N_6876,N_6702,N_6564);
nor U6877 (N_6877,N_6670,N_6587);
nor U6878 (N_6878,N_6679,N_6597);
xor U6879 (N_6879,N_6644,N_6608);
or U6880 (N_6880,N_6524,N_6550);
xor U6881 (N_6881,N_6594,N_6749);
and U6882 (N_6882,N_6585,N_6697);
nor U6883 (N_6883,N_6619,N_6747);
nor U6884 (N_6884,N_6587,N_6584);
nor U6885 (N_6885,N_6746,N_6738);
or U6886 (N_6886,N_6749,N_6519);
or U6887 (N_6887,N_6736,N_6708);
or U6888 (N_6888,N_6652,N_6608);
or U6889 (N_6889,N_6723,N_6715);
and U6890 (N_6890,N_6721,N_6641);
nand U6891 (N_6891,N_6668,N_6630);
nor U6892 (N_6892,N_6643,N_6743);
or U6893 (N_6893,N_6601,N_6629);
and U6894 (N_6894,N_6542,N_6625);
or U6895 (N_6895,N_6728,N_6521);
xnor U6896 (N_6896,N_6692,N_6717);
nor U6897 (N_6897,N_6555,N_6652);
nand U6898 (N_6898,N_6740,N_6623);
nand U6899 (N_6899,N_6682,N_6638);
xor U6900 (N_6900,N_6669,N_6716);
nor U6901 (N_6901,N_6608,N_6501);
or U6902 (N_6902,N_6613,N_6723);
nor U6903 (N_6903,N_6578,N_6683);
and U6904 (N_6904,N_6715,N_6641);
or U6905 (N_6905,N_6592,N_6656);
or U6906 (N_6906,N_6702,N_6698);
or U6907 (N_6907,N_6648,N_6633);
or U6908 (N_6908,N_6552,N_6557);
nor U6909 (N_6909,N_6555,N_6737);
or U6910 (N_6910,N_6572,N_6664);
or U6911 (N_6911,N_6597,N_6532);
nor U6912 (N_6912,N_6687,N_6535);
and U6913 (N_6913,N_6668,N_6639);
nor U6914 (N_6914,N_6646,N_6509);
xor U6915 (N_6915,N_6638,N_6571);
and U6916 (N_6916,N_6561,N_6711);
or U6917 (N_6917,N_6628,N_6677);
and U6918 (N_6918,N_6604,N_6715);
nand U6919 (N_6919,N_6654,N_6504);
and U6920 (N_6920,N_6558,N_6603);
nand U6921 (N_6921,N_6641,N_6542);
or U6922 (N_6922,N_6690,N_6678);
xor U6923 (N_6923,N_6589,N_6671);
nor U6924 (N_6924,N_6549,N_6596);
or U6925 (N_6925,N_6559,N_6524);
nand U6926 (N_6926,N_6587,N_6570);
xor U6927 (N_6927,N_6652,N_6506);
xnor U6928 (N_6928,N_6637,N_6707);
and U6929 (N_6929,N_6553,N_6571);
nand U6930 (N_6930,N_6620,N_6598);
nand U6931 (N_6931,N_6741,N_6530);
nor U6932 (N_6932,N_6720,N_6541);
or U6933 (N_6933,N_6662,N_6520);
xor U6934 (N_6934,N_6510,N_6688);
nand U6935 (N_6935,N_6516,N_6532);
or U6936 (N_6936,N_6705,N_6696);
nand U6937 (N_6937,N_6588,N_6621);
or U6938 (N_6938,N_6620,N_6541);
nor U6939 (N_6939,N_6525,N_6635);
nor U6940 (N_6940,N_6573,N_6588);
nor U6941 (N_6941,N_6604,N_6693);
nand U6942 (N_6942,N_6527,N_6627);
nor U6943 (N_6943,N_6748,N_6725);
or U6944 (N_6944,N_6716,N_6711);
xor U6945 (N_6945,N_6598,N_6665);
xnor U6946 (N_6946,N_6612,N_6518);
or U6947 (N_6947,N_6526,N_6598);
nor U6948 (N_6948,N_6737,N_6652);
nand U6949 (N_6949,N_6548,N_6604);
or U6950 (N_6950,N_6585,N_6635);
or U6951 (N_6951,N_6701,N_6573);
or U6952 (N_6952,N_6563,N_6527);
and U6953 (N_6953,N_6592,N_6713);
nor U6954 (N_6954,N_6643,N_6728);
nor U6955 (N_6955,N_6584,N_6734);
and U6956 (N_6956,N_6747,N_6550);
and U6957 (N_6957,N_6515,N_6653);
and U6958 (N_6958,N_6618,N_6679);
and U6959 (N_6959,N_6601,N_6697);
nand U6960 (N_6960,N_6696,N_6551);
nand U6961 (N_6961,N_6599,N_6521);
and U6962 (N_6962,N_6520,N_6629);
nor U6963 (N_6963,N_6747,N_6567);
nor U6964 (N_6964,N_6659,N_6656);
or U6965 (N_6965,N_6520,N_6640);
nand U6966 (N_6966,N_6647,N_6589);
or U6967 (N_6967,N_6719,N_6537);
nand U6968 (N_6968,N_6594,N_6708);
nand U6969 (N_6969,N_6598,N_6529);
and U6970 (N_6970,N_6503,N_6707);
or U6971 (N_6971,N_6597,N_6625);
xnor U6972 (N_6972,N_6675,N_6517);
xor U6973 (N_6973,N_6512,N_6738);
and U6974 (N_6974,N_6622,N_6735);
or U6975 (N_6975,N_6585,N_6738);
xnor U6976 (N_6976,N_6659,N_6714);
or U6977 (N_6977,N_6646,N_6639);
nor U6978 (N_6978,N_6718,N_6727);
nand U6979 (N_6979,N_6667,N_6657);
and U6980 (N_6980,N_6684,N_6541);
and U6981 (N_6981,N_6507,N_6576);
xor U6982 (N_6982,N_6650,N_6597);
and U6983 (N_6983,N_6739,N_6667);
or U6984 (N_6984,N_6654,N_6547);
nor U6985 (N_6985,N_6519,N_6544);
xnor U6986 (N_6986,N_6745,N_6610);
xor U6987 (N_6987,N_6717,N_6660);
nand U6988 (N_6988,N_6509,N_6592);
and U6989 (N_6989,N_6644,N_6556);
xor U6990 (N_6990,N_6634,N_6637);
nand U6991 (N_6991,N_6624,N_6724);
and U6992 (N_6992,N_6662,N_6581);
or U6993 (N_6993,N_6626,N_6660);
nand U6994 (N_6994,N_6543,N_6742);
nor U6995 (N_6995,N_6595,N_6694);
nand U6996 (N_6996,N_6569,N_6737);
and U6997 (N_6997,N_6640,N_6511);
or U6998 (N_6998,N_6661,N_6746);
and U6999 (N_6999,N_6624,N_6742);
xnor U7000 (N_7000,N_6971,N_6862);
and U7001 (N_7001,N_6963,N_6762);
xor U7002 (N_7002,N_6975,N_6968);
nor U7003 (N_7003,N_6863,N_6997);
xor U7004 (N_7004,N_6918,N_6754);
xnor U7005 (N_7005,N_6846,N_6869);
and U7006 (N_7006,N_6905,N_6803);
nor U7007 (N_7007,N_6893,N_6857);
and U7008 (N_7008,N_6945,N_6995);
and U7009 (N_7009,N_6937,N_6881);
nor U7010 (N_7010,N_6779,N_6976);
nand U7011 (N_7011,N_6960,N_6850);
xor U7012 (N_7012,N_6909,N_6777);
xnor U7013 (N_7013,N_6885,N_6994);
nor U7014 (N_7014,N_6787,N_6900);
nor U7015 (N_7015,N_6821,N_6864);
nor U7016 (N_7016,N_6922,N_6855);
and U7017 (N_7017,N_6987,N_6914);
nand U7018 (N_7018,N_6891,N_6983);
xor U7019 (N_7019,N_6956,N_6982);
xnor U7020 (N_7020,N_6886,N_6797);
or U7021 (N_7021,N_6770,N_6887);
nand U7022 (N_7022,N_6940,N_6890);
nand U7023 (N_7023,N_6888,N_6868);
nor U7024 (N_7024,N_6843,N_6782);
xor U7025 (N_7025,N_6932,N_6829);
nor U7026 (N_7026,N_6751,N_6841);
or U7027 (N_7027,N_6959,N_6839);
nor U7028 (N_7028,N_6854,N_6974);
and U7029 (N_7029,N_6783,N_6969);
nor U7030 (N_7030,N_6808,N_6773);
and U7031 (N_7031,N_6828,N_6876);
xnor U7032 (N_7032,N_6904,N_6800);
and U7033 (N_7033,N_6820,N_6965);
nor U7034 (N_7034,N_6830,N_6894);
nand U7035 (N_7035,N_6992,N_6840);
and U7036 (N_7036,N_6877,N_6906);
nand U7037 (N_7037,N_6798,N_6812);
xor U7038 (N_7038,N_6834,N_6842);
or U7039 (N_7039,N_6913,N_6757);
xor U7040 (N_7040,N_6756,N_6896);
nand U7041 (N_7041,N_6824,N_6813);
and U7042 (N_7042,N_6933,N_6851);
nand U7043 (N_7043,N_6935,N_6996);
nor U7044 (N_7044,N_6753,N_6921);
or U7045 (N_7045,N_6993,N_6815);
nor U7046 (N_7046,N_6871,N_6819);
and U7047 (N_7047,N_6837,N_6845);
xnor U7048 (N_7048,N_6925,N_6826);
nand U7049 (N_7049,N_6926,N_6929);
or U7050 (N_7050,N_6786,N_6832);
or U7051 (N_7051,N_6949,N_6912);
nor U7052 (N_7052,N_6818,N_6883);
and U7053 (N_7053,N_6985,N_6973);
and U7054 (N_7054,N_6953,N_6936);
or U7055 (N_7055,N_6989,N_6768);
xnor U7056 (N_7056,N_6774,N_6916);
nand U7057 (N_7057,N_6970,N_6990);
nand U7058 (N_7058,N_6991,N_6908);
or U7059 (N_7059,N_6972,N_6796);
and U7060 (N_7060,N_6814,N_6930);
nor U7061 (N_7061,N_6827,N_6811);
nor U7062 (N_7062,N_6875,N_6942);
xnor U7063 (N_7063,N_6898,N_6934);
or U7064 (N_7064,N_6957,N_6946);
nor U7065 (N_7065,N_6833,N_6810);
and U7066 (N_7066,N_6804,N_6785);
nor U7067 (N_7067,N_6999,N_6944);
and U7068 (N_7068,N_6984,N_6852);
nand U7069 (N_7069,N_6809,N_6859);
and U7070 (N_7070,N_6867,N_6941);
and U7071 (N_7071,N_6923,N_6790);
and U7072 (N_7072,N_6943,N_6853);
and U7073 (N_7073,N_6766,N_6761);
and U7074 (N_7074,N_6977,N_6924);
nand U7075 (N_7075,N_6865,N_6870);
and U7076 (N_7076,N_6895,N_6788);
nand U7077 (N_7077,N_6781,N_6831);
xnor U7078 (N_7078,N_6866,N_6901);
or U7079 (N_7079,N_6772,N_6806);
nor U7080 (N_7080,N_6759,N_6873);
nor U7081 (N_7081,N_6807,N_6849);
nor U7082 (N_7082,N_6817,N_6801);
or U7083 (N_7083,N_6775,N_6879);
and U7084 (N_7084,N_6795,N_6789);
xnor U7085 (N_7085,N_6917,N_6948);
nor U7086 (N_7086,N_6920,N_6836);
or U7087 (N_7087,N_6791,N_6799);
xnor U7088 (N_7088,N_6950,N_6882);
xor U7089 (N_7089,N_6771,N_6980);
or U7090 (N_7090,N_6765,N_6958);
xnor U7091 (N_7091,N_6897,N_6884);
nor U7092 (N_7092,N_6858,N_6928);
xor U7093 (N_7093,N_6915,N_6910);
nor U7094 (N_7094,N_6961,N_6793);
or U7095 (N_7095,N_6874,N_6880);
nor U7096 (N_7096,N_6760,N_6986);
nor U7097 (N_7097,N_6776,N_6805);
nand U7098 (N_7098,N_6794,N_6769);
nand U7099 (N_7099,N_6750,N_6872);
nor U7100 (N_7100,N_6954,N_6861);
nand U7101 (N_7101,N_6899,N_6998);
xnor U7102 (N_7102,N_6902,N_6767);
and U7103 (N_7103,N_6784,N_6878);
and U7104 (N_7104,N_6823,N_6802);
nand U7105 (N_7105,N_6938,N_6979);
or U7106 (N_7106,N_6955,N_6838);
xnor U7107 (N_7107,N_6927,N_6752);
nand U7108 (N_7108,N_6892,N_6981);
nor U7109 (N_7109,N_6763,N_6844);
nor U7110 (N_7110,N_6758,N_6856);
xnor U7111 (N_7111,N_6903,N_6911);
nor U7112 (N_7112,N_6835,N_6848);
or U7113 (N_7113,N_6978,N_6951);
or U7114 (N_7114,N_6778,N_6947);
and U7115 (N_7115,N_6816,N_6780);
or U7116 (N_7116,N_6847,N_6939);
or U7117 (N_7117,N_6966,N_6962);
or U7118 (N_7118,N_6860,N_6967);
xnor U7119 (N_7119,N_6792,N_6988);
nand U7120 (N_7120,N_6825,N_6931);
or U7121 (N_7121,N_6907,N_6919);
xnor U7122 (N_7122,N_6764,N_6822);
and U7123 (N_7123,N_6964,N_6952);
and U7124 (N_7124,N_6889,N_6755);
nor U7125 (N_7125,N_6986,N_6869);
or U7126 (N_7126,N_6940,N_6848);
nand U7127 (N_7127,N_6898,N_6860);
xnor U7128 (N_7128,N_6896,N_6816);
and U7129 (N_7129,N_6771,N_6968);
and U7130 (N_7130,N_6923,N_6918);
and U7131 (N_7131,N_6968,N_6900);
nand U7132 (N_7132,N_6965,N_6810);
and U7133 (N_7133,N_6804,N_6839);
nand U7134 (N_7134,N_6753,N_6999);
xnor U7135 (N_7135,N_6903,N_6910);
nor U7136 (N_7136,N_6849,N_6841);
or U7137 (N_7137,N_6936,N_6870);
nor U7138 (N_7138,N_6852,N_6848);
xor U7139 (N_7139,N_6838,N_6822);
xnor U7140 (N_7140,N_6942,N_6911);
or U7141 (N_7141,N_6811,N_6942);
or U7142 (N_7142,N_6811,N_6981);
and U7143 (N_7143,N_6868,N_6955);
or U7144 (N_7144,N_6960,N_6956);
and U7145 (N_7145,N_6910,N_6808);
nor U7146 (N_7146,N_6838,N_6842);
nor U7147 (N_7147,N_6931,N_6886);
nand U7148 (N_7148,N_6942,N_6923);
nor U7149 (N_7149,N_6758,N_6976);
or U7150 (N_7150,N_6920,N_6925);
or U7151 (N_7151,N_6821,N_6869);
and U7152 (N_7152,N_6756,N_6948);
xnor U7153 (N_7153,N_6874,N_6873);
nor U7154 (N_7154,N_6926,N_6881);
nor U7155 (N_7155,N_6916,N_6838);
nor U7156 (N_7156,N_6997,N_6862);
or U7157 (N_7157,N_6787,N_6908);
and U7158 (N_7158,N_6953,N_6995);
and U7159 (N_7159,N_6914,N_6985);
nand U7160 (N_7160,N_6811,N_6878);
nand U7161 (N_7161,N_6783,N_6764);
nor U7162 (N_7162,N_6953,N_6954);
or U7163 (N_7163,N_6834,N_6831);
or U7164 (N_7164,N_6824,N_6941);
xnor U7165 (N_7165,N_6895,N_6946);
nand U7166 (N_7166,N_6981,N_6983);
or U7167 (N_7167,N_6796,N_6783);
nand U7168 (N_7168,N_6810,N_6944);
or U7169 (N_7169,N_6937,N_6790);
or U7170 (N_7170,N_6983,N_6976);
or U7171 (N_7171,N_6861,N_6774);
nand U7172 (N_7172,N_6899,N_6909);
xor U7173 (N_7173,N_6997,N_6872);
or U7174 (N_7174,N_6900,N_6783);
nand U7175 (N_7175,N_6780,N_6877);
nor U7176 (N_7176,N_6907,N_6984);
nor U7177 (N_7177,N_6918,N_6834);
nor U7178 (N_7178,N_6788,N_6928);
nand U7179 (N_7179,N_6950,N_6939);
and U7180 (N_7180,N_6912,N_6924);
nor U7181 (N_7181,N_6790,N_6887);
nor U7182 (N_7182,N_6938,N_6754);
and U7183 (N_7183,N_6845,N_6978);
nand U7184 (N_7184,N_6958,N_6752);
or U7185 (N_7185,N_6987,N_6974);
xor U7186 (N_7186,N_6822,N_6863);
xnor U7187 (N_7187,N_6910,N_6835);
nand U7188 (N_7188,N_6952,N_6777);
xor U7189 (N_7189,N_6891,N_6914);
nor U7190 (N_7190,N_6925,N_6767);
xnor U7191 (N_7191,N_6870,N_6962);
and U7192 (N_7192,N_6991,N_6765);
and U7193 (N_7193,N_6760,N_6771);
and U7194 (N_7194,N_6923,N_6969);
and U7195 (N_7195,N_6876,N_6781);
nor U7196 (N_7196,N_6856,N_6977);
nor U7197 (N_7197,N_6953,N_6832);
or U7198 (N_7198,N_6754,N_6861);
xnor U7199 (N_7199,N_6950,N_6883);
nor U7200 (N_7200,N_6775,N_6961);
and U7201 (N_7201,N_6860,N_6828);
nand U7202 (N_7202,N_6946,N_6898);
or U7203 (N_7203,N_6866,N_6752);
nor U7204 (N_7204,N_6907,N_6899);
xnor U7205 (N_7205,N_6750,N_6876);
xnor U7206 (N_7206,N_6807,N_6835);
or U7207 (N_7207,N_6826,N_6831);
nand U7208 (N_7208,N_6766,N_6795);
and U7209 (N_7209,N_6926,N_6763);
nand U7210 (N_7210,N_6902,N_6956);
nor U7211 (N_7211,N_6976,N_6936);
nand U7212 (N_7212,N_6973,N_6986);
xor U7213 (N_7213,N_6931,N_6967);
or U7214 (N_7214,N_6821,N_6992);
nor U7215 (N_7215,N_6871,N_6905);
and U7216 (N_7216,N_6769,N_6913);
nand U7217 (N_7217,N_6912,N_6997);
and U7218 (N_7218,N_6959,N_6754);
or U7219 (N_7219,N_6751,N_6852);
and U7220 (N_7220,N_6939,N_6967);
nor U7221 (N_7221,N_6938,N_6785);
nand U7222 (N_7222,N_6900,N_6884);
and U7223 (N_7223,N_6767,N_6819);
or U7224 (N_7224,N_6975,N_6845);
xor U7225 (N_7225,N_6929,N_6918);
and U7226 (N_7226,N_6954,N_6768);
nor U7227 (N_7227,N_6953,N_6870);
nand U7228 (N_7228,N_6956,N_6828);
nand U7229 (N_7229,N_6835,N_6968);
nor U7230 (N_7230,N_6795,N_6833);
nor U7231 (N_7231,N_6890,N_6793);
nand U7232 (N_7232,N_6839,N_6879);
or U7233 (N_7233,N_6938,N_6861);
or U7234 (N_7234,N_6808,N_6863);
xor U7235 (N_7235,N_6852,N_6944);
xnor U7236 (N_7236,N_6750,N_6763);
xnor U7237 (N_7237,N_6866,N_6862);
or U7238 (N_7238,N_6944,N_6965);
and U7239 (N_7239,N_6873,N_6903);
and U7240 (N_7240,N_6937,N_6750);
nand U7241 (N_7241,N_6891,N_6966);
xor U7242 (N_7242,N_6846,N_6918);
nand U7243 (N_7243,N_6803,N_6765);
nor U7244 (N_7244,N_6907,N_6854);
xnor U7245 (N_7245,N_6950,N_6965);
and U7246 (N_7246,N_6945,N_6948);
nand U7247 (N_7247,N_6882,N_6793);
or U7248 (N_7248,N_6820,N_6783);
nor U7249 (N_7249,N_6918,N_6766);
nor U7250 (N_7250,N_7152,N_7026);
xor U7251 (N_7251,N_7000,N_7079);
nor U7252 (N_7252,N_7247,N_7175);
nand U7253 (N_7253,N_7093,N_7211);
nor U7254 (N_7254,N_7246,N_7006);
or U7255 (N_7255,N_7065,N_7146);
nor U7256 (N_7256,N_7237,N_7208);
and U7257 (N_7257,N_7126,N_7084);
xor U7258 (N_7258,N_7077,N_7060);
and U7259 (N_7259,N_7180,N_7119);
or U7260 (N_7260,N_7091,N_7103);
and U7261 (N_7261,N_7094,N_7241);
nand U7262 (N_7262,N_7234,N_7131);
or U7263 (N_7263,N_7020,N_7159);
xnor U7264 (N_7264,N_7117,N_7161);
and U7265 (N_7265,N_7043,N_7243);
xor U7266 (N_7266,N_7074,N_7036);
or U7267 (N_7267,N_7073,N_7014);
nor U7268 (N_7268,N_7068,N_7071);
and U7269 (N_7269,N_7013,N_7133);
nand U7270 (N_7270,N_7024,N_7156);
nand U7271 (N_7271,N_7238,N_7193);
and U7272 (N_7272,N_7029,N_7199);
nor U7273 (N_7273,N_7099,N_7142);
and U7274 (N_7274,N_7213,N_7169);
xor U7275 (N_7275,N_7039,N_7197);
xor U7276 (N_7276,N_7177,N_7053);
nor U7277 (N_7277,N_7127,N_7107);
and U7278 (N_7278,N_7108,N_7138);
and U7279 (N_7279,N_7087,N_7198);
or U7280 (N_7280,N_7100,N_7232);
and U7281 (N_7281,N_7139,N_7233);
or U7282 (N_7282,N_7166,N_7225);
or U7283 (N_7283,N_7002,N_7188);
nand U7284 (N_7284,N_7128,N_7012);
or U7285 (N_7285,N_7048,N_7104);
nor U7286 (N_7286,N_7248,N_7151);
or U7287 (N_7287,N_7185,N_7105);
and U7288 (N_7288,N_7003,N_7172);
nand U7289 (N_7289,N_7042,N_7049);
nand U7290 (N_7290,N_7196,N_7217);
and U7291 (N_7291,N_7192,N_7171);
nor U7292 (N_7292,N_7102,N_7052);
nor U7293 (N_7293,N_7222,N_7106);
or U7294 (N_7294,N_7207,N_7101);
nor U7295 (N_7295,N_7227,N_7044);
and U7296 (N_7296,N_7118,N_7130);
nand U7297 (N_7297,N_7057,N_7158);
and U7298 (N_7298,N_7230,N_7097);
and U7299 (N_7299,N_7219,N_7007);
or U7300 (N_7300,N_7150,N_7132);
nor U7301 (N_7301,N_7019,N_7096);
xnor U7302 (N_7302,N_7215,N_7113);
or U7303 (N_7303,N_7037,N_7178);
nand U7304 (N_7304,N_7210,N_7163);
nor U7305 (N_7305,N_7212,N_7228);
nand U7306 (N_7306,N_7083,N_7155);
and U7307 (N_7307,N_7162,N_7129);
and U7308 (N_7308,N_7027,N_7201);
or U7309 (N_7309,N_7203,N_7038);
or U7310 (N_7310,N_7009,N_7010);
or U7311 (N_7311,N_7125,N_7051);
nor U7312 (N_7312,N_7160,N_7229);
and U7313 (N_7313,N_7183,N_7147);
nor U7314 (N_7314,N_7045,N_7109);
nand U7315 (N_7315,N_7040,N_7056);
xnor U7316 (N_7316,N_7242,N_7184);
and U7317 (N_7317,N_7182,N_7022);
xor U7318 (N_7318,N_7124,N_7004);
nand U7319 (N_7319,N_7135,N_7218);
xnor U7320 (N_7320,N_7011,N_7194);
and U7321 (N_7321,N_7008,N_7224);
or U7322 (N_7322,N_7168,N_7174);
nand U7323 (N_7323,N_7157,N_7055);
nand U7324 (N_7324,N_7112,N_7016);
xnor U7325 (N_7325,N_7017,N_7145);
nor U7326 (N_7326,N_7110,N_7114);
nand U7327 (N_7327,N_7240,N_7186);
or U7328 (N_7328,N_7245,N_7078);
nor U7329 (N_7329,N_7081,N_7041);
nand U7330 (N_7330,N_7064,N_7220);
xnor U7331 (N_7331,N_7033,N_7115);
nor U7332 (N_7332,N_7095,N_7085);
nand U7333 (N_7333,N_7070,N_7216);
or U7334 (N_7334,N_7137,N_7058);
and U7335 (N_7335,N_7090,N_7062);
and U7336 (N_7336,N_7116,N_7173);
nand U7337 (N_7337,N_7120,N_7189);
xor U7338 (N_7338,N_7140,N_7195);
xor U7339 (N_7339,N_7167,N_7221);
xor U7340 (N_7340,N_7021,N_7059);
nor U7341 (N_7341,N_7206,N_7209);
nor U7342 (N_7342,N_7072,N_7050);
xor U7343 (N_7343,N_7214,N_7176);
nand U7344 (N_7344,N_7136,N_7165);
nor U7345 (N_7345,N_7231,N_7089);
nand U7346 (N_7346,N_7069,N_7067);
nor U7347 (N_7347,N_7144,N_7066);
nand U7348 (N_7348,N_7005,N_7149);
nand U7349 (N_7349,N_7153,N_7098);
xnor U7350 (N_7350,N_7028,N_7200);
xnor U7351 (N_7351,N_7204,N_7082);
xor U7352 (N_7352,N_7170,N_7080);
nand U7353 (N_7353,N_7123,N_7205);
or U7354 (N_7354,N_7025,N_7179);
xor U7355 (N_7355,N_7030,N_7244);
and U7356 (N_7356,N_7236,N_7046);
nor U7357 (N_7357,N_7035,N_7154);
nor U7358 (N_7358,N_7223,N_7034);
and U7359 (N_7359,N_7061,N_7023);
or U7360 (N_7360,N_7181,N_7202);
nand U7361 (N_7361,N_7063,N_7141);
nand U7362 (N_7362,N_7032,N_7191);
nor U7363 (N_7363,N_7047,N_7235);
nor U7364 (N_7364,N_7134,N_7143);
and U7365 (N_7365,N_7088,N_7121);
or U7366 (N_7366,N_7075,N_7239);
or U7367 (N_7367,N_7054,N_7018);
and U7368 (N_7368,N_7187,N_7148);
nand U7369 (N_7369,N_7001,N_7086);
xnor U7370 (N_7370,N_7190,N_7249);
nor U7371 (N_7371,N_7122,N_7031);
and U7372 (N_7372,N_7226,N_7076);
nor U7373 (N_7373,N_7092,N_7111);
or U7374 (N_7374,N_7015,N_7164);
and U7375 (N_7375,N_7058,N_7182);
nor U7376 (N_7376,N_7238,N_7119);
nand U7377 (N_7377,N_7134,N_7111);
xnor U7378 (N_7378,N_7091,N_7222);
or U7379 (N_7379,N_7186,N_7068);
or U7380 (N_7380,N_7214,N_7211);
and U7381 (N_7381,N_7193,N_7172);
nor U7382 (N_7382,N_7035,N_7008);
xor U7383 (N_7383,N_7025,N_7116);
nor U7384 (N_7384,N_7059,N_7237);
xor U7385 (N_7385,N_7068,N_7207);
nand U7386 (N_7386,N_7035,N_7072);
xnor U7387 (N_7387,N_7241,N_7124);
and U7388 (N_7388,N_7028,N_7137);
nand U7389 (N_7389,N_7106,N_7112);
xnor U7390 (N_7390,N_7004,N_7018);
xor U7391 (N_7391,N_7009,N_7191);
nand U7392 (N_7392,N_7028,N_7237);
nand U7393 (N_7393,N_7013,N_7143);
nor U7394 (N_7394,N_7083,N_7065);
nor U7395 (N_7395,N_7189,N_7016);
nor U7396 (N_7396,N_7045,N_7074);
or U7397 (N_7397,N_7203,N_7139);
xnor U7398 (N_7398,N_7140,N_7185);
nor U7399 (N_7399,N_7018,N_7097);
nand U7400 (N_7400,N_7085,N_7153);
nor U7401 (N_7401,N_7104,N_7004);
or U7402 (N_7402,N_7116,N_7175);
or U7403 (N_7403,N_7141,N_7155);
or U7404 (N_7404,N_7030,N_7069);
or U7405 (N_7405,N_7228,N_7025);
and U7406 (N_7406,N_7244,N_7111);
nor U7407 (N_7407,N_7063,N_7205);
nor U7408 (N_7408,N_7114,N_7072);
nor U7409 (N_7409,N_7178,N_7057);
or U7410 (N_7410,N_7241,N_7143);
and U7411 (N_7411,N_7006,N_7242);
xor U7412 (N_7412,N_7056,N_7146);
nor U7413 (N_7413,N_7243,N_7018);
xor U7414 (N_7414,N_7090,N_7225);
and U7415 (N_7415,N_7249,N_7219);
and U7416 (N_7416,N_7052,N_7243);
nor U7417 (N_7417,N_7220,N_7145);
nand U7418 (N_7418,N_7008,N_7222);
xnor U7419 (N_7419,N_7184,N_7016);
and U7420 (N_7420,N_7239,N_7235);
nand U7421 (N_7421,N_7191,N_7057);
and U7422 (N_7422,N_7076,N_7241);
xor U7423 (N_7423,N_7237,N_7042);
nand U7424 (N_7424,N_7038,N_7175);
or U7425 (N_7425,N_7039,N_7173);
and U7426 (N_7426,N_7138,N_7184);
nor U7427 (N_7427,N_7028,N_7202);
xnor U7428 (N_7428,N_7087,N_7240);
nand U7429 (N_7429,N_7070,N_7114);
and U7430 (N_7430,N_7171,N_7100);
and U7431 (N_7431,N_7111,N_7004);
nand U7432 (N_7432,N_7244,N_7102);
nand U7433 (N_7433,N_7099,N_7083);
nor U7434 (N_7434,N_7143,N_7073);
xnor U7435 (N_7435,N_7155,N_7128);
and U7436 (N_7436,N_7196,N_7101);
or U7437 (N_7437,N_7070,N_7149);
or U7438 (N_7438,N_7232,N_7205);
nand U7439 (N_7439,N_7159,N_7052);
and U7440 (N_7440,N_7132,N_7166);
nand U7441 (N_7441,N_7226,N_7173);
nor U7442 (N_7442,N_7034,N_7099);
nand U7443 (N_7443,N_7105,N_7022);
xor U7444 (N_7444,N_7192,N_7187);
nand U7445 (N_7445,N_7118,N_7041);
nor U7446 (N_7446,N_7146,N_7122);
nor U7447 (N_7447,N_7211,N_7009);
nand U7448 (N_7448,N_7243,N_7150);
nor U7449 (N_7449,N_7012,N_7176);
nand U7450 (N_7450,N_7211,N_7240);
nor U7451 (N_7451,N_7071,N_7011);
or U7452 (N_7452,N_7094,N_7078);
nor U7453 (N_7453,N_7108,N_7021);
and U7454 (N_7454,N_7249,N_7176);
nor U7455 (N_7455,N_7127,N_7063);
nor U7456 (N_7456,N_7001,N_7170);
and U7457 (N_7457,N_7071,N_7219);
xnor U7458 (N_7458,N_7019,N_7023);
nand U7459 (N_7459,N_7115,N_7072);
nor U7460 (N_7460,N_7058,N_7178);
nor U7461 (N_7461,N_7223,N_7072);
xor U7462 (N_7462,N_7080,N_7213);
or U7463 (N_7463,N_7171,N_7224);
xnor U7464 (N_7464,N_7151,N_7088);
or U7465 (N_7465,N_7044,N_7205);
xnor U7466 (N_7466,N_7169,N_7160);
or U7467 (N_7467,N_7129,N_7015);
xnor U7468 (N_7468,N_7178,N_7007);
nand U7469 (N_7469,N_7190,N_7058);
or U7470 (N_7470,N_7224,N_7099);
xnor U7471 (N_7471,N_7169,N_7086);
xnor U7472 (N_7472,N_7019,N_7083);
xnor U7473 (N_7473,N_7154,N_7162);
nor U7474 (N_7474,N_7147,N_7113);
and U7475 (N_7475,N_7043,N_7113);
xnor U7476 (N_7476,N_7014,N_7136);
nand U7477 (N_7477,N_7063,N_7189);
nand U7478 (N_7478,N_7011,N_7191);
and U7479 (N_7479,N_7071,N_7039);
or U7480 (N_7480,N_7081,N_7169);
nand U7481 (N_7481,N_7074,N_7008);
xor U7482 (N_7482,N_7200,N_7187);
or U7483 (N_7483,N_7045,N_7137);
xnor U7484 (N_7484,N_7118,N_7044);
or U7485 (N_7485,N_7208,N_7090);
xnor U7486 (N_7486,N_7152,N_7083);
nand U7487 (N_7487,N_7124,N_7182);
and U7488 (N_7488,N_7127,N_7026);
nand U7489 (N_7489,N_7137,N_7146);
xor U7490 (N_7490,N_7246,N_7130);
xnor U7491 (N_7491,N_7205,N_7169);
and U7492 (N_7492,N_7168,N_7157);
nor U7493 (N_7493,N_7005,N_7230);
and U7494 (N_7494,N_7108,N_7073);
and U7495 (N_7495,N_7105,N_7204);
nor U7496 (N_7496,N_7149,N_7137);
xor U7497 (N_7497,N_7235,N_7084);
or U7498 (N_7498,N_7011,N_7066);
or U7499 (N_7499,N_7056,N_7033);
and U7500 (N_7500,N_7490,N_7432);
nor U7501 (N_7501,N_7437,N_7403);
xor U7502 (N_7502,N_7347,N_7274);
and U7503 (N_7503,N_7445,N_7389);
nand U7504 (N_7504,N_7329,N_7325);
nand U7505 (N_7505,N_7472,N_7435);
nor U7506 (N_7506,N_7280,N_7380);
or U7507 (N_7507,N_7310,N_7302);
and U7508 (N_7508,N_7335,N_7273);
xnor U7509 (N_7509,N_7355,N_7478);
xnor U7510 (N_7510,N_7456,N_7311);
nand U7511 (N_7511,N_7486,N_7346);
xor U7512 (N_7512,N_7305,N_7365);
nand U7513 (N_7513,N_7284,N_7308);
nor U7514 (N_7514,N_7339,N_7290);
or U7515 (N_7515,N_7266,N_7261);
xor U7516 (N_7516,N_7301,N_7295);
nand U7517 (N_7517,N_7373,N_7444);
nand U7518 (N_7518,N_7425,N_7470);
nor U7519 (N_7519,N_7353,N_7326);
nor U7520 (N_7520,N_7477,N_7297);
or U7521 (N_7521,N_7336,N_7383);
nor U7522 (N_7522,N_7367,N_7372);
nand U7523 (N_7523,N_7277,N_7361);
or U7524 (N_7524,N_7420,N_7475);
and U7525 (N_7525,N_7312,N_7495);
or U7526 (N_7526,N_7322,N_7250);
or U7527 (N_7527,N_7251,N_7492);
or U7528 (N_7528,N_7263,N_7345);
nor U7529 (N_7529,N_7471,N_7344);
or U7530 (N_7530,N_7357,N_7438);
and U7531 (N_7531,N_7262,N_7315);
nor U7532 (N_7532,N_7334,N_7374);
and U7533 (N_7533,N_7417,N_7340);
and U7534 (N_7534,N_7466,N_7453);
nor U7535 (N_7535,N_7482,N_7451);
nand U7536 (N_7536,N_7410,N_7377);
or U7537 (N_7537,N_7309,N_7426);
xnor U7538 (N_7538,N_7396,N_7491);
xnor U7539 (N_7539,N_7256,N_7480);
xnor U7540 (N_7540,N_7378,N_7272);
and U7541 (N_7541,N_7441,N_7348);
nor U7542 (N_7542,N_7499,N_7293);
nor U7543 (N_7543,N_7342,N_7269);
nand U7544 (N_7544,N_7370,N_7300);
and U7545 (N_7545,N_7418,N_7321);
and U7546 (N_7546,N_7427,N_7257);
and U7547 (N_7547,N_7288,N_7488);
nand U7548 (N_7548,N_7497,N_7462);
nand U7549 (N_7549,N_7398,N_7366);
nand U7550 (N_7550,N_7494,N_7255);
nand U7551 (N_7551,N_7258,N_7327);
or U7552 (N_7552,N_7376,N_7406);
xor U7553 (N_7553,N_7292,N_7448);
nand U7554 (N_7554,N_7281,N_7413);
nor U7555 (N_7555,N_7415,N_7414);
nor U7556 (N_7556,N_7304,N_7333);
or U7557 (N_7557,N_7400,N_7464);
nor U7558 (N_7558,N_7287,N_7276);
and U7559 (N_7559,N_7351,N_7469);
and U7560 (N_7560,N_7375,N_7465);
xnor U7561 (N_7561,N_7449,N_7254);
nand U7562 (N_7562,N_7299,N_7401);
or U7563 (N_7563,N_7496,N_7397);
nand U7564 (N_7564,N_7419,N_7363);
xor U7565 (N_7565,N_7461,N_7384);
and U7566 (N_7566,N_7298,N_7433);
nor U7567 (N_7567,N_7473,N_7468);
or U7568 (N_7568,N_7393,N_7303);
nand U7569 (N_7569,N_7423,N_7289);
or U7570 (N_7570,N_7368,N_7364);
nand U7571 (N_7571,N_7404,N_7382);
xor U7572 (N_7572,N_7463,N_7493);
nor U7573 (N_7573,N_7307,N_7314);
or U7574 (N_7574,N_7442,N_7253);
nor U7575 (N_7575,N_7294,N_7362);
nor U7576 (N_7576,N_7324,N_7474);
xor U7577 (N_7577,N_7291,N_7411);
nand U7578 (N_7578,N_7429,N_7391);
nor U7579 (N_7579,N_7316,N_7369);
or U7580 (N_7580,N_7422,N_7479);
or U7581 (N_7581,N_7428,N_7407);
or U7582 (N_7582,N_7430,N_7436);
nand U7583 (N_7583,N_7271,N_7265);
and U7584 (N_7584,N_7350,N_7476);
nand U7585 (N_7585,N_7358,N_7412);
and U7586 (N_7586,N_7498,N_7330);
or U7587 (N_7587,N_7278,N_7359);
nand U7588 (N_7588,N_7343,N_7318);
nor U7589 (N_7589,N_7439,N_7447);
or U7590 (N_7590,N_7421,N_7483);
nor U7591 (N_7591,N_7431,N_7338);
xor U7592 (N_7592,N_7408,N_7328);
and U7593 (N_7593,N_7306,N_7268);
or U7594 (N_7594,N_7454,N_7450);
xnor U7595 (N_7595,N_7405,N_7352);
or U7596 (N_7596,N_7286,N_7388);
or U7597 (N_7597,N_7260,N_7481);
nand U7598 (N_7598,N_7455,N_7337);
nand U7599 (N_7599,N_7387,N_7296);
and U7600 (N_7600,N_7484,N_7489);
xor U7601 (N_7601,N_7341,N_7267);
xnor U7602 (N_7602,N_7385,N_7381);
nor U7603 (N_7603,N_7440,N_7457);
nor U7604 (N_7604,N_7424,N_7264);
nor U7605 (N_7605,N_7392,N_7459);
and U7606 (N_7606,N_7275,N_7416);
or U7607 (N_7607,N_7467,N_7331);
nor U7608 (N_7608,N_7446,N_7319);
nor U7609 (N_7609,N_7458,N_7356);
xnor U7610 (N_7610,N_7390,N_7434);
xnor U7611 (N_7611,N_7452,N_7460);
nor U7612 (N_7612,N_7379,N_7443);
or U7613 (N_7613,N_7402,N_7320);
or U7614 (N_7614,N_7394,N_7349);
and U7615 (N_7615,N_7409,N_7386);
and U7616 (N_7616,N_7270,N_7279);
nor U7617 (N_7617,N_7485,N_7313);
or U7618 (N_7618,N_7252,N_7317);
nand U7619 (N_7619,N_7283,N_7399);
or U7620 (N_7620,N_7332,N_7360);
and U7621 (N_7621,N_7395,N_7323);
or U7622 (N_7622,N_7487,N_7282);
nor U7623 (N_7623,N_7259,N_7354);
nor U7624 (N_7624,N_7371,N_7285);
xor U7625 (N_7625,N_7297,N_7449);
or U7626 (N_7626,N_7275,N_7378);
nand U7627 (N_7627,N_7396,N_7281);
nor U7628 (N_7628,N_7339,N_7250);
or U7629 (N_7629,N_7334,N_7403);
nand U7630 (N_7630,N_7301,N_7386);
nor U7631 (N_7631,N_7469,N_7490);
nand U7632 (N_7632,N_7495,N_7374);
and U7633 (N_7633,N_7348,N_7437);
or U7634 (N_7634,N_7413,N_7450);
xnor U7635 (N_7635,N_7459,N_7380);
nor U7636 (N_7636,N_7464,N_7284);
nand U7637 (N_7637,N_7490,N_7423);
nor U7638 (N_7638,N_7477,N_7499);
nand U7639 (N_7639,N_7330,N_7259);
nand U7640 (N_7640,N_7321,N_7389);
or U7641 (N_7641,N_7354,N_7297);
nand U7642 (N_7642,N_7428,N_7465);
or U7643 (N_7643,N_7377,N_7396);
nand U7644 (N_7644,N_7265,N_7341);
or U7645 (N_7645,N_7419,N_7308);
or U7646 (N_7646,N_7335,N_7323);
or U7647 (N_7647,N_7396,N_7486);
or U7648 (N_7648,N_7320,N_7289);
xor U7649 (N_7649,N_7405,N_7251);
and U7650 (N_7650,N_7324,N_7461);
nand U7651 (N_7651,N_7372,N_7259);
nand U7652 (N_7652,N_7324,N_7321);
and U7653 (N_7653,N_7260,N_7369);
and U7654 (N_7654,N_7332,N_7370);
nor U7655 (N_7655,N_7464,N_7422);
xnor U7656 (N_7656,N_7389,N_7402);
nor U7657 (N_7657,N_7301,N_7424);
and U7658 (N_7658,N_7399,N_7296);
and U7659 (N_7659,N_7290,N_7264);
and U7660 (N_7660,N_7467,N_7352);
or U7661 (N_7661,N_7386,N_7314);
and U7662 (N_7662,N_7484,N_7336);
and U7663 (N_7663,N_7488,N_7403);
nand U7664 (N_7664,N_7333,N_7483);
xor U7665 (N_7665,N_7394,N_7364);
xor U7666 (N_7666,N_7364,N_7280);
and U7667 (N_7667,N_7420,N_7311);
and U7668 (N_7668,N_7406,N_7325);
nor U7669 (N_7669,N_7470,N_7371);
nor U7670 (N_7670,N_7476,N_7401);
nand U7671 (N_7671,N_7404,N_7337);
xnor U7672 (N_7672,N_7361,N_7421);
or U7673 (N_7673,N_7451,N_7307);
and U7674 (N_7674,N_7275,N_7302);
and U7675 (N_7675,N_7496,N_7280);
xor U7676 (N_7676,N_7299,N_7284);
nor U7677 (N_7677,N_7457,N_7338);
and U7678 (N_7678,N_7367,N_7473);
xor U7679 (N_7679,N_7307,N_7354);
or U7680 (N_7680,N_7302,N_7264);
or U7681 (N_7681,N_7490,N_7439);
or U7682 (N_7682,N_7294,N_7439);
and U7683 (N_7683,N_7498,N_7471);
or U7684 (N_7684,N_7274,N_7428);
nand U7685 (N_7685,N_7295,N_7481);
and U7686 (N_7686,N_7318,N_7309);
or U7687 (N_7687,N_7320,N_7419);
xnor U7688 (N_7688,N_7251,N_7404);
or U7689 (N_7689,N_7458,N_7391);
nor U7690 (N_7690,N_7388,N_7306);
nand U7691 (N_7691,N_7355,N_7404);
nand U7692 (N_7692,N_7416,N_7474);
nor U7693 (N_7693,N_7306,N_7313);
and U7694 (N_7694,N_7388,N_7311);
xnor U7695 (N_7695,N_7267,N_7435);
nor U7696 (N_7696,N_7353,N_7354);
nand U7697 (N_7697,N_7333,N_7316);
nor U7698 (N_7698,N_7440,N_7306);
nand U7699 (N_7699,N_7485,N_7257);
nand U7700 (N_7700,N_7329,N_7385);
and U7701 (N_7701,N_7285,N_7389);
nand U7702 (N_7702,N_7365,N_7373);
nor U7703 (N_7703,N_7470,N_7411);
nand U7704 (N_7704,N_7324,N_7363);
nor U7705 (N_7705,N_7302,N_7306);
nor U7706 (N_7706,N_7443,N_7338);
and U7707 (N_7707,N_7458,N_7291);
xor U7708 (N_7708,N_7386,N_7271);
and U7709 (N_7709,N_7470,N_7283);
nor U7710 (N_7710,N_7465,N_7488);
and U7711 (N_7711,N_7255,N_7498);
nand U7712 (N_7712,N_7303,N_7293);
and U7713 (N_7713,N_7254,N_7453);
nand U7714 (N_7714,N_7297,N_7278);
and U7715 (N_7715,N_7482,N_7280);
nand U7716 (N_7716,N_7336,N_7417);
xor U7717 (N_7717,N_7327,N_7369);
nor U7718 (N_7718,N_7372,N_7348);
nor U7719 (N_7719,N_7329,N_7271);
xor U7720 (N_7720,N_7387,N_7428);
nand U7721 (N_7721,N_7353,N_7336);
xor U7722 (N_7722,N_7352,N_7324);
or U7723 (N_7723,N_7432,N_7291);
nand U7724 (N_7724,N_7429,N_7403);
or U7725 (N_7725,N_7455,N_7435);
nand U7726 (N_7726,N_7385,N_7362);
xnor U7727 (N_7727,N_7256,N_7427);
nor U7728 (N_7728,N_7283,N_7280);
nor U7729 (N_7729,N_7426,N_7253);
or U7730 (N_7730,N_7368,N_7251);
xor U7731 (N_7731,N_7364,N_7272);
and U7732 (N_7732,N_7274,N_7293);
or U7733 (N_7733,N_7414,N_7356);
xnor U7734 (N_7734,N_7404,N_7317);
xor U7735 (N_7735,N_7350,N_7342);
or U7736 (N_7736,N_7381,N_7396);
xnor U7737 (N_7737,N_7388,N_7299);
nor U7738 (N_7738,N_7462,N_7280);
nor U7739 (N_7739,N_7390,N_7466);
and U7740 (N_7740,N_7431,N_7426);
nor U7741 (N_7741,N_7272,N_7484);
xor U7742 (N_7742,N_7474,N_7421);
nor U7743 (N_7743,N_7303,N_7387);
nor U7744 (N_7744,N_7259,N_7285);
xnor U7745 (N_7745,N_7402,N_7463);
nand U7746 (N_7746,N_7480,N_7381);
nand U7747 (N_7747,N_7345,N_7357);
and U7748 (N_7748,N_7489,N_7458);
nor U7749 (N_7749,N_7273,N_7416);
xnor U7750 (N_7750,N_7658,N_7632);
nor U7751 (N_7751,N_7707,N_7645);
xor U7752 (N_7752,N_7605,N_7693);
or U7753 (N_7753,N_7612,N_7502);
nor U7754 (N_7754,N_7536,N_7634);
nor U7755 (N_7755,N_7582,N_7557);
and U7756 (N_7756,N_7747,N_7734);
or U7757 (N_7757,N_7699,N_7679);
nor U7758 (N_7758,N_7709,N_7508);
nand U7759 (N_7759,N_7712,N_7691);
and U7760 (N_7760,N_7588,N_7501);
nand U7761 (N_7761,N_7542,N_7677);
nor U7762 (N_7762,N_7676,N_7506);
nand U7763 (N_7763,N_7720,N_7638);
nor U7764 (N_7764,N_7597,N_7731);
nand U7765 (N_7765,N_7668,N_7581);
or U7766 (N_7766,N_7559,N_7655);
xor U7767 (N_7767,N_7606,N_7546);
or U7768 (N_7768,N_7579,N_7533);
or U7769 (N_7769,N_7613,N_7610);
nand U7770 (N_7770,N_7555,N_7721);
xor U7771 (N_7771,N_7578,N_7548);
and U7772 (N_7772,N_7526,N_7656);
and U7773 (N_7773,N_7552,N_7729);
and U7774 (N_7774,N_7585,N_7692);
and U7775 (N_7775,N_7637,N_7619);
and U7776 (N_7776,N_7620,N_7730);
xor U7777 (N_7777,N_7737,N_7618);
nand U7778 (N_7778,N_7544,N_7689);
and U7779 (N_7779,N_7512,N_7701);
nand U7780 (N_7780,N_7621,N_7703);
xnor U7781 (N_7781,N_7684,N_7617);
nand U7782 (N_7782,N_7696,N_7706);
nand U7783 (N_7783,N_7661,N_7690);
xnor U7784 (N_7784,N_7695,N_7517);
or U7785 (N_7785,N_7654,N_7674);
or U7786 (N_7786,N_7714,N_7500);
nor U7787 (N_7787,N_7504,N_7626);
nand U7788 (N_7788,N_7521,N_7593);
and U7789 (N_7789,N_7629,N_7739);
nor U7790 (N_7790,N_7598,N_7505);
xnor U7791 (N_7791,N_7697,N_7554);
and U7792 (N_7792,N_7568,N_7723);
xor U7793 (N_7793,N_7551,N_7733);
xor U7794 (N_7794,N_7599,N_7584);
nor U7795 (N_7795,N_7573,N_7673);
nand U7796 (N_7796,N_7567,N_7509);
nand U7797 (N_7797,N_7636,N_7681);
nand U7798 (N_7798,N_7607,N_7540);
or U7799 (N_7799,N_7622,N_7741);
xor U7800 (N_7800,N_7639,N_7534);
nand U7801 (N_7801,N_7550,N_7580);
and U7802 (N_7802,N_7510,N_7649);
nand U7803 (N_7803,N_7640,N_7662);
and U7804 (N_7804,N_7650,N_7678);
xnor U7805 (N_7805,N_7686,N_7575);
nand U7806 (N_7806,N_7672,N_7608);
and U7807 (N_7807,N_7563,N_7698);
nor U7808 (N_7808,N_7615,N_7694);
nand U7809 (N_7809,N_7528,N_7728);
nand U7810 (N_7810,N_7705,N_7735);
nor U7811 (N_7811,N_7713,N_7717);
or U7812 (N_7812,N_7623,N_7628);
nor U7813 (N_7813,N_7665,N_7744);
nor U7814 (N_7814,N_7601,N_7532);
or U7815 (N_7815,N_7547,N_7710);
xor U7816 (N_7816,N_7570,N_7561);
and U7817 (N_7817,N_7539,N_7715);
nand U7818 (N_7818,N_7543,N_7558);
xnor U7819 (N_7819,N_7519,N_7576);
and U7820 (N_7820,N_7560,N_7520);
nand U7821 (N_7821,N_7727,N_7651);
or U7822 (N_7822,N_7538,N_7587);
nor U7823 (N_7823,N_7600,N_7660);
nand U7824 (N_7824,N_7514,N_7515);
and U7825 (N_7825,N_7537,N_7726);
nor U7826 (N_7826,N_7704,N_7716);
nand U7827 (N_7827,N_7657,N_7648);
nand U7828 (N_7828,N_7609,N_7643);
xor U7829 (N_7829,N_7614,N_7602);
xnor U7830 (N_7830,N_7685,N_7591);
and U7831 (N_7831,N_7664,N_7738);
nand U7832 (N_7832,N_7522,N_7541);
or U7833 (N_7833,N_7667,N_7556);
xor U7834 (N_7834,N_7503,N_7574);
nor U7835 (N_7835,N_7518,N_7711);
nand U7836 (N_7836,N_7702,N_7740);
nor U7837 (N_7837,N_7652,N_7604);
nand U7838 (N_7838,N_7589,N_7524);
or U7839 (N_7839,N_7596,N_7683);
nor U7840 (N_7840,N_7616,N_7577);
and U7841 (N_7841,N_7687,N_7527);
xor U7842 (N_7842,N_7647,N_7653);
or U7843 (N_7843,N_7663,N_7513);
nand U7844 (N_7844,N_7611,N_7627);
or U7845 (N_7845,N_7669,N_7670);
or U7846 (N_7846,N_7564,N_7586);
nor U7847 (N_7847,N_7572,N_7562);
nand U7848 (N_7848,N_7624,N_7631);
or U7849 (N_7849,N_7745,N_7525);
xnor U7850 (N_7850,N_7633,N_7549);
xnor U7851 (N_7851,N_7749,N_7507);
nor U7852 (N_7852,N_7531,N_7724);
nand U7853 (N_7853,N_7523,N_7680);
nand U7854 (N_7854,N_7594,N_7571);
nand U7855 (N_7855,N_7688,N_7535);
and U7856 (N_7856,N_7644,N_7583);
nand U7857 (N_7857,N_7748,N_7732);
xnor U7858 (N_7858,N_7666,N_7566);
or U7859 (N_7859,N_7642,N_7722);
nor U7860 (N_7860,N_7565,N_7592);
nor U7861 (N_7861,N_7743,N_7516);
nor U7862 (N_7862,N_7553,N_7635);
nor U7863 (N_7863,N_7742,N_7625);
nor U7864 (N_7864,N_7630,N_7671);
nand U7865 (N_7865,N_7675,N_7595);
or U7866 (N_7866,N_7682,N_7659);
nand U7867 (N_7867,N_7719,N_7718);
nand U7868 (N_7868,N_7545,N_7511);
xor U7869 (N_7869,N_7641,N_7590);
xnor U7870 (N_7870,N_7646,N_7530);
xor U7871 (N_7871,N_7708,N_7529);
xor U7872 (N_7872,N_7746,N_7569);
xnor U7873 (N_7873,N_7725,N_7736);
xor U7874 (N_7874,N_7700,N_7603);
nor U7875 (N_7875,N_7716,N_7584);
and U7876 (N_7876,N_7587,N_7523);
nand U7877 (N_7877,N_7536,N_7711);
nor U7878 (N_7878,N_7544,N_7555);
and U7879 (N_7879,N_7526,N_7716);
nor U7880 (N_7880,N_7667,N_7742);
and U7881 (N_7881,N_7515,N_7573);
nand U7882 (N_7882,N_7716,N_7683);
xor U7883 (N_7883,N_7660,N_7632);
nor U7884 (N_7884,N_7520,N_7624);
xor U7885 (N_7885,N_7662,N_7637);
nor U7886 (N_7886,N_7540,N_7599);
nor U7887 (N_7887,N_7505,N_7679);
nor U7888 (N_7888,N_7729,N_7644);
nor U7889 (N_7889,N_7537,N_7632);
and U7890 (N_7890,N_7639,N_7673);
or U7891 (N_7891,N_7716,N_7736);
nand U7892 (N_7892,N_7728,N_7620);
nand U7893 (N_7893,N_7534,N_7717);
nand U7894 (N_7894,N_7671,N_7540);
nand U7895 (N_7895,N_7536,N_7522);
and U7896 (N_7896,N_7541,N_7658);
or U7897 (N_7897,N_7630,N_7583);
nand U7898 (N_7898,N_7636,N_7659);
nor U7899 (N_7899,N_7572,N_7728);
nor U7900 (N_7900,N_7615,N_7587);
or U7901 (N_7901,N_7542,N_7567);
nand U7902 (N_7902,N_7595,N_7565);
nand U7903 (N_7903,N_7643,N_7691);
nand U7904 (N_7904,N_7627,N_7723);
nor U7905 (N_7905,N_7574,N_7744);
and U7906 (N_7906,N_7500,N_7626);
xnor U7907 (N_7907,N_7556,N_7502);
and U7908 (N_7908,N_7746,N_7599);
or U7909 (N_7909,N_7681,N_7720);
and U7910 (N_7910,N_7614,N_7673);
nand U7911 (N_7911,N_7622,N_7684);
and U7912 (N_7912,N_7661,N_7534);
nand U7913 (N_7913,N_7634,N_7523);
or U7914 (N_7914,N_7529,N_7749);
xor U7915 (N_7915,N_7681,N_7605);
nand U7916 (N_7916,N_7552,N_7716);
xor U7917 (N_7917,N_7590,N_7642);
nand U7918 (N_7918,N_7543,N_7601);
nor U7919 (N_7919,N_7580,N_7661);
or U7920 (N_7920,N_7707,N_7554);
xor U7921 (N_7921,N_7747,N_7659);
nand U7922 (N_7922,N_7706,N_7595);
nand U7923 (N_7923,N_7581,N_7641);
or U7924 (N_7924,N_7568,N_7648);
or U7925 (N_7925,N_7659,N_7717);
xor U7926 (N_7926,N_7519,N_7659);
nand U7927 (N_7927,N_7544,N_7529);
nand U7928 (N_7928,N_7585,N_7595);
xor U7929 (N_7929,N_7526,N_7620);
nand U7930 (N_7930,N_7684,N_7563);
and U7931 (N_7931,N_7557,N_7722);
xnor U7932 (N_7932,N_7651,N_7631);
xor U7933 (N_7933,N_7696,N_7613);
nand U7934 (N_7934,N_7552,N_7715);
and U7935 (N_7935,N_7556,N_7576);
or U7936 (N_7936,N_7653,N_7592);
nand U7937 (N_7937,N_7683,N_7682);
and U7938 (N_7938,N_7711,N_7638);
xnor U7939 (N_7939,N_7694,N_7581);
nand U7940 (N_7940,N_7671,N_7529);
xnor U7941 (N_7941,N_7684,N_7646);
xor U7942 (N_7942,N_7709,N_7727);
and U7943 (N_7943,N_7539,N_7598);
or U7944 (N_7944,N_7621,N_7593);
and U7945 (N_7945,N_7735,N_7685);
nand U7946 (N_7946,N_7591,N_7505);
and U7947 (N_7947,N_7684,N_7636);
nor U7948 (N_7948,N_7620,N_7542);
or U7949 (N_7949,N_7736,N_7643);
or U7950 (N_7950,N_7603,N_7606);
and U7951 (N_7951,N_7681,N_7621);
and U7952 (N_7952,N_7626,N_7738);
nand U7953 (N_7953,N_7706,N_7620);
nor U7954 (N_7954,N_7648,N_7677);
or U7955 (N_7955,N_7712,N_7695);
nor U7956 (N_7956,N_7502,N_7529);
nand U7957 (N_7957,N_7710,N_7581);
nand U7958 (N_7958,N_7621,N_7690);
nand U7959 (N_7959,N_7664,N_7617);
xor U7960 (N_7960,N_7623,N_7647);
nor U7961 (N_7961,N_7515,N_7603);
nand U7962 (N_7962,N_7677,N_7703);
xor U7963 (N_7963,N_7589,N_7554);
xnor U7964 (N_7964,N_7545,N_7563);
nand U7965 (N_7965,N_7645,N_7504);
and U7966 (N_7966,N_7676,N_7566);
or U7967 (N_7967,N_7744,N_7708);
or U7968 (N_7968,N_7572,N_7506);
nand U7969 (N_7969,N_7727,N_7524);
nand U7970 (N_7970,N_7734,N_7703);
or U7971 (N_7971,N_7684,N_7654);
or U7972 (N_7972,N_7508,N_7637);
xor U7973 (N_7973,N_7723,N_7690);
or U7974 (N_7974,N_7711,N_7678);
nand U7975 (N_7975,N_7626,N_7677);
nor U7976 (N_7976,N_7565,N_7635);
and U7977 (N_7977,N_7700,N_7547);
and U7978 (N_7978,N_7535,N_7746);
or U7979 (N_7979,N_7597,N_7633);
nor U7980 (N_7980,N_7692,N_7512);
nor U7981 (N_7981,N_7711,N_7500);
xor U7982 (N_7982,N_7556,N_7564);
nor U7983 (N_7983,N_7647,N_7745);
and U7984 (N_7984,N_7603,N_7527);
and U7985 (N_7985,N_7529,N_7534);
and U7986 (N_7986,N_7562,N_7510);
xnor U7987 (N_7987,N_7651,N_7551);
and U7988 (N_7988,N_7593,N_7700);
or U7989 (N_7989,N_7653,N_7502);
xnor U7990 (N_7990,N_7542,N_7676);
nand U7991 (N_7991,N_7637,N_7501);
nor U7992 (N_7992,N_7606,N_7704);
nand U7993 (N_7993,N_7545,N_7556);
nor U7994 (N_7994,N_7719,N_7686);
xor U7995 (N_7995,N_7624,N_7633);
nor U7996 (N_7996,N_7624,N_7579);
nor U7997 (N_7997,N_7610,N_7652);
xnor U7998 (N_7998,N_7557,N_7727);
or U7999 (N_7999,N_7525,N_7563);
or U8000 (N_8000,N_7956,N_7966);
xor U8001 (N_8001,N_7981,N_7977);
and U8002 (N_8002,N_7826,N_7779);
nand U8003 (N_8003,N_7948,N_7907);
or U8004 (N_8004,N_7976,N_7855);
and U8005 (N_8005,N_7992,N_7880);
or U8006 (N_8006,N_7974,N_7849);
xor U8007 (N_8007,N_7886,N_7866);
and U8008 (N_8008,N_7854,N_7832);
and U8009 (N_8009,N_7877,N_7995);
nand U8010 (N_8010,N_7774,N_7908);
nor U8011 (N_8011,N_7798,N_7916);
nor U8012 (N_8012,N_7842,N_7949);
and U8013 (N_8013,N_7982,N_7864);
or U8014 (N_8014,N_7871,N_7758);
xor U8015 (N_8015,N_7996,N_7873);
nand U8016 (N_8016,N_7829,N_7891);
nor U8017 (N_8017,N_7904,N_7795);
and U8018 (N_8018,N_7923,N_7840);
xor U8019 (N_8019,N_7964,N_7994);
or U8020 (N_8020,N_7971,N_7884);
and U8021 (N_8021,N_7764,N_7847);
or U8022 (N_8022,N_7815,N_7984);
and U8023 (N_8023,N_7898,N_7761);
xnor U8024 (N_8024,N_7970,N_7801);
xnor U8025 (N_8025,N_7781,N_7818);
xor U8026 (N_8026,N_7934,N_7782);
xor U8027 (N_8027,N_7978,N_7867);
nand U8028 (N_8028,N_7786,N_7941);
nor U8029 (N_8029,N_7808,N_7835);
or U8030 (N_8030,N_7983,N_7915);
xor U8031 (N_8031,N_7980,N_7800);
and U8032 (N_8032,N_7892,N_7853);
nor U8033 (N_8033,N_7850,N_7828);
xnor U8034 (N_8034,N_7903,N_7888);
or U8035 (N_8035,N_7856,N_7794);
or U8036 (N_8036,N_7852,N_7767);
and U8037 (N_8037,N_7895,N_7857);
or U8038 (N_8038,N_7909,N_7804);
and U8039 (N_8039,N_7753,N_7940);
xnor U8040 (N_8040,N_7763,N_7851);
nand U8041 (N_8041,N_7897,N_7924);
or U8042 (N_8042,N_7929,N_7878);
xnor U8043 (N_8043,N_7845,N_7848);
and U8044 (N_8044,N_7822,N_7936);
nand U8045 (N_8045,N_7998,N_7975);
nand U8046 (N_8046,N_7811,N_7951);
nor U8047 (N_8047,N_7861,N_7947);
nand U8048 (N_8048,N_7963,N_7783);
or U8049 (N_8049,N_7799,N_7875);
and U8050 (N_8050,N_7931,N_7932);
xnor U8051 (N_8051,N_7942,N_7860);
or U8052 (N_8052,N_7921,N_7896);
or U8053 (N_8053,N_7912,N_7959);
nand U8054 (N_8054,N_7922,N_7760);
xor U8055 (N_8055,N_7913,N_7961);
or U8056 (N_8056,N_7930,N_7905);
nand U8057 (N_8057,N_7824,N_7838);
nand U8058 (N_8058,N_7890,N_7751);
xor U8059 (N_8059,N_7765,N_7759);
or U8060 (N_8060,N_7985,N_7846);
nand U8061 (N_8061,N_7754,N_7868);
or U8062 (N_8062,N_7991,N_7893);
and U8063 (N_8063,N_7986,N_7756);
xnor U8064 (N_8064,N_7881,N_7960);
and U8065 (N_8065,N_7920,N_7768);
and U8066 (N_8066,N_7870,N_7958);
nor U8067 (N_8067,N_7876,N_7973);
nand U8068 (N_8068,N_7772,N_7796);
nor U8069 (N_8069,N_7926,N_7967);
and U8070 (N_8070,N_7946,N_7938);
xor U8071 (N_8071,N_7831,N_7944);
and U8072 (N_8072,N_7787,N_7925);
xor U8073 (N_8073,N_7839,N_7836);
nand U8074 (N_8074,N_7843,N_7837);
nor U8075 (N_8075,N_7823,N_7919);
xor U8076 (N_8076,N_7957,N_7810);
nand U8077 (N_8077,N_7865,N_7834);
or U8078 (N_8078,N_7797,N_7972);
xor U8079 (N_8079,N_7937,N_7784);
nand U8080 (N_8080,N_7820,N_7894);
xnor U8081 (N_8081,N_7769,N_7803);
xor U8082 (N_8082,N_7918,N_7950);
xnor U8083 (N_8083,N_7819,N_7935);
or U8084 (N_8084,N_7841,N_7858);
nand U8085 (N_8085,N_7750,N_7790);
nand U8086 (N_8086,N_7954,N_7955);
and U8087 (N_8087,N_7993,N_7805);
xnor U8088 (N_8088,N_7862,N_7816);
or U8089 (N_8089,N_7806,N_7989);
and U8090 (N_8090,N_7785,N_7882);
or U8091 (N_8091,N_7863,N_7833);
nor U8092 (N_8092,N_7757,N_7911);
nand U8093 (N_8093,N_7945,N_7809);
xor U8094 (N_8094,N_7997,N_7817);
nand U8095 (N_8095,N_7889,N_7988);
nor U8096 (N_8096,N_7825,N_7821);
and U8097 (N_8097,N_7899,N_7969);
nand U8098 (N_8098,N_7939,N_7778);
nor U8099 (N_8099,N_7777,N_7812);
xnor U8100 (N_8100,N_7859,N_7814);
or U8101 (N_8101,N_7844,N_7900);
or U8102 (N_8102,N_7830,N_7914);
nor U8103 (N_8103,N_7766,N_7792);
nor U8104 (N_8104,N_7791,N_7965);
or U8105 (N_8105,N_7902,N_7901);
nor U8106 (N_8106,N_7990,N_7780);
xor U8107 (N_8107,N_7887,N_7879);
and U8108 (N_8108,N_7762,N_7793);
or U8109 (N_8109,N_7987,N_7979);
nor U8110 (N_8110,N_7910,N_7807);
and U8111 (N_8111,N_7999,N_7827);
xnor U8112 (N_8112,N_7968,N_7789);
nand U8113 (N_8113,N_7885,N_7813);
xor U8114 (N_8114,N_7775,N_7872);
and U8115 (N_8115,N_7928,N_7927);
or U8116 (N_8116,N_7952,N_7802);
nor U8117 (N_8117,N_7874,N_7943);
or U8118 (N_8118,N_7953,N_7906);
or U8119 (N_8119,N_7771,N_7883);
nor U8120 (N_8120,N_7773,N_7962);
xnor U8121 (N_8121,N_7776,N_7933);
xnor U8122 (N_8122,N_7755,N_7752);
or U8123 (N_8123,N_7770,N_7869);
xor U8124 (N_8124,N_7917,N_7788);
xnor U8125 (N_8125,N_7880,N_7919);
or U8126 (N_8126,N_7981,N_7952);
nor U8127 (N_8127,N_7776,N_7785);
and U8128 (N_8128,N_7889,N_7805);
and U8129 (N_8129,N_7785,N_7887);
nand U8130 (N_8130,N_7797,N_7813);
nand U8131 (N_8131,N_7807,N_7870);
or U8132 (N_8132,N_7922,N_7890);
and U8133 (N_8133,N_7847,N_7790);
nand U8134 (N_8134,N_7753,N_7788);
or U8135 (N_8135,N_7918,N_7845);
xnor U8136 (N_8136,N_7923,N_7962);
and U8137 (N_8137,N_7768,N_7872);
and U8138 (N_8138,N_7832,N_7907);
or U8139 (N_8139,N_7768,N_7854);
xor U8140 (N_8140,N_7816,N_7797);
nand U8141 (N_8141,N_7820,N_7807);
nor U8142 (N_8142,N_7939,N_7985);
and U8143 (N_8143,N_7922,N_7757);
and U8144 (N_8144,N_7895,N_7825);
nor U8145 (N_8145,N_7765,N_7789);
or U8146 (N_8146,N_7874,N_7857);
xnor U8147 (N_8147,N_7932,N_7997);
nor U8148 (N_8148,N_7907,N_7855);
nand U8149 (N_8149,N_7967,N_7755);
xnor U8150 (N_8150,N_7871,N_7953);
xnor U8151 (N_8151,N_7806,N_7925);
and U8152 (N_8152,N_7788,N_7975);
or U8153 (N_8153,N_7915,N_7989);
nor U8154 (N_8154,N_7961,N_7847);
or U8155 (N_8155,N_7918,N_7837);
xor U8156 (N_8156,N_7899,N_7876);
xnor U8157 (N_8157,N_7910,N_7975);
or U8158 (N_8158,N_7981,N_7961);
nor U8159 (N_8159,N_7997,N_7919);
nor U8160 (N_8160,N_7854,N_7866);
and U8161 (N_8161,N_7869,N_7777);
and U8162 (N_8162,N_7915,N_7804);
or U8163 (N_8163,N_7827,N_7959);
nand U8164 (N_8164,N_7914,N_7981);
and U8165 (N_8165,N_7796,N_7941);
or U8166 (N_8166,N_7937,N_7966);
xnor U8167 (N_8167,N_7965,N_7793);
and U8168 (N_8168,N_7838,N_7901);
or U8169 (N_8169,N_7807,N_7947);
or U8170 (N_8170,N_7964,N_7773);
nand U8171 (N_8171,N_7815,N_7885);
or U8172 (N_8172,N_7847,N_7976);
nor U8173 (N_8173,N_7998,N_7997);
nand U8174 (N_8174,N_7960,N_7775);
nand U8175 (N_8175,N_7878,N_7804);
xor U8176 (N_8176,N_7980,N_7993);
or U8177 (N_8177,N_7916,N_7790);
nand U8178 (N_8178,N_7819,N_7809);
and U8179 (N_8179,N_7860,N_7846);
or U8180 (N_8180,N_7979,N_7783);
xor U8181 (N_8181,N_7823,N_7953);
nand U8182 (N_8182,N_7810,N_7764);
and U8183 (N_8183,N_7753,N_7998);
xor U8184 (N_8184,N_7920,N_7759);
or U8185 (N_8185,N_7933,N_7858);
or U8186 (N_8186,N_7760,N_7960);
or U8187 (N_8187,N_7992,N_7984);
xor U8188 (N_8188,N_7984,N_7994);
nor U8189 (N_8189,N_7788,N_7835);
xor U8190 (N_8190,N_7961,N_7880);
nand U8191 (N_8191,N_7755,N_7902);
xnor U8192 (N_8192,N_7855,N_7755);
nor U8193 (N_8193,N_7923,N_7883);
or U8194 (N_8194,N_7932,N_7911);
and U8195 (N_8195,N_7886,N_7770);
and U8196 (N_8196,N_7885,N_7867);
nand U8197 (N_8197,N_7928,N_7848);
xnor U8198 (N_8198,N_7959,N_7819);
or U8199 (N_8199,N_7853,N_7880);
or U8200 (N_8200,N_7958,N_7764);
and U8201 (N_8201,N_7822,N_7947);
or U8202 (N_8202,N_7753,N_7924);
xnor U8203 (N_8203,N_7934,N_7767);
xnor U8204 (N_8204,N_7897,N_7757);
and U8205 (N_8205,N_7812,N_7936);
or U8206 (N_8206,N_7763,N_7819);
xor U8207 (N_8207,N_7881,N_7766);
xnor U8208 (N_8208,N_7816,N_7938);
xnor U8209 (N_8209,N_7995,N_7895);
nand U8210 (N_8210,N_7893,N_7964);
nor U8211 (N_8211,N_7947,N_7873);
xor U8212 (N_8212,N_7996,N_7750);
nand U8213 (N_8213,N_7979,N_7871);
nand U8214 (N_8214,N_7975,N_7908);
nor U8215 (N_8215,N_7806,N_7812);
nor U8216 (N_8216,N_7933,N_7847);
nand U8217 (N_8217,N_7880,N_7889);
or U8218 (N_8218,N_7982,N_7761);
and U8219 (N_8219,N_7849,N_7834);
nand U8220 (N_8220,N_7825,N_7832);
nor U8221 (N_8221,N_7901,N_7819);
nand U8222 (N_8222,N_7885,N_7958);
xnor U8223 (N_8223,N_7983,N_7899);
nor U8224 (N_8224,N_7944,N_7971);
xnor U8225 (N_8225,N_7920,N_7927);
and U8226 (N_8226,N_7864,N_7971);
nand U8227 (N_8227,N_7924,N_7888);
nand U8228 (N_8228,N_7857,N_7796);
and U8229 (N_8229,N_7785,N_7884);
and U8230 (N_8230,N_7828,N_7825);
nor U8231 (N_8231,N_7772,N_7756);
and U8232 (N_8232,N_7863,N_7921);
or U8233 (N_8233,N_7830,N_7772);
xor U8234 (N_8234,N_7753,N_7976);
nand U8235 (N_8235,N_7947,N_7998);
nand U8236 (N_8236,N_7830,N_7906);
and U8237 (N_8237,N_7927,N_7806);
xor U8238 (N_8238,N_7965,N_7933);
nor U8239 (N_8239,N_7984,N_7927);
and U8240 (N_8240,N_7801,N_7799);
and U8241 (N_8241,N_7876,N_7993);
and U8242 (N_8242,N_7826,N_7889);
or U8243 (N_8243,N_7972,N_7941);
and U8244 (N_8244,N_7901,N_7761);
xor U8245 (N_8245,N_7992,N_7923);
or U8246 (N_8246,N_7914,N_7911);
nor U8247 (N_8247,N_7841,N_7781);
nor U8248 (N_8248,N_7984,N_7908);
nand U8249 (N_8249,N_7871,N_7996);
xnor U8250 (N_8250,N_8094,N_8160);
xnor U8251 (N_8251,N_8027,N_8048);
and U8252 (N_8252,N_8185,N_8221);
and U8253 (N_8253,N_8034,N_8181);
nor U8254 (N_8254,N_8202,N_8071);
xor U8255 (N_8255,N_8206,N_8172);
and U8256 (N_8256,N_8062,N_8211);
nor U8257 (N_8257,N_8067,N_8164);
nor U8258 (N_8258,N_8014,N_8168);
xnor U8259 (N_8259,N_8163,N_8115);
xnor U8260 (N_8260,N_8131,N_8196);
nor U8261 (N_8261,N_8158,N_8199);
or U8262 (N_8262,N_8037,N_8056);
or U8263 (N_8263,N_8015,N_8002);
xor U8264 (N_8264,N_8183,N_8189);
nand U8265 (N_8265,N_8084,N_8234);
nor U8266 (N_8266,N_8069,N_8197);
nor U8267 (N_8267,N_8139,N_8247);
xor U8268 (N_8268,N_8046,N_8138);
xor U8269 (N_8269,N_8016,N_8060);
or U8270 (N_8270,N_8008,N_8063);
and U8271 (N_8271,N_8021,N_8153);
nand U8272 (N_8272,N_8082,N_8175);
xor U8273 (N_8273,N_8177,N_8148);
and U8274 (N_8274,N_8194,N_8118);
xnor U8275 (N_8275,N_8147,N_8210);
nor U8276 (N_8276,N_8242,N_8188);
xnor U8277 (N_8277,N_8077,N_8036);
nand U8278 (N_8278,N_8180,N_8142);
or U8279 (N_8279,N_8201,N_8162);
xor U8280 (N_8280,N_8150,N_8228);
or U8281 (N_8281,N_8100,N_8165);
nor U8282 (N_8282,N_8054,N_8076);
or U8283 (N_8283,N_8203,N_8184);
nor U8284 (N_8284,N_8246,N_8081);
nor U8285 (N_8285,N_8132,N_8135);
nor U8286 (N_8286,N_8151,N_8116);
xor U8287 (N_8287,N_8025,N_8230);
or U8288 (N_8288,N_8146,N_8149);
xor U8289 (N_8289,N_8134,N_8239);
nor U8290 (N_8290,N_8011,N_8238);
nor U8291 (N_8291,N_8170,N_8220);
nor U8292 (N_8292,N_8186,N_8087);
or U8293 (N_8293,N_8190,N_8061);
and U8294 (N_8294,N_8130,N_8001);
and U8295 (N_8295,N_8078,N_8167);
xnor U8296 (N_8296,N_8022,N_8026);
and U8297 (N_8297,N_8166,N_8227);
nor U8298 (N_8298,N_8216,N_8092);
nand U8299 (N_8299,N_8217,N_8129);
nor U8300 (N_8300,N_8058,N_8065);
nor U8301 (N_8301,N_8088,N_8178);
or U8302 (N_8302,N_8013,N_8137);
or U8303 (N_8303,N_8161,N_8109);
xor U8304 (N_8304,N_8004,N_8053);
nand U8305 (N_8305,N_8140,N_8112);
nor U8306 (N_8306,N_8072,N_8233);
nand U8307 (N_8307,N_8101,N_8017);
and U8308 (N_8308,N_8083,N_8113);
nor U8309 (N_8309,N_8219,N_8085);
or U8310 (N_8310,N_8191,N_8057);
nand U8311 (N_8311,N_8079,N_8218);
nand U8312 (N_8312,N_8075,N_8245);
and U8313 (N_8313,N_8144,N_8103);
and U8314 (N_8314,N_8223,N_8179);
and U8315 (N_8315,N_8225,N_8173);
nor U8316 (N_8316,N_8068,N_8044);
and U8317 (N_8317,N_8120,N_8157);
xor U8318 (N_8318,N_8169,N_8136);
nor U8319 (N_8319,N_8143,N_8198);
xnor U8320 (N_8320,N_8003,N_8192);
nor U8321 (N_8321,N_8000,N_8106);
nor U8322 (N_8322,N_8102,N_8123);
or U8323 (N_8323,N_8032,N_8193);
or U8324 (N_8324,N_8038,N_8125);
xnor U8325 (N_8325,N_8126,N_8237);
nor U8326 (N_8326,N_8099,N_8041);
nand U8327 (N_8327,N_8195,N_8096);
or U8328 (N_8328,N_8205,N_8119);
nor U8329 (N_8329,N_8128,N_8171);
or U8330 (N_8330,N_8204,N_8122);
and U8331 (N_8331,N_8007,N_8222);
nor U8332 (N_8332,N_8009,N_8226);
and U8333 (N_8333,N_8033,N_8066);
xor U8334 (N_8334,N_8070,N_8110);
nor U8335 (N_8335,N_8097,N_8224);
or U8336 (N_8336,N_8111,N_8093);
nor U8337 (N_8337,N_8209,N_8050);
or U8338 (N_8338,N_8154,N_8124);
nand U8339 (N_8339,N_8064,N_8145);
nand U8340 (N_8340,N_8086,N_8024);
xnor U8341 (N_8341,N_8010,N_8019);
or U8342 (N_8342,N_8020,N_8091);
and U8343 (N_8343,N_8040,N_8187);
xor U8344 (N_8344,N_8107,N_8030);
and U8345 (N_8345,N_8090,N_8244);
xnor U8346 (N_8346,N_8074,N_8127);
or U8347 (N_8347,N_8028,N_8049);
nand U8348 (N_8348,N_8200,N_8214);
or U8349 (N_8349,N_8159,N_8240);
or U8350 (N_8350,N_8243,N_8039);
nor U8351 (N_8351,N_8117,N_8005);
nor U8352 (N_8352,N_8182,N_8012);
nand U8353 (N_8353,N_8241,N_8047);
xnor U8354 (N_8354,N_8105,N_8059);
or U8355 (N_8355,N_8035,N_8029);
nand U8356 (N_8356,N_8235,N_8006);
xnor U8357 (N_8357,N_8018,N_8098);
nor U8358 (N_8358,N_8133,N_8045);
xnor U8359 (N_8359,N_8207,N_8073);
nor U8360 (N_8360,N_8232,N_8248);
and U8361 (N_8361,N_8104,N_8141);
nand U8362 (N_8362,N_8215,N_8152);
xnor U8363 (N_8363,N_8042,N_8155);
nand U8364 (N_8364,N_8208,N_8212);
xor U8365 (N_8365,N_8052,N_8080);
nor U8366 (N_8366,N_8236,N_8121);
nor U8367 (N_8367,N_8023,N_8108);
or U8368 (N_8368,N_8095,N_8055);
nor U8369 (N_8369,N_8249,N_8051);
nand U8370 (N_8370,N_8043,N_8089);
nand U8371 (N_8371,N_8031,N_8176);
and U8372 (N_8372,N_8213,N_8231);
nor U8373 (N_8373,N_8174,N_8114);
nor U8374 (N_8374,N_8229,N_8156);
or U8375 (N_8375,N_8022,N_8127);
nand U8376 (N_8376,N_8140,N_8234);
or U8377 (N_8377,N_8100,N_8159);
nand U8378 (N_8378,N_8239,N_8107);
xor U8379 (N_8379,N_8204,N_8020);
nor U8380 (N_8380,N_8087,N_8153);
nand U8381 (N_8381,N_8153,N_8024);
nor U8382 (N_8382,N_8053,N_8133);
xnor U8383 (N_8383,N_8231,N_8187);
nand U8384 (N_8384,N_8167,N_8031);
nand U8385 (N_8385,N_8055,N_8067);
xnor U8386 (N_8386,N_8074,N_8209);
and U8387 (N_8387,N_8203,N_8089);
nand U8388 (N_8388,N_8158,N_8001);
or U8389 (N_8389,N_8230,N_8136);
nor U8390 (N_8390,N_8084,N_8175);
xnor U8391 (N_8391,N_8168,N_8203);
nor U8392 (N_8392,N_8060,N_8008);
nand U8393 (N_8393,N_8033,N_8098);
xor U8394 (N_8394,N_8096,N_8103);
nand U8395 (N_8395,N_8024,N_8234);
or U8396 (N_8396,N_8153,N_8106);
and U8397 (N_8397,N_8085,N_8099);
nor U8398 (N_8398,N_8114,N_8108);
or U8399 (N_8399,N_8233,N_8179);
or U8400 (N_8400,N_8207,N_8008);
or U8401 (N_8401,N_8226,N_8135);
nor U8402 (N_8402,N_8023,N_8204);
nand U8403 (N_8403,N_8066,N_8106);
xor U8404 (N_8404,N_8248,N_8195);
nor U8405 (N_8405,N_8115,N_8248);
xor U8406 (N_8406,N_8097,N_8173);
xor U8407 (N_8407,N_8011,N_8097);
nand U8408 (N_8408,N_8004,N_8019);
nand U8409 (N_8409,N_8017,N_8181);
nand U8410 (N_8410,N_8054,N_8068);
and U8411 (N_8411,N_8156,N_8108);
and U8412 (N_8412,N_8021,N_8159);
nor U8413 (N_8413,N_8035,N_8197);
xnor U8414 (N_8414,N_8149,N_8170);
nor U8415 (N_8415,N_8080,N_8158);
and U8416 (N_8416,N_8215,N_8009);
or U8417 (N_8417,N_8098,N_8236);
nand U8418 (N_8418,N_8136,N_8149);
and U8419 (N_8419,N_8067,N_8030);
or U8420 (N_8420,N_8093,N_8164);
nor U8421 (N_8421,N_8172,N_8029);
nor U8422 (N_8422,N_8115,N_8249);
nand U8423 (N_8423,N_8217,N_8061);
xnor U8424 (N_8424,N_8066,N_8005);
and U8425 (N_8425,N_8118,N_8196);
nand U8426 (N_8426,N_8170,N_8049);
xor U8427 (N_8427,N_8223,N_8021);
nor U8428 (N_8428,N_8247,N_8088);
nor U8429 (N_8429,N_8032,N_8067);
nand U8430 (N_8430,N_8227,N_8187);
nor U8431 (N_8431,N_8011,N_8102);
nor U8432 (N_8432,N_8136,N_8140);
xor U8433 (N_8433,N_8217,N_8062);
or U8434 (N_8434,N_8111,N_8240);
or U8435 (N_8435,N_8180,N_8053);
nand U8436 (N_8436,N_8037,N_8244);
nand U8437 (N_8437,N_8172,N_8101);
nand U8438 (N_8438,N_8119,N_8133);
and U8439 (N_8439,N_8192,N_8221);
nand U8440 (N_8440,N_8205,N_8068);
and U8441 (N_8441,N_8033,N_8021);
xor U8442 (N_8442,N_8018,N_8221);
xor U8443 (N_8443,N_8024,N_8128);
nor U8444 (N_8444,N_8221,N_8146);
xnor U8445 (N_8445,N_8071,N_8049);
nor U8446 (N_8446,N_8198,N_8166);
xnor U8447 (N_8447,N_8189,N_8003);
nor U8448 (N_8448,N_8108,N_8196);
nand U8449 (N_8449,N_8178,N_8103);
and U8450 (N_8450,N_8213,N_8188);
nor U8451 (N_8451,N_8006,N_8079);
or U8452 (N_8452,N_8051,N_8127);
nand U8453 (N_8453,N_8061,N_8100);
or U8454 (N_8454,N_8184,N_8098);
nand U8455 (N_8455,N_8064,N_8246);
nand U8456 (N_8456,N_8100,N_8147);
or U8457 (N_8457,N_8127,N_8134);
nor U8458 (N_8458,N_8212,N_8249);
and U8459 (N_8459,N_8014,N_8097);
and U8460 (N_8460,N_8011,N_8075);
or U8461 (N_8461,N_8001,N_8152);
and U8462 (N_8462,N_8150,N_8134);
nand U8463 (N_8463,N_8096,N_8203);
and U8464 (N_8464,N_8068,N_8071);
nor U8465 (N_8465,N_8093,N_8114);
or U8466 (N_8466,N_8091,N_8058);
nand U8467 (N_8467,N_8119,N_8003);
xnor U8468 (N_8468,N_8188,N_8153);
or U8469 (N_8469,N_8055,N_8103);
or U8470 (N_8470,N_8223,N_8202);
and U8471 (N_8471,N_8051,N_8043);
or U8472 (N_8472,N_8055,N_8072);
nand U8473 (N_8473,N_8222,N_8155);
and U8474 (N_8474,N_8104,N_8190);
nand U8475 (N_8475,N_8048,N_8085);
nand U8476 (N_8476,N_8035,N_8170);
nand U8477 (N_8477,N_8093,N_8155);
nor U8478 (N_8478,N_8079,N_8071);
and U8479 (N_8479,N_8160,N_8065);
nor U8480 (N_8480,N_8050,N_8214);
and U8481 (N_8481,N_8009,N_8181);
and U8482 (N_8482,N_8167,N_8058);
nand U8483 (N_8483,N_8082,N_8167);
and U8484 (N_8484,N_8078,N_8071);
xnor U8485 (N_8485,N_8074,N_8227);
and U8486 (N_8486,N_8019,N_8198);
nand U8487 (N_8487,N_8120,N_8241);
nand U8488 (N_8488,N_8176,N_8014);
xnor U8489 (N_8489,N_8103,N_8188);
or U8490 (N_8490,N_8033,N_8163);
xnor U8491 (N_8491,N_8119,N_8149);
nor U8492 (N_8492,N_8136,N_8177);
and U8493 (N_8493,N_8181,N_8058);
nor U8494 (N_8494,N_8102,N_8087);
xnor U8495 (N_8495,N_8214,N_8117);
nand U8496 (N_8496,N_8059,N_8081);
or U8497 (N_8497,N_8246,N_8213);
xnor U8498 (N_8498,N_8107,N_8025);
or U8499 (N_8499,N_8163,N_8030);
nand U8500 (N_8500,N_8273,N_8349);
nor U8501 (N_8501,N_8301,N_8348);
nand U8502 (N_8502,N_8253,N_8486);
nor U8503 (N_8503,N_8326,N_8436);
and U8504 (N_8504,N_8464,N_8435);
nand U8505 (N_8505,N_8399,N_8261);
nor U8506 (N_8506,N_8434,N_8375);
nand U8507 (N_8507,N_8354,N_8458);
or U8508 (N_8508,N_8438,N_8479);
xor U8509 (N_8509,N_8318,N_8363);
or U8510 (N_8510,N_8310,N_8328);
nand U8511 (N_8511,N_8267,N_8400);
xor U8512 (N_8512,N_8335,N_8333);
nand U8513 (N_8513,N_8358,N_8446);
nor U8514 (N_8514,N_8304,N_8415);
or U8515 (N_8515,N_8497,N_8362);
nor U8516 (N_8516,N_8456,N_8380);
xor U8517 (N_8517,N_8414,N_8483);
xnor U8518 (N_8518,N_8347,N_8432);
nor U8519 (N_8519,N_8441,N_8272);
and U8520 (N_8520,N_8403,N_8313);
nand U8521 (N_8521,N_8448,N_8296);
nand U8522 (N_8522,N_8384,N_8379);
xnor U8523 (N_8523,N_8480,N_8365);
nor U8524 (N_8524,N_8281,N_8444);
and U8525 (N_8525,N_8445,N_8492);
nor U8526 (N_8526,N_8440,N_8406);
xnor U8527 (N_8527,N_8329,N_8312);
nor U8528 (N_8528,N_8316,N_8332);
and U8529 (N_8529,N_8300,N_8423);
nor U8530 (N_8530,N_8256,N_8370);
and U8531 (N_8531,N_8334,N_8465);
and U8532 (N_8532,N_8376,N_8342);
nor U8533 (N_8533,N_8346,N_8339);
nand U8534 (N_8534,N_8289,N_8297);
nor U8535 (N_8535,N_8343,N_8258);
nor U8536 (N_8536,N_8484,N_8449);
nor U8537 (N_8537,N_8425,N_8459);
xor U8538 (N_8538,N_8321,N_8340);
or U8539 (N_8539,N_8412,N_8386);
nor U8540 (N_8540,N_8292,N_8433);
nor U8541 (N_8541,N_8345,N_8426);
xor U8542 (N_8542,N_8481,N_8282);
nor U8543 (N_8543,N_8407,N_8271);
nor U8544 (N_8544,N_8311,N_8262);
nor U8545 (N_8545,N_8265,N_8417);
and U8546 (N_8546,N_8420,N_8495);
nor U8547 (N_8547,N_8361,N_8372);
and U8548 (N_8548,N_8302,N_8392);
and U8549 (N_8549,N_8390,N_8350);
nand U8550 (N_8550,N_8467,N_8295);
and U8551 (N_8551,N_8298,N_8266);
and U8552 (N_8552,N_8330,N_8315);
or U8553 (N_8553,N_8257,N_8286);
or U8554 (N_8554,N_8462,N_8453);
xnor U8555 (N_8555,N_8478,N_8381);
xor U8556 (N_8556,N_8367,N_8290);
and U8557 (N_8557,N_8250,N_8359);
xor U8558 (N_8558,N_8491,N_8439);
or U8559 (N_8559,N_8357,N_8387);
and U8560 (N_8560,N_8306,N_8396);
xnor U8561 (N_8561,N_8393,N_8490);
or U8562 (N_8562,N_8398,N_8450);
nor U8563 (N_8563,N_8410,N_8285);
or U8564 (N_8564,N_8428,N_8424);
and U8565 (N_8565,N_8251,N_8344);
and U8566 (N_8566,N_8309,N_8274);
or U8567 (N_8567,N_8499,N_8377);
xor U8568 (N_8568,N_8442,N_8320);
or U8569 (N_8569,N_8451,N_8287);
nand U8570 (N_8570,N_8457,N_8408);
xor U8571 (N_8571,N_8443,N_8284);
xnor U8572 (N_8572,N_8371,N_8356);
xor U8573 (N_8573,N_8402,N_8264);
or U8574 (N_8574,N_8404,N_8317);
and U8575 (N_8575,N_8291,N_8416);
xnor U8576 (N_8576,N_8489,N_8259);
nand U8577 (N_8577,N_8391,N_8485);
nand U8578 (N_8578,N_8283,N_8314);
or U8579 (N_8579,N_8252,N_8418);
and U8580 (N_8580,N_8482,N_8382);
or U8581 (N_8581,N_8411,N_8324);
or U8582 (N_8582,N_8496,N_8385);
nor U8583 (N_8583,N_8260,N_8364);
xnor U8584 (N_8584,N_8394,N_8460);
nor U8585 (N_8585,N_8255,N_8331);
or U8586 (N_8586,N_8336,N_8427);
and U8587 (N_8587,N_8498,N_8461);
xnor U8588 (N_8588,N_8337,N_8294);
or U8589 (N_8589,N_8308,N_8463);
or U8590 (N_8590,N_8299,N_8338);
or U8591 (N_8591,N_8369,N_8254);
or U8592 (N_8592,N_8405,N_8351);
nand U8593 (N_8593,N_8319,N_8341);
and U8594 (N_8594,N_8378,N_8327);
or U8595 (N_8595,N_8323,N_8383);
and U8596 (N_8596,N_8474,N_8360);
or U8597 (N_8597,N_8388,N_8275);
and U8598 (N_8598,N_8468,N_8279);
nand U8599 (N_8599,N_8303,N_8488);
nor U8600 (N_8600,N_8473,N_8397);
nor U8601 (N_8601,N_8419,N_8475);
or U8602 (N_8602,N_8494,N_8413);
or U8603 (N_8603,N_8263,N_8452);
nand U8604 (N_8604,N_8374,N_8447);
and U8605 (N_8605,N_8430,N_8278);
and U8606 (N_8606,N_8322,N_8325);
nand U8607 (N_8607,N_8401,N_8395);
nand U8608 (N_8608,N_8422,N_8389);
and U8609 (N_8609,N_8437,N_8276);
nor U8610 (N_8610,N_8429,N_8280);
nor U8611 (N_8611,N_8305,N_8270);
xnor U8612 (N_8612,N_8366,N_8269);
and U8613 (N_8613,N_8421,N_8493);
nand U8614 (N_8614,N_8288,N_8487);
or U8615 (N_8615,N_8409,N_8307);
or U8616 (N_8616,N_8431,N_8277);
xnor U8617 (N_8617,N_8455,N_8470);
xor U8618 (N_8618,N_8477,N_8352);
or U8619 (N_8619,N_8454,N_8472);
and U8620 (N_8620,N_8268,N_8355);
xor U8621 (N_8621,N_8466,N_8373);
nand U8622 (N_8622,N_8469,N_8476);
xnor U8623 (N_8623,N_8353,N_8368);
nand U8624 (N_8624,N_8471,N_8293);
nand U8625 (N_8625,N_8345,N_8316);
or U8626 (N_8626,N_8472,N_8379);
nand U8627 (N_8627,N_8496,N_8392);
nand U8628 (N_8628,N_8277,N_8335);
or U8629 (N_8629,N_8287,N_8349);
nor U8630 (N_8630,N_8462,N_8364);
nand U8631 (N_8631,N_8458,N_8408);
nor U8632 (N_8632,N_8474,N_8317);
xor U8633 (N_8633,N_8460,N_8412);
and U8634 (N_8634,N_8474,N_8274);
nand U8635 (N_8635,N_8462,N_8383);
or U8636 (N_8636,N_8319,N_8345);
nand U8637 (N_8637,N_8400,N_8375);
xor U8638 (N_8638,N_8462,N_8399);
nor U8639 (N_8639,N_8302,N_8257);
and U8640 (N_8640,N_8374,N_8475);
nand U8641 (N_8641,N_8470,N_8449);
xor U8642 (N_8642,N_8362,N_8296);
or U8643 (N_8643,N_8384,N_8436);
nor U8644 (N_8644,N_8284,N_8410);
nand U8645 (N_8645,N_8450,N_8432);
nand U8646 (N_8646,N_8497,N_8356);
xnor U8647 (N_8647,N_8306,N_8496);
nor U8648 (N_8648,N_8351,N_8319);
xor U8649 (N_8649,N_8377,N_8304);
nand U8650 (N_8650,N_8473,N_8482);
xnor U8651 (N_8651,N_8482,N_8317);
or U8652 (N_8652,N_8291,N_8488);
nor U8653 (N_8653,N_8283,N_8488);
xnor U8654 (N_8654,N_8316,N_8405);
and U8655 (N_8655,N_8298,N_8462);
nor U8656 (N_8656,N_8282,N_8492);
xnor U8657 (N_8657,N_8270,N_8418);
and U8658 (N_8658,N_8274,N_8294);
nor U8659 (N_8659,N_8347,N_8391);
and U8660 (N_8660,N_8457,N_8305);
or U8661 (N_8661,N_8446,N_8330);
or U8662 (N_8662,N_8446,N_8322);
nor U8663 (N_8663,N_8301,N_8419);
and U8664 (N_8664,N_8433,N_8430);
nor U8665 (N_8665,N_8308,N_8348);
nor U8666 (N_8666,N_8258,N_8362);
or U8667 (N_8667,N_8301,N_8291);
nor U8668 (N_8668,N_8257,N_8320);
and U8669 (N_8669,N_8395,N_8468);
and U8670 (N_8670,N_8330,N_8269);
and U8671 (N_8671,N_8385,N_8493);
and U8672 (N_8672,N_8303,N_8366);
xor U8673 (N_8673,N_8453,N_8313);
or U8674 (N_8674,N_8387,N_8301);
nor U8675 (N_8675,N_8411,N_8414);
xnor U8676 (N_8676,N_8289,N_8480);
and U8677 (N_8677,N_8496,N_8336);
and U8678 (N_8678,N_8336,N_8468);
or U8679 (N_8679,N_8323,N_8250);
and U8680 (N_8680,N_8479,N_8357);
or U8681 (N_8681,N_8259,N_8314);
or U8682 (N_8682,N_8468,N_8453);
and U8683 (N_8683,N_8492,N_8252);
or U8684 (N_8684,N_8336,N_8410);
xnor U8685 (N_8685,N_8339,N_8447);
nor U8686 (N_8686,N_8444,N_8490);
nor U8687 (N_8687,N_8399,N_8335);
xor U8688 (N_8688,N_8436,N_8250);
or U8689 (N_8689,N_8333,N_8478);
and U8690 (N_8690,N_8429,N_8277);
nand U8691 (N_8691,N_8398,N_8421);
and U8692 (N_8692,N_8459,N_8429);
nand U8693 (N_8693,N_8369,N_8430);
or U8694 (N_8694,N_8380,N_8462);
nor U8695 (N_8695,N_8406,N_8382);
nor U8696 (N_8696,N_8261,N_8328);
and U8697 (N_8697,N_8317,N_8435);
or U8698 (N_8698,N_8399,N_8345);
and U8699 (N_8699,N_8441,N_8490);
and U8700 (N_8700,N_8379,N_8407);
nor U8701 (N_8701,N_8412,N_8497);
xor U8702 (N_8702,N_8418,N_8341);
nor U8703 (N_8703,N_8403,N_8472);
and U8704 (N_8704,N_8392,N_8420);
and U8705 (N_8705,N_8326,N_8309);
nand U8706 (N_8706,N_8340,N_8437);
xnor U8707 (N_8707,N_8472,N_8363);
xnor U8708 (N_8708,N_8326,N_8355);
nor U8709 (N_8709,N_8445,N_8420);
xnor U8710 (N_8710,N_8373,N_8465);
and U8711 (N_8711,N_8257,N_8293);
and U8712 (N_8712,N_8435,N_8301);
or U8713 (N_8713,N_8299,N_8460);
or U8714 (N_8714,N_8357,N_8256);
and U8715 (N_8715,N_8449,N_8307);
or U8716 (N_8716,N_8475,N_8493);
nor U8717 (N_8717,N_8348,N_8312);
xor U8718 (N_8718,N_8255,N_8355);
nor U8719 (N_8719,N_8454,N_8345);
nor U8720 (N_8720,N_8472,N_8396);
and U8721 (N_8721,N_8416,N_8410);
and U8722 (N_8722,N_8497,N_8329);
and U8723 (N_8723,N_8356,N_8393);
xor U8724 (N_8724,N_8336,N_8302);
nor U8725 (N_8725,N_8376,N_8367);
nor U8726 (N_8726,N_8258,N_8422);
and U8727 (N_8727,N_8416,N_8253);
nor U8728 (N_8728,N_8317,N_8258);
and U8729 (N_8729,N_8250,N_8281);
xor U8730 (N_8730,N_8375,N_8432);
nor U8731 (N_8731,N_8445,N_8403);
or U8732 (N_8732,N_8328,N_8357);
xnor U8733 (N_8733,N_8303,N_8381);
and U8734 (N_8734,N_8288,N_8303);
xor U8735 (N_8735,N_8310,N_8305);
xnor U8736 (N_8736,N_8455,N_8457);
or U8737 (N_8737,N_8299,N_8491);
xor U8738 (N_8738,N_8311,N_8431);
and U8739 (N_8739,N_8349,N_8410);
xor U8740 (N_8740,N_8387,N_8382);
or U8741 (N_8741,N_8277,N_8304);
nand U8742 (N_8742,N_8433,N_8389);
nor U8743 (N_8743,N_8400,N_8313);
or U8744 (N_8744,N_8469,N_8354);
nand U8745 (N_8745,N_8263,N_8274);
or U8746 (N_8746,N_8260,N_8417);
nand U8747 (N_8747,N_8446,N_8291);
and U8748 (N_8748,N_8408,N_8422);
xor U8749 (N_8749,N_8311,N_8360);
or U8750 (N_8750,N_8559,N_8540);
nand U8751 (N_8751,N_8738,N_8502);
and U8752 (N_8752,N_8633,N_8687);
and U8753 (N_8753,N_8715,N_8577);
nor U8754 (N_8754,N_8599,N_8504);
xnor U8755 (N_8755,N_8629,N_8508);
or U8756 (N_8756,N_8509,N_8691);
xor U8757 (N_8757,N_8541,N_8544);
xnor U8758 (N_8758,N_8610,N_8628);
or U8759 (N_8759,N_8545,N_8594);
nand U8760 (N_8760,N_8620,N_8641);
nor U8761 (N_8761,N_8532,N_8636);
xnor U8762 (N_8762,N_8600,N_8713);
nor U8763 (N_8763,N_8548,N_8588);
and U8764 (N_8764,N_8646,N_8506);
xor U8765 (N_8765,N_8563,N_8745);
nand U8766 (N_8766,N_8717,N_8575);
xor U8767 (N_8767,N_8658,N_8688);
nand U8768 (N_8768,N_8520,N_8661);
and U8769 (N_8769,N_8573,N_8576);
nand U8770 (N_8770,N_8567,N_8719);
or U8771 (N_8771,N_8729,N_8511);
and U8772 (N_8772,N_8528,N_8693);
xnor U8773 (N_8773,N_8513,N_8530);
and U8774 (N_8774,N_8647,N_8521);
or U8775 (N_8775,N_8720,N_8624);
nand U8776 (N_8776,N_8663,N_8565);
or U8777 (N_8777,N_8527,N_8623);
xor U8778 (N_8778,N_8605,N_8664);
or U8779 (N_8779,N_8589,N_8615);
nand U8780 (N_8780,N_8604,N_8586);
or U8781 (N_8781,N_8700,N_8517);
nand U8782 (N_8782,N_8671,N_8710);
or U8783 (N_8783,N_8734,N_8564);
nor U8784 (N_8784,N_8744,N_8736);
xor U8785 (N_8785,N_8561,N_8674);
nor U8786 (N_8786,N_8602,N_8595);
xor U8787 (N_8787,N_8549,N_8670);
nor U8788 (N_8788,N_8657,N_8534);
or U8789 (N_8789,N_8731,N_8593);
nor U8790 (N_8790,N_8609,N_8660);
or U8791 (N_8791,N_8621,N_8676);
nand U8792 (N_8792,N_8737,N_8611);
nor U8793 (N_8793,N_8666,N_8578);
nand U8794 (N_8794,N_8617,N_8531);
nor U8795 (N_8795,N_8668,N_8742);
nor U8796 (N_8796,N_8603,N_8650);
or U8797 (N_8797,N_8568,N_8606);
or U8798 (N_8798,N_8550,N_8607);
or U8799 (N_8799,N_8644,N_8560);
or U8800 (N_8800,N_8716,N_8686);
and U8801 (N_8801,N_8536,N_8690);
nor U8802 (N_8802,N_8740,N_8672);
and U8803 (N_8803,N_8526,N_8743);
nor U8804 (N_8804,N_8659,N_8592);
xor U8805 (N_8805,N_8645,N_8537);
and U8806 (N_8806,N_8708,N_8634);
nand U8807 (N_8807,N_8590,N_8539);
or U8808 (N_8808,N_8709,N_8640);
nor U8809 (N_8809,N_8613,N_8630);
or U8810 (N_8810,N_8562,N_8656);
nor U8811 (N_8811,N_8639,N_8721);
nor U8812 (N_8812,N_8695,N_8648);
nand U8813 (N_8813,N_8678,N_8516);
nor U8814 (N_8814,N_8519,N_8701);
xnor U8815 (N_8815,N_8696,N_8748);
xnor U8816 (N_8816,N_8724,N_8677);
nand U8817 (N_8817,N_8582,N_8649);
nand U8818 (N_8818,N_8698,N_8705);
nand U8819 (N_8819,N_8538,N_8746);
nor U8820 (N_8820,N_8598,N_8553);
and U8821 (N_8821,N_8533,N_8706);
or U8822 (N_8822,N_8601,N_8591);
and U8823 (N_8823,N_8699,N_8570);
nor U8824 (N_8824,N_8529,N_8525);
and U8825 (N_8825,N_8718,N_8622);
nor U8826 (N_8826,N_8584,N_8684);
and U8827 (N_8827,N_8597,N_8707);
nand U8828 (N_8828,N_8714,N_8503);
or U8829 (N_8829,N_8667,N_8501);
nor U8830 (N_8830,N_8618,N_8711);
xnor U8831 (N_8831,N_8655,N_8524);
nand U8832 (N_8832,N_8518,N_8652);
nand U8833 (N_8833,N_8725,N_8683);
and U8834 (N_8834,N_8554,N_8510);
nand U8835 (N_8835,N_8583,N_8632);
nor U8836 (N_8836,N_8726,N_8739);
nor U8837 (N_8837,N_8523,N_8665);
xor U8838 (N_8838,N_8596,N_8585);
nor U8839 (N_8839,N_8619,N_8732);
or U8840 (N_8840,N_8728,N_8662);
nor U8841 (N_8841,N_8612,N_8733);
nand U8842 (N_8842,N_8542,N_8651);
and U8843 (N_8843,N_8653,N_8505);
nand U8844 (N_8844,N_8580,N_8638);
nand U8845 (N_8845,N_8723,N_8500);
nor U8846 (N_8846,N_8643,N_8626);
nand U8847 (N_8847,N_8625,N_8730);
nand U8848 (N_8848,N_8552,N_8551);
and U8849 (N_8849,N_8522,N_8703);
nor U8850 (N_8850,N_8543,N_8512);
xor U8851 (N_8851,N_8679,N_8692);
nand U8852 (N_8852,N_8555,N_8654);
xnor U8853 (N_8853,N_8581,N_8704);
xor U8854 (N_8854,N_8571,N_8569);
xor U8855 (N_8855,N_8749,N_8673);
nand U8856 (N_8856,N_8514,N_8557);
nor U8857 (N_8857,N_8702,N_8685);
nor U8858 (N_8858,N_8712,N_8547);
nand U8859 (N_8859,N_8587,N_8727);
and U8860 (N_8860,N_8697,N_8614);
or U8861 (N_8861,N_8642,N_8689);
xnor U8862 (N_8862,N_8566,N_8741);
or U8863 (N_8863,N_8579,N_8681);
or U8864 (N_8864,N_8546,N_8572);
xor U8865 (N_8865,N_8680,N_8558);
nand U8866 (N_8866,N_8608,N_8616);
nand U8867 (N_8867,N_8694,N_8722);
or U8868 (N_8868,N_8682,N_8635);
xor U8869 (N_8869,N_8556,N_8627);
or U8870 (N_8870,N_8675,N_8507);
xor U8871 (N_8871,N_8515,N_8669);
and U8872 (N_8872,N_8747,N_8574);
and U8873 (N_8873,N_8637,N_8735);
nor U8874 (N_8874,N_8535,N_8631);
nor U8875 (N_8875,N_8561,N_8659);
and U8876 (N_8876,N_8597,N_8534);
nor U8877 (N_8877,N_8655,N_8747);
nand U8878 (N_8878,N_8580,N_8720);
nor U8879 (N_8879,N_8624,N_8652);
nand U8880 (N_8880,N_8614,N_8535);
and U8881 (N_8881,N_8516,N_8690);
nor U8882 (N_8882,N_8747,N_8553);
nand U8883 (N_8883,N_8576,N_8529);
and U8884 (N_8884,N_8621,N_8602);
or U8885 (N_8885,N_8722,N_8606);
or U8886 (N_8886,N_8681,N_8646);
xor U8887 (N_8887,N_8728,N_8576);
nor U8888 (N_8888,N_8515,N_8711);
and U8889 (N_8889,N_8614,N_8501);
and U8890 (N_8890,N_8685,N_8509);
or U8891 (N_8891,N_8676,N_8702);
xnor U8892 (N_8892,N_8691,N_8527);
xnor U8893 (N_8893,N_8748,N_8621);
xnor U8894 (N_8894,N_8614,N_8645);
xnor U8895 (N_8895,N_8523,N_8708);
or U8896 (N_8896,N_8540,N_8740);
nand U8897 (N_8897,N_8507,N_8534);
or U8898 (N_8898,N_8602,N_8614);
nand U8899 (N_8899,N_8559,N_8712);
and U8900 (N_8900,N_8708,N_8603);
nand U8901 (N_8901,N_8663,N_8731);
and U8902 (N_8902,N_8520,N_8529);
nand U8903 (N_8903,N_8653,N_8536);
and U8904 (N_8904,N_8641,N_8592);
nand U8905 (N_8905,N_8581,N_8633);
xnor U8906 (N_8906,N_8579,N_8697);
or U8907 (N_8907,N_8663,N_8533);
and U8908 (N_8908,N_8647,N_8668);
xnor U8909 (N_8909,N_8590,N_8548);
and U8910 (N_8910,N_8741,N_8514);
nand U8911 (N_8911,N_8655,N_8694);
xor U8912 (N_8912,N_8655,N_8563);
nor U8913 (N_8913,N_8607,N_8500);
xnor U8914 (N_8914,N_8632,N_8571);
nor U8915 (N_8915,N_8658,N_8665);
and U8916 (N_8916,N_8642,N_8617);
nand U8917 (N_8917,N_8647,N_8626);
nand U8918 (N_8918,N_8738,N_8633);
and U8919 (N_8919,N_8722,N_8610);
xnor U8920 (N_8920,N_8595,N_8688);
and U8921 (N_8921,N_8643,N_8669);
or U8922 (N_8922,N_8505,N_8740);
nand U8923 (N_8923,N_8570,N_8597);
nand U8924 (N_8924,N_8663,N_8722);
or U8925 (N_8925,N_8732,N_8681);
and U8926 (N_8926,N_8599,N_8658);
nor U8927 (N_8927,N_8618,N_8557);
or U8928 (N_8928,N_8678,N_8622);
and U8929 (N_8929,N_8699,N_8624);
or U8930 (N_8930,N_8746,N_8690);
and U8931 (N_8931,N_8715,N_8610);
nand U8932 (N_8932,N_8622,N_8555);
nor U8933 (N_8933,N_8563,N_8643);
and U8934 (N_8934,N_8723,N_8521);
or U8935 (N_8935,N_8644,N_8661);
and U8936 (N_8936,N_8747,N_8717);
and U8937 (N_8937,N_8549,N_8664);
nand U8938 (N_8938,N_8553,N_8562);
nor U8939 (N_8939,N_8565,N_8508);
or U8940 (N_8940,N_8522,N_8537);
and U8941 (N_8941,N_8626,N_8679);
nor U8942 (N_8942,N_8591,N_8569);
nor U8943 (N_8943,N_8675,N_8617);
nor U8944 (N_8944,N_8558,N_8724);
and U8945 (N_8945,N_8517,N_8713);
and U8946 (N_8946,N_8562,N_8713);
nand U8947 (N_8947,N_8519,N_8679);
xnor U8948 (N_8948,N_8726,N_8519);
nor U8949 (N_8949,N_8642,N_8710);
or U8950 (N_8950,N_8686,N_8526);
xnor U8951 (N_8951,N_8650,N_8719);
nor U8952 (N_8952,N_8592,N_8729);
or U8953 (N_8953,N_8636,N_8670);
xor U8954 (N_8954,N_8545,N_8624);
and U8955 (N_8955,N_8505,N_8530);
nor U8956 (N_8956,N_8513,N_8694);
or U8957 (N_8957,N_8562,N_8500);
nand U8958 (N_8958,N_8677,N_8670);
and U8959 (N_8959,N_8660,N_8709);
or U8960 (N_8960,N_8689,N_8621);
nor U8961 (N_8961,N_8719,N_8625);
nand U8962 (N_8962,N_8722,N_8633);
or U8963 (N_8963,N_8613,N_8579);
nor U8964 (N_8964,N_8668,N_8596);
xnor U8965 (N_8965,N_8688,N_8714);
nor U8966 (N_8966,N_8502,N_8641);
or U8967 (N_8967,N_8728,N_8675);
or U8968 (N_8968,N_8516,N_8663);
nor U8969 (N_8969,N_8523,N_8731);
and U8970 (N_8970,N_8656,N_8739);
xor U8971 (N_8971,N_8563,N_8641);
nand U8972 (N_8972,N_8691,N_8631);
xor U8973 (N_8973,N_8738,N_8506);
or U8974 (N_8974,N_8657,N_8708);
or U8975 (N_8975,N_8517,N_8726);
or U8976 (N_8976,N_8670,N_8695);
or U8977 (N_8977,N_8580,N_8602);
and U8978 (N_8978,N_8510,N_8675);
or U8979 (N_8979,N_8579,N_8570);
and U8980 (N_8980,N_8543,N_8569);
and U8981 (N_8981,N_8601,N_8626);
nand U8982 (N_8982,N_8600,N_8531);
or U8983 (N_8983,N_8594,N_8608);
or U8984 (N_8984,N_8643,N_8697);
or U8985 (N_8985,N_8686,N_8629);
and U8986 (N_8986,N_8502,N_8596);
nand U8987 (N_8987,N_8502,N_8623);
xnor U8988 (N_8988,N_8698,N_8641);
nor U8989 (N_8989,N_8580,N_8659);
and U8990 (N_8990,N_8680,N_8732);
xor U8991 (N_8991,N_8572,N_8531);
and U8992 (N_8992,N_8645,N_8655);
and U8993 (N_8993,N_8626,N_8568);
or U8994 (N_8994,N_8500,N_8742);
nand U8995 (N_8995,N_8718,N_8706);
nand U8996 (N_8996,N_8561,N_8668);
xnor U8997 (N_8997,N_8638,N_8612);
nor U8998 (N_8998,N_8614,N_8576);
nor U8999 (N_8999,N_8682,N_8747);
and U9000 (N_9000,N_8981,N_8864);
or U9001 (N_9001,N_8897,N_8831);
and U9002 (N_9002,N_8996,N_8999);
nand U9003 (N_9003,N_8862,N_8966);
nand U9004 (N_9004,N_8881,N_8978);
xnor U9005 (N_9005,N_8816,N_8934);
nand U9006 (N_9006,N_8801,N_8988);
xor U9007 (N_9007,N_8766,N_8758);
nand U9008 (N_9008,N_8951,N_8783);
nor U9009 (N_9009,N_8891,N_8968);
and U9010 (N_9010,N_8770,N_8842);
xnor U9011 (N_9011,N_8798,N_8796);
nand U9012 (N_9012,N_8936,N_8892);
xnor U9013 (N_9013,N_8937,N_8850);
and U9014 (N_9014,N_8879,N_8789);
and U9015 (N_9015,N_8771,N_8808);
nand U9016 (N_9016,N_8753,N_8906);
nand U9017 (N_9017,N_8810,N_8956);
xor U9018 (N_9018,N_8839,N_8992);
and U9019 (N_9019,N_8953,N_8815);
or U9020 (N_9020,N_8822,N_8900);
xnor U9021 (N_9021,N_8994,N_8919);
and U9022 (N_9022,N_8792,N_8840);
nand U9023 (N_9023,N_8964,N_8991);
or U9024 (N_9024,N_8863,N_8969);
and U9025 (N_9025,N_8785,N_8977);
and U9026 (N_9026,N_8814,N_8846);
or U9027 (N_9027,N_8918,N_8800);
nor U9028 (N_9028,N_8779,N_8823);
and U9029 (N_9029,N_8847,N_8849);
nor U9030 (N_9030,N_8938,N_8843);
and U9031 (N_9031,N_8967,N_8835);
xnor U9032 (N_9032,N_8819,N_8837);
xor U9033 (N_9033,N_8914,N_8982);
xor U9034 (N_9034,N_8963,N_8760);
xnor U9035 (N_9035,N_8998,N_8921);
or U9036 (N_9036,N_8915,N_8876);
nor U9037 (N_9037,N_8941,N_8773);
nand U9038 (N_9038,N_8945,N_8909);
nor U9039 (N_9039,N_8916,N_8767);
and U9040 (N_9040,N_8948,N_8809);
and U9041 (N_9041,N_8777,N_8820);
nor U9042 (N_9042,N_8751,N_8857);
and U9043 (N_9043,N_8972,N_8954);
nand U9044 (N_9044,N_8889,N_8944);
nor U9045 (N_9045,N_8827,N_8973);
or U9046 (N_9046,N_8806,N_8959);
or U9047 (N_9047,N_8901,N_8917);
and U9048 (N_9048,N_8983,N_8899);
xnor U9049 (N_9049,N_8920,N_8828);
nor U9050 (N_9050,N_8926,N_8960);
xnor U9051 (N_9051,N_8946,N_8791);
xnor U9052 (N_9052,N_8790,N_8985);
nand U9053 (N_9053,N_8780,N_8979);
and U9054 (N_9054,N_8874,N_8860);
and U9055 (N_9055,N_8894,N_8905);
nor U9056 (N_9056,N_8765,N_8817);
nand U9057 (N_9057,N_8811,N_8883);
or U9058 (N_9058,N_8912,N_8976);
xor U9059 (N_9059,N_8872,N_8865);
nor U9060 (N_9060,N_8986,N_8995);
xnor U9061 (N_9061,N_8834,N_8805);
xor U9062 (N_9062,N_8768,N_8939);
xnor U9063 (N_9063,N_8825,N_8896);
or U9064 (N_9064,N_8804,N_8830);
or U9065 (N_9065,N_8778,N_8752);
nor U9066 (N_9066,N_8947,N_8975);
xor U9067 (N_9067,N_8755,N_8870);
nor U9068 (N_9068,N_8781,N_8833);
or U9069 (N_9069,N_8797,N_8772);
or U9070 (N_9070,N_8880,N_8756);
nor U9071 (N_9071,N_8826,N_8929);
xor U9072 (N_9072,N_8871,N_8885);
nor U9073 (N_9073,N_8869,N_8845);
or U9074 (N_9074,N_8861,N_8877);
and U9075 (N_9075,N_8793,N_8928);
nand U9076 (N_9076,N_8875,N_8787);
nor U9077 (N_9077,N_8930,N_8858);
xnor U9078 (N_9078,N_8931,N_8955);
and U9079 (N_9079,N_8990,N_8764);
nor U9080 (N_9080,N_8913,N_8952);
or U9081 (N_9081,N_8965,N_8878);
nor U9082 (N_9082,N_8813,N_8993);
and U9083 (N_9083,N_8759,N_8852);
nand U9084 (N_9084,N_8961,N_8898);
and U9085 (N_9085,N_8933,N_8868);
xor U9086 (N_9086,N_8924,N_8794);
nand U9087 (N_9087,N_8784,N_8786);
or U9088 (N_9088,N_8935,N_8859);
nor U9089 (N_9089,N_8855,N_8844);
nand U9090 (N_9090,N_8923,N_8775);
nand U9091 (N_9091,N_8754,N_8841);
nor U9092 (N_9092,N_8925,N_8895);
nand U9093 (N_9093,N_8927,N_8757);
xor U9094 (N_9094,N_8803,N_8949);
xnor U9095 (N_9095,N_8750,N_8854);
or U9096 (N_9096,N_8984,N_8971);
xnor U9097 (N_9097,N_8856,N_8886);
nor U9098 (N_9098,N_8873,N_8974);
and U9099 (N_9099,N_8890,N_8910);
or U9100 (N_9100,N_8997,N_8907);
and U9101 (N_9101,N_8818,N_8761);
nor U9102 (N_9102,N_8980,N_8902);
xnor U9103 (N_9103,N_8904,N_8987);
or U9104 (N_9104,N_8788,N_8957);
and U9105 (N_9105,N_8802,N_8888);
xnor U9106 (N_9106,N_8851,N_8884);
and U9107 (N_9107,N_8942,N_8763);
xor U9108 (N_9108,N_8943,N_8887);
or U9109 (N_9109,N_8807,N_8812);
nand U9110 (N_9110,N_8853,N_8911);
xor U9111 (N_9111,N_8824,N_8970);
or U9112 (N_9112,N_8903,N_8774);
nor U9113 (N_9113,N_8829,N_8848);
and U9114 (N_9114,N_8893,N_8882);
nand U9115 (N_9115,N_8799,N_8795);
nor U9116 (N_9116,N_8932,N_8836);
and U9117 (N_9117,N_8832,N_8769);
nor U9118 (N_9118,N_8866,N_8922);
nor U9119 (N_9119,N_8908,N_8958);
nand U9120 (N_9120,N_8762,N_8962);
nand U9121 (N_9121,N_8940,N_8821);
or U9122 (N_9122,N_8950,N_8867);
nor U9123 (N_9123,N_8776,N_8989);
and U9124 (N_9124,N_8838,N_8782);
and U9125 (N_9125,N_8756,N_8763);
nor U9126 (N_9126,N_8868,N_8889);
nand U9127 (N_9127,N_8761,N_8808);
or U9128 (N_9128,N_8862,N_8798);
or U9129 (N_9129,N_8857,N_8833);
xnor U9130 (N_9130,N_8751,N_8917);
and U9131 (N_9131,N_8802,N_8776);
or U9132 (N_9132,N_8848,N_8847);
and U9133 (N_9133,N_8777,N_8832);
nor U9134 (N_9134,N_8783,N_8797);
nor U9135 (N_9135,N_8899,N_8892);
or U9136 (N_9136,N_8914,N_8912);
nor U9137 (N_9137,N_8925,N_8755);
and U9138 (N_9138,N_8912,N_8881);
nor U9139 (N_9139,N_8752,N_8980);
nor U9140 (N_9140,N_8897,N_8919);
and U9141 (N_9141,N_8928,N_8785);
nand U9142 (N_9142,N_8898,N_8771);
and U9143 (N_9143,N_8864,N_8957);
xor U9144 (N_9144,N_8992,N_8796);
or U9145 (N_9145,N_8961,N_8855);
or U9146 (N_9146,N_8844,N_8960);
nand U9147 (N_9147,N_8788,N_8849);
xnor U9148 (N_9148,N_8962,N_8989);
nand U9149 (N_9149,N_8954,N_8927);
nand U9150 (N_9150,N_8842,N_8826);
and U9151 (N_9151,N_8965,N_8837);
nor U9152 (N_9152,N_8920,N_8814);
and U9153 (N_9153,N_8764,N_8847);
or U9154 (N_9154,N_8785,N_8787);
nor U9155 (N_9155,N_8884,N_8826);
xor U9156 (N_9156,N_8988,N_8823);
and U9157 (N_9157,N_8835,N_8842);
or U9158 (N_9158,N_8942,N_8984);
xnor U9159 (N_9159,N_8864,N_8826);
and U9160 (N_9160,N_8776,N_8941);
xor U9161 (N_9161,N_8953,N_8803);
nand U9162 (N_9162,N_8913,N_8767);
nand U9163 (N_9163,N_8823,N_8915);
nor U9164 (N_9164,N_8986,N_8949);
or U9165 (N_9165,N_8944,N_8971);
nor U9166 (N_9166,N_8764,N_8868);
nand U9167 (N_9167,N_8766,N_8969);
nor U9168 (N_9168,N_8851,N_8998);
nand U9169 (N_9169,N_8895,N_8990);
or U9170 (N_9170,N_8819,N_8753);
xnor U9171 (N_9171,N_8835,N_8961);
nor U9172 (N_9172,N_8798,N_8819);
nand U9173 (N_9173,N_8996,N_8786);
nor U9174 (N_9174,N_8810,N_8765);
nor U9175 (N_9175,N_8823,N_8934);
xnor U9176 (N_9176,N_8838,N_8893);
and U9177 (N_9177,N_8881,N_8999);
or U9178 (N_9178,N_8833,N_8780);
or U9179 (N_9179,N_8770,N_8793);
or U9180 (N_9180,N_8949,N_8752);
xor U9181 (N_9181,N_8815,N_8926);
nor U9182 (N_9182,N_8995,N_8793);
and U9183 (N_9183,N_8825,N_8865);
nand U9184 (N_9184,N_8854,N_8835);
xnor U9185 (N_9185,N_8972,N_8774);
nand U9186 (N_9186,N_8875,N_8796);
xor U9187 (N_9187,N_8778,N_8770);
or U9188 (N_9188,N_8825,N_8988);
nand U9189 (N_9189,N_8798,N_8922);
and U9190 (N_9190,N_8982,N_8977);
xnor U9191 (N_9191,N_8787,N_8814);
or U9192 (N_9192,N_8929,N_8914);
and U9193 (N_9193,N_8998,N_8829);
nand U9194 (N_9194,N_8866,N_8989);
nor U9195 (N_9195,N_8900,N_8845);
or U9196 (N_9196,N_8773,N_8832);
xor U9197 (N_9197,N_8891,N_8885);
nor U9198 (N_9198,N_8861,N_8883);
nor U9199 (N_9199,N_8752,N_8774);
and U9200 (N_9200,N_8803,N_8861);
nand U9201 (N_9201,N_8763,N_8879);
xor U9202 (N_9202,N_8981,N_8938);
xor U9203 (N_9203,N_8950,N_8827);
nor U9204 (N_9204,N_8827,N_8926);
and U9205 (N_9205,N_8764,N_8991);
xnor U9206 (N_9206,N_8901,N_8850);
xor U9207 (N_9207,N_8818,N_8910);
xor U9208 (N_9208,N_8778,N_8962);
xnor U9209 (N_9209,N_8899,N_8944);
xor U9210 (N_9210,N_8807,N_8951);
and U9211 (N_9211,N_8758,N_8776);
nand U9212 (N_9212,N_8988,N_8985);
xnor U9213 (N_9213,N_8818,N_8889);
and U9214 (N_9214,N_8981,N_8893);
xnor U9215 (N_9215,N_8787,N_8883);
xor U9216 (N_9216,N_8808,N_8872);
or U9217 (N_9217,N_8890,N_8812);
and U9218 (N_9218,N_8887,N_8795);
and U9219 (N_9219,N_8881,N_8852);
nor U9220 (N_9220,N_8765,N_8952);
nor U9221 (N_9221,N_8856,N_8905);
nand U9222 (N_9222,N_8890,N_8856);
nand U9223 (N_9223,N_8754,N_8786);
xnor U9224 (N_9224,N_8934,N_8952);
xnor U9225 (N_9225,N_8994,N_8781);
nor U9226 (N_9226,N_8877,N_8936);
xor U9227 (N_9227,N_8877,N_8945);
or U9228 (N_9228,N_8875,N_8960);
and U9229 (N_9229,N_8867,N_8833);
nor U9230 (N_9230,N_8887,N_8868);
or U9231 (N_9231,N_8851,N_8751);
nand U9232 (N_9232,N_8996,N_8773);
xnor U9233 (N_9233,N_8781,N_8982);
xor U9234 (N_9234,N_8774,N_8890);
xnor U9235 (N_9235,N_8762,N_8996);
and U9236 (N_9236,N_8840,N_8942);
xor U9237 (N_9237,N_8838,N_8891);
or U9238 (N_9238,N_8964,N_8955);
or U9239 (N_9239,N_8924,N_8839);
nand U9240 (N_9240,N_8787,N_8906);
nand U9241 (N_9241,N_8970,N_8779);
or U9242 (N_9242,N_8805,N_8989);
xnor U9243 (N_9243,N_8801,N_8996);
nor U9244 (N_9244,N_8965,N_8901);
xor U9245 (N_9245,N_8954,N_8844);
nand U9246 (N_9246,N_8757,N_8924);
and U9247 (N_9247,N_8863,N_8765);
and U9248 (N_9248,N_8751,N_8893);
nand U9249 (N_9249,N_8933,N_8988);
xor U9250 (N_9250,N_9239,N_9045);
or U9251 (N_9251,N_9039,N_9087);
nor U9252 (N_9252,N_9052,N_9155);
and U9253 (N_9253,N_9056,N_9013);
nand U9254 (N_9254,N_9125,N_9116);
or U9255 (N_9255,N_9195,N_9147);
xnor U9256 (N_9256,N_9191,N_9131);
or U9257 (N_9257,N_9219,N_9020);
or U9258 (N_9258,N_9236,N_9004);
xor U9259 (N_9259,N_9107,N_9229);
xor U9260 (N_9260,N_9213,N_9211);
nor U9261 (N_9261,N_9246,N_9225);
or U9262 (N_9262,N_9043,N_9210);
or U9263 (N_9263,N_9206,N_9145);
or U9264 (N_9264,N_9072,N_9134);
nand U9265 (N_9265,N_9033,N_9179);
nand U9266 (N_9266,N_9123,N_9159);
nand U9267 (N_9267,N_9241,N_9150);
or U9268 (N_9268,N_9140,N_9234);
xor U9269 (N_9269,N_9126,N_9129);
and U9270 (N_9270,N_9035,N_9040);
or U9271 (N_9271,N_9016,N_9009);
nor U9272 (N_9272,N_9231,N_9088);
or U9273 (N_9273,N_9201,N_9192);
nand U9274 (N_9274,N_9169,N_9008);
nand U9275 (N_9275,N_9074,N_9156);
or U9276 (N_9276,N_9012,N_9117);
nand U9277 (N_9277,N_9164,N_9180);
or U9278 (N_9278,N_9022,N_9160);
or U9279 (N_9279,N_9182,N_9063);
nand U9280 (N_9280,N_9217,N_9104);
xnor U9281 (N_9281,N_9103,N_9162);
xnor U9282 (N_9282,N_9200,N_9194);
nand U9283 (N_9283,N_9161,N_9207);
nor U9284 (N_9284,N_9077,N_9065);
and U9285 (N_9285,N_9142,N_9166);
nand U9286 (N_9286,N_9036,N_9174);
nand U9287 (N_9287,N_9235,N_9171);
xor U9288 (N_9288,N_9170,N_9027);
nand U9289 (N_9289,N_9054,N_9093);
and U9290 (N_9290,N_9069,N_9049);
nor U9291 (N_9291,N_9000,N_9078);
nand U9292 (N_9292,N_9220,N_9230);
xnor U9293 (N_9293,N_9098,N_9197);
nand U9294 (N_9294,N_9099,N_9202);
nand U9295 (N_9295,N_9173,N_9158);
or U9296 (N_9296,N_9190,N_9215);
xnor U9297 (N_9297,N_9238,N_9214);
xnor U9298 (N_9298,N_9151,N_9127);
nor U9299 (N_9299,N_9113,N_9044);
nor U9300 (N_9300,N_9095,N_9227);
nand U9301 (N_9301,N_9073,N_9122);
xnor U9302 (N_9302,N_9075,N_9153);
nor U9303 (N_9303,N_9080,N_9102);
nand U9304 (N_9304,N_9177,N_9055);
nand U9305 (N_9305,N_9030,N_9042);
nor U9306 (N_9306,N_9106,N_9165);
nand U9307 (N_9307,N_9146,N_9188);
nor U9308 (N_9308,N_9112,N_9224);
and U9309 (N_9309,N_9060,N_9248);
nand U9310 (N_9310,N_9081,N_9084);
or U9311 (N_9311,N_9071,N_9167);
nand U9312 (N_9312,N_9101,N_9244);
nor U9313 (N_9313,N_9133,N_9097);
and U9314 (N_9314,N_9168,N_9092);
nor U9315 (N_9315,N_9209,N_9006);
xnor U9316 (N_9316,N_9136,N_9110);
or U9317 (N_9317,N_9186,N_9070);
xor U9318 (N_9318,N_9066,N_9048);
or U9319 (N_9319,N_9120,N_9141);
and U9320 (N_9320,N_9083,N_9025);
nand U9321 (N_9321,N_9223,N_9187);
and U9322 (N_9322,N_9090,N_9059);
nand U9323 (N_9323,N_9181,N_9118);
nand U9324 (N_9324,N_9037,N_9011);
or U9325 (N_9325,N_9185,N_9094);
xnor U9326 (N_9326,N_9015,N_9163);
nand U9327 (N_9327,N_9024,N_9001);
nand U9328 (N_9328,N_9109,N_9061);
and U9329 (N_9329,N_9130,N_9137);
and U9330 (N_9330,N_9247,N_9047);
xor U9331 (N_9331,N_9029,N_9143);
or U9332 (N_9332,N_9124,N_9198);
and U9333 (N_9333,N_9237,N_9226);
xnor U9334 (N_9334,N_9062,N_9139);
or U9335 (N_9335,N_9135,N_9178);
nor U9336 (N_9336,N_9053,N_9208);
nand U9337 (N_9337,N_9100,N_9085);
and U9338 (N_9338,N_9058,N_9067);
xor U9339 (N_9339,N_9086,N_9076);
and U9340 (N_9340,N_9096,N_9019);
or U9341 (N_9341,N_9111,N_9157);
xor U9342 (N_9342,N_9216,N_9082);
and U9343 (N_9343,N_9014,N_9203);
nor U9344 (N_9344,N_9051,N_9046);
nand U9345 (N_9345,N_9149,N_9017);
nor U9346 (N_9346,N_9218,N_9172);
nand U9347 (N_9347,N_9023,N_9148);
and U9348 (N_9348,N_9119,N_9034);
nand U9349 (N_9349,N_9128,N_9057);
xnor U9350 (N_9350,N_9222,N_9064);
xnor U9351 (N_9351,N_9204,N_9007);
nand U9352 (N_9352,N_9249,N_9175);
nand U9353 (N_9353,N_9154,N_9221);
xnor U9354 (N_9354,N_9026,N_9183);
nor U9355 (N_9355,N_9232,N_9021);
or U9356 (N_9356,N_9184,N_9108);
nand U9357 (N_9357,N_9132,N_9152);
and U9358 (N_9358,N_9105,N_9068);
and U9359 (N_9359,N_9228,N_9196);
nand U9360 (N_9360,N_9193,N_9038);
or U9361 (N_9361,N_9028,N_9242);
or U9362 (N_9362,N_9114,N_9243);
and U9363 (N_9363,N_9003,N_9138);
nor U9364 (N_9364,N_9010,N_9005);
nand U9365 (N_9365,N_9089,N_9079);
and U9366 (N_9366,N_9050,N_9018);
and U9367 (N_9367,N_9144,N_9240);
nand U9368 (N_9368,N_9233,N_9245);
and U9369 (N_9369,N_9176,N_9121);
xnor U9370 (N_9370,N_9199,N_9115);
nor U9371 (N_9371,N_9002,N_9032);
and U9372 (N_9372,N_9041,N_9031);
and U9373 (N_9373,N_9091,N_9189);
xor U9374 (N_9374,N_9205,N_9212);
nor U9375 (N_9375,N_9223,N_9007);
or U9376 (N_9376,N_9210,N_9032);
and U9377 (N_9377,N_9052,N_9072);
or U9378 (N_9378,N_9102,N_9099);
nand U9379 (N_9379,N_9044,N_9171);
and U9380 (N_9380,N_9085,N_9136);
and U9381 (N_9381,N_9029,N_9015);
nor U9382 (N_9382,N_9231,N_9085);
or U9383 (N_9383,N_9119,N_9219);
xnor U9384 (N_9384,N_9102,N_9056);
or U9385 (N_9385,N_9040,N_9241);
and U9386 (N_9386,N_9244,N_9207);
and U9387 (N_9387,N_9082,N_9090);
or U9388 (N_9388,N_9067,N_9148);
and U9389 (N_9389,N_9111,N_9200);
nand U9390 (N_9390,N_9084,N_9091);
or U9391 (N_9391,N_9108,N_9149);
nor U9392 (N_9392,N_9003,N_9198);
nand U9393 (N_9393,N_9177,N_9078);
xnor U9394 (N_9394,N_9039,N_9025);
xor U9395 (N_9395,N_9077,N_9147);
and U9396 (N_9396,N_9107,N_9061);
xnor U9397 (N_9397,N_9221,N_9116);
nand U9398 (N_9398,N_9105,N_9020);
nand U9399 (N_9399,N_9221,N_9130);
nor U9400 (N_9400,N_9161,N_9048);
nand U9401 (N_9401,N_9116,N_9074);
and U9402 (N_9402,N_9212,N_9055);
and U9403 (N_9403,N_9108,N_9195);
and U9404 (N_9404,N_9236,N_9124);
nor U9405 (N_9405,N_9020,N_9153);
or U9406 (N_9406,N_9202,N_9051);
or U9407 (N_9407,N_9111,N_9235);
xor U9408 (N_9408,N_9228,N_9152);
xor U9409 (N_9409,N_9212,N_9154);
or U9410 (N_9410,N_9145,N_9047);
nor U9411 (N_9411,N_9143,N_9033);
and U9412 (N_9412,N_9052,N_9174);
nand U9413 (N_9413,N_9131,N_9152);
xor U9414 (N_9414,N_9235,N_9021);
and U9415 (N_9415,N_9042,N_9120);
nor U9416 (N_9416,N_9222,N_9137);
and U9417 (N_9417,N_9197,N_9007);
nand U9418 (N_9418,N_9021,N_9178);
or U9419 (N_9419,N_9195,N_9087);
or U9420 (N_9420,N_9142,N_9018);
nor U9421 (N_9421,N_9161,N_9216);
nand U9422 (N_9422,N_9065,N_9232);
or U9423 (N_9423,N_9128,N_9141);
xnor U9424 (N_9424,N_9190,N_9101);
and U9425 (N_9425,N_9001,N_9138);
nor U9426 (N_9426,N_9215,N_9138);
xnor U9427 (N_9427,N_9037,N_9038);
xnor U9428 (N_9428,N_9166,N_9128);
nand U9429 (N_9429,N_9094,N_9093);
or U9430 (N_9430,N_9193,N_9029);
and U9431 (N_9431,N_9243,N_9085);
and U9432 (N_9432,N_9210,N_9097);
xnor U9433 (N_9433,N_9116,N_9180);
nor U9434 (N_9434,N_9000,N_9065);
and U9435 (N_9435,N_9218,N_9206);
and U9436 (N_9436,N_9164,N_9156);
xor U9437 (N_9437,N_9241,N_9117);
nor U9438 (N_9438,N_9033,N_9155);
nand U9439 (N_9439,N_9013,N_9018);
nand U9440 (N_9440,N_9196,N_9092);
nand U9441 (N_9441,N_9158,N_9155);
and U9442 (N_9442,N_9056,N_9110);
and U9443 (N_9443,N_9129,N_9065);
nand U9444 (N_9444,N_9060,N_9228);
xnor U9445 (N_9445,N_9000,N_9132);
nor U9446 (N_9446,N_9048,N_9060);
nand U9447 (N_9447,N_9047,N_9021);
xnor U9448 (N_9448,N_9083,N_9078);
nor U9449 (N_9449,N_9214,N_9072);
nand U9450 (N_9450,N_9052,N_9181);
or U9451 (N_9451,N_9204,N_9073);
nor U9452 (N_9452,N_9143,N_9224);
or U9453 (N_9453,N_9169,N_9144);
or U9454 (N_9454,N_9193,N_9135);
nand U9455 (N_9455,N_9074,N_9041);
nor U9456 (N_9456,N_9061,N_9141);
nand U9457 (N_9457,N_9015,N_9076);
xnor U9458 (N_9458,N_9170,N_9098);
nor U9459 (N_9459,N_9126,N_9107);
or U9460 (N_9460,N_9181,N_9209);
and U9461 (N_9461,N_9080,N_9122);
nor U9462 (N_9462,N_9096,N_9086);
or U9463 (N_9463,N_9030,N_9159);
xnor U9464 (N_9464,N_9052,N_9111);
xnor U9465 (N_9465,N_9137,N_9124);
xnor U9466 (N_9466,N_9246,N_9182);
and U9467 (N_9467,N_9158,N_9114);
nor U9468 (N_9468,N_9060,N_9138);
nand U9469 (N_9469,N_9177,N_9206);
or U9470 (N_9470,N_9012,N_9131);
or U9471 (N_9471,N_9163,N_9150);
nor U9472 (N_9472,N_9223,N_9028);
or U9473 (N_9473,N_9153,N_9240);
or U9474 (N_9474,N_9054,N_9069);
and U9475 (N_9475,N_9197,N_9127);
xnor U9476 (N_9476,N_9240,N_9123);
nand U9477 (N_9477,N_9029,N_9105);
nand U9478 (N_9478,N_9168,N_9187);
nor U9479 (N_9479,N_9154,N_9165);
xnor U9480 (N_9480,N_9213,N_9130);
or U9481 (N_9481,N_9029,N_9068);
nor U9482 (N_9482,N_9014,N_9243);
or U9483 (N_9483,N_9106,N_9146);
nor U9484 (N_9484,N_9169,N_9182);
xnor U9485 (N_9485,N_9202,N_9243);
nand U9486 (N_9486,N_9069,N_9152);
and U9487 (N_9487,N_9097,N_9100);
and U9488 (N_9488,N_9155,N_9208);
and U9489 (N_9489,N_9046,N_9129);
xnor U9490 (N_9490,N_9008,N_9179);
or U9491 (N_9491,N_9126,N_9181);
nor U9492 (N_9492,N_9218,N_9099);
nor U9493 (N_9493,N_9196,N_9167);
nor U9494 (N_9494,N_9145,N_9175);
or U9495 (N_9495,N_9024,N_9025);
nor U9496 (N_9496,N_9122,N_9074);
xnor U9497 (N_9497,N_9108,N_9133);
nor U9498 (N_9498,N_9178,N_9125);
or U9499 (N_9499,N_9098,N_9020);
nor U9500 (N_9500,N_9423,N_9324);
nor U9501 (N_9501,N_9274,N_9397);
xnor U9502 (N_9502,N_9372,N_9365);
or U9503 (N_9503,N_9474,N_9347);
or U9504 (N_9504,N_9335,N_9447);
and U9505 (N_9505,N_9269,N_9430);
nor U9506 (N_9506,N_9484,N_9273);
xnor U9507 (N_9507,N_9344,N_9434);
xor U9508 (N_9508,N_9316,N_9407);
nand U9509 (N_9509,N_9464,N_9280);
nor U9510 (N_9510,N_9497,N_9440);
or U9511 (N_9511,N_9279,N_9353);
and U9512 (N_9512,N_9399,N_9450);
nor U9513 (N_9513,N_9482,N_9339);
xnor U9514 (N_9514,N_9322,N_9268);
or U9515 (N_9515,N_9251,N_9377);
nor U9516 (N_9516,N_9394,N_9432);
or U9517 (N_9517,N_9329,N_9479);
nor U9518 (N_9518,N_9414,N_9486);
nand U9519 (N_9519,N_9402,N_9388);
nor U9520 (N_9520,N_9313,N_9426);
or U9521 (N_9521,N_9328,N_9345);
and U9522 (N_9522,N_9356,N_9431);
nor U9523 (N_9523,N_9265,N_9258);
or U9524 (N_9524,N_9266,N_9462);
xnor U9525 (N_9525,N_9315,N_9254);
nand U9526 (N_9526,N_9460,N_9375);
nor U9527 (N_9527,N_9400,N_9470);
and U9528 (N_9528,N_9491,N_9255);
or U9529 (N_9529,N_9455,N_9459);
xor U9530 (N_9530,N_9391,N_9376);
nand U9531 (N_9531,N_9495,N_9342);
or U9532 (N_9532,N_9468,N_9349);
nand U9533 (N_9533,N_9308,N_9381);
nor U9534 (N_9534,N_9257,N_9272);
nor U9535 (N_9535,N_9469,N_9314);
and U9536 (N_9536,N_9261,N_9379);
or U9537 (N_9537,N_9312,N_9436);
nand U9538 (N_9538,N_9286,N_9318);
and U9539 (N_9539,N_9403,N_9362);
or U9540 (N_9540,N_9368,N_9374);
or U9541 (N_9541,N_9338,N_9435);
and U9542 (N_9542,N_9276,N_9300);
nor U9543 (N_9543,N_9350,N_9417);
and U9544 (N_9544,N_9478,N_9395);
xor U9545 (N_9545,N_9461,N_9310);
or U9546 (N_9546,N_9446,N_9492);
nand U9547 (N_9547,N_9343,N_9260);
nor U9548 (N_9548,N_9393,N_9369);
nor U9549 (N_9549,N_9442,N_9320);
and U9550 (N_9550,N_9360,N_9364);
or U9551 (N_9551,N_9443,N_9351);
or U9552 (N_9552,N_9404,N_9421);
nand U9553 (N_9553,N_9493,N_9444);
or U9554 (N_9554,N_9334,N_9454);
nor U9555 (N_9555,N_9389,N_9428);
xor U9556 (N_9556,N_9277,N_9285);
nor U9557 (N_9557,N_9311,N_9283);
nor U9558 (N_9558,N_9263,N_9458);
nor U9559 (N_9559,N_9386,N_9477);
and U9560 (N_9560,N_9437,N_9291);
and U9561 (N_9561,N_9467,N_9472);
nor U9562 (N_9562,N_9448,N_9326);
and U9563 (N_9563,N_9418,N_9358);
or U9564 (N_9564,N_9352,N_9262);
and U9565 (N_9565,N_9485,N_9433);
nand U9566 (N_9566,N_9259,N_9439);
or U9567 (N_9567,N_9333,N_9449);
xnor U9568 (N_9568,N_9411,N_9267);
xor U9569 (N_9569,N_9357,N_9294);
and U9570 (N_9570,N_9270,N_9271);
or U9571 (N_9571,N_9396,N_9410);
xnor U9572 (N_9572,N_9275,N_9496);
nor U9573 (N_9573,N_9494,N_9385);
xnor U9574 (N_9574,N_9302,N_9378);
nor U9575 (N_9575,N_9346,N_9336);
nand U9576 (N_9576,N_9292,N_9340);
nor U9577 (N_9577,N_9419,N_9405);
or U9578 (N_9578,N_9373,N_9409);
xor U9579 (N_9579,N_9489,N_9383);
and U9580 (N_9580,N_9398,N_9361);
xnor U9581 (N_9581,N_9288,N_9457);
and U9582 (N_9582,N_9284,N_9250);
nor U9583 (N_9583,N_9319,N_9264);
xor U9584 (N_9584,N_9427,N_9367);
xnor U9585 (N_9585,N_9330,N_9317);
or U9586 (N_9586,N_9281,N_9321);
or U9587 (N_9587,N_9382,N_9390);
xnor U9588 (N_9588,N_9278,N_9303);
or U9589 (N_9589,N_9476,N_9499);
and U9590 (N_9590,N_9453,N_9387);
or U9591 (N_9591,N_9256,N_9465);
nor U9592 (N_9592,N_9416,N_9293);
nor U9593 (N_9593,N_9392,N_9425);
and U9594 (N_9594,N_9498,N_9441);
xor U9595 (N_9595,N_9299,N_9384);
and U9596 (N_9596,N_9413,N_9354);
xor U9597 (N_9597,N_9355,N_9253);
xnor U9598 (N_9598,N_9420,N_9473);
xnor U9599 (N_9599,N_9296,N_9422);
and U9600 (N_9600,N_9323,N_9289);
xnor U9601 (N_9601,N_9456,N_9438);
xor U9602 (N_9602,N_9401,N_9483);
xnor U9603 (N_9603,N_9463,N_9406);
and U9604 (N_9604,N_9301,N_9487);
xor U9605 (N_9605,N_9370,N_9252);
nand U9606 (N_9606,N_9475,N_9471);
and U9607 (N_9607,N_9412,N_9305);
or U9608 (N_9608,N_9332,N_9366);
xor U9609 (N_9609,N_9408,N_9327);
and U9610 (N_9610,N_9287,N_9480);
and U9611 (N_9611,N_9331,N_9466);
nand U9612 (N_9612,N_9488,N_9282);
xnor U9613 (N_9613,N_9298,N_9337);
nand U9614 (N_9614,N_9325,N_9445);
nand U9615 (N_9615,N_9415,N_9424);
and U9616 (N_9616,N_9451,N_9297);
nor U9617 (N_9617,N_9307,N_9304);
nor U9618 (N_9618,N_9359,N_9306);
nor U9619 (N_9619,N_9348,N_9290);
xor U9620 (N_9620,N_9452,N_9371);
or U9621 (N_9621,N_9481,N_9490);
xor U9622 (N_9622,N_9341,N_9429);
nand U9623 (N_9623,N_9309,N_9380);
nor U9624 (N_9624,N_9295,N_9363);
and U9625 (N_9625,N_9266,N_9428);
or U9626 (N_9626,N_9442,N_9330);
nor U9627 (N_9627,N_9467,N_9318);
xnor U9628 (N_9628,N_9375,N_9381);
nand U9629 (N_9629,N_9434,N_9264);
nand U9630 (N_9630,N_9357,N_9419);
and U9631 (N_9631,N_9333,N_9337);
xnor U9632 (N_9632,N_9291,N_9376);
xor U9633 (N_9633,N_9301,N_9298);
nand U9634 (N_9634,N_9491,N_9472);
and U9635 (N_9635,N_9423,N_9269);
nor U9636 (N_9636,N_9387,N_9444);
and U9637 (N_9637,N_9255,N_9276);
and U9638 (N_9638,N_9378,N_9497);
xnor U9639 (N_9639,N_9468,N_9265);
and U9640 (N_9640,N_9370,N_9446);
nand U9641 (N_9641,N_9333,N_9488);
xnor U9642 (N_9642,N_9413,N_9493);
nand U9643 (N_9643,N_9477,N_9457);
nand U9644 (N_9644,N_9273,N_9491);
nor U9645 (N_9645,N_9472,N_9432);
xor U9646 (N_9646,N_9451,N_9313);
nand U9647 (N_9647,N_9395,N_9325);
and U9648 (N_9648,N_9316,N_9259);
xnor U9649 (N_9649,N_9258,N_9423);
and U9650 (N_9650,N_9362,N_9325);
nand U9651 (N_9651,N_9413,N_9346);
and U9652 (N_9652,N_9404,N_9340);
nand U9653 (N_9653,N_9252,N_9326);
xnor U9654 (N_9654,N_9292,N_9380);
and U9655 (N_9655,N_9476,N_9401);
xor U9656 (N_9656,N_9498,N_9275);
nor U9657 (N_9657,N_9332,N_9401);
nand U9658 (N_9658,N_9450,N_9493);
nand U9659 (N_9659,N_9405,N_9350);
or U9660 (N_9660,N_9392,N_9257);
xor U9661 (N_9661,N_9463,N_9493);
nor U9662 (N_9662,N_9275,N_9456);
nand U9663 (N_9663,N_9477,N_9449);
and U9664 (N_9664,N_9428,N_9286);
nand U9665 (N_9665,N_9452,N_9482);
xor U9666 (N_9666,N_9276,N_9265);
nand U9667 (N_9667,N_9439,N_9278);
or U9668 (N_9668,N_9343,N_9464);
and U9669 (N_9669,N_9355,N_9282);
or U9670 (N_9670,N_9441,N_9384);
or U9671 (N_9671,N_9487,N_9490);
nand U9672 (N_9672,N_9336,N_9401);
and U9673 (N_9673,N_9289,N_9251);
nor U9674 (N_9674,N_9324,N_9343);
and U9675 (N_9675,N_9323,N_9295);
and U9676 (N_9676,N_9382,N_9365);
nand U9677 (N_9677,N_9427,N_9414);
nor U9678 (N_9678,N_9418,N_9400);
xnor U9679 (N_9679,N_9416,N_9279);
xnor U9680 (N_9680,N_9298,N_9490);
or U9681 (N_9681,N_9369,N_9394);
nor U9682 (N_9682,N_9457,N_9435);
and U9683 (N_9683,N_9393,N_9449);
xor U9684 (N_9684,N_9343,N_9292);
and U9685 (N_9685,N_9417,N_9389);
xor U9686 (N_9686,N_9376,N_9486);
and U9687 (N_9687,N_9262,N_9484);
or U9688 (N_9688,N_9407,N_9497);
nor U9689 (N_9689,N_9318,N_9291);
or U9690 (N_9690,N_9494,N_9484);
nand U9691 (N_9691,N_9492,N_9350);
nor U9692 (N_9692,N_9326,N_9282);
nand U9693 (N_9693,N_9364,N_9404);
and U9694 (N_9694,N_9360,N_9473);
nor U9695 (N_9695,N_9420,N_9359);
xnor U9696 (N_9696,N_9335,N_9402);
and U9697 (N_9697,N_9336,N_9488);
nand U9698 (N_9698,N_9390,N_9469);
nand U9699 (N_9699,N_9475,N_9395);
nor U9700 (N_9700,N_9369,N_9392);
nand U9701 (N_9701,N_9488,N_9456);
nor U9702 (N_9702,N_9367,N_9300);
nand U9703 (N_9703,N_9360,N_9270);
or U9704 (N_9704,N_9455,N_9444);
nand U9705 (N_9705,N_9329,N_9264);
nor U9706 (N_9706,N_9402,N_9401);
nand U9707 (N_9707,N_9432,N_9294);
and U9708 (N_9708,N_9275,N_9323);
xnor U9709 (N_9709,N_9276,N_9281);
xnor U9710 (N_9710,N_9272,N_9317);
and U9711 (N_9711,N_9448,N_9370);
nor U9712 (N_9712,N_9281,N_9363);
or U9713 (N_9713,N_9279,N_9314);
nand U9714 (N_9714,N_9252,N_9490);
xor U9715 (N_9715,N_9347,N_9369);
xor U9716 (N_9716,N_9384,N_9495);
or U9717 (N_9717,N_9267,N_9425);
nor U9718 (N_9718,N_9257,N_9340);
nand U9719 (N_9719,N_9300,N_9413);
and U9720 (N_9720,N_9377,N_9366);
and U9721 (N_9721,N_9452,N_9348);
nor U9722 (N_9722,N_9335,N_9407);
nor U9723 (N_9723,N_9302,N_9289);
xor U9724 (N_9724,N_9449,N_9273);
nor U9725 (N_9725,N_9411,N_9362);
xnor U9726 (N_9726,N_9390,N_9480);
xnor U9727 (N_9727,N_9260,N_9312);
or U9728 (N_9728,N_9347,N_9397);
and U9729 (N_9729,N_9316,N_9262);
nor U9730 (N_9730,N_9345,N_9486);
nor U9731 (N_9731,N_9378,N_9274);
or U9732 (N_9732,N_9305,N_9453);
or U9733 (N_9733,N_9480,N_9362);
or U9734 (N_9734,N_9439,N_9497);
xnor U9735 (N_9735,N_9251,N_9313);
or U9736 (N_9736,N_9439,N_9479);
nand U9737 (N_9737,N_9495,N_9381);
xnor U9738 (N_9738,N_9482,N_9373);
or U9739 (N_9739,N_9439,N_9424);
or U9740 (N_9740,N_9333,N_9378);
xnor U9741 (N_9741,N_9498,N_9387);
nor U9742 (N_9742,N_9337,N_9299);
nor U9743 (N_9743,N_9257,N_9409);
nand U9744 (N_9744,N_9419,N_9476);
xnor U9745 (N_9745,N_9306,N_9332);
xnor U9746 (N_9746,N_9390,N_9295);
nor U9747 (N_9747,N_9352,N_9307);
and U9748 (N_9748,N_9252,N_9352);
and U9749 (N_9749,N_9358,N_9454);
or U9750 (N_9750,N_9670,N_9610);
nand U9751 (N_9751,N_9500,N_9517);
or U9752 (N_9752,N_9595,N_9544);
nand U9753 (N_9753,N_9512,N_9515);
nand U9754 (N_9754,N_9693,N_9746);
xnor U9755 (N_9755,N_9502,N_9716);
nor U9756 (N_9756,N_9576,N_9550);
nor U9757 (N_9757,N_9538,N_9501);
nor U9758 (N_9758,N_9700,N_9727);
xor U9759 (N_9759,N_9547,N_9667);
xor U9760 (N_9760,N_9702,N_9594);
nor U9761 (N_9761,N_9505,N_9589);
nor U9762 (N_9762,N_9634,N_9730);
nor U9763 (N_9763,N_9696,N_9587);
or U9764 (N_9764,N_9666,N_9642);
nand U9765 (N_9765,N_9749,N_9556);
xor U9766 (N_9766,N_9643,N_9518);
nand U9767 (N_9767,N_9560,N_9728);
and U9768 (N_9768,N_9664,N_9529);
xor U9769 (N_9769,N_9718,N_9729);
xor U9770 (N_9770,N_9720,N_9735);
xor U9771 (N_9771,N_9606,N_9504);
or U9772 (N_9772,N_9740,N_9654);
or U9773 (N_9773,N_9627,N_9508);
and U9774 (N_9774,N_9585,N_9733);
xor U9775 (N_9775,N_9710,N_9527);
or U9776 (N_9776,N_9579,N_9690);
nor U9777 (N_9777,N_9531,N_9588);
and U9778 (N_9778,N_9640,N_9566);
and U9779 (N_9779,N_9623,N_9682);
nand U9780 (N_9780,N_9598,N_9676);
and U9781 (N_9781,N_9692,N_9711);
or U9782 (N_9782,N_9680,N_9591);
xnor U9783 (N_9783,N_9668,N_9510);
or U9784 (N_9784,N_9705,N_9611);
nor U9785 (N_9785,N_9562,N_9715);
nor U9786 (N_9786,N_9632,N_9708);
nand U9787 (N_9787,N_9673,N_9524);
xor U9788 (N_9788,N_9563,N_9565);
xnor U9789 (N_9789,N_9537,N_9603);
or U9790 (N_9790,N_9635,N_9536);
or U9791 (N_9791,N_9613,N_9584);
or U9792 (N_9792,N_9561,N_9549);
nor U9793 (N_9793,N_9558,N_9726);
xnor U9794 (N_9794,N_9701,N_9590);
and U9795 (N_9795,N_9567,N_9638);
or U9796 (N_9796,N_9674,N_9507);
and U9797 (N_9797,N_9678,N_9521);
or U9798 (N_9798,N_9637,N_9636);
nor U9799 (N_9799,N_9712,N_9619);
xnor U9800 (N_9800,N_9514,N_9628);
and U9801 (N_9801,N_9543,N_9511);
nor U9802 (N_9802,N_9554,N_9742);
nand U9803 (N_9803,N_9652,N_9645);
xor U9804 (N_9804,N_9745,N_9631);
nor U9805 (N_9805,N_9719,N_9665);
xnor U9806 (N_9806,N_9723,N_9659);
xnor U9807 (N_9807,N_9699,N_9626);
xor U9808 (N_9808,N_9734,N_9681);
nor U9809 (N_9809,N_9675,N_9657);
and U9810 (N_9810,N_9703,N_9672);
nand U9811 (N_9811,N_9574,N_9630);
nor U9812 (N_9812,N_9540,N_9607);
or U9813 (N_9813,N_9622,N_9564);
xnor U9814 (N_9814,N_9533,N_9687);
and U9815 (N_9815,N_9620,N_9706);
xor U9816 (N_9816,N_9684,N_9572);
or U9817 (N_9817,N_9714,N_9707);
xor U9818 (N_9818,N_9597,N_9722);
nor U9819 (N_9819,N_9506,N_9557);
xor U9820 (N_9820,N_9534,N_9617);
nor U9821 (N_9821,N_9651,N_9614);
or U9822 (N_9822,N_9523,N_9581);
and U9823 (N_9823,N_9641,N_9609);
xnor U9824 (N_9824,N_9577,N_9525);
xnor U9825 (N_9825,N_9648,N_9522);
xnor U9826 (N_9826,N_9748,N_9644);
nand U9827 (N_9827,N_9592,N_9530);
or U9828 (N_9828,N_9671,N_9615);
nor U9829 (N_9829,N_9583,N_9503);
or U9830 (N_9830,N_9689,N_9526);
and U9831 (N_9831,N_9736,N_9513);
nand U9832 (N_9832,N_9647,N_9639);
nand U9833 (N_9833,N_9616,N_9688);
nor U9834 (N_9834,N_9509,N_9545);
xnor U9835 (N_9835,N_9605,N_9582);
or U9836 (N_9836,N_9731,N_9709);
nor U9837 (N_9837,N_9653,N_9516);
xnor U9838 (N_9838,N_9570,N_9571);
or U9839 (N_9839,N_9599,N_9621);
xor U9840 (N_9840,N_9629,N_9725);
nand U9841 (N_9841,N_9649,N_9656);
or U9842 (N_9842,N_9542,N_9698);
or U9843 (N_9843,N_9559,N_9552);
and U9844 (N_9844,N_9679,N_9669);
nor U9845 (N_9845,N_9553,N_9608);
nor U9846 (N_9846,N_9593,N_9743);
nand U9847 (N_9847,N_9633,N_9721);
nand U9848 (N_9848,N_9624,N_9650);
and U9849 (N_9849,N_9658,N_9578);
nor U9850 (N_9850,N_9655,N_9575);
nor U9851 (N_9851,N_9569,N_9618);
xnor U9852 (N_9852,N_9663,N_9535);
or U9853 (N_9853,N_9580,N_9738);
and U9854 (N_9854,N_9541,N_9697);
nand U9855 (N_9855,N_9685,N_9519);
nand U9856 (N_9856,N_9737,N_9532);
or U9857 (N_9857,N_9604,N_9717);
and U9858 (N_9858,N_9596,N_9612);
xor U9859 (N_9859,N_9695,N_9602);
and U9860 (N_9860,N_9683,N_9586);
nor U9861 (N_9861,N_9520,N_9694);
and U9862 (N_9862,N_9539,N_9741);
nor U9863 (N_9863,N_9691,N_9713);
nand U9864 (N_9864,N_9601,N_9661);
and U9865 (N_9865,N_9548,N_9646);
and U9866 (N_9866,N_9704,N_9747);
xnor U9867 (N_9867,N_9528,N_9662);
and U9868 (N_9868,N_9625,N_9739);
nand U9869 (N_9869,N_9600,N_9677);
nand U9870 (N_9870,N_9546,N_9744);
xnor U9871 (N_9871,N_9660,N_9686);
and U9872 (N_9872,N_9568,N_9555);
and U9873 (N_9873,N_9724,N_9551);
or U9874 (N_9874,N_9732,N_9573);
nor U9875 (N_9875,N_9536,N_9659);
and U9876 (N_9876,N_9634,N_9631);
or U9877 (N_9877,N_9563,N_9695);
and U9878 (N_9878,N_9667,N_9598);
xor U9879 (N_9879,N_9682,N_9730);
and U9880 (N_9880,N_9544,N_9603);
xnor U9881 (N_9881,N_9572,N_9686);
xnor U9882 (N_9882,N_9612,N_9517);
nand U9883 (N_9883,N_9686,N_9659);
or U9884 (N_9884,N_9685,N_9608);
nor U9885 (N_9885,N_9742,N_9749);
nand U9886 (N_9886,N_9635,N_9584);
and U9887 (N_9887,N_9540,N_9692);
nor U9888 (N_9888,N_9528,N_9639);
xnor U9889 (N_9889,N_9666,N_9744);
and U9890 (N_9890,N_9590,N_9650);
nor U9891 (N_9891,N_9612,N_9694);
or U9892 (N_9892,N_9662,N_9647);
nor U9893 (N_9893,N_9530,N_9721);
or U9894 (N_9894,N_9585,N_9601);
nand U9895 (N_9895,N_9674,N_9610);
and U9896 (N_9896,N_9700,N_9509);
and U9897 (N_9897,N_9556,N_9676);
or U9898 (N_9898,N_9527,N_9513);
nor U9899 (N_9899,N_9534,N_9614);
nor U9900 (N_9900,N_9749,N_9553);
or U9901 (N_9901,N_9600,N_9650);
xor U9902 (N_9902,N_9641,N_9564);
nor U9903 (N_9903,N_9715,N_9607);
and U9904 (N_9904,N_9644,N_9540);
or U9905 (N_9905,N_9592,N_9590);
or U9906 (N_9906,N_9597,N_9627);
nor U9907 (N_9907,N_9589,N_9565);
xor U9908 (N_9908,N_9736,N_9642);
or U9909 (N_9909,N_9556,N_9623);
nor U9910 (N_9910,N_9552,N_9519);
and U9911 (N_9911,N_9688,N_9503);
nand U9912 (N_9912,N_9732,N_9633);
nand U9913 (N_9913,N_9697,N_9737);
xor U9914 (N_9914,N_9742,N_9547);
xor U9915 (N_9915,N_9604,N_9570);
xor U9916 (N_9916,N_9732,N_9666);
nand U9917 (N_9917,N_9570,N_9694);
nand U9918 (N_9918,N_9653,N_9622);
nand U9919 (N_9919,N_9738,N_9717);
and U9920 (N_9920,N_9658,N_9641);
nand U9921 (N_9921,N_9614,N_9729);
and U9922 (N_9922,N_9716,N_9558);
nor U9923 (N_9923,N_9630,N_9575);
and U9924 (N_9924,N_9533,N_9578);
xor U9925 (N_9925,N_9627,N_9539);
and U9926 (N_9926,N_9573,N_9529);
xnor U9927 (N_9927,N_9649,N_9716);
xor U9928 (N_9928,N_9514,N_9569);
xor U9929 (N_9929,N_9580,N_9729);
or U9930 (N_9930,N_9515,N_9612);
and U9931 (N_9931,N_9624,N_9521);
xor U9932 (N_9932,N_9560,N_9743);
xnor U9933 (N_9933,N_9741,N_9746);
and U9934 (N_9934,N_9697,N_9664);
xnor U9935 (N_9935,N_9748,N_9630);
nand U9936 (N_9936,N_9695,N_9737);
and U9937 (N_9937,N_9623,N_9620);
and U9938 (N_9938,N_9736,N_9585);
and U9939 (N_9939,N_9596,N_9690);
and U9940 (N_9940,N_9688,N_9542);
nor U9941 (N_9941,N_9713,N_9600);
nand U9942 (N_9942,N_9630,N_9620);
xnor U9943 (N_9943,N_9605,N_9705);
nand U9944 (N_9944,N_9597,N_9686);
or U9945 (N_9945,N_9552,N_9664);
or U9946 (N_9946,N_9691,N_9612);
and U9947 (N_9947,N_9593,N_9503);
xnor U9948 (N_9948,N_9733,N_9746);
or U9949 (N_9949,N_9561,N_9694);
or U9950 (N_9950,N_9630,N_9549);
nor U9951 (N_9951,N_9641,N_9521);
or U9952 (N_9952,N_9728,N_9744);
or U9953 (N_9953,N_9747,N_9640);
nand U9954 (N_9954,N_9556,N_9674);
nand U9955 (N_9955,N_9628,N_9518);
or U9956 (N_9956,N_9570,N_9734);
and U9957 (N_9957,N_9747,N_9697);
and U9958 (N_9958,N_9531,N_9568);
or U9959 (N_9959,N_9574,N_9690);
or U9960 (N_9960,N_9625,N_9629);
nand U9961 (N_9961,N_9746,N_9711);
nand U9962 (N_9962,N_9743,N_9623);
or U9963 (N_9963,N_9628,N_9693);
and U9964 (N_9964,N_9549,N_9547);
nor U9965 (N_9965,N_9510,N_9564);
nor U9966 (N_9966,N_9561,N_9731);
or U9967 (N_9967,N_9514,N_9570);
nand U9968 (N_9968,N_9583,N_9599);
nor U9969 (N_9969,N_9733,N_9658);
xnor U9970 (N_9970,N_9683,N_9700);
or U9971 (N_9971,N_9625,N_9642);
nand U9972 (N_9972,N_9512,N_9534);
xor U9973 (N_9973,N_9613,N_9580);
and U9974 (N_9974,N_9597,N_9587);
nor U9975 (N_9975,N_9629,N_9736);
nand U9976 (N_9976,N_9604,N_9554);
or U9977 (N_9977,N_9522,N_9570);
nor U9978 (N_9978,N_9723,N_9713);
nand U9979 (N_9979,N_9585,N_9566);
and U9980 (N_9980,N_9704,N_9647);
xor U9981 (N_9981,N_9679,N_9562);
nand U9982 (N_9982,N_9604,N_9694);
nor U9983 (N_9983,N_9615,N_9589);
xor U9984 (N_9984,N_9699,N_9572);
or U9985 (N_9985,N_9657,N_9537);
xor U9986 (N_9986,N_9551,N_9556);
xnor U9987 (N_9987,N_9724,N_9671);
and U9988 (N_9988,N_9644,N_9503);
nand U9989 (N_9989,N_9524,N_9559);
nor U9990 (N_9990,N_9558,N_9530);
or U9991 (N_9991,N_9687,N_9523);
and U9992 (N_9992,N_9649,N_9603);
nand U9993 (N_9993,N_9525,N_9704);
or U9994 (N_9994,N_9651,N_9715);
xnor U9995 (N_9995,N_9671,N_9612);
xnor U9996 (N_9996,N_9659,N_9524);
nor U9997 (N_9997,N_9506,N_9735);
nor U9998 (N_9998,N_9587,N_9741);
and U9999 (N_9999,N_9632,N_9504);
xnor U10000 (N_10000,N_9836,N_9845);
or U10001 (N_10001,N_9877,N_9971);
xnor U10002 (N_10002,N_9761,N_9944);
nor U10003 (N_10003,N_9819,N_9928);
and U10004 (N_10004,N_9970,N_9922);
nor U10005 (N_10005,N_9856,N_9796);
nand U10006 (N_10006,N_9850,N_9778);
or U10007 (N_10007,N_9932,N_9783);
nor U10008 (N_10008,N_9875,N_9949);
or U10009 (N_10009,N_9827,N_9886);
or U10010 (N_10010,N_9948,N_9869);
nand U10011 (N_10011,N_9859,N_9938);
nand U10012 (N_10012,N_9941,N_9887);
and U10013 (N_10013,N_9864,N_9989);
xnor U10014 (N_10014,N_9773,N_9953);
or U10015 (N_10015,N_9884,N_9754);
xor U10016 (N_10016,N_9905,N_9935);
nor U10017 (N_10017,N_9772,N_9882);
or U10018 (N_10018,N_9914,N_9809);
and U10019 (N_10019,N_9865,N_9918);
and U10020 (N_10020,N_9911,N_9838);
nand U10021 (N_10021,N_9960,N_9867);
xnor U10022 (N_10022,N_9814,N_9893);
and U10023 (N_10023,N_9765,N_9832);
and U10024 (N_10024,N_9818,N_9753);
xor U10025 (N_10025,N_9876,N_9906);
xor U10026 (N_10026,N_9804,N_9786);
or U10027 (N_10027,N_9987,N_9752);
nor U10028 (N_10028,N_9966,N_9835);
or U10029 (N_10029,N_9931,N_9837);
and U10030 (N_10030,N_9985,N_9803);
or U10031 (N_10031,N_9756,N_9860);
nand U10032 (N_10032,N_9981,N_9942);
or U10033 (N_10033,N_9848,N_9828);
xnor U10034 (N_10034,N_9839,N_9947);
nand U10035 (N_10035,N_9961,N_9817);
xnor U10036 (N_10036,N_9833,N_9933);
nor U10037 (N_10037,N_9902,N_9924);
nand U10038 (N_10038,N_9993,N_9764);
or U10039 (N_10039,N_9842,N_9791);
nand U10040 (N_10040,N_9890,N_9991);
nand U10041 (N_10041,N_9849,N_9964);
or U10042 (N_10042,N_9959,N_9834);
or U10043 (N_10043,N_9811,N_9915);
or U10044 (N_10044,N_9852,N_9789);
xnor U10045 (N_10045,N_9760,N_9939);
nand U10046 (N_10046,N_9986,N_9896);
or U10047 (N_10047,N_9972,N_9984);
nand U10048 (N_10048,N_9978,N_9776);
and U10049 (N_10049,N_9841,N_9824);
and U10050 (N_10050,N_9908,N_9990);
nand U10051 (N_10051,N_9956,N_9815);
or U10052 (N_10052,N_9821,N_9775);
or U10053 (N_10053,N_9912,N_9995);
nand U10054 (N_10054,N_9976,N_9847);
and U10055 (N_10055,N_9957,N_9855);
xor U10056 (N_10056,N_9943,N_9913);
nor U10057 (N_10057,N_9806,N_9802);
nor U10058 (N_10058,N_9983,N_9897);
xnor U10059 (N_10059,N_9927,N_9858);
nand U10060 (N_10060,N_9881,N_9872);
nor U10061 (N_10061,N_9784,N_9785);
xnor U10062 (N_10062,N_9951,N_9862);
nor U10063 (N_10063,N_9854,N_9917);
xor U10064 (N_10064,N_9759,N_9926);
nand U10065 (N_10065,N_9788,N_9808);
xor U10066 (N_10066,N_9916,N_9816);
nand U10067 (N_10067,N_9929,N_9979);
nor U10068 (N_10068,N_9930,N_9768);
or U10069 (N_10069,N_9880,N_9940);
and U10070 (N_10070,N_9946,N_9812);
nand U10071 (N_10071,N_9750,N_9988);
xnor U10072 (N_10072,N_9919,N_9781);
and U10073 (N_10073,N_9969,N_9873);
or U10074 (N_10074,N_9888,N_9868);
nand U10075 (N_10075,N_9843,N_9771);
and U10076 (N_10076,N_9861,N_9779);
xnor U10077 (N_10077,N_9883,N_9997);
xnor U10078 (N_10078,N_9777,N_9826);
xor U10079 (N_10079,N_9851,N_9829);
nor U10080 (N_10080,N_9844,N_9879);
nor U10081 (N_10081,N_9797,N_9800);
nand U10082 (N_10082,N_9770,N_9866);
or U10083 (N_10083,N_9782,N_9977);
xnor U10084 (N_10084,N_9921,N_9822);
nor U10085 (N_10085,N_9954,N_9900);
xor U10086 (N_10086,N_9758,N_9965);
or U10087 (N_10087,N_9945,N_9901);
and U10088 (N_10088,N_9810,N_9885);
and U10089 (N_10089,N_9793,N_9767);
xnor U10090 (N_10090,N_9952,N_9955);
nand U10091 (N_10091,N_9975,N_9936);
xnor U10092 (N_10092,N_9820,N_9813);
nor U10093 (N_10093,N_9967,N_9958);
or U10094 (N_10094,N_9909,N_9973);
or U10095 (N_10095,N_9968,N_9755);
or U10096 (N_10096,N_9787,N_9762);
xnor U10097 (N_10097,N_9874,N_9889);
or U10098 (N_10098,N_9980,N_9853);
xnor U10099 (N_10099,N_9892,N_9891);
xnor U10100 (N_10100,N_9907,N_9790);
or U10101 (N_10101,N_9823,N_9805);
or U10102 (N_10102,N_9934,N_9903);
and U10103 (N_10103,N_9825,N_9925);
or U10104 (N_10104,N_9794,N_9831);
or U10105 (N_10105,N_9992,N_9780);
xor U10106 (N_10106,N_9795,N_9996);
xor U10107 (N_10107,N_9910,N_9870);
nor U10108 (N_10108,N_9863,N_9766);
nor U10109 (N_10109,N_9757,N_9871);
and U10110 (N_10110,N_9798,N_9963);
nor U10111 (N_10111,N_9998,N_9792);
and U10112 (N_10112,N_9878,N_9763);
nor U10113 (N_10113,N_9807,N_9846);
or U10114 (N_10114,N_9898,N_9840);
nand U10115 (N_10115,N_9751,N_9937);
nor U10116 (N_10116,N_9923,N_9857);
and U10117 (N_10117,N_9904,N_9994);
nor U10118 (N_10118,N_9801,N_9974);
nor U10119 (N_10119,N_9982,N_9962);
and U10120 (N_10120,N_9774,N_9920);
or U10121 (N_10121,N_9899,N_9999);
xor U10122 (N_10122,N_9895,N_9894);
nor U10123 (N_10123,N_9950,N_9799);
and U10124 (N_10124,N_9830,N_9769);
nand U10125 (N_10125,N_9834,N_9782);
xor U10126 (N_10126,N_9829,N_9884);
or U10127 (N_10127,N_9951,N_9874);
nand U10128 (N_10128,N_9951,N_9842);
and U10129 (N_10129,N_9787,N_9750);
xnor U10130 (N_10130,N_9840,N_9917);
and U10131 (N_10131,N_9842,N_9967);
and U10132 (N_10132,N_9816,N_9833);
or U10133 (N_10133,N_9976,N_9817);
and U10134 (N_10134,N_9794,N_9773);
and U10135 (N_10135,N_9803,N_9864);
nor U10136 (N_10136,N_9982,N_9994);
xnor U10137 (N_10137,N_9775,N_9892);
nor U10138 (N_10138,N_9840,N_9786);
or U10139 (N_10139,N_9786,N_9869);
xnor U10140 (N_10140,N_9831,N_9790);
nor U10141 (N_10141,N_9970,N_9895);
or U10142 (N_10142,N_9931,N_9874);
nand U10143 (N_10143,N_9820,N_9970);
nor U10144 (N_10144,N_9934,N_9864);
nand U10145 (N_10145,N_9945,N_9834);
and U10146 (N_10146,N_9804,N_9761);
nor U10147 (N_10147,N_9833,N_9786);
nor U10148 (N_10148,N_9922,N_9763);
nor U10149 (N_10149,N_9873,N_9811);
or U10150 (N_10150,N_9753,N_9930);
and U10151 (N_10151,N_9967,N_9872);
xnor U10152 (N_10152,N_9799,N_9856);
or U10153 (N_10153,N_9927,N_9811);
xor U10154 (N_10154,N_9958,N_9981);
nor U10155 (N_10155,N_9998,N_9751);
or U10156 (N_10156,N_9860,N_9833);
or U10157 (N_10157,N_9863,N_9751);
nand U10158 (N_10158,N_9848,N_9893);
nor U10159 (N_10159,N_9855,N_9883);
or U10160 (N_10160,N_9872,N_9950);
nor U10161 (N_10161,N_9996,N_9768);
and U10162 (N_10162,N_9784,N_9757);
nor U10163 (N_10163,N_9966,N_9801);
and U10164 (N_10164,N_9973,N_9925);
and U10165 (N_10165,N_9928,N_9861);
nor U10166 (N_10166,N_9800,N_9838);
nand U10167 (N_10167,N_9878,N_9998);
nor U10168 (N_10168,N_9943,N_9952);
or U10169 (N_10169,N_9797,N_9999);
and U10170 (N_10170,N_9841,N_9913);
xnor U10171 (N_10171,N_9978,N_9816);
nand U10172 (N_10172,N_9945,N_9951);
nor U10173 (N_10173,N_9927,N_9827);
and U10174 (N_10174,N_9849,N_9850);
nand U10175 (N_10175,N_9804,N_9933);
and U10176 (N_10176,N_9835,N_9928);
and U10177 (N_10177,N_9886,N_9980);
and U10178 (N_10178,N_9750,N_9880);
nor U10179 (N_10179,N_9928,N_9896);
or U10180 (N_10180,N_9807,N_9905);
or U10181 (N_10181,N_9828,N_9787);
xor U10182 (N_10182,N_9829,N_9899);
or U10183 (N_10183,N_9923,N_9906);
xor U10184 (N_10184,N_9964,N_9869);
or U10185 (N_10185,N_9805,N_9957);
nor U10186 (N_10186,N_9880,N_9885);
xor U10187 (N_10187,N_9950,N_9909);
xnor U10188 (N_10188,N_9903,N_9866);
nand U10189 (N_10189,N_9835,N_9880);
nor U10190 (N_10190,N_9930,N_9794);
nand U10191 (N_10191,N_9987,N_9779);
xnor U10192 (N_10192,N_9808,N_9917);
and U10193 (N_10193,N_9797,N_9994);
xor U10194 (N_10194,N_9960,N_9791);
and U10195 (N_10195,N_9866,N_9768);
xor U10196 (N_10196,N_9981,N_9882);
nand U10197 (N_10197,N_9786,N_9816);
xor U10198 (N_10198,N_9906,N_9825);
xor U10199 (N_10199,N_9915,N_9819);
or U10200 (N_10200,N_9776,N_9809);
nor U10201 (N_10201,N_9815,N_9996);
nand U10202 (N_10202,N_9824,N_9901);
or U10203 (N_10203,N_9931,N_9911);
and U10204 (N_10204,N_9981,N_9969);
or U10205 (N_10205,N_9942,N_9837);
nor U10206 (N_10206,N_9958,N_9872);
nand U10207 (N_10207,N_9771,N_9874);
or U10208 (N_10208,N_9781,N_9783);
xor U10209 (N_10209,N_9830,N_9798);
nand U10210 (N_10210,N_9957,N_9822);
xor U10211 (N_10211,N_9952,N_9858);
nand U10212 (N_10212,N_9813,N_9988);
nor U10213 (N_10213,N_9989,N_9792);
nor U10214 (N_10214,N_9808,N_9850);
xor U10215 (N_10215,N_9858,N_9959);
and U10216 (N_10216,N_9940,N_9852);
or U10217 (N_10217,N_9931,N_9838);
and U10218 (N_10218,N_9890,N_9827);
or U10219 (N_10219,N_9827,N_9968);
or U10220 (N_10220,N_9935,N_9944);
xor U10221 (N_10221,N_9916,N_9774);
and U10222 (N_10222,N_9808,N_9928);
nand U10223 (N_10223,N_9862,N_9970);
nor U10224 (N_10224,N_9782,N_9807);
and U10225 (N_10225,N_9890,N_9983);
and U10226 (N_10226,N_9923,N_9780);
or U10227 (N_10227,N_9868,N_9988);
and U10228 (N_10228,N_9765,N_9938);
and U10229 (N_10229,N_9771,N_9968);
xnor U10230 (N_10230,N_9810,N_9850);
nor U10231 (N_10231,N_9968,N_9759);
and U10232 (N_10232,N_9959,N_9828);
or U10233 (N_10233,N_9947,N_9967);
nor U10234 (N_10234,N_9993,N_9881);
nor U10235 (N_10235,N_9826,N_9864);
and U10236 (N_10236,N_9894,N_9767);
xnor U10237 (N_10237,N_9800,N_9774);
xnor U10238 (N_10238,N_9966,N_9980);
and U10239 (N_10239,N_9923,N_9896);
nor U10240 (N_10240,N_9785,N_9968);
xnor U10241 (N_10241,N_9968,N_9940);
nand U10242 (N_10242,N_9998,N_9905);
nand U10243 (N_10243,N_9976,N_9887);
nor U10244 (N_10244,N_9831,N_9784);
nand U10245 (N_10245,N_9858,N_9972);
nor U10246 (N_10246,N_9853,N_9784);
and U10247 (N_10247,N_9762,N_9911);
or U10248 (N_10248,N_9862,N_9867);
xnor U10249 (N_10249,N_9954,N_9770);
or U10250 (N_10250,N_10119,N_10238);
nor U10251 (N_10251,N_10089,N_10039);
or U10252 (N_10252,N_10033,N_10035);
nand U10253 (N_10253,N_10164,N_10014);
xor U10254 (N_10254,N_10012,N_10210);
nor U10255 (N_10255,N_10122,N_10180);
nor U10256 (N_10256,N_10112,N_10222);
or U10257 (N_10257,N_10129,N_10233);
nor U10258 (N_10258,N_10199,N_10030);
xor U10259 (N_10259,N_10105,N_10026);
nor U10260 (N_10260,N_10150,N_10141);
and U10261 (N_10261,N_10184,N_10193);
nand U10262 (N_10262,N_10246,N_10192);
xnor U10263 (N_10263,N_10103,N_10011);
or U10264 (N_10264,N_10007,N_10023);
xor U10265 (N_10265,N_10024,N_10102);
and U10266 (N_10266,N_10231,N_10044);
and U10267 (N_10267,N_10097,N_10005);
nor U10268 (N_10268,N_10076,N_10226);
and U10269 (N_10269,N_10168,N_10043);
and U10270 (N_10270,N_10050,N_10128);
nand U10271 (N_10271,N_10019,N_10195);
xnor U10272 (N_10272,N_10191,N_10104);
and U10273 (N_10273,N_10142,N_10127);
xor U10274 (N_10274,N_10126,N_10092);
nor U10275 (N_10275,N_10240,N_10037);
or U10276 (N_10276,N_10090,N_10158);
nand U10277 (N_10277,N_10218,N_10178);
nor U10278 (N_10278,N_10159,N_10230);
xnor U10279 (N_10279,N_10197,N_10063);
xor U10280 (N_10280,N_10227,N_10049);
nand U10281 (N_10281,N_10149,N_10068);
xnor U10282 (N_10282,N_10207,N_10031);
or U10283 (N_10283,N_10036,N_10046);
nor U10284 (N_10284,N_10066,N_10243);
nand U10285 (N_10285,N_10027,N_10125);
nor U10286 (N_10286,N_10048,N_10110);
nand U10287 (N_10287,N_10151,N_10144);
and U10288 (N_10288,N_10054,N_10091);
xor U10289 (N_10289,N_10139,N_10235);
nand U10290 (N_10290,N_10202,N_10015);
nor U10291 (N_10291,N_10166,N_10176);
nand U10292 (N_10292,N_10213,N_10081);
or U10293 (N_10293,N_10000,N_10003);
nor U10294 (N_10294,N_10200,N_10209);
and U10295 (N_10295,N_10140,N_10008);
xor U10296 (N_10296,N_10154,N_10071);
or U10297 (N_10297,N_10157,N_10225);
or U10298 (N_10298,N_10229,N_10211);
nand U10299 (N_10299,N_10188,N_10002);
or U10300 (N_10300,N_10244,N_10228);
and U10301 (N_10301,N_10161,N_10069);
nor U10302 (N_10302,N_10173,N_10083);
nor U10303 (N_10303,N_10143,N_10094);
nor U10304 (N_10304,N_10196,N_10101);
xor U10305 (N_10305,N_10237,N_10130);
and U10306 (N_10306,N_10169,N_10025);
or U10307 (N_10307,N_10241,N_10187);
nand U10308 (N_10308,N_10223,N_10152);
or U10309 (N_10309,N_10185,N_10113);
and U10310 (N_10310,N_10118,N_10174);
nor U10311 (N_10311,N_10239,N_10167);
or U10312 (N_10312,N_10057,N_10045);
nand U10313 (N_10313,N_10136,N_10131);
and U10314 (N_10314,N_10108,N_10189);
nor U10315 (N_10315,N_10114,N_10029);
or U10316 (N_10316,N_10182,N_10034);
nor U10317 (N_10317,N_10038,N_10117);
xnor U10318 (N_10318,N_10165,N_10042);
nor U10319 (N_10319,N_10206,N_10100);
or U10320 (N_10320,N_10056,N_10121);
nor U10321 (N_10321,N_10067,N_10055);
or U10322 (N_10322,N_10082,N_10053);
or U10323 (N_10323,N_10093,N_10147);
or U10324 (N_10324,N_10016,N_10132);
xnor U10325 (N_10325,N_10160,N_10249);
and U10326 (N_10326,N_10217,N_10059);
nand U10327 (N_10327,N_10021,N_10006);
or U10328 (N_10328,N_10107,N_10018);
nand U10329 (N_10329,N_10133,N_10074);
and U10330 (N_10330,N_10201,N_10077);
xnor U10331 (N_10331,N_10020,N_10181);
nand U10332 (N_10332,N_10153,N_10220);
or U10333 (N_10333,N_10017,N_10064);
xor U10334 (N_10334,N_10216,N_10028);
xnor U10335 (N_10335,N_10096,N_10203);
or U10336 (N_10336,N_10099,N_10177);
or U10337 (N_10337,N_10145,N_10080);
and U10338 (N_10338,N_10086,N_10009);
or U10339 (N_10339,N_10179,N_10190);
nand U10340 (N_10340,N_10098,N_10170);
or U10341 (N_10341,N_10032,N_10175);
xor U10342 (N_10342,N_10022,N_10214);
and U10343 (N_10343,N_10058,N_10224);
nor U10344 (N_10344,N_10109,N_10115);
nand U10345 (N_10345,N_10065,N_10242);
and U10346 (N_10346,N_10010,N_10052);
nand U10347 (N_10347,N_10212,N_10156);
nand U10348 (N_10348,N_10004,N_10137);
nor U10349 (N_10349,N_10116,N_10062);
xnor U10350 (N_10350,N_10051,N_10236);
nand U10351 (N_10351,N_10248,N_10111);
or U10352 (N_10352,N_10186,N_10106);
nand U10353 (N_10353,N_10155,N_10204);
nand U10354 (N_10354,N_10001,N_10171);
nor U10355 (N_10355,N_10061,N_10084);
xor U10356 (N_10356,N_10194,N_10162);
xnor U10357 (N_10357,N_10040,N_10060);
nand U10358 (N_10358,N_10087,N_10124);
or U10359 (N_10359,N_10148,N_10123);
nor U10360 (N_10360,N_10138,N_10013);
or U10361 (N_10361,N_10219,N_10234);
or U10362 (N_10362,N_10073,N_10135);
nand U10363 (N_10363,N_10075,N_10163);
and U10364 (N_10364,N_10247,N_10120);
nand U10365 (N_10365,N_10208,N_10221);
and U10366 (N_10366,N_10205,N_10041);
nand U10367 (N_10367,N_10172,N_10245);
nand U10368 (N_10368,N_10095,N_10085);
xnor U10369 (N_10369,N_10078,N_10183);
nand U10370 (N_10370,N_10047,N_10134);
nor U10371 (N_10371,N_10072,N_10070);
xnor U10372 (N_10372,N_10215,N_10198);
xnor U10373 (N_10373,N_10146,N_10088);
and U10374 (N_10374,N_10232,N_10079);
or U10375 (N_10375,N_10159,N_10083);
and U10376 (N_10376,N_10000,N_10042);
xor U10377 (N_10377,N_10030,N_10076);
and U10378 (N_10378,N_10192,N_10078);
nor U10379 (N_10379,N_10148,N_10186);
nor U10380 (N_10380,N_10072,N_10218);
nor U10381 (N_10381,N_10128,N_10184);
and U10382 (N_10382,N_10073,N_10208);
xor U10383 (N_10383,N_10194,N_10141);
nand U10384 (N_10384,N_10154,N_10183);
nor U10385 (N_10385,N_10062,N_10240);
nand U10386 (N_10386,N_10133,N_10045);
xor U10387 (N_10387,N_10157,N_10226);
xor U10388 (N_10388,N_10229,N_10214);
nor U10389 (N_10389,N_10175,N_10036);
nand U10390 (N_10390,N_10159,N_10105);
nor U10391 (N_10391,N_10183,N_10142);
nor U10392 (N_10392,N_10004,N_10094);
xor U10393 (N_10393,N_10029,N_10061);
nand U10394 (N_10394,N_10228,N_10167);
nor U10395 (N_10395,N_10097,N_10246);
and U10396 (N_10396,N_10108,N_10226);
xnor U10397 (N_10397,N_10084,N_10013);
or U10398 (N_10398,N_10085,N_10144);
xnor U10399 (N_10399,N_10119,N_10077);
xnor U10400 (N_10400,N_10028,N_10163);
or U10401 (N_10401,N_10249,N_10010);
nor U10402 (N_10402,N_10180,N_10205);
nand U10403 (N_10403,N_10166,N_10128);
xnor U10404 (N_10404,N_10082,N_10139);
xor U10405 (N_10405,N_10001,N_10135);
xnor U10406 (N_10406,N_10022,N_10137);
nor U10407 (N_10407,N_10021,N_10187);
nand U10408 (N_10408,N_10143,N_10128);
or U10409 (N_10409,N_10229,N_10245);
nand U10410 (N_10410,N_10069,N_10098);
nand U10411 (N_10411,N_10178,N_10012);
nor U10412 (N_10412,N_10091,N_10163);
xor U10413 (N_10413,N_10021,N_10126);
nor U10414 (N_10414,N_10244,N_10102);
nor U10415 (N_10415,N_10172,N_10066);
xor U10416 (N_10416,N_10100,N_10013);
or U10417 (N_10417,N_10223,N_10076);
nand U10418 (N_10418,N_10238,N_10163);
or U10419 (N_10419,N_10129,N_10075);
and U10420 (N_10420,N_10006,N_10022);
nand U10421 (N_10421,N_10021,N_10110);
nor U10422 (N_10422,N_10015,N_10108);
xnor U10423 (N_10423,N_10163,N_10207);
xor U10424 (N_10424,N_10219,N_10031);
and U10425 (N_10425,N_10142,N_10137);
nand U10426 (N_10426,N_10137,N_10051);
and U10427 (N_10427,N_10047,N_10079);
and U10428 (N_10428,N_10133,N_10090);
nor U10429 (N_10429,N_10155,N_10244);
or U10430 (N_10430,N_10235,N_10126);
or U10431 (N_10431,N_10144,N_10136);
and U10432 (N_10432,N_10244,N_10048);
or U10433 (N_10433,N_10247,N_10152);
nor U10434 (N_10434,N_10121,N_10172);
xor U10435 (N_10435,N_10153,N_10156);
xnor U10436 (N_10436,N_10126,N_10091);
and U10437 (N_10437,N_10218,N_10157);
or U10438 (N_10438,N_10002,N_10167);
xor U10439 (N_10439,N_10094,N_10072);
and U10440 (N_10440,N_10053,N_10116);
nand U10441 (N_10441,N_10162,N_10204);
or U10442 (N_10442,N_10127,N_10077);
nand U10443 (N_10443,N_10177,N_10073);
or U10444 (N_10444,N_10012,N_10246);
nand U10445 (N_10445,N_10006,N_10030);
or U10446 (N_10446,N_10088,N_10140);
nor U10447 (N_10447,N_10221,N_10210);
xnor U10448 (N_10448,N_10130,N_10052);
nand U10449 (N_10449,N_10155,N_10225);
nor U10450 (N_10450,N_10094,N_10024);
or U10451 (N_10451,N_10117,N_10051);
nor U10452 (N_10452,N_10147,N_10242);
xnor U10453 (N_10453,N_10001,N_10158);
and U10454 (N_10454,N_10217,N_10098);
xnor U10455 (N_10455,N_10174,N_10247);
or U10456 (N_10456,N_10246,N_10093);
nand U10457 (N_10457,N_10077,N_10166);
and U10458 (N_10458,N_10224,N_10025);
nor U10459 (N_10459,N_10114,N_10107);
nor U10460 (N_10460,N_10081,N_10238);
and U10461 (N_10461,N_10025,N_10248);
nor U10462 (N_10462,N_10098,N_10115);
xor U10463 (N_10463,N_10120,N_10072);
nand U10464 (N_10464,N_10085,N_10159);
xnor U10465 (N_10465,N_10128,N_10015);
xor U10466 (N_10466,N_10202,N_10128);
and U10467 (N_10467,N_10245,N_10169);
and U10468 (N_10468,N_10239,N_10100);
and U10469 (N_10469,N_10128,N_10162);
and U10470 (N_10470,N_10194,N_10150);
xnor U10471 (N_10471,N_10000,N_10080);
or U10472 (N_10472,N_10179,N_10108);
nor U10473 (N_10473,N_10050,N_10138);
xor U10474 (N_10474,N_10173,N_10248);
xor U10475 (N_10475,N_10225,N_10084);
nand U10476 (N_10476,N_10174,N_10170);
and U10477 (N_10477,N_10049,N_10044);
nand U10478 (N_10478,N_10001,N_10187);
or U10479 (N_10479,N_10194,N_10221);
and U10480 (N_10480,N_10017,N_10001);
nor U10481 (N_10481,N_10207,N_10013);
or U10482 (N_10482,N_10198,N_10021);
and U10483 (N_10483,N_10211,N_10223);
xor U10484 (N_10484,N_10005,N_10015);
and U10485 (N_10485,N_10123,N_10043);
nor U10486 (N_10486,N_10232,N_10049);
nor U10487 (N_10487,N_10042,N_10058);
nor U10488 (N_10488,N_10156,N_10118);
nor U10489 (N_10489,N_10103,N_10143);
or U10490 (N_10490,N_10034,N_10147);
nor U10491 (N_10491,N_10195,N_10229);
nand U10492 (N_10492,N_10098,N_10022);
nor U10493 (N_10493,N_10023,N_10238);
xor U10494 (N_10494,N_10146,N_10046);
and U10495 (N_10495,N_10008,N_10156);
nor U10496 (N_10496,N_10029,N_10062);
or U10497 (N_10497,N_10142,N_10201);
and U10498 (N_10498,N_10018,N_10166);
or U10499 (N_10499,N_10232,N_10186);
xnor U10500 (N_10500,N_10485,N_10464);
nand U10501 (N_10501,N_10286,N_10459);
or U10502 (N_10502,N_10265,N_10343);
xor U10503 (N_10503,N_10480,N_10405);
nand U10504 (N_10504,N_10386,N_10489);
and U10505 (N_10505,N_10374,N_10388);
or U10506 (N_10506,N_10360,N_10441);
or U10507 (N_10507,N_10442,N_10373);
xor U10508 (N_10508,N_10400,N_10425);
nor U10509 (N_10509,N_10288,N_10380);
or U10510 (N_10510,N_10298,N_10364);
or U10511 (N_10511,N_10435,N_10498);
and U10512 (N_10512,N_10267,N_10289);
nor U10513 (N_10513,N_10352,N_10372);
and U10514 (N_10514,N_10421,N_10273);
and U10515 (N_10515,N_10275,N_10439);
or U10516 (N_10516,N_10402,N_10471);
nand U10517 (N_10517,N_10350,N_10440);
and U10518 (N_10518,N_10340,N_10292);
nand U10519 (N_10519,N_10357,N_10495);
or U10520 (N_10520,N_10366,N_10406);
or U10521 (N_10521,N_10328,N_10318);
nor U10522 (N_10522,N_10469,N_10294);
nand U10523 (N_10523,N_10314,N_10279);
and U10524 (N_10524,N_10304,N_10346);
nand U10525 (N_10525,N_10334,N_10377);
nand U10526 (N_10526,N_10444,N_10413);
nor U10527 (N_10527,N_10256,N_10278);
xor U10528 (N_10528,N_10303,N_10270);
xnor U10529 (N_10529,N_10394,N_10453);
or U10530 (N_10530,N_10407,N_10452);
nand U10531 (N_10531,N_10282,N_10390);
and U10532 (N_10532,N_10269,N_10454);
and U10533 (N_10533,N_10306,N_10271);
xnor U10534 (N_10534,N_10255,N_10482);
xor U10535 (N_10535,N_10478,N_10359);
or U10536 (N_10536,N_10320,N_10381);
or U10537 (N_10537,N_10285,N_10477);
nor U10538 (N_10538,N_10443,N_10397);
or U10539 (N_10539,N_10266,N_10410);
or U10540 (N_10540,N_10347,N_10497);
nand U10541 (N_10541,N_10446,N_10492);
nor U10542 (N_10542,N_10378,N_10327);
xor U10543 (N_10543,N_10414,N_10335);
nor U10544 (N_10544,N_10309,N_10369);
or U10545 (N_10545,N_10488,N_10371);
nand U10546 (N_10546,N_10300,N_10392);
xor U10547 (N_10547,N_10457,N_10451);
xor U10548 (N_10548,N_10398,N_10305);
nand U10549 (N_10549,N_10365,N_10447);
xnor U10550 (N_10550,N_10481,N_10445);
and U10551 (N_10551,N_10431,N_10434);
or U10552 (N_10552,N_10436,N_10367);
xnor U10553 (N_10553,N_10412,N_10496);
xnor U10554 (N_10554,N_10424,N_10486);
xnor U10555 (N_10555,N_10264,N_10428);
and U10556 (N_10556,N_10301,N_10297);
or U10557 (N_10557,N_10409,N_10349);
nor U10558 (N_10558,N_10323,N_10472);
nand U10559 (N_10559,N_10423,N_10322);
nand U10560 (N_10560,N_10411,N_10448);
or U10561 (N_10561,N_10391,N_10355);
nor U10562 (N_10562,N_10313,N_10375);
or U10563 (N_10563,N_10430,N_10468);
nor U10564 (N_10564,N_10491,N_10465);
and U10565 (N_10565,N_10475,N_10499);
and U10566 (N_10566,N_10467,N_10438);
nor U10567 (N_10567,N_10476,N_10330);
nor U10568 (N_10568,N_10437,N_10268);
and U10569 (N_10569,N_10283,N_10383);
and U10570 (N_10570,N_10401,N_10474);
xor U10571 (N_10571,N_10325,N_10393);
nand U10572 (N_10572,N_10348,N_10466);
and U10573 (N_10573,N_10337,N_10455);
nor U10574 (N_10574,N_10420,N_10396);
nand U10575 (N_10575,N_10356,N_10295);
nand U10576 (N_10576,N_10338,N_10293);
and U10577 (N_10577,N_10362,N_10417);
or U10578 (N_10578,N_10326,N_10370);
or U10579 (N_10579,N_10274,N_10311);
nor U10580 (N_10580,N_10291,N_10277);
nand U10581 (N_10581,N_10345,N_10422);
nor U10582 (N_10582,N_10252,N_10382);
xnor U10583 (N_10583,N_10399,N_10351);
and U10584 (N_10584,N_10333,N_10368);
nand U10585 (N_10585,N_10259,N_10361);
and U10586 (N_10586,N_10262,N_10254);
nor U10587 (N_10587,N_10312,N_10354);
or U10588 (N_10588,N_10342,N_10456);
xnor U10589 (N_10589,N_10258,N_10329);
nor U10590 (N_10590,N_10257,N_10379);
xnor U10591 (N_10591,N_10403,N_10324);
or U10592 (N_10592,N_10263,N_10331);
nand U10593 (N_10593,N_10299,N_10260);
nor U10594 (N_10594,N_10363,N_10415);
nor U10595 (N_10595,N_10308,N_10416);
nand U10596 (N_10596,N_10408,N_10404);
nand U10597 (N_10597,N_10461,N_10449);
or U10598 (N_10598,N_10460,N_10272);
nand U10599 (N_10599,N_10358,N_10332);
or U10600 (N_10600,N_10494,N_10302);
and U10601 (N_10601,N_10384,N_10321);
xnor U10602 (N_10602,N_10389,N_10316);
and U10603 (N_10603,N_10341,N_10353);
or U10604 (N_10604,N_10261,N_10419);
xor U10605 (N_10605,N_10250,N_10296);
or U10606 (N_10606,N_10470,N_10310);
nor U10607 (N_10607,N_10287,N_10387);
nor U10608 (N_10608,N_10493,N_10385);
xnor U10609 (N_10609,N_10251,N_10376);
nand U10610 (N_10610,N_10479,N_10315);
or U10611 (N_10611,N_10433,N_10450);
nand U10612 (N_10612,N_10281,N_10462);
xor U10613 (N_10613,N_10473,N_10426);
nand U10614 (N_10614,N_10490,N_10484);
nand U10615 (N_10615,N_10458,N_10336);
nor U10616 (N_10616,N_10280,N_10317);
and U10617 (N_10617,N_10429,N_10344);
nor U10618 (N_10618,N_10339,N_10487);
and U10619 (N_10619,N_10253,N_10276);
nor U10620 (N_10620,N_10418,N_10290);
or U10621 (N_10621,N_10432,N_10427);
nor U10622 (N_10622,N_10319,N_10284);
or U10623 (N_10623,N_10483,N_10307);
and U10624 (N_10624,N_10395,N_10463);
nand U10625 (N_10625,N_10439,N_10448);
and U10626 (N_10626,N_10324,N_10363);
xor U10627 (N_10627,N_10386,N_10405);
or U10628 (N_10628,N_10340,N_10492);
and U10629 (N_10629,N_10426,N_10388);
nor U10630 (N_10630,N_10416,N_10476);
nand U10631 (N_10631,N_10380,N_10481);
and U10632 (N_10632,N_10324,N_10388);
nor U10633 (N_10633,N_10295,N_10487);
xnor U10634 (N_10634,N_10484,N_10274);
or U10635 (N_10635,N_10443,N_10411);
xor U10636 (N_10636,N_10333,N_10388);
and U10637 (N_10637,N_10380,N_10366);
and U10638 (N_10638,N_10283,N_10298);
nand U10639 (N_10639,N_10280,N_10394);
xnor U10640 (N_10640,N_10272,N_10353);
and U10641 (N_10641,N_10396,N_10435);
nor U10642 (N_10642,N_10267,N_10407);
and U10643 (N_10643,N_10305,N_10292);
or U10644 (N_10644,N_10452,N_10325);
and U10645 (N_10645,N_10479,N_10355);
nor U10646 (N_10646,N_10310,N_10392);
and U10647 (N_10647,N_10474,N_10302);
or U10648 (N_10648,N_10473,N_10453);
nor U10649 (N_10649,N_10417,N_10332);
nor U10650 (N_10650,N_10383,N_10397);
or U10651 (N_10651,N_10370,N_10389);
nor U10652 (N_10652,N_10284,N_10466);
and U10653 (N_10653,N_10327,N_10370);
xnor U10654 (N_10654,N_10360,N_10494);
nor U10655 (N_10655,N_10469,N_10263);
or U10656 (N_10656,N_10493,N_10305);
xor U10657 (N_10657,N_10488,N_10260);
or U10658 (N_10658,N_10464,N_10459);
and U10659 (N_10659,N_10432,N_10447);
and U10660 (N_10660,N_10351,N_10474);
or U10661 (N_10661,N_10470,N_10456);
nand U10662 (N_10662,N_10389,N_10323);
nor U10663 (N_10663,N_10437,N_10339);
nand U10664 (N_10664,N_10332,N_10439);
and U10665 (N_10665,N_10353,N_10261);
xnor U10666 (N_10666,N_10470,N_10381);
or U10667 (N_10667,N_10427,N_10480);
and U10668 (N_10668,N_10316,N_10328);
and U10669 (N_10669,N_10410,N_10480);
nand U10670 (N_10670,N_10275,N_10310);
xor U10671 (N_10671,N_10304,N_10366);
xnor U10672 (N_10672,N_10363,N_10399);
and U10673 (N_10673,N_10351,N_10419);
nor U10674 (N_10674,N_10379,N_10316);
nor U10675 (N_10675,N_10472,N_10308);
xor U10676 (N_10676,N_10454,N_10367);
or U10677 (N_10677,N_10386,N_10406);
or U10678 (N_10678,N_10487,N_10278);
and U10679 (N_10679,N_10295,N_10283);
or U10680 (N_10680,N_10435,N_10261);
nor U10681 (N_10681,N_10491,N_10255);
nand U10682 (N_10682,N_10466,N_10495);
xor U10683 (N_10683,N_10376,N_10321);
and U10684 (N_10684,N_10351,N_10477);
and U10685 (N_10685,N_10491,N_10454);
nand U10686 (N_10686,N_10486,N_10392);
nor U10687 (N_10687,N_10429,N_10372);
xnor U10688 (N_10688,N_10345,N_10352);
xnor U10689 (N_10689,N_10478,N_10270);
and U10690 (N_10690,N_10430,N_10263);
xnor U10691 (N_10691,N_10408,N_10290);
xor U10692 (N_10692,N_10255,N_10454);
xnor U10693 (N_10693,N_10465,N_10357);
or U10694 (N_10694,N_10400,N_10443);
or U10695 (N_10695,N_10331,N_10446);
xnor U10696 (N_10696,N_10335,N_10293);
nor U10697 (N_10697,N_10421,N_10349);
nor U10698 (N_10698,N_10371,N_10393);
xnor U10699 (N_10699,N_10457,N_10354);
and U10700 (N_10700,N_10465,N_10395);
nand U10701 (N_10701,N_10306,N_10274);
nor U10702 (N_10702,N_10321,N_10437);
and U10703 (N_10703,N_10317,N_10476);
or U10704 (N_10704,N_10350,N_10327);
xor U10705 (N_10705,N_10446,N_10286);
nor U10706 (N_10706,N_10307,N_10411);
nand U10707 (N_10707,N_10344,N_10321);
xnor U10708 (N_10708,N_10396,N_10393);
nor U10709 (N_10709,N_10424,N_10370);
nor U10710 (N_10710,N_10464,N_10359);
nand U10711 (N_10711,N_10417,N_10271);
or U10712 (N_10712,N_10491,N_10272);
xor U10713 (N_10713,N_10453,N_10387);
and U10714 (N_10714,N_10281,N_10385);
nor U10715 (N_10715,N_10303,N_10275);
or U10716 (N_10716,N_10430,N_10402);
nand U10717 (N_10717,N_10362,N_10496);
or U10718 (N_10718,N_10366,N_10375);
nand U10719 (N_10719,N_10334,N_10308);
and U10720 (N_10720,N_10352,N_10458);
nor U10721 (N_10721,N_10487,N_10478);
nor U10722 (N_10722,N_10457,N_10455);
xnor U10723 (N_10723,N_10274,N_10296);
nand U10724 (N_10724,N_10353,N_10356);
and U10725 (N_10725,N_10308,N_10420);
and U10726 (N_10726,N_10327,N_10402);
xor U10727 (N_10727,N_10402,N_10409);
or U10728 (N_10728,N_10353,N_10304);
xor U10729 (N_10729,N_10448,N_10404);
nand U10730 (N_10730,N_10384,N_10256);
or U10731 (N_10731,N_10353,N_10312);
nor U10732 (N_10732,N_10322,N_10281);
nand U10733 (N_10733,N_10307,N_10298);
nor U10734 (N_10734,N_10285,N_10499);
nor U10735 (N_10735,N_10301,N_10497);
nor U10736 (N_10736,N_10281,N_10356);
and U10737 (N_10737,N_10363,N_10266);
nor U10738 (N_10738,N_10425,N_10378);
nand U10739 (N_10739,N_10332,N_10260);
nor U10740 (N_10740,N_10304,N_10407);
xor U10741 (N_10741,N_10346,N_10356);
xor U10742 (N_10742,N_10317,N_10293);
nor U10743 (N_10743,N_10292,N_10307);
nand U10744 (N_10744,N_10320,N_10490);
or U10745 (N_10745,N_10421,N_10370);
or U10746 (N_10746,N_10401,N_10432);
and U10747 (N_10747,N_10482,N_10278);
xor U10748 (N_10748,N_10482,N_10418);
nor U10749 (N_10749,N_10435,N_10292);
and U10750 (N_10750,N_10577,N_10589);
or U10751 (N_10751,N_10534,N_10636);
xnor U10752 (N_10752,N_10653,N_10604);
nor U10753 (N_10753,N_10651,N_10718);
nand U10754 (N_10754,N_10678,N_10683);
or U10755 (N_10755,N_10500,N_10521);
nor U10756 (N_10756,N_10597,N_10606);
xnor U10757 (N_10757,N_10512,N_10705);
nor U10758 (N_10758,N_10626,N_10695);
xor U10759 (N_10759,N_10553,N_10572);
or U10760 (N_10760,N_10684,N_10689);
nand U10761 (N_10761,N_10704,N_10531);
nor U10762 (N_10762,N_10507,N_10586);
nor U10763 (N_10763,N_10628,N_10729);
xor U10764 (N_10764,N_10536,N_10733);
nand U10765 (N_10765,N_10532,N_10625);
or U10766 (N_10766,N_10746,N_10615);
xor U10767 (N_10767,N_10621,N_10595);
nand U10768 (N_10768,N_10730,N_10598);
nand U10769 (N_10769,N_10619,N_10697);
or U10770 (N_10770,N_10709,N_10554);
or U10771 (N_10771,N_10711,N_10647);
or U10772 (N_10772,N_10545,N_10745);
or U10773 (N_10773,N_10583,N_10638);
and U10774 (N_10774,N_10543,N_10740);
and U10775 (N_10775,N_10620,N_10713);
nor U10776 (N_10776,N_10668,N_10656);
and U10777 (N_10777,N_10748,N_10557);
nand U10778 (N_10778,N_10546,N_10722);
or U10779 (N_10779,N_10588,N_10666);
and U10780 (N_10780,N_10712,N_10514);
nand U10781 (N_10781,N_10661,N_10503);
nand U10782 (N_10782,N_10516,N_10721);
xnor U10783 (N_10783,N_10560,N_10582);
nand U10784 (N_10784,N_10573,N_10699);
or U10785 (N_10785,N_10631,N_10579);
xnor U10786 (N_10786,N_10735,N_10743);
and U10787 (N_10787,N_10665,N_10544);
xnor U10788 (N_10788,N_10526,N_10701);
and U10789 (N_10789,N_10502,N_10622);
nor U10790 (N_10790,N_10508,N_10564);
nor U10791 (N_10791,N_10708,N_10731);
or U10792 (N_10792,N_10535,N_10616);
xor U10793 (N_10793,N_10570,N_10732);
or U10794 (N_10794,N_10541,N_10617);
xnor U10795 (N_10795,N_10667,N_10677);
xnor U10796 (N_10796,N_10723,N_10674);
xnor U10797 (N_10797,N_10600,N_10727);
nor U10798 (N_10798,N_10585,N_10710);
nand U10799 (N_10799,N_10609,N_10645);
and U10800 (N_10800,N_10646,N_10660);
nand U10801 (N_10801,N_10726,N_10670);
xor U10802 (N_10802,N_10679,N_10565);
xor U10803 (N_10803,N_10613,N_10574);
xnor U10804 (N_10804,N_10703,N_10728);
nor U10805 (N_10805,N_10632,N_10618);
xor U10806 (N_10806,N_10691,N_10637);
and U10807 (N_10807,N_10652,N_10571);
or U10808 (N_10808,N_10644,N_10623);
xnor U10809 (N_10809,N_10608,N_10707);
and U10810 (N_10810,N_10686,N_10593);
or U10811 (N_10811,N_10737,N_10659);
xor U10812 (N_10812,N_10696,N_10717);
xor U10813 (N_10813,N_10720,N_10738);
and U10814 (N_10814,N_10603,N_10654);
nand U10815 (N_10815,N_10662,N_10657);
nand U10816 (N_10816,N_10513,N_10568);
nor U10817 (N_10817,N_10551,N_10555);
nand U10818 (N_10818,N_10675,N_10584);
nor U10819 (N_10819,N_10742,N_10518);
nor U10820 (N_10820,N_10639,N_10749);
nor U10821 (N_10821,N_10578,N_10538);
nand U10822 (N_10822,N_10702,N_10591);
or U10823 (N_10823,N_10673,N_10747);
and U10824 (N_10824,N_10611,N_10547);
or U10825 (N_10825,N_10529,N_10580);
or U10826 (N_10826,N_10641,N_10642);
xnor U10827 (N_10827,N_10655,N_10575);
nor U10828 (N_10828,N_10561,N_10627);
nand U10829 (N_10829,N_10511,N_10550);
nand U10830 (N_10830,N_10510,N_10537);
nand U10831 (N_10831,N_10607,N_10694);
and U10832 (N_10832,N_10596,N_10629);
and U10833 (N_10833,N_10592,N_10716);
nand U10834 (N_10834,N_10548,N_10681);
and U10835 (N_10835,N_10685,N_10515);
nand U10836 (N_10836,N_10624,N_10590);
or U10837 (N_10837,N_10599,N_10528);
and U10838 (N_10838,N_10663,N_10719);
or U10839 (N_10839,N_10552,N_10725);
nor U10840 (N_10840,N_10635,N_10739);
xnor U10841 (N_10841,N_10527,N_10688);
or U10842 (N_10842,N_10672,N_10525);
and U10843 (N_10843,N_10576,N_10601);
and U10844 (N_10844,N_10501,N_10505);
and U10845 (N_10845,N_10610,N_10676);
nor U10846 (N_10846,N_10680,N_10509);
nand U10847 (N_10847,N_10700,N_10633);
or U10848 (N_10848,N_10744,N_10736);
and U10849 (N_10849,N_10520,N_10690);
or U10850 (N_10850,N_10530,N_10715);
xnor U10851 (N_10851,N_10567,N_10698);
nor U10852 (N_10852,N_10558,N_10556);
and U10853 (N_10853,N_10594,N_10540);
or U10854 (N_10854,N_10539,N_10533);
nor U10855 (N_10855,N_10506,N_10741);
or U10856 (N_10856,N_10559,N_10669);
nor U10857 (N_10857,N_10602,N_10671);
xor U10858 (N_10858,N_10687,N_10612);
xnor U10859 (N_10859,N_10524,N_10587);
nand U10860 (N_10860,N_10648,N_10734);
or U10861 (N_10861,N_10649,N_10523);
xor U10862 (N_10862,N_10563,N_10614);
and U10863 (N_10863,N_10519,N_10658);
and U10864 (N_10864,N_10549,N_10566);
or U10865 (N_10865,N_10640,N_10569);
and U10866 (N_10866,N_10504,N_10581);
xor U10867 (N_10867,N_10724,N_10562);
nand U10868 (N_10868,N_10634,N_10706);
nor U10869 (N_10869,N_10714,N_10522);
nor U10870 (N_10870,N_10643,N_10605);
or U10871 (N_10871,N_10693,N_10517);
nand U10872 (N_10872,N_10682,N_10630);
and U10873 (N_10873,N_10542,N_10692);
xnor U10874 (N_10874,N_10664,N_10650);
nor U10875 (N_10875,N_10714,N_10592);
and U10876 (N_10876,N_10554,N_10583);
xnor U10877 (N_10877,N_10544,N_10617);
xor U10878 (N_10878,N_10646,N_10701);
and U10879 (N_10879,N_10730,N_10713);
nand U10880 (N_10880,N_10672,N_10728);
nor U10881 (N_10881,N_10648,N_10516);
nand U10882 (N_10882,N_10739,N_10522);
xor U10883 (N_10883,N_10533,N_10688);
or U10884 (N_10884,N_10636,N_10586);
xnor U10885 (N_10885,N_10512,N_10555);
nor U10886 (N_10886,N_10612,N_10721);
or U10887 (N_10887,N_10730,N_10602);
nor U10888 (N_10888,N_10722,N_10622);
or U10889 (N_10889,N_10577,N_10520);
or U10890 (N_10890,N_10625,N_10709);
xnor U10891 (N_10891,N_10605,N_10725);
and U10892 (N_10892,N_10712,N_10531);
or U10893 (N_10893,N_10512,N_10718);
xnor U10894 (N_10894,N_10743,N_10648);
nor U10895 (N_10895,N_10740,N_10723);
or U10896 (N_10896,N_10677,N_10717);
xor U10897 (N_10897,N_10704,N_10745);
nand U10898 (N_10898,N_10633,N_10723);
nor U10899 (N_10899,N_10672,N_10663);
nor U10900 (N_10900,N_10642,N_10528);
xnor U10901 (N_10901,N_10573,N_10533);
or U10902 (N_10902,N_10561,N_10597);
xor U10903 (N_10903,N_10616,N_10627);
nor U10904 (N_10904,N_10549,N_10595);
nand U10905 (N_10905,N_10668,N_10587);
nor U10906 (N_10906,N_10665,N_10628);
and U10907 (N_10907,N_10537,N_10738);
xnor U10908 (N_10908,N_10555,N_10670);
nor U10909 (N_10909,N_10645,N_10510);
or U10910 (N_10910,N_10670,N_10687);
or U10911 (N_10911,N_10618,N_10502);
nor U10912 (N_10912,N_10628,N_10626);
xnor U10913 (N_10913,N_10526,N_10557);
nor U10914 (N_10914,N_10607,N_10594);
nand U10915 (N_10915,N_10542,N_10684);
nor U10916 (N_10916,N_10624,N_10644);
xnor U10917 (N_10917,N_10511,N_10545);
nand U10918 (N_10918,N_10634,N_10749);
and U10919 (N_10919,N_10694,N_10624);
xor U10920 (N_10920,N_10594,N_10577);
or U10921 (N_10921,N_10650,N_10582);
nand U10922 (N_10922,N_10646,N_10554);
nand U10923 (N_10923,N_10574,N_10728);
nand U10924 (N_10924,N_10522,N_10692);
xor U10925 (N_10925,N_10710,N_10583);
and U10926 (N_10926,N_10557,N_10621);
and U10927 (N_10927,N_10552,N_10617);
nand U10928 (N_10928,N_10580,N_10616);
or U10929 (N_10929,N_10511,N_10540);
or U10930 (N_10930,N_10535,N_10517);
or U10931 (N_10931,N_10605,N_10736);
and U10932 (N_10932,N_10736,N_10623);
or U10933 (N_10933,N_10648,N_10649);
nand U10934 (N_10934,N_10505,N_10560);
nand U10935 (N_10935,N_10617,N_10633);
xor U10936 (N_10936,N_10732,N_10530);
or U10937 (N_10937,N_10593,N_10527);
nand U10938 (N_10938,N_10655,N_10519);
or U10939 (N_10939,N_10632,N_10661);
nor U10940 (N_10940,N_10654,N_10552);
nor U10941 (N_10941,N_10717,N_10663);
and U10942 (N_10942,N_10608,N_10635);
or U10943 (N_10943,N_10586,N_10549);
nor U10944 (N_10944,N_10527,N_10663);
and U10945 (N_10945,N_10588,N_10534);
or U10946 (N_10946,N_10558,N_10621);
xnor U10947 (N_10947,N_10659,N_10619);
nand U10948 (N_10948,N_10551,N_10536);
or U10949 (N_10949,N_10633,N_10537);
nand U10950 (N_10950,N_10508,N_10690);
or U10951 (N_10951,N_10545,N_10521);
nand U10952 (N_10952,N_10522,N_10510);
or U10953 (N_10953,N_10528,N_10596);
or U10954 (N_10954,N_10500,N_10658);
and U10955 (N_10955,N_10570,N_10514);
xor U10956 (N_10956,N_10688,N_10654);
xnor U10957 (N_10957,N_10655,N_10619);
and U10958 (N_10958,N_10621,N_10630);
nor U10959 (N_10959,N_10562,N_10659);
and U10960 (N_10960,N_10525,N_10513);
or U10961 (N_10961,N_10541,N_10573);
and U10962 (N_10962,N_10549,N_10539);
nand U10963 (N_10963,N_10540,N_10636);
nor U10964 (N_10964,N_10568,N_10562);
and U10965 (N_10965,N_10720,N_10510);
or U10966 (N_10966,N_10706,N_10628);
nand U10967 (N_10967,N_10538,N_10636);
or U10968 (N_10968,N_10728,N_10714);
nand U10969 (N_10969,N_10654,N_10535);
or U10970 (N_10970,N_10676,N_10595);
nor U10971 (N_10971,N_10551,N_10597);
and U10972 (N_10972,N_10511,N_10555);
nor U10973 (N_10973,N_10605,N_10710);
nand U10974 (N_10974,N_10719,N_10609);
or U10975 (N_10975,N_10615,N_10539);
xor U10976 (N_10976,N_10527,N_10607);
and U10977 (N_10977,N_10513,N_10550);
or U10978 (N_10978,N_10518,N_10668);
nor U10979 (N_10979,N_10625,N_10572);
nor U10980 (N_10980,N_10675,N_10544);
and U10981 (N_10981,N_10740,N_10550);
or U10982 (N_10982,N_10666,N_10506);
nand U10983 (N_10983,N_10622,N_10541);
nand U10984 (N_10984,N_10533,N_10740);
nand U10985 (N_10985,N_10668,N_10742);
nor U10986 (N_10986,N_10517,N_10541);
xnor U10987 (N_10987,N_10721,N_10566);
nor U10988 (N_10988,N_10534,N_10510);
nor U10989 (N_10989,N_10634,N_10656);
xnor U10990 (N_10990,N_10546,N_10651);
xor U10991 (N_10991,N_10703,N_10523);
or U10992 (N_10992,N_10566,N_10684);
nor U10993 (N_10993,N_10567,N_10723);
nand U10994 (N_10994,N_10677,N_10510);
nand U10995 (N_10995,N_10591,N_10516);
nand U10996 (N_10996,N_10684,N_10518);
nor U10997 (N_10997,N_10689,N_10505);
or U10998 (N_10998,N_10680,N_10643);
xor U10999 (N_10999,N_10679,N_10611);
or U11000 (N_11000,N_10829,N_10895);
xnor U11001 (N_11001,N_10921,N_10834);
and U11002 (N_11002,N_10854,N_10816);
and U11003 (N_11003,N_10795,N_10902);
or U11004 (N_11004,N_10917,N_10847);
and U11005 (N_11005,N_10856,N_10959);
xor U11006 (N_11006,N_10943,N_10791);
or U11007 (N_11007,N_10970,N_10956);
or U11008 (N_11008,N_10909,N_10877);
xor U11009 (N_11009,N_10842,N_10838);
and U11010 (N_11010,N_10860,N_10780);
nor U11011 (N_11011,N_10836,N_10910);
nor U11012 (N_11012,N_10813,N_10793);
or U11013 (N_11013,N_10951,N_10784);
or U11014 (N_11014,N_10881,N_10920);
nand U11015 (N_11015,N_10984,N_10769);
nor U11016 (N_11016,N_10789,N_10888);
or U11017 (N_11017,N_10996,N_10928);
or U11018 (N_11018,N_10983,N_10964);
xor U11019 (N_11019,N_10885,N_10971);
xor U11020 (N_11020,N_10782,N_10770);
and U11021 (N_11021,N_10999,N_10891);
nor U11022 (N_11022,N_10823,N_10764);
or U11023 (N_11023,N_10904,N_10805);
nor U11024 (N_11024,N_10967,N_10893);
nand U11025 (N_11025,N_10866,N_10945);
xor U11026 (N_11026,N_10905,N_10927);
and U11027 (N_11027,N_10901,N_10874);
xor U11028 (N_11028,N_10925,N_10892);
nor U11029 (N_11029,N_10840,N_10859);
xor U11030 (N_11030,N_10906,N_10852);
and U11031 (N_11031,N_10818,N_10792);
nor U11032 (N_11032,N_10988,N_10935);
nand U11033 (N_11033,N_10879,N_10760);
xnor U11034 (N_11034,N_10871,N_10875);
nor U11035 (N_11035,N_10837,N_10958);
or U11036 (N_11036,N_10946,N_10942);
nor U11037 (N_11037,N_10944,N_10977);
nand U11038 (N_11038,N_10978,N_10907);
nand U11039 (N_11039,N_10758,N_10973);
nand U11040 (N_11040,N_10765,N_10826);
and U11041 (N_11041,N_10822,N_10812);
nand U11042 (N_11042,N_10952,N_10884);
or U11043 (N_11043,N_10773,N_10912);
and U11044 (N_11044,N_10939,N_10987);
nor U11045 (N_11045,N_10807,N_10751);
and U11046 (N_11046,N_10811,N_10994);
and U11047 (N_11047,N_10940,N_10991);
and U11048 (N_11048,N_10843,N_10880);
nand U11049 (N_11049,N_10908,N_10766);
and U11050 (N_11050,N_10980,N_10899);
nand U11051 (N_11051,N_10771,N_10848);
nand U11052 (N_11052,N_10986,N_10915);
nor U11053 (N_11053,N_10786,N_10778);
and U11054 (N_11054,N_10981,N_10814);
nand U11055 (N_11055,N_10982,N_10998);
or U11056 (N_11056,N_10832,N_10897);
or U11057 (N_11057,N_10948,N_10775);
nor U11058 (N_11058,N_10916,N_10869);
nor U11059 (N_11059,N_10853,N_10867);
xnor U11060 (N_11060,N_10864,N_10754);
and U11061 (N_11061,N_10803,N_10955);
and U11062 (N_11062,N_10750,N_10845);
nand U11063 (N_11063,N_10878,N_10796);
xnor U11064 (N_11064,N_10933,N_10900);
or U11065 (N_11065,N_10756,N_10833);
xor U11066 (N_11066,N_10768,N_10835);
and U11067 (N_11067,N_10753,N_10930);
nand U11068 (N_11068,N_10993,N_10763);
nor U11069 (N_11069,N_10990,N_10911);
and U11070 (N_11070,N_10785,N_10972);
nor U11071 (N_11071,N_10886,N_10941);
nor U11072 (N_11072,N_10887,N_10932);
and U11073 (N_11073,N_10918,N_10827);
nand U11074 (N_11074,N_10808,N_10809);
and U11075 (N_11075,N_10868,N_10966);
nand U11076 (N_11076,N_10819,N_10790);
and U11077 (N_11077,N_10774,N_10776);
xnor U11078 (N_11078,N_10989,N_10851);
nand U11079 (N_11079,N_10979,N_10913);
or U11080 (N_11080,N_10938,N_10865);
nand U11081 (N_11081,N_10844,N_10922);
or U11082 (N_11082,N_10873,N_10855);
and U11083 (N_11083,N_10894,N_10762);
and U11084 (N_11084,N_10936,N_10947);
or U11085 (N_11085,N_10759,N_10883);
and U11086 (N_11086,N_10804,N_10962);
nand U11087 (N_11087,N_10872,N_10968);
and U11088 (N_11088,N_10882,N_10779);
xor U11089 (N_11089,N_10861,N_10755);
nand U11090 (N_11090,N_10963,N_10969);
or U11091 (N_11091,N_10924,N_10976);
nand U11092 (N_11092,N_10949,N_10934);
or U11093 (N_11093,N_10761,N_10849);
or U11094 (N_11094,N_10806,N_10799);
or U11095 (N_11095,N_10817,N_10820);
and U11096 (N_11096,N_10801,N_10794);
nand U11097 (N_11097,N_10997,N_10929);
and U11098 (N_11098,N_10890,N_10954);
or U11099 (N_11099,N_10846,N_10923);
nor U11100 (N_11100,N_10752,N_10858);
nand U11101 (N_11101,N_10757,N_10957);
xnor U11102 (N_11102,N_10876,N_10800);
and U11103 (N_11103,N_10931,N_10850);
or U11104 (N_11104,N_10815,N_10830);
and U11105 (N_11105,N_10995,N_10787);
and U11106 (N_11106,N_10767,N_10974);
nand U11107 (N_11107,N_10926,N_10825);
nor U11108 (N_11108,N_10870,N_10919);
nand U11109 (N_11109,N_10810,N_10788);
xnor U11110 (N_11110,N_10953,N_10965);
or U11111 (N_11111,N_10903,N_10828);
and U11112 (N_11112,N_10824,N_10898);
xor U11113 (N_11113,N_10896,N_10914);
nand U11114 (N_11114,N_10777,N_10950);
nand U11115 (N_11115,N_10772,N_10839);
nor U11116 (N_11116,N_10781,N_10862);
nor U11117 (N_11117,N_10857,N_10889);
and U11118 (N_11118,N_10992,N_10960);
and U11119 (N_11119,N_10961,N_10797);
xnor U11120 (N_11120,N_10798,N_10802);
nand U11121 (N_11121,N_10783,N_10975);
nand U11122 (N_11122,N_10985,N_10937);
nor U11123 (N_11123,N_10841,N_10863);
or U11124 (N_11124,N_10831,N_10821);
nor U11125 (N_11125,N_10945,N_10885);
xnor U11126 (N_11126,N_10858,N_10784);
nor U11127 (N_11127,N_10861,N_10857);
or U11128 (N_11128,N_10790,N_10944);
nor U11129 (N_11129,N_10851,N_10871);
xor U11130 (N_11130,N_10841,N_10933);
xor U11131 (N_11131,N_10874,N_10956);
nand U11132 (N_11132,N_10764,N_10900);
nand U11133 (N_11133,N_10980,N_10790);
and U11134 (N_11134,N_10987,N_10971);
nor U11135 (N_11135,N_10860,N_10947);
xor U11136 (N_11136,N_10874,N_10842);
nand U11137 (N_11137,N_10785,N_10773);
or U11138 (N_11138,N_10835,N_10759);
xnor U11139 (N_11139,N_10815,N_10829);
or U11140 (N_11140,N_10901,N_10917);
or U11141 (N_11141,N_10812,N_10916);
or U11142 (N_11142,N_10832,N_10753);
and U11143 (N_11143,N_10840,N_10972);
and U11144 (N_11144,N_10877,N_10939);
xor U11145 (N_11145,N_10819,N_10802);
or U11146 (N_11146,N_10798,N_10984);
and U11147 (N_11147,N_10837,N_10967);
nor U11148 (N_11148,N_10960,N_10839);
xnor U11149 (N_11149,N_10845,N_10810);
nor U11150 (N_11150,N_10972,N_10773);
xor U11151 (N_11151,N_10938,N_10921);
and U11152 (N_11152,N_10829,N_10752);
or U11153 (N_11153,N_10790,N_10900);
and U11154 (N_11154,N_10853,N_10840);
xor U11155 (N_11155,N_10962,N_10940);
xor U11156 (N_11156,N_10776,N_10957);
or U11157 (N_11157,N_10836,N_10794);
or U11158 (N_11158,N_10813,N_10993);
nand U11159 (N_11159,N_10868,N_10859);
nor U11160 (N_11160,N_10797,N_10821);
nor U11161 (N_11161,N_10776,N_10807);
nand U11162 (N_11162,N_10997,N_10815);
and U11163 (N_11163,N_10891,N_10913);
nor U11164 (N_11164,N_10821,N_10969);
nand U11165 (N_11165,N_10800,N_10885);
nor U11166 (N_11166,N_10870,N_10828);
and U11167 (N_11167,N_10999,N_10967);
nand U11168 (N_11168,N_10910,N_10859);
nor U11169 (N_11169,N_10907,N_10866);
or U11170 (N_11170,N_10987,N_10941);
xor U11171 (N_11171,N_10805,N_10900);
and U11172 (N_11172,N_10758,N_10883);
or U11173 (N_11173,N_10769,N_10829);
nor U11174 (N_11174,N_10844,N_10895);
nand U11175 (N_11175,N_10870,N_10897);
or U11176 (N_11176,N_10937,N_10765);
xnor U11177 (N_11177,N_10756,N_10898);
nor U11178 (N_11178,N_10786,N_10877);
nor U11179 (N_11179,N_10773,N_10834);
nand U11180 (N_11180,N_10973,N_10912);
nor U11181 (N_11181,N_10961,N_10912);
or U11182 (N_11182,N_10883,N_10897);
xor U11183 (N_11183,N_10805,N_10826);
xnor U11184 (N_11184,N_10918,N_10760);
nand U11185 (N_11185,N_10957,N_10949);
and U11186 (N_11186,N_10750,N_10929);
or U11187 (N_11187,N_10858,N_10872);
nand U11188 (N_11188,N_10926,N_10908);
nor U11189 (N_11189,N_10824,N_10808);
and U11190 (N_11190,N_10751,N_10801);
xor U11191 (N_11191,N_10989,N_10804);
nand U11192 (N_11192,N_10866,N_10883);
nor U11193 (N_11193,N_10890,N_10881);
xor U11194 (N_11194,N_10999,N_10803);
xnor U11195 (N_11195,N_10862,N_10865);
nand U11196 (N_11196,N_10831,N_10974);
nand U11197 (N_11197,N_10930,N_10807);
and U11198 (N_11198,N_10832,N_10913);
or U11199 (N_11199,N_10791,N_10897);
and U11200 (N_11200,N_10968,N_10994);
nand U11201 (N_11201,N_10915,N_10826);
nand U11202 (N_11202,N_10890,N_10877);
and U11203 (N_11203,N_10750,N_10792);
nand U11204 (N_11204,N_10951,N_10797);
or U11205 (N_11205,N_10873,N_10930);
or U11206 (N_11206,N_10817,N_10938);
xor U11207 (N_11207,N_10810,N_10860);
nor U11208 (N_11208,N_10962,N_10995);
nor U11209 (N_11209,N_10979,N_10788);
nand U11210 (N_11210,N_10875,N_10997);
and U11211 (N_11211,N_10764,N_10861);
nor U11212 (N_11212,N_10991,N_10946);
or U11213 (N_11213,N_10961,N_10891);
nor U11214 (N_11214,N_10833,N_10927);
xor U11215 (N_11215,N_10830,N_10914);
and U11216 (N_11216,N_10968,N_10996);
nand U11217 (N_11217,N_10773,N_10890);
or U11218 (N_11218,N_10950,N_10995);
and U11219 (N_11219,N_10900,N_10872);
nand U11220 (N_11220,N_10764,N_10760);
nand U11221 (N_11221,N_10867,N_10855);
and U11222 (N_11222,N_10870,N_10972);
xnor U11223 (N_11223,N_10958,N_10862);
or U11224 (N_11224,N_10812,N_10971);
nand U11225 (N_11225,N_10914,N_10845);
nor U11226 (N_11226,N_10935,N_10855);
and U11227 (N_11227,N_10949,N_10859);
xor U11228 (N_11228,N_10772,N_10970);
nor U11229 (N_11229,N_10885,N_10901);
xnor U11230 (N_11230,N_10923,N_10803);
and U11231 (N_11231,N_10971,N_10970);
nand U11232 (N_11232,N_10890,N_10803);
nand U11233 (N_11233,N_10966,N_10975);
or U11234 (N_11234,N_10777,N_10820);
or U11235 (N_11235,N_10874,N_10876);
and U11236 (N_11236,N_10927,N_10800);
xor U11237 (N_11237,N_10831,N_10818);
nor U11238 (N_11238,N_10790,N_10915);
nor U11239 (N_11239,N_10781,N_10858);
or U11240 (N_11240,N_10857,N_10836);
nor U11241 (N_11241,N_10942,N_10931);
or U11242 (N_11242,N_10901,N_10802);
nor U11243 (N_11243,N_10894,N_10891);
nand U11244 (N_11244,N_10909,N_10852);
nor U11245 (N_11245,N_10839,N_10790);
or U11246 (N_11246,N_10872,N_10940);
xnor U11247 (N_11247,N_10928,N_10880);
nor U11248 (N_11248,N_10979,N_10780);
nor U11249 (N_11249,N_10899,N_10837);
nand U11250 (N_11250,N_11138,N_11039);
and U11251 (N_11251,N_11143,N_11059);
xnor U11252 (N_11252,N_11158,N_11065);
or U11253 (N_11253,N_11246,N_11153);
nand U11254 (N_11254,N_11235,N_11102);
nand U11255 (N_11255,N_11096,N_11064);
xnor U11256 (N_11256,N_11201,N_11181);
or U11257 (N_11257,N_11193,N_11041);
and U11258 (N_11258,N_11042,N_11229);
nand U11259 (N_11259,N_11133,N_11047);
or U11260 (N_11260,N_11204,N_11233);
xnor U11261 (N_11261,N_11234,N_11018);
and U11262 (N_11262,N_11186,N_11076);
and U11263 (N_11263,N_11021,N_11142);
nor U11264 (N_11264,N_11090,N_11216);
and U11265 (N_11265,N_11182,N_11167);
nand U11266 (N_11266,N_11208,N_11245);
xnor U11267 (N_11267,N_11100,N_11173);
or U11268 (N_11268,N_11132,N_11134);
and U11269 (N_11269,N_11237,N_11110);
nor U11270 (N_11270,N_11077,N_11221);
and U11271 (N_11271,N_11147,N_11057);
xnor U11272 (N_11272,N_11152,N_11199);
and U11273 (N_11273,N_11044,N_11084);
or U11274 (N_11274,N_11004,N_11187);
or U11275 (N_11275,N_11247,N_11119);
nor U11276 (N_11276,N_11175,N_11121);
nand U11277 (N_11277,N_11050,N_11055);
nand U11278 (N_11278,N_11013,N_11011);
or U11279 (N_11279,N_11178,N_11014);
nor U11280 (N_11280,N_11239,N_11189);
xnor U11281 (N_11281,N_11070,N_11206);
nor U11282 (N_11282,N_11060,N_11176);
nand U11283 (N_11283,N_11174,N_11035);
nand U11284 (N_11284,N_11095,N_11051);
nor U11285 (N_11285,N_11067,N_11197);
xor U11286 (N_11286,N_11179,N_11217);
or U11287 (N_11287,N_11037,N_11194);
or U11288 (N_11288,N_11160,N_11108);
or U11289 (N_11289,N_11098,N_11107);
nor U11290 (N_11290,N_11029,N_11116);
nand U11291 (N_11291,N_11122,N_11205);
and U11292 (N_11292,N_11117,N_11017);
and U11293 (N_11293,N_11040,N_11080);
nor U11294 (N_11294,N_11180,N_11043);
xnor U11295 (N_11295,N_11151,N_11145);
or U11296 (N_11296,N_11113,N_11123);
or U11297 (N_11297,N_11222,N_11000);
nor U11298 (N_11298,N_11045,N_11156);
and U11299 (N_11299,N_11232,N_11196);
xnor U11300 (N_11300,N_11248,N_11219);
xor U11301 (N_11301,N_11089,N_11038);
xnor U11302 (N_11302,N_11169,N_11099);
xor U11303 (N_11303,N_11227,N_11088);
or U11304 (N_11304,N_11225,N_11114);
nand U11305 (N_11305,N_11028,N_11190);
nand U11306 (N_11306,N_11074,N_11104);
or U11307 (N_11307,N_11112,N_11052);
nand U11308 (N_11308,N_11048,N_11207);
nor U11309 (N_11309,N_11034,N_11185);
nor U11310 (N_11310,N_11071,N_11127);
nor U11311 (N_11311,N_11144,N_11009);
nor U11312 (N_11312,N_11023,N_11124);
xnor U11313 (N_11313,N_11027,N_11022);
nor U11314 (N_11314,N_11163,N_11129);
and U11315 (N_11315,N_11053,N_11137);
nor U11316 (N_11316,N_11103,N_11008);
or U11317 (N_11317,N_11202,N_11068);
nor U11318 (N_11318,N_11184,N_11168);
nor U11319 (N_11319,N_11192,N_11091);
and U11320 (N_11320,N_11230,N_11015);
nor U11321 (N_11321,N_11200,N_11125);
nor U11322 (N_11322,N_11061,N_11001);
or U11323 (N_11323,N_11036,N_11003);
and U11324 (N_11324,N_11213,N_11062);
nand U11325 (N_11325,N_11058,N_11170);
nand U11326 (N_11326,N_11162,N_11079);
xor U11327 (N_11327,N_11066,N_11243);
and U11328 (N_11328,N_11228,N_11082);
nor U11329 (N_11329,N_11120,N_11126);
or U11330 (N_11330,N_11092,N_11203);
and U11331 (N_11331,N_11073,N_11069);
nor U11332 (N_11332,N_11198,N_11083);
nor U11333 (N_11333,N_11210,N_11002);
nor U11334 (N_11334,N_11010,N_11249);
nand U11335 (N_11335,N_11244,N_11131);
nand U11336 (N_11336,N_11242,N_11109);
and U11337 (N_11337,N_11140,N_11072);
nor U11338 (N_11338,N_11086,N_11240);
and U11339 (N_11339,N_11209,N_11165);
nand U11340 (N_11340,N_11220,N_11155);
or U11341 (N_11341,N_11223,N_11172);
xnor U11342 (N_11342,N_11012,N_11106);
nor U11343 (N_11343,N_11211,N_11177);
and U11344 (N_11344,N_11195,N_11191);
or U11345 (N_11345,N_11136,N_11183);
xnor U11346 (N_11346,N_11157,N_11016);
and U11347 (N_11347,N_11161,N_11141);
and U11348 (N_11348,N_11007,N_11063);
and U11349 (N_11349,N_11171,N_11032);
nor U11350 (N_11350,N_11049,N_11081);
and U11351 (N_11351,N_11115,N_11130);
nand U11352 (N_11352,N_11212,N_11215);
or U11353 (N_11353,N_11166,N_11146);
and U11354 (N_11354,N_11236,N_11078);
xnor U11355 (N_11355,N_11164,N_11139);
nand U11356 (N_11356,N_11033,N_11094);
nand U11357 (N_11357,N_11024,N_11128);
and U11358 (N_11358,N_11241,N_11025);
xor U11359 (N_11359,N_11026,N_11075);
xnor U11360 (N_11360,N_11188,N_11020);
or U11361 (N_11361,N_11154,N_11105);
xnor U11362 (N_11362,N_11046,N_11006);
nand U11363 (N_11363,N_11231,N_11159);
or U11364 (N_11364,N_11224,N_11005);
nor U11365 (N_11365,N_11150,N_11226);
nand U11366 (N_11366,N_11054,N_11087);
or U11367 (N_11367,N_11101,N_11111);
and U11368 (N_11368,N_11238,N_11097);
xor U11369 (N_11369,N_11031,N_11218);
or U11370 (N_11370,N_11056,N_11148);
and U11371 (N_11371,N_11118,N_11085);
and U11372 (N_11372,N_11093,N_11030);
nand U11373 (N_11373,N_11019,N_11135);
xor U11374 (N_11374,N_11214,N_11149);
nor U11375 (N_11375,N_11084,N_11201);
and U11376 (N_11376,N_11235,N_11027);
nand U11377 (N_11377,N_11174,N_11039);
and U11378 (N_11378,N_11041,N_11156);
xnor U11379 (N_11379,N_11112,N_11097);
nor U11380 (N_11380,N_11003,N_11042);
xnor U11381 (N_11381,N_11206,N_11075);
nand U11382 (N_11382,N_11061,N_11017);
nand U11383 (N_11383,N_11092,N_11126);
xnor U11384 (N_11384,N_11054,N_11160);
or U11385 (N_11385,N_11110,N_11077);
and U11386 (N_11386,N_11226,N_11086);
nor U11387 (N_11387,N_11234,N_11038);
nand U11388 (N_11388,N_11221,N_11175);
nor U11389 (N_11389,N_11050,N_11210);
xnor U11390 (N_11390,N_11225,N_11167);
nand U11391 (N_11391,N_11169,N_11154);
nand U11392 (N_11392,N_11230,N_11090);
and U11393 (N_11393,N_11037,N_11066);
xnor U11394 (N_11394,N_11248,N_11001);
nand U11395 (N_11395,N_11126,N_11000);
or U11396 (N_11396,N_11219,N_11113);
nor U11397 (N_11397,N_11007,N_11098);
nand U11398 (N_11398,N_11059,N_11027);
nor U11399 (N_11399,N_11111,N_11239);
nand U11400 (N_11400,N_11130,N_11192);
nor U11401 (N_11401,N_11041,N_11105);
or U11402 (N_11402,N_11011,N_11019);
nor U11403 (N_11403,N_11232,N_11040);
and U11404 (N_11404,N_11045,N_11187);
nor U11405 (N_11405,N_11072,N_11206);
xor U11406 (N_11406,N_11086,N_11221);
xnor U11407 (N_11407,N_11194,N_11002);
or U11408 (N_11408,N_11146,N_11002);
nor U11409 (N_11409,N_11074,N_11091);
xor U11410 (N_11410,N_11233,N_11175);
nand U11411 (N_11411,N_11193,N_11050);
xor U11412 (N_11412,N_11158,N_11219);
or U11413 (N_11413,N_11017,N_11190);
nand U11414 (N_11414,N_11013,N_11054);
xor U11415 (N_11415,N_11198,N_11155);
nand U11416 (N_11416,N_11115,N_11226);
or U11417 (N_11417,N_11225,N_11206);
and U11418 (N_11418,N_11174,N_11112);
or U11419 (N_11419,N_11167,N_11031);
or U11420 (N_11420,N_11158,N_11085);
or U11421 (N_11421,N_11163,N_11069);
xor U11422 (N_11422,N_11201,N_11231);
xor U11423 (N_11423,N_11087,N_11019);
xor U11424 (N_11424,N_11009,N_11151);
and U11425 (N_11425,N_11109,N_11180);
nand U11426 (N_11426,N_11141,N_11046);
xor U11427 (N_11427,N_11042,N_11215);
nand U11428 (N_11428,N_11130,N_11132);
xor U11429 (N_11429,N_11167,N_11002);
nand U11430 (N_11430,N_11199,N_11140);
nor U11431 (N_11431,N_11229,N_11029);
xor U11432 (N_11432,N_11063,N_11052);
xnor U11433 (N_11433,N_11021,N_11075);
xor U11434 (N_11434,N_11124,N_11038);
or U11435 (N_11435,N_11226,N_11207);
xor U11436 (N_11436,N_11197,N_11187);
or U11437 (N_11437,N_11139,N_11200);
nor U11438 (N_11438,N_11159,N_11075);
xor U11439 (N_11439,N_11004,N_11102);
or U11440 (N_11440,N_11171,N_11125);
and U11441 (N_11441,N_11113,N_11197);
or U11442 (N_11442,N_11124,N_11056);
xnor U11443 (N_11443,N_11104,N_11041);
nor U11444 (N_11444,N_11021,N_11247);
and U11445 (N_11445,N_11138,N_11218);
or U11446 (N_11446,N_11202,N_11237);
and U11447 (N_11447,N_11100,N_11247);
or U11448 (N_11448,N_11218,N_11107);
or U11449 (N_11449,N_11122,N_11048);
nor U11450 (N_11450,N_11073,N_11164);
and U11451 (N_11451,N_11019,N_11010);
or U11452 (N_11452,N_11060,N_11241);
and U11453 (N_11453,N_11236,N_11146);
nand U11454 (N_11454,N_11008,N_11092);
and U11455 (N_11455,N_11192,N_11165);
xor U11456 (N_11456,N_11216,N_11141);
and U11457 (N_11457,N_11151,N_11182);
nand U11458 (N_11458,N_11099,N_11087);
or U11459 (N_11459,N_11153,N_11031);
or U11460 (N_11460,N_11208,N_11035);
and U11461 (N_11461,N_11181,N_11069);
and U11462 (N_11462,N_11069,N_11249);
or U11463 (N_11463,N_11194,N_11187);
nor U11464 (N_11464,N_11039,N_11028);
nand U11465 (N_11465,N_11190,N_11182);
nand U11466 (N_11466,N_11004,N_11091);
and U11467 (N_11467,N_11077,N_11003);
or U11468 (N_11468,N_11239,N_11114);
nor U11469 (N_11469,N_11013,N_11173);
nor U11470 (N_11470,N_11155,N_11056);
nand U11471 (N_11471,N_11007,N_11081);
nor U11472 (N_11472,N_11059,N_11205);
or U11473 (N_11473,N_11013,N_11104);
and U11474 (N_11474,N_11045,N_11072);
xor U11475 (N_11475,N_11059,N_11079);
nor U11476 (N_11476,N_11239,N_11044);
nor U11477 (N_11477,N_11233,N_11122);
nand U11478 (N_11478,N_11125,N_11184);
nor U11479 (N_11479,N_11127,N_11213);
and U11480 (N_11480,N_11082,N_11199);
and U11481 (N_11481,N_11091,N_11089);
xor U11482 (N_11482,N_11117,N_11247);
nor U11483 (N_11483,N_11071,N_11105);
or U11484 (N_11484,N_11010,N_11169);
and U11485 (N_11485,N_11245,N_11240);
nor U11486 (N_11486,N_11143,N_11177);
nor U11487 (N_11487,N_11156,N_11159);
nor U11488 (N_11488,N_11075,N_11192);
xor U11489 (N_11489,N_11114,N_11168);
or U11490 (N_11490,N_11153,N_11062);
xnor U11491 (N_11491,N_11113,N_11127);
nor U11492 (N_11492,N_11078,N_11032);
xor U11493 (N_11493,N_11190,N_11234);
xnor U11494 (N_11494,N_11189,N_11162);
and U11495 (N_11495,N_11205,N_11031);
nor U11496 (N_11496,N_11070,N_11038);
or U11497 (N_11497,N_11062,N_11065);
nor U11498 (N_11498,N_11095,N_11142);
xnor U11499 (N_11499,N_11113,N_11230);
xor U11500 (N_11500,N_11429,N_11420);
nand U11501 (N_11501,N_11282,N_11303);
nand U11502 (N_11502,N_11457,N_11460);
xnor U11503 (N_11503,N_11328,N_11325);
nor U11504 (N_11504,N_11427,N_11413);
nand U11505 (N_11505,N_11292,N_11466);
nand U11506 (N_11506,N_11480,N_11331);
nor U11507 (N_11507,N_11306,N_11456);
nand U11508 (N_11508,N_11266,N_11327);
xor U11509 (N_11509,N_11339,N_11349);
xnor U11510 (N_11510,N_11484,N_11297);
nand U11511 (N_11511,N_11486,N_11476);
or U11512 (N_11512,N_11468,N_11305);
nand U11513 (N_11513,N_11312,N_11462);
nor U11514 (N_11514,N_11489,N_11492);
xnor U11515 (N_11515,N_11357,N_11416);
and U11516 (N_11516,N_11419,N_11381);
or U11517 (N_11517,N_11388,N_11446);
xnor U11518 (N_11518,N_11285,N_11371);
or U11519 (N_11519,N_11481,N_11264);
nand U11520 (N_11520,N_11311,N_11370);
xor U11521 (N_11521,N_11400,N_11295);
or U11522 (N_11522,N_11404,N_11307);
or U11523 (N_11523,N_11324,N_11254);
xnor U11524 (N_11524,N_11342,N_11464);
or U11525 (N_11525,N_11380,N_11401);
nand U11526 (N_11526,N_11334,N_11428);
nor U11527 (N_11527,N_11274,N_11473);
xnor U11528 (N_11528,N_11436,N_11434);
and U11529 (N_11529,N_11362,N_11448);
xnor U11530 (N_11530,N_11403,N_11373);
or U11531 (N_11531,N_11316,N_11402);
nand U11532 (N_11532,N_11353,N_11343);
and U11533 (N_11533,N_11433,N_11412);
xnor U11534 (N_11534,N_11321,N_11344);
and U11535 (N_11535,N_11372,N_11273);
or U11536 (N_11536,N_11392,N_11320);
nand U11537 (N_11537,N_11252,N_11424);
and U11538 (N_11538,N_11435,N_11463);
xor U11539 (N_11539,N_11449,N_11439);
xor U11540 (N_11540,N_11317,N_11354);
nor U11541 (N_11541,N_11265,N_11315);
and U11542 (N_11542,N_11361,N_11386);
xor U11543 (N_11543,N_11368,N_11279);
xor U11544 (N_11544,N_11437,N_11425);
nor U11545 (N_11545,N_11387,N_11385);
nor U11546 (N_11546,N_11482,N_11499);
nor U11547 (N_11547,N_11330,N_11352);
nand U11548 (N_11548,N_11287,N_11491);
or U11549 (N_11549,N_11277,N_11258);
or U11550 (N_11550,N_11333,N_11391);
or U11551 (N_11551,N_11286,N_11470);
or U11552 (N_11552,N_11408,N_11399);
or U11553 (N_11553,N_11341,N_11300);
nand U11554 (N_11554,N_11421,N_11251);
or U11555 (N_11555,N_11418,N_11454);
and U11556 (N_11556,N_11423,N_11309);
xnor U11557 (N_11557,N_11291,N_11256);
and U11558 (N_11558,N_11494,N_11255);
and U11559 (N_11559,N_11363,N_11280);
xnor U11560 (N_11560,N_11467,N_11459);
nand U11561 (N_11561,N_11496,N_11493);
xnor U11562 (N_11562,N_11369,N_11472);
nand U11563 (N_11563,N_11374,N_11348);
nor U11564 (N_11564,N_11398,N_11445);
nand U11565 (N_11565,N_11313,N_11284);
nand U11566 (N_11566,N_11478,N_11319);
nor U11567 (N_11567,N_11278,N_11383);
nand U11568 (N_11568,N_11471,N_11294);
xnor U11569 (N_11569,N_11406,N_11411);
nor U11570 (N_11570,N_11422,N_11356);
or U11571 (N_11571,N_11393,N_11430);
xor U11572 (N_11572,N_11301,N_11323);
xor U11573 (N_11573,N_11453,N_11263);
nand U11574 (N_11574,N_11304,N_11440);
nor U11575 (N_11575,N_11497,N_11350);
nand U11576 (N_11576,N_11271,N_11367);
or U11577 (N_11577,N_11310,N_11272);
xor U11578 (N_11578,N_11415,N_11431);
and U11579 (N_11579,N_11336,N_11455);
or U11580 (N_11580,N_11340,N_11329);
nor U11581 (N_11581,N_11322,N_11358);
nand U11582 (N_11582,N_11298,N_11347);
xor U11583 (N_11583,N_11394,N_11337);
and U11584 (N_11584,N_11426,N_11396);
nand U11585 (N_11585,N_11346,N_11332);
nand U11586 (N_11586,N_11293,N_11268);
nand U11587 (N_11587,N_11269,N_11360);
xor U11588 (N_11588,N_11299,N_11442);
nor U11589 (N_11589,N_11366,N_11275);
or U11590 (N_11590,N_11465,N_11479);
and U11591 (N_11591,N_11417,N_11414);
nand U11592 (N_11592,N_11326,N_11338);
xnor U11593 (N_11593,N_11451,N_11405);
and U11594 (N_11594,N_11495,N_11270);
and U11595 (N_11595,N_11397,N_11382);
xor U11596 (N_11596,N_11461,N_11450);
xor U11597 (N_11597,N_11345,N_11296);
or U11598 (N_11598,N_11257,N_11377);
nor U11599 (N_11599,N_11260,N_11490);
nand U11600 (N_11600,N_11458,N_11314);
nand U11601 (N_11601,N_11355,N_11438);
or U11602 (N_11602,N_11250,N_11444);
and U11603 (N_11603,N_11390,N_11308);
nand U11604 (N_11604,N_11389,N_11432);
xnor U11605 (N_11605,N_11447,N_11487);
or U11606 (N_11606,N_11475,N_11488);
or U11607 (N_11607,N_11483,N_11375);
or U11608 (N_11608,N_11262,N_11477);
nor U11609 (N_11609,N_11498,N_11290);
xnor U11610 (N_11610,N_11379,N_11485);
nor U11611 (N_11611,N_11407,N_11410);
nor U11612 (N_11612,N_11365,N_11474);
nor U11613 (N_11613,N_11384,N_11351);
nor U11614 (N_11614,N_11409,N_11364);
xnor U11615 (N_11615,N_11359,N_11452);
nand U11616 (N_11616,N_11276,N_11335);
xnor U11617 (N_11617,N_11318,N_11253);
xor U11618 (N_11618,N_11288,N_11261);
and U11619 (N_11619,N_11259,N_11376);
nor U11620 (N_11620,N_11441,N_11469);
xor U11621 (N_11621,N_11443,N_11395);
nor U11622 (N_11622,N_11289,N_11267);
nand U11623 (N_11623,N_11283,N_11378);
nor U11624 (N_11624,N_11302,N_11281);
nand U11625 (N_11625,N_11337,N_11363);
or U11626 (N_11626,N_11415,N_11393);
or U11627 (N_11627,N_11428,N_11347);
nor U11628 (N_11628,N_11442,N_11276);
and U11629 (N_11629,N_11385,N_11494);
and U11630 (N_11630,N_11322,N_11478);
nor U11631 (N_11631,N_11434,N_11418);
nand U11632 (N_11632,N_11250,N_11369);
xnor U11633 (N_11633,N_11452,N_11318);
xnor U11634 (N_11634,N_11345,N_11469);
nand U11635 (N_11635,N_11456,N_11435);
and U11636 (N_11636,N_11426,N_11474);
nand U11637 (N_11637,N_11304,N_11327);
and U11638 (N_11638,N_11313,N_11461);
nand U11639 (N_11639,N_11251,N_11363);
and U11640 (N_11640,N_11354,N_11254);
nor U11641 (N_11641,N_11309,N_11354);
nand U11642 (N_11642,N_11364,N_11405);
nand U11643 (N_11643,N_11262,N_11320);
nand U11644 (N_11644,N_11312,N_11467);
xnor U11645 (N_11645,N_11484,N_11316);
xnor U11646 (N_11646,N_11310,N_11443);
nand U11647 (N_11647,N_11300,N_11337);
and U11648 (N_11648,N_11407,N_11394);
and U11649 (N_11649,N_11253,N_11315);
xnor U11650 (N_11650,N_11368,N_11372);
and U11651 (N_11651,N_11326,N_11330);
nand U11652 (N_11652,N_11435,N_11491);
xnor U11653 (N_11653,N_11388,N_11471);
xnor U11654 (N_11654,N_11420,N_11335);
xor U11655 (N_11655,N_11435,N_11441);
or U11656 (N_11656,N_11433,N_11356);
nor U11657 (N_11657,N_11476,N_11473);
nor U11658 (N_11658,N_11423,N_11341);
and U11659 (N_11659,N_11334,N_11495);
or U11660 (N_11660,N_11322,N_11274);
nand U11661 (N_11661,N_11311,N_11260);
nand U11662 (N_11662,N_11272,N_11410);
nor U11663 (N_11663,N_11292,N_11266);
nand U11664 (N_11664,N_11420,N_11447);
and U11665 (N_11665,N_11412,N_11336);
nand U11666 (N_11666,N_11477,N_11429);
xor U11667 (N_11667,N_11303,N_11269);
and U11668 (N_11668,N_11250,N_11435);
nor U11669 (N_11669,N_11359,N_11478);
or U11670 (N_11670,N_11337,N_11398);
and U11671 (N_11671,N_11492,N_11420);
nor U11672 (N_11672,N_11482,N_11290);
xor U11673 (N_11673,N_11355,N_11388);
or U11674 (N_11674,N_11392,N_11451);
or U11675 (N_11675,N_11400,N_11303);
and U11676 (N_11676,N_11393,N_11464);
and U11677 (N_11677,N_11353,N_11490);
or U11678 (N_11678,N_11316,N_11327);
nand U11679 (N_11679,N_11420,N_11302);
nor U11680 (N_11680,N_11398,N_11447);
or U11681 (N_11681,N_11276,N_11362);
and U11682 (N_11682,N_11251,N_11426);
xor U11683 (N_11683,N_11384,N_11445);
and U11684 (N_11684,N_11271,N_11402);
nand U11685 (N_11685,N_11325,N_11497);
xnor U11686 (N_11686,N_11436,N_11391);
nand U11687 (N_11687,N_11252,N_11353);
or U11688 (N_11688,N_11430,N_11394);
xnor U11689 (N_11689,N_11468,N_11423);
nor U11690 (N_11690,N_11260,N_11416);
nor U11691 (N_11691,N_11261,N_11359);
nand U11692 (N_11692,N_11462,N_11360);
and U11693 (N_11693,N_11456,N_11368);
xnor U11694 (N_11694,N_11477,N_11435);
xnor U11695 (N_11695,N_11448,N_11258);
nand U11696 (N_11696,N_11403,N_11449);
and U11697 (N_11697,N_11297,N_11496);
xor U11698 (N_11698,N_11351,N_11338);
xnor U11699 (N_11699,N_11481,N_11396);
and U11700 (N_11700,N_11460,N_11333);
nand U11701 (N_11701,N_11331,N_11489);
or U11702 (N_11702,N_11265,N_11384);
and U11703 (N_11703,N_11473,N_11360);
and U11704 (N_11704,N_11420,N_11460);
and U11705 (N_11705,N_11446,N_11427);
nand U11706 (N_11706,N_11280,N_11355);
xor U11707 (N_11707,N_11304,N_11486);
nor U11708 (N_11708,N_11288,N_11406);
or U11709 (N_11709,N_11423,N_11318);
nand U11710 (N_11710,N_11266,N_11305);
nor U11711 (N_11711,N_11466,N_11496);
or U11712 (N_11712,N_11255,N_11281);
or U11713 (N_11713,N_11470,N_11418);
nor U11714 (N_11714,N_11477,N_11389);
nor U11715 (N_11715,N_11356,N_11257);
or U11716 (N_11716,N_11481,N_11451);
and U11717 (N_11717,N_11304,N_11333);
nand U11718 (N_11718,N_11305,N_11398);
nand U11719 (N_11719,N_11470,N_11367);
xnor U11720 (N_11720,N_11311,N_11498);
or U11721 (N_11721,N_11325,N_11472);
xor U11722 (N_11722,N_11251,N_11268);
nor U11723 (N_11723,N_11420,N_11392);
and U11724 (N_11724,N_11421,N_11319);
and U11725 (N_11725,N_11470,N_11313);
xor U11726 (N_11726,N_11491,N_11474);
nor U11727 (N_11727,N_11269,N_11344);
and U11728 (N_11728,N_11472,N_11273);
nand U11729 (N_11729,N_11338,N_11458);
or U11730 (N_11730,N_11493,N_11259);
or U11731 (N_11731,N_11345,N_11262);
and U11732 (N_11732,N_11420,N_11353);
nand U11733 (N_11733,N_11416,N_11328);
and U11734 (N_11734,N_11288,N_11343);
or U11735 (N_11735,N_11372,N_11253);
xor U11736 (N_11736,N_11384,N_11358);
nor U11737 (N_11737,N_11375,N_11462);
or U11738 (N_11738,N_11350,N_11323);
xor U11739 (N_11739,N_11430,N_11457);
and U11740 (N_11740,N_11471,N_11492);
nand U11741 (N_11741,N_11294,N_11463);
or U11742 (N_11742,N_11450,N_11304);
nor U11743 (N_11743,N_11480,N_11349);
or U11744 (N_11744,N_11328,N_11323);
and U11745 (N_11745,N_11404,N_11382);
xnor U11746 (N_11746,N_11426,N_11493);
and U11747 (N_11747,N_11427,N_11276);
and U11748 (N_11748,N_11261,N_11414);
nor U11749 (N_11749,N_11451,N_11484);
nand U11750 (N_11750,N_11720,N_11561);
nor U11751 (N_11751,N_11658,N_11685);
nor U11752 (N_11752,N_11726,N_11701);
nand U11753 (N_11753,N_11553,N_11700);
or U11754 (N_11754,N_11689,N_11715);
and U11755 (N_11755,N_11646,N_11667);
nand U11756 (N_11756,N_11578,N_11501);
and U11757 (N_11757,N_11657,N_11545);
xor U11758 (N_11758,N_11632,N_11599);
nand U11759 (N_11759,N_11623,N_11564);
xnor U11760 (N_11760,N_11555,N_11749);
or U11761 (N_11761,N_11688,N_11741);
nor U11762 (N_11762,N_11571,N_11734);
and U11763 (N_11763,N_11538,N_11626);
xnor U11764 (N_11764,N_11709,N_11573);
nor U11765 (N_11765,N_11562,N_11697);
and U11766 (N_11766,N_11655,N_11597);
nor U11767 (N_11767,N_11733,N_11612);
nand U11768 (N_11768,N_11534,N_11523);
xor U11769 (N_11769,N_11677,N_11542);
and U11770 (N_11770,N_11708,N_11554);
or U11771 (N_11771,N_11508,N_11504);
and U11772 (N_11772,N_11699,N_11662);
xnor U11773 (N_11773,N_11645,N_11625);
nor U11774 (N_11774,N_11724,N_11746);
and U11775 (N_11775,N_11587,N_11703);
xor U11776 (N_11776,N_11702,N_11584);
xor U11777 (N_11777,N_11552,N_11514);
and U11778 (N_11778,N_11540,N_11513);
or U11779 (N_11779,N_11659,N_11560);
nand U11780 (N_11780,N_11500,N_11607);
and U11781 (N_11781,N_11506,N_11649);
nor U11782 (N_11782,N_11704,N_11651);
or U11783 (N_11783,N_11507,N_11574);
nand U11784 (N_11784,N_11664,N_11510);
nor U11785 (N_11785,N_11628,N_11515);
nand U11786 (N_11786,N_11524,N_11682);
xnor U11787 (N_11787,N_11712,N_11647);
nand U11788 (N_11788,N_11743,N_11692);
or U11789 (N_11789,N_11627,N_11648);
and U11790 (N_11790,N_11661,N_11609);
nand U11791 (N_11791,N_11603,N_11557);
or U11792 (N_11792,N_11714,N_11539);
nor U11793 (N_11793,N_11511,N_11517);
or U11794 (N_11794,N_11551,N_11678);
xor U11795 (N_11795,N_11617,N_11739);
and U11796 (N_11796,N_11644,N_11719);
xnor U11797 (N_11797,N_11669,N_11611);
and U11798 (N_11798,N_11532,N_11690);
nand U11799 (N_11799,N_11522,N_11722);
or U11800 (N_11800,N_11681,N_11550);
xnor U11801 (N_11801,N_11585,N_11672);
and U11802 (N_11802,N_11549,N_11530);
or U11803 (N_11803,N_11579,N_11694);
xnor U11804 (N_11804,N_11737,N_11591);
and U11805 (N_11805,N_11503,N_11558);
or U11806 (N_11806,N_11738,N_11728);
xnor U11807 (N_11807,N_11635,N_11721);
nand U11808 (N_11808,N_11680,N_11673);
and U11809 (N_11809,N_11521,N_11636);
and U11810 (N_11810,N_11687,N_11745);
xor U11811 (N_11811,N_11512,N_11605);
nor U11812 (N_11812,N_11706,N_11535);
xnor U11813 (N_11813,N_11653,N_11747);
or U11814 (N_11814,N_11595,N_11616);
and U11815 (N_11815,N_11543,N_11533);
xnor U11816 (N_11816,N_11707,N_11660);
nor U11817 (N_11817,N_11588,N_11637);
and U11818 (N_11818,N_11601,N_11589);
nand U11819 (N_11819,N_11537,N_11686);
and U11820 (N_11820,N_11711,N_11559);
nor U11821 (N_11821,N_11618,N_11520);
and U11822 (N_11822,N_11563,N_11547);
nand U11823 (N_11823,N_11735,N_11619);
or U11824 (N_11824,N_11730,N_11624);
nand U11825 (N_11825,N_11572,N_11602);
and U11826 (N_11826,N_11586,N_11710);
nand U11827 (N_11827,N_11525,N_11548);
nand U11828 (N_11828,N_11568,N_11723);
nand U11829 (N_11829,N_11505,N_11610);
nand U11830 (N_11830,N_11502,N_11717);
or U11831 (N_11831,N_11631,N_11598);
nor U11832 (N_11832,N_11670,N_11725);
nor U11833 (N_11833,N_11736,N_11665);
nor U11834 (N_11834,N_11582,N_11696);
or U11835 (N_11835,N_11519,N_11744);
nand U11836 (N_11836,N_11742,N_11639);
xnor U11837 (N_11837,N_11596,N_11705);
nor U11838 (N_11838,N_11570,N_11622);
nor U11839 (N_11839,N_11693,N_11666);
nand U11840 (N_11840,N_11630,N_11683);
nor U11841 (N_11841,N_11526,N_11629);
or U11842 (N_11842,N_11671,N_11592);
and U11843 (N_11843,N_11620,N_11528);
and U11844 (N_11844,N_11583,N_11727);
nand U11845 (N_11845,N_11748,N_11575);
or U11846 (N_11846,N_11527,N_11529);
nand U11847 (N_11847,N_11518,N_11642);
nor U11848 (N_11848,N_11674,N_11593);
or U11849 (N_11849,N_11641,N_11541);
or U11850 (N_11850,N_11581,N_11600);
xor U11851 (N_11851,N_11684,N_11713);
and U11852 (N_11852,N_11608,N_11732);
or U11853 (N_11853,N_11679,N_11615);
or U11854 (N_11854,N_11676,N_11590);
xor U11855 (N_11855,N_11729,N_11716);
xor U11856 (N_11856,N_11652,N_11531);
and U11857 (N_11857,N_11604,N_11613);
and U11858 (N_11858,N_11509,N_11567);
nor U11859 (N_11859,N_11544,N_11654);
xnor U11860 (N_11860,N_11580,N_11668);
or U11861 (N_11861,N_11576,N_11740);
xnor U11862 (N_11862,N_11566,N_11695);
or U11863 (N_11863,N_11638,N_11546);
nand U11864 (N_11864,N_11569,N_11640);
nand U11865 (N_11865,N_11606,N_11656);
and U11866 (N_11866,N_11633,N_11614);
nand U11867 (N_11867,N_11675,N_11634);
xnor U11868 (N_11868,N_11536,N_11577);
xnor U11869 (N_11869,N_11643,N_11698);
nor U11870 (N_11870,N_11718,N_11565);
xnor U11871 (N_11871,N_11556,N_11621);
nand U11872 (N_11872,N_11516,N_11663);
nor U11873 (N_11873,N_11691,N_11650);
nand U11874 (N_11874,N_11731,N_11594);
nor U11875 (N_11875,N_11645,N_11642);
nor U11876 (N_11876,N_11597,N_11594);
nand U11877 (N_11877,N_11508,N_11608);
and U11878 (N_11878,N_11539,N_11729);
nand U11879 (N_11879,N_11548,N_11614);
xor U11880 (N_11880,N_11550,N_11717);
nand U11881 (N_11881,N_11595,N_11657);
and U11882 (N_11882,N_11692,N_11575);
nor U11883 (N_11883,N_11564,N_11701);
nand U11884 (N_11884,N_11744,N_11717);
or U11885 (N_11885,N_11580,N_11570);
nor U11886 (N_11886,N_11658,N_11544);
nand U11887 (N_11887,N_11715,N_11625);
nand U11888 (N_11888,N_11504,N_11673);
nand U11889 (N_11889,N_11511,N_11696);
xnor U11890 (N_11890,N_11601,N_11596);
or U11891 (N_11891,N_11533,N_11618);
nor U11892 (N_11892,N_11520,N_11617);
and U11893 (N_11893,N_11621,N_11612);
nor U11894 (N_11894,N_11664,N_11636);
or U11895 (N_11895,N_11713,N_11673);
xnor U11896 (N_11896,N_11684,N_11655);
and U11897 (N_11897,N_11743,N_11586);
nor U11898 (N_11898,N_11699,N_11721);
or U11899 (N_11899,N_11588,N_11646);
nor U11900 (N_11900,N_11701,N_11581);
or U11901 (N_11901,N_11619,N_11683);
xnor U11902 (N_11902,N_11641,N_11658);
or U11903 (N_11903,N_11746,N_11550);
nor U11904 (N_11904,N_11612,N_11571);
or U11905 (N_11905,N_11623,N_11566);
or U11906 (N_11906,N_11559,N_11503);
and U11907 (N_11907,N_11525,N_11646);
xnor U11908 (N_11908,N_11612,N_11608);
nand U11909 (N_11909,N_11705,N_11679);
nand U11910 (N_11910,N_11605,N_11648);
xor U11911 (N_11911,N_11718,N_11538);
nand U11912 (N_11912,N_11722,N_11624);
and U11913 (N_11913,N_11543,N_11526);
nand U11914 (N_11914,N_11696,N_11726);
nor U11915 (N_11915,N_11609,N_11622);
or U11916 (N_11916,N_11541,N_11730);
xor U11917 (N_11917,N_11665,N_11670);
and U11918 (N_11918,N_11615,N_11602);
nor U11919 (N_11919,N_11583,N_11642);
or U11920 (N_11920,N_11730,N_11548);
nor U11921 (N_11921,N_11692,N_11606);
and U11922 (N_11922,N_11532,N_11620);
or U11923 (N_11923,N_11669,N_11593);
xor U11924 (N_11924,N_11528,N_11608);
or U11925 (N_11925,N_11617,N_11728);
and U11926 (N_11926,N_11729,N_11650);
xor U11927 (N_11927,N_11603,N_11737);
nand U11928 (N_11928,N_11514,N_11623);
nand U11929 (N_11929,N_11563,N_11697);
and U11930 (N_11930,N_11638,N_11733);
or U11931 (N_11931,N_11549,N_11653);
nor U11932 (N_11932,N_11651,N_11530);
nor U11933 (N_11933,N_11745,N_11698);
xor U11934 (N_11934,N_11516,N_11696);
nor U11935 (N_11935,N_11512,N_11700);
nor U11936 (N_11936,N_11572,N_11725);
xor U11937 (N_11937,N_11651,N_11554);
nor U11938 (N_11938,N_11713,N_11722);
xor U11939 (N_11939,N_11693,N_11692);
xor U11940 (N_11940,N_11561,N_11566);
and U11941 (N_11941,N_11566,N_11529);
nand U11942 (N_11942,N_11558,N_11549);
nand U11943 (N_11943,N_11578,N_11661);
xor U11944 (N_11944,N_11722,N_11580);
nor U11945 (N_11945,N_11730,N_11711);
or U11946 (N_11946,N_11623,N_11708);
xor U11947 (N_11947,N_11539,N_11746);
nand U11948 (N_11948,N_11692,N_11635);
xor U11949 (N_11949,N_11543,N_11514);
or U11950 (N_11950,N_11639,N_11670);
nand U11951 (N_11951,N_11572,N_11581);
and U11952 (N_11952,N_11734,N_11703);
nand U11953 (N_11953,N_11665,N_11590);
xor U11954 (N_11954,N_11523,N_11517);
xor U11955 (N_11955,N_11657,N_11566);
nor U11956 (N_11956,N_11727,N_11573);
xnor U11957 (N_11957,N_11652,N_11739);
and U11958 (N_11958,N_11562,N_11530);
xor U11959 (N_11959,N_11718,N_11518);
nor U11960 (N_11960,N_11711,N_11506);
nand U11961 (N_11961,N_11646,N_11527);
or U11962 (N_11962,N_11699,N_11684);
nand U11963 (N_11963,N_11537,N_11553);
or U11964 (N_11964,N_11546,N_11721);
nand U11965 (N_11965,N_11744,N_11625);
xnor U11966 (N_11966,N_11669,N_11518);
or U11967 (N_11967,N_11547,N_11520);
and U11968 (N_11968,N_11525,N_11628);
xor U11969 (N_11969,N_11630,N_11528);
xnor U11970 (N_11970,N_11681,N_11553);
xor U11971 (N_11971,N_11694,N_11575);
nor U11972 (N_11972,N_11641,N_11723);
xor U11973 (N_11973,N_11732,N_11735);
nand U11974 (N_11974,N_11501,N_11520);
and U11975 (N_11975,N_11596,N_11732);
nor U11976 (N_11976,N_11611,N_11726);
nand U11977 (N_11977,N_11591,N_11604);
nor U11978 (N_11978,N_11692,N_11710);
and U11979 (N_11979,N_11685,N_11559);
or U11980 (N_11980,N_11560,N_11714);
xor U11981 (N_11981,N_11603,N_11685);
xnor U11982 (N_11982,N_11644,N_11640);
and U11983 (N_11983,N_11619,N_11682);
nor U11984 (N_11984,N_11587,N_11607);
or U11985 (N_11985,N_11508,N_11573);
or U11986 (N_11986,N_11723,N_11637);
xnor U11987 (N_11987,N_11720,N_11527);
and U11988 (N_11988,N_11668,N_11627);
or U11989 (N_11989,N_11731,N_11646);
or U11990 (N_11990,N_11666,N_11562);
nand U11991 (N_11991,N_11623,N_11619);
and U11992 (N_11992,N_11530,N_11608);
or U11993 (N_11993,N_11559,N_11594);
or U11994 (N_11994,N_11680,N_11698);
xor U11995 (N_11995,N_11725,N_11630);
nor U11996 (N_11996,N_11706,N_11705);
and U11997 (N_11997,N_11590,N_11646);
or U11998 (N_11998,N_11723,N_11643);
xnor U11999 (N_11999,N_11588,N_11688);
xor U12000 (N_12000,N_11939,N_11905);
xnor U12001 (N_12001,N_11782,N_11924);
and U12002 (N_12002,N_11930,N_11890);
nand U12003 (N_12003,N_11759,N_11994);
and U12004 (N_12004,N_11790,N_11822);
or U12005 (N_12005,N_11838,N_11755);
and U12006 (N_12006,N_11835,N_11891);
and U12007 (N_12007,N_11920,N_11987);
and U12008 (N_12008,N_11981,N_11882);
xor U12009 (N_12009,N_11911,N_11916);
nor U12010 (N_12010,N_11873,N_11840);
xor U12011 (N_12011,N_11927,N_11800);
and U12012 (N_12012,N_11768,N_11899);
or U12013 (N_12013,N_11871,N_11766);
and U12014 (N_12014,N_11964,N_11820);
and U12015 (N_12015,N_11821,N_11763);
or U12016 (N_12016,N_11959,N_11761);
and U12017 (N_12017,N_11764,N_11844);
nor U12018 (N_12018,N_11791,N_11956);
or U12019 (N_12019,N_11945,N_11898);
nor U12020 (N_12020,N_11801,N_11825);
nand U12021 (N_12021,N_11892,N_11885);
nand U12022 (N_12022,N_11843,N_11813);
or U12023 (N_12023,N_11760,N_11807);
xor U12024 (N_12024,N_11826,N_11798);
xnor U12025 (N_12025,N_11802,N_11984);
xor U12026 (N_12026,N_11988,N_11917);
nor U12027 (N_12027,N_11827,N_11823);
and U12028 (N_12028,N_11753,N_11936);
and U12029 (N_12029,N_11864,N_11762);
xor U12030 (N_12030,N_11818,N_11976);
nand U12031 (N_12031,N_11856,N_11922);
nand U12032 (N_12032,N_11793,N_11982);
nand U12033 (N_12033,N_11947,N_11774);
xnor U12034 (N_12034,N_11852,N_11979);
nand U12035 (N_12035,N_11809,N_11817);
and U12036 (N_12036,N_11883,N_11999);
nor U12037 (N_12037,N_11886,N_11859);
and U12038 (N_12038,N_11752,N_11750);
or U12039 (N_12039,N_11880,N_11861);
nand U12040 (N_12040,N_11940,N_11929);
nand U12041 (N_12041,N_11867,N_11879);
or U12042 (N_12042,N_11816,N_11938);
xnor U12043 (N_12043,N_11847,N_11986);
nor U12044 (N_12044,N_11955,N_11837);
nand U12045 (N_12045,N_11773,N_11952);
or U12046 (N_12046,N_11977,N_11975);
and U12047 (N_12047,N_11978,N_11870);
and U12048 (N_12048,N_11908,N_11794);
nand U12049 (N_12049,N_11904,N_11901);
xor U12050 (N_12050,N_11829,N_11912);
and U12051 (N_12051,N_11770,N_11850);
and U12052 (N_12052,N_11784,N_11872);
xor U12053 (N_12053,N_11974,N_11810);
nand U12054 (N_12054,N_11765,N_11799);
and U12055 (N_12055,N_11998,N_11869);
and U12056 (N_12056,N_11878,N_11894);
xnor U12057 (N_12057,N_11913,N_11857);
nor U12058 (N_12058,N_11830,N_11854);
nand U12059 (N_12059,N_11781,N_11767);
xor U12060 (N_12060,N_11933,N_11923);
nand U12061 (N_12061,N_11954,N_11785);
nor U12062 (N_12062,N_11903,N_11973);
xnor U12063 (N_12063,N_11846,N_11941);
nor U12064 (N_12064,N_11960,N_11993);
nor U12065 (N_12065,N_11839,N_11831);
nor U12066 (N_12066,N_11786,N_11983);
nor U12067 (N_12067,N_11797,N_11972);
xnor U12068 (N_12068,N_11966,N_11814);
nand U12069 (N_12069,N_11906,N_11919);
and U12070 (N_12070,N_11851,N_11849);
or U12071 (N_12071,N_11868,N_11990);
or U12072 (N_12072,N_11992,N_11918);
nor U12073 (N_12073,N_11875,N_11946);
nor U12074 (N_12074,N_11949,N_11985);
or U12075 (N_12075,N_11863,N_11787);
nand U12076 (N_12076,N_11937,N_11965);
nand U12077 (N_12077,N_11788,N_11805);
or U12078 (N_12078,N_11848,N_11997);
xor U12079 (N_12079,N_11928,N_11914);
and U12080 (N_12080,N_11777,N_11907);
nor U12081 (N_12081,N_11811,N_11925);
nand U12082 (N_12082,N_11995,N_11775);
or U12083 (N_12083,N_11881,N_11935);
or U12084 (N_12084,N_11970,N_11845);
nand U12085 (N_12085,N_11751,N_11808);
nor U12086 (N_12086,N_11953,N_11833);
nor U12087 (N_12087,N_11803,N_11783);
or U12088 (N_12088,N_11971,N_11932);
xnor U12089 (N_12089,N_11866,N_11860);
or U12090 (N_12090,N_11921,N_11828);
nand U12091 (N_12091,N_11757,N_11944);
nand U12092 (N_12092,N_11934,N_11996);
and U12093 (N_12093,N_11910,N_11895);
and U12094 (N_12094,N_11957,N_11806);
and U12095 (N_12095,N_11961,N_11888);
and U12096 (N_12096,N_11776,N_11884);
nor U12097 (N_12097,N_11874,N_11980);
or U12098 (N_12098,N_11772,N_11769);
nand U12099 (N_12099,N_11841,N_11943);
nand U12100 (N_12100,N_11887,N_11942);
xnor U12101 (N_12101,N_11862,N_11950);
xnor U12102 (N_12102,N_11815,N_11758);
xnor U12103 (N_12103,N_11842,N_11963);
or U12104 (N_12104,N_11780,N_11756);
nand U12105 (N_12105,N_11969,N_11834);
nand U12106 (N_12106,N_11962,N_11836);
and U12107 (N_12107,N_11865,N_11991);
xnor U12108 (N_12108,N_11900,N_11804);
and U12109 (N_12109,N_11779,N_11948);
nor U12110 (N_12110,N_11967,N_11858);
nand U12111 (N_12111,N_11915,N_11771);
xnor U12112 (N_12112,N_11897,N_11889);
nor U12113 (N_12113,N_11796,N_11902);
or U12114 (N_12114,N_11853,N_11876);
or U12115 (N_12115,N_11968,N_11812);
nand U12116 (N_12116,N_11832,N_11951);
and U12117 (N_12117,N_11789,N_11958);
nor U12118 (N_12118,N_11893,N_11877);
xor U12119 (N_12119,N_11989,N_11896);
nor U12120 (N_12120,N_11792,N_11824);
nor U12121 (N_12121,N_11795,N_11754);
xnor U12122 (N_12122,N_11931,N_11926);
nand U12123 (N_12123,N_11819,N_11909);
nor U12124 (N_12124,N_11778,N_11855);
nor U12125 (N_12125,N_11795,N_11993);
or U12126 (N_12126,N_11836,N_11905);
nand U12127 (N_12127,N_11895,N_11841);
and U12128 (N_12128,N_11843,N_11997);
nor U12129 (N_12129,N_11866,N_11883);
or U12130 (N_12130,N_11880,N_11836);
or U12131 (N_12131,N_11812,N_11862);
or U12132 (N_12132,N_11974,N_11793);
xor U12133 (N_12133,N_11762,N_11995);
or U12134 (N_12134,N_11973,N_11792);
xnor U12135 (N_12135,N_11762,N_11902);
xor U12136 (N_12136,N_11760,N_11974);
or U12137 (N_12137,N_11998,N_11813);
xnor U12138 (N_12138,N_11987,N_11764);
nor U12139 (N_12139,N_11774,N_11812);
or U12140 (N_12140,N_11817,N_11767);
xor U12141 (N_12141,N_11928,N_11857);
nor U12142 (N_12142,N_11941,N_11965);
or U12143 (N_12143,N_11929,N_11834);
or U12144 (N_12144,N_11823,N_11915);
nor U12145 (N_12145,N_11859,N_11990);
nor U12146 (N_12146,N_11775,N_11881);
and U12147 (N_12147,N_11769,N_11996);
nand U12148 (N_12148,N_11892,N_11786);
xnor U12149 (N_12149,N_11857,N_11762);
xor U12150 (N_12150,N_11896,N_11978);
nand U12151 (N_12151,N_11874,N_11976);
xor U12152 (N_12152,N_11887,N_11842);
nand U12153 (N_12153,N_11766,N_11855);
nor U12154 (N_12154,N_11966,N_11886);
nand U12155 (N_12155,N_11815,N_11940);
and U12156 (N_12156,N_11795,N_11928);
and U12157 (N_12157,N_11949,N_11880);
nand U12158 (N_12158,N_11921,N_11985);
xnor U12159 (N_12159,N_11968,N_11849);
xnor U12160 (N_12160,N_11754,N_11963);
nor U12161 (N_12161,N_11924,N_11939);
xnor U12162 (N_12162,N_11923,N_11890);
xor U12163 (N_12163,N_11869,N_11949);
or U12164 (N_12164,N_11823,N_11758);
xnor U12165 (N_12165,N_11762,N_11805);
nand U12166 (N_12166,N_11926,N_11798);
or U12167 (N_12167,N_11876,N_11917);
and U12168 (N_12168,N_11919,N_11761);
nor U12169 (N_12169,N_11902,N_11753);
or U12170 (N_12170,N_11790,N_11986);
or U12171 (N_12171,N_11913,N_11989);
or U12172 (N_12172,N_11906,N_11872);
or U12173 (N_12173,N_11955,N_11797);
and U12174 (N_12174,N_11829,N_11826);
or U12175 (N_12175,N_11803,N_11958);
xor U12176 (N_12176,N_11849,N_11975);
nand U12177 (N_12177,N_11932,N_11988);
nand U12178 (N_12178,N_11837,N_11950);
xor U12179 (N_12179,N_11902,N_11997);
or U12180 (N_12180,N_11919,N_11800);
xor U12181 (N_12181,N_11787,N_11840);
xor U12182 (N_12182,N_11758,N_11886);
and U12183 (N_12183,N_11934,N_11902);
and U12184 (N_12184,N_11925,N_11873);
nor U12185 (N_12185,N_11765,N_11900);
nand U12186 (N_12186,N_11948,N_11879);
nand U12187 (N_12187,N_11810,N_11834);
nand U12188 (N_12188,N_11943,N_11905);
nor U12189 (N_12189,N_11879,N_11883);
xor U12190 (N_12190,N_11911,N_11870);
or U12191 (N_12191,N_11888,N_11824);
or U12192 (N_12192,N_11916,N_11985);
nor U12193 (N_12193,N_11772,N_11973);
and U12194 (N_12194,N_11759,N_11809);
nor U12195 (N_12195,N_11782,N_11952);
xor U12196 (N_12196,N_11980,N_11910);
xor U12197 (N_12197,N_11867,N_11969);
xnor U12198 (N_12198,N_11849,N_11985);
xnor U12199 (N_12199,N_11797,N_11771);
nand U12200 (N_12200,N_11965,N_11791);
and U12201 (N_12201,N_11935,N_11897);
xnor U12202 (N_12202,N_11862,N_11949);
and U12203 (N_12203,N_11974,N_11961);
and U12204 (N_12204,N_11925,N_11981);
xor U12205 (N_12205,N_11759,N_11821);
xnor U12206 (N_12206,N_11900,N_11815);
nor U12207 (N_12207,N_11955,N_11859);
and U12208 (N_12208,N_11987,N_11978);
nor U12209 (N_12209,N_11933,N_11857);
xnor U12210 (N_12210,N_11785,N_11752);
and U12211 (N_12211,N_11758,N_11782);
or U12212 (N_12212,N_11779,N_11919);
xor U12213 (N_12213,N_11983,N_11863);
nor U12214 (N_12214,N_11753,N_11860);
and U12215 (N_12215,N_11877,N_11923);
and U12216 (N_12216,N_11921,N_11840);
or U12217 (N_12217,N_11989,N_11981);
or U12218 (N_12218,N_11963,N_11892);
or U12219 (N_12219,N_11863,N_11946);
nand U12220 (N_12220,N_11853,N_11830);
or U12221 (N_12221,N_11874,N_11968);
nand U12222 (N_12222,N_11991,N_11786);
nand U12223 (N_12223,N_11818,N_11766);
nor U12224 (N_12224,N_11802,N_11969);
and U12225 (N_12225,N_11864,N_11969);
or U12226 (N_12226,N_11982,N_11846);
xor U12227 (N_12227,N_11873,N_11879);
nor U12228 (N_12228,N_11856,N_11796);
nand U12229 (N_12229,N_11894,N_11828);
or U12230 (N_12230,N_11944,N_11988);
xor U12231 (N_12231,N_11973,N_11865);
nor U12232 (N_12232,N_11895,N_11989);
nand U12233 (N_12233,N_11785,N_11889);
nor U12234 (N_12234,N_11923,N_11962);
nor U12235 (N_12235,N_11892,N_11777);
nor U12236 (N_12236,N_11844,N_11987);
nand U12237 (N_12237,N_11777,N_11766);
or U12238 (N_12238,N_11984,N_11884);
nand U12239 (N_12239,N_11866,N_11750);
nand U12240 (N_12240,N_11753,N_11851);
and U12241 (N_12241,N_11957,N_11776);
nand U12242 (N_12242,N_11784,N_11907);
xnor U12243 (N_12243,N_11837,N_11880);
or U12244 (N_12244,N_11840,N_11880);
or U12245 (N_12245,N_11785,N_11926);
and U12246 (N_12246,N_11806,N_11824);
nor U12247 (N_12247,N_11857,N_11753);
nor U12248 (N_12248,N_11831,N_11841);
nor U12249 (N_12249,N_11837,N_11865);
nor U12250 (N_12250,N_12038,N_12127);
and U12251 (N_12251,N_12194,N_12035);
xnor U12252 (N_12252,N_12243,N_12148);
nor U12253 (N_12253,N_12019,N_12175);
or U12254 (N_12254,N_12157,N_12152);
and U12255 (N_12255,N_12065,N_12133);
nand U12256 (N_12256,N_12217,N_12197);
nor U12257 (N_12257,N_12205,N_12054);
xor U12258 (N_12258,N_12072,N_12082);
or U12259 (N_12259,N_12031,N_12029);
and U12260 (N_12260,N_12055,N_12006);
or U12261 (N_12261,N_12095,N_12125);
nand U12262 (N_12262,N_12088,N_12172);
and U12263 (N_12263,N_12106,N_12027);
nor U12264 (N_12264,N_12060,N_12211);
xor U12265 (N_12265,N_12110,N_12153);
xnor U12266 (N_12266,N_12118,N_12180);
or U12267 (N_12267,N_12007,N_12092);
nand U12268 (N_12268,N_12015,N_12036);
or U12269 (N_12269,N_12142,N_12238);
or U12270 (N_12270,N_12213,N_12200);
or U12271 (N_12271,N_12132,N_12248);
nor U12272 (N_12272,N_12189,N_12201);
nand U12273 (N_12273,N_12138,N_12062);
nor U12274 (N_12274,N_12212,N_12122);
nand U12275 (N_12275,N_12028,N_12192);
nor U12276 (N_12276,N_12037,N_12024);
nor U12277 (N_12277,N_12202,N_12242);
xnor U12278 (N_12278,N_12168,N_12018);
nor U12279 (N_12279,N_12113,N_12171);
nor U12280 (N_12280,N_12050,N_12186);
xnor U12281 (N_12281,N_12061,N_12160);
xnor U12282 (N_12282,N_12081,N_12043);
and U12283 (N_12283,N_12139,N_12069);
nand U12284 (N_12284,N_12131,N_12239);
or U12285 (N_12285,N_12169,N_12049);
xor U12286 (N_12286,N_12170,N_12178);
xor U12287 (N_12287,N_12047,N_12233);
xnor U12288 (N_12288,N_12078,N_12063);
nor U12289 (N_12289,N_12151,N_12109);
and U12290 (N_12290,N_12058,N_12032);
xor U12291 (N_12291,N_12051,N_12102);
nor U12292 (N_12292,N_12030,N_12022);
or U12293 (N_12293,N_12227,N_12236);
and U12294 (N_12294,N_12206,N_12182);
nor U12295 (N_12295,N_12224,N_12098);
or U12296 (N_12296,N_12231,N_12135);
nand U12297 (N_12297,N_12146,N_12016);
nor U12298 (N_12298,N_12119,N_12101);
or U12299 (N_12299,N_12246,N_12126);
nor U12300 (N_12300,N_12056,N_12225);
nor U12301 (N_12301,N_12164,N_12241);
nor U12302 (N_12302,N_12130,N_12053);
nand U12303 (N_12303,N_12012,N_12108);
or U12304 (N_12304,N_12033,N_12144);
xor U12305 (N_12305,N_12188,N_12103);
or U12306 (N_12306,N_12181,N_12198);
nand U12307 (N_12307,N_12185,N_12222);
and U12308 (N_12308,N_12123,N_12045);
nand U12309 (N_12309,N_12196,N_12026);
nor U12310 (N_12310,N_12093,N_12048);
nor U12311 (N_12311,N_12149,N_12229);
nand U12312 (N_12312,N_12174,N_12204);
nand U12313 (N_12313,N_12064,N_12086);
or U12314 (N_12314,N_12013,N_12021);
xor U12315 (N_12315,N_12041,N_12011);
or U12316 (N_12316,N_12005,N_12116);
nand U12317 (N_12317,N_12025,N_12129);
nor U12318 (N_12318,N_12091,N_12074);
xnor U12319 (N_12319,N_12039,N_12176);
nand U12320 (N_12320,N_12190,N_12218);
nand U12321 (N_12321,N_12134,N_12184);
or U12322 (N_12322,N_12136,N_12140);
xor U12323 (N_12323,N_12166,N_12173);
or U12324 (N_12324,N_12111,N_12216);
or U12325 (N_12325,N_12124,N_12209);
or U12326 (N_12326,N_12014,N_12193);
xnor U12327 (N_12327,N_12099,N_12155);
nor U12328 (N_12328,N_12156,N_12002);
and U12329 (N_12329,N_12097,N_12158);
xnor U12330 (N_12330,N_12040,N_12167);
xor U12331 (N_12331,N_12080,N_12079);
and U12332 (N_12332,N_12208,N_12230);
nand U12333 (N_12333,N_12207,N_12247);
and U12334 (N_12334,N_12219,N_12066);
and U12335 (N_12335,N_12009,N_12187);
xnor U12336 (N_12336,N_12215,N_12141);
nand U12337 (N_12337,N_12143,N_12057);
xor U12338 (N_12338,N_12052,N_12232);
and U12339 (N_12339,N_12010,N_12068);
nand U12340 (N_12340,N_12203,N_12077);
nor U12341 (N_12341,N_12163,N_12100);
and U12342 (N_12342,N_12115,N_12067);
or U12343 (N_12343,N_12071,N_12161);
and U12344 (N_12344,N_12083,N_12183);
nor U12345 (N_12345,N_12165,N_12120);
nor U12346 (N_12346,N_12042,N_12044);
nor U12347 (N_12347,N_12087,N_12112);
and U12348 (N_12348,N_12179,N_12001);
and U12349 (N_12349,N_12128,N_12114);
nor U12350 (N_12350,N_12075,N_12199);
and U12351 (N_12351,N_12023,N_12245);
or U12352 (N_12352,N_12162,N_12000);
nand U12353 (N_12353,N_12220,N_12228);
nand U12354 (N_12354,N_12221,N_12147);
and U12355 (N_12355,N_12145,N_12076);
xor U12356 (N_12356,N_12223,N_12034);
nand U12357 (N_12357,N_12084,N_12214);
or U12358 (N_12358,N_12094,N_12177);
nand U12359 (N_12359,N_12073,N_12090);
xnor U12360 (N_12360,N_12249,N_12150);
nor U12361 (N_12361,N_12195,N_12240);
nor U12362 (N_12362,N_12159,N_12104);
and U12363 (N_12363,N_12226,N_12020);
and U12364 (N_12364,N_12154,N_12105);
and U12365 (N_12365,N_12107,N_12059);
nor U12366 (N_12366,N_12137,N_12004);
or U12367 (N_12367,N_12046,N_12234);
xnor U12368 (N_12368,N_12003,N_12096);
or U12369 (N_12369,N_12244,N_12191);
and U12370 (N_12370,N_12008,N_12017);
nand U12371 (N_12371,N_12089,N_12085);
xor U12372 (N_12372,N_12117,N_12210);
and U12373 (N_12373,N_12070,N_12235);
nor U12374 (N_12374,N_12237,N_12121);
nand U12375 (N_12375,N_12025,N_12075);
nor U12376 (N_12376,N_12204,N_12061);
nand U12377 (N_12377,N_12062,N_12192);
xor U12378 (N_12378,N_12015,N_12035);
nor U12379 (N_12379,N_12175,N_12219);
xor U12380 (N_12380,N_12247,N_12066);
xor U12381 (N_12381,N_12153,N_12135);
nand U12382 (N_12382,N_12098,N_12244);
nand U12383 (N_12383,N_12201,N_12053);
xnor U12384 (N_12384,N_12068,N_12200);
xor U12385 (N_12385,N_12106,N_12209);
or U12386 (N_12386,N_12006,N_12144);
xnor U12387 (N_12387,N_12168,N_12226);
nand U12388 (N_12388,N_12222,N_12221);
nand U12389 (N_12389,N_12078,N_12182);
nor U12390 (N_12390,N_12223,N_12051);
and U12391 (N_12391,N_12067,N_12035);
nand U12392 (N_12392,N_12236,N_12069);
and U12393 (N_12393,N_12039,N_12162);
or U12394 (N_12394,N_12147,N_12152);
nand U12395 (N_12395,N_12206,N_12098);
nand U12396 (N_12396,N_12220,N_12104);
nand U12397 (N_12397,N_12243,N_12064);
and U12398 (N_12398,N_12223,N_12220);
nor U12399 (N_12399,N_12124,N_12037);
or U12400 (N_12400,N_12092,N_12174);
nor U12401 (N_12401,N_12060,N_12241);
nand U12402 (N_12402,N_12070,N_12184);
nand U12403 (N_12403,N_12243,N_12084);
nor U12404 (N_12404,N_12014,N_12024);
xnor U12405 (N_12405,N_12170,N_12145);
xor U12406 (N_12406,N_12029,N_12249);
and U12407 (N_12407,N_12137,N_12099);
xor U12408 (N_12408,N_12040,N_12172);
and U12409 (N_12409,N_12233,N_12158);
nor U12410 (N_12410,N_12068,N_12168);
nand U12411 (N_12411,N_12016,N_12044);
nand U12412 (N_12412,N_12231,N_12065);
nand U12413 (N_12413,N_12242,N_12093);
xor U12414 (N_12414,N_12204,N_12194);
or U12415 (N_12415,N_12040,N_12119);
and U12416 (N_12416,N_12015,N_12237);
nand U12417 (N_12417,N_12126,N_12138);
nor U12418 (N_12418,N_12073,N_12027);
or U12419 (N_12419,N_12042,N_12172);
nor U12420 (N_12420,N_12119,N_12046);
nand U12421 (N_12421,N_12192,N_12210);
or U12422 (N_12422,N_12030,N_12117);
or U12423 (N_12423,N_12124,N_12159);
nor U12424 (N_12424,N_12136,N_12186);
and U12425 (N_12425,N_12044,N_12216);
or U12426 (N_12426,N_12005,N_12214);
nor U12427 (N_12427,N_12040,N_12019);
or U12428 (N_12428,N_12034,N_12092);
xor U12429 (N_12429,N_12083,N_12153);
or U12430 (N_12430,N_12134,N_12081);
and U12431 (N_12431,N_12056,N_12141);
xor U12432 (N_12432,N_12037,N_12081);
xnor U12433 (N_12433,N_12234,N_12237);
xor U12434 (N_12434,N_12188,N_12099);
nor U12435 (N_12435,N_12180,N_12060);
or U12436 (N_12436,N_12208,N_12184);
and U12437 (N_12437,N_12188,N_12125);
xnor U12438 (N_12438,N_12197,N_12234);
nand U12439 (N_12439,N_12021,N_12044);
or U12440 (N_12440,N_12015,N_12146);
nand U12441 (N_12441,N_12042,N_12063);
nand U12442 (N_12442,N_12012,N_12121);
nor U12443 (N_12443,N_12019,N_12079);
xor U12444 (N_12444,N_12234,N_12217);
nor U12445 (N_12445,N_12189,N_12230);
nand U12446 (N_12446,N_12225,N_12222);
and U12447 (N_12447,N_12093,N_12159);
xor U12448 (N_12448,N_12124,N_12106);
nand U12449 (N_12449,N_12090,N_12122);
and U12450 (N_12450,N_12201,N_12058);
nor U12451 (N_12451,N_12068,N_12157);
or U12452 (N_12452,N_12007,N_12137);
or U12453 (N_12453,N_12144,N_12028);
nor U12454 (N_12454,N_12136,N_12121);
and U12455 (N_12455,N_12222,N_12204);
and U12456 (N_12456,N_12052,N_12119);
nand U12457 (N_12457,N_12145,N_12048);
nand U12458 (N_12458,N_12182,N_12060);
and U12459 (N_12459,N_12016,N_12234);
nand U12460 (N_12460,N_12209,N_12064);
xnor U12461 (N_12461,N_12096,N_12012);
nand U12462 (N_12462,N_12107,N_12035);
or U12463 (N_12463,N_12144,N_12031);
xnor U12464 (N_12464,N_12105,N_12179);
or U12465 (N_12465,N_12048,N_12015);
nand U12466 (N_12466,N_12109,N_12087);
nor U12467 (N_12467,N_12082,N_12129);
xor U12468 (N_12468,N_12072,N_12095);
and U12469 (N_12469,N_12054,N_12003);
or U12470 (N_12470,N_12098,N_12147);
and U12471 (N_12471,N_12166,N_12152);
nand U12472 (N_12472,N_12008,N_12149);
nor U12473 (N_12473,N_12230,N_12055);
and U12474 (N_12474,N_12084,N_12195);
or U12475 (N_12475,N_12096,N_12161);
or U12476 (N_12476,N_12199,N_12198);
and U12477 (N_12477,N_12124,N_12242);
nand U12478 (N_12478,N_12180,N_12155);
and U12479 (N_12479,N_12101,N_12221);
xnor U12480 (N_12480,N_12224,N_12144);
xor U12481 (N_12481,N_12047,N_12198);
and U12482 (N_12482,N_12127,N_12196);
nor U12483 (N_12483,N_12240,N_12085);
or U12484 (N_12484,N_12248,N_12107);
xnor U12485 (N_12485,N_12138,N_12151);
xnor U12486 (N_12486,N_12006,N_12045);
nand U12487 (N_12487,N_12013,N_12119);
nor U12488 (N_12488,N_12061,N_12200);
and U12489 (N_12489,N_12078,N_12194);
nor U12490 (N_12490,N_12120,N_12212);
xor U12491 (N_12491,N_12041,N_12060);
nor U12492 (N_12492,N_12007,N_12249);
nor U12493 (N_12493,N_12006,N_12038);
or U12494 (N_12494,N_12211,N_12059);
or U12495 (N_12495,N_12122,N_12220);
nor U12496 (N_12496,N_12087,N_12018);
nor U12497 (N_12497,N_12104,N_12244);
nor U12498 (N_12498,N_12083,N_12236);
or U12499 (N_12499,N_12151,N_12113);
nand U12500 (N_12500,N_12459,N_12452);
or U12501 (N_12501,N_12496,N_12484);
nand U12502 (N_12502,N_12490,N_12485);
nor U12503 (N_12503,N_12364,N_12417);
nor U12504 (N_12504,N_12491,N_12268);
xor U12505 (N_12505,N_12399,N_12285);
and U12506 (N_12506,N_12426,N_12432);
xnor U12507 (N_12507,N_12316,N_12431);
xor U12508 (N_12508,N_12250,N_12380);
xor U12509 (N_12509,N_12407,N_12393);
and U12510 (N_12510,N_12287,N_12466);
or U12511 (N_12511,N_12328,N_12429);
nand U12512 (N_12512,N_12274,N_12296);
or U12513 (N_12513,N_12254,N_12412);
nand U12514 (N_12514,N_12474,N_12333);
xnor U12515 (N_12515,N_12464,N_12303);
nand U12516 (N_12516,N_12427,N_12422);
xnor U12517 (N_12517,N_12355,N_12444);
nand U12518 (N_12518,N_12286,N_12437);
nand U12519 (N_12519,N_12258,N_12343);
nand U12520 (N_12520,N_12414,N_12375);
or U12521 (N_12521,N_12454,N_12483);
or U12522 (N_12522,N_12262,N_12492);
or U12523 (N_12523,N_12310,N_12371);
nand U12524 (N_12524,N_12361,N_12433);
nor U12525 (N_12525,N_12338,N_12356);
nor U12526 (N_12526,N_12261,N_12334);
xnor U12527 (N_12527,N_12379,N_12415);
or U12528 (N_12528,N_12331,N_12383);
xor U12529 (N_12529,N_12386,N_12451);
nor U12530 (N_12530,N_12467,N_12298);
xnor U12531 (N_12531,N_12489,N_12397);
and U12532 (N_12532,N_12322,N_12267);
xnor U12533 (N_12533,N_12295,N_12344);
or U12534 (N_12534,N_12309,N_12275);
nand U12535 (N_12535,N_12456,N_12335);
or U12536 (N_12536,N_12299,N_12480);
and U12537 (N_12537,N_12495,N_12472);
and U12538 (N_12538,N_12291,N_12486);
xnor U12539 (N_12539,N_12403,N_12365);
and U12540 (N_12540,N_12392,N_12266);
nor U12541 (N_12541,N_12277,N_12319);
xor U12542 (N_12542,N_12406,N_12302);
or U12543 (N_12543,N_12455,N_12369);
nor U12544 (N_12544,N_12376,N_12305);
or U12545 (N_12545,N_12499,N_12362);
nor U12546 (N_12546,N_12411,N_12395);
nand U12547 (N_12547,N_12439,N_12493);
nand U12548 (N_12548,N_12280,N_12442);
and U12549 (N_12549,N_12294,N_12256);
and U12550 (N_12550,N_12446,N_12435);
or U12551 (N_12551,N_12325,N_12448);
xor U12552 (N_12552,N_12293,N_12445);
and U12553 (N_12553,N_12388,N_12283);
nor U12554 (N_12554,N_12312,N_12281);
nor U12555 (N_12555,N_12378,N_12471);
and U12556 (N_12556,N_12424,N_12374);
xnor U12557 (N_12557,N_12419,N_12423);
nor U12558 (N_12558,N_12473,N_12428);
xnor U12559 (N_12559,N_12263,N_12479);
nor U12560 (N_12560,N_12272,N_12478);
and U12561 (N_12561,N_12357,N_12438);
or U12562 (N_12562,N_12297,N_12373);
and U12563 (N_12563,N_12271,N_12408);
and U12564 (N_12564,N_12420,N_12337);
nor U12565 (N_12565,N_12264,N_12259);
xnor U12566 (N_12566,N_12385,N_12363);
nand U12567 (N_12567,N_12410,N_12339);
xnor U12568 (N_12568,N_12463,N_12487);
xnor U12569 (N_12569,N_12347,N_12260);
nand U12570 (N_12570,N_12346,N_12488);
and U12571 (N_12571,N_12269,N_12311);
or U12572 (N_12572,N_12358,N_12418);
and U12573 (N_12573,N_12327,N_12436);
and U12574 (N_12574,N_12391,N_12394);
and U12575 (N_12575,N_12306,N_12329);
nor U12576 (N_12576,N_12382,N_12400);
or U12577 (N_12577,N_12323,N_12341);
nor U12578 (N_12578,N_12458,N_12476);
nand U12579 (N_12579,N_12481,N_12387);
nor U12580 (N_12580,N_12255,N_12381);
nand U12581 (N_12581,N_12402,N_12340);
nand U12582 (N_12582,N_12440,N_12308);
xor U12583 (N_12583,N_12318,N_12390);
or U12584 (N_12584,N_12377,N_12320);
nand U12585 (N_12585,N_12300,N_12475);
or U12586 (N_12586,N_12434,N_12430);
or U12587 (N_12587,N_12470,N_12396);
nor U12588 (N_12588,N_12270,N_12352);
xor U12589 (N_12589,N_12497,N_12449);
nor U12590 (N_12590,N_12292,N_12416);
xnor U12591 (N_12591,N_12401,N_12413);
nor U12592 (N_12592,N_12317,N_12313);
xnor U12593 (N_12593,N_12304,N_12450);
nand U12594 (N_12594,N_12389,N_12477);
or U12595 (N_12595,N_12453,N_12350);
or U12596 (N_12596,N_12360,N_12421);
nand U12597 (N_12597,N_12307,N_12368);
nand U12598 (N_12598,N_12290,N_12409);
nand U12599 (N_12599,N_12342,N_12441);
xor U12600 (N_12600,N_12330,N_12469);
xnor U12601 (N_12601,N_12353,N_12354);
nor U12602 (N_12602,N_12443,N_12398);
nand U12603 (N_12603,N_12461,N_12348);
and U12604 (N_12604,N_12252,N_12460);
nand U12605 (N_12605,N_12498,N_12279);
nor U12606 (N_12606,N_12321,N_12253);
and U12607 (N_12607,N_12465,N_12482);
nand U12608 (N_12608,N_12314,N_12332);
nand U12609 (N_12609,N_12447,N_12372);
and U12610 (N_12610,N_12457,N_12289);
and U12611 (N_12611,N_12324,N_12494);
and U12612 (N_12612,N_12276,N_12284);
or U12613 (N_12613,N_12301,N_12351);
or U12614 (N_12614,N_12349,N_12405);
or U12615 (N_12615,N_12462,N_12367);
nor U12616 (N_12616,N_12366,N_12404);
nand U12617 (N_12617,N_12315,N_12326);
and U12618 (N_12618,N_12282,N_12468);
xor U12619 (N_12619,N_12278,N_12265);
and U12620 (N_12620,N_12370,N_12336);
and U12621 (N_12621,N_12288,N_12425);
xnor U12622 (N_12622,N_12273,N_12257);
nor U12623 (N_12623,N_12251,N_12345);
nand U12624 (N_12624,N_12384,N_12359);
nand U12625 (N_12625,N_12322,N_12416);
xor U12626 (N_12626,N_12291,N_12434);
xor U12627 (N_12627,N_12295,N_12393);
xor U12628 (N_12628,N_12424,N_12480);
xor U12629 (N_12629,N_12380,N_12488);
nor U12630 (N_12630,N_12497,N_12478);
and U12631 (N_12631,N_12334,N_12486);
nand U12632 (N_12632,N_12275,N_12354);
and U12633 (N_12633,N_12421,N_12372);
or U12634 (N_12634,N_12389,N_12430);
xor U12635 (N_12635,N_12385,N_12433);
nand U12636 (N_12636,N_12486,N_12451);
xor U12637 (N_12637,N_12318,N_12274);
and U12638 (N_12638,N_12446,N_12452);
xnor U12639 (N_12639,N_12341,N_12481);
or U12640 (N_12640,N_12336,N_12279);
nor U12641 (N_12641,N_12462,N_12296);
xor U12642 (N_12642,N_12350,N_12372);
or U12643 (N_12643,N_12443,N_12487);
xnor U12644 (N_12644,N_12294,N_12305);
nand U12645 (N_12645,N_12444,N_12396);
xor U12646 (N_12646,N_12351,N_12270);
nor U12647 (N_12647,N_12481,N_12323);
nor U12648 (N_12648,N_12342,N_12405);
nand U12649 (N_12649,N_12331,N_12477);
and U12650 (N_12650,N_12409,N_12444);
xnor U12651 (N_12651,N_12333,N_12291);
or U12652 (N_12652,N_12350,N_12263);
nor U12653 (N_12653,N_12268,N_12416);
nor U12654 (N_12654,N_12285,N_12434);
xnor U12655 (N_12655,N_12499,N_12357);
xnor U12656 (N_12656,N_12392,N_12419);
or U12657 (N_12657,N_12414,N_12391);
nor U12658 (N_12658,N_12330,N_12313);
and U12659 (N_12659,N_12296,N_12265);
and U12660 (N_12660,N_12321,N_12395);
nand U12661 (N_12661,N_12415,N_12471);
nor U12662 (N_12662,N_12356,N_12463);
or U12663 (N_12663,N_12369,N_12350);
and U12664 (N_12664,N_12429,N_12431);
nor U12665 (N_12665,N_12376,N_12394);
and U12666 (N_12666,N_12431,N_12402);
and U12667 (N_12667,N_12428,N_12303);
nor U12668 (N_12668,N_12286,N_12463);
or U12669 (N_12669,N_12316,N_12457);
and U12670 (N_12670,N_12444,N_12300);
or U12671 (N_12671,N_12340,N_12417);
xor U12672 (N_12672,N_12395,N_12436);
nor U12673 (N_12673,N_12498,N_12425);
nor U12674 (N_12674,N_12252,N_12255);
xnor U12675 (N_12675,N_12475,N_12389);
xor U12676 (N_12676,N_12264,N_12318);
xnor U12677 (N_12677,N_12281,N_12411);
nor U12678 (N_12678,N_12250,N_12344);
and U12679 (N_12679,N_12480,N_12265);
xnor U12680 (N_12680,N_12452,N_12337);
or U12681 (N_12681,N_12374,N_12311);
nand U12682 (N_12682,N_12379,N_12434);
xnor U12683 (N_12683,N_12412,N_12484);
and U12684 (N_12684,N_12490,N_12352);
xnor U12685 (N_12685,N_12271,N_12350);
nand U12686 (N_12686,N_12262,N_12258);
xor U12687 (N_12687,N_12373,N_12482);
and U12688 (N_12688,N_12337,N_12278);
xor U12689 (N_12689,N_12466,N_12293);
or U12690 (N_12690,N_12498,N_12270);
or U12691 (N_12691,N_12302,N_12445);
or U12692 (N_12692,N_12354,N_12277);
nor U12693 (N_12693,N_12472,N_12316);
xor U12694 (N_12694,N_12267,N_12462);
or U12695 (N_12695,N_12317,N_12272);
or U12696 (N_12696,N_12354,N_12365);
nand U12697 (N_12697,N_12399,N_12419);
or U12698 (N_12698,N_12381,N_12337);
nor U12699 (N_12699,N_12460,N_12315);
xnor U12700 (N_12700,N_12422,N_12267);
nand U12701 (N_12701,N_12272,N_12494);
nand U12702 (N_12702,N_12411,N_12453);
xor U12703 (N_12703,N_12371,N_12358);
nor U12704 (N_12704,N_12262,N_12480);
xor U12705 (N_12705,N_12455,N_12418);
or U12706 (N_12706,N_12384,N_12307);
xor U12707 (N_12707,N_12279,N_12345);
nor U12708 (N_12708,N_12321,N_12380);
xor U12709 (N_12709,N_12442,N_12395);
and U12710 (N_12710,N_12402,N_12474);
xnor U12711 (N_12711,N_12335,N_12296);
and U12712 (N_12712,N_12264,N_12258);
or U12713 (N_12713,N_12444,N_12356);
nand U12714 (N_12714,N_12360,N_12454);
nor U12715 (N_12715,N_12275,N_12355);
nand U12716 (N_12716,N_12305,N_12429);
nand U12717 (N_12717,N_12287,N_12383);
and U12718 (N_12718,N_12473,N_12385);
xnor U12719 (N_12719,N_12405,N_12334);
nor U12720 (N_12720,N_12468,N_12257);
nand U12721 (N_12721,N_12294,N_12365);
nor U12722 (N_12722,N_12367,N_12472);
nand U12723 (N_12723,N_12449,N_12452);
or U12724 (N_12724,N_12330,N_12435);
or U12725 (N_12725,N_12457,N_12402);
nand U12726 (N_12726,N_12299,N_12421);
nand U12727 (N_12727,N_12317,N_12353);
or U12728 (N_12728,N_12330,N_12399);
nor U12729 (N_12729,N_12295,N_12346);
and U12730 (N_12730,N_12306,N_12418);
or U12731 (N_12731,N_12480,N_12317);
nand U12732 (N_12732,N_12277,N_12471);
nor U12733 (N_12733,N_12271,N_12365);
and U12734 (N_12734,N_12295,N_12475);
and U12735 (N_12735,N_12437,N_12440);
nand U12736 (N_12736,N_12312,N_12419);
xnor U12737 (N_12737,N_12258,N_12407);
xnor U12738 (N_12738,N_12329,N_12250);
nor U12739 (N_12739,N_12302,N_12460);
xnor U12740 (N_12740,N_12495,N_12319);
xor U12741 (N_12741,N_12331,N_12452);
nor U12742 (N_12742,N_12444,N_12284);
or U12743 (N_12743,N_12259,N_12418);
xor U12744 (N_12744,N_12374,N_12375);
or U12745 (N_12745,N_12405,N_12424);
and U12746 (N_12746,N_12323,N_12450);
nand U12747 (N_12747,N_12253,N_12415);
and U12748 (N_12748,N_12259,N_12468);
xor U12749 (N_12749,N_12325,N_12476);
xor U12750 (N_12750,N_12633,N_12529);
xor U12751 (N_12751,N_12622,N_12691);
or U12752 (N_12752,N_12611,N_12711);
or U12753 (N_12753,N_12708,N_12664);
xnor U12754 (N_12754,N_12523,N_12697);
and U12755 (N_12755,N_12663,N_12726);
xor U12756 (N_12756,N_12609,N_12583);
or U12757 (N_12757,N_12690,N_12555);
nand U12758 (N_12758,N_12625,N_12548);
and U12759 (N_12759,N_12658,N_12530);
xor U12760 (N_12760,N_12674,N_12508);
xnor U12761 (N_12761,N_12607,N_12531);
and U12762 (N_12762,N_12619,N_12688);
and U12763 (N_12763,N_12541,N_12703);
and U12764 (N_12764,N_12594,N_12603);
nand U12765 (N_12765,N_12687,N_12610);
nand U12766 (N_12766,N_12627,N_12747);
or U12767 (N_12767,N_12665,N_12681);
and U12768 (N_12768,N_12623,N_12510);
xnor U12769 (N_12769,N_12731,N_12519);
xor U12770 (N_12770,N_12706,N_12589);
and U12771 (N_12771,N_12616,N_12536);
or U12772 (N_12772,N_12598,N_12678);
and U12773 (N_12773,N_12542,N_12538);
and U12774 (N_12774,N_12590,N_12582);
xor U12775 (N_12775,N_12528,N_12699);
xor U12776 (N_12776,N_12676,N_12653);
xor U12777 (N_12777,N_12683,N_12596);
and U12778 (N_12778,N_12550,N_12503);
or U12779 (N_12779,N_12651,N_12722);
nor U12780 (N_12780,N_12650,N_12615);
nand U12781 (N_12781,N_12739,N_12670);
nand U12782 (N_12782,N_12709,N_12558);
and U12783 (N_12783,N_12662,N_12743);
nor U12784 (N_12784,N_12626,N_12521);
or U12785 (N_12785,N_12617,N_12715);
and U12786 (N_12786,N_12642,N_12602);
and U12787 (N_12787,N_12639,N_12512);
nand U12788 (N_12788,N_12514,N_12685);
nand U12789 (N_12789,N_12559,N_12571);
or U12790 (N_12790,N_12696,N_12566);
xor U12791 (N_12791,N_12694,N_12608);
and U12792 (N_12792,N_12614,N_12680);
or U12793 (N_12793,N_12587,N_12570);
nand U12794 (N_12794,N_12671,N_12585);
or U12795 (N_12795,N_12723,N_12533);
and U12796 (N_12796,N_12733,N_12544);
nor U12797 (N_12797,N_12576,N_12744);
nand U12798 (N_12798,N_12700,N_12692);
xnor U12799 (N_12799,N_12669,N_12655);
nor U12800 (N_12800,N_12580,N_12612);
nor U12801 (N_12801,N_12600,N_12661);
xnor U12802 (N_12802,N_12727,N_12730);
nand U12803 (N_12803,N_12675,N_12704);
or U12804 (N_12804,N_12535,N_12736);
or U12805 (N_12805,N_12721,N_12748);
nand U12806 (N_12806,N_12673,N_12659);
nor U12807 (N_12807,N_12643,N_12513);
or U12808 (N_12808,N_12527,N_12599);
and U12809 (N_12809,N_12613,N_12562);
nor U12810 (N_12810,N_12644,N_12500);
or U12811 (N_12811,N_12557,N_12672);
or U12812 (N_12812,N_12586,N_12724);
xor U12813 (N_12813,N_12551,N_12720);
xnor U12814 (N_12814,N_12573,N_12537);
xnor U12815 (N_12815,N_12734,N_12705);
xor U12816 (N_12816,N_12618,N_12584);
xnor U12817 (N_12817,N_12595,N_12581);
xnor U12818 (N_12818,N_12682,N_12710);
nand U12819 (N_12819,N_12698,N_12631);
and U12820 (N_12820,N_12725,N_12547);
or U12821 (N_12821,N_12621,N_12501);
and U12822 (N_12822,N_12606,N_12546);
and U12823 (N_12823,N_12568,N_12506);
or U12824 (N_12824,N_12526,N_12677);
and U12825 (N_12825,N_12516,N_12630);
nor U12826 (N_12826,N_12718,N_12738);
xnor U12827 (N_12827,N_12620,N_12684);
or U12828 (N_12828,N_12540,N_12549);
or U12829 (N_12829,N_12657,N_12645);
nand U12830 (N_12830,N_12745,N_12648);
nand U12831 (N_12831,N_12746,N_12660);
xnor U12832 (N_12832,N_12554,N_12686);
and U12833 (N_12833,N_12517,N_12556);
xnor U12834 (N_12834,N_12668,N_12628);
xnor U12835 (N_12835,N_12509,N_12679);
nand U12836 (N_12836,N_12539,N_12532);
xnor U12837 (N_12837,N_12505,N_12564);
or U12838 (N_12838,N_12569,N_12735);
or U12839 (N_12839,N_12629,N_12636);
nor U12840 (N_12840,N_12729,N_12578);
xor U12841 (N_12841,N_12654,N_12565);
and U12842 (N_12842,N_12652,N_12553);
nor U12843 (N_12843,N_12646,N_12597);
or U12844 (N_12844,N_12577,N_12647);
xnor U12845 (N_12845,N_12511,N_12728);
or U12846 (N_12846,N_12716,N_12749);
nor U12847 (N_12847,N_12605,N_12552);
nand U12848 (N_12848,N_12522,N_12632);
or U12849 (N_12849,N_12575,N_12504);
nand U12850 (N_12850,N_12666,N_12579);
nand U12851 (N_12851,N_12635,N_12707);
nand U12852 (N_12852,N_12637,N_12534);
or U12853 (N_12853,N_12714,N_12701);
nand U12854 (N_12854,N_12561,N_12740);
or U12855 (N_12855,N_12717,N_12567);
xor U12856 (N_12856,N_12667,N_12737);
xor U12857 (N_12857,N_12574,N_12640);
or U12858 (N_12858,N_12591,N_12638);
and U12859 (N_12859,N_12588,N_12713);
and U12860 (N_12860,N_12712,N_12520);
nor U12861 (N_12861,N_12507,N_12502);
nand U12862 (N_12862,N_12545,N_12592);
xnor U12863 (N_12863,N_12695,N_12742);
and U12864 (N_12864,N_12702,N_12593);
nand U12865 (N_12865,N_12543,N_12563);
xnor U12866 (N_12866,N_12732,N_12604);
nand U12867 (N_12867,N_12689,N_12518);
nor U12868 (N_12868,N_12560,N_12649);
and U12869 (N_12869,N_12741,N_12634);
nand U12870 (N_12870,N_12656,N_12524);
and U12871 (N_12871,N_12624,N_12525);
xnor U12872 (N_12872,N_12515,N_12572);
xnor U12873 (N_12873,N_12601,N_12719);
nand U12874 (N_12874,N_12641,N_12693);
nor U12875 (N_12875,N_12514,N_12687);
nand U12876 (N_12876,N_12641,N_12684);
and U12877 (N_12877,N_12594,N_12572);
nand U12878 (N_12878,N_12605,N_12536);
or U12879 (N_12879,N_12657,N_12693);
nand U12880 (N_12880,N_12659,N_12582);
or U12881 (N_12881,N_12740,N_12582);
xor U12882 (N_12882,N_12509,N_12625);
nor U12883 (N_12883,N_12633,N_12596);
or U12884 (N_12884,N_12646,N_12541);
xor U12885 (N_12885,N_12588,N_12543);
or U12886 (N_12886,N_12599,N_12509);
and U12887 (N_12887,N_12542,N_12700);
or U12888 (N_12888,N_12611,N_12719);
nand U12889 (N_12889,N_12606,N_12518);
xnor U12890 (N_12890,N_12574,N_12628);
nand U12891 (N_12891,N_12715,N_12635);
nor U12892 (N_12892,N_12696,N_12642);
or U12893 (N_12893,N_12585,N_12651);
and U12894 (N_12894,N_12695,N_12673);
and U12895 (N_12895,N_12549,N_12738);
or U12896 (N_12896,N_12694,N_12580);
xor U12897 (N_12897,N_12714,N_12729);
nor U12898 (N_12898,N_12567,N_12628);
and U12899 (N_12899,N_12617,N_12719);
nand U12900 (N_12900,N_12725,N_12721);
xnor U12901 (N_12901,N_12629,N_12563);
and U12902 (N_12902,N_12732,N_12652);
nor U12903 (N_12903,N_12745,N_12576);
nor U12904 (N_12904,N_12709,N_12542);
nor U12905 (N_12905,N_12600,N_12657);
and U12906 (N_12906,N_12514,N_12621);
and U12907 (N_12907,N_12528,N_12715);
xor U12908 (N_12908,N_12705,N_12673);
or U12909 (N_12909,N_12556,N_12680);
or U12910 (N_12910,N_12707,N_12638);
nand U12911 (N_12911,N_12746,N_12585);
nor U12912 (N_12912,N_12521,N_12703);
or U12913 (N_12913,N_12583,N_12561);
and U12914 (N_12914,N_12651,N_12600);
nor U12915 (N_12915,N_12731,N_12532);
nor U12916 (N_12916,N_12713,N_12617);
or U12917 (N_12917,N_12682,N_12622);
and U12918 (N_12918,N_12500,N_12556);
xnor U12919 (N_12919,N_12628,N_12641);
and U12920 (N_12920,N_12722,N_12554);
or U12921 (N_12921,N_12618,N_12685);
xnor U12922 (N_12922,N_12585,N_12697);
xnor U12923 (N_12923,N_12691,N_12561);
xnor U12924 (N_12924,N_12673,N_12661);
or U12925 (N_12925,N_12627,N_12566);
nand U12926 (N_12926,N_12535,N_12562);
nand U12927 (N_12927,N_12538,N_12622);
nor U12928 (N_12928,N_12529,N_12735);
or U12929 (N_12929,N_12518,N_12545);
or U12930 (N_12930,N_12715,N_12533);
or U12931 (N_12931,N_12705,N_12522);
or U12932 (N_12932,N_12614,N_12502);
or U12933 (N_12933,N_12679,N_12577);
xnor U12934 (N_12934,N_12532,N_12502);
nand U12935 (N_12935,N_12651,N_12557);
and U12936 (N_12936,N_12722,N_12670);
nor U12937 (N_12937,N_12547,N_12620);
nand U12938 (N_12938,N_12581,N_12718);
xor U12939 (N_12939,N_12657,N_12570);
nor U12940 (N_12940,N_12561,N_12606);
and U12941 (N_12941,N_12523,N_12533);
xnor U12942 (N_12942,N_12735,N_12644);
nor U12943 (N_12943,N_12620,N_12694);
and U12944 (N_12944,N_12602,N_12681);
nand U12945 (N_12945,N_12539,N_12559);
nor U12946 (N_12946,N_12641,N_12614);
and U12947 (N_12947,N_12534,N_12666);
nand U12948 (N_12948,N_12744,N_12505);
nor U12949 (N_12949,N_12509,N_12640);
and U12950 (N_12950,N_12594,N_12524);
xnor U12951 (N_12951,N_12741,N_12626);
or U12952 (N_12952,N_12540,N_12736);
nor U12953 (N_12953,N_12681,N_12534);
xnor U12954 (N_12954,N_12726,N_12673);
and U12955 (N_12955,N_12689,N_12521);
nor U12956 (N_12956,N_12644,N_12661);
nor U12957 (N_12957,N_12629,N_12654);
xnor U12958 (N_12958,N_12712,N_12606);
nor U12959 (N_12959,N_12698,N_12704);
nor U12960 (N_12960,N_12742,N_12667);
xnor U12961 (N_12961,N_12688,N_12646);
nor U12962 (N_12962,N_12529,N_12640);
xor U12963 (N_12963,N_12575,N_12599);
and U12964 (N_12964,N_12583,N_12518);
nor U12965 (N_12965,N_12592,N_12589);
or U12966 (N_12966,N_12684,N_12582);
and U12967 (N_12967,N_12689,N_12516);
nand U12968 (N_12968,N_12627,N_12634);
nand U12969 (N_12969,N_12645,N_12519);
xnor U12970 (N_12970,N_12740,N_12587);
nand U12971 (N_12971,N_12569,N_12711);
xnor U12972 (N_12972,N_12587,N_12641);
and U12973 (N_12973,N_12517,N_12745);
xor U12974 (N_12974,N_12636,N_12747);
xor U12975 (N_12975,N_12502,N_12595);
and U12976 (N_12976,N_12559,N_12573);
nor U12977 (N_12977,N_12613,N_12731);
and U12978 (N_12978,N_12632,N_12648);
nor U12979 (N_12979,N_12504,N_12550);
nor U12980 (N_12980,N_12727,N_12543);
xnor U12981 (N_12981,N_12672,N_12652);
and U12982 (N_12982,N_12682,N_12731);
nor U12983 (N_12983,N_12598,N_12715);
and U12984 (N_12984,N_12732,N_12746);
xnor U12985 (N_12985,N_12725,N_12552);
nor U12986 (N_12986,N_12748,N_12681);
nor U12987 (N_12987,N_12645,N_12514);
and U12988 (N_12988,N_12510,N_12512);
nand U12989 (N_12989,N_12520,N_12570);
nand U12990 (N_12990,N_12734,N_12545);
or U12991 (N_12991,N_12724,N_12614);
or U12992 (N_12992,N_12621,N_12549);
nand U12993 (N_12993,N_12531,N_12695);
nor U12994 (N_12994,N_12673,N_12644);
nor U12995 (N_12995,N_12705,N_12685);
xor U12996 (N_12996,N_12691,N_12688);
xnor U12997 (N_12997,N_12664,N_12624);
nand U12998 (N_12998,N_12621,N_12711);
nand U12999 (N_12999,N_12719,N_12650);
xnor U13000 (N_13000,N_12830,N_12984);
or U13001 (N_13001,N_12951,N_12917);
xnor U13002 (N_13002,N_12787,N_12990);
nand U13003 (N_13003,N_12964,N_12821);
nor U13004 (N_13004,N_12818,N_12934);
or U13005 (N_13005,N_12947,N_12762);
nand U13006 (N_13006,N_12799,N_12824);
nor U13007 (N_13007,N_12876,N_12784);
or U13008 (N_13008,N_12781,N_12809);
and U13009 (N_13009,N_12893,N_12761);
xor U13010 (N_13010,N_12974,N_12980);
and U13011 (N_13011,N_12801,N_12771);
xnor U13012 (N_13012,N_12930,N_12849);
nand U13013 (N_13013,N_12802,N_12856);
nor U13014 (N_13014,N_12832,N_12941);
xor U13015 (N_13015,N_12891,N_12985);
nor U13016 (N_13016,N_12775,N_12776);
nand U13017 (N_13017,N_12932,N_12872);
nand U13018 (N_13018,N_12826,N_12953);
nand U13019 (N_13019,N_12966,N_12791);
nand U13020 (N_13020,N_12827,N_12940);
xnor U13021 (N_13021,N_12883,N_12925);
nor U13022 (N_13022,N_12845,N_12797);
nand U13023 (N_13023,N_12905,N_12881);
nand U13024 (N_13024,N_12897,N_12913);
nand U13025 (N_13025,N_12770,N_12839);
xor U13026 (N_13026,N_12877,N_12848);
and U13027 (N_13027,N_12935,N_12789);
nand U13028 (N_13028,N_12973,N_12998);
xor U13029 (N_13029,N_12810,N_12918);
or U13030 (N_13030,N_12769,N_12751);
nand U13031 (N_13031,N_12972,N_12907);
xnor U13032 (N_13032,N_12971,N_12884);
nand U13033 (N_13033,N_12798,N_12928);
and U13034 (N_13034,N_12960,N_12949);
and U13035 (N_13035,N_12785,N_12926);
or U13036 (N_13036,N_12908,N_12773);
and U13037 (N_13037,N_12921,N_12874);
nand U13038 (N_13038,N_12803,N_12774);
nand U13039 (N_13039,N_12860,N_12898);
and U13040 (N_13040,N_12983,N_12814);
xnor U13041 (N_13041,N_12887,N_12987);
xnor U13042 (N_13042,N_12758,N_12844);
and U13043 (N_13043,N_12914,N_12952);
or U13044 (N_13044,N_12796,N_12944);
and U13045 (N_13045,N_12836,N_12833);
xnor U13046 (N_13046,N_12764,N_12962);
nor U13047 (N_13047,N_12878,N_12882);
xnor U13048 (N_13048,N_12869,N_12841);
nand U13049 (N_13049,N_12837,N_12904);
nand U13050 (N_13050,N_12923,N_12950);
nand U13051 (N_13051,N_12939,N_12788);
nand U13052 (N_13052,N_12760,N_12819);
or U13053 (N_13053,N_12942,N_12880);
nor U13054 (N_13054,N_12840,N_12790);
nor U13055 (N_13055,N_12992,N_12910);
nor U13056 (N_13056,N_12865,N_12954);
nand U13057 (N_13057,N_12995,N_12823);
xnor U13058 (N_13058,N_12864,N_12922);
nor U13059 (N_13059,N_12975,N_12750);
xor U13060 (N_13060,N_12871,N_12970);
or U13061 (N_13061,N_12831,N_12903);
nand U13062 (N_13062,N_12912,N_12936);
and U13063 (N_13063,N_12779,N_12828);
and U13064 (N_13064,N_12806,N_12804);
nor U13065 (N_13065,N_12780,N_12755);
nand U13066 (N_13066,N_12994,N_12902);
xor U13067 (N_13067,N_12885,N_12817);
and U13068 (N_13068,N_12782,N_12858);
and U13069 (N_13069,N_12896,N_12768);
and U13070 (N_13070,N_12899,N_12752);
nand U13071 (N_13071,N_12900,N_12997);
or U13072 (N_13072,N_12846,N_12948);
nand U13073 (N_13073,N_12868,N_12906);
xnor U13074 (N_13074,N_12759,N_12820);
nor U13075 (N_13075,N_12777,N_12863);
nor U13076 (N_13076,N_12870,N_12911);
or U13077 (N_13077,N_12958,N_12772);
nor U13078 (N_13078,N_12886,N_12982);
nor U13079 (N_13079,N_12875,N_12786);
nor U13080 (N_13080,N_12978,N_12757);
xnor U13081 (N_13081,N_12976,N_12853);
nand U13082 (N_13082,N_12927,N_12961);
xor U13083 (N_13083,N_12919,N_12873);
nand U13084 (N_13084,N_12816,N_12901);
xnor U13085 (N_13085,N_12767,N_12879);
nor U13086 (N_13086,N_12993,N_12959);
or U13087 (N_13087,N_12800,N_12920);
xor U13088 (N_13088,N_12909,N_12890);
and U13089 (N_13089,N_12945,N_12999);
xnor U13090 (N_13090,N_12829,N_12867);
xnor U13091 (N_13091,N_12924,N_12822);
nand U13092 (N_13092,N_12979,N_12929);
nand U13093 (N_13093,N_12812,N_12847);
nor U13094 (N_13094,N_12965,N_12756);
xnor U13095 (N_13095,N_12857,N_12811);
xor U13096 (N_13096,N_12783,N_12895);
or U13097 (N_13097,N_12946,N_12795);
or U13098 (N_13098,N_12838,N_12753);
nand U13099 (N_13099,N_12859,N_12843);
or U13100 (N_13100,N_12861,N_12937);
xnor U13101 (N_13101,N_12807,N_12989);
nand U13102 (N_13102,N_12852,N_12825);
nand U13103 (N_13103,N_12834,N_12805);
nor U13104 (N_13104,N_12792,N_12778);
xnor U13105 (N_13105,N_12991,N_12808);
xor U13106 (N_13106,N_12854,N_12938);
or U13107 (N_13107,N_12815,N_12986);
xnor U13108 (N_13108,N_12754,N_12855);
xor U13109 (N_13109,N_12842,N_12977);
and U13110 (N_13110,N_12969,N_12793);
and U13111 (N_13111,N_12916,N_12894);
nor U13112 (N_13112,N_12835,N_12943);
and U13113 (N_13113,N_12956,N_12931);
nor U13114 (N_13114,N_12996,N_12933);
xnor U13115 (N_13115,N_12967,N_12968);
and U13116 (N_13116,N_12889,N_12851);
nor U13117 (N_13117,N_12892,N_12955);
xnor U13118 (N_13118,N_12988,N_12766);
nand U13119 (N_13119,N_12763,N_12850);
and U13120 (N_13120,N_12765,N_12915);
nor U13121 (N_13121,N_12981,N_12888);
nor U13122 (N_13122,N_12794,N_12862);
nor U13123 (N_13123,N_12866,N_12957);
nor U13124 (N_13124,N_12813,N_12963);
xor U13125 (N_13125,N_12853,N_12825);
nand U13126 (N_13126,N_12838,N_12980);
nand U13127 (N_13127,N_12871,N_12978);
xor U13128 (N_13128,N_12880,N_12852);
and U13129 (N_13129,N_12939,N_12883);
or U13130 (N_13130,N_12751,N_12773);
or U13131 (N_13131,N_12779,N_12932);
nand U13132 (N_13132,N_12750,N_12816);
and U13133 (N_13133,N_12819,N_12954);
xnor U13134 (N_13134,N_12843,N_12901);
and U13135 (N_13135,N_12757,N_12761);
nand U13136 (N_13136,N_12996,N_12953);
nor U13137 (N_13137,N_12940,N_12837);
or U13138 (N_13138,N_12821,N_12782);
xnor U13139 (N_13139,N_12946,N_12768);
nand U13140 (N_13140,N_12837,N_12793);
nand U13141 (N_13141,N_12926,N_12968);
xnor U13142 (N_13142,N_12842,N_12991);
or U13143 (N_13143,N_12983,N_12991);
xnor U13144 (N_13144,N_12830,N_12758);
xor U13145 (N_13145,N_12789,N_12827);
xnor U13146 (N_13146,N_12786,N_12880);
xor U13147 (N_13147,N_12905,N_12788);
nand U13148 (N_13148,N_12839,N_12964);
xnor U13149 (N_13149,N_12893,N_12786);
or U13150 (N_13150,N_12929,N_12846);
nor U13151 (N_13151,N_12975,N_12871);
xor U13152 (N_13152,N_12851,N_12778);
xnor U13153 (N_13153,N_12884,N_12953);
and U13154 (N_13154,N_12813,N_12823);
and U13155 (N_13155,N_12990,N_12903);
xnor U13156 (N_13156,N_12794,N_12839);
xor U13157 (N_13157,N_12874,N_12888);
or U13158 (N_13158,N_12856,N_12919);
xnor U13159 (N_13159,N_12997,N_12820);
nand U13160 (N_13160,N_12965,N_12893);
nand U13161 (N_13161,N_12762,N_12933);
nor U13162 (N_13162,N_12877,N_12883);
nor U13163 (N_13163,N_12846,N_12898);
nand U13164 (N_13164,N_12813,N_12888);
and U13165 (N_13165,N_12959,N_12919);
or U13166 (N_13166,N_12782,N_12914);
or U13167 (N_13167,N_12874,N_12814);
or U13168 (N_13168,N_12862,N_12886);
xnor U13169 (N_13169,N_12824,N_12907);
xor U13170 (N_13170,N_12966,N_12954);
nor U13171 (N_13171,N_12803,N_12901);
nor U13172 (N_13172,N_12836,N_12852);
xor U13173 (N_13173,N_12912,N_12872);
nand U13174 (N_13174,N_12878,N_12994);
and U13175 (N_13175,N_12914,N_12937);
xor U13176 (N_13176,N_12868,N_12756);
nor U13177 (N_13177,N_12995,N_12793);
or U13178 (N_13178,N_12815,N_12854);
nor U13179 (N_13179,N_12821,N_12999);
xnor U13180 (N_13180,N_12882,N_12989);
and U13181 (N_13181,N_12830,N_12757);
xor U13182 (N_13182,N_12913,N_12886);
xnor U13183 (N_13183,N_12845,N_12894);
or U13184 (N_13184,N_12937,N_12923);
xor U13185 (N_13185,N_12939,N_12841);
xnor U13186 (N_13186,N_12996,N_12803);
nor U13187 (N_13187,N_12824,N_12976);
xnor U13188 (N_13188,N_12958,N_12933);
and U13189 (N_13189,N_12856,N_12986);
or U13190 (N_13190,N_12996,N_12955);
xor U13191 (N_13191,N_12919,N_12774);
or U13192 (N_13192,N_12759,N_12854);
or U13193 (N_13193,N_12922,N_12965);
xor U13194 (N_13194,N_12844,N_12843);
and U13195 (N_13195,N_12947,N_12942);
or U13196 (N_13196,N_12921,N_12846);
nor U13197 (N_13197,N_12826,N_12942);
nor U13198 (N_13198,N_12791,N_12879);
nand U13199 (N_13199,N_12820,N_12907);
xor U13200 (N_13200,N_12760,N_12992);
and U13201 (N_13201,N_12958,N_12904);
and U13202 (N_13202,N_12916,N_12793);
nand U13203 (N_13203,N_12796,N_12854);
xor U13204 (N_13204,N_12964,N_12934);
nand U13205 (N_13205,N_12849,N_12875);
or U13206 (N_13206,N_12835,N_12972);
nor U13207 (N_13207,N_12911,N_12857);
nand U13208 (N_13208,N_12944,N_12841);
nor U13209 (N_13209,N_12761,N_12824);
xnor U13210 (N_13210,N_12987,N_12755);
xor U13211 (N_13211,N_12777,N_12911);
nand U13212 (N_13212,N_12764,N_12923);
and U13213 (N_13213,N_12774,N_12785);
xor U13214 (N_13214,N_12793,N_12972);
xor U13215 (N_13215,N_12807,N_12802);
xor U13216 (N_13216,N_12838,N_12993);
xnor U13217 (N_13217,N_12808,N_12990);
xor U13218 (N_13218,N_12985,N_12835);
nor U13219 (N_13219,N_12941,N_12961);
xnor U13220 (N_13220,N_12887,N_12895);
or U13221 (N_13221,N_12808,N_12974);
xnor U13222 (N_13222,N_12944,N_12822);
nand U13223 (N_13223,N_12998,N_12886);
nor U13224 (N_13224,N_12927,N_12783);
xor U13225 (N_13225,N_12763,N_12780);
and U13226 (N_13226,N_12788,N_12754);
and U13227 (N_13227,N_12774,N_12899);
nor U13228 (N_13228,N_12823,N_12952);
nand U13229 (N_13229,N_12946,N_12822);
and U13230 (N_13230,N_12937,N_12892);
xnor U13231 (N_13231,N_12960,N_12763);
or U13232 (N_13232,N_12836,N_12840);
nor U13233 (N_13233,N_12999,N_12890);
nor U13234 (N_13234,N_12968,N_12939);
xnor U13235 (N_13235,N_12913,N_12816);
nor U13236 (N_13236,N_12760,N_12806);
nor U13237 (N_13237,N_12986,N_12885);
and U13238 (N_13238,N_12866,N_12823);
xor U13239 (N_13239,N_12981,N_12908);
nor U13240 (N_13240,N_12975,N_12955);
or U13241 (N_13241,N_12863,N_12881);
or U13242 (N_13242,N_12797,N_12904);
and U13243 (N_13243,N_12978,N_12846);
and U13244 (N_13244,N_12752,N_12796);
nor U13245 (N_13245,N_12908,N_12759);
nor U13246 (N_13246,N_12801,N_12911);
nand U13247 (N_13247,N_12929,N_12837);
or U13248 (N_13248,N_12872,N_12981);
nor U13249 (N_13249,N_12917,N_12932);
xor U13250 (N_13250,N_13072,N_13167);
xor U13251 (N_13251,N_13173,N_13092);
nor U13252 (N_13252,N_13114,N_13018);
nand U13253 (N_13253,N_13143,N_13170);
and U13254 (N_13254,N_13098,N_13206);
nor U13255 (N_13255,N_13148,N_13020);
or U13256 (N_13256,N_13154,N_13108);
and U13257 (N_13257,N_13125,N_13116);
nand U13258 (N_13258,N_13014,N_13202);
or U13259 (N_13259,N_13063,N_13193);
xnor U13260 (N_13260,N_13045,N_13019);
nand U13261 (N_13261,N_13142,N_13231);
xor U13262 (N_13262,N_13129,N_13022);
or U13263 (N_13263,N_13100,N_13248);
nor U13264 (N_13264,N_13032,N_13039);
xnor U13265 (N_13265,N_13210,N_13025);
xnor U13266 (N_13266,N_13091,N_13223);
nor U13267 (N_13267,N_13102,N_13026);
or U13268 (N_13268,N_13205,N_13106);
nor U13269 (N_13269,N_13049,N_13064);
and U13270 (N_13270,N_13220,N_13186);
or U13271 (N_13271,N_13191,N_13222);
or U13272 (N_13272,N_13164,N_13194);
xnor U13273 (N_13273,N_13077,N_13118);
xnor U13274 (N_13274,N_13126,N_13141);
nor U13275 (N_13275,N_13239,N_13120);
nand U13276 (N_13276,N_13041,N_13089);
nor U13277 (N_13277,N_13134,N_13009);
or U13278 (N_13278,N_13211,N_13216);
nand U13279 (N_13279,N_13030,N_13152);
xnor U13280 (N_13280,N_13215,N_13068);
and U13281 (N_13281,N_13157,N_13035);
nor U13282 (N_13282,N_13112,N_13228);
nor U13283 (N_13283,N_13247,N_13158);
nand U13284 (N_13284,N_13123,N_13176);
nor U13285 (N_13285,N_13209,N_13015);
nand U13286 (N_13286,N_13117,N_13055);
and U13287 (N_13287,N_13136,N_13227);
nor U13288 (N_13288,N_13048,N_13180);
nand U13289 (N_13289,N_13096,N_13185);
nand U13290 (N_13290,N_13017,N_13175);
nor U13291 (N_13291,N_13007,N_13225);
or U13292 (N_13292,N_13047,N_13240);
nand U13293 (N_13293,N_13145,N_13012);
and U13294 (N_13294,N_13011,N_13031);
or U13295 (N_13295,N_13213,N_13188);
nand U13296 (N_13296,N_13084,N_13044);
or U13297 (N_13297,N_13065,N_13082);
nand U13298 (N_13298,N_13107,N_13203);
nor U13299 (N_13299,N_13110,N_13199);
xnor U13300 (N_13300,N_13241,N_13121);
and U13301 (N_13301,N_13172,N_13128);
nor U13302 (N_13302,N_13074,N_13224);
and U13303 (N_13303,N_13062,N_13200);
and U13304 (N_13304,N_13183,N_13001);
nand U13305 (N_13305,N_13027,N_13171);
nand U13306 (N_13306,N_13060,N_13093);
nor U13307 (N_13307,N_13156,N_13086);
nand U13308 (N_13308,N_13088,N_13005);
and U13309 (N_13309,N_13137,N_13085);
nand U13310 (N_13310,N_13103,N_13124);
xor U13311 (N_13311,N_13201,N_13232);
xnor U13312 (N_13312,N_13021,N_13204);
and U13313 (N_13313,N_13003,N_13073);
and U13314 (N_13314,N_13040,N_13132);
nor U13315 (N_13315,N_13138,N_13244);
nand U13316 (N_13316,N_13246,N_13229);
xor U13317 (N_13317,N_13008,N_13029);
xnor U13318 (N_13318,N_13174,N_13245);
or U13319 (N_13319,N_13097,N_13131);
xor U13320 (N_13320,N_13067,N_13076);
xnor U13321 (N_13321,N_13002,N_13161);
nand U13322 (N_13322,N_13000,N_13197);
nand U13323 (N_13323,N_13184,N_13198);
and U13324 (N_13324,N_13237,N_13218);
or U13325 (N_13325,N_13070,N_13160);
nand U13326 (N_13326,N_13178,N_13075);
and U13327 (N_13327,N_13033,N_13207);
nor U13328 (N_13328,N_13226,N_13046);
nor U13329 (N_13329,N_13155,N_13151);
xnor U13330 (N_13330,N_13150,N_13105);
and U13331 (N_13331,N_13036,N_13187);
nand U13332 (N_13332,N_13104,N_13140);
or U13333 (N_13333,N_13119,N_13006);
nand U13334 (N_13334,N_13249,N_13080);
xor U13335 (N_13335,N_13052,N_13078);
nand U13336 (N_13336,N_13234,N_13190);
or U13337 (N_13337,N_13168,N_13004);
or U13338 (N_13338,N_13010,N_13149);
nor U13339 (N_13339,N_13056,N_13037);
or U13340 (N_13340,N_13057,N_13162);
nor U13341 (N_13341,N_13212,N_13139);
or U13342 (N_13342,N_13179,N_13111);
and U13343 (N_13343,N_13230,N_13053);
xnor U13344 (N_13344,N_13133,N_13034);
or U13345 (N_13345,N_13066,N_13233);
nand U13346 (N_13346,N_13109,N_13189);
xor U13347 (N_13347,N_13169,N_13028);
or U13348 (N_13348,N_13165,N_13113);
nand U13349 (N_13349,N_13196,N_13051);
or U13350 (N_13350,N_13221,N_13115);
xnor U13351 (N_13351,N_13024,N_13130);
xnor U13352 (N_13352,N_13094,N_13192);
nor U13353 (N_13353,N_13050,N_13087);
and U13354 (N_13354,N_13090,N_13016);
xnor U13355 (N_13355,N_13127,N_13147);
nand U13356 (N_13356,N_13058,N_13043);
nor U13357 (N_13357,N_13054,N_13195);
xor U13358 (N_13358,N_13235,N_13081);
nand U13359 (N_13359,N_13079,N_13023);
nor U13360 (N_13360,N_13182,N_13242);
nand U13361 (N_13361,N_13146,N_13238);
nand U13362 (N_13362,N_13159,N_13208);
and U13363 (N_13363,N_13071,N_13099);
xnor U13364 (N_13364,N_13042,N_13061);
or U13365 (N_13365,N_13219,N_13153);
and U13366 (N_13366,N_13217,N_13083);
and U13367 (N_13367,N_13214,N_13095);
or U13368 (N_13368,N_13177,N_13236);
or U13369 (N_13369,N_13069,N_13038);
nor U13370 (N_13370,N_13243,N_13181);
nand U13371 (N_13371,N_13163,N_13144);
nor U13372 (N_13372,N_13166,N_13101);
xor U13373 (N_13373,N_13122,N_13135);
nand U13374 (N_13374,N_13013,N_13059);
nand U13375 (N_13375,N_13216,N_13207);
nor U13376 (N_13376,N_13074,N_13117);
xor U13377 (N_13377,N_13146,N_13093);
xor U13378 (N_13378,N_13191,N_13127);
nand U13379 (N_13379,N_13027,N_13191);
or U13380 (N_13380,N_13095,N_13101);
and U13381 (N_13381,N_13058,N_13149);
or U13382 (N_13382,N_13081,N_13182);
nand U13383 (N_13383,N_13234,N_13090);
nand U13384 (N_13384,N_13166,N_13198);
nand U13385 (N_13385,N_13008,N_13110);
nor U13386 (N_13386,N_13124,N_13001);
nand U13387 (N_13387,N_13011,N_13198);
nor U13388 (N_13388,N_13239,N_13025);
nand U13389 (N_13389,N_13065,N_13173);
and U13390 (N_13390,N_13088,N_13091);
nand U13391 (N_13391,N_13075,N_13077);
and U13392 (N_13392,N_13153,N_13230);
xnor U13393 (N_13393,N_13192,N_13043);
nor U13394 (N_13394,N_13106,N_13097);
or U13395 (N_13395,N_13139,N_13142);
and U13396 (N_13396,N_13192,N_13213);
nor U13397 (N_13397,N_13235,N_13230);
or U13398 (N_13398,N_13086,N_13167);
or U13399 (N_13399,N_13244,N_13142);
nand U13400 (N_13400,N_13215,N_13092);
xor U13401 (N_13401,N_13238,N_13199);
and U13402 (N_13402,N_13108,N_13157);
nor U13403 (N_13403,N_13056,N_13147);
nand U13404 (N_13404,N_13036,N_13129);
xnor U13405 (N_13405,N_13171,N_13071);
nor U13406 (N_13406,N_13176,N_13067);
and U13407 (N_13407,N_13081,N_13050);
nor U13408 (N_13408,N_13023,N_13057);
nand U13409 (N_13409,N_13069,N_13154);
nor U13410 (N_13410,N_13075,N_13194);
nand U13411 (N_13411,N_13103,N_13097);
nand U13412 (N_13412,N_13230,N_13193);
and U13413 (N_13413,N_13226,N_13043);
and U13414 (N_13414,N_13117,N_13030);
or U13415 (N_13415,N_13162,N_13139);
or U13416 (N_13416,N_13194,N_13161);
or U13417 (N_13417,N_13247,N_13104);
nor U13418 (N_13418,N_13077,N_13205);
nand U13419 (N_13419,N_13230,N_13130);
and U13420 (N_13420,N_13074,N_13028);
nor U13421 (N_13421,N_13115,N_13016);
nand U13422 (N_13422,N_13194,N_13040);
and U13423 (N_13423,N_13165,N_13096);
xor U13424 (N_13424,N_13101,N_13224);
nand U13425 (N_13425,N_13027,N_13077);
nor U13426 (N_13426,N_13056,N_13139);
xnor U13427 (N_13427,N_13033,N_13009);
nand U13428 (N_13428,N_13123,N_13145);
nand U13429 (N_13429,N_13048,N_13193);
nand U13430 (N_13430,N_13092,N_13098);
and U13431 (N_13431,N_13023,N_13084);
nor U13432 (N_13432,N_13238,N_13015);
xnor U13433 (N_13433,N_13100,N_13185);
nand U13434 (N_13434,N_13123,N_13205);
nand U13435 (N_13435,N_13243,N_13163);
xor U13436 (N_13436,N_13162,N_13166);
and U13437 (N_13437,N_13110,N_13177);
and U13438 (N_13438,N_13180,N_13196);
and U13439 (N_13439,N_13044,N_13060);
xor U13440 (N_13440,N_13060,N_13229);
and U13441 (N_13441,N_13201,N_13196);
nor U13442 (N_13442,N_13213,N_13111);
or U13443 (N_13443,N_13224,N_13241);
nand U13444 (N_13444,N_13234,N_13147);
or U13445 (N_13445,N_13056,N_13114);
nand U13446 (N_13446,N_13083,N_13175);
xnor U13447 (N_13447,N_13174,N_13147);
nand U13448 (N_13448,N_13170,N_13072);
or U13449 (N_13449,N_13072,N_13204);
xor U13450 (N_13450,N_13201,N_13035);
nand U13451 (N_13451,N_13168,N_13182);
xnor U13452 (N_13452,N_13070,N_13224);
xnor U13453 (N_13453,N_13104,N_13042);
and U13454 (N_13454,N_13119,N_13033);
nand U13455 (N_13455,N_13157,N_13097);
or U13456 (N_13456,N_13208,N_13088);
nand U13457 (N_13457,N_13046,N_13058);
and U13458 (N_13458,N_13107,N_13132);
xor U13459 (N_13459,N_13222,N_13150);
nor U13460 (N_13460,N_13050,N_13203);
xnor U13461 (N_13461,N_13031,N_13142);
and U13462 (N_13462,N_13150,N_13060);
or U13463 (N_13463,N_13032,N_13080);
or U13464 (N_13464,N_13083,N_13202);
nand U13465 (N_13465,N_13208,N_13059);
nand U13466 (N_13466,N_13129,N_13126);
or U13467 (N_13467,N_13216,N_13167);
or U13468 (N_13468,N_13171,N_13187);
xnor U13469 (N_13469,N_13017,N_13025);
and U13470 (N_13470,N_13112,N_13150);
and U13471 (N_13471,N_13013,N_13062);
nand U13472 (N_13472,N_13202,N_13031);
nor U13473 (N_13473,N_13180,N_13003);
xnor U13474 (N_13474,N_13067,N_13222);
nand U13475 (N_13475,N_13119,N_13176);
xnor U13476 (N_13476,N_13223,N_13191);
nand U13477 (N_13477,N_13072,N_13183);
and U13478 (N_13478,N_13141,N_13012);
xnor U13479 (N_13479,N_13030,N_13239);
xnor U13480 (N_13480,N_13129,N_13206);
nor U13481 (N_13481,N_13064,N_13229);
or U13482 (N_13482,N_13070,N_13018);
and U13483 (N_13483,N_13160,N_13032);
and U13484 (N_13484,N_13210,N_13004);
nand U13485 (N_13485,N_13140,N_13204);
xor U13486 (N_13486,N_13212,N_13221);
xor U13487 (N_13487,N_13154,N_13217);
and U13488 (N_13488,N_13128,N_13002);
nand U13489 (N_13489,N_13014,N_13046);
or U13490 (N_13490,N_13176,N_13068);
and U13491 (N_13491,N_13090,N_13166);
xor U13492 (N_13492,N_13044,N_13080);
nand U13493 (N_13493,N_13088,N_13038);
and U13494 (N_13494,N_13035,N_13151);
and U13495 (N_13495,N_13110,N_13023);
nand U13496 (N_13496,N_13186,N_13216);
or U13497 (N_13497,N_13189,N_13247);
xnor U13498 (N_13498,N_13141,N_13130);
nor U13499 (N_13499,N_13003,N_13149);
or U13500 (N_13500,N_13487,N_13410);
nand U13501 (N_13501,N_13302,N_13390);
nor U13502 (N_13502,N_13460,N_13256);
nor U13503 (N_13503,N_13472,N_13342);
nand U13504 (N_13504,N_13369,N_13471);
nor U13505 (N_13505,N_13399,N_13290);
nand U13506 (N_13506,N_13397,N_13400);
xnor U13507 (N_13507,N_13337,N_13269);
or U13508 (N_13508,N_13424,N_13451);
or U13509 (N_13509,N_13359,N_13395);
nand U13510 (N_13510,N_13270,N_13458);
or U13511 (N_13511,N_13352,N_13417);
xnor U13512 (N_13512,N_13478,N_13447);
xor U13513 (N_13513,N_13278,N_13364);
or U13514 (N_13514,N_13455,N_13426);
xnor U13515 (N_13515,N_13363,N_13316);
xnor U13516 (N_13516,N_13354,N_13419);
or U13517 (N_13517,N_13402,N_13493);
nor U13518 (N_13518,N_13298,N_13261);
and U13519 (N_13519,N_13432,N_13409);
or U13520 (N_13520,N_13465,N_13325);
nand U13521 (N_13521,N_13257,N_13279);
xor U13522 (N_13522,N_13449,N_13283);
and U13523 (N_13523,N_13481,N_13489);
nand U13524 (N_13524,N_13355,N_13469);
xor U13525 (N_13525,N_13299,N_13334);
xnor U13526 (N_13526,N_13300,N_13414);
nand U13527 (N_13527,N_13382,N_13450);
nor U13528 (N_13528,N_13368,N_13340);
nand U13529 (N_13529,N_13293,N_13281);
xnor U13530 (N_13530,N_13420,N_13306);
and U13531 (N_13531,N_13254,N_13291);
or U13532 (N_13532,N_13467,N_13305);
and U13533 (N_13533,N_13366,N_13333);
and U13534 (N_13534,N_13464,N_13332);
xor U13535 (N_13535,N_13266,N_13486);
and U13536 (N_13536,N_13386,N_13385);
and U13537 (N_13537,N_13444,N_13327);
xor U13538 (N_13538,N_13427,N_13470);
xor U13539 (N_13539,N_13383,N_13372);
and U13540 (N_13540,N_13362,N_13413);
nor U13541 (N_13541,N_13408,N_13287);
xor U13542 (N_13542,N_13285,N_13379);
nor U13543 (N_13543,N_13341,N_13428);
or U13544 (N_13544,N_13466,N_13259);
nand U13545 (N_13545,N_13274,N_13365);
and U13546 (N_13546,N_13457,N_13477);
xnor U13547 (N_13547,N_13423,N_13326);
or U13548 (N_13548,N_13335,N_13388);
or U13549 (N_13549,N_13317,N_13349);
or U13550 (N_13550,N_13391,N_13485);
or U13551 (N_13551,N_13344,N_13310);
nand U13552 (N_13552,N_13462,N_13314);
or U13553 (N_13553,N_13301,N_13461);
and U13554 (N_13554,N_13289,N_13253);
nand U13555 (N_13555,N_13267,N_13482);
nor U13556 (N_13556,N_13357,N_13348);
or U13557 (N_13557,N_13422,N_13393);
xor U13558 (N_13558,N_13294,N_13430);
or U13559 (N_13559,N_13268,N_13491);
xor U13560 (N_13560,N_13282,N_13381);
xor U13561 (N_13561,N_13396,N_13418);
xnor U13562 (N_13562,N_13387,N_13350);
nand U13563 (N_13563,N_13288,N_13492);
nand U13564 (N_13564,N_13483,N_13251);
xnor U13565 (N_13565,N_13436,N_13304);
nor U13566 (N_13566,N_13415,N_13263);
and U13567 (N_13567,N_13404,N_13272);
or U13568 (N_13568,N_13262,N_13318);
or U13569 (N_13569,N_13429,N_13371);
nand U13570 (N_13570,N_13438,N_13403);
and U13571 (N_13571,N_13330,N_13474);
nor U13572 (N_13572,N_13360,N_13373);
xnor U13573 (N_13573,N_13412,N_13280);
nand U13574 (N_13574,N_13277,N_13361);
nand U13575 (N_13575,N_13498,N_13490);
and U13576 (N_13576,N_13452,N_13319);
or U13577 (N_13577,N_13339,N_13445);
nor U13578 (N_13578,N_13434,N_13459);
xnor U13579 (N_13579,N_13320,N_13435);
nand U13580 (N_13580,N_13497,N_13384);
xnor U13581 (N_13581,N_13421,N_13475);
nor U13582 (N_13582,N_13303,N_13440);
and U13583 (N_13583,N_13358,N_13297);
or U13584 (N_13584,N_13416,N_13377);
and U13585 (N_13585,N_13343,N_13367);
nor U13586 (N_13586,N_13463,N_13442);
and U13587 (N_13587,N_13380,N_13324);
xnor U13588 (N_13588,N_13456,N_13411);
xnor U13589 (N_13589,N_13284,N_13338);
and U13590 (N_13590,N_13315,N_13295);
and U13591 (N_13591,N_13292,N_13441);
nor U13592 (N_13592,N_13378,N_13311);
nand U13593 (N_13593,N_13286,N_13323);
xor U13594 (N_13594,N_13374,N_13394);
nor U13595 (N_13595,N_13405,N_13271);
nand U13596 (N_13596,N_13331,N_13389);
and U13597 (N_13597,N_13479,N_13264);
nor U13598 (N_13598,N_13370,N_13488);
or U13599 (N_13599,N_13431,N_13407);
nor U13600 (N_13600,N_13401,N_13496);
xnor U13601 (N_13601,N_13476,N_13322);
nand U13602 (N_13602,N_13453,N_13439);
nor U13603 (N_13603,N_13329,N_13313);
nor U13604 (N_13604,N_13468,N_13437);
and U13605 (N_13605,N_13308,N_13260);
and U13606 (N_13606,N_13406,N_13265);
xnor U13607 (N_13607,N_13376,N_13321);
nand U13608 (N_13608,N_13375,N_13307);
nor U13609 (N_13609,N_13347,N_13328);
or U13610 (N_13610,N_13309,N_13255);
xnor U13611 (N_13611,N_13345,N_13480);
nand U13612 (N_13612,N_13346,N_13484);
nor U13613 (N_13613,N_13425,N_13433);
nor U13614 (N_13614,N_13312,N_13454);
and U13615 (N_13615,N_13336,N_13273);
nor U13616 (N_13616,N_13353,N_13392);
xor U13617 (N_13617,N_13258,N_13473);
nor U13618 (N_13618,N_13275,N_13446);
and U13619 (N_13619,N_13252,N_13448);
and U13620 (N_13620,N_13296,N_13276);
or U13621 (N_13621,N_13351,N_13495);
xor U13622 (N_13622,N_13356,N_13494);
nand U13623 (N_13623,N_13398,N_13499);
nand U13624 (N_13624,N_13443,N_13250);
or U13625 (N_13625,N_13466,N_13329);
xor U13626 (N_13626,N_13479,N_13306);
nand U13627 (N_13627,N_13491,N_13398);
nand U13628 (N_13628,N_13466,N_13409);
nor U13629 (N_13629,N_13483,N_13454);
xnor U13630 (N_13630,N_13481,N_13300);
xnor U13631 (N_13631,N_13255,N_13482);
and U13632 (N_13632,N_13387,N_13252);
or U13633 (N_13633,N_13382,N_13470);
or U13634 (N_13634,N_13306,N_13330);
or U13635 (N_13635,N_13449,N_13291);
or U13636 (N_13636,N_13311,N_13307);
xor U13637 (N_13637,N_13385,N_13282);
or U13638 (N_13638,N_13316,N_13306);
nor U13639 (N_13639,N_13269,N_13263);
nand U13640 (N_13640,N_13428,N_13402);
nor U13641 (N_13641,N_13306,N_13317);
nor U13642 (N_13642,N_13258,N_13470);
nor U13643 (N_13643,N_13382,N_13468);
and U13644 (N_13644,N_13400,N_13496);
xor U13645 (N_13645,N_13388,N_13337);
nand U13646 (N_13646,N_13285,N_13310);
xor U13647 (N_13647,N_13434,N_13469);
nor U13648 (N_13648,N_13287,N_13311);
xnor U13649 (N_13649,N_13408,N_13316);
nand U13650 (N_13650,N_13449,N_13259);
nand U13651 (N_13651,N_13255,N_13432);
nand U13652 (N_13652,N_13359,N_13421);
and U13653 (N_13653,N_13369,N_13290);
nor U13654 (N_13654,N_13303,N_13302);
or U13655 (N_13655,N_13352,N_13373);
and U13656 (N_13656,N_13446,N_13394);
or U13657 (N_13657,N_13371,N_13377);
and U13658 (N_13658,N_13255,N_13268);
nand U13659 (N_13659,N_13319,N_13253);
nand U13660 (N_13660,N_13366,N_13295);
xnor U13661 (N_13661,N_13395,N_13282);
nor U13662 (N_13662,N_13474,N_13494);
or U13663 (N_13663,N_13489,N_13439);
and U13664 (N_13664,N_13439,N_13446);
nand U13665 (N_13665,N_13324,N_13386);
nand U13666 (N_13666,N_13367,N_13299);
or U13667 (N_13667,N_13470,N_13413);
and U13668 (N_13668,N_13393,N_13312);
nor U13669 (N_13669,N_13410,N_13463);
nor U13670 (N_13670,N_13298,N_13482);
nor U13671 (N_13671,N_13341,N_13337);
nor U13672 (N_13672,N_13372,N_13306);
xnor U13673 (N_13673,N_13417,N_13330);
and U13674 (N_13674,N_13461,N_13257);
or U13675 (N_13675,N_13387,N_13311);
or U13676 (N_13676,N_13275,N_13497);
or U13677 (N_13677,N_13362,N_13359);
nand U13678 (N_13678,N_13311,N_13259);
xor U13679 (N_13679,N_13278,N_13341);
nand U13680 (N_13680,N_13386,N_13478);
nand U13681 (N_13681,N_13388,N_13406);
nor U13682 (N_13682,N_13325,N_13318);
and U13683 (N_13683,N_13300,N_13304);
nand U13684 (N_13684,N_13428,N_13292);
xor U13685 (N_13685,N_13332,N_13290);
nand U13686 (N_13686,N_13309,N_13486);
and U13687 (N_13687,N_13331,N_13271);
nand U13688 (N_13688,N_13385,N_13436);
and U13689 (N_13689,N_13428,N_13493);
nor U13690 (N_13690,N_13425,N_13281);
nor U13691 (N_13691,N_13453,N_13271);
or U13692 (N_13692,N_13351,N_13325);
nor U13693 (N_13693,N_13267,N_13299);
and U13694 (N_13694,N_13289,N_13393);
or U13695 (N_13695,N_13459,N_13338);
and U13696 (N_13696,N_13287,N_13318);
xor U13697 (N_13697,N_13253,N_13330);
nand U13698 (N_13698,N_13487,N_13473);
and U13699 (N_13699,N_13304,N_13493);
or U13700 (N_13700,N_13486,N_13462);
xor U13701 (N_13701,N_13264,N_13254);
nor U13702 (N_13702,N_13305,N_13252);
nor U13703 (N_13703,N_13442,N_13424);
and U13704 (N_13704,N_13286,N_13390);
nor U13705 (N_13705,N_13331,N_13320);
nor U13706 (N_13706,N_13427,N_13376);
or U13707 (N_13707,N_13474,N_13461);
and U13708 (N_13708,N_13293,N_13363);
nand U13709 (N_13709,N_13381,N_13251);
nor U13710 (N_13710,N_13341,N_13283);
nor U13711 (N_13711,N_13356,N_13384);
and U13712 (N_13712,N_13463,N_13280);
nor U13713 (N_13713,N_13364,N_13372);
and U13714 (N_13714,N_13310,N_13429);
and U13715 (N_13715,N_13277,N_13371);
xnor U13716 (N_13716,N_13315,N_13480);
nor U13717 (N_13717,N_13433,N_13399);
and U13718 (N_13718,N_13289,N_13489);
nor U13719 (N_13719,N_13394,N_13326);
nor U13720 (N_13720,N_13321,N_13345);
nand U13721 (N_13721,N_13375,N_13391);
nand U13722 (N_13722,N_13383,N_13311);
or U13723 (N_13723,N_13296,N_13317);
nand U13724 (N_13724,N_13494,N_13464);
nand U13725 (N_13725,N_13403,N_13395);
nor U13726 (N_13726,N_13263,N_13417);
nand U13727 (N_13727,N_13316,N_13432);
nand U13728 (N_13728,N_13490,N_13473);
nor U13729 (N_13729,N_13485,N_13264);
or U13730 (N_13730,N_13420,N_13483);
nand U13731 (N_13731,N_13481,N_13437);
nor U13732 (N_13732,N_13363,N_13420);
and U13733 (N_13733,N_13403,N_13277);
and U13734 (N_13734,N_13279,N_13255);
nor U13735 (N_13735,N_13272,N_13405);
xnor U13736 (N_13736,N_13325,N_13352);
or U13737 (N_13737,N_13346,N_13356);
nor U13738 (N_13738,N_13261,N_13308);
nor U13739 (N_13739,N_13399,N_13487);
or U13740 (N_13740,N_13299,N_13250);
nand U13741 (N_13741,N_13360,N_13480);
or U13742 (N_13742,N_13474,N_13393);
nor U13743 (N_13743,N_13428,N_13266);
or U13744 (N_13744,N_13410,N_13368);
or U13745 (N_13745,N_13370,N_13432);
and U13746 (N_13746,N_13433,N_13328);
nor U13747 (N_13747,N_13410,N_13396);
xnor U13748 (N_13748,N_13451,N_13461);
nor U13749 (N_13749,N_13318,N_13491);
nor U13750 (N_13750,N_13748,N_13566);
xor U13751 (N_13751,N_13568,N_13604);
and U13752 (N_13752,N_13690,N_13679);
or U13753 (N_13753,N_13639,N_13734);
or U13754 (N_13754,N_13707,N_13630);
and U13755 (N_13755,N_13557,N_13590);
xnor U13756 (N_13756,N_13747,N_13550);
xor U13757 (N_13757,N_13562,N_13695);
nor U13758 (N_13758,N_13537,N_13737);
xor U13759 (N_13759,N_13588,N_13688);
and U13760 (N_13760,N_13549,N_13569);
and U13761 (N_13761,N_13720,N_13623);
xor U13762 (N_13762,N_13703,N_13656);
or U13763 (N_13763,N_13522,N_13647);
xor U13764 (N_13764,N_13591,N_13560);
or U13765 (N_13765,N_13666,N_13663);
xor U13766 (N_13766,N_13519,N_13581);
xnor U13767 (N_13767,N_13685,N_13683);
and U13768 (N_13768,N_13572,N_13744);
nor U13769 (N_13769,N_13536,N_13555);
nand U13770 (N_13770,N_13578,N_13520);
xnor U13771 (N_13771,N_13680,N_13514);
and U13772 (N_13772,N_13634,N_13657);
and U13773 (N_13773,N_13582,N_13697);
nand U13774 (N_13774,N_13548,N_13619);
nand U13775 (N_13775,N_13704,N_13711);
or U13776 (N_13776,N_13606,N_13573);
nand U13777 (N_13777,N_13509,N_13551);
or U13778 (N_13778,N_13714,N_13521);
nand U13779 (N_13779,N_13628,N_13529);
or U13780 (N_13780,N_13513,N_13653);
nand U13781 (N_13781,N_13501,N_13559);
nor U13782 (N_13782,N_13601,N_13561);
and U13783 (N_13783,N_13611,N_13727);
and U13784 (N_13784,N_13625,N_13741);
xor U13785 (N_13785,N_13694,N_13698);
xnor U13786 (N_13786,N_13651,N_13618);
xnor U13787 (N_13787,N_13570,N_13615);
nor U13788 (N_13788,N_13696,N_13652);
xor U13789 (N_13789,N_13546,N_13621);
xnor U13790 (N_13790,N_13543,N_13511);
or U13791 (N_13791,N_13641,N_13700);
nor U13792 (N_13792,N_13508,N_13580);
nand U13793 (N_13793,N_13595,N_13556);
nand U13794 (N_13794,N_13575,N_13567);
or U13795 (N_13795,N_13667,N_13669);
nor U13796 (N_13796,N_13563,N_13665);
xnor U13797 (N_13797,N_13583,N_13502);
nor U13798 (N_13798,N_13503,N_13539);
nor U13799 (N_13799,N_13574,N_13723);
nand U13800 (N_13800,N_13544,N_13662);
or U13801 (N_13801,N_13609,N_13594);
and U13802 (N_13802,N_13620,N_13589);
or U13803 (N_13803,N_13646,N_13693);
nor U13804 (N_13804,N_13612,N_13719);
nor U13805 (N_13805,N_13532,N_13614);
xnor U13806 (N_13806,N_13541,N_13616);
or U13807 (N_13807,N_13728,N_13661);
nor U13808 (N_13808,N_13730,N_13565);
or U13809 (N_13809,N_13731,N_13689);
nor U13810 (N_13810,N_13733,N_13554);
or U13811 (N_13811,N_13523,N_13642);
nand U13812 (N_13812,N_13505,N_13673);
nor U13813 (N_13813,N_13596,N_13712);
and U13814 (N_13814,N_13736,N_13650);
and U13815 (N_13815,N_13743,N_13678);
or U13816 (N_13816,N_13558,N_13664);
or U13817 (N_13817,N_13713,N_13699);
xor U13818 (N_13818,N_13674,N_13709);
xnor U13819 (N_13819,N_13708,N_13597);
xnor U13820 (N_13820,N_13524,N_13626);
nor U13821 (N_13821,N_13553,N_13638);
nor U13822 (N_13822,N_13517,N_13655);
or U13823 (N_13823,N_13538,N_13610);
and U13824 (N_13824,N_13593,N_13605);
nor U13825 (N_13825,N_13691,N_13585);
nand U13826 (N_13826,N_13617,N_13608);
or U13827 (N_13827,N_13645,N_13671);
nand U13828 (N_13828,N_13518,N_13643);
nor U13829 (N_13829,N_13571,N_13746);
xor U13830 (N_13830,N_13721,N_13510);
nand U13831 (N_13831,N_13710,N_13516);
and U13832 (N_13832,N_13705,N_13716);
or U13833 (N_13833,N_13528,N_13670);
xnor U13834 (N_13834,N_13542,N_13624);
nand U13835 (N_13835,N_13715,N_13701);
nor U13836 (N_13836,N_13668,N_13598);
and U13837 (N_13837,N_13592,N_13512);
xor U13838 (N_13838,N_13735,N_13675);
xor U13839 (N_13839,N_13672,N_13692);
and U13840 (N_13840,N_13603,N_13681);
xor U13841 (N_13841,N_13729,N_13545);
xor U13842 (N_13842,N_13660,N_13649);
xnor U13843 (N_13843,N_13749,N_13726);
and U13844 (N_13844,N_13530,N_13635);
or U13845 (N_13845,N_13507,N_13525);
nand U13846 (N_13846,N_13640,N_13722);
nand U13847 (N_13847,N_13535,N_13632);
or U13848 (N_13848,N_13587,N_13740);
and U13849 (N_13849,N_13506,N_13725);
xor U13850 (N_13850,N_13627,N_13677);
or U13851 (N_13851,N_13552,N_13648);
or U13852 (N_13852,N_13724,N_13659);
and U13853 (N_13853,N_13629,N_13658);
and U13854 (N_13854,N_13607,N_13584);
nand U13855 (N_13855,N_13577,N_13739);
nand U13856 (N_13856,N_13742,N_13676);
and U13857 (N_13857,N_13576,N_13684);
xor U13858 (N_13858,N_13526,N_13636);
nor U13859 (N_13859,N_13531,N_13633);
nor U13860 (N_13860,N_13547,N_13602);
and U13861 (N_13861,N_13599,N_13533);
and U13862 (N_13862,N_13644,N_13682);
or U13863 (N_13863,N_13732,N_13500);
or U13864 (N_13864,N_13718,N_13613);
nand U13865 (N_13865,N_13515,N_13586);
xor U13866 (N_13866,N_13631,N_13579);
or U13867 (N_13867,N_13540,N_13738);
or U13868 (N_13868,N_13702,N_13706);
nor U13869 (N_13869,N_13534,N_13527);
and U13870 (N_13870,N_13687,N_13654);
xnor U13871 (N_13871,N_13600,N_13686);
nand U13872 (N_13872,N_13637,N_13504);
nand U13873 (N_13873,N_13564,N_13622);
and U13874 (N_13874,N_13745,N_13717);
or U13875 (N_13875,N_13663,N_13682);
or U13876 (N_13876,N_13541,N_13677);
nor U13877 (N_13877,N_13591,N_13501);
or U13878 (N_13878,N_13632,N_13685);
nand U13879 (N_13879,N_13626,N_13676);
and U13880 (N_13880,N_13687,N_13686);
or U13881 (N_13881,N_13538,N_13639);
nor U13882 (N_13882,N_13693,N_13503);
and U13883 (N_13883,N_13716,N_13616);
nand U13884 (N_13884,N_13574,N_13686);
and U13885 (N_13885,N_13748,N_13519);
xor U13886 (N_13886,N_13538,N_13629);
nor U13887 (N_13887,N_13527,N_13617);
nor U13888 (N_13888,N_13545,N_13650);
nand U13889 (N_13889,N_13690,N_13547);
nor U13890 (N_13890,N_13531,N_13606);
and U13891 (N_13891,N_13705,N_13727);
and U13892 (N_13892,N_13505,N_13557);
nand U13893 (N_13893,N_13612,N_13504);
and U13894 (N_13894,N_13733,N_13671);
xor U13895 (N_13895,N_13599,N_13633);
or U13896 (N_13896,N_13597,N_13575);
xnor U13897 (N_13897,N_13517,N_13642);
nor U13898 (N_13898,N_13596,N_13645);
and U13899 (N_13899,N_13613,N_13713);
nor U13900 (N_13900,N_13508,N_13579);
nor U13901 (N_13901,N_13598,N_13736);
nand U13902 (N_13902,N_13714,N_13517);
nor U13903 (N_13903,N_13613,N_13580);
and U13904 (N_13904,N_13644,N_13521);
nand U13905 (N_13905,N_13740,N_13555);
xnor U13906 (N_13906,N_13701,N_13519);
nor U13907 (N_13907,N_13592,N_13726);
nor U13908 (N_13908,N_13583,N_13573);
and U13909 (N_13909,N_13554,N_13547);
nor U13910 (N_13910,N_13745,N_13638);
nand U13911 (N_13911,N_13703,N_13662);
nor U13912 (N_13912,N_13600,N_13646);
xnor U13913 (N_13913,N_13704,N_13567);
nand U13914 (N_13914,N_13603,N_13575);
xor U13915 (N_13915,N_13713,N_13619);
xnor U13916 (N_13916,N_13600,N_13572);
nand U13917 (N_13917,N_13657,N_13670);
xnor U13918 (N_13918,N_13735,N_13656);
nor U13919 (N_13919,N_13629,N_13730);
xor U13920 (N_13920,N_13621,N_13679);
or U13921 (N_13921,N_13564,N_13637);
and U13922 (N_13922,N_13676,N_13642);
or U13923 (N_13923,N_13670,N_13597);
nor U13924 (N_13924,N_13582,N_13679);
nor U13925 (N_13925,N_13641,N_13628);
nand U13926 (N_13926,N_13640,N_13516);
or U13927 (N_13927,N_13602,N_13601);
and U13928 (N_13928,N_13553,N_13578);
nand U13929 (N_13929,N_13553,N_13635);
xor U13930 (N_13930,N_13738,N_13707);
and U13931 (N_13931,N_13609,N_13607);
nor U13932 (N_13932,N_13547,N_13541);
or U13933 (N_13933,N_13580,N_13661);
or U13934 (N_13934,N_13714,N_13590);
xor U13935 (N_13935,N_13641,N_13745);
xnor U13936 (N_13936,N_13707,N_13523);
nand U13937 (N_13937,N_13731,N_13718);
xor U13938 (N_13938,N_13748,N_13662);
nor U13939 (N_13939,N_13548,N_13701);
nand U13940 (N_13940,N_13630,N_13721);
xnor U13941 (N_13941,N_13601,N_13678);
or U13942 (N_13942,N_13685,N_13561);
and U13943 (N_13943,N_13559,N_13705);
nor U13944 (N_13944,N_13630,N_13526);
or U13945 (N_13945,N_13573,N_13535);
xnor U13946 (N_13946,N_13731,N_13593);
nand U13947 (N_13947,N_13641,N_13604);
or U13948 (N_13948,N_13553,N_13735);
or U13949 (N_13949,N_13687,N_13595);
xor U13950 (N_13950,N_13681,N_13655);
nor U13951 (N_13951,N_13691,N_13570);
and U13952 (N_13952,N_13540,N_13619);
nand U13953 (N_13953,N_13613,N_13570);
nor U13954 (N_13954,N_13701,N_13588);
and U13955 (N_13955,N_13604,N_13714);
nor U13956 (N_13956,N_13568,N_13741);
nand U13957 (N_13957,N_13702,N_13583);
and U13958 (N_13958,N_13626,N_13573);
and U13959 (N_13959,N_13509,N_13552);
and U13960 (N_13960,N_13548,N_13633);
nor U13961 (N_13961,N_13738,N_13734);
nor U13962 (N_13962,N_13563,N_13607);
xor U13963 (N_13963,N_13591,N_13527);
or U13964 (N_13964,N_13730,N_13737);
and U13965 (N_13965,N_13737,N_13686);
or U13966 (N_13966,N_13585,N_13670);
nand U13967 (N_13967,N_13667,N_13623);
nor U13968 (N_13968,N_13671,N_13734);
and U13969 (N_13969,N_13671,N_13712);
and U13970 (N_13970,N_13562,N_13676);
nand U13971 (N_13971,N_13589,N_13551);
nor U13972 (N_13972,N_13638,N_13535);
or U13973 (N_13973,N_13697,N_13683);
and U13974 (N_13974,N_13560,N_13727);
and U13975 (N_13975,N_13691,N_13643);
xor U13976 (N_13976,N_13652,N_13580);
nor U13977 (N_13977,N_13605,N_13679);
nand U13978 (N_13978,N_13576,N_13534);
and U13979 (N_13979,N_13548,N_13663);
and U13980 (N_13980,N_13549,N_13701);
nand U13981 (N_13981,N_13696,N_13599);
and U13982 (N_13982,N_13579,N_13593);
nand U13983 (N_13983,N_13500,N_13561);
xor U13984 (N_13984,N_13514,N_13506);
and U13985 (N_13985,N_13652,N_13574);
xor U13986 (N_13986,N_13524,N_13587);
nand U13987 (N_13987,N_13729,N_13739);
or U13988 (N_13988,N_13656,N_13741);
and U13989 (N_13989,N_13664,N_13603);
xnor U13990 (N_13990,N_13560,N_13559);
nand U13991 (N_13991,N_13662,N_13597);
nor U13992 (N_13992,N_13717,N_13540);
xor U13993 (N_13993,N_13657,N_13648);
or U13994 (N_13994,N_13699,N_13574);
xnor U13995 (N_13995,N_13580,N_13700);
and U13996 (N_13996,N_13589,N_13680);
or U13997 (N_13997,N_13689,N_13553);
nand U13998 (N_13998,N_13645,N_13699);
nor U13999 (N_13999,N_13507,N_13726);
or U14000 (N_14000,N_13857,N_13993);
nand U14001 (N_14001,N_13998,N_13860);
xor U14002 (N_14002,N_13936,N_13995);
or U14003 (N_14003,N_13957,N_13808);
and U14004 (N_14004,N_13846,N_13985);
xor U14005 (N_14005,N_13844,N_13773);
nor U14006 (N_14006,N_13818,N_13793);
nand U14007 (N_14007,N_13812,N_13832);
nand U14008 (N_14008,N_13990,N_13837);
xor U14009 (N_14009,N_13884,N_13786);
nor U14010 (N_14010,N_13902,N_13790);
and U14011 (N_14011,N_13777,N_13839);
xnor U14012 (N_14012,N_13804,N_13999);
nor U14013 (N_14013,N_13827,N_13881);
and U14014 (N_14014,N_13983,N_13918);
nand U14015 (N_14015,N_13771,N_13965);
and U14016 (N_14016,N_13824,N_13893);
and U14017 (N_14017,N_13778,N_13756);
nor U14018 (N_14018,N_13866,N_13976);
xor U14019 (N_14019,N_13895,N_13770);
nor U14020 (N_14020,N_13916,N_13810);
nand U14021 (N_14021,N_13903,N_13766);
nand U14022 (N_14022,N_13755,N_13809);
or U14023 (N_14023,N_13831,N_13800);
xor U14024 (N_14024,N_13845,N_13926);
or U14025 (N_14025,N_13940,N_13872);
xnor U14026 (N_14026,N_13888,N_13750);
or U14027 (N_14027,N_13795,N_13987);
nor U14028 (N_14028,N_13937,N_13996);
nand U14029 (N_14029,N_13819,N_13973);
or U14030 (N_14030,N_13885,N_13972);
and U14031 (N_14031,N_13967,N_13910);
nor U14032 (N_14032,N_13823,N_13991);
or U14033 (N_14033,N_13864,N_13782);
nand U14034 (N_14034,N_13939,N_13779);
nand U14035 (N_14035,N_13858,N_13801);
nand U14036 (N_14036,N_13751,N_13761);
nor U14037 (N_14037,N_13970,N_13963);
or U14038 (N_14038,N_13891,N_13988);
nor U14039 (N_14039,N_13989,N_13925);
and U14040 (N_14040,N_13835,N_13856);
and U14041 (N_14041,N_13933,N_13941);
nor U14042 (N_14042,N_13960,N_13799);
and U14043 (N_14043,N_13909,N_13964);
and U14044 (N_14044,N_13994,N_13838);
and U14045 (N_14045,N_13877,N_13861);
and U14046 (N_14046,N_13843,N_13982);
nand U14047 (N_14047,N_13915,N_13968);
xnor U14048 (N_14048,N_13871,N_13934);
or U14049 (N_14049,N_13978,N_13797);
or U14050 (N_14050,N_13875,N_13919);
xor U14051 (N_14051,N_13772,N_13953);
nor U14052 (N_14052,N_13896,N_13904);
xnor U14053 (N_14053,N_13956,N_13883);
xor U14054 (N_14054,N_13950,N_13813);
and U14055 (N_14055,N_13851,N_13792);
and U14056 (N_14056,N_13788,N_13874);
and U14057 (N_14057,N_13791,N_13959);
or U14058 (N_14058,N_13892,N_13894);
xor U14059 (N_14059,N_13986,N_13769);
nor U14060 (N_14060,N_13927,N_13913);
and U14061 (N_14061,N_13762,N_13898);
and U14062 (N_14062,N_13820,N_13815);
and U14063 (N_14063,N_13997,N_13863);
xnor U14064 (N_14064,N_13981,N_13974);
and U14065 (N_14065,N_13803,N_13979);
or U14066 (N_14066,N_13805,N_13833);
nand U14067 (N_14067,N_13911,N_13840);
and U14068 (N_14068,N_13900,N_13811);
and U14069 (N_14069,N_13971,N_13943);
or U14070 (N_14070,N_13876,N_13764);
nor U14071 (N_14071,N_13935,N_13930);
and U14072 (N_14072,N_13841,N_13855);
nor U14073 (N_14073,N_13754,N_13865);
nand U14074 (N_14074,N_13859,N_13775);
nand U14075 (N_14075,N_13869,N_13908);
or U14076 (N_14076,N_13853,N_13905);
or U14077 (N_14077,N_13873,N_13944);
nor U14078 (N_14078,N_13868,N_13946);
nor U14079 (N_14079,N_13802,N_13980);
xor U14080 (N_14080,N_13961,N_13862);
nor U14081 (N_14081,N_13958,N_13969);
and U14082 (N_14082,N_13879,N_13922);
or U14083 (N_14083,N_13951,N_13829);
nor U14084 (N_14084,N_13848,N_13757);
nand U14085 (N_14085,N_13882,N_13784);
xor U14086 (N_14086,N_13901,N_13752);
xor U14087 (N_14087,N_13984,N_13758);
xor U14088 (N_14088,N_13947,N_13952);
and U14089 (N_14089,N_13899,N_13854);
nand U14090 (N_14090,N_13796,N_13938);
and U14091 (N_14091,N_13850,N_13966);
and U14092 (N_14092,N_13849,N_13912);
or U14093 (N_14093,N_13867,N_13920);
and U14094 (N_14094,N_13924,N_13928);
nor U14095 (N_14095,N_13794,N_13753);
nor U14096 (N_14096,N_13760,N_13774);
and U14097 (N_14097,N_13817,N_13945);
nand U14098 (N_14098,N_13962,N_13787);
or U14099 (N_14099,N_13917,N_13826);
xor U14100 (N_14100,N_13781,N_13886);
xnor U14101 (N_14101,N_13768,N_13798);
or U14102 (N_14102,N_13834,N_13906);
and U14103 (N_14103,N_13763,N_13931);
nand U14104 (N_14104,N_13932,N_13907);
and U14105 (N_14105,N_13816,N_13890);
xor U14106 (N_14106,N_13765,N_13948);
xor U14107 (N_14107,N_13767,N_13975);
nand U14108 (N_14108,N_13825,N_13949);
and U14109 (N_14109,N_13785,N_13992);
and U14110 (N_14110,N_13897,N_13852);
and U14111 (N_14111,N_13806,N_13814);
nor U14112 (N_14112,N_13821,N_13914);
and U14113 (N_14113,N_13783,N_13887);
and U14114 (N_14114,N_13942,N_13955);
nand U14115 (N_14115,N_13889,N_13954);
nand U14116 (N_14116,N_13870,N_13842);
and U14117 (N_14117,N_13847,N_13878);
or U14118 (N_14118,N_13921,N_13923);
xnor U14119 (N_14119,N_13828,N_13780);
xor U14120 (N_14120,N_13776,N_13789);
or U14121 (N_14121,N_13929,N_13830);
xor U14122 (N_14122,N_13836,N_13977);
and U14123 (N_14123,N_13822,N_13759);
and U14124 (N_14124,N_13807,N_13880);
nand U14125 (N_14125,N_13864,N_13955);
xor U14126 (N_14126,N_13808,N_13857);
nor U14127 (N_14127,N_13948,N_13929);
nor U14128 (N_14128,N_13863,N_13759);
or U14129 (N_14129,N_13782,N_13863);
and U14130 (N_14130,N_13870,N_13997);
xnor U14131 (N_14131,N_13818,N_13820);
and U14132 (N_14132,N_13913,N_13760);
nor U14133 (N_14133,N_13905,N_13983);
and U14134 (N_14134,N_13796,N_13795);
xor U14135 (N_14135,N_13822,N_13977);
nand U14136 (N_14136,N_13755,N_13981);
nand U14137 (N_14137,N_13767,N_13917);
nand U14138 (N_14138,N_13908,N_13777);
or U14139 (N_14139,N_13807,N_13769);
nor U14140 (N_14140,N_13885,N_13845);
nand U14141 (N_14141,N_13813,N_13861);
and U14142 (N_14142,N_13895,N_13846);
nand U14143 (N_14143,N_13825,N_13876);
or U14144 (N_14144,N_13900,N_13893);
nor U14145 (N_14145,N_13848,N_13985);
nand U14146 (N_14146,N_13892,N_13817);
nand U14147 (N_14147,N_13959,N_13796);
nand U14148 (N_14148,N_13921,N_13955);
nor U14149 (N_14149,N_13836,N_13960);
nor U14150 (N_14150,N_13867,N_13930);
xnor U14151 (N_14151,N_13810,N_13851);
or U14152 (N_14152,N_13917,N_13925);
nor U14153 (N_14153,N_13836,N_13832);
nor U14154 (N_14154,N_13905,N_13942);
xnor U14155 (N_14155,N_13786,N_13765);
nor U14156 (N_14156,N_13779,N_13821);
nor U14157 (N_14157,N_13940,N_13910);
and U14158 (N_14158,N_13969,N_13949);
xnor U14159 (N_14159,N_13988,N_13858);
nor U14160 (N_14160,N_13883,N_13868);
nor U14161 (N_14161,N_13961,N_13782);
nor U14162 (N_14162,N_13962,N_13968);
nand U14163 (N_14163,N_13853,N_13823);
xor U14164 (N_14164,N_13811,N_13860);
nand U14165 (N_14165,N_13885,N_13788);
nand U14166 (N_14166,N_13878,N_13953);
and U14167 (N_14167,N_13943,N_13812);
nor U14168 (N_14168,N_13925,N_13843);
or U14169 (N_14169,N_13903,N_13758);
nand U14170 (N_14170,N_13851,N_13991);
and U14171 (N_14171,N_13895,N_13806);
and U14172 (N_14172,N_13916,N_13906);
or U14173 (N_14173,N_13993,N_13932);
and U14174 (N_14174,N_13907,N_13803);
or U14175 (N_14175,N_13928,N_13915);
nor U14176 (N_14176,N_13845,N_13957);
xor U14177 (N_14177,N_13942,N_13819);
nand U14178 (N_14178,N_13786,N_13950);
and U14179 (N_14179,N_13952,N_13863);
xor U14180 (N_14180,N_13788,N_13987);
or U14181 (N_14181,N_13826,N_13875);
and U14182 (N_14182,N_13754,N_13822);
xor U14183 (N_14183,N_13917,N_13817);
xor U14184 (N_14184,N_13798,N_13859);
or U14185 (N_14185,N_13997,N_13884);
nor U14186 (N_14186,N_13790,N_13802);
nand U14187 (N_14187,N_13838,N_13893);
xor U14188 (N_14188,N_13952,N_13813);
xor U14189 (N_14189,N_13885,N_13851);
and U14190 (N_14190,N_13766,N_13894);
xor U14191 (N_14191,N_13992,N_13990);
and U14192 (N_14192,N_13760,N_13825);
or U14193 (N_14193,N_13987,N_13926);
xor U14194 (N_14194,N_13976,N_13846);
nor U14195 (N_14195,N_13947,N_13967);
or U14196 (N_14196,N_13985,N_13822);
nor U14197 (N_14197,N_13776,N_13781);
nand U14198 (N_14198,N_13960,N_13776);
xnor U14199 (N_14199,N_13786,N_13879);
nand U14200 (N_14200,N_13866,N_13993);
and U14201 (N_14201,N_13827,N_13770);
or U14202 (N_14202,N_13974,N_13920);
nand U14203 (N_14203,N_13761,N_13941);
or U14204 (N_14204,N_13789,N_13860);
nor U14205 (N_14205,N_13957,N_13771);
and U14206 (N_14206,N_13812,N_13975);
or U14207 (N_14207,N_13973,N_13764);
nor U14208 (N_14208,N_13945,N_13832);
xnor U14209 (N_14209,N_13773,N_13919);
xor U14210 (N_14210,N_13979,N_13843);
or U14211 (N_14211,N_13892,N_13794);
nor U14212 (N_14212,N_13936,N_13780);
and U14213 (N_14213,N_13824,N_13892);
nand U14214 (N_14214,N_13960,N_13811);
nor U14215 (N_14215,N_13785,N_13991);
xnor U14216 (N_14216,N_13820,N_13908);
or U14217 (N_14217,N_13769,N_13844);
xnor U14218 (N_14218,N_13828,N_13822);
nor U14219 (N_14219,N_13817,N_13932);
xor U14220 (N_14220,N_13854,N_13790);
xor U14221 (N_14221,N_13972,N_13903);
and U14222 (N_14222,N_13796,N_13961);
or U14223 (N_14223,N_13953,N_13795);
nand U14224 (N_14224,N_13779,N_13893);
xor U14225 (N_14225,N_13859,N_13846);
nor U14226 (N_14226,N_13914,N_13777);
nor U14227 (N_14227,N_13936,N_13896);
or U14228 (N_14228,N_13943,N_13893);
nor U14229 (N_14229,N_13949,N_13833);
nor U14230 (N_14230,N_13989,N_13876);
nor U14231 (N_14231,N_13789,N_13888);
nand U14232 (N_14232,N_13971,N_13803);
nor U14233 (N_14233,N_13831,N_13933);
nand U14234 (N_14234,N_13989,N_13768);
and U14235 (N_14235,N_13796,N_13800);
xor U14236 (N_14236,N_13872,N_13820);
and U14237 (N_14237,N_13930,N_13817);
nand U14238 (N_14238,N_13922,N_13925);
nor U14239 (N_14239,N_13904,N_13946);
nand U14240 (N_14240,N_13915,N_13797);
or U14241 (N_14241,N_13912,N_13957);
and U14242 (N_14242,N_13858,N_13900);
and U14243 (N_14243,N_13974,N_13857);
nor U14244 (N_14244,N_13988,N_13959);
and U14245 (N_14245,N_13762,N_13928);
or U14246 (N_14246,N_13803,N_13781);
or U14247 (N_14247,N_13827,N_13909);
or U14248 (N_14248,N_13862,N_13813);
xnor U14249 (N_14249,N_13908,N_13990);
nand U14250 (N_14250,N_14209,N_14180);
and U14251 (N_14251,N_14065,N_14092);
nor U14252 (N_14252,N_14116,N_14201);
or U14253 (N_14253,N_14082,N_14156);
or U14254 (N_14254,N_14060,N_14127);
and U14255 (N_14255,N_14228,N_14208);
nor U14256 (N_14256,N_14139,N_14203);
or U14257 (N_14257,N_14004,N_14131);
nand U14258 (N_14258,N_14165,N_14054);
nand U14259 (N_14259,N_14021,N_14126);
nor U14260 (N_14260,N_14171,N_14159);
or U14261 (N_14261,N_14006,N_14176);
nor U14262 (N_14262,N_14026,N_14140);
and U14263 (N_14263,N_14245,N_14213);
or U14264 (N_14264,N_14145,N_14058);
xnor U14265 (N_14265,N_14078,N_14133);
nand U14266 (N_14266,N_14177,N_14040);
and U14267 (N_14267,N_14226,N_14023);
xnor U14268 (N_14268,N_14050,N_14205);
nor U14269 (N_14269,N_14034,N_14161);
or U14270 (N_14270,N_14076,N_14233);
and U14271 (N_14271,N_14020,N_14094);
nand U14272 (N_14272,N_14220,N_14243);
nand U14273 (N_14273,N_14013,N_14168);
xnor U14274 (N_14274,N_14137,N_14059);
xor U14275 (N_14275,N_14148,N_14120);
nor U14276 (N_14276,N_14005,N_14083);
xnor U14277 (N_14277,N_14108,N_14158);
nor U14278 (N_14278,N_14000,N_14167);
nor U14279 (N_14279,N_14093,N_14008);
xor U14280 (N_14280,N_14028,N_14182);
nor U14281 (N_14281,N_14101,N_14244);
or U14282 (N_14282,N_14135,N_14218);
nor U14283 (N_14283,N_14194,N_14051);
and U14284 (N_14284,N_14068,N_14104);
nand U14285 (N_14285,N_14019,N_14121);
nor U14286 (N_14286,N_14045,N_14240);
xnor U14287 (N_14287,N_14200,N_14009);
or U14288 (N_14288,N_14085,N_14112);
and U14289 (N_14289,N_14173,N_14081);
nor U14290 (N_14290,N_14061,N_14149);
nor U14291 (N_14291,N_14105,N_14232);
nand U14292 (N_14292,N_14039,N_14215);
and U14293 (N_14293,N_14113,N_14190);
nand U14294 (N_14294,N_14248,N_14099);
nand U14295 (N_14295,N_14166,N_14214);
nand U14296 (N_14296,N_14064,N_14098);
nor U14297 (N_14297,N_14151,N_14091);
and U14298 (N_14298,N_14185,N_14241);
and U14299 (N_14299,N_14206,N_14152);
or U14300 (N_14300,N_14236,N_14238);
and U14301 (N_14301,N_14041,N_14077);
or U14302 (N_14302,N_14056,N_14191);
nor U14303 (N_14303,N_14016,N_14202);
nand U14304 (N_14304,N_14002,N_14169);
nor U14305 (N_14305,N_14038,N_14037);
nand U14306 (N_14306,N_14010,N_14178);
nand U14307 (N_14307,N_14119,N_14162);
or U14308 (N_14308,N_14219,N_14193);
nand U14309 (N_14309,N_14029,N_14181);
xnor U14310 (N_14310,N_14007,N_14087);
xor U14311 (N_14311,N_14079,N_14199);
or U14312 (N_14312,N_14142,N_14147);
xnor U14313 (N_14313,N_14097,N_14103);
nand U14314 (N_14314,N_14227,N_14216);
nand U14315 (N_14315,N_14192,N_14183);
or U14316 (N_14316,N_14170,N_14231);
or U14317 (N_14317,N_14035,N_14141);
xnor U14318 (N_14318,N_14046,N_14044);
nor U14319 (N_14319,N_14164,N_14117);
and U14320 (N_14320,N_14242,N_14128);
xnor U14321 (N_14321,N_14249,N_14211);
and U14322 (N_14322,N_14033,N_14017);
or U14323 (N_14323,N_14100,N_14184);
nand U14324 (N_14324,N_14247,N_14110);
xor U14325 (N_14325,N_14143,N_14073);
xnor U14326 (N_14326,N_14042,N_14221);
nand U14327 (N_14327,N_14053,N_14025);
nor U14328 (N_14328,N_14003,N_14130);
xor U14329 (N_14329,N_14111,N_14123);
or U14330 (N_14330,N_14230,N_14048);
nor U14331 (N_14331,N_14057,N_14114);
nor U14332 (N_14332,N_14052,N_14070);
nand U14333 (N_14333,N_14102,N_14155);
and U14334 (N_14334,N_14090,N_14204);
nor U14335 (N_14335,N_14012,N_14172);
nand U14336 (N_14336,N_14237,N_14154);
and U14337 (N_14337,N_14031,N_14197);
nor U14338 (N_14338,N_14179,N_14001);
or U14339 (N_14339,N_14062,N_14174);
xor U14340 (N_14340,N_14049,N_14136);
or U14341 (N_14341,N_14234,N_14217);
nor U14342 (N_14342,N_14067,N_14187);
nand U14343 (N_14343,N_14160,N_14235);
or U14344 (N_14344,N_14144,N_14088);
or U14345 (N_14345,N_14022,N_14080);
nor U14346 (N_14346,N_14129,N_14118);
and U14347 (N_14347,N_14089,N_14207);
and U14348 (N_14348,N_14163,N_14095);
or U14349 (N_14349,N_14134,N_14246);
and U14350 (N_14350,N_14015,N_14069);
nor U14351 (N_14351,N_14225,N_14096);
and U14352 (N_14352,N_14224,N_14212);
or U14353 (N_14353,N_14071,N_14109);
and U14354 (N_14354,N_14124,N_14072);
nand U14355 (N_14355,N_14063,N_14222);
and U14356 (N_14356,N_14122,N_14014);
and U14357 (N_14357,N_14107,N_14229);
nor U14358 (N_14358,N_14157,N_14210);
nand U14359 (N_14359,N_14074,N_14066);
and U14360 (N_14360,N_14198,N_14043);
xnor U14361 (N_14361,N_14153,N_14036);
nand U14362 (N_14362,N_14084,N_14018);
nor U14363 (N_14363,N_14146,N_14189);
or U14364 (N_14364,N_14150,N_14106);
or U14365 (N_14365,N_14024,N_14196);
xor U14366 (N_14366,N_14027,N_14175);
nor U14367 (N_14367,N_14075,N_14011);
and U14368 (N_14368,N_14188,N_14055);
nor U14369 (N_14369,N_14086,N_14030);
xor U14370 (N_14370,N_14115,N_14223);
xnor U14371 (N_14371,N_14132,N_14125);
or U14372 (N_14372,N_14186,N_14138);
and U14373 (N_14373,N_14239,N_14032);
xnor U14374 (N_14374,N_14047,N_14195);
nor U14375 (N_14375,N_14055,N_14155);
nand U14376 (N_14376,N_14069,N_14077);
nand U14377 (N_14377,N_14199,N_14096);
or U14378 (N_14378,N_14135,N_14132);
and U14379 (N_14379,N_14033,N_14052);
xnor U14380 (N_14380,N_14113,N_14075);
and U14381 (N_14381,N_14140,N_14086);
xor U14382 (N_14382,N_14238,N_14198);
nand U14383 (N_14383,N_14059,N_14121);
nand U14384 (N_14384,N_14035,N_14011);
and U14385 (N_14385,N_14215,N_14019);
nor U14386 (N_14386,N_14165,N_14090);
nor U14387 (N_14387,N_14042,N_14025);
or U14388 (N_14388,N_14176,N_14080);
and U14389 (N_14389,N_14163,N_14099);
and U14390 (N_14390,N_14089,N_14063);
xnor U14391 (N_14391,N_14047,N_14166);
or U14392 (N_14392,N_14172,N_14214);
or U14393 (N_14393,N_14057,N_14094);
xnor U14394 (N_14394,N_14139,N_14120);
nor U14395 (N_14395,N_14127,N_14227);
or U14396 (N_14396,N_14043,N_14050);
nor U14397 (N_14397,N_14107,N_14238);
nor U14398 (N_14398,N_14134,N_14038);
nor U14399 (N_14399,N_14093,N_14157);
nor U14400 (N_14400,N_14069,N_14043);
nand U14401 (N_14401,N_14131,N_14164);
xor U14402 (N_14402,N_14059,N_14044);
xnor U14403 (N_14403,N_14082,N_14100);
and U14404 (N_14404,N_14114,N_14229);
or U14405 (N_14405,N_14144,N_14007);
and U14406 (N_14406,N_14172,N_14077);
xnor U14407 (N_14407,N_14046,N_14239);
xor U14408 (N_14408,N_14118,N_14178);
and U14409 (N_14409,N_14172,N_14209);
xnor U14410 (N_14410,N_14083,N_14023);
nand U14411 (N_14411,N_14043,N_14032);
or U14412 (N_14412,N_14121,N_14226);
or U14413 (N_14413,N_14028,N_14136);
or U14414 (N_14414,N_14007,N_14100);
nor U14415 (N_14415,N_14223,N_14104);
xor U14416 (N_14416,N_14195,N_14238);
nor U14417 (N_14417,N_14210,N_14130);
xnor U14418 (N_14418,N_14147,N_14073);
nor U14419 (N_14419,N_14034,N_14134);
and U14420 (N_14420,N_14170,N_14094);
xor U14421 (N_14421,N_14025,N_14236);
nand U14422 (N_14422,N_14146,N_14007);
xnor U14423 (N_14423,N_14040,N_14239);
and U14424 (N_14424,N_14054,N_14006);
xnor U14425 (N_14425,N_14064,N_14113);
or U14426 (N_14426,N_14167,N_14150);
or U14427 (N_14427,N_14194,N_14146);
xnor U14428 (N_14428,N_14092,N_14108);
nand U14429 (N_14429,N_14050,N_14099);
or U14430 (N_14430,N_14220,N_14042);
nor U14431 (N_14431,N_14010,N_14047);
nor U14432 (N_14432,N_14248,N_14174);
xor U14433 (N_14433,N_14133,N_14091);
nand U14434 (N_14434,N_14123,N_14166);
nor U14435 (N_14435,N_14132,N_14106);
xor U14436 (N_14436,N_14145,N_14008);
and U14437 (N_14437,N_14152,N_14047);
or U14438 (N_14438,N_14042,N_14084);
and U14439 (N_14439,N_14200,N_14122);
nand U14440 (N_14440,N_14053,N_14034);
xnor U14441 (N_14441,N_14076,N_14023);
and U14442 (N_14442,N_14037,N_14191);
and U14443 (N_14443,N_14153,N_14051);
xnor U14444 (N_14444,N_14017,N_14092);
xnor U14445 (N_14445,N_14008,N_14070);
or U14446 (N_14446,N_14058,N_14035);
nand U14447 (N_14447,N_14037,N_14053);
or U14448 (N_14448,N_14192,N_14245);
and U14449 (N_14449,N_14172,N_14197);
xor U14450 (N_14450,N_14197,N_14174);
nor U14451 (N_14451,N_14162,N_14135);
nor U14452 (N_14452,N_14001,N_14038);
and U14453 (N_14453,N_14095,N_14074);
xor U14454 (N_14454,N_14039,N_14020);
nand U14455 (N_14455,N_14146,N_14064);
or U14456 (N_14456,N_14099,N_14226);
nor U14457 (N_14457,N_14175,N_14070);
and U14458 (N_14458,N_14134,N_14088);
or U14459 (N_14459,N_14191,N_14024);
or U14460 (N_14460,N_14054,N_14172);
nand U14461 (N_14461,N_14015,N_14032);
nor U14462 (N_14462,N_14193,N_14083);
xor U14463 (N_14463,N_14156,N_14215);
or U14464 (N_14464,N_14216,N_14015);
nand U14465 (N_14465,N_14065,N_14247);
and U14466 (N_14466,N_14013,N_14098);
and U14467 (N_14467,N_14071,N_14229);
or U14468 (N_14468,N_14177,N_14201);
nand U14469 (N_14469,N_14119,N_14221);
nand U14470 (N_14470,N_14220,N_14194);
or U14471 (N_14471,N_14162,N_14016);
or U14472 (N_14472,N_14216,N_14105);
nor U14473 (N_14473,N_14011,N_14030);
or U14474 (N_14474,N_14246,N_14247);
nor U14475 (N_14475,N_14235,N_14233);
nand U14476 (N_14476,N_14116,N_14179);
nor U14477 (N_14477,N_14137,N_14249);
nor U14478 (N_14478,N_14161,N_14025);
nand U14479 (N_14479,N_14232,N_14041);
or U14480 (N_14480,N_14145,N_14246);
and U14481 (N_14481,N_14010,N_14229);
nor U14482 (N_14482,N_14121,N_14225);
xor U14483 (N_14483,N_14141,N_14046);
nand U14484 (N_14484,N_14214,N_14044);
and U14485 (N_14485,N_14059,N_14012);
nor U14486 (N_14486,N_14062,N_14124);
nand U14487 (N_14487,N_14094,N_14192);
nor U14488 (N_14488,N_14104,N_14187);
xnor U14489 (N_14489,N_14119,N_14100);
or U14490 (N_14490,N_14162,N_14107);
and U14491 (N_14491,N_14150,N_14247);
xor U14492 (N_14492,N_14077,N_14192);
xnor U14493 (N_14493,N_14206,N_14126);
and U14494 (N_14494,N_14233,N_14125);
nand U14495 (N_14495,N_14171,N_14151);
and U14496 (N_14496,N_14132,N_14034);
nand U14497 (N_14497,N_14157,N_14058);
nand U14498 (N_14498,N_14049,N_14114);
and U14499 (N_14499,N_14142,N_14084);
and U14500 (N_14500,N_14298,N_14378);
and U14501 (N_14501,N_14467,N_14440);
nor U14502 (N_14502,N_14287,N_14497);
or U14503 (N_14503,N_14261,N_14426);
or U14504 (N_14504,N_14420,N_14358);
nand U14505 (N_14505,N_14297,N_14371);
and U14506 (N_14506,N_14390,N_14409);
xor U14507 (N_14507,N_14485,N_14385);
and U14508 (N_14508,N_14353,N_14416);
or U14509 (N_14509,N_14293,N_14320);
nand U14510 (N_14510,N_14269,N_14337);
or U14511 (N_14511,N_14423,N_14427);
and U14512 (N_14512,N_14363,N_14252);
or U14513 (N_14513,N_14498,N_14254);
xor U14514 (N_14514,N_14274,N_14352);
nor U14515 (N_14515,N_14400,N_14301);
or U14516 (N_14516,N_14311,N_14266);
nor U14517 (N_14517,N_14288,N_14442);
xnor U14518 (N_14518,N_14418,N_14435);
or U14519 (N_14519,N_14333,N_14495);
nand U14520 (N_14520,N_14398,N_14460);
and U14521 (N_14521,N_14391,N_14429);
or U14522 (N_14522,N_14468,N_14472);
or U14523 (N_14523,N_14313,N_14268);
nand U14524 (N_14524,N_14312,N_14493);
or U14525 (N_14525,N_14372,N_14331);
nor U14526 (N_14526,N_14306,N_14368);
and U14527 (N_14527,N_14470,N_14258);
nor U14528 (N_14528,N_14439,N_14402);
nor U14529 (N_14529,N_14308,N_14291);
xor U14530 (N_14530,N_14373,N_14351);
nand U14531 (N_14531,N_14355,N_14335);
nor U14532 (N_14532,N_14316,N_14421);
nand U14533 (N_14533,N_14336,N_14449);
nand U14534 (N_14534,N_14419,N_14469);
nand U14535 (N_14535,N_14341,N_14284);
or U14536 (N_14536,N_14422,N_14270);
nor U14537 (N_14537,N_14477,N_14319);
or U14538 (N_14538,N_14272,N_14366);
nand U14539 (N_14539,N_14453,N_14417);
xnor U14540 (N_14540,N_14326,N_14434);
nor U14541 (N_14541,N_14486,N_14489);
xnor U14542 (N_14542,N_14443,N_14410);
or U14543 (N_14543,N_14299,N_14340);
nand U14544 (N_14544,N_14359,N_14323);
nor U14545 (N_14545,N_14476,N_14310);
and U14546 (N_14546,N_14413,N_14321);
nor U14547 (N_14547,N_14357,N_14492);
nor U14548 (N_14548,N_14346,N_14380);
nand U14549 (N_14549,N_14496,N_14264);
nand U14550 (N_14550,N_14322,N_14295);
and U14551 (N_14551,N_14432,N_14389);
nand U14552 (N_14552,N_14479,N_14354);
xor U14553 (N_14553,N_14394,N_14275);
and U14554 (N_14554,N_14456,N_14415);
and U14555 (N_14555,N_14464,N_14364);
nor U14556 (N_14556,N_14392,N_14414);
or U14557 (N_14557,N_14474,N_14330);
or U14558 (N_14558,N_14289,N_14280);
and U14559 (N_14559,N_14370,N_14339);
or U14560 (N_14560,N_14437,N_14487);
xnor U14561 (N_14561,N_14307,N_14428);
and U14562 (N_14562,N_14447,N_14296);
and U14563 (N_14563,N_14475,N_14405);
xor U14564 (N_14564,N_14488,N_14267);
or U14565 (N_14565,N_14325,N_14494);
and U14566 (N_14566,N_14360,N_14404);
nand U14567 (N_14567,N_14256,N_14290);
or U14568 (N_14568,N_14292,N_14436);
nand U14569 (N_14569,N_14463,N_14384);
nand U14570 (N_14570,N_14318,N_14441);
nor U14571 (N_14571,N_14431,N_14455);
nor U14572 (N_14572,N_14406,N_14396);
nor U14573 (N_14573,N_14309,N_14263);
or U14574 (N_14574,N_14257,N_14304);
or U14575 (N_14575,N_14315,N_14303);
and U14576 (N_14576,N_14327,N_14262);
nor U14577 (N_14577,N_14490,N_14438);
xor U14578 (N_14578,N_14278,N_14273);
nand U14579 (N_14579,N_14491,N_14407);
and U14580 (N_14580,N_14411,N_14412);
nand U14581 (N_14581,N_14328,N_14347);
or U14582 (N_14582,N_14334,N_14349);
xnor U14583 (N_14583,N_14343,N_14369);
or U14584 (N_14584,N_14361,N_14381);
xnor U14585 (N_14585,N_14271,N_14260);
and U14586 (N_14586,N_14379,N_14403);
xor U14587 (N_14587,N_14365,N_14458);
and U14588 (N_14588,N_14374,N_14387);
nor U14589 (N_14589,N_14450,N_14338);
xor U14590 (N_14590,N_14300,N_14277);
nand U14591 (N_14591,N_14281,N_14383);
and U14592 (N_14592,N_14285,N_14459);
xor U14593 (N_14593,N_14377,N_14481);
or U14594 (N_14594,N_14433,N_14342);
xnor U14595 (N_14595,N_14283,N_14276);
xor U14596 (N_14596,N_14305,N_14345);
xnor U14597 (N_14597,N_14484,N_14465);
nand U14598 (N_14598,N_14317,N_14452);
or U14599 (N_14599,N_14265,N_14253);
or U14600 (N_14600,N_14448,N_14457);
or U14601 (N_14601,N_14473,N_14302);
nand U14602 (N_14602,N_14444,N_14499);
xnor U14603 (N_14603,N_14279,N_14362);
nor U14604 (N_14604,N_14401,N_14375);
xor U14605 (N_14605,N_14356,N_14255);
and U14606 (N_14606,N_14397,N_14399);
nand U14607 (N_14607,N_14329,N_14382);
and U14608 (N_14608,N_14430,N_14259);
or U14609 (N_14609,N_14348,N_14466);
xor U14610 (N_14610,N_14408,N_14367);
or U14611 (N_14611,N_14250,N_14451);
and U14612 (N_14612,N_14332,N_14251);
xnor U14613 (N_14613,N_14480,N_14386);
and U14614 (N_14614,N_14388,N_14478);
nand U14615 (N_14615,N_14314,N_14324);
nor U14616 (N_14616,N_14344,N_14393);
xnor U14617 (N_14617,N_14294,N_14483);
or U14618 (N_14618,N_14446,N_14454);
xnor U14619 (N_14619,N_14424,N_14286);
nand U14620 (N_14620,N_14461,N_14482);
xor U14621 (N_14621,N_14376,N_14350);
nand U14622 (N_14622,N_14425,N_14462);
nand U14623 (N_14623,N_14282,N_14445);
nand U14624 (N_14624,N_14395,N_14471);
xor U14625 (N_14625,N_14481,N_14269);
nor U14626 (N_14626,N_14333,N_14272);
xnor U14627 (N_14627,N_14410,N_14361);
nand U14628 (N_14628,N_14353,N_14357);
xor U14629 (N_14629,N_14343,N_14408);
and U14630 (N_14630,N_14280,N_14279);
xnor U14631 (N_14631,N_14336,N_14367);
xor U14632 (N_14632,N_14469,N_14439);
xor U14633 (N_14633,N_14293,N_14298);
nor U14634 (N_14634,N_14414,N_14283);
and U14635 (N_14635,N_14454,N_14331);
or U14636 (N_14636,N_14351,N_14450);
and U14637 (N_14637,N_14406,N_14259);
or U14638 (N_14638,N_14291,N_14370);
and U14639 (N_14639,N_14373,N_14287);
nand U14640 (N_14640,N_14329,N_14365);
or U14641 (N_14641,N_14345,N_14376);
nand U14642 (N_14642,N_14452,N_14357);
nand U14643 (N_14643,N_14458,N_14491);
nand U14644 (N_14644,N_14314,N_14445);
xnor U14645 (N_14645,N_14400,N_14434);
or U14646 (N_14646,N_14382,N_14390);
nand U14647 (N_14647,N_14252,N_14442);
xnor U14648 (N_14648,N_14302,N_14279);
xor U14649 (N_14649,N_14313,N_14388);
and U14650 (N_14650,N_14305,N_14395);
nor U14651 (N_14651,N_14342,N_14336);
and U14652 (N_14652,N_14316,N_14344);
nor U14653 (N_14653,N_14477,N_14357);
nand U14654 (N_14654,N_14472,N_14442);
nand U14655 (N_14655,N_14490,N_14409);
or U14656 (N_14656,N_14378,N_14371);
and U14657 (N_14657,N_14451,N_14284);
and U14658 (N_14658,N_14291,N_14348);
nand U14659 (N_14659,N_14498,N_14395);
and U14660 (N_14660,N_14468,N_14271);
or U14661 (N_14661,N_14296,N_14433);
or U14662 (N_14662,N_14438,N_14301);
or U14663 (N_14663,N_14469,N_14343);
and U14664 (N_14664,N_14285,N_14333);
nand U14665 (N_14665,N_14342,N_14434);
xnor U14666 (N_14666,N_14358,N_14446);
or U14667 (N_14667,N_14395,N_14366);
nand U14668 (N_14668,N_14458,N_14405);
xor U14669 (N_14669,N_14255,N_14312);
or U14670 (N_14670,N_14387,N_14379);
or U14671 (N_14671,N_14487,N_14476);
or U14672 (N_14672,N_14298,N_14364);
nor U14673 (N_14673,N_14384,N_14478);
and U14674 (N_14674,N_14392,N_14335);
or U14675 (N_14675,N_14462,N_14450);
nor U14676 (N_14676,N_14293,N_14474);
nor U14677 (N_14677,N_14417,N_14404);
nor U14678 (N_14678,N_14279,N_14329);
or U14679 (N_14679,N_14288,N_14463);
nor U14680 (N_14680,N_14434,N_14362);
and U14681 (N_14681,N_14297,N_14274);
nand U14682 (N_14682,N_14273,N_14258);
and U14683 (N_14683,N_14275,N_14310);
and U14684 (N_14684,N_14487,N_14373);
or U14685 (N_14685,N_14446,N_14260);
or U14686 (N_14686,N_14324,N_14497);
nor U14687 (N_14687,N_14474,N_14375);
nor U14688 (N_14688,N_14318,N_14442);
and U14689 (N_14689,N_14494,N_14316);
nor U14690 (N_14690,N_14334,N_14278);
and U14691 (N_14691,N_14404,N_14286);
nand U14692 (N_14692,N_14321,N_14472);
nor U14693 (N_14693,N_14430,N_14440);
and U14694 (N_14694,N_14478,N_14273);
nand U14695 (N_14695,N_14321,N_14442);
xor U14696 (N_14696,N_14392,N_14300);
xor U14697 (N_14697,N_14404,N_14401);
or U14698 (N_14698,N_14381,N_14345);
nand U14699 (N_14699,N_14476,N_14414);
xnor U14700 (N_14700,N_14310,N_14489);
and U14701 (N_14701,N_14451,N_14348);
nor U14702 (N_14702,N_14268,N_14264);
and U14703 (N_14703,N_14377,N_14270);
xor U14704 (N_14704,N_14342,N_14295);
nor U14705 (N_14705,N_14407,N_14498);
xor U14706 (N_14706,N_14420,N_14492);
or U14707 (N_14707,N_14366,N_14279);
nor U14708 (N_14708,N_14425,N_14469);
or U14709 (N_14709,N_14355,N_14310);
xnor U14710 (N_14710,N_14439,N_14316);
or U14711 (N_14711,N_14386,N_14437);
nor U14712 (N_14712,N_14475,N_14467);
nor U14713 (N_14713,N_14381,N_14259);
nand U14714 (N_14714,N_14294,N_14285);
nor U14715 (N_14715,N_14367,N_14384);
nor U14716 (N_14716,N_14445,N_14252);
and U14717 (N_14717,N_14294,N_14422);
or U14718 (N_14718,N_14403,N_14482);
and U14719 (N_14719,N_14398,N_14363);
nor U14720 (N_14720,N_14320,N_14332);
or U14721 (N_14721,N_14252,N_14289);
nand U14722 (N_14722,N_14496,N_14406);
xnor U14723 (N_14723,N_14314,N_14261);
nand U14724 (N_14724,N_14443,N_14415);
xor U14725 (N_14725,N_14368,N_14280);
nand U14726 (N_14726,N_14492,N_14263);
nand U14727 (N_14727,N_14305,N_14410);
xnor U14728 (N_14728,N_14402,N_14420);
and U14729 (N_14729,N_14257,N_14481);
nor U14730 (N_14730,N_14482,N_14324);
xnor U14731 (N_14731,N_14363,N_14274);
and U14732 (N_14732,N_14296,N_14283);
or U14733 (N_14733,N_14307,N_14427);
xnor U14734 (N_14734,N_14312,N_14302);
or U14735 (N_14735,N_14329,N_14389);
and U14736 (N_14736,N_14288,N_14318);
or U14737 (N_14737,N_14339,N_14265);
and U14738 (N_14738,N_14311,N_14321);
xor U14739 (N_14739,N_14480,N_14483);
xnor U14740 (N_14740,N_14414,N_14315);
xor U14741 (N_14741,N_14415,N_14353);
or U14742 (N_14742,N_14255,N_14329);
xnor U14743 (N_14743,N_14455,N_14468);
nor U14744 (N_14744,N_14255,N_14432);
and U14745 (N_14745,N_14256,N_14398);
nor U14746 (N_14746,N_14270,N_14486);
nand U14747 (N_14747,N_14430,N_14359);
and U14748 (N_14748,N_14472,N_14257);
nor U14749 (N_14749,N_14365,N_14325);
or U14750 (N_14750,N_14522,N_14702);
or U14751 (N_14751,N_14723,N_14692);
nor U14752 (N_14752,N_14517,N_14675);
nor U14753 (N_14753,N_14715,N_14547);
and U14754 (N_14754,N_14706,N_14623);
nor U14755 (N_14755,N_14591,N_14653);
nor U14756 (N_14756,N_14681,N_14589);
nand U14757 (N_14757,N_14611,N_14663);
and U14758 (N_14758,N_14534,N_14540);
and U14759 (N_14759,N_14575,N_14695);
or U14760 (N_14760,N_14531,N_14701);
xnor U14761 (N_14761,N_14552,N_14605);
xnor U14762 (N_14762,N_14713,N_14501);
and U14763 (N_14763,N_14543,N_14510);
or U14764 (N_14764,N_14674,N_14544);
and U14765 (N_14765,N_14724,N_14705);
and U14766 (N_14766,N_14731,N_14728);
or U14767 (N_14767,N_14580,N_14603);
or U14768 (N_14768,N_14505,N_14683);
or U14769 (N_14769,N_14631,N_14635);
or U14770 (N_14770,N_14642,N_14610);
nand U14771 (N_14771,N_14722,N_14703);
and U14772 (N_14772,N_14573,N_14585);
and U14773 (N_14773,N_14600,N_14710);
or U14774 (N_14774,N_14648,N_14684);
xor U14775 (N_14775,N_14595,N_14525);
nor U14776 (N_14776,N_14618,N_14739);
nand U14777 (N_14777,N_14545,N_14570);
or U14778 (N_14778,N_14614,N_14546);
and U14779 (N_14779,N_14554,N_14716);
or U14780 (N_14780,N_14569,N_14574);
xor U14781 (N_14781,N_14732,N_14500);
or U14782 (N_14782,N_14519,N_14561);
or U14783 (N_14783,N_14551,N_14572);
nor U14784 (N_14784,N_14733,N_14620);
nor U14785 (N_14785,N_14596,N_14530);
or U14786 (N_14786,N_14597,N_14639);
xor U14787 (N_14787,N_14735,N_14646);
nor U14788 (N_14788,N_14749,N_14748);
nor U14789 (N_14789,N_14521,N_14711);
nand U14790 (N_14790,N_14700,N_14557);
nand U14791 (N_14791,N_14651,N_14526);
or U14792 (N_14792,N_14677,N_14654);
nand U14793 (N_14793,N_14661,N_14649);
and U14794 (N_14794,N_14588,N_14587);
xor U14795 (N_14795,N_14687,N_14602);
nor U14796 (N_14796,N_14568,N_14613);
and U14797 (N_14797,N_14532,N_14536);
xor U14798 (N_14798,N_14523,N_14625);
and U14799 (N_14799,N_14657,N_14582);
or U14800 (N_14800,N_14662,N_14609);
or U14801 (N_14801,N_14528,N_14515);
or U14802 (N_14802,N_14563,N_14529);
xnor U14803 (N_14803,N_14607,N_14690);
nand U14804 (N_14804,N_14694,N_14542);
or U14805 (N_14805,N_14747,N_14727);
nand U14806 (N_14806,N_14558,N_14745);
or U14807 (N_14807,N_14619,N_14698);
and U14808 (N_14808,N_14640,N_14627);
or U14809 (N_14809,N_14629,N_14678);
or U14810 (N_14810,N_14506,N_14718);
or U14811 (N_14811,N_14664,N_14579);
xnor U14812 (N_14812,N_14553,N_14559);
nand U14813 (N_14813,N_14616,N_14746);
xnor U14814 (N_14814,N_14686,N_14508);
nor U14815 (N_14815,N_14633,N_14599);
xnor U14816 (N_14816,N_14697,N_14673);
nand U14817 (N_14817,N_14509,N_14571);
nand U14818 (N_14818,N_14712,N_14670);
xnor U14819 (N_14819,N_14556,N_14576);
nand U14820 (N_14820,N_14527,N_14583);
nor U14821 (N_14821,N_14626,N_14606);
and U14822 (N_14822,N_14699,N_14518);
or U14823 (N_14823,N_14688,N_14656);
nand U14824 (N_14824,N_14666,N_14691);
xor U14825 (N_14825,N_14562,N_14566);
xnor U14826 (N_14826,N_14630,N_14617);
nand U14827 (N_14827,N_14689,N_14734);
and U14828 (N_14828,N_14507,N_14720);
and U14829 (N_14829,N_14516,N_14560);
or U14830 (N_14830,N_14512,N_14520);
xor U14831 (N_14831,N_14502,N_14730);
and U14832 (N_14832,N_14696,N_14541);
xor U14833 (N_14833,N_14660,N_14671);
and U14834 (N_14834,N_14593,N_14628);
or U14835 (N_14835,N_14637,N_14638);
or U14836 (N_14836,N_14578,N_14717);
xor U14837 (N_14837,N_14707,N_14709);
xor U14838 (N_14838,N_14565,N_14719);
nor U14839 (N_14839,N_14511,N_14622);
nand U14840 (N_14840,N_14743,N_14721);
xor U14841 (N_14841,N_14704,N_14669);
nand U14842 (N_14842,N_14612,N_14598);
nor U14843 (N_14843,N_14655,N_14685);
nor U14844 (N_14844,N_14645,N_14592);
nor U14845 (N_14845,N_14736,N_14641);
xor U14846 (N_14846,N_14659,N_14535);
xnor U14847 (N_14847,N_14584,N_14567);
or U14848 (N_14848,N_14555,N_14524);
nor U14849 (N_14849,N_14676,N_14726);
or U14850 (N_14850,N_14740,N_14634);
nor U14851 (N_14851,N_14714,N_14608);
xnor U14852 (N_14852,N_14550,N_14621);
xor U14853 (N_14853,N_14725,N_14643);
nor U14854 (N_14854,N_14590,N_14514);
and U14855 (N_14855,N_14538,N_14665);
nand U14856 (N_14856,N_14658,N_14744);
xor U14857 (N_14857,N_14564,N_14668);
nand U14858 (N_14858,N_14737,N_14615);
and U14859 (N_14859,N_14644,N_14679);
or U14860 (N_14860,N_14680,N_14672);
nor U14861 (N_14861,N_14537,N_14581);
xnor U14862 (N_14862,N_14741,N_14594);
or U14863 (N_14863,N_14549,N_14650);
or U14864 (N_14864,N_14708,N_14738);
nand U14865 (N_14865,N_14729,N_14586);
nand U14866 (N_14866,N_14513,N_14577);
xnor U14867 (N_14867,N_14548,N_14742);
nand U14868 (N_14868,N_14693,N_14632);
xor U14869 (N_14869,N_14539,N_14647);
or U14870 (N_14870,N_14682,N_14503);
and U14871 (N_14871,N_14604,N_14652);
xor U14872 (N_14872,N_14533,N_14636);
or U14873 (N_14873,N_14624,N_14601);
or U14874 (N_14874,N_14504,N_14667);
nor U14875 (N_14875,N_14716,N_14526);
and U14876 (N_14876,N_14632,N_14515);
or U14877 (N_14877,N_14538,N_14585);
nor U14878 (N_14878,N_14612,N_14533);
nor U14879 (N_14879,N_14643,N_14645);
nand U14880 (N_14880,N_14554,N_14516);
xor U14881 (N_14881,N_14718,N_14569);
xor U14882 (N_14882,N_14655,N_14526);
or U14883 (N_14883,N_14619,N_14719);
xor U14884 (N_14884,N_14682,N_14623);
xor U14885 (N_14885,N_14548,N_14562);
or U14886 (N_14886,N_14528,N_14681);
nand U14887 (N_14887,N_14586,N_14675);
and U14888 (N_14888,N_14601,N_14604);
xor U14889 (N_14889,N_14603,N_14622);
and U14890 (N_14890,N_14674,N_14500);
xor U14891 (N_14891,N_14556,N_14666);
or U14892 (N_14892,N_14631,N_14548);
or U14893 (N_14893,N_14598,N_14625);
nor U14894 (N_14894,N_14667,N_14709);
nor U14895 (N_14895,N_14690,N_14709);
nor U14896 (N_14896,N_14660,N_14576);
and U14897 (N_14897,N_14721,N_14706);
nor U14898 (N_14898,N_14589,N_14697);
xnor U14899 (N_14899,N_14577,N_14647);
and U14900 (N_14900,N_14578,N_14551);
xor U14901 (N_14901,N_14633,N_14630);
nand U14902 (N_14902,N_14593,N_14604);
xnor U14903 (N_14903,N_14734,N_14590);
nor U14904 (N_14904,N_14679,N_14582);
and U14905 (N_14905,N_14590,N_14693);
or U14906 (N_14906,N_14626,N_14633);
nor U14907 (N_14907,N_14523,N_14630);
nand U14908 (N_14908,N_14704,N_14541);
xnor U14909 (N_14909,N_14507,N_14739);
nand U14910 (N_14910,N_14521,N_14678);
xnor U14911 (N_14911,N_14548,N_14529);
nor U14912 (N_14912,N_14578,N_14715);
nand U14913 (N_14913,N_14701,N_14638);
or U14914 (N_14914,N_14749,N_14662);
or U14915 (N_14915,N_14563,N_14631);
nand U14916 (N_14916,N_14683,N_14632);
or U14917 (N_14917,N_14717,N_14608);
nand U14918 (N_14918,N_14668,N_14535);
xnor U14919 (N_14919,N_14589,N_14546);
or U14920 (N_14920,N_14562,N_14545);
or U14921 (N_14921,N_14585,N_14565);
and U14922 (N_14922,N_14615,N_14511);
or U14923 (N_14923,N_14620,N_14664);
or U14924 (N_14924,N_14697,N_14723);
xnor U14925 (N_14925,N_14686,N_14524);
nor U14926 (N_14926,N_14596,N_14638);
nand U14927 (N_14927,N_14572,N_14532);
nor U14928 (N_14928,N_14541,N_14667);
nand U14929 (N_14929,N_14582,N_14501);
and U14930 (N_14930,N_14640,N_14737);
nor U14931 (N_14931,N_14524,N_14715);
nand U14932 (N_14932,N_14528,N_14656);
and U14933 (N_14933,N_14535,N_14728);
nor U14934 (N_14934,N_14610,N_14736);
xor U14935 (N_14935,N_14524,N_14742);
or U14936 (N_14936,N_14661,N_14683);
nand U14937 (N_14937,N_14730,N_14682);
nand U14938 (N_14938,N_14563,N_14503);
nand U14939 (N_14939,N_14687,N_14627);
nor U14940 (N_14940,N_14575,N_14749);
xor U14941 (N_14941,N_14593,N_14539);
or U14942 (N_14942,N_14603,N_14591);
or U14943 (N_14943,N_14613,N_14693);
xor U14944 (N_14944,N_14526,N_14571);
or U14945 (N_14945,N_14602,N_14739);
and U14946 (N_14946,N_14543,N_14578);
and U14947 (N_14947,N_14686,N_14600);
nor U14948 (N_14948,N_14640,N_14583);
nand U14949 (N_14949,N_14636,N_14669);
and U14950 (N_14950,N_14704,N_14553);
nor U14951 (N_14951,N_14650,N_14508);
nor U14952 (N_14952,N_14643,N_14603);
xnor U14953 (N_14953,N_14591,N_14657);
and U14954 (N_14954,N_14747,N_14596);
or U14955 (N_14955,N_14614,N_14728);
or U14956 (N_14956,N_14651,N_14503);
nand U14957 (N_14957,N_14618,N_14683);
xor U14958 (N_14958,N_14594,N_14664);
xnor U14959 (N_14959,N_14621,N_14700);
or U14960 (N_14960,N_14711,N_14500);
nor U14961 (N_14961,N_14703,N_14700);
nand U14962 (N_14962,N_14518,N_14743);
or U14963 (N_14963,N_14548,N_14564);
nand U14964 (N_14964,N_14738,N_14589);
or U14965 (N_14965,N_14616,N_14638);
xor U14966 (N_14966,N_14728,N_14638);
xnor U14967 (N_14967,N_14746,N_14598);
or U14968 (N_14968,N_14512,N_14658);
nor U14969 (N_14969,N_14569,N_14669);
or U14970 (N_14970,N_14586,N_14517);
nand U14971 (N_14971,N_14619,N_14516);
xor U14972 (N_14972,N_14582,N_14619);
nand U14973 (N_14973,N_14607,N_14661);
xor U14974 (N_14974,N_14604,N_14713);
nor U14975 (N_14975,N_14613,N_14684);
xnor U14976 (N_14976,N_14622,N_14662);
and U14977 (N_14977,N_14623,N_14527);
and U14978 (N_14978,N_14501,N_14554);
nand U14979 (N_14979,N_14692,N_14687);
nand U14980 (N_14980,N_14522,N_14679);
nor U14981 (N_14981,N_14644,N_14721);
nand U14982 (N_14982,N_14514,N_14728);
xor U14983 (N_14983,N_14715,N_14573);
xnor U14984 (N_14984,N_14640,N_14607);
and U14985 (N_14985,N_14704,N_14649);
nor U14986 (N_14986,N_14602,N_14608);
or U14987 (N_14987,N_14683,N_14602);
or U14988 (N_14988,N_14527,N_14589);
nor U14989 (N_14989,N_14672,N_14589);
nor U14990 (N_14990,N_14705,N_14581);
nor U14991 (N_14991,N_14697,N_14748);
xor U14992 (N_14992,N_14727,N_14683);
xnor U14993 (N_14993,N_14508,N_14529);
nor U14994 (N_14994,N_14608,N_14660);
nand U14995 (N_14995,N_14724,N_14603);
xnor U14996 (N_14996,N_14572,N_14550);
and U14997 (N_14997,N_14512,N_14580);
nand U14998 (N_14998,N_14625,N_14618);
nand U14999 (N_14999,N_14596,N_14700);
or UO_0 (O_0,N_14763,N_14895);
nor UO_1 (O_1,N_14782,N_14794);
nand UO_2 (O_2,N_14831,N_14841);
or UO_3 (O_3,N_14828,N_14897);
or UO_4 (O_4,N_14864,N_14881);
nor UO_5 (O_5,N_14844,N_14961);
and UO_6 (O_6,N_14790,N_14944);
nor UO_7 (O_7,N_14914,N_14820);
nand UO_8 (O_8,N_14862,N_14918);
nor UO_9 (O_9,N_14755,N_14769);
nand UO_10 (O_10,N_14832,N_14974);
or UO_11 (O_11,N_14754,N_14967);
nor UO_12 (O_12,N_14929,N_14946);
and UO_13 (O_13,N_14893,N_14761);
nor UO_14 (O_14,N_14951,N_14882);
xnor UO_15 (O_15,N_14938,N_14924);
nor UO_16 (O_16,N_14861,N_14783);
xnor UO_17 (O_17,N_14953,N_14969);
xnor UO_18 (O_18,N_14982,N_14936);
nor UO_19 (O_19,N_14837,N_14856);
xor UO_20 (O_20,N_14973,N_14793);
xnor UO_21 (O_21,N_14989,N_14826);
xor UO_22 (O_22,N_14788,N_14883);
xnor UO_23 (O_23,N_14891,N_14752);
and UO_24 (O_24,N_14968,N_14771);
xor UO_25 (O_25,N_14906,N_14853);
xor UO_26 (O_26,N_14994,N_14834);
or UO_27 (O_27,N_14770,N_14902);
nand UO_28 (O_28,N_14935,N_14979);
xnor UO_29 (O_29,N_14933,N_14781);
nand UO_30 (O_30,N_14768,N_14889);
nor UO_31 (O_31,N_14996,N_14907);
nand UO_32 (O_32,N_14865,N_14877);
nor UO_33 (O_33,N_14803,N_14869);
or UO_34 (O_34,N_14776,N_14960);
or UO_35 (O_35,N_14899,N_14972);
nand UO_36 (O_36,N_14812,N_14981);
nand UO_37 (O_37,N_14821,N_14927);
nor UO_38 (O_38,N_14758,N_14926);
xor UO_39 (O_39,N_14859,N_14913);
nand UO_40 (O_40,N_14798,N_14995);
xor UO_41 (O_41,N_14930,N_14810);
nand UO_42 (O_42,N_14833,N_14966);
xnor UO_43 (O_43,N_14908,N_14779);
or UO_44 (O_44,N_14945,N_14774);
or UO_45 (O_45,N_14845,N_14958);
nor UO_46 (O_46,N_14800,N_14934);
nand UO_47 (O_47,N_14898,N_14963);
nor UO_48 (O_48,N_14848,N_14786);
nor UO_49 (O_49,N_14764,N_14809);
or UO_50 (O_50,N_14939,N_14797);
nor UO_51 (O_51,N_14796,N_14984);
nor UO_52 (O_52,N_14923,N_14959);
nand UO_53 (O_53,N_14816,N_14855);
or UO_54 (O_54,N_14920,N_14993);
nor UO_55 (O_55,N_14854,N_14785);
and UO_56 (O_56,N_14954,N_14866);
nand UO_57 (O_57,N_14840,N_14992);
nor UO_58 (O_58,N_14948,N_14870);
or UO_59 (O_59,N_14896,N_14756);
nor UO_60 (O_60,N_14892,N_14750);
or UO_61 (O_61,N_14991,N_14884);
nor UO_62 (O_62,N_14876,N_14775);
and UO_63 (O_63,N_14957,N_14911);
nor UO_64 (O_64,N_14767,N_14947);
xor UO_65 (O_65,N_14814,N_14867);
xnor UO_66 (O_66,N_14941,N_14807);
and UO_67 (O_67,N_14880,N_14751);
and UO_68 (O_68,N_14928,N_14910);
or UO_69 (O_69,N_14852,N_14952);
nand UO_70 (O_70,N_14795,N_14792);
or UO_71 (O_71,N_14773,N_14825);
or UO_72 (O_72,N_14894,N_14903);
xnor UO_73 (O_73,N_14842,N_14888);
nor UO_74 (O_74,N_14805,N_14789);
xnor UO_75 (O_75,N_14839,N_14931);
xor UO_76 (O_76,N_14824,N_14819);
or UO_77 (O_77,N_14971,N_14818);
or UO_78 (O_78,N_14940,N_14872);
xor UO_79 (O_79,N_14858,N_14843);
and UO_80 (O_80,N_14823,N_14829);
nand UO_81 (O_81,N_14804,N_14806);
and UO_82 (O_82,N_14977,N_14846);
and UO_83 (O_83,N_14922,N_14937);
and UO_84 (O_84,N_14916,N_14791);
nand UO_85 (O_85,N_14799,N_14813);
and UO_86 (O_86,N_14904,N_14850);
xnor UO_87 (O_87,N_14879,N_14925);
or UO_88 (O_88,N_14975,N_14900);
and UO_89 (O_89,N_14919,N_14836);
and UO_90 (O_90,N_14849,N_14838);
and UO_91 (O_91,N_14827,N_14987);
or UO_92 (O_92,N_14873,N_14983);
nand UO_93 (O_93,N_14878,N_14874);
nor UO_94 (O_94,N_14965,N_14871);
or UO_95 (O_95,N_14777,N_14988);
nand UO_96 (O_96,N_14921,N_14976);
or UO_97 (O_97,N_14980,N_14905);
and UO_98 (O_98,N_14885,N_14999);
nand UO_99 (O_99,N_14990,N_14998);
or UO_100 (O_100,N_14970,N_14890);
xor UO_101 (O_101,N_14863,N_14997);
and UO_102 (O_102,N_14753,N_14955);
or UO_103 (O_103,N_14942,N_14964);
or UO_104 (O_104,N_14986,N_14943);
and UO_105 (O_105,N_14802,N_14917);
nand UO_106 (O_106,N_14857,N_14817);
nor UO_107 (O_107,N_14801,N_14808);
nand UO_108 (O_108,N_14978,N_14860);
nand UO_109 (O_109,N_14830,N_14887);
xor UO_110 (O_110,N_14787,N_14912);
xnor UO_111 (O_111,N_14780,N_14778);
or UO_112 (O_112,N_14962,N_14762);
xnor UO_113 (O_113,N_14760,N_14847);
nor UO_114 (O_114,N_14886,N_14765);
nor UO_115 (O_115,N_14766,N_14851);
nand UO_116 (O_116,N_14811,N_14985);
nand UO_117 (O_117,N_14949,N_14784);
xnor UO_118 (O_118,N_14757,N_14868);
nor UO_119 (O_119,N_14822,N_14950);
xnor UO_120 (O_120,N_14956,N_14932);
nor UO_121 (O_121,N_14875,N_14909);
nor UO_122 (O_122,N_14901,N_14915);
and UO_123 (O_123,N_14835,N_14759);
xnor UO_124 (O_124,N_14815,N_14772);
nand UO_125 (O_125,N_14788,N_14782);
and UO_126 (O_126,N_14926,N_14894);
nand UO_127 (O_127,N_14898,N_14907);
nor UO_128 (O_128,N_14944,N_14844);
nor UO_129 (O_129,N_14784,N_14788);
and UO_130 (O_130,N_14757,N_14890);
or UO_131 (O_131,N_14865,N_14846);
and UO_132 (O_132,N_14906,N_14939);
xor UO_133 (O_133,N_14759,N_14755);
and UO_134 (O_134,N_14909,N_14881);
and UO_135 (O_135,N_14768,N_14990);
or UO_136 (O_136,N_14991,N_14849);
nand UO_137 (O_137,N_14909,N_14811);
and UO_138 (O_138,N_14812,N_14787);
or UO_139 (O_139,N_14811,N_14782);
and UO_140 (O_140,N_14797,N_14903);
and UO_141 (O_141,N_14844,N_14984);
or UO_142 (O_142,N_14979,N_14776);
xnor UO_143 (O_143,N_14974,N_14890);
nand UO_144 (O_144,N_14799,N_14777);
nor UO_145 (O_145,N_14966,N_14979);
nor UO_146 (O_146,N_14779,N_14932);
or UO_147 (O_147,N_14915,N_14774);
and UO_148 (O_148,N_14901,N_14937);
nand UO_149 (O_149,N_14785,N_14863);
xnor UO_150 (O_150,N_14922,N_14790);
and UO_151 (O_151,N_14830,N_14910);
nor UO_152 (O_152,N_14831,N_14918);
nor UO_153 (O_153,N_14879,N_14791);
and UO_154 (O_154,N_14846,N_14787);
nor UO_155 (O_155,N_14759,N_14932);
nor UO_156 (O_156,N_14843,N_14938);
and UO_157 (O_157,N_14914,N_14940);
xnor UO_158 (O_158,N_14950,N_14848);
nand UO_159 (O_159,N_14882,N_14959);
and UO_160 (O_160,N_14909,N_14896);
nand UO_161 (O_161,N_14850,N_14755);
nand UO_162 (O_162,N_14782,N_14892);
xnor UO_163 (O_163,N_14914,N_14811);
nand UO_164 (O_164,N_14859,N_14990);
or UO_165 (O_165,N_14872,N_14811);
nand UO_166 (O_166,N_14803,N_14976);
or UO_167 (O_167,N_14997,N_14865);
nor UO_168 (O_168,N_14975,N_14790);
nor UO_169 (O_169,N_14915,N_14762);
nor UO_170 (O_170,N_14918,N_14806);
xor UO_171 (O_171,N_14799,N_14790);
nor UO_172 (O_172,N_14929,N_14821);
or UO_173 (O_173,N_14937,N_14997);
nor UO_174 (O_174,N_14840,N_14969);
nor UO_175 (O_175,N_14911,N_14861);
or UO_176 (O_176,N_14885,N_14837);
nor UO_177 (O_177,N_14865,N_14977);
xor UO_178 (O_178,N_14860,N_14955);
xor UO_179 (O_179,N_14805,N_14943);
xor UO_180 (O_180,N_14968,N_14845);
nand UO_181 (O_181,N_14971,N_14839);
xnor UO_182 (O_182,N_14887,N_14995);
nor UO_183 (O_183,N_14958,N_14993);
nand UO_184 (O_184,N_14916,N_14855);
xnor UO_185 (O_185,N_14902,N_14954);
nor UO_186 (O_186,N_14891,N_14917);
and UO_187 (O_187,N_14878,N_14800);
and UO_188 (O_188,N_14801,N_14789);
and UO_189 (O_189,N_14960,N_14916);
nand UO_190 (O_190,N_14758,N_14978);
xor UO_191 (O_191,N_14948,N_14982);
nand UO_192 (O_192,N_14794,N_14836);
and UO_193 (O_193,N_14856,N_14962);
nand UO_194 (O_194,N_14978,N_14809);
and UO_195 (O_195,N_14966,N_14867);
and UO_196 (O_196,N_14801,N_14782);
nor UO_197 (O_197,N_14784,N_14969);
or UO_198 (O_198,N_14880,N_14776);
nand UO_199 (O_199,N_14806,N_14760);
and UO_200 (O_200,N_14957,N_14796);
nand UO_201 (O_201,N_14811,N_14930);
xnor UO_202 (O_202,N_14784,N_14812);
nand UO_203 (O_203,N_14853,N_14898);
and UO_204 (O_204,N_14764,N_14980);
and UO_205 (O_205,N_14823,N_14844);
or UO_206 (O_206,N_14976,N_14787);
nand UO_207 (O_207,N_14930,N_14987);
or UO_208 (O_208,N_14782,N_14799);
nor UO_209 (O_209,N_14971,N_14767);
nor UO_210 (O_210,N_14987,N_14870);
or UO_211 (O_211,N_14951,N_14866);
nor UO_212 (O_212,N_14835,N_14994);
and UO_213 (O_213,N_14915,N_14850);
and UO_214 (O_214,N_14754,N_14848);
or UO_215 (O_215,N_14819,N_14999);
nand UO_216 (O_216,N_14845,N_14758);
or UO_217 (O_217,N_14772,N_14943);
nor UO_218 (O_218,N_14900,N_14869);
xnor UO_219 (O_219,N_14962,N_14946);
nand UO_220 (O_220,N_14944,N_14983);
nor UO_221 (O_221,N_14976,N_14911);
nand UO_222 (O_222,N_14786,N_14912);
nand UO_223 (O_223,N_14932,N_14750);
nand UO_224 (O_224,N_14904,N_14805);
and UO_225 (O_225,N_14828,N_14809);
nand UO_226 (O_226,N_14771,N_14820);
xnor UO_227 (O_227,N_14778,N_14847);
nor UO_228 (O_228,N_14907,N_14847);
xnor UO_229 (O_229,N_14878,N_14756);
nand UO_230 (O_230,N_14804,N_14769);
nor UO_231 (O_231,N_14870,N_14851);
and UO_232 (O_232,N_14922,N_14926);
or UO_233 (O_233,N_14819,N_14959);
and UO_234 (O_234,N_14887,N_14764);
nor UO_235 (O_235,N_14957,N_14901);
nand UO_236 (O_236,N_14948,N_14760);
xnor UO_237 (O_237,N_14787,N_14999);
or UO_238 (O_238,N_14980,N_14940);
nand UO_239 (O_239,N_14951,N_14815);
nand UO_240 (O_240,N_14870,N_14822);
or UO_241 (O_241,N_14981,N_14777);
nand UO_242 (O_242,N_14969,N_14911);
and UO_243 (O_243,N_14811,N_14776);
and UO_244 (O_244,N_14810,N_14866);
xnor UO_245 (O_245,N_14862,N_14819);
or UO_246 (O_246,N_14918,N_14764);
or UO_247 (O_247,N_14914,N_14828);
xnor UO_248 (O_248,N_14942,N_14941);
and UO_249 (O_249,N_14825,N_14961);
nor UO_250 (O_250,N_14927,N_14907);
nor UO_251 (O_251,N_14994,N_14982);
xnor UO_252 (O_252,N_14828,N_14996);
and UO_253 (O_253,N_14874,N_14877);
or UO_254 (O_254,N_14789,N_14857);
nand UO_255 (O_255,N_14942,N_14798);
or UO_256 (O_256,N_14766,N_14957);
xnor UO_257 (O_257,N_14851,N_14849);
or UO_258 (O_258,N_14908,N_14763);
xnor UO_259 (O_259,N_14906,N_14965);
or UO_260 (O_260,N_14823,N_14894);
or UO_261 (O_261,N_14954,N_14986);
and UO_262 (O_262,N_14791,N_14932);
or UO_263 (O_263,N_14878,N_14873);
nand UO_264 (O_264,N_14824,N_14903);
and UO_265 (O_265,N_14983,N_14799);
nand UO_266 (O_266,N_14884,N_14961);
and UO_267 (O_267,N_14881,N_14891);
nor UO_268 (O_268,N_14934,N_14768);
nand UO_269 (O_269,N_14893,N_14882);
xnor UO_270 (O_270,N_14991,N_14904);
xnor UO_271 (O_271,N_14896,N_14951);
xnor UO_272 (O_272,N_14997,N_14926);
and UO_273 (O_273,N_14834,N_14891);
xor UO_274 (O_274,N_14957,N_14765);
and UO_275 (O_275,N_14826,N_14785);
nand UO_276 (O_276,N_14854,N_14831);
xnor UO_277 (O_277,N_14832,N_14925);
xnor UO_278 (O_278,N_14808,N_14999);
or UO_279 (O_279,N_14788,N_14764);
nor UO_280 (O_280,N_14900,N_14855);
or UO_281 (O_281,N_14897,N_14823);
xor UO_282 (O_282,N_14867,N_14979);
nand UO_283 (O_283,N_14982,N_14793);
nand UO_284 (O_284,N_14795,N_14754);
nand UO_285 (O_285,N_14751,N_14993);
or UO_286 (O_286,N_14938,N_14792);
xnor UO_287 (O_287,N_14971,N_14841);
or UO_288 (O_288,N_14929,N_14936);
xor UO_289 (O_289,N_14844,N_14879);
xnor UO_290 (O_290,N_14981,N_14824);
nor UO_291 (O_291,N_14917,N_14919);
and UO_292 (O_292,N_14984,N_14946);
or UO_293 (O_293,N_14920,N_14795);
or UO_294 (O_294,N_14785,N_14970);
nand UO_295 (O_295,N_14822,N_14929);
xnor UO_296 (O_296,N_14860,N_14782);
nor UO_297 (O_297,N_14758,N_14847);
and UO_298 (O_298,N_14778,N_14920);
nor UO_299 (O_299,N_14769,N_14831);
xor UO_300 (O_300,N_14899,N_14921);
and UO_301 (O_301,N_14982,N_14877);
or UO_302 (O_302,N_14807,N_14891);
xor UO_303 (O_303,N_14959,N_14801);
nand UO_304 (O_304,N_14780,N_14983);
and UO_305 (O_305,N_14810,N_14952);
xnor UO_306 (O_306,N_14794,N_14925);
and UO_307 (O_307,N_14849,N_14953);
and UO_308 (O_308,N_14846,N_14888);
nand UO_309 (O_309,N_14852,N_14768);
nand UO_310 (O_310,N_14841,N_14902);
and UO_311 (O_311,N_14971,N_14898);
xor UO_312 (O_312,N_14876,N_14871);
and UO_313 (O_313,N_14953,N_14777);
or UO_314 (O_314,N_14889,N_14995);
or UO_315 (O_315,N_14933,N_14779);
nand UO_316 (O_316,N_14869,N_14952);
nand UO_317 (O_317,N_14843,N_14840);
and UO_318 (O_318,N_14916,N_14934);
or UO_319 (O_319,N_14977,N_14827);
xor UO_320 (O_320,N_14971,N_14873);
and UO_321 (O_321,N_14933,N_14809);
xnor UO_322 (O_322,N_14814,N_14850);
and UO_323 (O_323,N_14994,N_14772);
nor UO_324 (O_324,N_14923,N_14794);
and UO_325 (O_325,N_14846,N_14812);
or UO_326 (O_326,N_14966,N_14800);
or UO_327 (O_327,N_14892,N_14964);
or UO_328 (O_328,N_14888,N_14824);
nand UO_329 (O_329,N_14759,N_14943);
or UO_330 (O_330,N_14976,N_14771);
or UO_331 (O_331,N_14961,N_14895);
xor UO_332 (O_332,N_14856,N_14903);
nor UO_333 (O_333,N_14863,N_14826);
nand UO_334 (O_334,N_14913,N_14901);
xnor UO_335 (O_335,N_14925,N_14758);
and UO_336 (O_336,N_14948,N_14778);
nor UO_337 (O_337,N_14788,N_14904);
or UO_338 (O_338,N_14788,N_14840);
nor UO_339 (O_339,N_14896,N_14822);
xnor UO_340 (O_340,N_14784,N_14927);
nand UO_341 (O_341,N_14793,N_14895);
xor UO_342 (O_342,N_14833,N_14981);
nor UO_343 (O_343,N_14957,N_14878);
xor UO_344 (O_344,N_14891,N_14901);
xnor UO_345 (O_345,N_14998,N_14757);
or UO_346 (O_346,N_14852,N_14835);
nand UO_347 (O_347,N_14936,N_14907);
xor UO_348 (O_348,N_14842,N_14786);
nor UO_349 (O_349,N_14890,N_14954);
or UO_350 (O_350,N_14822,N_14836);
nor UO_351 (O_351,N_14916,N_14976);
nor UO_352 (O_352,N_14937,N_14787);
nand UO_353 (O_353,N_14802,N_14797);
xor UO_354 (O_354,N_14767,N_14996);
or UO_355 (O_355,N_14951,N_14838);
or UO_356 (O_356,N_14868,N_14845);
nor UO_357 (O_357,N_14782,N_14757);
xor UO_358 (O_358,N_14895,N_14970);
or UO_359 (O_359,N_14921,N_14964);
and UO_360 (O_360,N_14981,N_14854);
xor UO_361 (O_361,N_14910,N_14920);
or UO_362 (O_362,N_14890,N_14896);
nor UO_363 (O_363,N_14765,N_14842);
and UO_364 (O_364,N_14838,N_14832);
nor UO_365 (O_365,N_14804,N_14943);
and UO_366 (O_366,N_14751,N_14828);
nor UO_367 (O_367,N_14945,N_14841);
or UO_368 (O_368,N_14869,N_14873);
or UO_369 (O_369,N_14854,N_14786);
and UO_370 (O_370,N_14996,N_14841);
and UO_371 (O_371,N_14797,N_14787);
nor UO_372 (O_372,N_14785,N_14758);
xnor UO_373 (O_373,N_14948,N_14937);
nand UO_374 (O_374,N_14990,N_14978);
and UO_375 (O_375,N_14784,N_14965);
or UO_376 (O_376,N_14772,N_14938);
nor UO_377 (O_377,N_14791,N_14995);
nand UO_378 (O_378,N_14871,N_14914);
or UO_379 (O_379,N_14810,N_14988);
nand UO_380 (O_380,N_14877,N_14853);
xor UO_381 (O_381,N_14788,N_14806);
nand UO_382 (O_382,N_14861,N_14781);
and UO_383 (O_383,N_14960,N_14961);
or UO_384 (O_384,N_14889,N_14847);
or UO_385 (O_385,N_14803,N_14867);
nand UO_386 (O_386,N_14934,N_14822);
nor UO_387 (O_387,N_14891,N_14813);
nand UO_388 (O_388,N_14898,N_14831);
xnor UO_389 (O_389,N_14773,N_14914);
nand UO_390 (O_390,N_14758,N_14876);
nor UO_391 (O_391,N_14830,N_14829);
nand UO_392 (O_392,N_14856,N_14893);
xnor UO_393 (O_393,N_14789,N_14858);
nor UO_394 (O_394,N_14761,N_14983);
nor UO_395 (O_395,N_14964,N_14867);
nand UO_396 (O_396,N_14818,N_14824);
and UO_397 (O_397,N_14777,N_14865);
nor UO_398 (O_398,N_14920,N_14818);
or UO_399 (O_399,N_14769,N_14994);
or UO_400 (O_400,N_14943,N_14896);
nor UO_401 (O_401,N_14979,N_14921);
nor UO_402 (O_402,N_14827,N_14956);
nand UO_403 (O_403,N_14807,N_14783);
nor UO_404 (O_404,N_14966,N_14874);
nor UO_405 (O_405,N_14974,N_14948);
and UO_406 (O_406,N_14792,N_14960);
nor UO_407 (O_407,N_14944,N_14840);
nand UO_408 (O_408,N_14776,N_14949);
or UO_409 (O_409,N_14974,N_14874);
nand UO_410 (O_410,N_14996,N_14924);
nor UO_411 (O_411,N_14814,N_14991);
nand UO_412 (O_412,N_14805,N_14869);
or UO_413 (O_413,N_14948,N_14960);
nand UO_414 (O_414,N_14990,N_14830);
xor UO_415 (O_415,N_14789,N_14927);
nor UO_416 (O_416,N_14801,N_14982);
and UO_417 (O_417,N_14968,N_14805);
or UO_418 (O_418,N_14872,N_14865);
or UO_419 (O_419,N_14860,N_14952);
and UO_420 (O_420,N_14934,N_14966);
and UO_421 (O_421,N_14959,N_14928);
nor UO_422 (O_422,N_14776,N_14833);
or UO_423 (O_423,N_14909,N_14882);
or UO_424 (O_424,N_14825,N_14932);
nor UO_425 (O_425,N_14974,N_14937);
or UO_426 (O_426,N_14800,N_14828);
or UO_427 (O_427,N_14982,N_14802);
or UO_428 (O_428,N_14938,N_14902);
xnor UO_429 (O_429,N_14972,N_14918);
xor UO_430 (O_430,N_14766,N_14785);
nor UO_431 (O_431,N_14843,N_14929);
nand UO_432 (O_432,N_14998,N_14774);
nand UO_433 (O_433,N_14871,N_14774);
or UO_434 (O_434,N_14842,N_14949);
or UO_435 (O_435,N_14891,N_14994);
or UO_436 (O_436,N_14945,N_14973);
xor UO_437 (O_437,N_14982,N_14973);
xnor UO_438 (O_438,N_14763,N_14792);
and UO_439 (O_439,N_14978,N_14836);
nand UO_440 (O_440,N_14893,N_14835);
nor UO_441 (O_441,N_14782,N_14785);
xor UO_442 (O_442,N_14937,N_14931);
xor UO_443 (O_443,N_14897,N_14791);
or UO_444 (O_444,N_14853,N_14817);
nand UO_445 (O_445,N_14998,N_14786);
xor UO_446 (O_446,N_14823,N_14758);
xor UO_447 (O_447,N_14925,N_14843);
and UO_448 (O_448,N_14970,N_14981);
xnor UO_449 (O_449,N_14882,N_14783);
nand UO_450 (O_450,N_14901,N_14834);
nor UO_451 (O_451,N_14928,N_14985);
or UO_452 (O_452,N_14750,N_14985);
nor UO_453 (O_453,N_14831,N_14931);
and UO_454 (O_454,N_14843,N_14766);
and UO_455 (O_455,N_14903,N_14869);
nand UO_456 (O_456,N_14879,N_14838);
xnor UO_457 (O_457,N_14984,N_14983);
or UO_458 (O_458,N_14821,N_14984);
xor UO_459 (O_459,N_14777,N_14825);
nand UO_460 (O_460,N_14973,N_14805);
and UO_461 (O_461,N_14974,N_14959);
nor UO_462 (O_462,N_14915,N_14769);
nor UO_463 (O_463,N_14958,N_14992);
nor UO_464 (O_464,N_14807,N_14780);
or UO_465 (O_465,N_14994,N_14813);
nand UO_466 (O_466,N_14831,N_14837);
nor UO_467 (O_467,N_14783,N_14963);
xnor UO_468 (O_468,N_14973,N_14755);
and UO_469 (O_469,N_14957,N_14880);
nand UO_470 (O_470,N_14914,N_14874);
nor UO_471 (O_471,N_14826,N_14906);
xnor UO_472 (O_472,N_14872,N_14755);
nand UO_473 (O_473,N_14844,N_14755);
xnor UO_474 (O_474,N_14879,N_14800);
xor UO_475 (O_475,N_14769,N_14972);
and UO_476 (O_476,N_14829,N_14960);
xnor UO_477 (O_477,N_14832,N_14783);
and UO_478 (O_478,N_14807,N_14828);
xor UO_479 (O_479,N_14854,N_14979);
nand UO_480 (O_480,N_14830,N_14750);
xnor UO_481 (O_481,N_14909,N_14980);
and UO_482 (O_482,N_14819,N_14829);
nand UO_483 (O_483,N_14841,N_14864);
or UO_484 (O_484,N_14869,N_14752);
or UO_485 (O_485,N_14760,N_14827);
xor UO_486 (O_486,N_14880,N_14780);
and UO_487 (O_487,N_14843,N_14894);
and UO_488 (O_488,N_14958,N_14820);
nand UO_489 (O_489,N_14836,N_14970);
and UO_490 (O_490,N_14973,N_14861);
xnor UO_491 (O_491,N_14890,N_14897);
and UO_492 (O_492,N_14909,N_14859);
or UO_493 (O_493,N_14852,N_14948);
xnor UO_494 (O_494,N_14865,N_14797);
xnor UO_495 (O_495,N_14787,N_14883);
xnor UO_496 (O_496,N_14927,N_14767);
and UO_497 (O_497,N_14861,N_14924);
nor UO_498 (O_498,N_14773,N_14926);
nand UO_499 (O_499,N_14802,N_14825);
or UO_500 (O_500,N_14761,N_14810);
nand UO_501 (O_501,N_14800,N_14958);
nor UO_502 (O_502,N_14915,N_14838);
xor UO_503 (O_503,N_14983,N_14947);
xnor UO_504 (O_504,N_14849,N_14924);
and UO_505 (O_505,N_14992,N_14972);
and UO_506 (O_506,N_14798,N_14882);
and UO_507 (O_507,N_14955,N_14957);
or UO_508 (O_508,N_14905,N_14787);
xnor UO_509 (O_509,N_14759,N_14924);
or UO_510 (O_510,N_14953,N_14834);
xor UO_511 (O_511,N_14805,N_14858);
or UO_512 (O_512,N_14983,N_14867);
and UO_513 (O_513,N_14788,N_14917);
nor UO_514 (O_514,N_14891,N_14852);
or UO_515 (O_515,N_14970,N_14818);
xor UO_516 (O_516,N_14940,N_14935);
nor UO_517 (O_517,N_14765,N_14846);
or UO_518 (O_518,N_14765,N_14774);
nor UO_519 (O_519,N_14815,N_14838);
or UO_520 (O_520,N_14917,N_14768);
nor UO_521 (O_521,N_14984,N_14805);
and UO_522 (O_522,N_14945,N_14919);
nand UO_523 (O_523,N_14793,N_14972);
and UO_524 (O_524,N_14789,N_14827);
or UO_525 (O_525,N_14794,N_14875);
and UO_526 (O_526,N_14919,N_14853);
nor UO_527 (O_527,N_14914,N_14760);
and UO_528 (O_528,N_14768,N_14758);
xor UO_529 (O_529,N_14944,N_14996);
nand UO_530 (O_530,N_14993,N_14936);
nand UO_531 (O_531,N_14995,N_14861);
xnor UO_532 (O_532,N_14852,N_14821);
or UO_533 (O_533,N_14983,N_14786);
xor UO_534 (O_534,N_14824,N_14894);
and UO_535 (O_535,N_14795,N_14977);
nor UO_536 (O_536,N_14755,N_14796);
nand UO_537 (O_537,N_14765,N_14992);
or UO_538 (O_538,N_14761,N_14819);
nor UO_539 (O_539,N_14816,N_14853);
and UO_540 (O_540,N_14902,N_14955);
or UO_541 (O_541,N_14790,N_14776);
and UO_542 (O_542,N_14856,N_14789);
nor UO_543 (O_543,N_14940,N_14830);
xnor UO_544 (O_544,N_14855,N_14813);
or UO_545 (O_545,N_14934,N_14833);
nor UO_546 (O_546,N_14847,N_14973);
xnor UO_547 (O_547,N_14852,N_14901);
xnor UO_548 (O_548,N_14990,N_14887);
and UO_549 (O_549,N_14805,N_14773);
and UO_550 (O_550,N_14985,N_14993);
and UO_551 (O_551,N_14976,N_14936);
nor UO_552 (O_552,N_14974,N_14780);
nor UO_553 (O_553,N_14768,N_14835);
nand UO_554 (O_554,N_14864,N_14895);
or UO_555 (O_555,N_14951,N_14755);
and UO_556 (O_556,N_14769,N_14876);
and UO_557 (O_557,N_14919,N_14808);
nand UO_558 (O_558,N_14841,N_14928);
and UO_559 (O_559,N_14916,N_14759);
xor UO_560 (O_560,N_14847,N_14768);
and UO_561 (O_561,N_14756,N_14997);
and UO_562 (O_562,N_14896,N_14855);
or UO_563 (O_563,N_14815,N_14842);
nand UO_564 (O_564,N_14894,N_14772);
or UO_565 (O_565,N_14908,N_14918);
and UO_566 (O_566,N_14987,N_14929);
and UO_567 (O_567,N_14808,N_14784);
and UO_568 (O_568,N_14936,N_14751);
or UO_569 (O_569,N_14863,N_14913);
and UO_570 (O_570,N_14813,N_14915);
and UO_571 (O_571,N_14987,N_14778);
nor UO_572 (O_572,N_14916,N_14905);
nand UO_573 (O_573,N_14994,N_14997);
nand UO_574 (O_574,N_14896,N_14801);
or UO_575 (O_575,N_14753,N_14851);
nor UO_576 (O_576,N_14863,N_14897);
and UO_577 (O_577,N_14938,N_14927);
and UO_578 (O_578,N_14822,N_14947);
and UO_579 (O_579,N_14756,N_14837);
xnor UO_580 (O_580,N_14757,N_14853);
xnor UO_581 (O_581,N_14913,N_14786);
nand UO_582 (O_582,N_14810,N_14991);
or UO_583 (O_583,N_14758,N_14836);
xnor UO_584 (O_584,N_14763,N_14851);
or UO_585 (O_585,N_14765,N_14917);
xor UO_586 (O_586,N_14981,N_14924);
or UO_587 (O_587,N_14956,N_14773);
xnor UO_588 (O_588,N_14877,N_14931);
nor UO_589 (O_589,N_14765,N_14916);
xor UO_590 (O_590,N_14771,N_14951);
nor UO_591 (O_591,N_14878,N_14796);
xor UO_592 (O_592,N_14799,N_14752);
xnor UO_593 (O_593,N_14984,N_14929);
xor UO_594 (O_594,N_14992,N_14919);
or UO_595 (O_595,N_14845,N_14960);
and UO_596 (O_596,N_14965,N_14843);
xnor UO_597 (O_597,N_14780,N_14845);
nand UO_598 (O_598,N_14983,N_14814);
and UO_599 (O_599,N_14858,N_14891);
nor UO_600 (O_600,N_14847,N_14858);
and UO_601 (O_601,N_14910,N_14977);
xnor UO_602 (O_602,N_14752,N_14936);
or UO_603 (O_603,N_14910,N_14788);
nor UO_604 (O_604,N_14801,N_14772);
or UO_605 (O_605,N_14856,N_14998);
nand UO_606 (O_606,N_14757,N_14968);
and UO_607 (O_607,N_14985,N_14827);
xor UO_608 (O_608,N_14795,N_14991);
and UO_609 (O_609,N_14795,N_14888);
or UO_610 (O_610,N_14770,N_14814);
and UO_611 (O_611,N_14840,N_14923);
and UO_612 (O_612,N_14879,N_14878);
xor UO_613 (O_613,N_14827,N_14919);
or UO_614 (O_614,N_14930,N_14753);
or UO_615 (O_615,N_14803,N_14913);
xnor UO_616 (O_616,N_14791,N_14867);
nor UO_617 (O_617,N_14806,N_14792);
and UO_618 (O_618,N_14955,N_14752);
nor UO_619 (O_619,N_14828,N_14979);
nor UO_620 (O_620,N_14842,N_14824);
nor UO_621 (O_621,N_14998,N_14941);
and UO_622 (O_622,N_14905,N_14789);
nor UO_623 (O_623,N_14951,N_14839);
and UO_624 (O_624,N_14901,N_14758);
nand UO_625 (O_625,N_14875,N_14813);
nand UO_626 (O_626,N_14871,N_14938);
and UO_627 (O_627,N_14779,N_14985);
and UO_628 (O_628,N_14876,N_14778);
nand UO_629 (O_629,N_14852,N_14797);
nor UO_630 (O_630,N_14931,N_14949);
or UO_631 (O_631,N_14866,N_14904);
xnor UO_632 (O_632,N_14910,N_14986);
and UO_633 (O_633,N_14803,N_14766);
nor UO_634 (O_634,N_14960,N_14828);
and UO_635 (O_635,N_14854,N_14925);
and UO_636 (O_636,N_14949,N_14823);
xnor UO_637 (O_637,N_14848,N_14959);
nand UO_638 (O_638,N_14782,N_14905);
nor UO_639 (O_639,N_14894,N_14878);
and UO_640 (O_640,N_14828,N_14798);
and UO_641 (O_641,N_14973,N_14817);
nor UO_642 (O_642,N_14774,N_14983);
and UO_643 (O_643,N_14981,N_14861);
or UO_644 (O_644,N_14889,N_14927);
xnor UO_645 (O_645,N_14827,N_14953);
or UO_646 (O_646,N_14799,N_14988);
nor UO_647 (O_647,N_14935,N_14924);
or UO_648 (O_648,N_14930,N_14945);
or UO_649 (O_649,N_14994,N_14971);
xnor UO_650 (O_650,N_14807,N_14785);
nor UO_651 (O_651,N_14829,N_14994);
xnor UO_652 (O_652,N_14841,N_14791);
xor UO_653 (O_653,N_14825,N_14879);
nor UO_654 (O_654,N_14861,N_14909);
xnor UO_655 (O_655,N_14918,N_14924);
or UO_656 (O_656,N_14954,N_14822);
xnor UO_657 (O_657,N_14963,N_14753);
and UO_658 (O_658,N_14779,N_14805);
xnor UO_659 (O_659,N_14976,N_14811);
xnor UO_660 (O_660,N_14785,N_14931);
and UO_661 (O_661,N_14773,N_14890);
nand UO_662 (O_662,N_14993,N_14945);
and UO_663 (O_663,N_14928,N_14866);
and UO_664 (O_664,N_14844,N_14947);
xor UO_665 (O_665,N_14936,N_14792);
and UO_666 (O_666,N_14971,N_14752);
nand UO_667 (O_667,N_14933,N_14824);
and UO_668 (O_668,N_14966,N_14951);
or UO_669 (O_669,N_14899,N_14955);
nand UO_670 (O_670,N_14962,N_14879);
nor UO_671 (O_671,N_14969,N_14802);
or UO_672 (O_672,N_14787,N_14941);
and UO_673 (O_673,N_14751,N_14825);
or UO_674 (O_674,N_14966,N_14827);
nor UO_675 (O_675,N_14984,N_14760);
or UO_676 (O_676,N_14771,N_14873);
nand UO_677 (O_677,N_14763,N_14879);
and UO_678 (O_678,N_14898,N_14883);
nand UO_679 (O_679,N_14983,N_14936);
and UO_680 (O_680,N_14896,N_14849);
nor UO_681 (O_681,N_14991,N_14897);
and UO_682 (O_682,N_14806,N_14835);
or UO_683 (O_683,N_14829,N_14781);
nand UO_684 (O_684,N_14809,N_14872);
nand UO_685 (O_685,N_14966,N_14981);
xnor UO_686 (O_686,N_14957,N_14923);
nor UO_687 (O_687,N_14894,N_14898);
nor UO_688 (O_688,N_14757,N_14795);
nor UO_689 (O_689,N_14861,N_14897);
nand UO_690 (O_690,N_14822,N_14878);
or UO_691 (O_691,N_14835,N_14929);
xor UO_692 (O_692,N_14775,N_14793);
nor UO_693 (O_693,N_14793,N_14958);
nor UO_694 (O_694,N_14797,N_14943);
xnor UO_695 (O_695,N_14777,N_14966);
or UO_696 (O_696,N_14845,N_14900);
or UO_697 (O_697,N_14793,N_14935);
or UO_698 (O_698,N_14903,N_14913);
xnor UO_699 (O_699,N_14807,N_14879);
nand UO_700 (O_700,N_14999,N_14881);
and UO_701 (O_701,N_14858,N_14996);
and UO_702 (O_702,N_14984,N_14880);
nand UO_703 (O_703,N_14890,N_14916);
nor UO_704 (O_704,N_14931,N_14838);
or UO_705 (O_705,N_14857,N_14796);
nor UO_706 (O_706,N_14859,N_14753);
xor UO_707 (O_707,N_14862,N_14987);
and UO_708 (O_708,N_14865,N_14931);
nand UO_709 (O_709,N_14912,N_14870);
nand UO_710 (O_710,N_14877,N_14983);
and UO_711 (O_711,N_14759,N_14963);
xor UO_712 (O_712,N_14839,N_14972);
xnor UO_713 (O_713,N_14949,N_14764);
nor UO_714 (O_714,N_14859,N_14823);
and UO_715 (O_715,N_14830,N_14871);
xor UO_716 (O_716,N_14996,N_14751);
or UO_717 (O_717,N_14785,N_14872);
and UO_718 (O_718,N_14836,N_14896);
xnor UO_719 (O_719,N_14943,N_14967);
and UO_720 (O_720,N_14816,N_14859);
xnor UO_721 (O_721,N_14982,N_14978);
nand UO_722 (O_722,N_14844,N_14964);
xnor UO_723 (O_723,N_14900,N_14762);
nor UO_724 (O_724,N_14911,N_14986);
nand UO_725 (O_725,N_14815,N_14983);
or UO_726 (O_726,N_14870,N_14975);
nand UO_727 (O_727,N_14814,N_14977);
or UO_728 (O_728,N_14956,N_14886);
or UO_729 (O_729,N_14881,N_14914);
nor UO_730 (O_730,N_14775,N_14911);
or UO_731 (O_731,N_14961,N_14807);
or UO_732 (O_732,N_14881,N_14861);
xor UO_733 (O_733,N_14831,N_14883);
nand UO_734 (O_734,N_14861,N_14969);
and UO_735 (O_735,N_14905,N_14780);
and UO_736 (O_736,N_14772,N_14930);
and UO_737 (O_737,N_14914,N_14958);
or UO_738 (O_738,N_14924,N_14887);
and UO_739 (O_739,N_14971,N_14824);
xnor UO_740 (O_740,N_14973,N_14803);
xor UO_741 (O_741,N_14883,N_14980);
or UO_742 (O_742,N_14754,N_14949);
or UO_743 (O_743,N_14949,N_14773);
or UO_744 (O_744,N_14979,N_14888);
and UO_745 (O_745,N_14886,N_14933);
nor UO_746 (O_746,N_14755,N_14789);
or UO_747 (O_747,N_14836,N_14994);
xor UO_748 (O_748,N_14934,N_14798);
xnor UO_749 (O_749,N_14895,N_14992);
and UO_750 (O_750,N_14771,N_14818);
xor UO_751 (O_751,N_14902,N_14953);
xor UO_752 (O_752,N_14866,N_14789);
nand UO_753 (O_753,N_14791,N_14751);
nor UO_754 (O_754,N_14862,N_14776);
or UO_755 (O_755,N_14883,N_14760);
nand UO_756 (O_756,N_14952,N_14766);
nand UO_757 (O_757,N_14796,N_14959);
and UO_758 (O_758,N_14775,N_14947);
and UO_759 (O_759,N_14887,N_14991);
or UO_760 (O_760,N_14777,N_14839);
xor UO_761 (O_761,N_14983,N_14978);
nand UO_762 (O_762,N_14800,N_14977);
xor UO_763 (O_763,N_14917,N_14928);
nand UO_764 (O_764,N_14959,N_14898);
nand UO_765 (O_765,N_14753,N_14957);
and UO_766 (O_766,N_14938,N_14841);
nand UO_767 (O_767,N_14858,N_14767);
nand UO_768 (O_768,N_14834,N_14988);
or UO_769 (O_769,N_14973,N_14884);
nor UO_770 (O_770,N_14807,N_14837);
nor UO_771 (O_771,N_14834,N_14844);
xnor UO_772 (O_772,N_14813,N_14949);
or UO_773 (O_773,N_14885,N_14844);
or UO_774 (O_774,N_14955,N_14870);
nand UO_775 (O_775,N_14940,N_14819);
xnor UO_776 (O_776,N_14802,N_14936);
nand UO_777 (O_777,N_14930,N_14973);
xor UO_778 (O_778,N_14951,N_14924);
or UO_779 (O_779,N_14926,N_14895);
and UO_780 (O_780,N_14910,N_14770);
xnor UO_781 (O_781,N_14988,N_14977);
nand UO_782 (O_782,N_14895,N_14776);
nand UO_783 (O_783,N_14804,N_14899);
xor UO_784 (O_784,N_14950,N_14889);
xnor UO_785 (O_785,N_14786,N_14961);
xnor UO_786 (O_786,N_14754,N_14888);
nor UO_787 (O_787,N_14938,N_14758);
and UO_788 (O_788,N_14928,N_14999);
or UO_789 (O_789,N_14814,N_14889);
nand UO_790 (O_790,N_14999,N_14812);
nor UO_791 (O_791,N_14962,N_14890);
nand UO_792 (O_792,N_14792,N_14757);
xor UO_793 (O_793,N_14965,N_14931);
and UO_794 (O_794,N_14929,N_14808);
xnor UO_795 (O_795,N_14781,N_14995);
nor UO_796 (O_796,N_14861,N_14872);
or UO_797 (O_797,N_14891,N_14790);
nor UO_798 (O_798,N_14876,N_14817);
nand UO_799 (O_799,N_14814,N_14868);
nor UO_800 (O_800,N_14958,N_14853);
xnor UO_801 (O_801,N_14861,N_14826);
nand UO_802 (O_802,N_14965,N_14954);
nand UO_803 (O_803,N_14829,N_14912);
or UO_804 (O_804,N_14914,N_14888);
nor UO_805 (O_805,N_14778,N_14995);
xnor UO_806 (O_806,N_14922,N_14770);
xor UO_807 (O_807,N_14902,N_14900);
xnor UO_808 (O_808,N_14995,N_14775);
and UO_809 (O_809,N_14949,N_14886);
nand UO_810 (O_810,N_14868,N_14927);
or UO_811 (O_811,N_14949,N_14888);
or UO_812 (O_812,N_14787,N_14875);
nand UO_813 (O_813,N_14968,N_14981);
xnor UO_814 (O_814,N_14786,N_14914);
or UO_815 (O_815,N_14864,N_14752);
nand UO_816 (O_816,N_14978,N_14906);
or UO_817 (O_817,N_14895,N_14876);
and UO_818 (O_818,N_14768,N_14783);
nor UO_819 (O_819,N_14953,N_14900);
nor UO_820 (O_820,N_14841,N_14817);
nand UO_821 (O_821,N_14984,N_14751);
and UO_822 (O_822,N_14850,N_14799);
or UO_823 (O_823,N_14960,N_14876);
and UO_824 (O_824,N_14988,N_14950);
or UO_825 (O_825,N_14938,N_14799);
nand UO_826 (O_826,N_14770,N_14789);
or UO_827 (O_827,N_14782,N_14796);
or UO_828 (O_828,N_14845,N_14874);
xor UO_829 (O_829,N_14785,N_14839);
xnor UO_830 (O_830,N_14847,N_14765);
xnor UO_831 (O_831,N_14923,N_14888);
xor UO_832 (O_832,N_14980,N_14804);
nand UO_833 (O_833,N_14865,N_14824);
or UO_834 (O_834,N_14803,N_14886);
nor UO_835 (O_835,N_14977,N_14773);
and UO_836 (O_836,N_14985,N_14988);
xor UO_837 (O_837,N_14791,N_14962);
xor UO_838 (O_838,N_14756,N_14892);
or UO_839 (O_839,N_14872,N_14909);
and UO_840 (O_840,N_14963,N_14972);
nand UO_841 (O_841,N_14862,N_14956);
nand UO_842 (O_842,N_14996,N_14915);
nand UO_843 (O_843,N_14904,N_14819);
and UO_844 (O_844,N_14754,N_14789);
or UO_845 (O_845,N_14967,N_14938);
or UO_846 (O_846,N_14863,N_14990);
nand UO_847 (O_847,N_14980,N_14836);
or UO_848 (O_848,N_14871,N_14929);
or UO_849 (O_849,N_14930,N_14853);
nor UO_850 (O_850,N_14841,N_14924);
xor UO_851 (O_851,N_14755,N_14813);
xnor UO_852 (O_852,N_14972,N_14854);
and UO_853 (O_853,N_14869,N_14818);
or UO_854 (O_854,N_14990,N_14852);
xnor UO_855 (O_855,N_14866,N_14775);
or UO_856 (O_856,N_14784,N_14796);
nor UO_857 (O_857,N_14872,N_14784);
nor UO_858 (O_858,N_14922,N_14866);
nor UO_859 (O_859,N_14797,N_14949);
or UO_860 (O_860,N_14850,N_14867);
nand UO_861 (O_861,N_14924,N_14820);
nor UO_862 (O_862,N_14884,N_14830);
nor UO_863 (O_863,N_14827,N_14845);
nor UO_864 (O_864,N_14889,N_14907);
nand UO_865 (O_865,N_14926,N_14821);
or UO_866 (O_866,N_14815,N_14798);
xnor UO_867 (O_867,N_14764,N_14957);
and UO_868 (O_868,N_14870,N_14841);
and UO_869 (O_869,N_14785,N_14829);
or UO_870 (O_870,N_14872,N_14902);
xor UO_871 (O_871,N_14943,N_14868);
xnor UO_872 (O_872,N_14885,N_14979);
nor UO_873 (O_873,N_14816,N_14782);
xor UO_874 (O_874,N_14943,N_14922);
or UO_875 (O_875,N_14912,N_14795);
xor UO_876 (O_876,N_14769,N_14931);
nand UO_877 (O_877,N_14823,N_14888);
nor UO_878 (O_878,N_14763,N_14903);
nand UO_879 (O_879,N_14917,N_14925);
or UO_880 (O_880,N_14965,N_14940);
nor UO_881 (O_881,N_14857,N_14772);
xnor UO_882 (O_882,N_14849,N_14916);
and UO_883 (O_883,N_14964,N_14848);
or UO_884 (O_884,N_14971,N_14861);
xor UO_885 (O_885,N_14975,N_14863);
or UO_886 (O_886,N_14908,N_14958);
xor UO_887 (O_887,N_14978,N_14904);
and UO_888 (O_888,N_14976,N_14872);
nor UO_889 (O_889,N_14801,N_14864);
xor UO_890 (O_890,N_14841,N_14986);
nor UO_891 (O_891,N_14897,N_14821);
nor UO_892 (O_892,N_14773,N_14879);
and UO_893 (O_893,N_14800,N_14806);
and UO_894 (O_894,N_14957,N_14886);
xor UO_895 (O_895,N_14874,N_14973);
and UO_896 (O_896,N_14879,N_14954);
nor UO_897 (O_897,N_14889,N_14798);
nand UO_898 (O_898,N_14835,N_14990);
nand UO_899 (O_899,N_14821,N_14825);
xor UO_900 (O_900,N_14831,N_14840);
or UO_901 (O_901,N_14842,N_14790);
xnor UO_902 (O_902,N_14808,N_14764);
and UO_903 (O_903,N_14841,N_14845);
nand UO_904 (O_904,N_14890,N_14925);
xor UO_905 (O_905,N_14989,N_14803);
nor UO_906 (O_906,N_14867,N_14777);
nor UO_907 (O_907,N_14759,N_14905);
and UO_908 (O_908,N_14807,N_14937);
and UO_909 (O_909,N_14855,N_14967);
and UO_910 (O_910,N_14943,N_14826);
and UO_911 (O_911,N_14938,N_14879);
or UO_912 (O_912,N_14863,N_14850);
xnor UO_913 (O_913,N_14944,N_14779);
xnor UO_914 (O_914,N_14887,N_14983);
nor UO_915 (O_915,N_14845,N_14884);
nand UO_916 (O_916,N_14857,N_14897);
nand UO_917 (O_917,N_14791,N_14939);
and UO_918 (O_918,N_14866,N_14819);
or UO_919 (O_919,N_14879,N_14897);
or UO_920 (O_920,N_14970,N_14929);
nand UO_921 (O_921,N_14913,N_14988);
nor UO_922 (O_922,N_14890,N_14939);
nand UO_923 (O_923,N_14769,N_14951);
and UO_924 (O_924,N_14915,N_14976);
and UO_925 (O_925,N_14915,N_14750);
and UO_926 (O_926,N_14817,N_14821);
and UO_927 (O_927,N_14772,N_14891);
and UO_928 (O_928,N_14801,N_14930);
nand UO_929 (O_929,N_14902,N_14903);
nor UO_930 (O_930,N_14795,N_14918);
xnor UO_931 (O_931,N_14770,N_14751);
nor UO_932 (O_932,N_14874,N_14829);
nand UO_933 (O_933,N_14766,N_14764);
nor UO_934 (O_934,N_14788,N_14983);
xor UO_935 (O_935,N_14787,N_14928);
nor UO_936 (O_936,N_14938,N_14955);
xor UO_937 (O_937,N_14860,N_14779);
or UO_938 (O_938,N_14818,N_14828);
nor UO_939 (O_939,N_14986,N_14800);
nor UO_940 (O_940,N_14969,N_14964);
and UO_941 (O_941,N_14912,N_14785);
nand UO_942 (O_942,N_14773,N_14893);
and UO_943 (O_943,N_14797,N_14904);
and UO_944 (O_944,N_14835,N_14824);
nor UO_945 (O_945,N_14855,N_14914);
nor UO_946 (O_946,N_14819,N_14864);
or UO_947 (O_947,N_14947,N_14919);
xnor UO_948 (O_948,N_14900,N_14989);
nor UO_949 (O_949,N_14884,N_14888);
nand UO_950 (O_950,N_14836,N_14812);
nand UO_951 (O_951,N_14862,N_14996);
or UO_952 (O_952,N_14786,N_14811);
xnor UO_953 (O_953,N_14765,N_14870);
xnor UO_954 (O_954,N_14852,N_14757);
or UO_955 (O_955,N_14997,N_14882);
and UO_956 (O_956,N_14962,N_14923);
nand UO_957 (O_957,N_14818,N_14838);
nor UO_958 (O_958,N_14784,N_14858);
and UO_959 (O_959,N_14901,N_14851);
nand UO_960 (O_960,N_14999,N_14807);
nor UO_961 (O_961,N_14920,N_14940);
xor UO_962 (O_962,N_14771,N_14875);
xnor UO_963 (O_963,N_14860,N_14907);
or UO_964 (O_964,N_14786,N_14975);
xor UO_965 (O_965,N_14812,N_14970);
or UO_966 (O_966,N_14855,N_14954);
and UO_967 (O_967,N_14825,N_14992);
and UO_968 (O_968,N_14910,N_14890);
and UO_969 (O_969,N_14825,N_14904);
xnor UO_970 (O_970,N_14911,N_14974);
or UO_971 (O_971,N_14894,N_14820);
xor UO_972 (O_972,N_14986,N_14812);
or UO_973 (O_973,N_14765,N_14789);
nand UO_974 (O_974,N_14818,N_14832);
nand UO_975 (O_975,N_14944,N_14995);
nor UO_976 (O_976,N_14905,N_14876);
nor UO_977 (O_977,N_14908,N_14882);
nor UO_978 (O_978,N_14783,N_14811);
or UO_979 (O_979,N_14944,N_14824);
nor UO_980 (O_980,N_14788,N_14947);
nor UO_981 (O_981,N_14946,N_14772);
nand UO_982 (O_982,N_14943,N_14931);
or UO_983 (O_983,N_14812,N_14822);
nor UO_984 (O_984,N_14812,N_14808);
nor UO_985 (O_985,N_14953,N_14830);
nor UO_986 (O_986,N_14768,N_14819);
nand UO_987 (O_987,N_14797,N_14911);
and UO_988 (O_988,N_14937,N_14777);
or UO_989 (O_989,N_14872,N_14988);
or UO_990 (O_990,N_14952,N_14935);
xor UO_991 (O_991,N_14762,N_14956);
nor UO_992 (O_992,N_14829,N_14833);
and UO_993 (O_993,N_14987,N_14802);
nand UO_994 (O_994,N_14982,N_14795);
nand UO_995 (O_995,N_14966,N_14819);
or UO_996 (O_996,N_14904,N_14947);
or UO_997 (O_997,N_14913,N_14909);
or UO_998 (O_998,N_14776,N_14782);
or UO_999 (O_999,N_14985,N_14778);
xor UO_1000 (O_1000,N_14774,N_14968);
and UO_1001 (O_1001,N_14797,N_14750);
and UO_1002 (O_1002,N_14750,N_14860);
and UO_1003 (O_1003,N_14765,N_14806);
or UO_1004 (O_1004,N_14911,N_14922);
nand UO_1005 (O_1005,N_14815,N_14986);
nor UO_1006 (O_1006,N_14752,N_14905);
and UO_1007 (O_1007,N_14831,N_14972);
or UO_1008 (O_1008,N_14779,N_14901);
xnor UO_1009 (O_1009,N_14985,N_14826);
and UO_1010 (O_1010,N_14841,N_14754);
nand UO_1011 (O_1011,N_14927,N_14764);
nand UO_1012 (O_1012,N_14786,N_14873);
or UO_1013 (O_1013,N_14975,N_14850);
or UO_1014 (O_1014,N_14902,N_14985);
nor UO_1015 (O_1015,N_14966,N_14954);
nand UO_1016 (O_1016,N_14784,N_14859);
xnor UO_1017 (O_1017,N_14961,N_14881);
nor UO_1018 (O_1018,N_14993,N_14962);
nor UO_1019 (O_1019,N_14757,N_14856);
nand UO_1020 (O_1020,N_14995,N_14914);
xor UO_1021 (O_1021,N_14979,N_14998);
xor UO_1022 (O_1022,N_14873,N_14931);
xnor UO_1023 (O_1023,N_14934,N_14876);
nand UO_1024 (O_1024,N_14753,N_14867);
nand UO_1025 (O_1025,N_14932,N_14945);
or UO_1026 (O_1026,N_14751,N_14824);
xor UO_1027 (O_1027,N_14966,N_14807);
nand UO_1028 (O_1028,N_14759,N_14827);
xnor UO_1029 (O_1029,N_14976,N_14944);
xnor UO_1030 (O_1030,N_14854,N_14913);
nand UO_1031 (O_1031,N_14915,N_14908);
nor UO_1032 (O_1032,N_14838,N_14969);
and UO_1033 (O_1033,N_14864,N_14887);
xor UO_1034 (O_1034,N_14807,N_14836);
nor UO_1035 (O_1035,N_14951,N_14854);
nand UO_1036 (O_1036,N_14895,N_14809);
or UO_1037 (O_1037,N_14991,N_14883);
xor UO_1038 (O_1038,N_14757,N_14985);
and UO_1039 (O_1039,N_14878,N_14916);
xnor UO_1040 (O_1040,N_14811,N_14873);
or UO_1041 (O_1041,N_14851,N_14900);
and UO_1042 (O_1042,N_14899,N_14850);
or UO_1043 (O_1043,N_14966,N_14886);
xor UO_1044 (O_1044,N_14974,N_14865);
nor UO_1045 (O_1045,N_14837,N_14812);
nand UO_1046 (O_1046,N_14855,N_14847);
nor UO_1047 (O_1047,N_14935,N_14977);
and UO_1048 (O_1048,N_14898,N_14995);
nand UO_1049 (O_1049,N_14919,N_14817);
and UO_1050 (O_1050,N_14804,N_14939);
nand UO_1051 (O_1051,N_14949,N_14908);
xnor UO_1052 (O_1052,N_14847,N_14820);
nor UO_1053 (O_1053,N_14872,N_14922);
and UO_1054 (O_1054,N_14918,N_14836);
nor UO_1055 (O_1055,N_14868,N_14896);
nor UO_1056 (O_1056,N_14946,N_14828);
xnor UO_1057 (O_1057,N_14770,N_14911);
nand UO_1058 (O_1058,N_14767,N_14884);
and UO_1059 (O_1059,N_14963,N_14939);
or UO_1060 (O_1060,N_14788,N_14807);
nand UO_1061 (O_1061,N_14784,N_14915);
or UO_1062 (O_1062,N_14873,N_14972);
and UO_1063 (O_1063,N_14828,N_14844);
and UO_1064 (O_1064,N_14991,N_14963);
or UO_1065 (O_1065,N_14763,N_14797);
xor UO_1066 (O_1066,N_14892,N_14791);
xnor UO_1067 (O_1067,N_14927,N_14796);
or UO_1068 (O_1068,N_14868,N_14968);
or UO_1069 (O_1069,N_14787,N_14767);
or UO_1070 (O_1070,N_14771,N_14791);
xor UO_1071 (O_1071,N_14794,N_14882);
xor UO_1072 (O_1072,N_14882,N_14923);
and UO_1073 (O_1073,N_14927,N_14986);
xor UO_1074 (O_1074,N_14801,N_14859);
nor UO_1075 (O_1075,N_14976,N_14829);
xnor UO_1076 (O_1076,N_14856,N_14753);
nand UO_1077 (O_1077,N_14983,N_14843);
nand UO_1078 (O_1078,N_14920,N_14876);
nand UO_1079 (O_1079,N_14834,N_14797);
nor UO_1080 (O_1080,N_14864,N_14797);
and UO_1081 (O_1081,N_14786,N_14995);
xnor UO_1082 (O_1082,N_14959,N_14816);
and UO_1083 (O_1083,N_14819,N_14952);
nor UO_1084 (O_1084,N_14970,N_14884);
or UO_1085 (O_1085,N_14864,N_14949);
xor UO_1086 (O_1086,N_14947,N_14865);
or UO_1087 (O_1087,N_14797,N_14810);
or UO_1088 (O_1088,N_14756,N_14950);
xnor UO_1089 (O_1089,N_14756,N_14916);
nor UO_1090 (O_1090,N_14797,N_14849);
and UO_1091 (O_1091,N_14799,N_14985);
nor UO_1092 (O_1092,N_14872,N_14776);
or UO_1093 (O_1093,N_14889,N_14751);
nor UO_1094 (O_1094,N_14827,N_14938);
xnor UO_1095 (O_1095,N_14977,N_14813);
nor UO_1096 (O_1096,N_14947,N_14939);
and UO_1097 (O_1097,N_14815,N_14904);
and UO_1098 (O_1098,N_14763,N_14931);
xnor UO_1099 (O_1099,N_14941,N_14922);
and UO_1100 (O_1100,N_14851,N_14798);
and UO_1101 (O_1101,N_14793,N_14888);
nor UO_1102 (O_1102,N_14856,N_14922);
and UO_1103 (O_1103,N_14765,N_14868);
and UO_1104 (O_1104,N_14775,N_14897);
or UO_1105 (O_1105,N_14930,N_14864);
or UO_1106 (O_1106,N_14840,N_14955);
nor UO_1107 (O_1107,N_14796,N_14930);
nor UO_1108 (O_1108,N_14895,N_14826);
or UO_1109 (O_1109,N_14963,N_14857);
and UO_1110 (O_1110,N_14887,N_14805);
and UO_1111 (O_1111,N_14859,N_14905);
and UO_1112 (O_1112,N_14864,N_14959);
nor UO_1113 (O_1113,N_14778,N_14817);
nand UO_1114 (O_1114,N_14991,N_14842);
nor UO_1115 (O_1115,N_14783,N_14902);
or UO_1116 (O_1116,N_14870,N_14973);
or UO_1117 (O_1117,N_14904,N_14827);
or UO_1118 (O_1118,N_14765,N_14777);
or UO_1119 (O_1119,N_14848,N_14852);
or UO_1120 (O_1120,N_14991,N_14967);
nand UO_1121 (O_1121,N_14868,N_14998);
or UO_1122 (O_1122,N_14905,N_14893);
xor UO_1123 (O_1123,N_14804,N_14999);
nand UO_1124 (O_1124,N_14869,N_14789);
nor UO_1125 (O_1125,N_14977,N_14755);
and UO_1126 (O_1126,N_14761,N_14789);
and UO_1127 (O_1127,N_14809,N_14936);
nor UO_1128 (O_1128,N_14783,N_14949);
and UO_1129 (O_1129,N_14919,N_14968);
and UO_1130 (O_1130,N_14825,N_14816);
nand UO_1131 (O_1131,N_14767,N_14950);
and UO_1132 (O_1132,N_14752,N_14862);
nor UO_1133 (O_1133,N_14915,N_14814);
or UO_1134 (O_1134,N_14879,N_14889);
xor UO_1135 (O_1135,N_14854,N_14867);
or UO_1136 (O_1136,N_14844,N_14966);
and UO_1137 (O_1137,N_14981,N_14990);
nor UO_1138 (O_1138,N_14750,N_14755);
and UO_1139 (O_1139,N_14903,N_14868);
nor UO_1140 (O_1140,N_14996,N_14953);
and UO_1141 (O_1141,N_14815,N_14945);
or UO_1142 (O_1142,N_14909,N_14792);
or UO_1143 (O_1143,N_14838,N_14984);
nand UO_1144 (O_1144,N_14871,N_14959);
or UO_1145 (O_1145,N_14905,N_14976);
nand UO_1146 (O_1146,N_14966,N_14989);
xnor UO_1147 (O_1147,N_14892,N_14770);
nand UO_1148 (O_1148,N_14822,N_14935);
or UO_1149 (O_1149,N_14882,N_14838);
or UO_1150 (O_1150,N_14757,N_14865);
nor UO_1151 (O_1151,N_14779,N_14812);
or UO_1152 (O_1152,N_14881,N_14884);
or UO_1153 (O_1153,N_14890,N_14817);
xor UO_1154 (O_1154,N_14799,N_14956);
or UO_1155 (O_1155,N_14775,N_14776);
and UO_1156 (O_1156,N_14960,N_14911);
and UO_1157 (O_1157,N_14814,N_14870);
or UO_1158 (O_1158,N_14927,N_14752);
xnor UO_1159 (O_1159,N_14855,N_14801);
nor UO_1160 (O_1160,N_14881,N_14760);
nand UO_1161 (O_1161,N_14874,N_14847);
xnor UO_1162 (O_1162,N_14928,N_14810);
or UO_1163 (O_1163,N_14829,N_14832);
nor UO_1164 (O_1164,N_14888,N_14782);
nor UO_1165 (O_1165,N_14847,N_14946);
nor UO_1166 (O_1166,N_14868,N_14961);
or UO_1167 (O_1167,N_14890,N_14850);
nand UO_1168 (O_1168,N_14819,N_14944);
or UO_1169 (O_1169,N_14994,N_14937);
or UO_1170 (O_1170,N_14770,N_14853);
nand UO_1171 (O_1171,N_14823,N_14872);
xnor UO_1172 (O_1172,N_14859,N_14824);
xnor UO_1173 (O_1173,N_14997,N_14912);
xnor UO_1174 (O_1174,N_14803,N_14819);
xnor UO_1175 (O_1175,N_14781,N_14914);
nand UO_1176 (O_1176,N_14959,N_14884);
xor UO_1177 (O_1177,N_14974,N_14989);
and UO_1178 (O_1178,N_14982,N_14853);
xnor UO_1179 (O_1179,N_14928,N_14979);
and UO_1180 (O_1180,N_14753,N_14910);
xnor UO_1181 (O_1181,N_14788,N_14887);
or UO_1182 (O_1182,N_14793,N_14963);
nand UO_1183 (O_1183,N_14773,N_14992);
nor UO_1184 (O_1184,N_14995,N_14953);
and UO_1185 (O_1185,N_14968,N_14803);
or UO_1186 (O_1186,N_14771,N_14898);
nand UO_1187 (O_1187,N_14915,N_14977);
and UO_1188 (O_1188,N_14789,N_14759);
or UO_1189 (O_1189,N_14750,N_14870);
nand UO_1190 (O_1190,N_14962,N_14988);
xor UO_1191 (O_1191,N_14763,N_14873);
or UO_1192 (O_1192,N_14897,N_14764);
or UO_1193 (O_1193,N_14985,N_14907);
nand UO_1194 (O_1194,N_14962,N_14867);
or UO_1195 (O_1195,N_14874,N_14997);
or UO_1196 (O_1196,N_14972,N_14860);
xor UO_1197 (O_1197,N_14984,N_14966);
or UO_1198 (O_1198,N_14903,N_14859);
or UO_1199 (O_1199,N_14801,N_14938);
nand UO_1200 (O_1200,N_14962,N_14937);
or UO_1201 (O_1201,N_14780,N_14828);
xnor UO_1202 (O_1202,N_14892,N_14990);
and UO_1203 (O_1203,N_14978,N_14973);
and UO_1204 (O_1204,N_14895,N_14849);
xnor UO_1205 (O_1205,N_14972,N_14978);
nand UO_1206 (O_1206,N_14995,N_14759);
nand UO_1207 (O_1207,N_14783,N_14803);
and UO_1208 (O_1208,N_14891,N_14818);
or UO_1209 (O_1209,N_14837,N_14966);
xor UO_1210 (O_1210,N_14979,N_14768);
and UO_1211 (O_1211,N_14787,N_14978);
or UO_1212 (O_1212,N_14837,N_14851);
and UO_1213 (O_1213,N_14898,N_14779);
and UO_1214 (O_1214,N_14900,N_14973);
nor UO_1215 (O_1215,N_14902,N_14766);
nand UO_1216 (O_1216,N_14860,N_14862);
and UO_1217 (O_1217,N_14929,N_14972);
and UO_1218 (O_1218,N_14949,N_14847);
nor UO_1219 (O_1219,N_14858,N_14882);
nand UO_1220 (O_1220,N_14777,N_14941);
nand UO_1221 (O_1221,N_14905,N_14781);
or UO_1222 (O_1222,N_14992,N_14807);
nand UO_1223 (O_1223,N_14990,N_14857);
or UO_1224 (O_1224,N_14975,N_14892);
xor UO_1225 (O_1225,N_14941,N_14846);
nor UO_1226 (O_1226,N_14847,N_14975);
and UO_1227 (O_1227,N_14798,N_14831);
nor UO_1228 (O_1228,N_14900,N_14946);
or UO_1229 (O_1229,N_14832,N_14795);
nand UO_1230 (O_1230,N_14805,N_14988);
and UO_1231 (O_1231,N_14973,N_14966);
xor UO_1232 (O_1232,N_14836,N_14789);
and UO_1233 (O_1233,N_14810,N_14804);
or UO_1234 (O_1234,N_14782,N_14820);
nand UO_1235 (O_1235,N_14839,N_14755);
xor UO_1236 (O_1236,N_14845,N_14812);
xor UO_1237 (O_1237,N_14950,N_14991);
and UO_1238 (O_1238,N_14886,N_14922);
xnor UO_1239 (O_1239,N_14877,N_14757);
nor UO_1240 (O_1240,N_14913,N_14911);
or UO_1241 (O_1241,N_14885,N_14904);
and UO_1242 (O_1242,N_14808,N_14767);
xnor UO_1243 (O_1243,N_14866,N_14882);
nand UO_1244 (O_1244,N_14830,N_14753);
nand UO_1245 (O_1245,N_14857,N_14952);
and UO_1246 (O_1246,N_14752,N_14774);
or UO_1247 (O_1247,N_14948,N_14897);
and UO_1248 (O_1248,N_14895,N_14799);
nand UO_1249 (O_1249,N_14958,N_14973);
nand UO_1250 (O_1250,N_14991,N_14945);
nand UO_1251 (O_1251,N_14932,N_14766);
xor UO_1252 (O_1252,N_14877,N_14978);
or UO_1253 (O_1253,N_14898,N_14999);
and UO_1254 (O_1254,N_14915,N_14911);
xor UO_1255 (O_1255,N_14951,N_14829);
xnor UO_1256 (O_1256,N_14885,N_14853);
xnor UO_1257 (O_1257,N_14835,N_14980);
nand UO_1258 (O_1258,N_14787,N_14755);
xnor UO_1259 (O_1259,N_14928,N_14902);
xnor UO_1260 (O_1260,N_14799,N_14928);
or UO_1261 (O_1261,N_14919,N_14986);
or UO_1262 (O_1262,N_14976,N_14925);
nor UO_1263 (O_1263,N_14821,N_14905);
xnor UO_1264 (O_1264,N_14861,N_14989);
nand UO_1265 (O_1265,N_14999,N_14843);
or UO_1266 (O_1266,N_14776,N_14886);
nand UO_1267 (O_1267,N_14926,N_14838);
nor UO_1268 (O_1268,N_14979,N_14997);
and UO_1269 (O_1269,N_14815,N_14984);
nor UO_1270 (O_1270,N_14832,N_14943);
or UO_1271 (O_1271,N_14835,N_14951);
and UO_1272 (O_1272,N_14852,N_14759);
xnor UO_1273 (O_1273,N_14865,N_14909);
and UO_1274 (O_1274,N_14981,N_14805);
nand UO_1275 (O_1275,N_14900,N_14925);
nand UO_1276 (O_1276,N_14884,N_14803);
nand UO_1277 (O_1277,N_14958,N_14923);
and UO_1278 (O_1278,N_14753,N_14925);
nor UO_1279 (O_1279,N_14846,N_14950);
and UO_1280 (O_1280,N_14888,N_14971);
nor UO_1281 (O_1281,N_14881,N_14902);
or UO_1282 (O_1282,N_14968,N_14811);
nand UO_1283 (O_1283,N_14935,N_14986);
and UO_1284 (O_1284,N_14808,N_14896);
or UO_1285 (O_1285,N_14994,N_14999);
nor UO_1286 (O_1286,N_14989,N_14789);
nand UO_1287 (O_1287,N_14771,N_14997);
and UO_1288 (O_1288,N_14781,N_14907);
or UO_1289 (O_1289,N_14874,N_14768);
and UO_1290 (O_1290,N_14968,N_14997);
or UO_1291 (O_1291,N_14953,N_14819);
xor UO_1292 (O_1292,N_14761,N_14766);
nor UO_1293 (O_1293,N_14884,N_14805);
nor UO_1294 (O_1294,N_14865,N_14935);
nor UO_1295 (O_1295,N_14833,N_14882);
nand UO_1296 (O_1296,N_14873,N_14986);
xnor UO_1297 (O_1297,N_14963,N_14899);
nand UO_1298 (O_1298,N_14962,N_14955);
nand UO_1299 (O_1299,N_14831,N_14928);
and UO_1300 (O_1300,N_14998,N_14912);
nand UO_1301 (O_1301,N_14814,N_14809);
xnor UO_1302 (O_1302,N_14969,N_14773);
or UO_1303 (O_1303,N_14885,N_14991);
and UO_1304 (O_1304,N_14931,N_14773);
nor UO_1305 (O_1305,N_14937,N_14806);
nor UO_1306 (O_1306,N_14941,N_14808);
xnor UO_1307 (O_1307,N_14769,N_14933);
nor UO_1308 (O_1308,N_14974,N_14894);
nor UO_1309 (O_1309,N_14897,N_14935);
or UO_1310 (O_1310,N_14870,N_14983);
nand UO_1311 (O_1311,N_14959,N_14779);
or UO_1312 (O_1312,N_14926,N_14968);
nor UO_1313 (O_1313,N_14768,N_14854);
and UO_1314 (O_1314,N_14871,N_14767);
nor UO_1315 (O_1315,N_14988,N_14821);
nand UO_1316 (O_1316,N_14989,N_14760);
nor UO_1317 (O_1317,N_14811,N_14965);
xnor UO_1318 (O_1318,N_14819,N_14848);
and UO_1319 (O_1319,N_14817,N_14932);
nand UO_1320 (O_1320,N_14812,N_14918);
and UO_1321 (O_1321,N_14855,N_14794);
and UO_1322 (O_1322,N_14775,N_14952);
or UO_1323 (O_1323,N_14841,N_14823);
xnor UO_1324 (O_1324,N_14888,N_14812);
nand UO_1325 (O_1325,N_14819,N_14975);
nor UO_1326 (O_1326,N_14961,N_14874);
and UO_1327 (O_1327,N_14753,N_14885);
and UO_1328 (O_1328,N_14866,N_14847);
nand UO_1329 (O_1329,N_14842,N_14791);
nand UO_1330 (O_1330,N_14893,N_14860);
or UO_1331 (O_1331,N_14814,N_14901);
nor UO_1332 (O_1332,N_14799,N_14766);
or UO_1333 (O_1333,N_14863,N_14983);
or UO_1334 (O_1334,N_14897,N_14893);
xor UO_1335 (O_1335,N_14839,N_14793);
xor UO_1336 (O_1336,N_14970,N_14971);
xor UO_1337 (O_1337,N_14754,N_14919);
xor UO_1338 (O_1338,N_14861,N_14829);
or UO_1339 (O_1339,N_14916,N_14794);
nand UO_1340 (O_1340,N_14980,N_14821);
nand UO_1341 (O_1341,N_14786,N_14982);
xor UO_1342 (O_1342,N_14845,N_14976);
nand UO_1343 (O_1343,N_14955,N_14852);
nand UO_1344 (O_1344,N_14784,N_14846);
xor UO_1345 (O_1345,N_14862,N_14979);
xor UO_1346 (O_1346,N_14798,N_14892);
nand UO_1347 (O_1347,N_14799,N_14757);
and UO_1348 (O_1348,N_14888,N_14840);
nor UO_1349 (O_1349,N_14850,N_14771);
and UO_1350 (O_1350,N_14964,N_14949);
xor UO_1351 (O_1351,N_14906,N_14766);
xnor UO_1352 (O_1352,N_14758,N_14805);
nor UO_1353 (O_1353,N_14810,N_14783);
nand UO_1354 (O_1354,N_14998,N_14864);
nand UO_1355 (O_1355,N_14795,N_14796);
or UO_1356 (O_1356,N_14873,N_14866);
xnor UO_1357 (O_1357,N_14828,N_14947);
nand UO_1358 (O_1358,N_14974,N_14992);
xnor UO_1359 (O_1359,N_14770,N_14768);
nor UO_1360 (O_1360,N_14793,N_14801);
xnor UO_1361 (O_1361,N_14926,N_14995);
nand UO_1362 (O_1362,N_14880,N_14793);
nor UO_1363 (O_1363,N_14971,N_14805);
and UO_1364 (O_1364,N_14785,N_14937);
xnor UO_1365 (O_1365,N_14936,N_14810);
and UO_1366 (O_1366,N_14942,N_14983);
and UO_1367 (O_1367,N_14989,N_14852);
nand UO_1368 (O_1368,N_14959,N_14992);
or UO_1369 (O_1369,N_14874,N_14882);
or UO_1370 (O_1370,N_14958,N_14956);
nor UO_1371 (O_1371,N_14820,N_14916);
and UO_1372 (O_1372,N_14860,N_14766);
nor UO_1373 (O_1373,N_14898,N_14875);
xnor UO_1374 (O_1374,N_14932,N_14890);
and UO_1375 (O_1375,N_14850,N_14786);
xnor UO_1376 (O_1376,N_14985,N_14781);
or UO_1377 (O_1377,N_14779,N_14917);
xor UO_1378 (O_1378,N_14797,N_14906);
or UO_1379 (O_1379,N_14977,N_14753);
nand UO_1380 (O_1380,N_14860,N_14751);
or UO_1381 (O_1381,N_14992,N_14822);
and UO_1382 (O_1382,N_14804,N_14882);
nor UO_1383 (O_1383,N_14776,N_14951);
and UO_1384 (O_1384,N_14864,N_14768);
and UO_1385 (O_1385,N_14767,N_14873);
and UO_1386 (O_1386,N_14906,N_14958);
nand UO_1387 (O_1387,N_14853,N_14810);
or UO_1388 (O_1388,N_14814,N_14833);
and UO_1389 (O_1389,N_14849,N_14788);
nand UO_1390 (O_1390,N_14815,N_14761);
xnor UO_1391 (O_1391,N_14976,N_14884);
xnor UO_1392 (O_1392,N_14883,N_14964);
or UO_1393 (O_1393,N_14760,N_14874);
xor UO_1394 (O_1394,N_14954,N_14911);
nor UO_1395 (O_1395,N_14988,N_14855);
nand UO_1396 (O_1396,N_14994,N_14853);
or UO_1397 (O_1397,N_14956,N_14970);
or UO_1398 (O_1398,N_14844,N_14842);
and UO_1399 (O_1399,N_14917,N_14961);
xor UO_1400 (O_1400,N_14884,N_14863);
and UO_1401 (O_1401,N_14785,N_14925);
or UO_1402 (O_1402,N_14765,N_14783);
and UO_1403 (O_1403,N_14883,N_14949);
and UO_1404 (O_1404,N_14903,N_14942);
or UO_1405 (O_1405,N_14883,N_14885);
and UO_1406 (O_1406,N_14964,N_14800);
nand UO_1407 (O_1407,N_14829,N_14854);
or UO_1408 (O_1408,N_14822,N_14944);
nand UO_1409 (O_1409,N_14995,N_14874);
and UO_1410 (O_1410,N_14878,N_14780);
nand UO_1411 (O_1411,N_14847,N_14770);
and UO_1412 (O_1412,N_14775,N_14815);
xnor UO_1413 (O_1413,N_14763,N_14756);
and UO_1414 (O_1414,N_14935,N_14996);
and UO_1415 (O_1415,N_14872,N_14807);
and UO_1416 (O_1416,N_14909,N_14817);
xor UO_1417 (O_1417,N_14993,N_14995);
nor UO_1418 (O_1418,N_14907,N_14978);
and UO_1419 (O_1419,N_14889,N_14858);
nand UO_1420 (O_1420,N_14833,N_14878);
nor UO_1421 (O_1421,N_14939,N_14971);
and UO_1422 (O_1422,N_14750,N_14858);
nand UO_1423 (O_1423,N_14752,N_14973);
and UO_1424 (O_1424,N_14801,N_14917);
nand UO_1425 (O_1425,N_14870,N_14762);
or UO_1426 (O_1426,N_14850,N_14973);
xor UO_1427 (O_1427,N_14978,N_14765);
nor UO_1428 (O_1428,N_14798,N_14850);
or UO_1429 (O_1429,N_14896,N_14986);
xnor UO_1430 (O_1430,N_14861,N_14940);
and UO_1431 (O_1431,N_14815,N_14814);
nor UO_1432 (O_1432,N_14943,N_14836);
nand UO_1433 (O_1433,N_14783,N_14867);
or UO_1434 (O_1434,N_14906,N_14828);
xor UO_1435 (O_1435,N_14988,N_14882);
nor UO_1436 (O_1436,N_14993,N_14789);
or UO_1437 (O_1437,N_14840,N_14800);
nor UO_1438 (O_1438,N_14950,N_14838);
and UO_1439 (O_1439,N_14791,N_14966);
xor UO_1440 (O_1440,N_14913,N_14804);
nand UO_1441 (O_1441,N_14774,N_14817);
or UO_1442 (O_1442,N_14805,N_14826);
nor UO_1443 (O_1443,N_14793,N_14836);
or UO_1444 (O_1444,N_14990,N_14958);
xnor UO_1445 (O_1445,N_14960,N_14910);
nor UO_1446 (O_1446,N_14785,N_14903);
and UO_1447 (O_1447,N_14813,N_14919);
or UO_1448 (O_1448,N_14788,N_14801);
xor UO_1449 (O_1449,N_14998,N_14984);
nor UO_1450 (O_1450,N_14949,N_14806);
and UO_1451 (O_1451,N_14837,N_14872);
nor UO_1452 (O_1452,N_14833,N_14961);
nand UO_1453 (O_1453,N_14811,N_14936);
nor UO_1454 (O_1454,N_14985,N_14947);
and UO_1455 (O_1455,N_14962,N_14899);
nor UO_1456 (O_1456,N_14810,N_14820);
xnor UO_1457 (O_1457,N_14798,N_14898);
or UO_1458 (O_1458,N_14876,N_14847);
and UO_1459 (O_1459,N_14983,N_14900);
nand UO_1460 (O_1460,N_14977,N_14815);
or UO_1461 (O_1461,N_14978,N_14887);
nand UO_1462 (O_1462,N_14963,N_14815);
nor UO_1463 (O_1463,N_14943,N_14885);
nand UO_1464 (O_1464,N_14760,N_14791);
or UO_1465 (O_1465,N_14948,N_14901);
xnor UO_1466 (O_1466,N_14918,N_14945);
xor UO_1467 (O_1467,N_14986,N_14811);
and UO_1468 (O_1468,N_14986,N_14957);
and UO_1469 (O_1469,N_14810,N_14790);
nor UO_1470 (O_1470,N_14790,N_14987);
xnor UO_1471 (O_1471,N_14789,N_14782);
nor UO_1472 (O_1472,N_14935,N_14841);
nand UO_1473 (O_1473,N_14823,N_14906);
xor UO_1474 (O_1474,N_14752,N_14923);
xnor UO_1475 (O_1475,N_14867,N_14938);
and UO_1476 (O_1476,N_14791,N_14858);
or UO_1477 (O_1477,N_14800,N_14846);
and UO_1478 (O_1478,N_14938,N_14840);
and UO_1479 (O_1479,N_14825,N_14941);
nand UO_1480 (O_1480,N_14863,N_14750);
nand UO_1481 (O_1481,N_14969,N_14925);
or UO_1482 (O_1482,N_14949,N_14865);
xnor UO_1483 (O_1483,N_14857,N_14836);
or UO_1484 (O_1484,N_14774,N_14820);
nor UO_1485 (O_1485,N_14780,N_14847);
and UO_1486 (O_1486,N_14817,N_14873);
xnor UO_1487 (O_1487,N_14845,N_14990);
or UO_1488 (O_1488,N_14903,N_14880);
and UO_1489 (O_1489,N_14908,N_14991);
or UO_1490 (O_1490,N_14842,N_14963);
xnor UO_1491 (O_1491,N_14816,N_14762);
xor UO_1492 (O_1492,N_14965,N_14975);
or UO_1493 (O_1493,N_14824,N_14923);
xor UO_1494 (O_1494,N_14852,N_14824);
nor UO_1495 (O_1495,N_14814,N_14785);
or UO_1496 (O_1496,N_14900,N_14977);
nor UO_1497 (O_1497,N_14789,N_14834);
and UO_1498 (O_1498,N_14790,N_14812);
and UO_1499 (O_1499,N_14847,N_14831);
or UO_1500 (O_1500,N_14754,N_14836);
nor UO_1501 (O_1501,N_14770,N_14890);
and UO_1502 (O_1502,N_14794,N_14969);
or UO_1503 (O_1503,N_14967,N_14935);
xor UO_1504 (O_1504,N_14830,N_14954);
or UO_1505 (O_1505,N_14954,N_14756);
nor UO_1506 (O_1506,N_14932,N_14819);
nand UO_1507 (O_1507,N_14812,N_14757);
xor UO_1508 (O_1508,N_14863,N_14845);
xor UO_1509 (O_1509,N_14862,N_14804);
nand UO_1510 (O_1510,N_14829,N_14973);
xor UO_1511 (O_1511,N_14956,N_14842);
xnor UO_1512 (O_1512,N_14864,N_14877);
nand UO_1513 (O_1513,N_14846,N_14752);
and UO_1514 (O_1514,N_14933,N_14898);
nand UO_1515 (O_1515,N_14944,N_14977);
or UO_1516 (O_1516,N_14804,N_14953);
nor UO_1517 (O_1517,N_14847,N_14809);
or UO_1518 (O_1518,N_14995,N_14770);
xnor UO_1519 (O_1519,N_14877,N_14869);
xnor UO_1520 (O_1520,N_14825,N_14838);
xor UO_1521 (O_1521,N_14947,N_14898);
xor UO_1522 (O_1522,N_14978,N_14807);
nor UO_1523 (O_1523,N_14867,N_14810);
and UO_1524 (O_1524,N_14923,N_14989);
nand UO_1525 (O_1525,N_14933,N_14890);
nand UO_1526 (O_1526,N_14967,N_14897);
xnor UO_1527 (O_1527,N_14781,N_14965);
nor UO_1528 (O_1528,N_14883,N_14987);
nor UO_1529 (O_1529,N_14870,N_14834);
or UO_1530 (O_1530,N_14874,N_14879);
nor UO_1531 (O_1531,N_14994,N_14958);
and UO_1532 (O_1532,N_14827,N_14925);
or UO_1533 (O_1533,N_14910,N_14817);
or UO_1534 (O_1534,N_14943,N_14915);
xor UO_1535 (O_1535,N_14982,N_14933);
nand UO_1536 (O_1536,N_14759,N_14824);
nand UO_1537 (O_1537,N_14910,N_14849);
nor UO_1538 (O_1538,N_14906,N_14789);
or UO_1539 (O_1539,N_14794,N_14826);
and UO_1540 (O_1540,N_14847,N_14757);
nor UO_1541 (O_1541,N_14795,N_14985);
xor UO_1542 (O_1542,N_14822,N_14969);
nand UO_1543 (O_1543,N_14901,N_14844);
and UO_1544 (O_1544,N_14817,N_14885);
xnor UO_1545 (O_1545,N_14818,N_14853);
nor UO_1546 (O_1546,N_14805,N_14792);
nand UO_1547 (O_1547,N_14770,N_14884);
nor UO_1548 (O_1548,N_14928,N_14757);
xor UO_1549 (O_1549,N_14934,N_14846);
nor UO_1550 (O_1550,N_14833,N_14843);
nor UO_1551 (O_1551,N_14756,N_14911);
xor UO_1552 (O_1552,N_14896,N_14889);
nor UO_1553 (O_1553,N_14940,N_14768);
nand UO_1554 (O_1554,N_14951,N_14912);
xnor UO_1555 (O_1555,N_14988,N_14879);
or UO_1556 (O_1556,N_14819,N_14771);
xor UO_1557 (O_1557,N_14798,N_14997);
or UO_1558 (O_1558,N_14914,N_14843);
nand UO_1559 (O_1559,N_14934,N_14991);
or UO_1560 (O_1560,N_14750,N_14788);
and UO_1561 (O_1561,N_14960,N_14851);
nor UO_1562 (O_1562,N_14940,N_14758);
nand UO_1563 (O_1563,N_14764,N_14833);
nor UO_1564 (O_1564,N_14915,N_14981);
nor UO_1565 (O_1565,N_14810,N_14980);
nor UO_1566 (O_1566,N_14962,N_14952);
xor UO_1567 (O_1567,N_14765,N_14897);
nor UO_1568 (O_1568,N_14886,N_14885);
and UO_1569 (O_1569,N_14921,N_14756);
and UO_1570 (O_1570,N_14952,N_14757);
nand UO_1571 (O_1571,N_14942,N_14890);
nand UO_1572 (O_1572,N_14854,N_14992);
nand UO_1573 (O_1573,N_14970,N_14776);
nand UO_1574 (O_1574,N_14995,N_14938);
and UO_1575 (O_1575,N_14756,N_14854);
and UO_1576 (O_1576,N_14879,N_14758);
xor UO_1577 (O_1577,N_14829,N_14848);
nand UO_1578 (O_1578,N_14874,N_14753);
nand UO_1579 (O_1579,N_14928,N_14972);
and UO_1580 (O_1580,N_14844,N_14921);
and UO_1581 (O_1581,N_14862,N_14784);
xor UO_1582 (O_1582,N_14928,N_14953);
nor UO_1583 (O_1583,N_14805,N_14800);
or UO_1584 (O_1584,N_14837,N_14925);
and UO_1585 (O_1585,N_14789,N_14963);
or UO_1586 (O_1586,N_14965,N_14936);
nor UO_1587 (O_1587,N_14957,N_14898);
or UO_1588 (O_1588,N_14932,N_14903);
or UO_1589 (O_1589,N_14932,N_14967);
and UO_1590 (O_1590,N_14880,N_14832);
nor UO_1591 (O_1591,N_14817,N_14993);
and UO_1592 (O_1592,N_14844,N_14903);
nor UO_1593 (O_1593,N_14764,N_14840);
nand UO_1594 (O_1594,N_14895,N_14925);
nor UO_1595 (O_1595,N_14931,N_14806);
or UO_1596 (O_1596,N_14803,N_14931);
nand UO_1597 (O_1597,N_14887,N_14910);
nor UO_1598 (O_1598,N_14819,N_14946);
nor UO_1599 (O_1599,N_14807,N_14855);
nand UO_1600 (O_1600,N_14993,N_14756);
nor UO_1601 (O_1601,N_14869,N_14817);
xnor UO_1602 (O_1602,N_14824,N_14862);
and UO_1603 (O_1603,N_14826,N_14773);
nor UO_1604 (O_1604,N_14931,N_14859);
or UO_1605 (O_1605,N_14898,N_14950);
nor UO_1606 (O_1606,N_14898,N_14909);
xnor UO_1607 (O_1607,N_14962,N_14935);
nand UO_1608 (O_1608,N_14854,N_14921);
or UO_1609 (O_1609,N_14973,N_14767);
nor UO_1610 (O_1610,N_14925,N_14816);
or UO_1611 (O_1611,N_14958,N_14917);
or UO_1612 (O_1612,N_14859,N_14973);
nand UO_1613 (O_1613,N_14788,N_14949);
and UO_1614 (O_1614,N_14750,N_14865);
or UO_1615 (O_1615,N_14807,N_14932);
or UO_1616 (O_1616,N_14874,N_14962);
or UO_1617 (O_1617,N_14780,N_14959);
nand UO_1618 (O_1618,N_14977,N_14765);
and UO_1619 (O_1619,N_14909,N_14893);
xnor UO_1620 (O_1620,N_14882,N_14808);
or UO_1621 (O_1621,N_14804,N_14854);
and UO_1622 (O_1622,N_14769,N_14782);
xor UO_1623 (O_1623,N_14815,N_14818);
and UO_1624 (O_1624,N_14827,N_14757);
or UO_1625 (O_1625,N_14959,N_14774);
xor UO_1626 (O_1626,N_14993,N_14765);
or UO_1627 (O_1627,N_14991,N_14921);
or UO_1628 (O_1628,N_14934,N_14849);
or UO_1629 (O_1629,N_14900,N_14894);
and UO_1630 (O_1630,N_14822,N_14875);
or UO_1631 (O_1631,N_14785,N_14894);
nor UO_1632 (O_1632,N_14836,N_14872);
nor UO_1633 (O_1633,N_14968,N_14815);
or UO_1634 (O_1634,N_14842,N_14847);
or UO_1635 (O_1635,N_14926,N_14814);
or UO_1636 (O_1636,N_14815,N_14940);
nor UO_1637 (O_1637,N_14937,N_14859);
nand UO_1638 (O_1638,N_14975,N_14802);
and UO_1639 (O_1639,N_14989,N_14830);
nor UO_1640 (O_1640,N_14780,N_14801);
xor UO_1641 (O_1641,N_14884,N_14896);
xnor UO_1642 (O_1642,N_14821,N_14936);
and UO_1643 (O_1643,N_14849,N_14984);
nor UO_1644 (O_1644,N_14758,N_14911);
xor UO_1645 (O_1645,N_14982,N_14819);
nor UO_1646 (O_1646,N_14997,N_14758);
or UO_1647 (O_1647,N_14979,N_14755);
nor UO_1648 (O_1648,N_14793,N_14815);
or UO_1649 (O_1649,N_14884,N_14913);
nor UO_1650 (O_1650,N_14917,N_14898);
nand UO_1651 (O_1651,N_14876,N_14816);
xnor UO_1652 (O_1652,N_14888,N_14905);
nor UO_1653 (O_1653,N_14866,N_14811);
and UO_1654 (O_1654,N_14776,N_14803);
and UO_1655 (O_1655,N_14924,N_14915);
nand UO_1656 (O_1656,N_14763,N_14971);
nor UO_1657 (O_1657,N_14836,N_14820);
xnor UO_1658 (O_1658,N_14819,N_14990);
nor UO_1659 (O_1659,N_14854,N_14825);
nand UO_1660 (O_1660,N_14855,N_14793);
nor UO_1661 (O_1661,N_14792,N_14869);
or UO_1662 (O_1662,N_14903,N_14831);
or UO_1663 (O_1663,N_14880,N_14932);
or UO_1664 (O_1664,N_14898,N_14952);
xnor UO_1665 (O_1665,N_14839,N_14949);
or UO_1666 (O_1666,N_14846,N_14867);
nor UO_1667 (O_1667,N_14832,N_14991);
and UO_1668 (O_1668,N_14904,N_14861);
xnor UO_1669 (O_1669,N_14799,N_14926);
nor UO_1670 (O_1670,N_14826,N_14857);
xor UO_1671 (O_1671,N_14766,N_14835);
xor UO_1672 (O_1672,N_14884,N_14909);
nor UO_1673 (O_1673,N_14787,N_14959);
and UO_1674 (O_1674,N_14796,N_14753);
nand UO_1675 (O_1675,N_14836,N_14826);
or UO_1676 (O_1676,N_14804,N_14835);
nand UO_1677 (O_1677,N_14966,N_14831);
xor UO_1678 (O_1678,N_14867,N_14990);
xnor UO_1679 (O_1679,N_14893,N_14936);
nor UO_1680 (O_1680,N_14818,N_14782);
xnor UO_1681 (O_1681,N_14919,N_14881);
nor UO_1682 (O_1682,N_14922,N_14871);
nor UO_1683 (O_1683,N_14759,N_14875);
nand UO_1684 (O_1684,N_14892,N_14818);
nor UO_1685 (O_1685,N_14872,N_14798);
and UO_1686 (O_1686,N_14964,N_14966);
or UO_1687 (O_1687,N_14847,N_14865);
and UO_1688 (O_1688,N_14820,N_14824);
nor UO_1689 (O_1689,N_14975,N_14833);
nand UO_1690 (O_1690,N_14906,N_14824);
nor UO_1691 (O_1691,N_14973,N_14917);
nor UO_1692 (O_1692,N_14927,N_14949);
nand UO_1693 (O_1693,N_14785,N_14786);
xor UO_1694 (O_1694,N_14934,N_14925);
and UO_1695 (O_1695,N_14914,N_14952);
nor UO_1696 (O_1696,N_14812,N_14805);
nand UO_1697 (O_1697,N_14752,N_14907);
nand UO_1698 (O_1698,N_14852,N_14833);
nor UO_1699 (O_1699,N_14877,N_14967);
nand UO_1700 (O_1700,N_14909,N_14870);
xnor UO_1701 (O_1701,N_14899,N_14959);
or UO_1702 (O_1702,N_14763,N_14821);
and UO_1703 (O_1703,N_14864,N_14974);
nor UO_1704 (O_1704,N_14767,N_14917);
nand UO_1705 (O_1705,N_14839,N_14825);
or UO_1706 (O_1706,N_14752,N_14977);
or UO_1707 (O_1707,N_14974,N_14789);
nor UO_1708 (O_1708,N_14805,N_14864);
nor UO_1709 (O_1709,N_14999,N_14966);
xnor UO_1710 (O_1710,N_14981,N_14816);
xnor UO_1711 (O_1711,N_14792,N_14955);
xor UO_1712 (O_1712,N_14893,N_14964);
or UO_1713 (O_1713,N_14774,N_14758);
and UO_1714 (O_1714,N_14766,N_14756);
and UO_1715 (O_1715,N_14981,N_14938);
nand UO_1716 (O_1716,N_14769,N_14787);
nand UO_1717 (O_1717,N_14757,N_14967);
xor UO_1718 (O_1718,N_14953,N_14951);
nand UO_1719 (O_1719,N_14856,N_14769);
or UO_1720 (O_1720,N_14883,N_14842);
nand UO_1721 (O_1721,N_14935,N_14766);
nor UO_1722 (O_1722,N_14982,N_14816);
nand UO_1723 (O_1723,N_14777,N_14812);
xor UO_1724 (O_1724,N_14972,N_14872);
or UO_1725 (O_1725,N_14811,N_14969);
or UO_1726 (O_1726,N_14986,N_14818);
or UO_1727 (O_1727,N_14974,N_14768);
nor UO_1728 (O_1728,N_14839,N_14934);
xor UO_1729 (O_1729,N_14908,N_14804);
xnor UO_1730 (O_1730,N_14987,N_14982);
or UO_1731 (O_1731,N_14787,N_14838);
nand UO_1732 (O_1732,N_14888,N_14936);
or UO_1733 (O_1733,N_14941,N_14879);
and UO_1734 (O_1734,N_14777,N_14826);
nand UO_1735 (O_1735,N_14908,N_14983);
or UO_1736 (O_1736,N_14841,N_14807);
nor UO_1737 (O_1737,N_14794,N_14820);
nor UO_1738 (O_1738,N_14909,N_14789);
and UO_1739 (O_1739,N_14904,N_14802);
xnor UO_1740 (O_1740,N_14862,N_14855);
or UO_1741 (O_1741,N_14898,N_14835);
or UO_1742 (O_1742,N_14918,N_14828);
nand UO_1743 (O_1743,N_14942,N_14973);
xor UO_1744 (O_1744,N_14981,N_14994);
and UO_1745 (O_1745,N_14964,N_14775);
xnor UO_1746 (O_1746,N_14968,N_14751);
xnor UO_1747 (O_1747,N_14844,N_14953);
or UO_1748 (O_1748,N_14814,N_14934);
nor UO_1749 (O_1749,N_14935,N_14970);
and UO_1750 (O_1750,N_14751,N_14779);
and UO_1751 (O_1751,N_14861,N_14987);
xor UO_1752 (O_1752,N_14964,N_14791);
nand UO_1753 (O_1753,N_14907,N_14905);
nand UO_1754 (O_1754,N_14862,N_14923);
or UO_1755 (O_1755,N_14928,N_14978);
and UO_1756 (O_1756,N_14889,N_14952);
and UO_1757 (O_1757,N_14821,N_14983);
or UO_1758 (O_1758,N_14856,N_14909);
or UO_1759 (O_1759,N_14856,N_14843);
nor UO_1760 (O_1760,N_14899,N_14900);
or UO_1761 (O_1761,N_14844,N_14793);
nor UO_1762 (O_1762,N_14969,N_14832);
xor UO_1763 (O_1763,N_14882,N_14896);
nand UO_1764 (O_1764,N_14897,N_14866);
nand UO_1765 (O_1765,N_14771,N_14940);
nand UO_1766 (O_1766,N_14998,N_14785);
nor UO_1767 (O_1767,N_14806,N_14773);
nand UO_1768 (O_1768,N_14787,N_14882);
xor UO_1769 (O_1769,N_14898,N_14794);
or UO_1770 (O_1770,N_14999,N_14796);
nand UO_1771 (O_1771,N_14876,N_14925);
and UO_1772 (O_1772,N_14983,N_14868);
xor UO_1773 (O_1773,N_14923,N_14753);
or UO_1774 (O_1774,N_14938,N_14766);
nor UO_1775 (O_1775,N_14950,N_14769);
xnor UO_1776 (O_1776,N_14926,N_14817);
nand UO_1777 (O_1777,N_14850,N_14901);
nand UO_1778 (O_1778,N_14973,N_14892);
xor UO_1779 (O_1779,N_14891,N_14948);
nand UO_1780 (O_1780,N_14753,N_14879);
nor UO_1781 (O_1781,N_14897,N_14870);
or UO_1782 (O_1782,N_14935,N_14889);
xnor UO_1783 (O_1783,N_14917,N_14889);
or UO_1784 (O_1784,N_14806,N_14816);
or UO_1785 (O_1785,N_14951,N_14791);
or UO_1786 (O_1786,N_14974,N_14970);
nor UO_1787 (O_1787,N_14801,N_14940);
xnor UO_1788 (O_1788,N_14997,N_14907);
and UO_1789 (O_1789,N_14819,N_14816);
nor UO_1790 (O_1790,N_14985,N_14874);
nor UO_1791 (O_1791,N_14850,N_14817);
nand UO_1792 (O_1792,N_14889,N_14968);
nand UO_1793 (O_1793,N_14804,N_14864);
nand UO_1794 (O_1794,N_14884,N_14967);
nand UO_1795 (O_1795,N_14955,N_14768);
and UO_1796 (O_1796,N_14777,N_14987);
and UO_1797 (O_1797,N_14756,N_14994);
or UO_1798 (O_1798,N_14800,N_14978);
nor UO_1799 (O_1799,N_14898,N_14974);
nor UO_1800 (O_1800,N_14779,N_14973);
nand UO_1801 (O_1801,N_14844,N_14888);
xnor UO_1802 (O_1802,N_14818,N_14953);
xor UO_1803 (O_1803,N_14780,N_14997);
or UO_1804 (O_1804,N_14928,N_14935);
nand UO_1805 (O_1805,N_14950,N_14956);
nand UO_1806 (O_1806,N_14807,N_14928);
nand UO_1807 (O_1807,N_14875,N_14842);
and UO_1808 (O_1808,N_14951,N_14772);
or UO_1809 (O_1809,N_14809,N_14910);
or UO_1810 (O_1810,N_14981,N_14837);
nand UO_1811 (O_1811,N_14901,N_14793);
or UO_1812 (O_1812,N_14888,N_14803);
nand UO_1813 (O_1813,N_14932,N_14758);
nor UO_1814 (O_1814,N_14888,N_14993);
and UO_1815 (O_1815,N_14914,N_14812);
nand UO_1816 (O_1816,N_14819,N_14937);
nand UO_1817 (O_1817,N_14801,N_14763);
nor UO_1818 (O_1818,N_14805,N_14951);
and UO_1819 (O_1819,N_14792,N_14823);
nand UO_1820 (O_1820,N_14929,N_14882);
xor UO_1821 (O_1821,N_14924,N_14945);
or UO_1822 (O_1822,N_14873,N_14845);
nand UO_1823 (O_1823,N_14900,N_14932);
and UO_1824 (O_1824,N_14828,N_14827);
xor UO_1825 (O_1825,N_14882,N_14873);
xor UO_1826 (O_1826,N_14799,N_14800);
xnor UO_1827 (O_1827,N_14903,N_14971);
and UO_1828 (O_1828,N_14819,N_14900);
and UO_1829 (O_1829,N_14919,N_14863);
nor UO_1830 (O_1830,N_14897,N_14826);
and UO_1831 (O_1831,N_14817,N_14776);
nor UO_1832 (O_1832,N_14751,N_14832);
nand UO_1833 (O_1833,N_14860,N_14923);
nand UO_1834 (O_1834,N_14836,N_14780);
nand UO_1835 (O_1835,N_14780,N_14994);
or UO_1836 (O_1836,N_14889,N_14946);
and UO_1837 (O_1837,N_14917,N_14860);
and UO_1838 (O_1838,N_14894,N_14788);
nor UO_1839 (O_1839,N_14767,N_14765);
nor UO_1840 (O_1840,N_14894,N_14955);
or UO_1841 (O_1841,N_14924,N_14927);
and UO_1842 (O_1842,N_14817,N_14998);
xor UO_1843 (O_1843,N_14871,N_14859);
xor UO_1844 (O_1844,N_14995,N_14917);
and UO_1845 (O_1845,N_14792,N_14802);
nand UO_1846 (O_1846,N_14832,N_14777);
nand UO_1847 (O_1847,N_14948,N_14753);
nor UO_1848 (O_1848,N_14910,N_14814);
nor UO_1849 (O_1849,N_14904,N_14757);
and UO_1850 (O_1850,N_14909,N_14813);
nand UO_1851 (O_1851,N_14816,N_14869);
nand UO_1852 (O_1852,N_14971,N_14972);
nor UO_1853 (O_1853,N_14993,N_14793);
and UO_1854 (O_1854,N_14978,N_14923);
xnor UO_1855 (O_1855,N_14791,N_14985);
or UO_1856 (O_1856,N_14939,N_14929);
and UO_1857 (O_1857,N_14881,N_14791);
nand UO_1858 (O_1858,N_14985,N_14824);
and UO_1859 (O_1859,N_14956,N_14919);
xnor UO_1860 (O_1860,N_14754,N_14779);
xor UO_1861 (O_1861,N_14977,N_14953);
nor UO_1862 (O_1862,N_14987,N_14764);
or UO_1863 (O_1863,N_14961,N_14824);
and UO_1864 (O_1864,N_14761,N_14858);
and UO_1865 (O_1865,N_14832,N_14853);
and UO_1866 (O_1866,N_14993,N_14931);
and UO_1867 (O_1867,N_14911,N_14907);
nor UO_1868 (O_1868,N_14825,N_14836);
and UO_1869 (O_1869,N_14893,N_14837);
nor UO_1870 (O_1870,N_14784,N_14864);
and UO_1871 (O_1871,N_14981,N_14806);
nor UO_1872 (O_1872,N_14960,N_14890);
xnor UO_1873 (O_1873,N_14945,N_14961);
and UO_1874 (O_1874,N_14857,N_14853);
nor UO_1875 (O_1875,N_14879,N_14999);
nor UO_1876 (O_1876,N_14757,N_14783);
nor UO_1877 (O_1877,N_14879,N_14776);
nor UO_1878 (O_1878,N_14841,N_14827);
xnor UO_1879 (O_1879,N_14916,N_14766);
nand UO_1880 (O_1880,N_14911,N_14857);
and UO_1881 (O_1881,N_14830,N_14763);
xnor UO_1882 (O_1882,N_14815,N_14819);
or UO_1883 (O_1883,N_14769,N_14817);
or UO_1884 (O_1884,N_14934,N_14945);
and UO_1885 (O_1885,N_14852,N_14983);
xor UO_1886 (O_1886,N_14892,N_14861);
and UO_1887 (O_1887,N_14759,N_14843);
nor UO_1888 (O_1888,N_14806,N_14789);
nor UO_1889 (O_1889,N_14914,N_14998);
and UO_1890 (O_1890,N_14888,N_14950);
nand UO_1891 (O_1891,N_14765,N_14796);
xor UO_1892 (O_1892,N_14961,N_14975);
and UO_1893 (O_1893,N_14948,N_14915);
nand UO_1894 (O_1894,N_14895,N_14850);
or UO_1895 (O_1895,N_14977,N_14859);
and UO_1896 (O_1896,N_14878,N_14896);
xor UO_1897 (O_1897,N_14755,N_14889);
or UO_1898 (O_1898,N_14765,N_14976);
or UO_1899 (O_1899,N_14815,N_14790);
and UO_1900 (O_1900,N_14817,N_14995);
nor UO_1901 (O_1901,N_14790,N_14957);
or UO_1902 (O_1902,N_14828,N_14878);
nor UO_1903 (O_1903,N_14913,N_14796);
and UO_1904 (O_1904,N_14799,N_14847);
or UO_1905 (O_1905,N_14939,N_14914);
nor UO_1906 (O_1906,N_14903,N_14773);
nand UO_1907 (O_1907,N_14768,N_14932);
or UO_1908 (O_1908,N_14941,N_14781);
nand UO_1909 (O_1909,N_14831,N_14870);
or UO_1910 (O_1910,N_14905,N_14824);
and UO_1911 (O_1911,N_14759,N_14832);
xor UO_1912 (O_1912,N_14987,N_14822);
nand UO_1913 (O_1913,N_14982,N_14809);
and UO_1914 (O_1914,N_14811,N_14991);
or UO_1915 (O_1915,N_14979,N_14751);
nor UO_1916 (O_1916,N_14851,N_14752);
nor UO_1917 (O_1917,N_14804,N_14805);
xor UO_1918 (O_1918,N_14989,N_14950);
nor UO_1919 (O_1919,N_14814,N_14992);
or UO_1920 (O_1920,N_14848,N_14988);
or UO_1921 (O_1921,N_14775,N_14774);
nand UO_1922 (O_1922,N_14763,N_14951);
xor UO_1923 (O_1923,N_14891,N_14902);
nand UO_1924 (O_1924,N_14791,N_14778);
nand UO_1925 (O_1925,N_14771,N_14934);
or UO_1926 (O_1926,N_14953,N_14856);
and UO_1927 (O_1927,N_14788,N_14809);
xnor UO_1928 (O_1928,N_14885,N_14788);
or UO_1929 (O_1929,N_14993,N_14889);
nor UO_1930 (O_1930,N_14967,N_14787);
nand UO_1931 (O_1931,N_14933,N_14984);
nand UO_1932 (O_1932,N_14991,N_14975);
and UO_1933 (O_1933,N_14811,N_14861);
xor UO_1934 (O_1934,N_14904,N_14786);
xor UO_1935 (O_1935,N_14852,N_14758);
nand UO_1936 (O_1936,N_14967,N_14904);
nor UO_1937 (O_1937,N_14876,N_14811);
or UO_1938 (O_1938,N_14857,N_14918);
and UO_1939 (O_1939,N_14843,N_14798);
nor UO_1940 (O_1940,N_14989,N_14976);
nor UO_1941 (O_1941,N_14838,N_14896);
and UO_1942 (O_1942,N_14895,N_14908);
or UO_1943 (O_1943,N_14891,N_14768);
or UO_1944 (O_1944,N_14912,N_14970);
xor UO_1945 (O_1945,N_14849,N_14752);
nand UO_1946 (O_1946,N_14863,N_14876);
nor UO_1947 (O_1947,N_14841,N_14922);
or UO_1948 (O_1948,N_14778,N_14903);
nor UO_1949 (O_1949,N_14773,N_14758);
nor UO_1950 (O_1950,N_14964,N_14902);
and UO_1951 (O_1951,N_14909,N_14908);
nor UO_1952 (O_1952,N_14767,N_14998);
nand UO_1953 (O_1953,N_14942,N_14794);
nor UO_1954 (O_1954,N_14933,N_14913);
nand UO_1955 (O_1955,N_14924,N_14966);
nor UO_1956 (O_1956,N_14838,N_14819);
or UO_1957 (O_1957,N_14946,N_14757);
or UO_1958 (O_1958,N_14923,N_14772);
nor UO_1959 (O_1959,N_14903,N_14879);
and UO_1960 (O_1960,N_14814,N_14755);
or UO_1961 (O_1961,N_14931,N_14880);
and UO_1962 (O_1962,N_14907,N_14868);
and UO_1963 (O_1963,N_14853,N_14783);
and UO_1964 (O_1964,N_14764,N_14760);
nor UO_1965 (O_1965,N_14991,N_14796);
xnor UO_1966 (O_1966,N_14940,N_14877);
nor UO_1967 (O_1967,N_14980,N_14917);
nor UO_1968 (O_1968,N_14921,N_14780);
or UO_1969 (O_1969,N_14844,N_14985);
or UO_1970 (O_1970,N_14896,N_14765);
xor UO_1971 (O_1971,N_14823,N_14909);
or UO_1972 (O_1972,N_14782,N_14989);
and UO_1973 (O_1973,N_14855,N_14843);
xnor UO_1974 (O_1974,N_14866,N_14999);
nand UO_1975 (O_1975,N_14781,N_14769);
and UO_1976 (O_1976,N_14835,N_14867);
nor UO_1977 (O_1977,N_14996,N_14871);
nand UO_1978 (O_1978,N_14868,N_14957);
nand UO_1979 (O_1979,N_14940,N_14783);
and UO_1980 (O_1980,N_14922,N_14925);
nand UO_1981 (O_1981,N_14976,N_14947);
or UO_1982 (O_1982,N_14964,N_14861);
and UO_1983 (O_1983,N_14767,N_14829);
or UO_1984 (O_1984,N_14899,N_14928);
and UO_1985 (O_1985,N_14894,N_14849);
or UO_1986 (O_1986,N_14788,N_14799);
nand UO_1987 (O_1987,N_14856,N_14969);
or UO_1988 (O_1988,N_14758,N_14945);
nand UO_1989 (O_1989,N_14929,N_14758);
or UO_1990 (O_1990,N_14824,N_14800);
nor UO_1991 (O_1991,N_14936,N_14927);
nand UO_1992 (O_1992,N_14926,N_14793);
nand UO_1993 (O_1993,N_14953,N_14992);
and UO_1994 (O_1994,N_14760,N_14975);
nand UO_1995 (O_1995,N_14793,N_14832);
xor UO_1996 (O_1996,N_14765,N_14945);
nand UO_1997 (O_1997,N_14753,N_14974);
xnor UO_1998 (O_1998,N_14983,N_14771);
or UO_1999 (O_1999,N_14816,N_14793);
endmodule