module basic_750_5000_1000_2_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2504,N_2505,N_2506,N_2507,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2553,N_2554,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2565,N_2566,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2584,N_2585,N_2586,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2595,N_2596,N_2597,N_2598,N_2599,N_2601,N_2602,N_2603,N_2604,N_2605,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2618,N_2619,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2629,N_2630,N_2631,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2644,N_2645,N_2647,N_2648,N_2650,N_2651,N_2652,N_2653,N_2654,N_2656,N_2657,N_2658,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2668,N_2669,N_2672,N_2673,N_2674,N_2675,N_2678,N_2679,N_2680,N_2681,N_2682,N_2684,N_2685,N_2686,N_2687,N_2689,N_2691,N_2692,N_2694,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2707,N_2708,N_2709,N_2710,N_2712,N_2713,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2728,N_2729,N_2730,N_2732,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2757,N_2759,N_2760,N_2763,N_2766,N_2767,N_2768,N_2769,N_2771,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2786,N_2788,N_2789,N_2794,N_2795,N_2796,N_2797,N_2798,N_2800,N_2801,N_2802,N_2804,N_2806,N_2807,N_2808,N_2809,N_2810,N_2812,N_2813,N_2814,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2838,N_2839,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2850,N_2852,N_2854,N_2855,N_2856,N_2858,N_2859,N_2861,N_2862,N_2863,N_2864,N_2865,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2874,N_2875,N_2876,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2891,N_2892,N_2893,N_2894,N_2895,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2907,N_2911,N_2912,N_2913,N_2914,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2936,N_2937,N_2938,N_2939,N_2940,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2961,N_2962,N_2964,N_2966,N_2968,N_2969,N_2970,N_2971,N_2973,N_2974,N_2975,N_2976,N_2977,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2987,N_2989,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2999,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3012,N_3013,N_3014,N_3015,N_3017,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3034,N_3035,N_3036,N_3037,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3047,N_3048,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3060,N_3061,N_3062,N_3063,N_3064,N_3067,N_3068,N_3069,N_3070,N_3072,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3084,N_3085,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3116,N_3117,N_3118,N_3119,N_3120,N_3122,N_3125,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3144,N_3146,N_3147,N_3148,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3179,N_3180,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3207,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3224,N_3225,N_3227,N_3228,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3255,N_3256,N_3257,N_3258,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3291,N_3292,N_3293,N_3294,N_3295,N_3297,N_3298,N_3299,N_3300,N_3301,N_3303,N_3304,N_3305,N_3306,N_3309,N_3310,N_3311,N_3312,N_3314,N_3315,N_3317,N_3318,N_3319,N_3320,N_3323,N_3325,N_3327,N_3329,N_3330,N_3331,N_3332,N_3334,N_3336,N_3337,N_3338,N_3339,N_3340,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3349,N_3350,N_3351,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3362,N_3363,N_3364,N_3365,N_3367,N_3369,N_3370,N_3372,N_3373,N_3374,N_3375,N_3376,N_3379,N_3381,N_3382,N_3383,N_3384,N_3386,N_3388,N_3389,N_3390,N_3391,N_3393,N_3394,N_3395,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3411,N_3412,N_3413,N_3414,N_3417,N_3418,N_3420,N_3422,N_3423,N_3424,N_3427,N_3428,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3441,N_3442,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3469,N_3470,N_3472,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3486,N_3488,N_3489,N_3490,N_3491,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3501,N_3502,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3542,N_3543,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3558,N_3559,N_3561,N_3563,N_3564,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3578,N_3579,N_3580,N_3582,N_3583,N_3584,N_3585,N_3586,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3598,N_3599,N_3601,N_3602,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3611,N_3614,N_3616,N_3618,N_3619,N_3620,N_3621,N_3623,N_3624,N_3625,N_3628,N_3629,N_3630,N_3632,N_3633,N_3634,N_3635,N_3637,N_3638,N_3639,N_3640,N_3641,N_3643,N_3645,N_3646,N_3647,N_3648,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3669,N_3670,N_3672,N_3673,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3682,N_3684,N_3685,N_3687,N_3689,N_3690,N_3691,N_3692,N_3694,N_3697,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3706,N_3707,N_3708,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3719,N_3720,N_3721,N_3722,N_3723,N_3725,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3761,N_3762,N_3763,N_3764,N_3765,N_3767,N_3768,N_3769,N_3772,N_3775,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3802,N_3804,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3829,N_3831,N_3833,N_3834,N_3835,N_3837,N_3838,N_3839,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3861,N_3862,N_3863,N_3864,N_3865,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3880,N_3881,N_3882,N_3883,N_3884,N_3887,N_3888,N_3890,N_3891,N_3892,N_3894,N_3897,N_3899,N_3900,N_3901,N_3902,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3920,N_3921,N_3922,N_3923,N_3924,N_3926,N_3927,N_3928,N_3929,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3947,N_3948,N_3949,N_3950,N_3951,N_3955,N_3956,N_3957,N_3958,N_3959,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3983,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3993,N_3994,N_3995,N_3996,N_3998,N_3999,N_4001,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4014,N_4015,N_4016,N_4017,N_4019,N_4020,N_4023,N_4025,N_4026,N_4027,N_4028,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4043,N_4044,N_4045,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4077,N_4078,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4088,N_4092,N_4093,N_4094,N_4095,N_4096,N_4098,N_4099,N_4100,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4109,N_4111,N_4112,N_4113,N_4116,N_4118,N_4119,N_4121,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4142,N_4143,N_4144,N_4145,N_4146,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4158,N_4159,N_4161,N_4162,N_4163,N_4165,N_4166,N_4167,N_4168,N_4172,N_4173,N_4175,N_4176,N_4177,N_4178,N_4180,N_4181,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4219,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4228,N_4229,N_4231,N_4232,N_4233,N_4235,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4247,N_4248,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4262,N_4263,N_4266,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4275,N_4276,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4290,N_4291,N_4293,N_4294,N_4296,N_4298,N_4299,N_4300,N_4302,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4326,N_4328,N_4329,N_4330,N_4331,N_4334,N_4335,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4352,N_4353,N_4354,N_4355,N_4357,N_4358,N_4359,N_4360,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4373,N_4374,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4385,N_4386,N_4387,N_4389,N_4390,N_4391,N_4392,N_4393,N_4395,N_4396,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4408,N_4409,N_4411,N_4412,N_4413,N_4415,N_4416,N_4417,N_4418,N_4419,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4441,N_4443,N_4444,N_4446,N_4447,N_4448,N_4449,N_4451,N_4453,N_4454,N_4455,N_4457,N_4458,N_4459,N_4460,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4479,N_4480,N_4481,N_4483,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4501,N_4503,N_4504,N_4505,N_4506,N_4507,N_4509,N_4511,N_4512,N_4514,N_4516,N_4517,N_4518,N_4519,N_4520,N_4523,N_4527,N_4528,N_4530,N_4531,N_4532,N_4533,N_4535,N_4537,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4550,N_4551,N_4552,N_4553,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4572,N_4574,N_4575,N_4577,N_4578,N_4579,N_4580,N_4581,N_4583,N_4585,N_4586,N_4587,N_4589,N_4590,N_4591,N_4592,N_4595,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4635,N_4636,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4652,N_4653,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4663,N_4664,N_4665,N_4666,N_4667,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4680,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4706,N_4707,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4720,N_4722,N_4723,N_4725,N_4726,N_4728,N_4729,N_4730,N_4731,N_4732,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4744,N_4745,N_4747,N_4748,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4765,N_4766,N_4768,N_4770,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4789,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4800,N_4801,N_4802,N_4803,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4813,N_4816,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4845,N_4847,N_4848,N_4852,N_4854,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4874,N_4875,N_4876,N_4877,N_4879,N_4880,N_4881,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4893,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4915,N_4916,N_4917,N_4920,N_4921,N_4922,N_4923,N_4927,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4938,N_4939,N_4942,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4961,N_4962,N_4963,N_4964,N_4965,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4993,N_4994,N_4995,N_4997,N_4998,N_4999;
or U0 (N_0,In_713,In_26);
nor U1 (N_1,In_659,In_614);
nand U2 (N_2,In_197,In_147);
nor U3 (N_3,In_339,In_608);
and U4 (N_4,In_628,In_86);
and U5 (N_5,In_350,In_437);
or U6 (N_6,In_349,In_128);
or U7 (N_7,In_430,In_66);
nor U8 (N_8,In_553,In_367);
nor U9 (N_9,In_621,In_448);
nor U10 (N_10,In_85,In_48);
and U11 (N_11,In_491,In_724);
and U12 (N_12,In_657,In_172);
nand U13 (N_13,In_573,In_215);
or U14 (N_14,In_120,In_509);
and U15 (N_15,In_81,In_551);
nor U16 (N_16,In_370,In_527);
nand U17 (N_17,In_597,In_188);
nand U18 (N_18,In_598,In_412);
nor U19 (N_19,In_739,In_166);
and U20 (N_20,In_203,In_378);
and U21 (N_21,In_285,In_7);
nor U22 (N_22,In_744,In_136);
nor U23 (N_23,In_70,In_90);
nor U24 (N_24,In_315,In_391);
nand U25 (N_25,In_632,In_725);
nor U26 (N_26,In_112,In_645);
or U27 (N_27,In_497,In_195);
nor U28 (N_28,In_8,In_101);
nor U29 (N_29,In_208,In_624);
and U30 (N_30,In_358,In_150);
nand U31 (N_31,In_173,In_189);
nand U32 (N_32,In_351,In_244);
and U33 (N_33,In_305,In_229);
nand U34 (N_34,In_561,In_319);
and U35 (N_35,In_545,In_143);
nand U36 (N_36,In_424,In_380);
nor U37 (N_37,In_606,In_239);
nor U38 (N_38,In_209,In_673);
nor U39 (N_39,In_276,In_626);
and U40 (N_40,In_248,In_465);
and U41 (N_41,In_408,In_581);
nor U42 (N_42,In_114,In_536);
and U43 (N_43,In_646,In_306);
and U44 (N_44,In_529,In_694);
or U45 (N_45,In_613,In_359);
nor U46 (N_46,In_219,In_261);
nand U47 (N_47,In_51,In_660);
xor U48 (N_48,In_392,In_630);
and U49 (N_49,In_11,In_455);
and U50 (N_50,In_309,In_299);
nand U51 (N_51,In_242,In_201);
nor U52 (N_52,In_708,In_584);
nand U53 (N_53,In_560,In_320);
and U54 (N_54,In_31,In_583);
and U55 (N_55,In_363,In_328);
nor U56 (N_56,In_726,In_185);
or U57 (N_57,In_125,In_35);
nor U58 (N_58,In_282,In_199);
nand U59 (N_59,In_293,In_549);
and U60 (N_60,In_207,In_383);
or U61 (N_61,In_280,In_490);
or U62 (N_62,In_36,In_37);
nor U63 (N_63,In_684,In_402);
or U64 (N_64,In_460,In_464);
nor U65 (N_65,In_458,In_258);
or U66 (N_66,In_662,In_601);
or U67 (N_67,In_685,In_97);
or U68 (N_68,In_555,In_291);
nor U69 (N_69,In_138,In_187);
nand U70 (N_70,In_322,In_177);
or U71 (N_71,In_451,In_107);
or U72 (N_72,In_577,In_418);
or U73 (N_73,In_29,In_655);
nand U74 (N_74,In_272,In_206);
or U75 (N_75,In_661,In_87);
nand U76 (N_76,In_170,In_155);
nand U77 (N_77,In_712,In_263);
and U78 (N_78,In_699,In_308);
or U79 (N_79,In_44,In_639);
or U80 (N_80,In_108,In_268);
nor U81 (N_81,In_670,In_605);
and U82 (N_82,In_434,In_323);
or U83 (N_83,In_116,In_281);
or U84 (N_84,In_579,In_297);
nand U85 (N_85,In_274,In_352);
or U86 (N_86,In_401,In_679);
nand U87 (N_87,In_337,In_167);
nor U88 (N_88,In_611,In_296);
or U89 (N_89,In_362,In_0);
or U90 (N_90,In_531,In_431);
and U91 (N_91,In_225,In_250);
nand U92 (N_92,In_43,In_516);
nand U93 (N_93,In_84,In_278);
or U94 (N_94,In_525,In_519);
and U95 (N_95,In_311,In_449);
nor U96 (N_96,In_444,In_702);
or U97 (N_97,In_39,In_106);
or U98 (N_98,In_571,In_474);
nor U99 (N_99,In_393,In_638);
or U100 (N_100,In_53,In_538);
nand U101 (N_101,In_603,In_60);
nand U102 (N_102,In_144,In_433);
nand U103 (N_103,In_663,In_379);
or U104 (N_104,In_650,In_493);
nor U105 (N_105,In_158,In_316);
and U106 (N_106,In_552,In_484);
or U107 (N_107,In_71,In_740);
and U108 (N_108,In_677,In_422);
or U109 (N_109,In_238,In_686);
or U110 (N_110,In_79,In_676);
nand U111 (N_111,In_723,In_404);
or U112 (N_112,In_477,In_748);
nor U113 (N_113,In_57,In_135);
and U114 (N_114,In_175,In_115);
or U115 (N_115,In_169,In_427);
nand U116 (N_116,In_194,In_667);
nand U117 (N_117,In_18,In_591);
and U118 (N_118,In_544,In_151);
and U119 (N_119,In_452,In_534);
nor U120 (N_120,In_221,In_196);
or U121 (N_121,In_176,In_365);
nor U122 (N_122,In_508,In_664);
or U123 (N_123,In_42,In_181);
nor U124 (N_124,In_313,In_63);
or U125 (N_125,In_501,In_683);
and U126 (N_126,In_256,In_616);
nand U127 (N_127,In_644,In_356);
nor U128 (N_128,In_453,In_473);
nor U129 (N_129,In_257,In_241);
nor U130 (N_130,In_535,In_333);
nand U131 (N_131,In_533,In_40);
nand U132 (N_132,In_139,In_668);
and U133 (N_133,In_524,In_526);
nand U134 (N_134,In_706,In_27);
and U135 (N_135,In_692,In_127);
nor U136 (N_136,In_178,In_335);
and U137 (N_137,In_475,In_680);
nand U138 (N_138,In_675,In_634);
and U139 (N_139,In_565,In_441);
and U140 (N_140,In_374,In_592);
nand U141 (N_141,In_216,In_495);
nand U142 (N_142,In_749,In_658);
nand U143 (N_143,In_625,In_19);
nand U144 (N_144,In_481,In_466);
and U145 (N_145,In_721,In_741);
nor U146 (N_146,In_714,In_480);
nand U147 (N_147,In_722,In_394);
or U148 (N_148,In_249,In_20);
and U149 (N_149,In_503,In_469);
nand U150 (N_150,In_204,In_697);
nand U151 (N_151,In_618,In_34);
nand U152 (N_152,In_129,In_252);
nand U153 (N_153,In_377,In_550);
xor U154 (N_154,In_647,In_558);
nor U155 (N_155,In_354,In_499);
nand U156 (N_156,In_361,In_425);
nor U157 (N_157,In_303,In_576);
nor U158 (N_158,In_153,In_532);
nand U159 (N_159,In_198,In_310);
or U160 (N_160,In_472,In_78);
nor U161 (N_161,In_275,In_720);
nand U162 (N_162,In_651,In_498);
or U163 (N_163,In_91,In_397);
nand U164 (N_164,In_58,In_271);
and U165 (N_165,In_142,In_6);
or U166 (N_166,In_403,In_727);
and U167 (N_167,In_376,In_134);
nand U168 (N_168,In_717,In_557);
nor U169 (N_169,In_510,In_23);
or U170 (N_170,In_222,In_156);
and U171 (N_171,In_506,In_578);
nor U172 (N_172,In_384,In_145);
and U173 (N_173,In_575,In_746);
and U174 (N_174,In_286,In_245);
nand U175 (N_175,In_15,In_386);
and U176 (N_176,In_61,In_615);
nor U177 (N_177,In_92,In_543);
or U178 (N_178,In_318,In_223);
and U179 (N_179,In_334,In_183);
or U180 (N_180,In_179,In_604);
nor U181 (N_181,In_126,In_390);
or U182 (N_182,In_637,In_231);
nand U183 (N_183,In_232,In_600);
or U184 (N_184,In_117,In_653);
nor U185 (N_185,In_416,In_633);
or U186 (N_186,In_360,In_489);
nand U187 (N_187,In_1,In_317);
and U188 (N_188,In_695,In_69);
nand U189 (N_189,In_17,In_331);
or U190 (N_190,In_612,In_277);
or U191 (N_191,In_273,In_13);
and U192 (N_192,In_307,In_342);
nor U193 (N_193,In_113,In_696);
and U194 (N_194,In_121,In_468);
nand U195 (N_195,In_345,In_288);
nor U196 (N_196,In_554,In_287);
and U197 (N_197,In_617,In_5);
and U198 (N_198,In_716,In_414);
or U199 (N_199,In_643,In_410);
and U200 (N_200,In_507,In_709);
nand U201 (N_201,In_654,In_338);
or U202 (N_202,In_398,In_240);
nor U203 (N_203,In_505,In_283);
nand U204 (N_204,In_364,In_629);
or U205 (N_205,In_210,In_385);
nand U206 (N_206,In_711,In_109);
nor U207 (N_207,In_419,In_269);
and U208 (N_208,In_411,In_75);
or U209 (N_209,In_649,In_47);
or U210 (N_210,In_341,In_159);
nand U211 (N_211,In_295,In_666);
and U212 (N_212,In_407,In_171);
nor U213 (N_213,In_214,In_89);
nor U214 (N_214,In_73,In_96);
and U215 (N_215,In_80,In_672);
or U216 (N_216,In_168,In_191);
nor U217 (N_217,In_259,In_574);
and U218 (N_218,In_517,In_470);
nor U219 (N_219,In_719,In_132);
nor U220 (N_220,In_326,In_230);
or U221 (N_221,In_487,In_438);
and U222 (N_222,In_366,In_314);
or U223 (N_223,In_457,In_212);
and U224 (N_224,In_165,In_648);
nor U225 (N_225,In_104,In_200);
nand U226 (N_226,In_137,In_486);
or U227 (N_227,In_246,In_547);
or U228 (N_228,In_68,In_494);
nand U229 (N_229,In_327,In_562);
nor U230 (N_230,In_389,In_436);
and U231 (N_231,In_270,In_442);
or U232 (N_232,In_671,In_255);
nor U233 (N_233,In_528,In_559);
nor U234 (N_234,In_67,In_146);
nand U235 (N_235,In_602,In_461);
or U236 (N_236,In_154,In_599);
nand U237 (N_237,In_440,In_49);
or U238 (N_238,In_710,In_371);
or U239 (N_239,In_678,In_110);
or U240 (N_240,In_747,In_704);
nand U241 (N_241,In_237,In_570);
and U242 (N_242,In_690,In_152);
nor U243 (N_243,In_149,In_707);
nor U244 (N_244,In_742,In_635);
or U245 (N_245,In_445,In_735);
or U246 (N_246,In_729,In_698);
nor U247 (N_247,In_622,In_140);
nor U248 (N_248,In_406,In_641);
nand U249 (N_249,In_540,In_568);
and U250 (N_250,In_290,In_102);
or U251 (N_251,In_343,In_467);
nor U252 (N_252,In_582,In_479);
xnor U253 (N_253,In_236,In_593);
nor U254 (N_254,In_546,In_82);
and U255 (N_255,In_567,In_462);
or U256 (N_256,In_55,In_164);
or U257 (N_257,In_521,In_426);
nand U258 (N_258,In_174,In_45);
nor U259 (N_259,In_566,In_131);
nand U260 (N_260,In_631,In_347);
nor U261 (N_261,In_141,In_300);
nand U262 (N_262,In_450,In_627);
or U263 (N_263,In_88,In_21);
nand U264 (N_264,In_569,In_265);
and U265 (N_265,In_375,In_428);
nand U266 (N_266,In_728,In_294);
nand U267 (N_267,In_542,In_148);
nor U268 (N_268,In_511,In_218);
and U269 (N_269,In_301,In_476);
or U270 (N_270,In_731,In_24);
and U271 (N_271,In_284,In_656);
or U272 (N_272,In_530,In_330);
or U273 (N_273,In_485,In_224);
and U274 (N_274,In_163,In_56);
or U275 (N_275,In_32,In_190);
and U276 (N_276,In_737,In_59);
nor U277 (N_277,In_496,In_267);
nor U278 (N_278,In_266,In_429);
or U279 (N_279,In_522,In_417);
nand U280 (N_280,In_325,In_421);
or U281 (N_281,In_10,In_595);
or U282 (N_282,In_46,In_681);
nand U283 (N_283,In_703,In_329);
and U284 (N_284,In_298,In_304);
nor U285 (N_285,In_217,In_64);
nor U286 (N_286,In_381,In_353);
or U287 (N_287,In_745,In_700);
or U288 (N_288,In_83,In_368);
nand U289 (N_289,In_609,In_435);
or U290 (N_290,In_541,In_483);
and U291 (N_291,In_587,In_563);
nand U292 (N_292,In_103,In_213);
and U293 (N_293,In_701,In_718);
nor U294 (N_294,In_346,In_588);
and U295 (N_295,In_580,In_420);
or U296 (N_296,In_409,In_733);
or U297 (N_297,In_607,In_693);
and U298 (N_298,In_93,In_520);
and U299 (N_299,In_564,In_344);
nand U300 (N_300,In_220,In_292);
or U301 (N_301,In_691,In_471);
and U302 (N_302,In_399,In_705);
nor U303 (N_303,In_537,In_193);
or U304 (N_304,In_28,In_373);
and U305 (N_305,In_72,In_518);
nor U306 (N_306,In_369,In_4);
nor U307 (N_307,In_254,In_596);
and U308 (N_308,In_205,In_251);
and U309 (N_309,In_16,In_133);
or U310 (N_310,In_357,In_715);
or U311 (N_311,In_227,In_478);
nor U312 (N_312,In_732,In_119);
and U313 (N_313,In_515,In_123);
and U314 (N_314,In_415,In_99);
xor U315 (N_315,In_423,In_182);
nor U316 (N_316,In_105,In_395);
nor U317 (N_317,In_226,In_652);
nor U318 (N_318,In_264,In_548);
nand U319 (N_319,In_157,In_689);
and U320 (N_320,In_100,In_279);
nand U321 (N_321,In_556,In_340);
nor U322 (N_322,In_233,In_572);
and U323 (N_323,In_22,In_50);
nand U324 (N_324,In_388,In_160);
and U325 (N_325,In_253,In_589);
nand U326 (N_326,In_124,In_669);
or U327 (N_327,In_454,In_594);
nor U328 (N_328,In_202,In_432);
nor U329 (N_329,In_180,In_586);
or U330 (N_330,In_736,In_623);
nor U331 (N_331,In_482,In_38);
nand U332 (N_332,In_41,In_439);
and U333 (N_333,In_400,In_504);
nand U334 (N_334,In_289,In_523);
nand U335 (N_335,In_65,In_76);
nand U336 (N_336,In_492,In_321);
xnor U337 (N_337,In_640,In_162);
nor U338 (N_338,In_585,In_54);
nor U339 (N_339,In_122,In_2);
nor U340 (N_340,In_446,In_642);
and U341 (N_341,In_62,In_33);
or U342 (N_342,In_95,In_312);
nor U343 (N_343,In_161,In_98);
or U344 (N_344,In_665,In_459);
nand U345 (N_345,In_738,In_247);
or U346 (N_346,In_262,In_77);
or U347 (N_347,In_30,In_687);
and U348 (N_348,In_513,In_324);
and U349 (N_349,In_456,In_502);
nor U350 (N_350,In_3,In_512);
or U351 (N_351,In_14,In_382);
nor U352 (N_352,In_405,In_620);
or U353 (N_353,In_211,In_192);
or U354 (N_354,In_302,In_730);
and U355 (N_355,In_9,In_118);
or U356 (N_356,In_186,In_743);
nor U357 (N_357,In_355,In_463);
and U358 (N_358,In_130,In_514);
nand U359 (N_359,In_688,In_74);
and U360 (N_360,In_610,In_336);
nor U361 (N_361,In_235,In_94);
nor U362 (N_362,In_25,In_413);
and U363 (N_363,In_260,In_488);
and U364 (N_364,In_234,In_387);
nand U365 (N_365,In_228,In_619);
and U366 (N_366,In_12,In_682);
or U367 (N_367,In_396,In_348);
and U368 (N_368,In_539,In_332);
nor U369 (N_369,In_734,In_372);
nor U370 (N_370,In_243,In_443);
nand U371 (N_371,In_184,In_52);
nor U372 (N_372,In_636,In_111);
and U373 (N_373,In_590,In_447);
and U374 (N_374,In_674,In_500);
nor U375 (N_375,In_433,In_135);
and U376 (N_376,In_117,In_706);
or U377 (N_377,In_275,In_386);
or U378 (N_378,In_367,In_466);
nor U379 (N_379,In_407,In_488);
nand U380 (N_380,In_86,In_401);
or U381 (N_381,In_652,In_377);
nand U382 (N_382,In_394,In_450);
and U383 (N_383,In_697,In_303);
nor U384 (N_384,In_674,In_394);
and U385 (N_385,In_677,In_157);
or U386 (N_386,In_403,In_651);
nand U387 (N_387,In_346,In_673);
nor U388 (N_388,In_117,In_319);
nor U389 (N_389,In_654,In_603);
nor U390 (N_390,In_459,In_733);
or U391 (N_391,In_678,In_470);
nor U392 (N_392,In_565,In_155);
nor U393 (N_393,In_527,In_461);
or U394 (N_394,In_250,In_48);
and U395 (N_395,In_427,In_476);
nand U396 (N_396,In_434,In_113);
or U397 (N_397,In_604,In_251);
and U398 (N_398,In_286,In_425);
and U399 (N_399,In_424,In_299);
nor U400 (N_400,In_432,In_252);
and U401 (N_401,In_340,In_527);
or U402 (N_402,In_659,In_619);
and U403 (N_403,In_200,In_269);
nand U404 (N_404,In_59,In_485);
nor U405 (N_405,In_395,In_719);
nor U406 (N_406,In_702,In_733);
nand U407 (N_407,In_329,In_262);
nor U408 (N_408,In_544,In_33);
and U409 (N_409,In_209,In_236);
nor U410 (N_410,In_198,In_722);
or U411 (N_411,In_176,In_71);
nor U412 (N_412,In_497,In_233);
nor U413 (N_413,In_267,In_650);
nor U414 (N_414,In_558,In_626);
xnor U415 (N_415,In_6,In_45);
and U416 (N_416,In_485,In_725);
or U417 (N_417,In_57,In_546);
nand U418 (N_418,In_609,In_16);
xor U419 (N_419,In_498,In_315);
or U420 (N_420,In_13,In_163);
nor U421 (N_421,In_477,In_83);
or U422 (N_422,In_246,In_244);
nor U423 (N_423,In_335,In_560);
and U424 (N_424,In_477,In_452);
nand U425 (N_425,In_149,In_559);
or U426 (N_426,In_395,In_275);
nor U427 (N_427,In_643,In_283);
nand U428 (N_428,In_232,In_291);
nand U429 (N_429,In_597,In_351);
nand U430 (N_430,In_423,In_111);
or U431 (N_431,In_54,In_624);
and U432 (N_432,In_741,In_317);
nand U433 (N_433,In_479,In_153);
or U434 (N_434,In_586,In_164);
nand U435 (N_435,In_316,In_687);
and U436 (N_436,In_159,In_16);
or U437 (N_437,In_354,In_168);
nand U438 (N_438,In_332,In_143);
nor U439 (N_439,In_360,In_8);
nand U440 (N_440,In_354,In_276);
and U441 (N_441,In_572,In_435);
nand U442 (N_442,In_431,In_356);
or U443 (N_443,In_2,In_259);
nand U444 (N_444,In_136,In_411);
and U445 (N_445,In_274,In_169);
and U446 (N_446,In_154,In_679);
nand U447 (N_447,In_720,In_381);
nand U448 (N_448,In_153,In_81);
and U449 (N_449,In_563,In_477);
and U450 (N_450,In_651,In_642);
or U451 (N_451,In_308,In_566);
and U452 (N_452,In_8,In_309);
and U453 (N_453,In_389,In_581);
nand U454 (N_454,In_366,In_0);
or U455 (N_455,In_628,In_250);
nor U456 (N_456,In_372,In_217);
nor U457 (N_457,In_121,In_651);
or U458 (N_458,In_352,In_510);
or U459 (N_459,In_265,In_313);
and U460 (N_460,In_128,In_588);
nand U461 (N_461,In_348,In_361);
nand U462 (N_462,In_62,In_328);
nor U463 (N_463,In_158,In_399);
nand U464 (N_464,In_539,In_709);
nand U465 (N_465,In_86,In_205);
and U466 (N_466,In_348,In_295);
nand U467 (N_467,In_412,In_702);
and U468 (N_468,In_408,In_178);
nand U469 (N_469,In_44,In_389);
nand U470 (N_470,In_200,In_244);
nor U471 (N_471,In_732,In_590);
and U472 (N_472,In_26,In_561);
xnor U473 (N_473,In_61,In_688);
or U474 (N_474,In_29,In_545);
nor U475 (N_475,In_646,In_735);
nor U476 (N_476,In_211,In_709);
or U477 (N_477,In_357,In_167);
nand U478 (N_478,In_110,In_368);
or U479 (N_479,In_77,In_654);
nor U480 (N_480,In_121,In_23);
and U481 (N_481,In_374,In_364);
nand U482 (N_482,In_186,In_448);
nand U483 (N_483,In_513,In_625);
nand U484 (N_484,In_183,In_748);
and U485 (N_485,In_270,In_154);
and U486 (N_486,In_559,In_696);
nor U487 (N_487,In_249,In_27);
nand U488 (N_488,In_610,In_506);
xor U489 (N_489,In_180,In_219);
and U490 (N_490,In_72,In_665);
nor U491 (N_491,In_670,In_547);
or U492 (N_492,In_572,In_175);
and U493 (N_493,In_680,In_284);
nor U494 (N_494,In_243,In_107);
nand U495 (N_495,In_41,In_414);
or U496 (N_496,In_83,In_259);
nand U497 (N_497,In_738,In_151);
and U498 (N_498,In_748,In_349);
nor U499 (N_499,In_278,In_386);
and U500 (N_500,In_137,In_731);
nor U501 (N_501,In_560,In_374);
or U502 (N_502,In_7,In_116);
nor U503 (N_503,In_532,In_229);
nor U504 (N_504,In_664,In_457);
nor U505 (N_505,In_603,In_2);
or U506 (N_506,In_393,In_41);
and U507 (N_507,In_467,In_135);
or U508 (N_508,In_406,In_378);
or U509 (N_509,In_333,In_690);
or U510 (N_510,In_626,In_634);
or U511 (N_511,In_522,In_41);
nor U512 (N_512,In_368,In_2);
nor U513 (N_513,In_284,In_410);
nor U514 (N_514,In_413,In_470);
and U515 (N_515,In_74,In_497);
nand U516 (N_516,In_364,In_691);
nand U517 (N_517,In_91,In_684);
and U518 (N_518,In_718,In_406);
or U519 (N_519,In_649,In_501);
and U520 (N_520,In_60,In_486);
nor U521 (N_521,In_337,In_51);
nor U522 (N_522,In_391,In_282);
or U523 (N_523,In_321,In_202);
nand U524 (N_524,In_538,In_319);
nand U525 (N_525,In_463,In_346);
or U526 (N_526,In_345,In_210);
nor U527 (N_527,In_418,In_359);
nor U528 (N_528,In_365,In_656);
or U529 (N_529,In_580,In_720);
and U530 (N_530,In_212,In_489);
and U531 (N_531,In_204,In_642);
nor U532 (N_532,In_446,In_349);
or U533 (N_533,In_600,In_527);
nor U534 (N_534,In_406,In_627);
or U535 (N_535,In_730,In_631);
and U536 (N_536,In_538,In_81);
or U537 (N_537,In_20,In_521);
or U538 (N_538,In_567,In_218);
and U539 (N_539,In_553,In_190);
or U540 (N_540,In_254,In_240);
or U541 (N_541,In_539,In_50);
and U542 (N_542,In_379,In_234);
nor U543 (N_543,In_604,In_737);
or U544 (N_544,In_458,In_218);
nand U545 (N_545,In_84,In_599);
and U546 (N_546,In_356,In_649);
nor U547 (N_547,In_121,In_228);
and U548 (N_548,In_477,In_58);
nand U549 (N_549,In_295,In_219);
or U550 (N_550,In_375,In_102);
or U551 (N_551,In_53,In_317);
or U552 (N_552,In_72,In_292);
nand U553 (N_553,In_544,In_71);
nor U554 (N_554,In_309,In_19);
nor U555 (N_555,In_706,In_452);
or U556 (N_556,In_679,In_722);
or U557 (N_557,In_46,In_605);
or U558 (N_558,In_257,In_670);
and U559 (N_559,In_480,In_28);
nand U560 (N_560,In_91,In_568);
nor U561 (N_561,In_230,In_258);
or U562 (N_562,In_162,In_728);
nor U563 (N_563,In_619,In_686);
nor U564 (N_564,In_301,In_490);
nand U565 (N_565,In_190,In_499);
and U566 (N_566,In_499,In_708);
nand U567 (N_567,In_642,In_621);
and U568 (N_568,In_304,In_278);
nor U569 (N_569,In_264,In_14);
or U570 (N_570,In_144,In_551);
and U571 (N_571,In_703,In_88);
and U572 (N_572,In_58,In_724);
or U573 (N_573,In_410,In_644);
nor U574 (N_574,In_173,In_406);
nor U575 (N_575,In_369,In_158);
and U576 (N_576,In_162,In_638);
nor U577 (N_577,In_78,In_608);
xor U578 (N_578,In_675,In_641);
nor U579 (N_579,In_448,In_595);
or U580 (N_580,In_446,In_616);
nor U581 (N_581,In_310,In_373);
and U582 (N_582,In_355,In_559);
and U583 (N_583,In_295,In_367);
or U584 (N_584,In_415,In_35);
nor U585 (N_585,In_171,In_523);
nand U586 (N_586,In_372,In_635);
and U587 (N_587,In_614,In_414);
nor U588 (N_588,In_598,In_439);
and U589 (N_589,In_261,In_92);
or U590 (N_590,In_454,In_690);
nand U591 (N_591,In_315,In_622);
or U592 (N_592,In_559,In_315);
nor U593 (N_593,In_651,In_553);
nor U594 (N_594,In_577,In_331);
or U595 (N_595,In_74,In_451);
or U596 (N_596,In_699,In_320);
and U597 (N_597,In_92,In_707);
nand U598 (N_598,In_616,In_300);
and U599 (N_599,In_244,In_510);
nand U600 (N_600,In_453,In_702);
nor U601 (N_601,In_47,In_644);
or U602 (N_602,In_61,In_438);
nor U603 (N_603,In_398,In_630);
nand U604 (N_604,In_490,In_324);
nand U605 (N_605,In_671,In_82);
nand U606 (N_606,In_104,In_155);
or U607 (N_607,In_652,In_685);
and U608 (N_608,In_156,In_720);
or U609 (N_609,In_43,In_423);
and U610 (N_610,In_8,In_317);
nand U611 (N_611,In_229,In_22);
nand U612 (N_612,In_634,In_515);
nand U613 (N_613,In_58,In_530);
nor U614 (N_614,In_642,In_21);
or U615 (N_615,In_48,In_146);
nand U616 (N_616,In_185,In_623);
and U617 (N_617,In_205,In_206);
or U618 (N_618,In_379,In_396);
and U619 (N_619,In_307,In_289);
nor U620 (N_620,In_634,In_123);
or U621 (N_621,In_72,In_67);
nand U622 (N_622,In_478,In_114);
nor U623 (N_623,In_686,In_252);
or U624 (N_624,In_714,In_345);
and U625 (N_625,In_447,In_83);
nor U626 (N_626,In_314,In_575);
nand U627 (N_627,In_55,In_277);
and U628 (N_628,In_338,In_238);
nand U629 (N_629,In_126,In_72);
or U630 (N_630,In_228,In_744);
nor U631 (N_631,In_644,In_695);
nand U632 (N_632,In_639,In_631);
nor U633 (N_633,In_628,In_472);
nand U634 (N_634,In_328,In_576);
or U635 (N_635,In_172,In_134);
and U636 (N_636,In_674,In_596);
and U637 (N_637,In_728,In_564);
nor U638 (N_638,In_85,In_88);
nand U639 (N_639,In_320,In_555);
nand U640 (N_640,In_383,In_347);
and U641 (N_641,In_486,In_502);
and U642 (N_642,In_230,In_69);
and U643 (N_643,In_71,In_733);
or U644 (N_644,In_459,In_698);
or U645 (N_645,In_202,In_418);
or U646 (N_646,In_7,In_746);
nand U647 (N_647,In_694,In_736);
nand U648 (N_648,In_99,In_228);
or U649 (N_649,In_42,In_444);
nor U650 (N_650,In_696,In_638);
nor U651 (N_651,In_468,In_718);
and U652 (N_652,In_95,In_581);
or U653 (N_653,In_597,In_205);
nor U654 (N_654,In_440,In_29);
and U655 (N_655,In_108,In_577);
nor U656 (N_656,In_647,In_148);
xor U657 (N_657,In_40,In_631);
nand U658 (N_658,In_157,In_691);
and U659 (N_659,In_156,In_639);
or U660 (N_660,In_185,In_563);
and U661 (N_661,In_122,In_681);
or U662 (N_662,In_98,In_154);
nand U663 (N_663,In_211,In_528);
nor U664 (N_664,In_742,In_368);
or U665 (N_665,In_59,In_641);
or U666 (N_666,In_456,In_297);
nor U667 (N_667,In_461,In_648);
or U668 (N_668,In_624,In_301);
and U669 (N_669,In_365,In_282);
nand U670 (N_670,In_586,In_543);
and U671 (N_671,In_149,In_736);
or U672 (N_672,In_403,In_99);
or U673 (N_673,In_135,In_516);
or U674 (N_674,In_725,In_446);
and U675 (N_675,In_421,In_712);
nand U676 (N_676,In_655,In_182);
and U677 (N_677,In_585,In_656);
or U678 (N_678,In_648,In_670);
nor U679 (N_679,In_388,In_397);
nor U680 (N_680,In_421,In_244);
nand U681 (N_681,In_490,In_283);
or U682 (N_682,In_358,In_25);
nand U683 (N_683,In_472,In_35);
or U684 (N_684,In_258,In_440);
and U685 (N_685,In_102,In_431);
or U686 (N_686,In_733,In_254);
or U687 (N_687,In_423,In_297);
or U688 (N_688,In_87,In_85);
nor U689 (N_689,In_166,In_718);
and U690 (N_690,In_447,In_537);
nor U691 (N_691,In_606,In_276);
or U692 (N_692,In_201,In_4);
nor U693 (N_693,In_206,In_65);
nor U694 (N_694,In_674,In_460);
nand U695 (N_695,In_427,In_175);
nor U696 (N_696,In_683,In_434);
or U697 (N_697,In_349,In_332);
or U698 (N_698,In_347,In_93);
nand U699 (N_699,In_225,In_42);
and U700 (N_700,In_499,In_439);
nand U701 (N_701,In_643,In_359);
nand U702 (N_702,In_516,In_553);
or U703 (N_703,In_133,In_66);
and U704 (N_704,In_438,In_265);
nor U705 (N_705,In_410,In_337);
nor U706 (N_706,In_41,In_202);
or U707 (N_707,In_293,In_632);
or U708 (N_708,In_630,In_680);
and U709 (N_709,In_265,In_329);
nand U710 (N_710,In_478,In_562);
nand U711 (N_711,In_57,In_134);
and U712 (N_712,In_293,In_117);
and U713 (N_713,In_92,In_357);
and U714 (N_714,In_420,In_455);
and U715 (N_715,In_584,In_511);
nand U716 (N_716,In_372,In_205);
nor U717 (N_717,In_597,In_209);
or U718 (N_718,In_525,In_47);
nand U719 (N_719,In_234,In_633);
or U720 (N_720,In_577,In_524);
nor U721 (N_721,In_721,In_243);
or U722 (N_722,In_430,In_736);
and U723 (N_723,In_31,In_257);
and U724 (N_724,In_85,In_439);
and U725 (N_725,In_344,In_29);
and U726 (N_726,In_217,In_357);
nor U727 (N_727,In_66,In_7);
and U728 (N_728,In_330,In_671);
and U729 (N_729,In_195,In_533);
nand U730 (N_730,In_78,In_584);
or U731 (N_731,In_172,In_706);
and U732 (N_732,In_187,In_230);
nand U733 (N_733,In_230,In_99);
or U734 (N_734,In_490,In_645);
and U735 (N_735,In_84,In_1);
nor U736 (N_736,In_270,In_559);
nor U737 (N_737,In_732,In_730);
or U738 (N_738,In_548,In_585);
or U739 (N_739,In_488,In_147);
or U740 (N_740,In_114,In_646);
nand U741 (N_741,In_505,In_569);
or U742 (N_742,In_524,In_306);
or U743 (N_743,In_387,In_78);
nor U744 (N_744,In_64,In_284);
or U745 (N_745,In_595,In_601);
xnor U746 (N_746,In_255,In_446);
nand U747 (N_747,In_335,In_448);
nor U748 (N_748,In_397,In_699);
nor U749 (N_749,In_274,In_99);
and U750 (N_750,In_291,In_243);
nor U751 (N_751,In_323,In_512);
nor U752 (N_752,In_711,In_624);
and U753 (N_753,In_229,In_344);
nand U754 (N_754,In_222,In_296);
and U755 (N_755,In_137,In_208);
and U756 (N_756,In_593,In_250);
nor U757 (N_757,In_129,In_415);
nand U758 (N_758,In_632,In_703);
nor U759 (N_759,In_272,In_623);
and U760 (N_760,In_630,In_556);
or U761 (N_761,In_202,In_244);
or U762 (N_762,In_455,In_230);
nor U763 (N_763,In_687,In_735);
nor U764 (N_764,In_596,In_458);
or U765 (N_765,In_76,In_152);
and U766 (N_766,In_668,In_14);
and U767 (N_767,In_532,In_681);
nor U768 (N_768,In_186,In_744);
nor U769 (N_769,In_299,In_40);
nor U770 (N_770,In_555,In_545);
or U771 (N_771,In_484,In_399);
and U772 (N_772,In_605,In_357);
and U773 (N_773,In_586,In_401);
or U774 (N_774,In_658,In_253);
or U775 (N_775,In_668,In_404);
nor U776 (N_776,In_118,In_412);
or U777 (N_777,In_9,In_406);
and U778 (N_778,In_127,In_437);
or U779 (N_779,In_201,In_734);
or U780 (N_780,In_11,In_91);
and U781 (N_781,In_457,In_115);
or U782 (N_782,In_543,In_69);
and U783 (N_783,In_126,In_516);
nor U784 (N_784,In_206,In_259);
nand U785 (N_785,In_112,In_175);
and U786 (N_786,In_643,In_352);
nand U787 (N_787,In_645,In_206);
nand U788 (N_788,In_333,In_488);
nor U789 (N_789,In_135,In_325);
or U790 (N_790,In_131,In_390);
and U791 (N_791,In_328,In_372);
and U792 (N_792,In_418,In_345);
and U793 (N_793,In_678,In_159);
or U794 (N_794,In_628,In_515);
or U795 (N_795,In_524,In_276);
nor U796 (N_796,In_236,In_99);
nor U797 (N_797,In_654,In_156);
and U798 (N_798,In_601,In_20);
nand U799 (N_799,In_673,In_544);
nor U800 (N_800,In_290,In_142);
nor U801 (N_801,In_8,In_254);
nand U802 (N_802,In_489,In_475);
nor U803 (N_803,In_148,In_491);
or U804 (N_804,In_693,In_272);
or U805 (N_805,In_221,In_219);
nand U806 (N_806,In_85,In_258);
nand U807 (N_807,In_709,In_688);
or U808 (N_808,In_613,In_77);
or U809 (N_809,In_699,In_630);
or U810 (N_810,In_352,In_219);
or U811 (N_811,In_125,In_200);
and U812 (N_812,In_679,In_504);
nand U813 (N_813,In_670,In_490);
and U814 (N_814,In_625,In_709);
and U815 (N_815,In_477,In_157);
and U816 (N_816,In_303,In_228);
nor U817 (N_817,In_48,In_401);
or U818 (N_818,In_142,In_522);
or U819 (N_819,In_705,In_165);
nor U820 (N_820,In_516,In_390);
nand U821 (N_821,In_402,In_67);
nand U822 (N_822,In_652,In_128);
nand U823 (N_823,In_661,In_171);
and U824 (N_824,In_152,In_151);
and U825 (N_825,In_454,In_715);
nand U826 (N_826,In_154,In_73);
nand U827 (N_827,In_724,In_651);
and U828 (N_828,In_526,In_558);
and U829 (N_829,In_105,In_211);
nor U830 (N_830,In_647,In_408);
nand U831 (N_831,In_56,In_427);
nor U832 (N_832,In_219,In_99);
nand U833 (N_833,In_301,In_538);
nor U834 (N_834,In_638,In_734);
nand U835 (N_835,In_576,In_477);
and U836 (N_836,In_487,In_356);
nor U837 (N_837,In_329,In_159);
or U838 (N_838,In_578,In_432);
or U839 (N_839,In_445,In_195);
or U840 (N_840,In_18,In_398);
nand U841 (N_841,In_629,In_407);
and U842 (N_842,In_264,In_566);
nor U843 (N_843,In_116,In_691);
and U844 (N_844,In_99,In_683);
and U845 (N_845,In_695,In_512);
nand U846 (N_846,In_301,In_452);
nand U847 (N_847,In_193,In_335);
nor U848 (N_848,In_731,In_53);
or U849 (N_849,In_91,In_199);
and U850 (N_850,In_219,In_21);
or U851 (N_851,In_749,In_57);
nand U852 (N_852,In_322,In_694);
nor U853 (N_853,In_652,In_186);
or U854 (N_854,In_657,In_65);
and U855 (N_855,In_741,In_354);
or U856 (N_856,In_43,In_457);
and U857 (N_857,In_370,In_79);
nor U858 (N_858,In_620,In_567);
nor U859 (N_859,In_572,In_465);
nand U860 (N_860,In_602,In_586);
or U861 (N_861,In_360,In_463);
and U862 (N_862,In_235,In_229);
and U863 (N_863,In_674,In_437);
nor U864 (N_864,In_56,In_109);
nand U865 (N_865,In_613,In_363);
nand U866 (N_866,In_288,In_146);
nand U867 (N_867,In_14,In_20);
xor U868 (N_868,In_241,In_498);
nand U869 (N_869,In_726,In_521);
nand U870 (N_870,In_659,In_407);
and U871 (N_871,In_267,In_704);
or U872 (N_872,In_439,In_535);
and U873 (N_873,In_718,In_636);
nor U874 (N_874,In_568,In_195);
and U875 (N_875,In_54,In_337);
nor U876 (N_876,In_184,In_570);
xnor U877 (N_877,In_459,In_455);
nor U878 (N_878,In_305,In_142);
nand U879 (N_879,In_88,In_112);
and U880 (N_880,In_713,In_380);
nand U881 (N_881,In_428,In_611);
or U882 (N_882,In_555,In_413);
or U883 (N_883,In_416,In_84);
and U884 (N_884,In_12,In_559);
or U885 (N_885,In_441,In_517);
nand U886 (N_886,In_303,In_632);
nand U887 (N_887,In_437,In_279);
nand U888 (N_888,In_681,In_593);
and U889 (N_889,In_651,In_720);
nand U890 (N_890,In_595,In_165);
nand U891 (N_891,In_319,In_599);
nor U892 (N_892,In_628,In_222);
nor U893 (N_893,In_191,In_351);
nand U894 (N_894,In_226,In_143);
or U895 (N_895,In_23,In_27);
nand U896 (N_896,In_419,In_73);
nand U897 (N_897,In_70,In_158);
and U898 (N_898,In_410,In_256);
xor U899 (N_899,In_331,In_429);
or U900 (N_900,In_167,In_282);
or U901 (N_901,In_134,In_521);
xor U902 (N_902,In_122,In_608);
and U903 (N_903,In_510,In_241);
nor U904 (N_904,In_548,In_295);
nor U905 (N_905,In_409,In_515);
and U906 (N_906,In_215,In_156);
or U907 (N_907,In_186,In_101);
nor U908 (N_908,In_142,In_109);
nor U909 (N_909,In_77,In_643);
or U910 (N_910,In_203,In_230);
nand U911 (N_911,In_452,In_155);
nor U912 (N_912,In_522,In_436);
nor U913 (N_913,In_738,In_608);
nor U914 (N_914,In_115,In_435);
nor U915 (N_915,In_537,In_657);
and U916 (N_916,In_241,In_369);
or U917 (N_917,In_731,In_291);
or U918 (N_918,In_311,In_180);
or U919 (N_919,In_727,In_523);
nand U920 (N_920,In_233,In_12);
and U921 (N_921,In_177,In_109);
and U922 (N_922,In_224,In_630);
or U923 (N_923,In_243,In_219);
nor U924 (N_924,In_625,In_65);
nor U925 (N_925,In_278,In_532);
or U926 (N_926,In_631,In_281);
nand U927 (N_927,In_460,In_424);
and U928 (N_928,In_308,In_228);
and U929 (N_929,In_168,In_525);
nor U930 (N_930,In_727,In_391);
and U931 (N_931,In_675,In_86);
or U932 (N_932,In_25,In_197);
and U933 (N_933,In_683,In_535);
nor U934 (N_934,In_636,In_414);
and U935 (N_935,In_53,In_600);
xor U936 (N_936,In_548,In_28);
and U937 (N_937,In_535,In_698);
and U938 (N_938,In_465,In_580);
nand U939 (N_939,In_319,In_435);
or U940 (N_940,In_133,In_155);
nand U941 (N_941,In_313,In_137);
and U942 (N_942,In_607,In_7);
nand U943 (N_943,In_261,In_422);
nand U944 (N_944,In_598,In_45);
nor U945 (N_945,In_269,In_607);
nand U946 (N_946,In_75,In_436);
or U947 (N_947,In_676,In_95);
nand U948 (N_948,In_246,In_452);
nand U949 (N_949,In_101,In_15);
nand U950 (N_950,In_137,In_129);
or U951 (N_951,In_538,In_110);
or U952 (N_952,In_49,In_458);
xor U953 (N_953,In_295,In_89);
and U954 (N_954,In_192,In_179);
nand U955 (N_955,In_321,In_505);
or U956 (N_956,In_181,In_618);
or U957 (N_957,In_391,In_604);
and U958 (N_958,In_511,In_294);
and U959 (N_959,In_329,In_558);
nor U960 (N_960,In_318,In_654);
nor U961 (N_961,In_649,In_555);
and U962 (N_962,In_502,In_663);
or U963 (N_963,In_100,In_668);
or U964 (N_964,In_140,In_333);
and U965 (N_965,In_356,In_502);
or U966 (N_966,In_394,In_5);
nand U967 (N_967,In_527,In_566);
and U968 (N_968,In_398,In_596);
nand U969 (N_969,In_380,In_506);
or U970 (N_970,In_320,In_156);
nand U971 (N_971,In_680,In_249);
or U972 (N_972,In_520,In_112);
xnor U973 (N_973,In_434,In_404);
and U974 (N_974,In_505,In_429);
nor U975 (N_975,In_479,In_426);
nand U976 (N_976,In_332,In_304);
nor U977 (N_977,In_740,In_588);
and U978 (N_978,In_272,In_294);
or U979 (N_979,In_246,In_303);
and U980 (N_980,In_44,In_197);
nor U981 (N_981,In_53,In_216);
and U982 (N_982,In_641,In_49);
or U983 (N_983,In_427,In_464);
or U984 (N_984,In_357,In_182);
and U985 (N_985,In_22,In_546);
nor U986 (N_986,In_283,In_634);
nand U987 (N_987,In_568,In_411);
nor U988 (N_988,In_527,In_155);
and U989 (N_989,In_286,In_162);
and U990 (N_990,In_704,In_9);
and U991 (N_991,In_74,In_695);
nor U992 (N_992,In_188,In_705);
or U993 (N_993,In_329,In_441);
or U994 (N_994,In_702,In_142);
nor U995 (N_995,In_419,In_67);
nor U996 (N_996,In_330,In_217);
and U997 (N_997,In_40,In_295);
nand U998 (N_998,In_717,In_85);
nand U999 (N_999,In_288,In_513);
or U1000 (N_1000,In_311,In_584);
or U1001 (N_1001,In_572,In_246);
and U1002 (N_1002,In_402,In_660);
or U1003 (N_1003,In_512,In_33);
nor U1004 (N_1004,In_172,In_235);
and U1005 (N_1005,In_105,In_263);
or U1006 (N_1006,In_226,In_539);
nor U1007 (N_1007,In_310,In_541);
or U1008 (N_1008,In_388,In_324);
nor U1009 (N_1009,In_171,In_453);
nand U1010 (N_1010,In_240,In_653);
nand U1011 (N_1011,In_589,In_157);
xnor U1012 (N_1012,In_616,In_9);
nand U1013 (N_1013,In_377,In_303);
or U1014 (N_1014,In_680,In_405);
and U1015 (N_1015,In_289,In_741);
nand U1016 (N_1016,In_748,In_440);
and U1017 (N_1017,In_410,In_506);
nor U1018 (N_1018,In_174,In_256);
and U1019 (N_1019,In_714,In_172);
and U1020 (N_1020,In_45,In_152);
and U1021 (N_1021,In_7,In_351);
xnor U1022 (N_1022,In_542,In_618);
nand U1023 (N_1023,In_11,In_102);
and U1024 (N_1024,In_641,In_93);
and U1025 (N_1025,In_344,In_158);
nor U1026 (N_1026,In_592,In_53);
nand U1027 (N_1027,In_304,In_135);
xor U1028 (N_1028,In_68,In_116);
and U1029 (N_1029,In_729,In_556);
nand U1030 (N_1030,In_521,In_352);
nand U1031 (N_1031,In_583,In_90);
and U1032 (N_1032,In_386,In_26);
nor U1033 (N_1033,In_92,In_286);
and U1034 (N_1034,In_440,In_378);
or U1035 (N_1035,In_214,In_188);
nand U1036 (N_1036,In_682,In_451);
and U1037 (N_1037,In_617,In_638);
or U1038 (N_1038,In_584,In_89);
nor U1039 (N_1039,In_282,In_464);
nor U1040 (N_1040,In_187,In_154);
nand U1041 (N_1041,In_258,In_27);
nand U1042 (N_1042,In_375,In_32);
and U1043 (N_1043,In_374,In_731);
and U1044 (N_1044,In_530,In_239);
or U1045 (N_1045,In_425,In_86);
or U1046 (N_1046,In_574,In_385);
nand U1047 (N_1047,In_143,In_717);
and U1048 (N_1048,In_114,In_128);
nor U1049 (N_1049,In_675,In_708);
and U1050 (N_1050,In_416,In_464);
or U1051 (N_1051,In_4,In_551);
and U1052 (N_1052,In_614,In_702);
nor U1053 (N_1053,In_215,In_605);
nand U1054 (N_1054,In_484,In_407);
and U1055 (N_1055,In_159,In_326);
and U1056 (N_1056,In_634,In_655);
nor U1057 (N_1057,In_395,In_517);
or U1058 (N_1058,In_42,In_678);
nand U1059 (N_1059,In_389,In_444);
nand U1060 (N_1060,In_158,In_88);
or U1061 (N_1061,In_649,In_25);
or U1062 (N_1062,In_466,In_680);
nand U1063 (N_1063,In_587,In_669);
nor U1064 (N_1064,In_636,In_562);
nor U1065 (N_1065,In_172,In_322);
nor U1066 (N_1066,In_573,In_177);
or U1067 (N_1067,In_703,In_312);
nor U1068 (N_1068,In_746,In_530);
nand U1069 (N_1069,In_613,In_492);
nor U1070 (N_1070,In_445,In_295);
and U1071 (N_1071,In_492,In_712);
or U1072 (N_1072,In_569,In_607);
nand U1073 (N_1073,In_584,In_714);
nor U1074 (N_1074,In_687,In_51);
nand U1075 (N_1075,In_88,In_199);
nor U1076 (N_1076,In_537,In_606);
nand U1077 (N_1077,In_236,In_147);
and U1078 (N_1078,In_626,In_228);
and U1079 (N_1079,In_89,In_489);
or U1080 (N_1080,In_212,In_631);
nor U1081 (N_1081,In_737,In_491);
or U1082 (N_1082,In_404,In_216);
and U1083 (N_1083,In_515,In_243);
nand U1084 (N_1084,In_411,In_497);
nand U1085 (N_1085,In_651,In_619);
or U1086 (N_1086,In_544,In_269);
nor U1087 (N_1087,In_303,In_332);
nor U1088 (N_1088,In_286,In_653);
nor U1089 (N_1089,In_460,In_715);
and U1090 (N_1090,In_643,In_575);
and U1091 (N_1091,In_310,In_731);
or U1092 (N_1092,In_399,In_295);
nor U1093 (N_1093,In_440,In_327);
and U1094 (N_1094,In_173,In_733);
nor U1095 (N_1095,In_350,In_589);
or U1096 (N_1096,In_380,In_149);
and U1097 (N_1097,In_166,In_62);
or U1098 (N_1098,In_668,In_51);
and U1099 (N_1099,In_169,In_46);
or U1100 (N_1100,In_76,In_264);
and U1101 (N_1101,In_486,In_624);
nor U1102 (N_1102,In_33,In_625);
or U1103 (N_1103,In_529,In_396);
nand U1104 (N_1104,In_219,In_14);
nor U1105 (N_1105,In_108,In_735);
and U1106 (N_1106,In_593,In_327);
or U1107 (N_1107,In_220,In_471);
or U1108 (N_1108,In_121,In_593);
and U1109 (N_1109,In_91,In_582);
or U1110 (N_1110,In_232,In_437);
nand U1111 (N_1111,In_532,In_101);
and U1112 (N_1112,In_372,In_281);
and U1113 (N_1113,In_735,In_307);
nand U1114 (N_1114,In_711,In_80);
and U1115 (N_1115,In_592,In_652);
and U1116 (N_1116,In_153,In_318);
and U1117 (N_1117,In_454,In_274);
or U1118 (N_1118,In_456,In_584);
xnor U1119 (N_1119,In_9,In_703);
nor U1120 (N_1120,In_349,In_607);
nand U1121 (N_1121,In_395,In_557);
and U1122 (N_1122,In_135,In_186);
or U1123 (N_1123,In_26,In_180);
nand U1124 (N_1124,In_484,In_247);
nor U1125 (N_1125,In_235,In_384);
or U1126 (N_1126,In_182,In_475);
and U1127 (N_1127,In_597,In_572);
and U1128 (N_1128,In_377,In_64);
nand U1129 (N_1129,In_354,In_616);
xnor U1130 (N_1130,In_690,In_254);
nor U1131 (N_1131,In_202,In_601);
or U1132 (N_1132,In_631,In_100);
and U1133 (N_1133,In_25,In_263);
or U1134 (N_1134,In_644,In_720);
nor U1135 (N_1135,In_707,In_666);
nor U1136 (N_1136,In_397,In_525);
and U1137 (N_1137,In_581,In_486);
nand U1138 (N_1138,In_274,In_308);
nand U1139 (N_1139,In_93,In_734);
nor U1140 (N_1140,In_357,In_589);
nor U1141 (N_1141,In_501,In_227);
and U1142 (N_1142,In_265,In_456);
nand U1143 (N_1143,In_440,In_504);
nor U1144 (N_1144,In_452,In_119);
or U1145 (N_1145,In_525,In_473);
or U1146 (N_1146,In_45,In_194);
nand U1147 (N_1147,In_122,In_214);
nor U1148 (N_1148,In_700,In_473);
or U1149 (N_1149,In_493,In_118);
or U1150 (N_1150,In_88,In_446);
nand U1151 (N_1151,In_121,In_36);
or U1152 (N_1152,In_191,In_249);
nor U1153 (N_1153,In_399,In_731);
and U1154 (N_1154,In_11,In_691);
or U1155 (N_1155,In_228,In_417);
nor U1156 (N_1156,In_54,In_451);
nor U1157 (N_1157,In_21,In_123);
or U1158 (N_1158,In_663,In_395);
nand U1159 (N_1159,In_457,In_101);
or U1160 (N_1160,In_548,In_684);
and U1161 (N_1161,In_460,In_707);
nor U1162 (N_1162,In_13,In_70);
and U1163 (N_1163,In_679,In_627);
nor U1164 (N_1164,In_397,In_148);
and U1165 (N_1165,In_189,In_315);
or U1166 (N_1166,In_84,In_646);
and U1167 (N_1167,In_148,In_124);
or U1168 (N_1168,In_746,In_561);
or U1169 (N_1169,In_364,In_158);
or U1170 (N_1170,In_575,In_106);
nand U1171 (N_1171,In_92,In_168);
and U1172 (N_1172,In_583,In_17);
nand U1173 (N_1173,In_440,In_544);
nor U1174 (N_1174,In_170,In_287);
nor U1175 (N_1175,In_217,In_239);
and U1176 (N_1176,In_82,In_419);
and U1177 (N_1177,In_525,In_613);
nor U1178 (N_1178,In_678,In_666);
nor U1179 (N_1179,In_250,In_402);
or U1180 (N_1180,In_529,In_186);
nor U1181 (N_1181,In_82,In_272);
nand U1182 (N_1182,In_212,In_362);
or U1183 (N_1183,In_36,In_242);
and U1184 (N_1184,In_145,In_665);
nor U1185 (N_1185,In_737,In_490);
or U1186 (N_1186,In_713,In_582);
and U1187 (N_1187,In_716,In_54);
or U1188 (N_1188,In_333,In_98);
or U1189 (N_1189,In_429,In_262);
or U1190 (N_1190,In_303,In_481);
nor U1191 (N_1191,In_501,In_518);
or U1192 (N_1192,In_184,In_60);
or U1193 (N_1193,In_393,In_149);
or U1194 (N_1194,In_118,In_23);
xor U1195 (N_1195,In_388,In_29);
or U1196 (N_1196,In_420,In_287);
or U1197 (N_1197,In_308,In_533);
nor U1198 (N_1198,In_666,In_470);
or U1199 (N_1199,In_288,In_119);
or U1200 (N_1200,In_361,In_168);
nor U1201 (N_1201,In_318,In_353);
or U1202 (N_1202,In_610,In_44);
and U1203 (N_1203,In_406,In_436);
nand U1204 (N_1204,In_207,In_250);
nand U1205 (N_1205,In_57,In_94);
or U1206 (N_1206,In_390,In_384);
and U1207 (N_1207,In_102,In_559);
nor U1208 (N_1208,In_73,In_244);
nor U1209 (N_1209,In_132,In_446);
nand U1210 (N_1210,In_614,In_472);
and U1211 (N_1211,In_80,In_375);
and U1212 (N_1212,In_550,In_502);
nand U1213 (N_1213,In_0,In_301);
nor U1214 (N_1214,In_582,In_611);
or U1215 (N_1215,In_735,In_536);
nor U1216 (N_1216,In_636,In_500);
or U1217 (N_1217,In_200,In_601);
nand U1218 (N_1218,In_631,In_699);
nand U1219 (N_1219,In_460,In_561);
or U1220 (N_1220,In_460,In_224);
or U1221 (N_1221,In_147,In_545);
nand U1222 (N_1222,In_430,In_221);
nand U1223 (N_1223,In_319,In_286);
nand U1224 (N_1224,In_554,In_341);
or U1225 (N_1225,In_714,In_154);
and U1226 (N_1226,In_209,In_223);
nor U1227 (N_1227,In_711,In_117);
or U1228 (N_1228,In_326,In_266);
or U1229 (N_1229,In_369,In_584);
or U1230 (N_1230,In_236,In_50);
or U1231 (N_1231,In_231,In_480);
and U1232 (N_1232,In_270,In_106);
nor U1233 (N_1233,In_400,In_219);
nand U1234 (N_1234,In_340,In_723);
nor U1235 (N_1235,In_572,In_580);
nor U1236 (N_1236,In_68,In_130);
or U1237 (N_1237,In_429,In_253);
xor U1238 (N_1238,In_141,In_15);
nand U1239 (N_1239,In_141,In_485);
nor U1240 (N_1240,In_503,In_638);
nand U1241 (N_1241,In_354,In_46);
and U1242 (N_1242,In_136,In_748);
nand U1243 (N_1243,In_393,In_445);
or U1244 (N_1244,In_11,In_634);
and U1245 (N_1245,In_192,In_465);
nand U1246 (N_1246,In_327,In_437);
nand U1247 (N_1247,In_10,In_422);
or U1248 (N_1248,In_166,In_648);
and U1249 (N_1249,In_648,In_203);
and U1250 (N_1250,In_561,In_450);
or U1251 (N_1251,In_60,In_621);
nand U1252 (N_1252,In_678,In_530);
nor U1253 (N_1253,In_210,In_275);
nor U1254 (N_1254,In_5,In_197);
nor U1255 (N_1255,In_281,In_288);
or U1256 (N_1256,In_423,In_463);
or U1257 (N_1257,In_543,In_231);
or U1258 (N_1258,In_145,In_474);
nand U1259 (N_1259,In_430,In_699);
nand U1260 (N_1260,In_45,In_98);
or U1261 (N_1261,In_451,In_45);
or U1262 (N_1262,In_658,In_156);
nand U1263 (N_1263,In_615,In_288);
nor U1264 (N_1264,In_697,In_146);
nand U1265 (N_1265,In_671,In_749);
and U1266 (N_1266,In_541,In_689);
nor U1267 (N_1267,In_585,In_325);
and U1268 (N_1268,In_179,In_18);
or U1269 (N_1269,In_744,In_481);
xor U1270 (N_1270,In_41,In_140);
or U1271 (N_1271,In_192,In_628);
nor U1272 (N_1272,In_165,In_179);
nand U1273 (N_1273,In_72,In_297);
and U1274 (N_1274,In_79,In_618);
nand U1275 (N_1275,In_135,In_499);
nand U1276 (N_1276,In_8,In_575);
and U1277 (N_1277,In_672,In_185);
and U1278 (N_1278,In_98,In_479);
nor U1279 (N_1279,In_294,In_570);
and U1280 (N_1280,In_643,In_134);
nor U1281 (N_1281,In_19,In_472);
and U1282 (N_1282,In_83,In_601);
nor U1283 (N_1283,In_425,In_435);
or U1284 (N_1284,In_564,In_617);
or U1285 (N_1285,In_345,In_148);
or U1286 (N_1286,In_659,In_577);
nand U1287 (N_1287,In_115,In_745);
nor U1288 (N_1288,In_171,In_71);
nand U1289 (N_1289,In_430,In_16);
or U1290 (N_1290,In_268,In_437);
nand U1291 (N_1291,In_178,In_305);
nor U1292 (N_1292,In_714,In_158);
nor U1293 (N_1293,In_70,In_143);
nand U1294 (N_1294,In_518,In_140);
and U1295 (N_1295,In_529,In_294);
nor U1296 (N_1296,In_695,In_387);
nand U1297 (N_1297,In_326,In_518);
and U1298 (N_1298,In_119,In_604);
nand U1299 (N_1299,In_505,In_257);
and U1300 (N_1300,In_196,In_669);
and U1301 (N_1301,In_708,In_617);
nor U1302 (N_1302,In_150,In_284);
and U1303 (N_1303,In_400,In_689);
or U1304 (N_1304,In_728,In_485);
nor U1305 (N_1305,In_57,In_214);
and U1306 (N_1306,In_42,In_71);
and U1307 (N_1307,In_593,In_318);
nand U1308 (N_1308,In_494,In_433);
nor U1309 (N_1309,In_643,In_492);
and U1310 (N_1310,In_130,In_160);
nor U1311 (N_1311,In_280,In_176);
and U1312 (N_1312,In_296,In_171);
or U1313 (N_1313,In_333,In_230);
nor U1314 (N_1314,In_617,In_192);
nand U1315 (N_1315,In_23,In_126);
and U1316 (N_1316,In_267,In_5);
or U1317 (N_1317,In_102,In_232);
nand U1318 (N_1318,In_547,In_181);
and U1319 (N_1319,In_70,In_676);
nor U1320 (N_1320,In_385,In_34);
nand U1321 (N_1321,In_595,In_671);
or U1322 (N_1322,In_235,In_724);
nand U1323 (N_1323,In_186,In_392);
or U1324 (N_1324,In_444,In_693);
nor U1325 (N_1325,In_743,In_557);
and U1326 (N_1326,In_696,In_374);
xnor U1327 (N_1327,In_12,In_681);
and U1328 (N_1328,In_673,In_341);
and U1329 (N_1329,In_138,In_294);
nand U1330 (N_1330,In_287,In_483);
or U1331 (N_1331,In_310,In_316);
and U1332 (N_1332,In_123,In_485);
nand U1333 (N_1333,In_604,In_594);
or U1334 (N_1334,In_61,In_339);
nand U1335 (N_1335,In_148,In_63);
nand U1336 (N_1336,In_440,In_46);
nor U1337 (N_1337,In_161,In_310);
nor U1338 (N_1338,In_424,In_561);
or U1339 (N_1339,In_218,In_484);
and U1340 (N_1340,In_522,In_619);
nand U1341 (N_1341,In_418,In_7);
nor U1342 (N_1342,In_706,In_523);
nand U1343 (N_1343,In_579,In_619);
or U1344 (N_1344,In_651,In_733);
nand U1345 (N_1345,In_84,In_367);
nand U1346 (N_1346,In_477,In_24);
nand U1347 (N_1347,In_260,In_303);
nor U1348 (N_1348,In_570,In_537);
nand U1349 (N_1349,In_36,In_89);
and U1350 (N_1350,In_662,In_190);
or U1351 (N_1351,In_194,In_728);
and U1352 (N_1352,In_283,In_35);
nand U1353 (N_1353,In_550,In_263);
nand U1354 (N_1354,In_596,In_664);
nor U1355 (N_1355,In_373,In_732);
nand U1356 (N_1356,In_353,In_119);
and U1357 (N_1357,In_25,In_712);
nor U1358 (N_1358,In_680,In_564);
or U1359 (N_1359,In_144,In_348);
nor U1360 (N_1360,In_614,In_239);
or U1361 (N_1361,In_355,In_215);
and U1362 (N_1362,In_594,In_399);
or U1363 (N_1363,In_508,In_686);
or U1364 (N_1364,In_223,In_28);
and U1365 (N_1365,In_600,In_189);
and U1366 (N_1366,In_276,In_139);
and U1367 (N_1367,In_341,In_358);
nor U1368 (N_1368,In_411,In_274);
and U1369 (N_1369,In_269,In_130);
and U1370 (N_1370,In_298,In_535);
or U1371 (N_1371,In_206,In_249);
and U1372 (N_1372,In_465,In_464);
nor U1373 (N_1373,In_493,In_236);
and U1374 (N_1374,In_574,In_31);
and U1375 (N_1375,In_603,In_700);
and U1376 (N_1376,In_170,In_364);
nand U1377 (N_1377,In_235,In_389);
or U1378 (N_1378,In_20,In_481);
nor U1379 (N_1379,In_601,In_227);
or U1380 (N_1380,In_214,In_464);
or U1381 (N_1381,In_607,In_622);
and U1382 (N_1382,In_215,In_616);
and U1383 (N_1383,In_676,In_630);
nand U1384 (N_1384,In_527,In_7);
nor U1385 (N_1385,In_578,In_596);
nor U1386 (N_1386,In_139,In_421);
nand U1387 (N_1387,In_178,In_194);
nand U1388 (N_1388,In_749,In_663);
nand U1389 (N_1389,In_713,In_640);
nor U1390 (N_1390,In_186,In_53);
or U1391 (N_1391,In_552,In_593);
and U1392 (N_1392,In_473,In_64);
nor U1393 (N_1393,In_77,In_309);
and U1394 (N_1394,In_713,In_335);
nor U1395 (N_1395,In_387,In_606);
nor U1396 (N_1396,In_586,In_449);
nor U1397 (N_1397,In_45,In_72);
nand U1398 (N_1398,In_573,In_612);
or U1399 (N_1399,In_630,In_626);
nand U1400 (N_1400,In_494,In_403);
and U1401 (N_1401,In_80,In_616);
nand U1402 (N_1402,In_514,In_468);
and U1403 (N_1403,In_726,In_648);
nor U1404 (N_1404,In_79,In_608);
nor U1405 (N_1405,In_273,In_435);
nor U1406 (N_1406,In_72,In_391);
and U1407 (N_1407,In_588,In_707);
and U1408 (N_1408,In_355,In_296);
or U1409 (N_1409,In_153,In_332);
and U1410 (N_1410,In_161,In_534);
and U1411 (N_1411,In_745,In_284);
or U1412 (N_1412,In_270,In_138);
nor U1413 (N_1413,In_61,In_255);
and U1414 (N_1414,In_705,In_208);
nor U1415 (N_1415,In_715,In_320);
nand U1416 (N_1416,In_54,In_88);
nor U1417 (N_1417,In_218,In_59);
and U1418 (N_1418,In_653,In_222);
nand U1419 (N_1419,In_1,In_383);
nand U1420 (N_1420,In_491,In_164);
nand U1421 (N_1421,In_356,In_598);
nor U1422 (N_1422,In_334,In_107);
or U1423 (N_1423,In_99,In_504);
nand U1424 (N_1424,In_599,In_685);
or U1425 (N_1425,In_482,In_634);
nor U1426 (N_1426,In_430,In_612);
and U1427 (N_1427,In_445,In_263);
and U1428 (N_1428,In_11,In_229);
or U1429 (N_1429,In_151,In_474);
and U1430 (N_1430,In_123,In_149);
and U1431 (N_1431,In_547,In_537);
and U1432 (N_1432,In_30,In_543);
nor U1433 (N_1433,In_610,In_15);
or U1434 (N_1434,In_394,In_108);
nor U1435 (N_1435,In_596,In_60);
and U1436 (N_1436,In_280,In_181);
nand U1437 (N_1437,In_731,In_605);
and U1438 (N_1438,In_2,In_264);
nor U1439 (N_1439,In_380,In_263);
or U1440 (N_1440,In_168,In_79);
or U1441 (N_1441,In_639,In_92);
or U1442 (N_1442,In_360,In_66);
or U1443 (N_1443,In_377,In_24);
nand U1444 (N_1444,In_144,In_213);
and U1445 (N_1445,In_671,In_109);
nand U1446 (N_1446,In_502,In_531);
nor U1447 (N_1447,In_196,In_609);
nor U1448 (N_1448,In_51,In_671);
nor U1449 (N_1449,In_426,In_640);
and U1450 (N_1450,In_380,In_359);
or U1451 (N_1451,In_439,In_236);
and U1452 (N_1452,In_170,In_308);
or U1453 (N_1453,In_317,In_87);
and U1454 (N_1454,In_324,In_18);
nor U1455 (N_1455,In_320,In_652);
nor U1456 (N_1456,In_631,In_376);
nand U1457 (N_1457,In_117,In_312);
or U1458 (N_1458,In_327,In_588);
nor U1459 (N_1459,In_582,In_372);
or U1460 (N_1460,In_495,In_50);
and U1461 (N_1461,In_216,In_399);
and U1462 (N_1462,In_610,In_548);
and U1463 (N_1463,In_99,In_31);
xnor U1464 (N_1464,In_272,In_565);
or U1465 (N_1465,In_579,In_491);
or U1466 (N_1466,In_366,In_420);
or U1467 (N_1467,In_639,In_309);
nor U1468 (N_1468,In_33,In_446);
and U1469 (N_1469,In_504,In_146);
and U1470 (N_1470,In_367,In_406);
nor U1471 (N_1471,In_368,In_450);
or U1472 (N_1472,In_74,In_559);
and U1473 (N_1473,In_49,In_635);
nand U1474 (N_1474,In_266,In_699);
or U1475 (N_1475,In_586,In_671);
or U1476 (N_1476,In_256,In_53);
and U1477 (N_1477,In_71,In_654);
or U1478 (N_1478,In_99,In_715);
and U1479 (N_1479,In_657,In_332);
nand U1480 (N_1480,In_63,In_379);
nor U1481 (N_1481,In_581,In_636);
and U1482 (N_1482,In_364,In_125);
nor U1483 (N_1483,In_655,In_514);
nor U1484 (N_1484,In_468,In_575);
nor U1485 (N_1485,In_78,In_511);
nand U1486 (N_1486,In_247,In_579);
and U1487 (N_1487,In_345,In_497);
and U1488 (N_1488,In_693,In_172);
or U1489 (N_1489,In_584,In_258);
nor U1490 (N_1490,In_50,In_513);
or U1491 (N_1491,In_140,In_280);
nor U1492 (N_1492,In_636,In_276);
and U1493 (N_1493,In_85,In_710);
or U1494 (N_1494,In_460,In_67);
nand U1495 (N_1495,In_239,In_294);
and U1496 (N_1496,In_256,In_697);
or U1497 (N_1497,In_738,In_381);
nor U1498 (N_1498,In_680,In_539);
nand U1499 (N_1499,In_495,In_404);
nor U1500 (N_1500,In_660,In_648);
nor U1501 (N_1501,In_266,In_39);
or U1502 (N_1502,In_102,In_574);
nor U1503 (N_1503,In_156,In_345);
and U1504 (N_1504,In_124,In_516);
nand U1505 (N_1505,In_251,In_472);
nor U1506 (N_1506,In_9,In_235);
nand U1507 (N_1507,In_292,In_525);
nand U1508 (N_1508,In_135,In_386);
or U1509 (N_1509,In_601,In_247);
and U1510 (N_1510,In_95,In_472);
or U1511 (N_1511,In_76,In_419);
nor U1512 (N_1512,In_53,In_455);
and U1513 (N_1513,In_734,In_194);
or U1514 (N_1514,In_602,In_408);
nor U1515 (N_1515,In_380,In_180);
and U1516 (N_1516,In_79,In_733);
nor U1517 (N_1517,In_246,In_239);
nand U1518 (N_1518,In_448,In_681);
or U1519 (N_1519,In_652,In_548);
or U1520 (N_1520,In_433,In_66);
and U1521 (N_1521,In_150,In_555);
and U1522 (N_1522,In_79,In_584);
nand U1523 (N_1523,In_98,In_694);
nand U1524 (N_1524,In_51,In_369);
nor U1525 (N_1525,In_516,In_58);
nor U1526 (N_1526,In_175,In_554);
or U1527 (N_1527,In_590,In_196);
nand U1528 (N_1528,In_721,In_358);
xor U1529 (N_1529,In_387,In_616);
nand U1530 (N_1530,In_362,In_683);
nor U1531 (N_1531,In_340,In_124);
and U1532 (N_1532,In_299,In_125);
or U1533 (N_1533,In_221,In_103);
nor U1534 (N_1534,In_576,In_296);
nor U1535 (N_1535,In_276,In_404);
nand U1536 (N_1536,In_195,In_705);
or U1537 (N_1537,In_20,In_47);
or U1538 (N_1538,In_23,In_305);
nand U1539 (N_1539,In_79,In_117);
or U1540 (N_1540,In_148,In_709);
or U1541 (N_1541,In_701,In_263);
or U1542 (N_1542,In_372,In_384);
nand U1543 (N_1543,In_467,In_507);
nor U1544 (N_1544,In_595,In_745);
or U1545 (N_1545,In_88,In_500);
nor U1546 (N_1546,In_172,In_643);
nand U1547 (N_1547,In_276,In_16);
nor U1548 (N_1548,In_234,In_703);
or U1549 (N_1549,In_186,In_249);
or U1550 (N_1550,In_548,In_708);
and U1551 (N_1551,In_182,In_425);
nor U1552 (N_1552,In_486,In_343);
nor U1553 (N_1553,In_680,In_275);
nand U1554 (N_1554,In_494,In_185);
nand U1555 (N_1555,In_321,In_443);
and U1556 (N_1556,In_500,In_383);
or U1557 (N_1557,In_509,In_287);
and U1558 (N_1558,In_427,In_479);
nand U1559 (N_1559,In_501,In_706);
and U1560 (N_1560,In_649,In_102);
nor U1561 (N_1561,In_663,In_641);
nor U1562 (N_1562,In_179,In_180);
nand U1563 (N_1563,In_647,In_136);
nand U1564 (N_1564,In_512,In_319);
nand U1565 (N_1565,In_188,In_41);
or U1566 (N_1566,In_37,In_123);
nor U1567 (N_1567,In_452,In_407);
and U1568 (N_1568,In_287,In_555);
nor U1569 (N_1569,In_561,In_683);
nor U1570 (N_1570,In_657,In_69);
and U1571 (N_1571,In_537,In_184);
nor U1572 (N_1572,In_469,In_138);
nand U1573 (N_1573,In_22,In_19);
nor U1574 (N_1574,In_8,In_38);
nand U1575 (N_1575,In_119,In_349);
nand U1576 (N_1576,In_436,In_283);
and U1577 (N_1577,In_108,In_706);
or U1578 (N_1578,In_363,In_126);
and U1579 (N_1579,In_315,In_263);
and U1580 (N_1580,In_581,In_422);
and U1581 (N_1581,In_424,In_436);
or U1582 (N_1582,In_10,In_266);
and U1583 (N_1583,In_406,In_88);
nand U1584 (N_1584,In_461,In_495);
or U1585 (N_1585,In_334,In_157);
and U1586 (N_1586,In_61,In_236);
and U1587 (N_1587,In_648,In_210);
nand U1588 (N_1588,In_327,In_89);
xnor U1589 (N_1589,In_466,In_424);
nand U1590 (N_1590,In_119,In_37);
nor U1591 (N_1591,In_483,In_357);
and U1592 (N_1592,In_718,In_502);
nor U1593 (N_1593,In_111,In_369);
and U1594 (N_1594,In_278,In_464);
nor U1595 (N_1595,In_620,In_616);
nor U1596 (N_1596,In_487,In_344);
and U1597 (N_1597,In_114,In_212);
or U1598 (N_1598,In_445,In_690);
and U1599 (N_1599,In_471,In_407);
or U1600 (N_1600,In_187,In_37);
and U1601 (N_1601,In_120,In_280);
nand U1602 (N_1602,In_311,In_479);
nand U1603 (N_1603,In_633,In_36);
and U1604 (N_1604,In_411,In_645);
and U1605 (N_1605,In_90,In_474);
nor U1606 (N_1606,In_384,In_424);
nor U1607 (N_1607,In_563,In_675);
and U1608 (N_1608,In_163,In_351);
and U1609 (N_1609,In_196,In_434);
and U1610 (N_1610,In_431,In_627);
nand U1611 (N_1611,In_690,In_325);
xor U1612 (N_1612,In_200,In_453);
nand U1613 (N_1613,In_379,In_217);
or U1614 (N_1614,In_558,In_448);
and U1615 (N_1615,In_703,In_110);
nand U1616 (N_1616,In_611,In_393);
and U1617 (N_1617,In_137,In_693);
nand U1618 (N_1618,In_357,In_741);
nand U1619 (N_1619,In_173,In_473);
or U1620 (N_1620,In_271,In_667);
or U1621 (N_1621,In_190,In_486);
or U1622 (N_1622,In_603,In_610);
nand U1623 (N_1623,In_732,In_238);
nor U1624 (N_1624,In_94,In_455);
nand U1625 (N_1625,In_485,In_170);
and U1626 (N_1626,In_209,In_53);
nor U1627 (N_1627,In_525,In_421);
and U1628 (N_1628,In_102,In_57);
and U1629 (N_1629,In_532,In_677);
nand U1630 (N_1630,In_241,In_568);
nand U1631 (N_1631,In_33,In_442);
nand U1632 (N_1632,In_380,In_71);
nand U1633 (N_1633,In_97,In_76);
or U1634 (N_1634,In_340,In_165);
and U1635 (N_1635,In_121,In_432);
nor U1636 (N_1636,In_279,In_562);
nand U1637 (N_1637,In_714,In_639);
or U1638 (N_1638,In_210,In_593);
or U1639 (N_1639,In_445,In_145);
and U1640 (N_1640,In_5,In_345);
nand U1641 (N_1641,In_167,In_399);
and U1642 (N_1642,In_352,In_130);
nand U1643 (N_1643,In_212,In_40);
and U1644 (N_1644,In_64,In_282);
nand U1645 (N_1645,In_642,In_548);
nand U1646 (N_1646,In_267,In_408);
nand U1647 (N_1647,In_83,In_536);
or U1648 (N_1648,In_532,In_160);
and U1649 (N_1649,In_522,In_699);
nor U1650 (N_1650,In_471,In_532);
nor U1651 (N_1651,In_297,In_523);
nor U1652 (N_1652,In_238,In_721);
nand U1653 (N_1653,In_140,In_409);
or U1654 (N_1654,In_30,In_473);
nor U1655 (N_1655,In_132,In_573);
nor U1656 (N_1656,In_120,In_576);
and U1657 (N_1657,In_178,In_338);
and U1658 (N_1658,In_612,In_170);
and U1659 (N_1659,In_556,In_578);
and U1660 (N_1660,In_30,In_104);
or U1661 (N_1661,In_482,In_519);
and U1662 (N_1662,In_708,In_716);
or U1663 (N_1663,In_614,In_699);
nor U1664 (N_1664,In_411,In_321);
and U1665 (N_1665,In_566,In_652);
nand U1666 (N_1666,In_63,In_310);
and U1667 (N_1667,In_299,In_133);
nand U1668 (N_1668,In_610,In_487);
or U1669 (N_1669,In_93,In_318);
or U1670 (N_1670,In_387,In_709);
and U1671 (N_1671,In_198,In_545);
nor U1672 (N_1672,In_511,In_440);
nor U1673 (N_1673,In_383,In_360);
xor U1674 (N_1674,In_597,In_450);
and U1675 (N_1675,In_424,In_211);
nor U1676 (N_1676,In_565,In_288);
nor U1677 (N_1677,In_610,In_18);
nand U1678 (N_1678,In_231,In_723);
nand U1679 (N_1679,In_399,In_67);
nor U1680 (N_1680,In_613,In_535);
and U1681 (N_1681,In_112,In_189);
nor U1682 (N_1682,In_675,In_658);
nor U1683 (N_1683,In_157,In_250);
nand U1684 (N_1684,In_287,In_142);
or U1685 (N_1685,In_579,In_724);
nor U1686 (N_1686,In_23,In_145);
nand U1687 (N_1687,In_608,In_682);
or U1688 (N_1688,In_386,In_180);
and U1689 (N_1689,In_372,In_617);
nor U1690 (N_1690,In_407,In_675);
or U1691 (N_1691,In_374,In_25);
nor U1692 (N_1692,In_395,In_491);
and U1693 (N_1693,In_745,In_145);
and U1694 (N_1694,In_285,In_403);
and U1695 (N_1695,In_611,In_263);
or U1696 (N_1696,In_460,In_721);
nor U1697 (N_1697,In_328,In_15);
nand U1698 (N_1698,In_397,In_423);
or U1699 (N_1699,In_386,In_733);
or U1700 (N_1700,In_46,In_717);
and U1701 (N_1701,In_100,In_542);
nand U1702 (N_1702,In_300,In_77);
or U1703 (N_1703,In_361,In_40);
or U1704 (N_1704,In_708,In_304);
nor U1705 (N_1705,In_183,In_523);
or U1706 (N_1706,In_223,In_105);
and U1707 (N_1707,In_219,In_427);
or U1708 (N_1708,In_92,In_515);
nand U1709 (N_1709,In_265,In_291);
nand U1710 (N_1710,In_381,In_560);
nand U1711 (N_1711,In_631,In_629);
and U1712 (N_1712,In_420,In_398);
xor U1713 (N_1713,In_719,In_496);
nor U1714 (N_1714,In_563,In_179);
and U1715 (N_1715,In_574,In_287);
and U1716 (N_1716,In_510,In_738);
and U1717 (N_1717,In_391,In_716);
nor U1718 (N_1718,In_648,In_606);
or U1719 (N_1719,In_728,In_695);
nor U1720 (N_1720,In_422,In_191);
and U1721 (N_1721,In_93,In_344);
nand U1722 (N_1722,In_91,In_131);
and U1723 (N_1723,In_546,In_7);
nor U1724 (N_1724,In_73,In_68);
and U1725 (N_1725,In_544,In_482);
or U1726 (N_1726,In_151,In_113);
nor U1727 (N_1727,In_441,In_639);
or U1728 (N_1728,In_13,In_378);
nand U1729 (N_1729,In_538,In_221);
nand U1730 (N_1730,In_175,In_636);
and U1731 (N_1731,In_588,In_246);
and U1732 (N_1732,In_291,In_691);
or U1733 (N_1733,In_393,In_429);
or U1734 (N_1734,In_12,In_204);
nor U1735 (N_1735,In_224,In_678);
and U1736 (N_1736,In_239,In_430);
xnor U1737 (N_1737,In_586,In_577);
and U1738 (N_1738,In_275,In_96);
or U1739 (N_1739,In_147,In_441);
nand U1740 (N_1740,In_470,In_46);
or U1741 (N_1741,In_701,In_304);
nor U1742 (N_1742,In_576,In_267);
and U1743 (N_1743,In_560,In_347);
nand U1744 (N_1744,In_136,In_719);
or U1745 (N_1745,In_414,In_366);
nor U1746 (N_1746,In_644,In_1);
and U1747 (N_1747,In_13,In_417);
xor U1748 (N_1748,In_624,In_359);
nand U1749 (N_1749,In_39,In_490);
or U1750 (N_1750,In_150,In_105);
nand U1751 (N_1751,In_625,In_216);
or U1752 (N_1752,In_284,In_460);
or U1753 (N_1753,In_58,In_91);
nand U1754 (N_1754,In_659,In_138);
and U1755 (N_1755,In_62,In_394);
or U1756 (N_1756,In_508,In_447);
and U1757 (N_1757,In_496,In_285);
nor U1758 (N_1758,In_109,In_422);
nor U1759 (N_1759,In_271,In_70);
or U1760 (N_1760,In_617,In_186);
and U1761 (N_1761,In_380,In_536);
or U1762 (N_1762,In_202,In_116);
nand U1763 (N_1763,In_9,In_175);
or U1764 (N_1764,In_278,In_185);
and U1765 (N_1765,In_445,In_368);
xnor U1766 (N_1766,In_146,In_281);
or U1767 (N_1767,In_174,In_326);
or U1768 (N_1768,In_583,In_106);
nor U1769 (N_1769,In_503,In_244);
or U1770 (N_1770,In_338,In_497);
and U1771 (N_1771,In_59,In_718);
nand U1772 (N_1772,In_675,In_469);
or U1773 (N_1773,In_140,In_555);
or U1774 (N_1774,In_410,In_689);
nand U1775 (N_1775,In_589,In_429);
nand U1776 (N_1776,In_511,In_293);
nor U1777 (N_1777,In_9,In_552);
and U1778 (N_1778,In_137,In_421);
nand U1779 (N_1779,In_66,In_275);
nand U1780 (N_1780,In_619,In_637);
nor U1781 (N_1781,In_535,In_58);
nand U1782 (N_1782,In_54,In_260);
nor U1783 (N_1783,In_460,In_192);
or U1784 (N_1784,In_545,In_569);
and U1785 (N_1785,In_334,In_232);
and U1786 (N_1786,In_176,In_239);
or U1787 (N_1787,In_206,In_19);
or U1788 (N_1788,In_272,In_220);
nand U1789 (N_1789,In_552,In_153);
nor U1790 (N_1790,In_388,In_557);
and U1791 (N_1791,In_50,In_18);
nor U1792 (N_1792,In_743,In_108);
nand U1793 (N_1793,In_433,In_366);
and U1794 (N_1794,In_500,In_60);
and U1795 (N_1795,In_734,In_416);
nand U1796 (N_1796,In_338,In_711);
nand U1797 (N_1797,In_202,In_305);
nor U1798 (N_1798,In_426,In_420);
nor U1799 (N_1799,In_109,In_499);
nand U1800 (N_1800,In_475,In_39);
or U1801 (N_1801,In_572,In_104);
and U1802 (N_1802,In_104,In_652);
and U1803 (N_1803,In_386,In_538);
xor U1804 (N_1804,In_180,In_400);
nor U1805 (N_1805,In_503,In_651);
nor U1806 (N_1806,In_468,In_527);
nor U1807 (N_1807,In_4,In_706);
nor U1808 (N_1808,In_342,In_127);
nand U1809 (N_1809,In_704,In_328);
or U1810 (N_1810,In_334,In_274);
nand U1811 (N_1811,In_696,In_124);
nor U1812 (N_1812,In_544,In_589);
xnor U1813 (N_1813,In_259,In_284);
nor U1814 (N_1814,In_202,In_218);
nor U1815 (N_1815,In_603,In_669);
or U1816 (N_1816,In_254,In_396);
nor U1817 (N_1817,In_606,In_351);
or U1818 (N_1818,In_352,In_541);
and U1819 (N_1819,In_62,In_259);
nor U1820 (N_1820,In_164,In_495);
nor U1821 (N_1821,In_472,In_664);
or U1822 (N_1822,In_378,In_382);
or U1823 (N_1823,In_357,In_17);
nand U1824 (N_1824,In_570,In_351);
nand U1825 (N_1825,In_374,In_742);
and U1826 (N_1826,In_370,In_6);
or U1827 (N_1827,In_302,In_273);
or U1828 (N_1828,In_122,In_72);
and U1829 (N_1829,In_577,In_661);
and U1830 (N_1830,In_226,In_102);
nor U1831 (N_1831,In_254,In_652);
nor U1832 (N_1832,In_581,In_286);
nand U1833 (N_1833,In_391,In_603);
xor U1834 (N_1834,In_346,In_439);
and U1835 (N_1835,In_122,In_501);
nor U1836 (N_1836,In_672,In_333);
or U1837 (N_1837,In_213,In_419);
and U1838 (N_1838,In_15,In_673);
or U1839 (N_1839,In_108,In_481);
nor U1840 (N_1840,In_86,In_270);
and U1841 (N_1841,In_516,In_521);
and U1842 (N_1842,In_133,In_231);
and U1843 (N_1843,In_616,In_200);
and U1844 (N_1844,In_147,In_203);
nor U1845 (N_1845,In_490,In_309);
and U1846 (N_1846,In_76,In_727);
nand U1847 (N_1847,In_429,In_395);
or U1848 (N_1848,In_63,In_382);
or U1849 (N_1849,In_645,In_270);
nor U1850 (N_1850,In_714,In_664);
nand U1851 (N_1851,In_176,In_414);
nor U1852 (N_1852,In_22,In_106);
nand U1853 (N_1853,In_659,In_177);
nand U1854 (N_1854,In_440,In_380);
nand U1855 (N_1855,In_546,In_383);
nand U1856 (N_1856,In_670,In_586);
nand U1857 (N_1857,In_380,In_484);
nor U1858 (N_1858,In_580,In_565);
nand U1859 (N_1859,In_595,In_549);
nand U1860 (N_1860,In_204,In_60);
nand U1861 (N_1861,In_408,In_603);
or U1862 (N_1862,In_731,In_707);
nor U1863 (N_1863,In_126,In_534);
or U1864 (N_1864,In_591,In_240);
or U1865 (N_1865,In_576,In_592);
and U1866 (N_1866,In_450,In_655);
nand U1867 (N_1867,In_517,In_167);
nand U1868 (N_1868,In_710,In_485);
nand U1869 (N_1869,In_748,In_660);
nand U1870 (N_1870,In_13,In_503);
xor U1871 (N_1871,In_28,In_587);
xor U1872 (N_1872,In_39,In_85);
nor U1873 (N_1873,In_574,In_170);
or U1874 (N_1874,In_446,In_348);
or U1875 (N_1875,In_646,In_370);
or U1876 (N_1876,In_111,In_477);
or U1877 (N_1877,In_80,In_335);
nor U1878 (N_1878,In_659,In_371);
nand U1879 (N_1879,In_701,In_486);
or U1880 (N_1880,In_337,In_717);
nand U1881 (N_1881,In_84,In_2);
and U1882 (N_1882,In_182,In_289);
nor U1883 (N_1883,In_382,In_631);
nand U1884 (N_1884,In_385,In_244);
or U1885 (N_1885,In_207,In_616);
nor U1886 (N_1886,In_359,In_234);
nand U1887 (N_1887,In_696,In_360);
nand U1888 (N_1888,In_736,In_122);
nor U1889 (N_1889,In_687,In_437);
or U1890 (N_1890,In_357,In_248);
or U1891 (N_1891,In_672,In_100);
nor U1892 (N_1892,In_398,In_3);
nor U1893 (N_1893,In_420,In_600);
nand U1894 (N_1894,In_720,In_696);
and U1895 (N_1895,In_327,In_524);
or U1896 (N_1896,In_367,In_401);
or U1897 (N_1897,In_553,In_609);
or U1898 (N_1898,In_428,In_297);
nor U1899 (N_1899,In_713,In_400);
nor U1900 (N_1900,In_615,In_220);
nor U1901 (N_1901,In_641,In_145);
and U1902 (N_1902,In_268,In_174);
nand U1903 (N_1903,In_400,In_534);
and U1904 (N_1904,In_552,In_728);
or U1905 (N_1905,In_187,In_622);
nor U1906 (N_1906,In_436,In_244);
or U1907 (N_1907,In_210,In_644);
or U1908 (N_1908,In_737,In_264);
or U1909 (N_1909,In_495,In_743);
nand U1910 (N_1910,In_394,In_675);
xnor U1911 (N_1911,In_498,In_723);
and U1912 (N_1912,In_177,In_440);
or U1913 (N_1913,In_234,In_416);
nor U1914 (N_1914,In_149,In_447);
nor U1915 (N_1915,In_466,In_644);
and U1916 (N_1916,In_489,In_733);
nor U1917 (N_1917,In_41,In_653);
nand U1918 (N_1918,In_671,In_180);
and U1919 (N_1919,In_289,In_559);
nand U1920 (N_1920,In_588,In_452);
or U1921 (N_1921,In_113,In_311);
nor U1922 (N_1922,In_545,In_38);
nor U1923 (N_1923,In_721,In_36);
and U1924 (N_1924,In_171,In_3);
nand U1925 (N_1925,In_515,In_41);
and U1926 (N_1926,In_470,In_328);
or U1927 (N_1927,In_134,In_266);
or U1928 (N_1928,In_402,In_478);
nand U1929 (N_1929,In_326,In_446);
nand U1930 (N_1930,In_569,In_66);
or U1931 (N_1931,In_468,In_492);
nor U1932 (N_1932,In_450,In_452);
and U1933 (N_1933,In_573,In_187);
nand U1934 (N_1934,In_127,In_110);
xor U1935 (N_1935,In_456,In_717);
nand U1936 (N_1936,In_283,In_578);
or U1937 (N_1937,In_84,In_731);
or U1938 (N_1938,In_222,In_434);
or U1939 (N_1939,In_684,In_22);
or U1940 (N_1940,In_63,In_549);
or U1941 (N_1941,In_616,In_348);
nor U1942 (N_1942,In_581,In_477);
nor U1943 (N_1943,In_354,In_11);
nand U1944 (N_1944,In_448,In_467);
or U1945 (N_1945,In_165,In_397);
nor U1946 (N_1946,In_473,In_728);
nand U1947 (N_1947,In_647,In_289);
and U1948 (N_1948,In_210,In_208);
xor U1949 (N_1949,In_118,In_346);
or U1950 (N_1950,In_127,In_412);
or U1951 (N_1951,In_743,In_81);
nand U1952 (N_1952,In_165,In_362);
and U1953 (N_1953,In_197,In_143);
nand U1954 (N_1954,In_69,In_523);
and U1955 (N_1955,In_614,In_228);
nor U1956 (N_1956,In_479,In_195);
and U1957 (N_1957,In_66,In_54);
nand U1958 (N_1958,In_484,In_549);
and U1959 (N_1959,In_353,In_670);
or U1960 (N_1960,In_320,In_247);
or U1961 (N_1961,In_676,In_668);
and U1962 (N_1962,In_376,In_559);
and U1963 (N_1963,In_236,In_641);
nor U1964 (N_1964,In_341,In_582);
or U1965 (N_1965,In_622,In_624);
nor U1966 (N_1966,In_83,In_59);
nand U1967 (N_1967,In_234,In_308);
nand U1968 (N_1968,In_19,In_124);
or U1969 (N_1969,In_648,In_293);
and U1970 (N_1970,In_122,In_343);
and U1971 (N_1971,In_245,In_418);
and U1972 (N_1972,In_688,In_378);
nand U1973 (N_1973,In_423,In_298);
nor U1974 (N_1974,In_651,In_365);
or U1975 (N_1975,In_89,In_275);
nand U1976 (N_1976,In_207,In_286);
nand U1977 (N_1977,In_196,In_556);
nand U1978 (N_1978,In_154,In_3);
and U1979 (N_1979,In_443,In_318);
nor U1980 (N_1980,In_53,In_418);
or U1981 (N_1981,In_55,In_425);
or U1982 (N_1982,In_67,In_627);
and U1983 (N_1983,In_563,In_188);
and U1984 (N_1984,In_533,In_484);
nand U1985 (N_1985,In_362,In_538);
and U1986 (N_1986,In_529,In_498);
nor U1987 (N_1987,In_91,In_312);
nor U1988 (N_1988,In_95,In_375);
nand U1989 (N_1989,In_35,In_386);
and U1990 (N_1990,In_377,In_492);
or U1991 (N_1991,In_3,In_178);
nor U1992 (N_1992,In_104,In_664);
nand U1993 (N_1993,In_614,In_505);
nor U1994 (N_1994,In_547,In_48);
or U1995 (N_1995,In_582,In_380);
nand U1996 (N_1996,In_333,In_609);
nand U1997 (N_1997,In_238,In_2);
nand U1998 (N_1998,In_177,In_169);
and U1999 (N_1999,In_136,In_264);
or U2000 (N_2000,In_463,In_659);
or U2001 (N_2001,In_97,In_133);
or U2002 (N_2002,In_10,In_381);
or U2003 (N_2003,In_445,In_312);
and U2004 (N_2004,In_653,In_556);
nor U2005 (N_2005,In_87,In_510);
nor U2006 (N_2006,In_608,In_173);
nor U2007 (N_2007,In_727,In_159);
and U2008 (N_2008,In_466,In_587);
nand U2009 (N_2009,In_627,In_444);
nor U2010 (N_2010,In_115,In_635);
nand U2011 (N_2011,In_312,In_174);
nor U2012 (N_2012,In_237,In_578);
and U2013 (N_2013,In_708,In_259);
nor U2014 (N_2014,In_51,In_187);
or U2015 (N_2015,In_381,In_155);
and U2016 (N_2016,In_442,In_269);
or U2017 (N_2017,In_239,In_644);
nor U2018 (N_2018,In_522,In_351);
nand U2019 (N_2019,In_645,In_15);
nor U2020 (N_2020,In_495,In_437);
nand U2021 (N_2021,In_585,In_127);
nor U2022 (N_2022,In_305,In_636);
nand U2023 (N_2023,In_215,In_328);
or U2024 (N_2024,In_689,In_425);
nor U2025 (N_2025,In_130,In_0);
and U2026 (N_2026,In_452,In_568);
nor U2027 (N_2027,In_263,In_286);
and U2028 (N_2028,In_87,In_350);
nand U2029 (N_2029,In_297,In_267);
xnor U2030 (N_2030,In_387,In_438);
nand U2031 (N_2031,In_442,In_183);
or U2032 (N_2032,In_464,In_540);
nand U2033 (N_2033,In_184,In_396);
nor U2034 (N_2034,In_608,In_684);
and U2035 (N_2035,In_212,In_519);
xor U2036 (N_2036,In_317,In_30);
nand U2037 (N_2037,In_325,In_514);
or U2038 (N_2038,In_193,In_737);
nand U2039 (N_2039,In_587,In_18);
nand U2040 (N_2040,In_379,In_332);
nand U2041 (N_2041,In_414,In_342);
nor U2042 (N_2042,In_317,In_702);
nand U2043 (N_2043,In_701,In_350);
and U2044 (N_2044,In_306,In_695);
nor U2045 (N_2045,In_374,In_529);
and U2046 (N_2046,In_71,In_263);
nor U2047 (N_2047,In_184,In_213);
and U2048 (N_2048,In_675,In_684);
nand U2049 (N_2049,In_652,In_559);
nand U2050 (N_2050,In_597,In_665);
nor U2051 (N_2051,In_377,In_544);
nor U2052 (N_2052,In_502,In_540);
or U2053 (N_2053,In_629,In_644);
nand U2054 (N_2054,In_703,In_631);
and U2055 (N_2055,In_159,In_7);
nand U2056 (N_2056,In_129,In_596);
nor U2057 (N_2057,In_379,In_210);
or U2058 (N_2058,In_634,In_599);
and U2059 (N_2059,In_51,In_70);
nand U2060 (N_2060,In_595,In_683);
nor U2061 (N_2061,In_103,In_112);
and U2062 (N_2062,In_458,In_696);
nor U2063 (N_2063,In_737,In_743);
nand U2064 (N_2064,In_581,In_629);
nand U2065 (N_2065,In_586,In_556);
or U2066 (N_2066,In_623,In_174);
and U2067 (N_2067,In_98,In_430);
or U2068 (N_2068,In_424,In_330);
nor U2069 (N_2069,In_355,In_278);
and U2070 (N_2070,In_314,In_241);
or U2071 (N_2071,In_193,In_157);
and U2072 (N_2072,In_160,In_66);
and U2073 (N_2073,In_503,In_269);
nand U2074 (N_2074,In_484,In_323);
nand U2075 (N_2075,In_74,In_540);
nand U2076 (N_2076,In_259,In_41);
nand U2077 (N_2077,In_447,In_229);
or U2078 (N_2078,In_665,In_105);
or U2079 (N_2079,In_311,In_602);
nand U2080 (N_2080,In_500,In_541);
and U2081 (N_2081,In_627,In_686);
or U2082 (N_2082,In_9,In_747);
nor U2083 (N_2083,In_159,In_65);
nor U2084 (N_2084,In_636,In_380);
nand U2085 (N_2085,In_145,In_15);
nor U2086 (N_2086,In_119,In_717);
and U2087 (N_2087,In_311,In_119);
or U2088 (N_2088,In_609,In_634);
and U2089 (N_2089,In_274,In_157);
nand U2090 (N_2090,In_6,In_254);
nor U2091 (N_2091,In_304,In_325);
nor U2092 (N_2092,In_52,In_588);
nand U2093 (N_2093,In_725,In_721);
xor U2094 (N_2094,In_105,In_207);
or U2095 (N_2095,In_623,In_88);
or U2096 (N_2096,In_101,In_475);
or U2097 (N_2097,In_506,In_406);
nor U2098 (N_2098,In_229,In_408);
nand U2099 (N_2099,In_529,In_284);
and U2100 (N_2100,In_694,In_495);
nand U2101 (N_2101,In_324,In_219);
and U2102 (N_2102,In_250,In_369);
or U2103 (N_2103,In_244,In_748);
nand U2104 (N_2104,In_7,In_362);
or U2105 (N_2105,In_54,In_249);
and U2106 (N_2106,In_199,In_745);
nand U2107 (N_2107,In_650,In_172);
and U2108 (N_2108,In_510,In_420);
nor U2109 (N_2109,In_281,In_629);
and U2110 (N_2110,In_597,In_138);
nand U2111 (N_2111,In_237,In_581);
nor U2112 (N_2112,In_596,In_65);
or U2113 (N_2113,In_507,In_574);
and U2114 (N_2114,In_727,In_546);
or U2115 (N_2115,In_574,In_713);
nor U2116 (N_2116,In_97,In_531);
and U2117 (N_2117,In_564,In_98);
nand U2118 (N_2118,In_531,In_193);
nand U2119 (N_2119,In_538,In_440);
and U2120 (N_2120,In_540,In_79);
nand U2121 (N_2121,In_196,In_577);
and U2122 (N_2122,In_129,In_263);
nor U2123 (N_2123,In_571,In_161);
nor U2124 (N_2124,In_722,In_424);
nor U2125 (N_2125,In_495,In_719);
or U2126 (N_2126,In_593,In_68);
or U2127 (N_2127,In_156,In_107);
nor U2128 (N_2128,In_680,In_388);
or U2129 (N_2129,In_638,In_642);
and U2130 (N_2130,In_198,In_58);
or U2131 (N_2131,In_388,In_419);
or U2132 (N_2132,In_601,In_720);
nor U2133 (N_2133,In_77,In_144);
and U2134 (N_2134,In_8,In_310);
or U2135 (N_2135,In_235,In_668);
nand U2136 (N_2136,In_9,In_115);
nand U2137 (N_2137,In_427,In_223);
or U2138 (N_2138,In_95,In_466);
and U2139 (N_2139,In_744,In_429);
nor U2140 (N_2140,In_535,In_192);
nor U2141 (N_2141,In_258,In_519);
nand U2142 (N_2142,In_663,In_433);
nand U2143 (N_2143,In_294,In_118);
and U2144 (N_2144,In_286,In_577);
nor U2145 (N_2145,In_340,In_168);
nor U2146 (N_2146,In_69,In_586);
or U2147 (N_2147,In_98,In_301);
or U2148 (N_2148,In_32,In_652);
nand U2149 (N_2149,In_74,In_265);
and U2150 (N_2150,In_34,In_333);
nand U2151 (N_2151,In_182,In_557);
nor U2152 (N_2152,In_189,In_363);
and U2153 (N_2153,In_56,In_474);
and U2154 (N_2154,In_727,In_673);
nand U2155 (N_2155,In_205,In_105);
nand U2156 (N_2156,In_280,In_685);
nor U2157 (N_2157,In_175,In_151);
xor U2158 (N_2158,In_443,In_720);
nand U2159 (N_2159,In_307,In_595);
or U2160 (N_2160,In_56,In_558);
or U2161 (N_2161,In_71,In_390);
or U2162 (N_2162,In_84,In_259);
and U2163 (N_2163,In_165,In_223);
nor U2164 (N_2164,In_158,In_626);
or U2165 (N_2165,In_541,In_123);
or U2166 (N_2166,In_445,In_733);
nor U2167 (N_2167,In_631,In_745);
or U2168 (N_2168,In_291,In_481);
or U2169 (N_2169,In_602,In_710);
or U2170 (N_2170,In_447,In_1);
or U2171 (N_2171,In_598,In_566);
nor U2172 (N_2172,In_44,In_137);
or U2173 (N_2173,In_665,In_726);
and U2174 (N_2174,In_697,In_405);
nor U2175 (N_2175,In_219,In_434);
nand U2176 (N_2176,In_282,In_278);
nand U2177 (N_2177,In_743,In_67);
and U2178 (N_2178,In_567,In_312);
and U2179 (N_2179,In_383,In_617);
nand U2180 (N_2180,In_147,In_576);
nand U2181 (N_2181,In_278,In_251);
nor U2182 (N_2182,In_555,In_219);
and U2183 (N_2183,In_545,In_634);
nand U2184 (N_2184,In_10,In_612);
and U2185 (N_2185,In_547,In_346);
or U2186 (N_2186,In_105,In_49);
nand U2187 (N_2187,In_112,In_504);
and U2188 (N_2188,In_49,In_20);
nand U2189 (N_2189,In_659,In_242);
nand U2190 (N_2190,In_123,In_35);
or U2191 (N_2191,In_64,In_444);
and U2192 (N_2192,In_350,In_588);
nor U2193 (N_2193,In_143,In_48);
nor U2194 (N_2194,In_602,In_53);
or U2195 (N_2195,In_425,In_415);
or U2196 (N_2196,In_249,In_74);
nand U2197 (N_2197,In_595,In_614);
and U2198 (N_2198,In_586,In_582);
nor U2199 (N_2199,In_640,In_617);
and U2200 (N_2200,In_427,In_629);
nor U2201 (N_2201,In_512,In_551);
nor U2202 (N_2202,In_137,In_625);
and U2203 (N_2203,In_19,In_742);
or U2204 (N_2204,In_167,In_684);
or U2205 (N_2205,In_196,In_641);
and U2206 (N_2206,In_265,In_220);
and U2207 (N_2207,In_193,In_24);
and U2208 (N_2208,In_152,In_626);
nor U2209 (N_2209,In_393,In_69);
nor U2210 (N_2210,In_77,In_66);
or U2211 (N_2211,In_495,In_521);
nor U2212 (N_2212,In_620,In_115);
nand U2213 (N_2213,In_196,In_20);
nand U2214 (N_2214,In_118,In_92);
nand U2215 (N_2215,In_329,In_560);
or U2216 (N_2216,In_643,In_280);
nor U2217 (N_2217,In_400,In_135);
nor U2218 (N_2218,In_383,In_15);
and U2219 (N_2219,In_456,In_4);
xnor U2220 (N_2220,In_157,In_460);
nand U2221 (N_2221,In_608,In_127);
and U2222 (N_2222,In_537,In_62);
nor U2223 (N_2223,In_41,In_627);
and U2224 (N_2224,In_174,In_411);
and U2225 (N_2225,In_623,In_341);
xnor U2226 (N_2226,In_669,In_375);
nor U2227 (N_2227,In_719,In_251);
and U2228 (N_2228,In_711,In_103);
or U2229 (N_2229,In_624,In_94);
or U2230 (N_2230,In_660,In_441);
nand U2231 (N_2231,In_79,In_73);
and U2232 (N_2232,In_404,In_115);
nand U2233 (N_2233,In_220,In_289);
or U2234 (N_2234,In_520,In_301);
nand U2235 (N_2235,In_654,In_26);
and U2236 (N_2236,In_196,In_333);
or U2237 (N_2237,In_549,In_214);
and U2238 (N_2238,In_644,In_700);
nor U2239 (N_2239,In_648,In_719);
nand U2240 (N_2240,In_558,In_486);
nor U2241 (N_2241,In_520,In_676);
nand U2242 (N_2242,In_373,In_705);
nor U2243 (N_2243,In_537,In_213);
nand U2244 (N_2244,In_247,In_690);
and U2245 (N_2245,In_522,In_542);
nand U2246 (N_2246,In_387,In_58);
nand U2247 (N_2247,In_12,In_299);
nor U2248 (N_2248,In_35,In_185);
or U2249 (N_2249,In_104,In_325);
nor U2250 (N_2250,In_416,In_29);
or U2251 (N_2251,In_723,In_493);
or U2252 (N_2252,In_55,In_517);
or U2253 (N_2253,In_469,In_227);
or U2254 (N_2254,In_516,In_215);
or U2255 (N_2255,In_14,In_283);
nand U2256 (N_2256,In_357,In_265);
nand U2257 (N_2257,In_99,In_371);
nand U2258 (N_2258,In_333,In_264);
nor U2259 (N_2259,In_48,In_81);
or U2260 (N_2260,In_444,In_115);
and U2261 (N_2261,In_623,In_321);
nand U2262 (N_2262,In_355,In_121);
and U2263 (N_2263,In_552,In_23);
nor U2264 (N_2264,In_712,In_150);
nand U2265 (N_2265,In_741,In_366);
nor U2266 (N_2266,In_418,In_171);
nand U2267 (N_2267,In_399,In_265);
nor U2268 (N_2268,In_301,In_143);
nor U2269 (N_2269,In_9,In_37);
or U2270 (N_2270,In_36,In_158);
nor U2271 (N_2271,In_518,In_225);
and U2272 (N_2272,In_741,In_716);
nor U2273 (N_2273,In_7,In_143);
nand U2274 (N_2274,In_324,In_93);
nand U2275 (N_2275,In_501,In_265);
nor U2276 (N_2276,In_136,In_428);
nor U2277 (N_2277,In_298,In_280);
nand U2278 (N_2278,In_443,In_700);
nand U2279 (N_2279,In_193,In_391);
and U2280 (N_2280,In_290,In_534);
nor U2281 (N_2281,In_527,In_634);
nor U2282 (N_2282,In_547,In_570);
nor U2283 (N_2283,In_171,In_248);
or U2284 (N_2284,In_59,In_359);
nor U2285 (N_2285,In_618,In_21);
and U2286 (N_2286,In_748,In_670);
and U2287 (N_2287,In_472,In_261);
nand U2288 (N_2288,In_127,In_147);
nand U2289 (N_2289,In_407,In_93);
or U2290 (N_2290,In_14,In_596);
and U2291 (N_2291,In_112,In_499);
or U2292 (N_2292,In_527,In_617);
nand U2293 (N_2293,In_241,In_680);
or U2294 (N_2294,In_291,In_318);
nor U2295 (N_2295,In_214,In_408);
nand U2296 (N_2296,In_479,In_22);
and U2297 (N_2297,In_522,In_137);
nand U2298 (N_2298,In_185,In_394);
and U2299 (N_2299,In_100,In_88);
or U2300 (N_2300,In_677,In_245);
and U2301 (N_2301,In_532,In_63);
nand U2302 (N_2302,In_503,In_337);
nand U2303 (N_2303,In_628,In_364);
nand U2304 (N_2304,In_103,In_569);
nand U2305 (N_2305,In_150,In_328);
or U2306 (N_2306,In_227,In_480);
or U2307 (N_2307,In_721,In_540);
or U2308 (N_2308,In_133,In_409);
nor U2309 (N_2309,In_555,In_430);
and U2310 (N_2310,In_534,In_103);
and U2311 (N_2311,In_179,In_136);
nor U2312 (N_2312,In_207,In_629);
nand U2313 (N_2313,In_738,In_571);
nor U2314 (N_2314,In_86,In_393);
nand U2315 (N_2315,In_505,In_648);
nand U2316 (N_2316,In_514,In_601);
and U2317 (N_2317,In_299,In_579);
or U2318 (N_2318,In_649,In_723);
nor U2319 (N_2319,In_317,In_536);
nand U2320 (N_2320,In_697,In_339);
and U2321 (N_2321,In_734,In_720);
or U2322 (N_2322,In_621,In_101);
and U2323 (N_2323,In_125,In_55);
and U2324 (N_2324,In_523,In_347);
nand U2325 (N_2325,In_281,In_189);
or U2326 (N_2326,In_298,In_8);
and U2327 (N_2327,In_50,In_200);
nor U2328 (N_2328,In_76,In_654);
and U2329 (N_2329,In_294,In_626);
and U2330 (N_2330,In_353,In_739);
or U2331 (N_2331,In_67,In_154);
or U2332 (N_2332,In_413,In_637);
nand U2333 (N_2333,In_496,In_124);
and U2334 (N_2334,In_519,In_303);
or U2335 (N_2335,In_596,In_220);
or U2336 (N_2336,In_735,In_683);
or U2337 (N_2337,In_124,In_642);
nor U2338 (N_2338,In_91,In_613);
nor U2339 (N_2339,In_563,In_441);
and U2340 (N_2340,In_611,In_150);
nor U2341 (N_2341,In_472,In_602);
nor U2342 (N_2342,In_482,In_137);
and U2343 (N_2343,In_367,In_105);
and U2344 (N_2344,In_554,In_43);
and U2345 (N_2345,In_733,In_327);
nand U2346 (N_2346,In_304,In_507);
nor U2347 (N_2347,In_26,In_314);
nor U2348 (N_2348,In_46,In_673);
or U2349 (N_2349,In_634,In_577);
and U2350 (N_2350,In_560,In_727);
and U2351 (N_2351,In_504,In_66);
nand U2352 (N_2352,In_458,In_450);
and U2353 (N_2353,In_636,In_360);
nor U2354 (N_2354,In_612,In_533);
nand U2355 (N_2355,In_576,In_15);
nand U2356 (N_2356,In_366,In_81);
nor U2357 (N_2357,In_481,In_146);
nand U2358 (N_2358,In_625,In_79);
nor U2359 (N_2359,In_585,In_371);
nand U2360 (N_2360,In_124,In_70);
or U2361 (N_2361,In_695,In_685);
or U2362 (N_2362,In_648,In_715);
and U2363 (N_2363,In_575,In_490);
xor U2364 (N_2364,In_447,In_7);
nand U2365 (N_2365,In_397,In_682);
nand U2366 (N_2366,In_25,In_439);
and U2367 (N_2367,In_332,In_321);
nand U2368 (N_2368,In_256,In_428);
and U2369 (N_2369,In_574,In_79);
nor U2370 (N_2370,In_741,In_19);
nor U2371 (N_2371,In_455,In_695);
or U2372 (N_2372,In_559,In_333);
nor U2373 (N_2373,In_258,In_89);
xnor U2374 (N_2374,In_274,In_281);
or U2375 (N_2375,In_64,In_263);
nor U2376 (N_2376,In_749,In_465);
and U2377 (N_2377,In_427,In_154);
and U2378 (N_2378,In_532,In_435);
or U2379 (N_2379,In_649,In_179);
and U2380 (N_2380,In_252,In_292);
nand U2381 (N_2381,In_31,In_620);
and U2382 (N_2382,In_413,In_530);
and U2383 (N_2383,In_37,In_152);
and U2384 (N_2384,In_252,In_290);
nor U2385 (N_2385,In_62,In_324);
xor U2386 (N_2386,In_383,In_656);
and U2387 (N_2387,In_409,In_362);
or U2388 (N_2388,In_562,In_378);
and U2389 (N_2389,In_721,In_643);
or U2390 (N_2390,In_590,In_207);
and U2391 (N_2391,In_453,In_393);
and U2392 (N_2392,In_152,In_253);
or U2393 (N_2393,In_138,In_372);
or U2394 (N_2394,In_734,In_143);
or U2395 (N_2395,In_375,In_172);
or U2396 (N_2396,In_659,In_601);
and U2397 (N_2397,In_565,In_187);
and U2398 (N_2398,In_587,In_492);
nor U2399 (N_2399,In_567,In_334);
nor U2400 (N_2400,In_262,In_119);
nor U2401 (N_2401,In_77,In_606);
nand U2402 (N_2402,In_523,In_206);
nand U2403 (N_2403,In_442,In_102);
nor U2404 (N_2404,In_721,In_583);
nand U2405 (N_2405,In_626,In_588);
and U2406 (N_2406,In_27,In_568);
nand U2407 (N_2407,In_231,In_746);
nand U2408 (N_2408,In_104,In_276);
nand U2409 (N_2409,In_724,In_572);
or U2410 (N_2410,In_167,In_575);
and U2411 (N_2411,In_22,In_310);
or U2412 (N_2412,In_312,In_164);
nor U2413 (N_2413,In_33,In_620);
or U2414 (N_2414,In_381,In_314);
nand U2415 (N_2415,In_41,In_672);
nand U2416 (N_2416,In_729,In_697);
nor U2417 (N_2417,In_617,In_156);
nor U2418 (N_2418,In_518,In_137);
nand U2419 (N_2419,In_120,In_202);
nor U2420 (N_2420,In_71,In_438);
or U2421 (N_2421,In_155,In_427);
and U2422 (N_2422,In_603,In_429);
or U2423 (N_2423,In_385,In_417);
nor U2424 (N_2424,In_293,In_365);
nor U2425 (N_2425,In_735,In_681);
nand U2426 (N_2426,In_104,In_145);
or U2427 (N_2427,In_88,In_604);
nor U2428 (N_2428,In_741,In_587);
nor U2429 (N_2429,In_687,In_119);
or U2430 (N_2430,In_592,In_616);
and U2431 (N_2431,In_166,In_480);
nand U2432 (N_2432,In_631,In_412);
nand U2433 (N_2433,In_562,In_549);
nor U2434 (N_2434,In_349,In_397);
or U2435 (N_2435,In_691,In_488);
or U2436 (N_2436,In_260,In_417);
nor U2437 (N_2437,In_57,In_420);
and U2438 (N_2438,In_518,In_682);
nor U2439 (N_2439,In_308,In_538);
nand U2440 (N_2440,In_453,In_300);
or U2441 (N_2441,In_482,In_113);
nor U2442 (N_2442,In_210,In_505);
nand U2443 (N_2443,In_309,In_141);
nand U2444 (N_2444,In_736,In_591);
nor U2445 (N_2445,In_71,In_720);
or U2446 (N_2446,In_51,In_288);
or U2447 (N_2447,In_457,In_181);
or U2448 (N_2448,In_700,In_164);
and U2449 (N_2449,In_200,In_344);
nand U2450 (N_2450,In_420,In_673);
or U2451 (N_2451,In_686,In_111);
nand U2452 (N_2452,In_397,In_381);
or U2453 (N_2453,In_423,In_573);
nor U2454 (N_2454,In_60,In_746);
nor U2455 (N_2455,In_738,In_256);
nand U2456 (N_2456,In_738,In_345);
and U2457 (N_2457,In_403,In_0);
nor U2458 (N_2458,In_245,In_516);
or U2459 (N_2459,In_695,In_339);
nor U2460 (N_2460,In_365,In_225);
or U2461 (N_2461,In_632,In_221);
nand U2462 (N_2462,In_420,In_523);
or U2463 (N_2463,In_337,In_446);
nand U2464 (N_2464,In_560,In_108);
or U2465 (N_2465,In_92,In_160);
and U2466 (N_2466,In_729,In_159);
and U2467 (N_2467,In_313,In_728);
nor U2468 (N_2468,In_268,In_543);
and U2469 (N_2469,In_281,In_330);
or U2470 (N_2470,In_541,In_425);
or U2471 (N_2471,In_82,In_749);
nor U2472 (N_2472,In_178,In_426);
nand U2473 (N_2473,In_697,In_186);
nand U2474 (N_2474,In_405,In_138);
and U2475 (N_2475,In_672,In_465);
and U2476 (N_2476,In_485,In_701);
or U2477 (N_2477,In_478,In_575);
and U2478 (N_2478,In_462,In_491);
and U2479 (N_2479,In_167,In_577);
nor U2480 (N_2480,In_550,In_65);
nand U2481 (N_2481,In_196,In_729);
or U2482 (N_2482,In_95,In_415);
nor U2483 (N_2483,In_460,In_280);
nand U2484 (N_2484,In_437,In_434);
nor U2485 (N_2485,In_328,In_68);
or U2486 (N_2486,In_103,In_350);
nor U2487 (N_2487,In_72,In_419);
and U2488 (N_2488,In_587,In_126);
and U2489 (N_2489,In_630,In_135);
nand U2490 (N_2490,In_132,In_170);
and U2491 (N_2491,In_484,In_575);
or U2492 (N_2492,In_699,In_111);
and U2493 (N_2493,In_610,In_560);
nand U2494 (N_2494,In_671,In_717);
xnor U2495 (N_2495,In_277,In_326);
nor U2496 (N_2496,In_480,In_375);
or U2497 (N_2497,In_477,In_248);
and U2498 (N_2498,In_121,In_602);
or U2499 (N_2499,In_39,In_437);
or U2500 (N_2500,N_651,N_2217);
nand U2501 (N_2501,N_69,N_1629);
nand U2502 (N_2502,N_2208,N_2048);
nand U2503 (N_2503,N_2398,N_916);
xor U2504 (N_2504,N_914,N_2431);
nand U2505 (N_2505,N_62,N_921);
or U2506 (N_2506,N_875,N_360);
nand U2507 (N_2507,N_1748,N_1651);
nor U2508 (N_2508,N_695,N_981);
nand U2509 (N_2509,N_624,N_2414);
or U2510 (N_2510,N_1751,N_17);
nand U2511 (N_2511,N_190,N_110);
nand U2512 (N_2512,N_619,N_195);
nand U2513 (N_2513,N_2311,N_741);
nor U2514 (N_2514,N_577,N_1574);
nor U2515 (N_2515,N_2413,N_1541);
and U2516 (N_2516,N_955,N_917);
nor U2517 (N_2517,N_1167,N_544);
nor U2518 (N_2518,N_400,N_1068);
or U2519 (N_2519,N_1017,N_1140);
and U2520 (N_2520,N_1846,N_1203);
or U2521 (N_2521,N_563,N_1159);
nand U2522 (N_2522,N_1654,N_2106);
nand U2523 (N_2523,N_1549,N_1301);
and U2524 (N_2524,N_517,N_1190);
or U2525 (N_2525,N_2293,N_1216);
and U2526 (N_2526,N_1682,N_642);
and U2527 (N_2527,N_1362,N_494);
and U2528 (N_2528,N_1117,N_1094);
nor U2529 (N_2529,N_1200,N_1835);
and U2530 (N_2530,N_1186,N_209);
nand U2531 (N_2531,N_2103,N_15);
or U2532 (N_2532,N_1533,N_594);
nand U2533 (N_2533,N_1185,N_808);
and U2534 (N_2534,N_1432,N_724);
nor U2535 (N_2535,N_1838,N_1197);
nand U2536 (N_2536,N_899,N_1223);
nand U2537 (N_2537,N_627,N_3);
nor U2538 (N_2538,N_933,N_227);
nand U2539 (N_2539,N_1022,N_971);
or U2540 (N_2540,N_529,N_1287);
and U2541 (N_2541,N_2484,N_1779);
or U2542 (N_2542,N_1647,N_2185);
or U2543 (N_2543,N_882,N_1799);
nand U2544 (N_2544,N_519,N_1026);
and U2545 (N_2545,N_837,N_1305);
and U2546 (N_2546,N_1812,N_784);
nand U2547 (N_2547,N_202,N_2055);
nor U2548 (N_2548,N_1340,N_1980);
nand U2549 (N_2549,N_632,N_339);
or U2550 (N_2550,N_2120,N_622);
and U2551 (N_2551,N_1826,N_1614);
nor U2552 (N_2552,N_1282,N_946);
and U2553 (N_2553,N_950,N_1323);
nand U2554 (N_2554,N_363,N_1283);
or U2555 (N_2555,N_450,N_1037);
nand U2556 (N_2556,N_2189,N_351);
and U2557 (N_2557,N_1859,N_1767);
nor U2558 (N_2558,N_252,N_1130);
nand U2559 (N_2559,N_2335,N_731);
and U2560 (N_2560,N_1095,N_1688);
or U2561 (N_2561,N_247,N_1844);
nor U2562 (N_2562,N_1039,N_2029);
and U2563 (N_2563,N_2118,N_1866);
nand U2564 (N_2564,N_222,N_1448);
nor U2565 (N_2565,N_1243,N_2099);
or U2566 (N_2566,N_616,N_930);
and U2567 (N_2567,N_614,N_2463);
and U2568 (N_2568,N_565,N_1394);
nor U2569 (N_2569,N_2421,N_1319);
and U2570 (N_2570,N_1630,N_962);
nand U2571 (N_2571,N_1255,N_0);
or U2572 (N_2572,N_1373,N_1357);
nor U2573 (N_2573,N_151,N_282);
nand U2574 (N_2574,N_1108,N_1723);
and U2575 (N_2575,N_1031,N_894);
or U2576 (N_2576,N_1825,N_1518);
nor U2577 (N_2577,N_1011,N_136);
nor U2578 (N_2578,N_1579,N_1910);
or U2579 (N_2579,N_860,N_57);
and U2580 (N_2580,N_211,N_2296);
and U2581 (N_2581,N_569,N_2127);
nand U2582 (N_2582,N_698,N_1953);
nor U2583 (N_2583,N_150,N_1211);
nor U2584 (N_2584,N_1551,N_602);
nor U2585 (N_2585,N_653,N_114);
or U2586 (N_2586,N_809,N_1959);
and U2587 (N_2587,N_1388,N_270);
nor U2588 (N_2588,N_421,N_835);
and U2589 (N_2589,N_2038,N_604);
or U2590 (N_2590,N_1438,N_2188);
or U2591 (N_2591,N_109,N_1450);
or U2592 (N_2592,N_2134,N_1155);
or U2593 (N_2593,N_1643,N_1033);
or U2594 (N_2594,N_1034,N_1585);
and U2595 (N_2595,N_975,N_2126);
nand U2596 (N_2596,N_2301,N_343);
nor U2597 (N_2597,N_21,N_1027);
nor U2598 (N_2598,N_856,N_1868);
or U2599 (N_2599,N_672,N_838);
nand U2600 (N_2600,N_2012,N_24);
and U2601 (N_2601,N_1934,N_1891);
or U2602 (N_2602,N_1106,N_883);
and U2603 (N_2603,N_306,N_559);
nor U2604 (N_2604,N_797,N_1435);
nor U2605 (N_2605,N_201,N_302);
nor U2606 (N_2606,N_116,N_1047);
xor U2607 (N_2607,N_999,N_754);
or U2608 (N_2608,N_1046,N_2112);
nand U2609 (N_2609,N_64,N_684);
nand U2610 (N_2610,N_1119,N_582);
or U2611 (N_2611,N_716,N_1493);
or U2612 (N_2612,N_271,N_1831);
and U2613 (N_2613,N_53,N_2137);
and U2614 (N_2614,N_285,N_1770);
nor U2615 (N_2615,N_726,N_2409);
nand U2616 (N_2616,N_97,N_682);
or U2617 (N_2617,N_1753,N_314);
and U2618 (N_2618,N_1995,N_196);
nor U2619 (N_2619,N_954,N_1171);
nand U2620 (N_2620,N_1136,N_1138);
nand U2621 (N_2621,N_1750,N_501);
nor U2622 (N_2622,N_348,N_800);
and U2623 (N_2623,N_75,N_1987);
or U2624 (N_2624,N_973,N_979);
nand U2625 (N_2625,N_2437,N_1338);
or U2626 (N_2626,N_1152,N_1871);
and U2627 (N_2627,N_2128,N_1102);
nand U2628 (N_2628,N_841,N_2042);
or U2629 (N_2629,N_1019,N_2322);
nor U2630 (N_2630,N_74,N_958);
nor U2631 (N_2631,N_350,N_1942);
nand U2632 (N_2632,N_1917,N_1150);
nand U2633 (N_2633,N_2101,N_405);
nor U2634 (N_2634,N_948,N_493);
nor U2635 (N_2635,N_1856,N_1949);
or U2636 (N_2636,N_2385,N_681);
or U2637 (N_2637,N_783,N_850);
or U2638 (N_2638,N_481,N_2034);
and U2639 (N_2639,N_479,N_2320);
and U2640 (N_2640,N_2058,N_1928);
and U2641 (N_2641,N_2054,N_488);
nor U2642 (N_2642,N_94,N_1086);
nand U2643 (N_2643,N_669,N_1659);
or U2644 (N_2644,N_857,N_2190);
and U2645 (N_2645,N_1091,N_1121);
nor U2646 (N_2646,N_492,N_2419);
or U2647 (N_2647,N_2132,N_2346);
nor U2648 (N_2648,N_35,N_1653);
nand U2649 (N_2649,N_1342,N_1001);
and U2650 (N_2650,N_647,N_1529);
nor U2651 (N_2651,N_1510,N_1116);
nand U2652 (N_2652,N_2473,N_1423);
or U2653 (N_2653,N_2420,N_192);
or U2654 (N_2654,N_1872,N_2019);
and U2655 (N_2655,N_18,N_1097);
nor U2656 (N_2656,N_1073,N_819);
and U2657 (N_2657,N_1007,N_58);
or U2658 (N_2658,N_375,N_2098);
or U2659 (N_2659,N_1578,N_2192);
nand U2660 (N_2660,N_1970,N_1466);
and U2661 (N_2661,N_660,N_1505);
and U2662 (N_2662,N_522,N_2018);
and U2663 (N_2663,N_1530,N_1110);
and U2664 (N_2664,N_248,N_1479);
and U2665 (N_2665,N_277,N_2003);
and U2666 (N_2666,N_2364,N_1271);
nand U2667 (N_2667,N_1237,N_1326);
nand U2668 (N_2668,N_1259,N_1372);
nor U2669 (N_2669,N_2025,N_1898);
nor U2670 (N_2670,N_701,N_1410);
nor U2671 (N_2671,N_1904,N_118);
and U2672 (N_2672,N_1576,N_1849);
nor U2673 (N_2673,N_1367,N_336);
nor U2674 (N_2674,N_1727,N_297);
nor U2675 (N_2675,N_1419,N_499);
and U2676 (N_2676,N_2040,N_359);
or U2677 (N_2677,N_1177,N_1991);
nor U2678 (N_2678,N_312,N_1424);
nor U2679 (N_2679,N_2044,N_2314);
and U2680 (N_2680,N_154,N_1407);
nand U2681 (N_2681,N_2016,N_1355);
and U2682 (N_2682,N_1157,N_2418);
nand U2683 (N_2683,N_1523,N_2388);
nand U2684 (N_2684,N_2139,N_652);
and U2685 (N_2685,N_2352,N_1266);
nand U2686 (N_2686,N_551,N_890);
xnor U2687 (N_2687,N_1238,N_2417);
and U2688 (N_2688,N_465,N_251);
or U2689 (N_2689,N_2154,N_1884);
nand U2690 (N_2690,N_1621,N_147);
nor U2691 (N_2691,N_729,N_609);
or U2692 (N_2692,N_1181,N_1620);
nand U2693 (N_2693,N_985,N_1382);
and U2694 (N_2694,N_1343,N_900);
or U2695 (N_2695,N_1596,N_199);
and U2696 (N_2696,N_1484,N_2173);
nor U2697 (N_2697,N_520,N_2367);
nand U2698 (N_2698,N_152,N_1933);
nor U2699 (N_2699,N_2408,N_61);
or U2700 (N_2700,N_286,N_1650);
or U2701 (N_2701,N_765,N_2156);
nand U2702 (N_2702,N_203,N_239);
nor U2703 (N_2703,N_1636,N_1896);
or U2704 (N_2704,N_2474,N_1416);
or U2705 (N_2705,N_1724,N_743);
nand U2706 (N_2706,N_969,N_1199);
and U2707 (N_2707,N_2261,N_1060);
and U2708 (N_2708,N_2422,N_1522);
nand U2709 (N_2709,N_2109,N_36);
nand U2710 (N_2710,N_2002,N_2215);
nand U2711 (N_2711,N_929,N_238);
and U2712 (N_2712,N_399,N_1024);
and U2713 (N_2713,N_2292,N_1145);
nor U2714 (N_2714,N_266,N_361);
or U2715 (N_2715,N_710,N_1858);
nand U2716 (N_2716,N_1789,N_2465);
nor U2717 (N_2717,N_483,N_1344);
nand U2718 (N_2718,N_1721,N_46);
and U2719 (N_2719,N_554,N_1464);
nand U2720 (N_2720,N_54,N_1137);
and U2721 (N_2721,N_156,N_1778);
nor U2722 (N_2722,N_323,N_1716);
nand U2723 (N_2723,N_1187,N_37);
nor U2724 (N_2724,N_1881,N_810);
and U2725 (N_2725,N_281,N_1729);
nor U2726 (N_2726,N_1469,N_1916);
and U2727 (N_2727,N_589,N_597);
and U2728 (N_2728,N_730,N_81);
nand U2729 (N_2729,N_305,N_1125);
nand U2730 (N_2730,N_1863,N_2080);
or U2731 (N_2731,N_1314,N_993);
and U2732 (N_2732,N_2186,N_1712);
nor U2733 (N_2733,N_2359,N_853);
nor U2734 (N_2734,N_1945,N_854);
or U2735 (N_2735,N_245,N_1132);
nor U2736 (N_2736,N_489,N_472);
nand U2737 (N_2737,N_1417,N_524);
or U2738 (N_2738,N_1536,N_980);
nor U2739 (N_2739,N_163,N_903);
and U2740 (N_2740,N_1127,N_2248);
or U2741 (N_2741,N_1892,N_388);
nor U2742 (N_2742,N_51,N_249);
nor U2743 (N_2743,N_1428,N_732);
or U2744 (N_2744,N_1514,N_1865);
or U2745 (N_2745,N_223,N_744);
nand U2746 (N_2746,N_1504,N_1524);
nand U2747 (N_2747,N_1371,N_2165);
nor U2748 (N_2748,N_2466,N_462);
and U2749 (N_2749,N_1590,N_1085);
and U2750 (N_2750,N_1817,N_570);
and U2751 (N_2751,N_1874,N_2035);
nor U2752 (N_2752,N_1957,N_148);
nor U2753 (N_2753,N_1074,N_78);
and U2754 (N_2754,N_785,N_1985);
nand U2755 (N_2755,N_791,N_1101);
or U2756 (N_2756,N_947,N_1239);
nor U2757 (N_2757,N_1718,N_1507);
or U2758 (N_2758,N_2303,N_2274);
or U2759 (N_2759,N_25,N_2271);
or U2760 (N_2760,N_2395,N_231);
or U2761 (N_2761,N_1333,N_2260);
nor U2762 (N_2762,N_2280,N_1719);
nand U2763 (N_2763,N_530,N_1383);
nand U2764 (N_2764,N_214,N_1252);
or U2765 (N_2765,N_383,N_2207);
or U2766 (N_2766,N_1409,N_1456);
or U2767 (N_2767,N_1104,N_892);
and U2768 (N_2768,N_2488,N_1893);
and U2769 (N_2769,N_1114,N_2230);
nor U2770 (N_2770,N_556,N_576);
or U2771 (N_2771,N_2443,N_1618);
and U2772 (N_2772,N_250,N_258);
and U2773 (N_2773,N_1531,N_30);
or U2774 (N_2774,N_628,N_1854);
or U2775 (N_2775,N_2200,N_584);
or U2776 (N_2776,N_2066,N_2047);
xor U2777 (N_2777,N_1544,N_1349);
or U2778 (N_2778,N_432,N_1441);
nand U2779 (N_2779,N_1758,N_1907);
and U2780 (N_2780,N_2023,N_912);
nand U2781 (N_2781,N_531,N_2449);
or U2782 (N_2782,N_2494,N_1694);
nand U2783 (N_2783,N_1747,N_1284);
and U2784 (N_2784,N_218,N_2353);
or U2785 (N_2785,N_1490,N_1453);
and U2786 (N_2786,N_1064,N_583);
or U2787 (N_2787,N_120,N_2141);
nor U2788 (N_2788,N_702,N_1781);
nor U2789 (N_2789,N_446,N_645);
nand U2790 (N_2790,N_2272,N_873);
nand U2791 (N_2791,N_1973,N_187);
nor U2792 (N_2792,N_244,N_1281);
or U2793 (N_2793,N_2072,N_952);
nand U2794 (N_2794,N_371,N_2355);
nand U2795 (N_2795,N_1304,N_2255);
or U2796 (N_2796,N_2124,N_1044);
nor U2797 (N_2797,N_2262,N_2094);
and U2798 (N_2798,N_573,N_1374);
xor U2799 (N_2799,N_591,N_2433);
xor U2800 (N_2800,N_1816,N_289);
or U2801 (N_2801,N_1852,N_1092);
nor U2802 (N_2802,N_1061,N_232);
or U2803 (N_2803,N_2425,N_2224);
or U2804 (N_2804,N_572,N_1886);
or U2805 (N_2805,N_67,N_104);
or U2806 (N_2806,N_739,N_2448);
and U2807 (N_2807,N_2107,N_978);
or U2808 (N_2808,N_753,N_759);
or U2809 (N_2809,N_737,N_2178);
nand U2810 (N_2810,N_32,N_221);
nand U2811 (N_2811,N_2116,N_851);
nand U2812 (N_2812,N_1545,N_1677);
or U2813 (N_2813,N_1288,N_68);
or U2814 (N_2814,N_1290,N_953);
nand U2815 (N_2815,N_1609,N_2252);
nor U2816 (N_2816,N_2194,N_1774);
nor U2817 (N_2817,N_131,N_637);
nor U2818 (N_2818,N_2450,N_1353);
nand U2819 (N_2819,N_374,N_599);
nor U2820 (N_2820,N_2462,N_884);
nor U2821 (N_2821,N_697,N_910);
nor U2822 (N_2822,N_1588,N_1974);
nor U2823 (N_2823,N_1978,N_1295);
and U2824 (N_2824,N_1124,N_299);
and U2825 (N_2825,N_1543,N_172);
nand U2826 (N_2826,N_2010,N_2022);
nor U2827 (N_2827,N_2181,N_1807);
nand U2828 (N_2828,N_618,N_667);
or U2829 (N_2829,N_1002,N_1425);
or U2830 (N_2830,N_878,N_2356);
nor U2831 (N_2831,N_2377,N_352);
or U2832 (N_2832,N_1316,N_1567);
nor U2833 (N_2833,N_1954,N_1745);
and U2834 (N_2834,N_2380,N_656);
nor U2835 (N_2835,N_1746,N_1813);
and U2836 (N_2836,N_1502,N_1553);
or U2837 (N_2837,N_960,N_1274);
nand U2838 (N_2838,N_580,N_1468);
nor U2839 (N_2839,N_2053,N_1947);
nor U2840 (N_2840,N_2161,N_770);
nand U2841 (N_2841,N_2267,N_265);
nor U2842 (N_2842,N_1840,N_1582);
nor U2843 (N_2843,N_1146,N_1939);
and U2844 (N_2844,N_1418,N_847);
and U2845 (N_2845,N_1597,N_1538);
nor U2846 (N_2846,N_1356,N_2083);
nand U2847 (N_2847,N_1525,N_1912);
nand U2848 (N_2848,N_1222,N_1296);
and U2849 (N_2849,N_474,N_2240);
nor U2850 (N_2850,N_309,N_558);
nor U2851 (N_2851,N_325,N_2275);
nand U2852 (N_2852,N_1380,N_1776);
and U2853 (N_2853,N_1678,N_128);
nand U2854 (N_2854,N_1657,N_1246);
nand U2855 (N_2855,N_210,N_834);
nor U2856 (N_2856,N_145,N_112);
or U2857 (N_2857,N_1078,N_1847);
or U2858 (N_2858,N_1406,N_123);
nor U2859 (N_2859,N_468,N_1532);
nor U2860 (N_2860,N_381,N_1370);
nor U2861 (N_2861,N_422,N_1098);
nand U2862 (N_2862,N_500,N_1873);
nor U2863 (N_2863,N_1477,N_1164);
or U2864 (N_2864,N_1756,N_2321);
and U2865 (N_2865,N_2316,N_262);
or U2866 (N_2866,N_2069,N_2416);
nor U2867 (N_2867,N_863,N_419);
or U2868 (N_2868,N_457,N_1233);
or U2869 (N_2869,N_2237,N_799);
nand U2870 (N_2870,N_2043,N_2489);
and U2871 (N_2871,N_842,N_220);
nor U2872 (N_2872,N_294,N_1128);
nand U2873 (N_2873,N_1149,N_263);
xnor U2874 (N_2874,N_922,N_1701);
or U2875 (N_2875,N_1900,N_44);
and U2876 (N_2876,N_442,N_2070);
nand U2877 (N_2877,N_2176,N_427);
and U2878 (N_2878,N_1075,N_938);
nor U2879 (N_2879,N_1911,N_877);
or U2880 (N_2880,N_611,N_226);
nor U2881 (N_2881,N_1503,N_485);
and U2882 (N_2882,N_241,N_855);
nand U2883 (N_2883,N_1669,N_1648);
nand U2884 (N_2884,N_1683,N_1244);
nor U2885 (N_2885,N_1172,N_414);
nor U2886 (N_2886,N_1264,N_1800);
nand U2887 (N_2887,N_2197,N_2330);
nand U2888 (N_2888,N_2285,N_2245);
or U2889 (N_2889,N_1635,N_678);
nor U2890 (N_2890,N_2193,N_194);
nand U2891 (N_2891,N_2305,N_607);
and U2892 (N_2892,N_1249,N_2382);
nor U2893 (N_2893,N_1598,N_2470);
or U2894 (N_2894,N_418,N_1231);
nand U2895 (N_2895,N_259,N_1696);
or U2896 (N_2896,N_1170,N_28);
nand U2897 (N_2897,N_2009,N_332);
nand U2898 (N_2898,N_1497,N_122);
and U2899 (N_2899,N_1500,N_516);
nor U2900 (N_2900,N_1315,N_2436);
nand U2901 (N_2901,N_2148,N_1668);
nor U2902 (N_2902,N_2423,N_1035);
and U2903 (N_2903,N_1625,N_893);
or U2904 (N_2904,N_1345,N_101);
nand U2905 (N_2905,N_1496,N_1710);
and U2906 (N_2906,N_936,N_1462);
or U2907 (N_2907,N_2348,N_2461);
nand U2908 (N_2908,N_165,N_2084);
and U2909 (N_2909,N_1563,N_1686);
or U2910 (N_2910,N_549,N_924);
and U2911 (N_2911,N_648,N_2307);
nand U2912 (N_2912,N_2059,N_1783);
nor U2913 (N_2913,N_1176,N_1824);
and U2914 (N_2914,N_1773,N_1310);
and U2915 (N_2915,N_2028,N_269);
or U2916 (N_2916,N_2362,N_2087);
and U2917 (N_2917,N_366,N_340);
nor U2918 (N_2918,N_92,N_578);
or U2919 (N_2919,N_1294,N_1229);
or U2920 (N_2920,N_1183,N_2037);
nor U2921 (N_2921,N_2326,N_1053);
and U2922 (N_2922,N_548,N_1883);
nand U2923 (N_2923,N_840,N_789);
nor U2924 (N_2924,N_1960,N_2140);
and U2925 (N_2925,N_200,N_1969);
or U2926 (N_2926,N_510,N_1550);
or U2927 (N_2927,N_2343,N_66);
or U2928 (N_2928,N_859,N_934);
nor U2929 (N_2929,N_717,N_1811);
nor U2930 (N_2930,N_2389,N_1944);
and U2931 (N_2931,N_1709,N_1988);
or U2932 (N_2932,N_692,N_1058);
nand U2933 (N_2933,N_1218,N_1548);
and U2934 (N_2934,N_475,N_180);
or U2935 (N_2935,N_80,N_1919);
nor U2936 (N_2936,N_2187,N_2300);
nand U2937 (N_2937,N_2399,N_267);
and U2938 (N_2938,N_1365,N_923);
and U2939 (N_2939,N_2306,N_720);
or U2940 (N_2940,N_2478,N_1242);
and U2941 (N_2941,N_575,N_1535);
nor U2942 (N_2942,N_2276,N_385);
or U2943 (N_2943,N_2096,N_2136);
and U2944 (N_2944,N_1154,N_1030);
nand U2945 (N_2945,N_23,N_159);
or U2946 (N_2946,N_1335,N_1923);
or U2947 (N_2947,N_1722,N_86);
nand U2948 (N_2948,N_2499,N_2457);
and U2949 (N_2949,N_2481,N_816);
or U2950 (N_2950,N_1762,N_1470);
and U2951 (N_2951,N_1426,N_2073);
and U2952 (N_2952,N_1742,N_480);
or U2953 (N_2953,N_2130,N_1188);
nand U2954 (N_2954,N_1903,N_1473);
or U2955 (N_2955,N_193,N_288);
and U2956 (N_2956,N_149,N_1660);
nand U2957 (N_2957,N_567,N_1921);
or U2958 (N_2958,N_1449,N_760);
or U2959 (N_2959,N_949,N_689);
and U2960 (N_2960,N_1454,N_404);
nand U2961 (N_2961,N_915,N_2400);
nor U2962 (N_2962,N_694,N_2368);
or U2963 (N_2963,N_76,N_503);
nor U2964 (N_2964,N_2404,N_646);
and U2965 (N_2965,N_2319,N_9);
and U2966 (N_2966,N_945,N_177);
or U2967 (N_2967,N_1126,N_658);
nand U2968 (N_2968,N_362,N_1077);
nor U2969 (N_2969,N_1279,N_1918);
nor U2970 (N_2970,N_1516,N_1072);
and U2971 (N_2971,N_4,N_1993);
nand U2972 (N_2972,N_1836,N_1994);
xor U2973 (N_2973,N_1699,N_603);
nand U2974 (N_2974,N_1880,N_1775);
xnor U2975 (N_2975,N_229,N_16);
nand U2976 (N_2976,N_1434,N_2150);
nor U2977 (N_2977,N_1666,N_1619);
nor U2978 (N_2978,N_392,N_866);
or U2979 (N_2979,N_1693,N_1850);
nor U2980 (N_2980,N_509,N_2282);
and U2981 (N_2981,N_1623,N_96);
nor U2982 (N_2982,N_768,N_515);
and U2983 (N_2983,N_1705,N_1320);
or U2984 (N_2984,N_1595,N_1757);
nor U2985 (N_2985,N_905,N_77);
nand U2986 (N_2986,N_967,N_696);
nor U2987 (N_2987,N_763,N_690);
or U2988 (N_2988,N_566,N_1391);
nor U2989 (N_2989,N_2220,N_1814);
nor U2990 (N_2990,N_2244,N_382);
or U2991 (N_2991,N_674,N_1050);
nor U2992 (N_2992,N_941,N_11);
or U2993 (N_2993,N_2317,N_469);
nor U2994 (N_2994,N_862,N_511);
or U2995 (N_2995,N_1005,N_1214);
or U2996 (N_2996,N_542,N_1366);
and U2997 (N_2997,N_293,N_755);
nand U2998 (N_2998,N_639,N_1572);
nand U2999 (N_2999,N_1429,N_1889);
or U3000 (N_3000,N_812,N_358);
and U3001 (N_3001,N_849,N_2138);
and U3002 (N_3002,N_869,N_1070);
nand U3003 (N_3003,N_843,N_787);
nor U3004 (N_3004,N_2027,N_2341);
nand U3005 (N_3005,N_1788,N_219);
or U3006 (N_3006,N_1634,N_2151);
and U3007 (N_3007,N_1809,N_2487);
or U3008 (N_3008,N_740,N_2020);
nor U3009 (N_3009,N_1556,N_1166);
nor U3010 (N_3010,N_911,N_505);
or U3011 (N_3011,N_240,N_1581);
and U3012 (N_3012,N_761,N_395);
nand U3013 (N_3013,N_1546,N_1224);
nor U3014 (N_3014,N_107,N_1573);
nor U3015 (N_3015,N_396,N_2256);
or U3016 (N_3016,N_773,N_355);
nand U3017 (N_3017,N_13,N_1300);
nor U3018 (N_3018,N_1822,N_1265);
nor U3019 (N_3019,N_665,N_1626);
and U3020 (N_3020,N_1478,N_919);
or U3021 (N_3021,N_389,N_2226);
nor U3022 (N_3022,N_514,N_1272);
nand U3023 (N_3023,N_1890,N_2381);
and U3024 (N_3024,N_1703,N_1768);
nor U3025 (N_3025,N_1471,N_135);
and U3026 (N_3026,N_2135,N_749);
nand U3027 (N_3027,N_2172,N_944);
or U3028 (N_3028,N_370,N_2295);
nor U3029 (N_3029,N_811,N_2229);
nand U3030 (N_3030,N_1793,N_1631);
and U3031 (N_3031,N_47,N_1839);
and U3032 (N_3032,N_2331,N_2195);
or U3033 (N_3033,N_188,N_426);
and U3034 (N_3034,N_1489,N_2251);
or U3035 (N_3035,N_545,N_2403);
nor U3036 (N_3036,N_1054,N_1830);
nand U3037 (N_3037,N_1899,N_1559);
nand U3038 (N_3038,N_1139,N_2065);
or U3039 (N_3039,N_2045,N_605);
nor U3040 (N_3040,N_541,N_380);
nand U3041 (N_3041,N_2479,N_1946);
and U3042 (N_3042,N_2142,N_1133);
and U3043 (N_3043,N_216,N_560);
nand U3044 (N_3044,N_617,N_2081);
nand U3045 (N_3045,N_538,N_631);
nand U3046 (N_3046,N_2050,N_867);
nand U3047 (N_3047,N_1965,N_992);
or U3048 (N_3048,N_1875,N_1346);
and U3049 (N_3049,N_1726,N_1105);
or U3050 (N_3050,N_2266,N_935);
nand U3051 (N_3051,N_471,N_2498);
or U3052 (N_3052,N_2328,N_1602);
and U3053 (N_3053,N_1460,N_502);
nand U3054 (N_3054,N_160,N_99);
nor U3055 (N_3055,N_2014,N_1400);
and U3056 (N_3056,N_1385,N_974);
or U3057 (N_3057,N_585,N_1179);
nor U3058 (N_3058,N_595,N_127);
and U3059 (N_3059,N_178,N_2432);
nor U3060 (N_3060,N_175,N_1601);
and U3061 (N_3061,N_1853,N_2253);
nor U3062 (N_3062,N_87,N_12);
or U3063 (N_3063,N_727,N_896);
nor U3064 (N_3064,N_1240,N_824);
and U3065 (N_3065,N_778,N_1180);
and U3066 (N_3066,N_902,N_844);
and U3067 (N_3067,N_307,N_2338);
nand U3068 (N_3068,N_1488,N_723);
nand U3069 (N_3069,N_762,N_413);
or U3070 (N_3070,N_1398,N_2199);
and U3071 (N_3071,N_623,N_2204);
or U3072 (N_3072,N_2218,N_1810);
and U3073 (N_3073,N_1205,N_2075);
nor U3074 (N_3074,N_7,N_212);
nor U3075 (N_3075,N_447,N_1143);
and U3076 (N_3076,N_996,N_476);
or U3077 (N_3077,N_1512,N_564);
and U3078 (N_3078,N_998,N_100);
nand U3079 (N_3079,N_1163,N_184);
or U3080 (N_3080,N_1129,N_1941);
or U3081 (N_3081,N_1867,N_146);
and U3082 (N_3082,N_1797,N_1175);
nor U3083 (N_3083,N_1733,N_1887);
nand U3084 (N_3084,N_858,N_185);
nor U3085 (N_3085,N_677,N_1079);
nand U3086 (N_3086,N_1616,N_1691);
and U3087 (N_3087,N_1041,N_2052);
nor U3088 (N_3088,N_2491,N_806);
nor U3089 (N_3089,N_1029,N_1379);
or U3090 (N_3090,N_871,N_2164);
or U3091 (N_3091,N_206,N_437);
nand U3092 (N_3092,N_527,N_2225);
and U3093 (N_3093,N_2036,N_168);
or U3094 (N_3094,N_1162,N_1120);
or U3095 (N_3095,N_2451,N_794);
nand U3096 (N_3096,N_1720,N_189);
nor U3097 (N_3097,N_608,N_673);
nor U3098 (N_3098,N_2011,N_2041);
and U3099 (N_3099,N_1818,N_455);
and U3100 (N_3100,N_587,N_2211);
or U3101 (N_3101,N_640,N_913);
or U3102 (N_3102,N_95,N_331);
nor U3103 (N_3103,N_2435,N_176);
or U3104 (N_3104,N_2082,N_452);
or U3105 (N_3105,N_2079,N_571);
and U3106 (N_3106,N_635,N_2004);
and U3107 (N_3107,N_330,N_273);
nor U3108 (N_3108,N_406,N_661);
nand U3109 (N_3109,N_10,N_103);
nand U3110 (N_3110,N_296,N_1439);
or U3111 (N_3111,N_1908,N_456);
and U3112 (N_3112,N_2097,N_1055);
or U3113 (N_3113,N_1906,N_88);
nor U3114 (N_3114,N_1526,N_543);
nand U3115 (N_3115,N_1697,N_828);
nand U3116 (N_3116,N_574,N_984);
or U3117 (N_3117,N_712,N_85);
or U3118 (N_3118,N_1317,N_881);
nand U3119 (N_3119,N_461,N_2205);
and U3120 (N_3120,N_1065,N_1990);
and U3121 (N_3121,N_813,N_213);
and U3122 (N_3122,N_173,N_1608);
or U3123 (N_3123,N_1245,N_874);
nor U3124 (N_3124,N_2269,N_1735);
nor U3125 (N_3125,N_1006,N_1178);
and U3126 (N_3126,N_1191,N_182);
nor U3127 (N_3127,N_1772,N_1981);
nor U3128 (N_3128,N_1832,N_2203);
or U3129 (N_3129,N_2455,N_79);
xor U3130 (N_3130,N_781,N_2119);
or U3131 (N_3131,N_650,N_140);
or U3132 (N_3132,N_279,N_237);
or U3133 (N_3133,N_1675,N_592);
nor U3134 (N_3134,N_792,N_52);
or U3135 (N_3135,N_728,N_1212);
nand U3136 (N_3136,N_322,N_2250);
and U3137 (N_3137,N_1979,N_451);
or U3138 (N_3138,N_1633,N_1465);
nor U3139 (N_3139,N_1967,N_2486);
and U3140 (N_3140,N_2,N_73);
or U3141 (N_3141,N_1665,N_1823);
nand U3142 (N_3142,N_2201,N_326);
nor U3143 (N_3143,N_1909,N_1494);
nand U3144 (N_3144,N_119,N_1671);
nand U3145 (N_3145,N_1637,N_1741);
nor U3146 (N_3146,N_137,N_1415);
and U3147 (N_3147,N_303,N_2146);
or U3148 (N_3148,N_43,N_1263);
and U3149 (N_3149,N_1071,N_839);
nand U3150 (N_3150,N_2227,N_198);
or U3151 (N_3151,N_2223,N_552);
nor U3152 (N_3152,N_497,N_415);
nand U3153 (N_3153,N_1584,N_2108);
or U3154 (N_3154,N_711,N_1225);
and U3155 (N_3155,N_1040,N_532);
nor U3156 (N_3156,N_793,N_1248);
nand U3157 (N_3157,N_1790,N_1377);
or U3158 (N_3158,N_2264,N_1256);
nand U3159 (N_3159,N_1732,N_1226);
or U3160 (N_3160,N_2074,N_1194);
or U3161 (N_3161,N_1291,N_1642);
nor U3162 (N_3162,N_1607,N_2149);
and U3163 (N_3163,N_983,N_1293);
or U3164 (N_3164,N_144,N_1336);
or U3165 (N_3165,N_320,N_2249);
and U3166 (N_3166,N_1151,N_72);
nand U3167 (N_3167,N_169,N_1848);
or U3168 (N_3168,N_886,N_968);
or U3169 (N_3169,N_920,N_2017);
nand U3170 (N_3170,N_1297,N_2236);
nand U3171 (N_3171,N_823,N_394);
nor U3172 (N_3172,N_1932,N_2143);
or U3173 (N_3173,N_721,N_2387);
and U3174 (N_3174,N_2391,N_1413);
nand U3175 (N_3175,N_1028,N_822);
and U3176 (N_3176,N_436,N_1842);
nor U3177 (N_3177,N_706,N_412);
nor U3178 (N_3178,N_1680,N_1737);
and U3179 (N_3179,N_2370,N_818);
nand U3180 (N_3180,N_2033,N_671);
and U3181 (N_3181,N_416,N_1307);
nor U3182 (N_3182,N_2376,N_1445);
and U3183 (N_3183,N_1327,N_2000);
nor U3184 (N_3184,N_2221,N_133);
nand U3185 (N_3185,N_1324,N_290);
or U3186 (N_3186,N_1442,N_534);
and U3187 (N_3187,N_1645,N_420);
and U3188 (N_3188,N_1100,N_547);
or U3189 (N_3189,N_801,N_1977);
or U3190 (N_3190,N_490,N_1059);
nand U3191 (N_3191,N_1498,N_2412);
or U3192 (N_3192,N_1395,N_1217);
nor U3193 (N_3193,N_1655,N_1676);
nor U3194 (N_3194,N_1784,N_2342);
nand U3195 (N_3195,N_1986,N_1613);
nor U3196 (N_3196,N_1667,N_1463);
nor U3197 (N_3197,N_1016,N_40);
nand U3198 (N_3198,N_2242,N_5);
or U3199 (N_3199,N_1013,N_1707);
and U3200 (N_3200,N_1661,N_1329);
xnor U3201 (N_3201,N_1996,N_1902);
or U3202 (N_3202,N_304,N_1968);
nand U3203 (N_3203,N_1443,N_1348);
and U3204 (N_3204,N_1571,N_1330);
nor U3205 (N_3205,N_736,N_525);
nor U3206 (N_3206,N_478,N_1971);
or U3207 (N_3207,N_496,N_276);
nand U3208 (N_3208,N_615,N_464);
and U3209 (N_3209,N_1051,N_709);
and U3210 (N_3210,N_2235,N_1706);
nor U3211 (N_3211,N_1437,N_610);
or U3212 (N_3212,N_428,N_2123);
nor U3213 (N_3213,N_1656,N_1664);
and U3214 (N_3214,N_313,N_429);
nand U3215 (N_3215,N_292,N_1583);
or U3216 (N_3216,N_454,N_1213);
and U3217 (N_3217,N_1440,N_142);
nand U3218 (N_3218,N_440,N_1714);
or U3219 (N_3219,N_1787,N_14);
nor U3220 (N_3220,N_2458,N_1989);
nand U3221 (N_3221,N_1331,N_1802);
and U3222 (N_3222,N_410,N_1638);
and U3223 (N_3223,N_1924,N_1487);
nand U3224 (N_3224,N_2209,N_1966);
nand U3225 (N_3225,N_1698,N_889);
nor U3226 (N_3226,N_588,N_2323);
and U3227 (N_3227,N_2405,N_756);
nor U3228 (N_3228,N_2234,N_780);
nor U3229 (N_3229,N_891,N_581);
nand U3230 (N_3230,N_1080,N_174);
nor U3231 (N_3231,N_2438,N_1587);
or U3232 (N_3232,N_1632,N_2392);
or U3233 (N_3233,N_300,N_1730);
nand U3234 (N_3234,N_1515,N_1738);
and U3235 (N_3235,N_718,N_865);
nand U3236 (N_3236,N_1358,N_308);
xor U3237 (N_3237,N_1014,N_2460);
nand U3238 (N_3238,N_1486,N_1794);
and U3239 (N_3239,N_1131,N_2496);
nand U3240 (N_3240,N_1564,N_704);
or U3241 (N_3241,N_1568,N_668);
nor U3242 (N_3242,N_338,N_83);
nand U3243 (N_3243,N_1082,N_1600);
nand U3244 (N_3244,N_1278,N_2171);
nand U3245 (N_3245,N_2363,N_1458);
and U3246 (N_3246,N_1209,N_1628);
or U3247 (N_3247,N_2283,N_1804);
nor U3248 (N_3248,N_134,N_521);
nand U3249 (N_3249,N_1173,N_2198);
and U3250 (N_3250,N_1234,N_324);
or U3251 (N_3251,N_926,N_283);
and U3252 (N_3252,N_1045,N_439);
nand U3253 (N_3253,N_539,N_1640);
nand U3254 (N_3254,N_482,N_1935);
and U3255 (N_3255,N_431,N_33);
or U3256 (N_3256,N_141,N_807);
nand U3257 (N_3257,N_972,N_1594);
and U3258 (N_3258,N_345,N_2456);
or U3259 (N_3259,N_1257,N_1685);
or U3260 (N_3260,N_1396,N_379);
or U3261 (N_3261,N_2430,N_555);
and U3262 (N_3262,N_1427,N_102);
nand U3263 (N_3263,N_2060,N_2440);
xnor U3264 (N_3264,N_1558,N_1519);
or U3265 (N_3265,N_1926,N_1000);
or U3266 (N_3266,N_1270,N_204);
and U3267 (N_3267,N_341,N_321);
or U3268 (N_3268,N_663,N_928);
nand U3269 (N_3269,N_272,N_2078);
and U3270 (N_3270,N_63,N_491);
nor U3271 (N_3271,N_714,N_1032);
nor U3272 (N_3272,N_586,N_2031);
and U3273 (N_3273,N_2333,N_815);
nand U3274 (N_3274,N_208,N_990);
nor U3275 (N_3275,N_814,N_657);
or U3276 (N_3276,N_1795,N_666);
nand U3277 (N_3277,N_636,N_1043);
nand U3278 (N_3278,N_1649,N_459);
nor U3279 (N_3279,N_2427,N_1056);
or U3280 (N_3280,N_2129,N_1261);
nand U3281 (N_3281,N_1408,N_1734);
nand U3282 (N_3282,N_1090,N_2424);
or U3283 (N_3283,N_1267,N_2071);
nand U3284 (N_3284,N_1639,N_1715);
nand U3285 (N_3285,N_504,N_1036);
nand U3286 (N_3286,N_2160,N_1207);
and U3287 (N_3287,N_1158,N_2288);
nand U3288 (N_3288,N_925,N_536);
and U3289 (N_3289,N_703,N_513);
or U3290 (N_3290,N_1452,N_2063);
or U3291 (N_3291,N_1864,N_1885);
or U3292 (N_3292,N_275,N_310);
nand U3293 (N_3293,N_2015,N_613);
or U3294 (N_3294,N_1540,N_22);
or U3295 (N_3295,N_45,N_215);
or U3296 (N_3296,N_378,N_879);
and U3297 (N_3297,N_1360,N_1397);
or U3298 (N_3298,N_39,N_8);
or U3299 (N_3299,N_2476,N_2085);
nand U3300 (N_3300,N_986,N_1455);
nor U3301 (N_3301,N_764,N_2162);
nor U3302 (N_3302,N_278,N_1375);
or U3303 (N_3303,N_779,N_1870);
and U3304 (N_3304,N_1679,N_1201);
nand U3305 (N_3305,N_1480,N_2334);
nand U3306 (N_3306,N_1312,N_523);
nor U3307 (N_3307,N_2243,N_676);
nand U3308 (N_3308,N_1087,N_2360);
and U3309 (N_3309,N_138,N_2469);
nor U3310 (N_3310,N_590,N_1421);
or U3311 (N_3311,N_1447,N_1165);
nor U3312 (N_3312,N_991,N_20);
or U3313 (N_3313,N_1389,N_1042);
nand U3314 (N_3314,N_334,N_1658);
and U3315 (N_3315,N_2429,N_2110);
and U3316 (N_3316,N_643,N_1785);
and U3317 (N_3317,N_827,N_393);
and U3318 (N_3318,N_833,N_1940);
nor U3319 (N_3319,N_2354,N_115);
and U3320 (N_3320,N_1401,N_2313);
nand U3321 (N_3321,N_1376,N_1766);
or U3322 (N_3322,N_1792,N_1328);
or U3323 (N_3323,N_444,N_466);
and U3324 (N_3324,N_1736,N_2325);
nor U3325 (N_3325,N_1093,N_1569);
and U3326 (N_3326,N_1081,N_742);
or U3327 (N_3327,N_932,N_225);
or U3328 (N_3328,N_391,N_2182);
and U3329 (N_3329,N_746,N_649);
nand U3330 (N_3330,N_620,N_153);
nor U3331 (N_3331,N_1253,N_171);
nand U3332 (N_3332,N_2021,N_1901);
and U3333 (N_3333,N_1915,N_2086);
nor U3334 (N_3334,N_264,N_1309);
or U3335 (N_3335,N_157,N_2411);
nand U3336 (N_3336,N_55,N_1202);
nor U3337 (N_3337,N_2434,N_568);
and U3338 (N_3338,N_1765,N_1862);
nor U3339 (N_3339,N_1118,N_880);
and U3340 (N_3340,N_1704,N_1860);
or U3341 (N_3341,N_318,N_1204);
nor U3342 (N_3342,N_1057,N_357);
nor U3343 (N_3343,N_1869,N_2344);
or U3344 (N_3344,N_1711,N_725);
or U3345 (N_3345,N_257,N_1021);
nand U3346 (N_3346,N_458,N_1821);
or U3347 (N_3347,N_644,N_2375);
or U3348 (N_3348,N_1210,N_1008);
or U3349 (N_3349,N_425,N_2241);
nand U3350 (N_3350,N_2299,N_596);
nor U3351 (N_3351,N_2485,N_390);
nor U3352 (N_3352,N_2336,N_1459);
and U3353 (N_3353,N_2068,N_2308);
and U3354 (N_3354,N_561,N_376);
nor U3355 (N_3355,N_1517,N_1876);
nor U3356 (N_3356,N_1198,N_2144);
or U3357 (N_3357,N_887,N_1227);
nand U3358 (N_3358,N_750,N_738);
and U3359 (N_3359,N_885,N_158);
and U3360 (N_3360,N_1963,N_2294);
nor U3361 (N_3361,N_1184,N_301);
nor U3362 (N_3362,N_2401,N_2180);
nor U3363 (N_3363,N_528,N_876);
or U3364 (N_3364,N_2361,N_638);
nand U3365 (N_3365,N_274,N_1700);
nand U3366 (N_3366,N_1364,N_2428);
nor U3367 (N_3367,N_1339,N_1052);
nand U3368 (N_3368,N_829,N_1702);
nand U3369 (N_3369,N_748,N_907);
and U3370 (N_3370,N_268,N_675);
nor U3371 (N_3371,N_751,N_2206);
or U3372 (N_3372,N_435,N_349);
and U3373 (N_3373,N_1230,N_1168);
or U3374 (N_3374,N_626,N_1586);
and U3375 (N_3375,N_601,N_852);
nand U3376 (N_3376,N_82,N_1405);
nand U3377 (N_3377,N_291,N_2030);
nor U3378 (N_3378,N_1857,N_2006);
or U3379 (N_3379,N_1402,N_1539);
nor U3380 (N_3380,N_1936,N_775);
nor U3381 (N_3381,N_964,N_2452);
nor U3382 (N_3382,N_1589,N_1829);
or U3383 (N_3383,N_1561,N_139);
and U3384 (N_3384,N_93,N_316);
and U3385 (N_3385,N_1289,N_1764);
nand U3386 (N_3386,N_2046,N_2170);
nand U3387 (N_3387,N_1599,N_2371);
nor U3388 (N_3388,N_1018,N_49);
or U3389 (N_3389,N_233,N_217);
or U3390 (N_3390,N_2263,N_2238);
nor U3391 (N_3391,N_2365,N_1352);
nand U3392 (N_3392,N_2402,N_1235);
nand U3393 (N_3393,N_2369,N_1067);
nand U3394 (N_3394,N_1951,N_2477);
or U3395 (N_3395,N_161,N_126);
nand U3396 (N_3396,N_2386,N_512);
nand U3397 (N_3397,N_970,N_2159);
nor U3398 (N_3398,N_347,N_1436);
nand U3399 (N_3399,N_2383,N_1298);
and U3400 (N_3400,N_1808,N_1731);
and U3401 (N_3401,N_2179,N_1580);
nor U3402 (N_3402,N_1277,N_1378);
and U3403 (N_3403,N_1752,N_2393);
nand U3404 (N_3404,N_409,N_353);
or U3405 (N_3405,N_2088,N_6);
nand U3406 (N_3406,N_2349,N_1948);
and U3407 (N_3407,N_2026,N_2133);
nor U3408 (N_3408,N_1369,N_155);
nor U3409 (N_3409,N_2459,N_1147);
and U3410 (N_3410,N_1363,N_550);
nand U3411 (N_3411,N_60,N_1341);
nor U3412 (N_3412,N_1048,N_1313);
and U3413 (N_3413,N_1461,N_1492);
and U3414 (N_3414,N_625,N_2394);
nor U3415 (N_3415,N_228,N_1777);
and U3416 (N_3416,N_2286,N_2092);
nor U3417 (N_3417,N_888,N_1771);
nor U3418 (N_3418,N_2324,N_1189);
nor U3419 (N_3419,N_664,N_1109);
and U3420 (N_3420,N_1913,N_745);
or U3421 (N_3421,N_733,N_1182);
and U3422 (N_3422,N_1761,N_1390);
nand U3423 (N_3423,N_2340,N_2147);
nor U3424 (N_3424,N_298,N_484);
and U3425 (N_3425,N_2468,N_403);
nand U3426 (N_3426,N_1012,N_1689);
nor U3427 (N_3427,N_411,N_1605);
and U3428 (N_3428,N_1302,N_942);
nor U3429 (N_3429,N_2183,N_1624);
nor U3430 (N_3430,N_988,N_836);
nand U3431 (N_3431,N_498,N_1387);
or U3432 (N_3432,N_1010,N_287);
or U3433 (N_3433,N_2373,N_1828);
and U3434 (N_3434,N_908,N_1566);
nor U3435 (N_3435,N_1196,N_600);
or U3436 (N_3436,N_1318,N_1221);
nand U3437 (N_3437,N_795,N_1557);
and U3438 (N_3438,N_342,N_734);
nand U3439 (N_3439,N_445,N_1843);
or U3440 (N_3440,N_956,N_621);
or U3441 (N_3441,N_629,N_1905);
and U3442 (N_3442,N_2228,N_2077);
and U3443 (N_3443,N_2122,N_1325);
or U3444 (N_3444,N_2472,N_2265);
nor U3445 (N_3445,N_1483,N_1481);
or U3446 (N_3446,N_508,N_861);
nand U3447 (N_3447,N_1513,N_1174);
and U3448 (N_3448,N_2426,N_864);
nand U3449 (N_3449,N_982,N_1806);
nor U3450 (N_3450,N_170,N_433);
nor U3451 (N_3451,N_2454,N_708);
and U3452 (N_3452,N_2374,N_2093);
nand U3453 (N_3453,N_1135,N_2214);
nand U3454 (N_3454,N_845,N_1292);
and U3455 (N_3455,N_1153,N_2222);
and U3456 (N_3456,N_2057,N_2483);
and U3457 (N_3457,N_767,N_254);
or U3458 (N_3458,N_2257,N_1083);
and U3459 (N_3459,N_2005,N_2013);
or U3460 (N_3460,N_1276,N_1251);
or U3461 (N_3461,N_940,N_344);
nor U3462 (N_3462,N_1354,N_1386);
or U3463 (N_3463,N_747,N_2125);
and U3464 (N_3464,N_1673,N_166);
or U3465 (N_3465,N_1520,N_1552);
or U3466 (N_3466,N_1956,N_735);
or U3467 (N_3467,N_1791,N_2439);
nor U3468 (N_3468,N_470,N_1160);
or U3469 (N_3469,N_699,N_1422);
or U3470 (N_3470,N_98,N_377);
or U3471 (N_3471,N_965,N_2410);
nor U3472 (N_3472,N_1615,N_38);
and U3473 (N_3473,N_966,N_872);
and U3474 (N_3474,N_2384,N_2372);
and U3475 (N_3475,N_2270,N_486);
and U3476 (N_3476,N_130,N_951);
nor U3477 (N_3477,N_846,N_2309);
or U3478 (N_3478,N_230,N_831);
xnor U3479 (N_3479,N_989,N_997);
or U3480 (N_3480,N_1801,N_802);
nor U3481 (N_3481,N_398,N_579);
nor U3482 (N_3482,N_2298,N_790);
nor U3483 (N_3483,N_2121,N_2480);
and U3484 (N_3484,N_31,N_19);
nand U3485 (N_3485,N_34,N_1740);
nor U3486 (N_3486,N_84,N_2104);
or U3487 (N_3487,N_367,N_1269);
and U3488 (N_3488,N_26,N_2495);
or U3489 (N_3489,N_1937,N_408);
or U3490 (N_3490,N_453,N_788);
or U3491 (N_3491,N_987,N_438);
and U3492 (N_3492,N_1099,N_994);
nand U3493 (N_3493,N_1511,N_125);
and U3494 (N_3494,N_507,N_715);
or U3495 (N_3495,N_1931,N_557);
or U3496 (N_3496,N_2239,N_1652);
nand U3497 (N_3497,N_1115,N_401);
and U3498 (N_3498,N_2445,N_825);
and U3499 (N_3499,N_959,N_832);
or U3500 (N_3500,N_995,N_1308);
and U3501 (N_3501,N_904,N_757);
and U3502 (N_3502,N_1122,N_1897);
nor U3503 (N_3503,N_1961,N_59);
and U3504 (N_3504,N_506,N_655);
and U3505 (N_3505,N_1141,N_670);
or U3506 (N_3506,N_1878,N_1321);
and U3507 (N_3507,N_1743,N_1475);
nand U3508 (N_3508,N_1351,N_1144);
xor U3509 (N_3509,N_179,N_1684);
nor U3510 (N_3510,N_1236,N_2155);
or U3511 (N_3511,N_2067,N_1384);
nand U3512 (N_3512,N_804,N_2213);
or U3513 (N_3513,N_1976,N_1695);
nand U3514 (N_3514,N_1411,N_261);
nor U3515 (N_3515,N_2318,N_1322);
or U3516 (N_3516,N_2281,N_473);
or U3517 (N_3517,N_1681,N_124);
nand U3518 (N_3518,N_688,N_1009);
nand U3519 (N_3519,N_460,N_417);
or U3520 (N_3520,N_2441,N_1570);
nor U3521 (N_3521,N_1610,N_2278);
nor U3522 (N_3522,N_111,N_1920);
or U3523 (N_3523,N_868,N_633);
and U3524 (N_3524,N_2202,N_2007);
nand U3525 (N_3525,N_1641,N_1412);
or U3526 (N_3526,N_1084,N_1076);
or U3527 (N_3527,N_2464,N_1984);
and U3528 (N_3528,N_1861,N_826);
and U3529 (N_3529,N_796,N_2158);
or U3530 (N_3530,N_805,N_777);
xor U3531 (N_3531,N_540,N_1992);
or U3532 (N_3532,N_1997,N_1837);
nand U3533 (N_3533,N_1952,N_1049);
nand U3534 (N_3534,N_2114,N_1467);
nand U3535 (N_3535,N_1780,N_1604);
and U3536 (N_3536,N_691,N_2113);
and U3537 (N_3537,N_1528,N_2231);
and U3538 (N_3538,N_1708,N_2032);
or U3539 (N_3539,N_1560,N_1299);
or U3540 (N_3540,N_129,N_295);
or U3541 (N_3541,N_1798,N_963);
nand U3542 (N_3542,N_205,N_197);
and U3543 (N_3543,N_1334,N_2117);
and U3544 (N_3544,N_224,N_1687);
and U3545 (N_3545,N_337,N_1303);
or U3546 (N_3546,N_1565,N_448);
and U3547 (N_3547,N_909,N_2492);
nand U3548 (N_3548,N_2100,N_1112);
or U3549 (N_3549,N_1537,N_918);
and U3550 (N_3550,N_533,N_2167);
or U3551 (N_3551,N_424,N_327);
nand U3552 (N_3552,N_384,N_1805);
and U3553 (N_3553,N_713,N_1827);
nor U3554 (N_3554,N_1914,N_1020);
and U3555 (N_3555,N_654,N_1123);
nand U3556 (N_3556,N_333,N_1420);
and U3557 (N_3557,N_1472,N_895);
nor U3558 (N_3558,N_1219,N_553);
or U3559 (N_3559,N_2312,N_467);
nor U3560 (N_3560,N_1069,N_2329);
or U3561 (N_3561,N_373,N_1476);
nand U3562 (N_3562,N_662,N_256);
nand U3563 (N_3563,N_2490,N_772);
or U3564 (N_3564,N_319,N_1922);
nand U3565 (N_3565,N_2157,N_2062);
and U3566 (N_3566,N_2259,N_927);
nand U3567 (N_3567,N_2315,N_1474);
or U3568 (N_3568,N_191,N_758);
nor U3569 (N_3569,N_1820,N_848);
and U3570 (N_3570,N_2049,N_937);
and U3571 (N_3571,N_242,N_1403);
nand U3572 (N_3572,N_1501,N_526);
nor U3573 (N_3573,N_1430,N_90);
nor U3574 (N_3574,N_372,N_255);
nand U3575 (N_3575,N_1845,N_2304);
and U3576 (N_3576,N_260,N_407);
nor U3577 (N_3577,N_2279,N_719);
nor U3578 (N_3578,N_679,N_2453);
nand U3579 (N_3579,N_1534,N_2219);
or U3580 (N_3580,N_1062,N_253);
or U3581 (N_3581,N_1268,N_2482);
nand U3582 (N_3582,N_1361,N_387);
nor U3583 (N_3583,N_1763,N_183);
nor U3584 (N_3584,N_1485,N_817);
nor U3585 (N_3585,N_1499,N_368);
nor U3586 (N_3586,N_1622,N_2442);
or U3587 (N_3587,N_1575,N_943);
or U3588 (N_3588,N_535,N_1414);
or U3589 (N_3589,N_776,N_1692);
nor U3590 (N_3590,N_463,N_1088);
or U3591 (N_3591,N_1491,N_477);
nand U3592 (N_3592,N_1208,N_1554);
and U3593 (N_3593,N_1717,N_2064);
or U3594 (N_3594,N_1003,N_1958);
or U3595 (N_3595,N_1950,N_2008);
and U3596 (N_3596,N_1431,N_356);
nand U3597 (N_3597,N_2191,N_1286);
or U3598 (N_3598,N_364,N_495);
or U3599 (N_3599,N_1627,N_1521);
or U3600 (N_3600,N_1206,N_1577);
and U3601 (N_3601,N_2232,N_1096);
or U3602 (N_3602,N_1392,N_820);
or U3603 (N_3603,N_2357,N_1280);
xor U3604 (N_3604,N_630,N_606);
and U3605 (N_3605,N_2153,N_771);
and U3606 (N_3606,N_1606,N_1254);
nand U3607 (N_3607,N_1195,N_898);
and U3608 (N_3608,N_1593,N_1381);
and U3609 (N_3609,N_683,N_1508);
nor U3610 (N_3610,N_1247,N_1399);
nor U3611 (N_3611,N_2145,N_2390);
nand U3612 (N_3612,N_2310,N_328);
and U3613 (N_3613,N_1929,N_1023);
nor U3614 (N_3614,N_1879,N_1611);
and U3615 (N_3615,N_117,N_1547);
nor U3616 (N_3616,N_1851,N_2246);
or U3617 (N_3617,N_680,N_782);
nand U3618 (N_3618,N_181,N_2339);
or U3619 (N_3619,N_1142,N_162);
nor U3620 (N_3620,N_386,N_1894);
nor U3621 (N_3621,N_2366,N_1134);
and U3622 (N_3622,N_2493,N_1258);
and U3623 (N_3623,N_1111,N_1509);
or U3624 (N_3624,N_1662,N_2024);
nor U3625 (N_3625,N_2247,N_518);
and U3626 (N_3626,N_280,N_1404);
nor U3627 (N_3627,N_2115,N_1250);
nand U3628 (N_3628,N_1749,N_1982);
xor U3629 (N_3629,N_132,N_423);
nand U3630 (N_3630,N_2152,N_186);
and U3631 (N_3631,N_1215,N_1451);
and U3632 (N_3632,N_1089,N_443);
nor U3633 (N_3633,N_2379,N_1148);
and U3634 (N_3634,N_1562,N_1156);
and U3635 (N_3635,N_65,N_1260);
nor U3636 (N_3636,N_1769,N_2105);
nor U3637 (N_3637,N_234,N_1964);
nand U3638 (N_3638,N_91,N_2284);
nor U3639 (N_3639,N_2358,N_1782);
nor U3640 (N_3640,N_1,N_70);
or U3641 (N_3641,N_1446,N_2163);
nand U3642 (N_3642,N_1306,N_1592);
and U3643 (N_3643,N_766,N_1495);
nand U3644 (N_3644,N_50,N_1803);
and U3645 (N_3645,N_106,N_1015);
nand U3646 (N_3646,N_798,N_2177);
nand U3647 (N_3647,N_1457,N_2168);
or U3648 (N_3648,N_2397,N_1955);
nor U3649 (N_3649,N_687,N_685);
nor U3650 (N_3650,N_2345,N_1796);
nand U3651 (N_3651,N_2169,N_1161);
and U3652 (N_3652,N_1759,N_487);
and U3653 (N_3653,N_1938,N_2212);
or U3654 (N_3654,N_2289,N_901);
and U3655 (N_3655,N_2175,N_1925);
and U3656 (N_3656,N_2444,N_1744);
nand U3657 (N_3657,N_2102,N_1882);
or U3658 (N_3658,N_207,N_1368);
nand U3659 (N_3659,N_335,N_1359);
or U3660 (N_3660,N_705,N_2277);
nand U3661 (N_3661,N_2327,N_113);
nand U3662 (N_3662,N_1285,N_2378);
nand U3663 (N_3663,N_2051,N_1962);
nand U3664 (N_3664,N_284,N_1103);
nor U3665 (N_3665,N_641,N_2351);
or U3666 (N_3666,N_41,N_537);
nand U3667 (N_3667,N_906,N_108);
nand U3668 (N_3668,N_2258,N_1983);
nand U3669 (N_3669,N_830,N_430);
xnor U3670 (N_3670,N_243,N_2001);
or U3671 (N_3671,N_449,N_1527);
nor U3672 (N_3672,N_329,N_1591);
nand U3673 (N_3673,N_1025,N_48);
or U3674 (N_3674,N_1350,N_1113);
nand U3675 (N_3675,N_1725,N_2166);
or U3676 (N_3676,N_1332,N_1482);
nand U3677 (N_3677,N_1617,N_786);
or U3678 (N_3678,N_1192,N_1728);
nand U3679 (N_3679,N_2447,N_2347);
nor U3680 (N_3680,N_562,N_402);
nor U3681 (N_3681,N_1262,N_2396);
or U3682 (N_3682,N_774,N_2089);
xor U3683 (N_3683,N_346,N_121);
and U3684 (N_3684,N_1690,N_1220);
or U3685 (N_3685,N_2090,N_612);
nand U3686 (N_3686,N_1877,N_1393);
nand U3687 (N_3687,N_1241,N_1834);
and U3688 (N_3688,N_2475,N_1004);
nor U3689 (N_3689,N_1311,N_2406);
nor U3690 (N_3690,N_546,N_2291);
nor U3691 (N_3691,N_700,N_29);
nor U3692 (N_3692,N_1275,N_1755);
and U3693 (N_3693,N_2210,N_1506);
or U3694 (N_3694,N_2233,N_235);
and U3695 (N_3695,N_1169,N_311);
or U3696 (N_3696,N_2297,N_977);
nor U3697 (N_3697,N_1713,N_1855);
nand U3698 (N_3698,N_2196,N_659);
and U3699 (N_3699,N_2287,N_1066);
nor U3700 (N_3700,N_1943,N_1674);
and U3701 (N_3701,N_434,N_2254);
nor U3702 (N_3702,N_803,N_1433);
or U3703 (N_3703,N_769,N_1646);
or U3704 (N_3704,N_598,N_105);
nand U3705 (N_3705,N_821,N_441);
and U3706 (N_3706,N_2061,N_707);
and U3707 (N_3707,N_2471,N_164);
nand U3708 (N_3708,N_1972,N_2467);
or U3709 (N_3709,N_2131,N_1841);
or U3710 (N_3710,N_365,N_1063);
nand U3711 (N_3711,N_2056,N_1670);
nor U3712 (N_3712,N_236,N_1999);
and U3713 (N_3713,N_1815,N_1193);
nand U3714 (N_3714,N_246,N_2446);
nand U3715 (N_3715,N_686,N_1888);
and U3716 (N_3716,N_143,N_1612);
or U3717 (N_3717,N_2273,N_1644);
and U3718 (N_3718,N_2039,N_1786);
nor U3719 (N_3719,N_897,N_1038);
and U3720 (N_3720,N_931,N_1739);
and U3721 (N_3721,N_2216,N_1347);
and U3722 (N_3722,N_317,N_354);
nor U3723 (N_3723,N_2111,N_722);
or U3724 (N_3724,N_957,N_1819);
and U3725 (N_3725,N_369,N_1975);
nand U3726 (N_3726,N_2076,N_2332);
nor U3727 (N_3727,N_27,N_2497);
and U3728 (N_3728,N_2268,N_752);
nor U3729 (N_3729,N_89,N_2302);
nand U3730 (N_3730,N_42,N_961);
or U3731 (N_3731,N_634,N_2337);
and U3732 (N_3732,N_2407,N_2415);
nor U3733 (N_3733,N_1273,N_1542);
nand U3734 (N_3734,N_2184,N_1760);
nor U3735 (N_3735,N_2095,N_71);
and U3736 (N_3736,N_397,N_1895);
nand U3737 (N_3737,N_2350,N_1603);
nand U3738 (N_3738,N_1444,N_1663);
nor U3739 (N_3739,N_693,N_593);
or U3740 (N_3740,N_167,N_1927);
and U3741 (N_3741,N_1232,N_2174);
nor U3742 (N_3742,N_2091,N_56);
nand U3743 (N_3743,N_315,N_1555);
nor U3744 (N_3744,N_1754,N_976);
nor U3745 (N_3745,N_870,N_1833);
nand U3746 (N_3746,N_2290,N_1337);
or U3747 (N_3747,N_1930,N_1228);
nand U3748 (N_3748,N_1672,N_939);
nand U3749 (N_3749,N_1107,N_1998);
nand U3750 (N_3750,N_853,N_1078);
nand U3751 (N_3751,N_2240,N_1156);
or U3752 (N_3752,N_1862,N_84);
nor U3753 (N_3753,N_687,N_726);
nor U3754 (N_3754,N_2058,N_1752);
xnor U3755 (N_3755,N_319,N_162);
nor U3756 (N_3756,N_1914,N_1179);
or U3757 (N_3757,N_958,N_2261);
or U3758 (N_3758,N_1804,N_551);
nand U3759 (N_3759,N_430,N_1872);
nand U3760 (N_3760,N_1663,N_92);
and U3761 (N_3761,N_201,N_2464);
nor U3762 (N_3762,N_81,N_959);
or U3763 (N_3763,N_1394,N_225);
nor U3764 (N_3764,N_2197,N_690);
and U3765 (N_3765,N_1592,N_2083);
or U3766 (N_3766,N_1999,N_1394);
nor U3767 (N_3767,N_335,N_2438);
nand U3768 (N_3768,N_1631,N_339);
or U3769 (N_3769,N_1033,N_2116);
nor U3770 (N_3770,N_292,N_223);
or U3771 (N_3771,N_2304,N_822);
and U3772 (N_3772,N_758,N_2323);
or U3773 (N_3773,N_2312,N_670);
and U3774 (N_3774,N_1369,N_570);
nand U3775 (N_3775,N_339,N_2241);
or U3776 (N_3776,N_1409,N_345);
and U3777 (N_3777,N_1177,N_1396);
or U3778 (N_3778,N_145,N_2466);
nand U3779 (N_3779,N_1668,N_1740);
or U3780 (N_3780,N_1607,N_1829);
or U3781 (N_3781,N_641,N_1972);
and U3782 (N_3782,N_1863,N_138);
nand U3783 (N_3783,N_1277,N_1314);
nor U3784 (N_3784,N_82,N_2426);
or U3785 (N_3785,N_4,N_1575);
nor U3786 (N_3786,N_1898,N_136);
nor U3787 (N_3787,N_246,N_1849);
nor U3788 (N_3788,N_257,N_2292);
xnor U3789 (N_3789,N_2103,N_588);
nand U3790 (N_3790,N_122,N_1982);
nand U3791 (N_3791,N_486,N_640);
nand U3792 (N_3792,N_71,N_1877);
nor U3793 (N_3793,N_278,N_1778);
nor U3794 (N_3794,N_245,N_971);
or U3795 (N_3795,N_1185,N_720);
and U3796 (N_3796,N_1727,N_942);
and U3797 (N_3797,N_757,N_1815);
or U3798 (N_3798,N_2350,N_726);
and U3799 (N_3799,N_962,N_1830);
nor U3800 (N_3800,N_796,N_10);
or U3801 (N_3801,N_963,N_1);
or U3802 (N_3802,N_1646,N_101);
nor U3803 (N_3803,N_1277,N_1889);
and U3804 (N_3804,N_1850,N_2057);
or U3805 (N_3805,N_508,N_2316);
nand U3806 (N_3806,N_1037,N_753);
and U3807 (N_3807,N_2049,N_2394);
or U3808 (N_3808,N_1468,N_927);
or U3809 (N_3809,N_306,N_1293);
nand U3810 (N_3810,N_1376,N_1608);
and U3811 (N_3811,N_510,N_1369);
or U3812 (N_3812,N_1937,N_1604);
or U3813 (N_3813,N_799,N_1522);
or U3814 (N_3814,N_1860,N_448);
nand U3815 (N_3815,N_1168,N_2488);
or U3816 (N_3816,N_1806,N_1547);
nor U3817 (N_3817,N_283,N_2005);
xor U3818 (N_3818,N_1490,N_1020);
nand U3819 (N_3819,N_354,N_1220);
and U3820 (N_3820,N_2154,N_1346);
nor U3821 (N_3821,N_1450,N_1301);
nor U3822 (N_3822,N_574,N_1315);
or U3823 (N_3823,N_266,N_955);
or U3824 (N_3824,N_2223,N_775);
nor U3825 (N_3825,N_2031,N_1419);
xnor U3826 (N_3826,N_2351,N_1758);
or U3827 (N_3827,N_592,N_1633);
nand U3828 (N_3828,N_754,N_1917);
and U3829 (N_3829,N_465,N_2062);
nor U3830 (N_3830,N_377,N_1120);
nor U3831 (N_3831,N_20,N_422);
nor U3832 (N_3832,N_2319,N_426);
nand U3833 (N_3833,N_19,N_2219);
or U3834 (N_3834,N_1870,N_1948);
and U3835 (N_3835,N_893,N_2158);
and U3836 (N_3836,N_739,N_21);
nand U3837 (N_3837,N_1744,N_2206);
and U3838 (N_3838,N_679,N_2347);
nor U3839 (N_3839,N_1686,N_2447);
and U3840 (N_3840,N_1449,N_1525);
nor U3841 (N_3841,N_1419,N_1819);
nor U3842 (N_3842,N_1760,N_796);
or U3843 (N_3843,N_649,N_1739);
nand U3844 (N_3844,N_1560,N_1692);
or U3845 (N_3845,N_792,N_762);
or U3846 (N_3846,N_1230,N_353);
and U3847 (N_3847,N_404,N_1461);
nand U3848 (N_3848,N_1592,N_2490);
nor U3849 (N_3849,N_1953,N_850);
and U3850 (N_3850,N_413,N_1395);
nor U3851 (N_3851,N_1363,N_873);
and U3852 (N_3852,N_1956,N_1401);
nand U3853 (N_3853,N_1643,N_415);
nor U3854 (N_3854,N_64,N_105);
nand U3855 (N_3855,N_1855,N_2112);
nor U3856 (N_3856,N_2375,N_1901);
nand U3857 (N_3857,N_1318,N_2181);
or U3858 (N_3858,N_2455,N_979);
nand U3859 (N_3859,N_1867,N_526);
nor U3860 (N_3860,N_304,N_2445);
and U3861 (N_3861,N_12,N_2336);
and U3862 (N_3862,N_1988,N_997);
and U3863 (N_3863,N_991,N_2156);
nor U3864 (N_3864,N_1944,N_355);
and U3865 (N_3865,N_2395,N_15);
nor U3866 (N_3866,N_809,N_1923);
nand U3867 (N_3867,N_1570,N_1165);
nor U3868 (N_3868,N_1810,N_559);
nor U3869 (N_3869,N_269,N_2165);
nand U3870 (N_3870,N_1390,N_597);
or U3871 (N_3871,N_143,N_1296);
or U3872 (N_3872,N_1580,N_256);
and U3873 (N_3873,N_2489,N_54);
nand U3874 (N_3874,N_100,N_1785);
nand U3875 (N_3875,N_860,N_842);
nand U3876 (N_3876,N_1643,N_1350);
nor U3877 (N_3877,N_1832,N_1757);
and U3878 (N_3878,N_2165,N_1627);
nor U3879 (N_3879,N_189,N_1789);
nand U3880 (N_3880,N_2440,N_1259);
or U3881 (N_3881,N_2207,N_238);
or U3882 (N_3882,N_1778,N_1060);
or U3883 (N_3883,N_2149,N_2278);
nand U3884 (N_3884,N_1906,N_623);
nand U3885 (N_3885,N_223,N_1577);
nor U3886 (N_3886,N_1775,N_358);
nand U3887 (N_3887,N_1589,N_2107);
and U3888 (N_3888,N_2333,N_1527);
nor U3889 (N_3889,N_1817,N_696);
and U3890 (N_3890,N_2010,N_1673);
or U3891 (N_3891,N_327,N_562);
nor U3892 (N_3892,N_1589,N_1907);
nand U3893 (N_3893,N_1962,N_647);
nand U3894 (N_3894,N_1773,N_2457);
and U3895 (N_3895,N_1431,N_458);
or U3896 (N_3896,N_1495,N_2444);
or U3897 (N_3897,N_2238,N_2234);
nor U3898 (N_3898,N_682,N_802);
nor U3899 (N_3899,N_393,N_724);
xor U3900 (N_3900,N_1172,N_997);
and U3901 (N_3901,N_2034,N_1587);
nor U3902 (N_3902,N_2330,N_721);
nand U3903 (N_3903,N_50,N_2448);
nand U3904 (N_3904,N_1293,N_986);
nor U3905 (N_3905,N_1439,N_1413);
and U3906 (N_3906,N_506,N_1835);
nor U3907 (N_3907,N_1952,N_524);
and U3908 (N_3908,N_267,N_405);
nand U3909 (N_3909,N_1633,N_650);
or U3910 (N_3910,N_2432,N_1585);
nand U3911 (N_3911,N_2453,N_962);
nor U3912 (N_3912,N_701,N_278);
nand U3913 (N_3913,N_600,N_786);
nand U3914 (N_3914,N_770,N_704);
nor U3915 (N_3915,N_1602,N_469);
nor U3916 (N_3916,N_430,N_2416);
or U3917 (N_3917,N_1571,N_1399);
or U3918 (N_3918,N_1196,N_1520);
and U3919 (N_3919,N_1658,N_2156);
nand U3920 (N_3920,N_516,N_2333);
or U3921 (N_3921,N_1990,N_2312);
or U3922 (N_3922,N_1855,N_672);
nor U3923 (N_3923,N_2038,N_865);
and U3924 (N_3924,N_541,N_391);
nor U3925 (N_3925,N_938,N_92);
and U3926 (N_3926,N_1453,N_2459);
and U3927 (N_3927,N_2058,N_187);
or U3928 (N_3928,N_1779,N_1892);
or U3929 (N_3929,N_1283,N_949);
nor U3930 (N_3930,N_1820,N_1755);
nand U3931 (N_3931,N_1149,N_363);
nor U3932 (N_3932,N_2365,N_644);
nand U3933 (N_3933,N_1647,N_1549);
nand U3934 (N_3934,N_1071,N_2017);
nor U3935 (N_3935,N_2256,N_562);
nand U3936 (N_3936,N_2397,N_977);
nand U3937 (N_3937,N_1894,N_2243);
or U3938 (N_3938,N_298,N_1721);
nor U3939 (N_3939,N_2215,N_1615);
nand U3940 (N_3940,N_1565,N_839);
nand U3941 (N_3941,N_2323,N_464);
or U3942 (N_3942,N_1043,N_398);
and U3943 (N_3943,N_646,N_1820);
nor U3944 (N_3944,N_806,N_2384);
nand U3945 (N_3945,N_2193,N_883);
nand U3946 (N_3946,N_1398,N_1992);
nor U3947 (N_3947,N_1298,N_736);
or U3948 (N_3948,N_2369,N_1462);
nand U3949 (N_3949,N_1482,N_2174);
nand U3950 (N_3950,N_289,N_1168);
nand U3951 (N_3951,N_39,N_1242);
and U3952 (N_3952,N_1742,N_2489);
nand U3953 (N_3953,N_1746,N_2435);
or U3954 (N_3954,N_1129,N_310);
nand U3955 (N_3955,N_1827,N_594);
and U3956 (N_3956,N_335,N_1046);
nand U3957 (N_3957,N_1876,N_2308);
or U3958 (N_3958,N_823,N_1495);
nand U3959 (N_3959,N_1166,N_2473);
nor U3960 (N_3960,N_1942,N_812);
and U3961 (N_3961,N_2318,N_145);
nor U3962 (N_3962,N_1925,N_88);
nand U3963 (N_3963,N_1487,N_599);
and U3964 (N_3964,N_1696,N_1451);
and U3965 (N_3965,N_2067,N_1614);
nand U3966 (N_3966,N_204,N_752);
and U3967 (N_3967,N_1291,N_1666);
nand U3968 (N_3968,N_1264,N_2035);
nor U3969 (N_3969,N_647,N_291);
nand U3970 (N_3970,N_585,N_2268);
nand U3971 (N_3971,N_886,N_1630);
nor U3972 (N_3972,N_2178,N_2232);
or U3973 (N_3973,N_2200,N_722);
nand U3974 (N_3974,N_2066,N_1435);
nor U3975 (N_3975,N_2205,N_699);
or U3976 (N_3976,N_289,N_216);
or U3977 (N_3977,N_974,N_750);
or U3978 (N_3978,N_2276,N_1803);
nor U3979 (N_3979,N_676,N_1981);
nor U3980 (N_3980,N_2414,N_153);
or U3981 (N_3981,N_2488,N_1862);
nor U3982 (N_3982,N_403,N_699);
or U3983 (N_3983,N_1904,N_1765);
nand U3984 (N_3984,N_1995,N_503);
and U3985 (N_3985,N_985,N_1908);
or U3986 (N_3986,N_1921,N_1111);
nand U3987 (N_3987,N_767,N_1099);
nor U3988 (N_3988,N_359,N_2483);
and U3989 (N_3989,N_1130,N_441);
nand U3990 (N_3990,N_2290,N_153);
nand U3991 (N_3991,N_1899,N_2261);
xnor U3992 (N_3992,N_933,N_865);
nand U3993 (N_3993,N_132,N_2398);
nor U3994 (N_3994,N_2405,N_1957);
and U3995 (N_3995,N_543,N_1634);
and U3996 (N_3996,N_1749,N_1790);
or U3997 (N_3997,N_983,N_2245);
nand U3998 (N_3998,N_2020,N_1958);
nor U3999 (N_3999,N_1135,N_775);
and U4000 (N_4000,N_2172,N_1658);
or U4001 (N_4001,N_1443,N_1796);
and U4002 (N_4002,N_1772,N_2145);
nand U4003 (N_4003,N_2256,N_870);
or U4004 (N_4004,N_2333,N_730);
nor U4005 (N_4005,N_401,N_678);
or U4006 (N_4006,N_1616,N_289);
nor U4007 (N_4007,N_776,N_2420);
nor U4008 (N_4008,N_1490,N_841);
nand U4009 (N_4009,N_909,N_836);
or U4010 (N_4010,N_69,N_1927);
nand U4011 (N_4011,N_2137,N_1709);
nor U4012 (N_4012,N_1693,N_678);
and U4013 (N_4013,N_1439,N_738);
or U4014 (N_4014,N_1736,N_1512);
nor U4015 (N_4015,N_1035,N_854);
and U4016 (N_4016,N_1919,N_1304);
nand U4017 (N_4017,N_17,N_2416);
nand U4018 (N_4018,N_11,N_187);
nand U4019 (N_4019,N_1613,N_350);
and U4020 (N_4020,N_800,N_1002);
nand U4021 (N_4021,N_1377,N_1700);
or U4022 (N_4022,N_195,N_1021);
nor U4023 (N_4023,N_1974,N_529);
and U4024 (N_4024,N_1954,N_2202);
or U4025 (N_4025,N_914,N_875);
nand U4026 (N_4026,N_1939,N_1552);
nor U4027 (N_4027,N_649,N_1455);
or U4028 (N_4028,N_1884,N_922);
nand U4029 (N_4029,N_1441,N_278);
and U4030 (N_4030,N_2034,N_1269);
nor U4031 (N_4031,N_2439,N_1145);
nor U4032 (N_4032,N_2145,N_1883);
or U4033 (N_4033,N_709,N_2139);
nor U4034 (N_4034,N_551,N_2216);
nor U4035 (N_4035,N_181,N_220);
nand U4036 (N_4036,N_528,N_1826);
or U4037 (N_4037,N_1866,N_1700);
or U4038 (N_4038,N_2166,N_219);
or U4039 (N_4039,N_2112,N_783);
or U4040 (N_4040,N_1316,N_206);
nand U4041 (N_4041,N_1762,N_736);
nand U4042 (N_4042,N_1705,N_2148);
or U4043 (N_4043,N_587,N_1122);
and U4044 (N_4044,N_1161,N_1297);
nand U4045 (N_4045,N_2499,N_552);
nand U4046 (N_4046,N_2412,N_954);
or U4047 (N_4047,N_1430,N_1850);
and U4048 (N_4048,N_95,N_190);
or U4049 (N_4049,N_1410,N_845);
nand U4050 (N_4050,N_2159,N_1850);
and U4051 (N_4051,N_232,N_832);
and U4052 (N_4052,N_817,N_2356);
and U4053 (N_4053,N_1542,N_1219);
nand U4054 (N_4054,N_2241,N_2467);
and U4055 (N_4055,N_1120,N_951);
or U4056 (N_4056,N_395,N_828);
and U4057 (N_4057,N_2440,N_13);
nor U4058 (N_4058,N_1266,N_139);
nor U4059 (N_4059,N_81,N_2395);
or U4060 (N_4060,N_260,N_1073);
and U4061 (N_4061,N_367,N_1990);
nor U4062 (N_4062,N_126,N_2409);
nor U4063 (N_4063,N_2238,N_1903);
or U4064 (N_4064,N_1774,N_695);
and U4065 (N_4065,N_1449,N_1350);
nand U4066 (N_4066,N_2477,N_1056);
and U4067 (N_4067,N_2085,N_222);
or U4068 (N_4068,N_487,N_2290);
nor U4069 (N_4069,N_472,N_2478);
and U4070 (N_4070,N_2381,N_1710);
nor U4071 (N_4071,N_1358,N_370);
or U4072 (N_4072,N_745,N_234);
and U4073 (N_4073,N_1858,N_1281);
and U4074 (N_4074,N_837,N_209);
and U4075 (N_4075,N_699,N_2369);
or U4076 (N_4076,N_1097,N_1512);
nor U4077 (N_4077,N_384,N_1297);
and U4078 (N_4078,N_1195,N_1031);
nand U4079 (N_4079,N_249,N_911);
or U4080 (N_4080,N_166,N_1926);
and U4081 (N_4081,N_1839,N_484);
or U4082 (N_4082,N_1405,N_1402);
nor U4083 (N_4083,N_867,N_1251);
nor U4084 (N_4084,N_169,N_1653);
nand U4085 (N_4085,N_446,N_1801);
nor U4086 (N_4086,N_605,N_697);
and U4087 (N_4087,N_1518,N_2057);
nor U4088 (N_4088,N_834,N_1296);
nor U4089 (N_4089,N_1870,N_1622);
and U4090 (N_4090,N_2257,N_1429);
nor U4091 (N_4091,N_870,N_1184);
or U4092 (N_4092,N_395,N_1265);
or U4093 (N_4093,N_1204,N_2400);
nand U4094 (N_4094,N_1783,N_934);
and U4095 (N_4095,N_284,N_890);
or U4096 (N_4096,N_1068,N_1678);
nor U4097 (N_4097,N_2080,N_194);
nand U4098 (N_4098,N_1931,N_655);
nand U4099 (N_4099,N_1192,N_1460);
nand U4100 (N_4100,N_11,N_673);
nor U4101 (N_4101,N_53,N_281);
nor U4102 (N_4102,N_2031,N_817);
nand U4103 (N_4103,N_520,N_437);
or U4104 (N_4104,N_1568,N_2476);
or U4105 (N_4105,N_1128,N_1604);
nor U4106 (N_4106,N_1689,N_1170);
nand U4107 (N_4107,N_751,N_1964);
or U4108 (N_4108,N_2354,N_1334);
or U4109 (N_4109,N_1898,N_2288);
nor U4110 (N_4110,N_372,N_1594);
and U4111 (N_4111,N_1483,N_2073);
and U4112 (N_4112,N_225,N_733);
and U4113 (N_4113,N_2162,N_325);
and U4114 (N_4114,N_768,N_2124);
or U4115 (N_4115,N_1952,N_1997);
and U4116 (N_4116,N_428,N_692);
or U4117 (N_4117,N_1000,N_1431);
nor U4118 (N_4118,N_1339,N_1922);
and U4119 (N_4119,N_2139,N_2253);
nand U4120 (N_4120,N_55,N_1859);
nor U4121 (N_4121,N_994,N_2348);
nand U4122 (N_4122,N_210,N_748);
nor U4123 (N_4123,N_1489,N_197);
nand U4124 (N_4124,N_725,N_580);
nor U4125 (N_4125,N_368,N_1098);
nand U4126 (N_4126,N_1300,N_38);
nand U4127 (N_4127,N_1177,N_1144);
nor U4128 (N_4128,N_1598,N_2367);
and U4129 (N_4129,N_656,N_593);
nand U4130 (N_4130,N_1197,N_608);
and U4131 (N_4131,N_933,N_1882);
and U4132 (N_4132,N_1486,N_2275);
nor U4133 (N_4133,N_1273,N_870);
or U4134 (N_4134,N_206,N_596);
nor U4135 (N_4135,N_1123,N_2143);
and U4136 (N_4136,N_1998,N_129);
and U4137 (N_4137,N_769,N_1441);
or U4138 (N_4138,N_1156,N_1314);
xor U4139 (N_4139,N_210,N_747);
nor U4140 (N_4140,N_1568,N_1222);
or U4141 (N_4141,N_225,N_1324);
nor U4142 (N_4142,N_1068,N_229);
nor U4143 (N_4143,N_1628,N_192);
nand U4144 (N_4144,N_1700,N_620);
and U4145 (N_4145,N_1329,N_528);
nor U4146 (N_4146,N_901,N_1168);
and U4147 (N_4147,N_579,N_1054);
or U4148 (N_4148,N_367,N_1190);
nor U4149 (N_4149,N_1272,N_125);
and U4150 (N_4150,N_871,N_286);
nand U4151 (N_4151,N_1246,N_67);
and U4152 (N_4152,N_2209,N_2340);
or U4153 (N_4153,N_220,N_1448);
nor U4154 (N_4154,N_1433,N_1891);
or U4155 (N_4155,N_406,N_1022);
and U4156 (N_4156,N_280,N_1107);
or U4157 (N_4157,N_1438,N_1095);
or U4158 (N_4158,N_105,N_864);
or U4159 (N_4159,N_11,N_2178);
and U4160 (N_4160,N_1228,N_1642);
nor U4161 (N_4161,N_2314,N_1053);
nor U4162 (N_4162,N_1791,N_1534);
and U4163 (N_4163,N_279,N_2271);
nand U4164 (N_4164,N_2258,N_1536);
or U4165 (N_4165,N_299,N_811);
nand U4166 (N_4166,N_1140,N_1285);
and U4167 (N_4167,N_930,N_428);
nand U4168 (N_4168,N_1648,N_1787);
nor U4169 (N_4169,N_1718,N_2318);
nor U4170 (N_4170,N_858,N_2404);
or U4171 (N_4171,N_923,N_303);
or U4172 (N_4172,N_1197,N_2336);
nand U4173 (N_4173,N_109,N_599);
and U4174 (N_4174,N_638,N_2274);
or U4175 (N_4175,N_515,N_1788);
nand U4176 (N_4176,N_1622,N_574);
nand U4177 (N_4177,N_1023,N_2459);
or U4178 (N_4178,N_2272,N_42);
nand U4179 (N_4179,N_1156,N_1407);
and U4180 (N_4180,N_253,N_351);
nor U4181 (N_4181,N_1158,N_1499);
nand U4182 (N_4182,N_1758,N_38);
nor U4183 (N_4183,N_2412,N_1645);
or U4184 (N_4184,N_2271,N_2056);
and U4185 (N_4185,N_1629,N_1136);
and U4186 (N_4186,N_1589,N_1360);
nor U4187 (N_4187,N_464,N_1747);
nor U4188 (N_4188,N_1189,N_2337);
and U4189 (N_4189,N_912,N_1427);
nand U4190 (N_4190,N_702,N_2407);
nor U4191 (N_4191,N_688,N_88);
nand U4192 (N_4192,N_371,N_729);
or U4193 (N_4193,N_646,N_124);
or U4194 (N_4194,N_970,N_826);
nand U4195 (N_4195,N_2350,N_1679);
or U4196 (N_4196,N_281,N_1352);
nand U4197 (N_4197,N_514,N_1424);
nand U4198 (N_4198,N_600,N_1583);
and U4199 (N_4199,N_1513,N_744);
nor U4200 (N_4200,N_658,N_1054);
nand U4201 (N_4201,N_89,N_2052);
and U4202 (N_4202,N_1364,N_487);
nand U4203 (N_4203,N_2218,N_776);
or U4204 (N_4204,N_517,N_1884);
nand U4205 (N_4205,N_1016,N_1279);
and U4206 (N_4206,N_1207,N_2408);
or U4207 (N_4207,N_269,N_959);
and U4208 (N_4208,N_1336,N_1246);
nand U4209 (N_4209,N_1223,N_441);
xnor U4210 (N_4210,N_2266,N_1179);
nor U4211 (N_4211,N_800,N_90);
and U4212 (N_4212,N_1648,N_2454);
nor U4213 (N_4213,N_469,N_1714);
and U4214 (N_4214,N_721,N_2073);
nand U4215 (N_4215,N_2019,N_1060);
nand U4216 (N_4216,N_890,N_1229);
nor U4217 (N_4217,N_1056,N_2209);
or U4218 (N_4218,N_1759,N_1609);
nand U4219 (N_4219,N_182,N_1842);
or U4220 (N_4220,N_2373,N_509);
and U4221 (N_4221,N_2234,N_1321);
nor U4222 (N_4222,N_670,N_1322);
nor U4223 (N_4223,N_112,N_612);
or U4224 (N_4224,N_558,N_1515);
or U4225 (N_4225,N_196,N_268);
nor U4226 (N_4226,N_394,N_612);
or U4227 (N_4227,N_1712,N_1046);
or U4228 (N_4228,N_1770,N_1368);
or U4229 (N_4229,N_1607,N_2060);
or U4230 (N_4230,N_114,N_365);
and U4231 (N_4231,N_73,N_2198);
nand U4232 (N_4232,N_876,N_167);
and U4233 (N_4233,N_341,N_496);
nor U4234 (N_4234,N_1641,N_1079);
and U4235 (N_4235,N_560,N_344);
nand U4236 (N_4236,N_2238,N_79);
nand U4237 (N_4237,N_1202,N_1090);
nor U4238 (N_4238,N_1410,N_2091);
nor U4239 (N_4239,N_1063,N_301);
or U4240 (N_4240,N_184,N_1269);
nand U4241 (N_4241,N_881,N_290);
nor U4242 (N_4242,N_618,N_1350);
or U4243 (N_4243,N_1054,N_2120);
nor U4244 (N_4244,N_1712,N_604);
or U4245 (N_4245,N_173,N_277);
and U4246 (N_4246,N_2339,N_131);
nand U4247 (N_4247,N_119,N_389);
nor U4248 (N_4248,N_567,N_1224);
nand U4249 (N_4249,N_1662,N_1189);
nand U4250 (N_4250,N_438,N_717);
or U4251 (N_4251,N_226,N_1860);
and U4252 (N_4252,N_21,N_310);
nand U4253 (N_4253,N_2005,N_309);
nand U4254 (N_4254,N_663,N_853);
nand U4255 (N_4255,N_1950,N_377);
and U4256 (N_4256,N_1260,N_2209);
nor U4257 (N_4257,N_2497,N_1841);
and U4258 (N_4258,N_2450,N_196);
or U4259 (N_4259,N_1830,N_1475);
and U4260 (N_4260,N_992,N_1934);
and U4261 (N_4261,N_2085,N_2453);
nor U4262 (N_4262,N_500,N_309);
and U4263 (N_4263,N_154,N_1049);
and U4264 (N_4264,N_2244,N_233);
and U4265 (N_4265,N_766,N_776);
or U4266 (N_4266,N_1381,N_1931);
or U4267 (N_4267,N_1033,N_1918);
nor U4268 (N_4268,N_2393,N_2181);
or U4269 (N_4269,N_373,N_449);
nor U4270 (N_4270,N_2400,N_817);
and U4271 (N_4271,N_1743,N_1995);
nand U4272 (N_4272,N_136,N_1456);
and U4273 (N_4273,N_1226,N_2310);
or U4274 (N_4274,N_648,N_1340);
nor U4275 (N_4275,N_970,N_1721);
or U4276 (N_4276,N_350,N_1589);
and U4277 (N_4277,N_894,N_1381);
nand U4278 (N_4278,N_1566,N_781);
nor U4279 (N_4279,N_1709,N_2265);
nand U4280 (N_4280,N_2478,N_1538);
nand U4281 (N_4281,N_1027,N_1357);
nand U4282 (N_4282,N_1861,N_1897);
nor U4283 (N_4283,N_2031,N_298);
nor U4284 (N_4284,N_2263,N_301);
or U4285 (N_4285,N_1228,N_2333);
nand U4286 (N_4286,N_1652,N_2131);
or U4287 (N_4287,N_110,N_1192);
nand U4288 (N_4288,N_511,N_1202);
or U4289 (N_4289,N_2088,N_2153);
or U4290 (N_4290,N_1544,N_626);
or U4291 (N_4291,N_458,N_1605);
nand U4292 (N_4292,N_73,N_1866);
or U4293 (N_4293,N_1072,N_464);
or U4294 (N_4294,N_372,N_2393);
nand U4295 (N_4295,N_718,N_2018);
nor U4296 (N_4296,N_1679,N_1886);
and U4297 (N_4297,N_37,N_1841);
or U4298 (N_4298,N_412,N_486);
nand U4299 (N_4299,N_721,N_1311);
nand U4300 (N_4300,N_153,N_157);
nand U4301 (N_4301,N_2134,N_1505);
and U4302 (N_4302,N_588,N_1443);
nand U4303 (N_4303,N_1846,N_1239);
nor U4304 (N_4304,N_1598,N_565);
and U4305 (N_4305,N_1087,N_764);
nor U4306 (N_4306,N_1291,N_1688);
nor U4307 (N_4307,N_882,N_936);
and U4308 (N_4308,N_666,N_1994);
nor U4309 (N_4309,N_1396,N_1131);
and U4310 (N_4310,N_1514,N_2377);
nand U4311 (N_4311,N_1367,N_294);
or U4312 (N_4312,N_76,N_2432);
nor U4313 (N_4313,N_324,N_160);
and U4314 (N_4314,N_1189,N_463);
or U4315 (N_4315,N_604,N_1432);
nor U4316 (N_4316,N_1449,N_1347);
and U4317 (N_4317,N_76,N_136);
xnor U4318 (N_4318,N_738,N_2334);
nor U4319 (N_4319,N_1982,N_895);
and U4320 (N_4320,N_2058,N_1780);
and U4321 (N_4321,N_949,N_2258);
and U4322 (N_4322,N_790,N_1613);
nand U4323 (N_4323,N_314,N_1065);
nor U4324 (N_4324,N_2060,N_1339);
or U4325 (N_4325,N_445,N_258);
nor U4326 (N_4326,N_1559,N_1450);
and U4327 (N_4327,N_745,N_1361);
or U4328 (N_4328,N_1971,N_1757);
and U4329 (N_4329,N_1866,N_882);
and U4330 (N_4330,N_2222,N_639);
nand U4331 (N_4331,N_1801,N_149);
or U4332 (N_4332,N_2273,N_181);
and U4333 (N_4333,N_18,N_1082);
or U4334 (N_4334,N_1,N_613);
nor U4335 (N_4335,N_564,N_2156);
and U4336 (N_4336,N_1511,N_224);
nand U4337 (N_4337,N_397,N_808);
or U4338 (N_4338,N_228,N_1325);
and U4339 (N_4339,N_2227,N_39);
nor U4340 (N_4340,N_2166,N_1611);
or U4341 (N_4341,N_1251,N_1288);
or U4342 (N_4342,N_2419,N_582);
and U4343 (N_4343,N_338,N_2171);
or U4344 (N_4344,N_2413,N_229);
nor U4345 (N_4345,N_1078,N_1361);
nand U4346 (N_4346,N_2025,N_2065);
and U4347 (N_4347,N_1350,N_1877);
and U4348 (N_4348,N_913,N_1708);
and U4349 (N_4349,N_1400,N_591);
xnor U4350 (N_4350,N_878,N_1268);
nor U4351 (N_4351,N_1666,N_799);
and U4352 (N_4352,N_1134,N_1121);
or U4353 (N_4353,N_514,N_1641);
nor U4354 (N_4354,N_1545,N_1080);
nand U4355 (N_4355,N_372,N_2480);
and U4356 (N_4356,N_988,N_1082);
nand U4357 (N_4357,N_2203,N_58);
nand U4358 (N_4358,N_287,N_498);
or U4359 (N_4359,N_2080,N_1578);
nor U4360 (N_4360,N_1011,N_249);
nand U4361 (N_4361,N_1625,N_378);
nand U4362 (N_4362,N_571,N_326);
nor U4363 (N_4363,N_1887,N_2141);
nor U4364 (N_4364,N_2353,N_1265);
nand U4365 (N_4365,N_1840,N_583);
nor U4366 (N_4366,N_139,N_1409);
nor U4367 (N_4367,N_36,N_221);
and U4368 (N_4368,N_661,N_903);
nand U4369 (N_4369,N_2486,N_1085);
nand U4370 (N_4370,N_964,N_1255);
or U4371 (N_4371,N_1943,N_2137);
or U4372 (N_4372,N_1431,N_126);
nand U4373 (N_4373,N_1221,N_2019);
or U4374 (N_4374,N_1827,N_1120);
or U4375 (N_4375,N_1586,N_957);
or U4376 (N_4376,N_178,N_871);
and U4377 (N_4377,N_692,N_68);
nor U4378 (N_4378,N_1742,N_1409);
nand U4379 (N_4379,N_322,N_1182);
and U4380 (N_4380,N_1256,N_271);
or U4381 (N_4381,N_1521,N_202);
or U4382 (N_4382,N_110,N_1137);
nand U4383 (N_4383,N_144,N_1563);
or U4384 (N_4384,N_1727,N_366);
and U4385 (N_4385,N_1625,N_1289);
nor U4386 (N_4386,N_259,N_443);
or U4387 (N_4387,N_432,N_846);
or U4388 (N_4388,N_646,N_1818);
and U4389 (N_4389,N_1364,N_2363);
and U4390 (N_4390,N_1964,N_487);
and U4391 (N_4391,N_2172,N_1665);
nand U4392 (N_4392,N_839,N_1998);
and U4393 (N_4393,N_1154,N_1333);
nand U4394 (N_4394,N_343,N_1976);
nor U4395 (N_4395,N_17,N_371);
or U4396 (N_4396,N_1594,N_708);
or U4397 (N_4397,N_890,N_858);
and U4398 (N_4398,N_306,N_671);
and U4399 (N_4399,N_2165,N_822);
nor U4400 (N_4400,N_1416,N_1441);
and U4401 (N_4401,N_1691,N_1217);
or U4402 (N_4402,N_382,N_410);
or U4403 (N_4403,N_771,N_967);
or U4404 (N_4404,N_1769,N_34);
or U4405 (N_4405,N_1268,N_2137);
nor U4406 (N_4406,N_945,N_1269);
and U4407 (N_4407,N_331,N_1315);
nand U4408 (N_4408,N_72,N_2173);
and U4409 (N_4409,N_1379,N_2378);
or U4410 (N_4410,N_88,N_193);
or U4411 (N_4411,N_2153,N_305);
or U4412 (N_4412,N_1155,N_585);
or U4413 (N_4413,N_2318,N_221);
nand U4414 (N_4414,N_797,N_121);
or U4415 (N_4415,N_1152,N_633);
and U4416 (N_4416,N_269,N_392);
nor U4417 (N_4417,N_2270,N_1988);
and U4418 (N_4418,N_2093,N_167);
and U4419 (N_4419,N_1928,N_249);
or U4420 (N_4420,N_2405,N_2475);
nand U4421 (N_4421,N_2292,N_1009);
nand U4422 (N_4422,N_1700,N_1093);
and U4423 (N_4423,N_594,N_2041);
or U4424 (N_4424,N_382,N_748);
nand U4425 (N_4425,N_695,N_66);
or U4426 (N_4426,N_1325,N_699);
and U4427 (N_4427,N_1978,N_130);
and U4428 (N_4428,N_156,N_1051);
nor U4429 (N_4429,N_2153,N_1935);
or U4430 (N_4430,N_1002,N_1188);
nand U4431 (N_4431,N_444,N_454);
xor U4432 (N_4432,N_1510,N_1900);
or U4433 (N_4433,N_72,N_2158);
nor U4434 (N_4434,N_1937,N_1110);
nand U4435 (N_4435,N_909,N_2141);
nand U4436 (N_4436,N_2023,N_191);
nor U4437 (N_4437,N_2224,N_1327);
or U4438 (N_4438,N_1358,N_1168);
or U4439 (N_4439,N_1105,N_2426);
or U4440 (N_4440,N_2188,N_1136);
and U4441 (N_4441,N_1806,N_2493);
nor U4442 (N_4442,N_2087,N_2172);
or U4443 (N_4443,N_1013,N_1798);
nand U4444 (N_4444,N_1455,N_1189);
nand U4445 (N_4445,N_1947,N_628);
nor U4446 (N_4446,N_952,N_2227);
nor U4447 (N_4447,N_764,N_1065);
and U4448 (N_4448,N_2460,N_613);
or U4449 (N_4449,N_1199,N_2402);
or U4450 (N_4450,N_892,N_1714);
or U4451 (N_4451,N_1248,N_1409);
or U4452 (N_4452,N_1839,N_1561);
and U4453 (N_4453,N_545,N_457);
nand U4454 (N_4454,N_621,N_397);
nor U4455 (N_4455,N_1310,N_2058);
and U4456 (N_4456,N_432,N_830);
or U4457 (N_4457,N_1282,N_2481);
and U4458 (N_4458,N_2423,N_1416);
nand U4459 (N_4459,N_1067,N_2259);
nor U4460 (N_4460,N_1384,N_642);
xor U4461 (N_4461,N_1761,N_109);
nand U4462 (N_4462,N_2225,N_856);
and U4463 (N_4463,N_55,N_2392);
and U4464 (N_4464,N_116,N_2415);
nor U4465 (N_4465,N_577,N_1965);
nand U4466 (N_4466,N_166,N_1290);
nor U4467 (N_4467,N_1492,N_2032);
and U4468 (N_4468,N_379,N_2154);
and U4469 (N_4469,N_489,N_958);
nor U4470 (N_4470,N_1933,N_2365);
or U4471 (N_4471,N_2071,N_1132);
and U4472 (N_4472,N_1585,N_1909);
nand U4473 (N_4473,N_403,N_784);
and U4474 (N_4474,N_2134,N_1897);
nand U4475 (N_4475,N_12,N_1309);
xor U4476 (N_4476,N_1583,N_1821);
nand U4477 (N_4477,N_1502,N_1537);
and U4478 (N_4478,N_294,N_940);
nand U4479 (N_4479,N_1980,N_1855);
and U4480 (N_4480,N_2099,N_301);
and U4481 (N_4481,N_1430,N_347);
or U4482 (N_4482,N_1716,N_703);
nand U4483 (N_4483,N_1454,N_2462);
nand U4484 (N_4484,N_804,N_1903);
and U4485 (N_4485,N_1077,N_1108);
nand U4486 (N_4486,N_1500,N_1237);
nor U4487 (N_4487,N_662,N_1172);
nor U4488 (N_4488,N_1612,N_2382);
nor U4489 (N_4489,N_2304,N_2109);
nand U4490 (N_4490,N_1863,N_266);
or U4491 (N_4491,N_1633,N_744);
or U4492 (N_4492,N_933,N_1234);
or U4493 (N_4493,N_2150,N_2295);
nand U4494 (N_4494,N_2430,N_1291);
nor U4495 (N_4495,N_606,N_1849);
and U4496 (N_4496,N_2194,N_1416);
and U4497 (N_4497,N_1437,N_2291);
nor U4498 (N_4498,N_537,N_405);
or U4499 (N_4499,N_987,N_1037);
xnor U4500 (N_4500,N_211,N_878);
or U4501 (N_4501,N_362,N_2477);
nor U4502 (N_4502,N_94,N_1754);
nor U4503 (N_4503,N_2077,N_1230);
nand U4504 (N_4504,N_1273,N_1548);
and U4505 (N_4505,N_783,N_550);
nor U4506 (N_4506,N_347,N_275);
or U4507 (N_4507,N_1463,N_992);
nor U4508 (N_4508,N_523,N_1302);
nor U4509 (N_4509,N_1652,N_1641);
nand U4510 (N_4510,N_353,N_2188);
or U4511 (N_4511,N_275,N_891);
nor U4512 (N_4512,N_1321,N_1357);
nand U4513 (N_4513,N_2361,N_2312);
nor U4514 (N_4514,N_578,N_1144);
nor U4515 (N_4515,N_1019,N_1920);
or U4516 (N_4516,N_682,N_805);
or U4517 (N_4517,N_1875,N_1846);
nand U4518 (N_4518,N_1718,N_876);
nor U4519 (N_4519,N_688,N_1948);
or U4520 (N_4520,N_1313,N_2240);
and U4521 (N_4521,N_2113,N_211);
nand U4522 (N_4522,N_88,N_463);
or U4523 (N_4523,N_2471,N_1561);
or U4524 (N_4524,N_1041,N_2248);
nand U4525 (N_4525,N_1052,N_2129);
and U4526 (N_4526,N_2196,N_1522);
nor U4527 (N_4527,N_281,N_654);
and U4528 (N_4528,N_1565,N_927);
nor U4529 (N_4529,N_2289,N_2300);
nand U4530 (N_4530,N_2317,N_1390);
nor U4531 (N_4531,N_879,N_157);
nor U4532 (N_4532,N_1683,N_2332);
and U4533 (N_4533,N_1602,N_2307);
nand U4534 (N_4534,N_1546,N_2137);
nor U4535 (N_4535,N_752,N_1724);
nor U4536 (N_4536,N_257,N_951);
or U4537 (N_4537,N_2173,N_1785);
nor U4538 (N_4538,N_1882,N_1307);
nand U4539 (N_4539,N_1204,N_955);
or U4540 (N_4540,N_2497,N_2168);
nor U4541 (N_4541,N_1790,N_1850);
nor U4542 (N_4542,N_2048,N_383);
and U4543 (N_4543,N_2465,N_2033);
and U4544 (N_4544,N_1766,N_441);
nand U4545 (N_4545,N_1476,N_121);
or U4546 (N_4546,N_271,N_1131);
or U4547 (N_4547,N_174,N_801);
nand U4548 (N_4548,N_696,N_1877);
nand U4549 (N_4549,N_312,N_1185);
or U4550 (N_4550,N_2383,N_1887);
and U4551 (N_4551,N_1752,N_704);
nor U4552 (N_4552,N_259,N_2256);
nand U4553 (N_4553,N_1980,N_318);
and U4554 (N_4554,N_2316,N_1817);
and U4555 (N_4555,N_1565,N_49);
nand U4556 (N_4556,N_1236,N_2476);
nand U4557 (N_4557,N_1676,N_669);
nand U4558 (N_4558,N_2083,N_1532);
or U4559 (N_4559,N_1160,N_850);
or U4560 (N_4560,N_1962,N_1981);
and U4561 (N_4561,N_486,N_971);
or U4562 (N_4562,N_2347,N_2409);
nor U4563 (N_4563,N_1822,N_160);
nor U4564 (N_4564,N_2486,N_2068);
or U4565 (N_4565,N_680,N_2075);
nand U4566 (N_4566,N_1382,N_753);
or U4567 (N_4567,N_2347,N_1496);
and U4568 (N_4568,N_1680,N_447);
nand U4569 (N_4569,N_2437,N_1473);
and U4570 (N_4570,N_1271,N_813);
nand U4571 (N_4571,N_512,N_784);
or U4572 (N_4572,N_1482,N_587);
or U4573 (N_4573,N_775,N_1488);
nand U4574 (N_4574,N_2477,N_1886);
or U4575 (N_4575,N_1706,N_892);
nor U4576 (N_4576,N_2368,N_2082);
nor U4577 (N_4577,N_1383,N_1149);
nor U4578 (N_4578,N_630,N_1123);
or U4579 (N_4579,N_611,N_189);
and U4580 (N_4580,N_9,N_1747);
and U4581 (N_4581,N_2221,N_934);
xor U4582 (N_4582,N_1226,N_1961);
and U4583 (N_4583,N_2437,N_372);
nand U4584 (N_4584,N_1712,N_1298);
nor U4585 (N_4585,N_2454,N_446);
nand U4586 (N_4586,N_2111,N_459);
and U4587 (N_4587,N_2484,N_104);
nor U4588 (N_4588,N_1331,N_1555);
and U4589 (N_4589,N_187,N_175);
nor U4590 (N_4590,N_1079,N_886);
nor U4591 (N_4591,N_1159,N_1822);
and U4592 (N_4592,N_40,N_539);
nand U4593 (N_4593,N_2087,N_571);
nand U4594 (N_4594,N_484,N_1739);
nand U4595 (N_4595,N_620,N_1359);
and U4596 (N_4596,N_2252,N_1507);
or U4597 (N_4597,N_274,N_2005);
nand U4598 (N_4598,N_494,N_2100);
nand U4599 (N_4599,N_1782,N_1765);
nand U4600 (N_4600,N_1124,N_2209);
and U4601 (N_4601,N_1145,N_998);
or U4602 (N_4602,N_2481,N_1397);
and U4603 (N_4603,N_2088,N_1104);
nor U4604 (N_4604,N_747,N_2458);
nand U4605 (N_4605,N_38,N_2026);
nand U4606 (N_4606,N_955,N_2172);
nor U4607 (N_4607,N_2206,N_960);
or U4608 (N_4608,N_666,N_1735);
and U4609 (N_4609,N_194,N_382);
nor U4610 (N_4610,N_2060,N_1408);
nor U4611 (N_4611,N_85,N_1260);
or U4612 (N_4612,N_434,N_802);
nor U4613 (N_4613,N_1996,N_2004);
nand U4614 (N_4614,N_1670,N_625);
and U4615 (N_4615,N_1525,N_1340);
nor U4616 (N_4616,N_1960,N_840);
and U4617 (N_4617,N_1481,N_1805);
and U4618 (N_4618,N_920,N_646);
or U4619 (N_4619,N_2104,N_1784);
and U4620 (N_4620,N_1399,N_629);
or U4621 (N_4621,N_1608,N_422);
and U4622 (N_4622,N_2218,N_282);
nand U4623 (N_4623,N_1647,N_1288);
nor U4624 (N_4624,N_660,N_1355);
and U4625 (N_4625,N_1172,N_1841);
and U4626 (N_4626,N_1467,N_379);
or U4627 (N_4627,N_2286,N_1034);
nand U4628 (N_4628,N_2432,N_1285);
and U4629 (N_4629,N_10,N_24);
or U4630 (N_4630,N_1104,N_1391);
xor U4631 (N_4631,N_345,N_1262);
nor U4632 (N_4632,N_426,N_1097);
nor U4633 (N_4633,N_525,N_1334);
nor U4634 (N_4634,N_669,N_1414);
and U4635 (N_4635,N_101,N_734);
xnor U4636 (N_4636,N_994,N_858);
nand U4637 (N_4637,N_2183,N_1236);
and U4638 (N_4638,N_2078,N_325);
nor U4639 (N_4639,N_1900,N_973);
or U4640 (N_4640,N_75,N_791);
nand U4641 (N_4641,N_2460,N_1640);
and U4642 (N_4642,N_1071,N_1846);
or U4643 (N_4643,N_1620,N_1161);
or U4644 (N_4644,N_2049,N_2010);
nor U4645 (N_4645,N_1132,N_2462);
nor U4646 (N_4646,N_2293,N_1278);
or U4647 (N_4647,N_686,N_1905);
and U4648 (N_4648,N_1580,N_1375);
and U4649 (N_4649,N_1467,N_1113);
nand U4650 (N_4650,N_173,N_2084);
nand U4651 (N_4651,N_649,N_317);
nand U4652 (N_4652,N_308,N_803);
nand U4653 (N_4653,N_731,N_1634);
nor U4654 (N_4654,N_512,N_2018);
nor U4655 (N_4655,N_955,N_2250);
nand U4656 (N_4656,N_2489,N_323);
xnor U4657 (N_4657,N_2275,N_2149);
nand U4658 (N_4658,N_235,N_2269);
nand U4659 (N_4659,N_1036,N_303);
and U4660 (N_4660,N_1938,N_1838);
nor U4661 (N_4661,N_556,N_1751);
nand U4662 (N_4662,N_1163,N_163);
nor U4663 (N_4663,N_1202,N_2432);
nand U4664 (N_4664,N_1368,N_179);
nand U4665 (N_4665,N_1841,N_1890);
and U4666 (N_4666,N_2171,N_1281);
nand U4667 (N_4667,N_1902,N_788);
nor U4668 (N_4668,N_891,N_393);
or U4669 (N_4669,N_1173,N_724);
nand U4670 (N_4670,N_2163,N_2201);
nor U4671 (N_4671,N_1292,N_2369);
and U4672 (N_4672,N_251,N_1833);
nor U4673 (N_4673,N_180,N_565);
or U4674 (N_4674,N_1722,N_1000);
nor U4675 (N_4675,N_665,N_1197);
nand U4676 (N_4676,N_319,N_250);
nor U4677 (N_4677,N_2444,N_524);
nor U4678 (N_4678,N_1680,N_1045);
xor U4679 (N_4679,N_124,N_1860);
nor U4680 (N_4680,N_548,N_1779);
nor U4681 (N_4681,N_2383,N_1109);
and U4682 (N_4682,N_1152,N_248);
nor U4683 (N_4683,N_268,N_719);
nor U4684 (N_4684,N_1898,N_450);
nand U4685 (N_4685,N_1276,N_2121);
or U4686 (N_4686,N_381,N_306);
nor U4687 (N_4687,N_1279,N_735);
and U4688 (N_4688,N_283,N_646);
or U4689 (N_4689,N_2341,N_1471);
and U4690 (N_4690,N_1265,N_2046);
nand U4691 (N_4691,N_559,N_894);
and U4692 (N_4692,N_2322,N_2193);
and U4693 (N_4693,N_2358,N_1842);
or U4694 (N_4694,N_124,N_1049);
nor U4695 (N_4695,N_0,N_619);
nand U4696 (N_4696,N_907,N_1256);
or U4697 (N_4697,N_1129,N_1803);
nor U4698 (N_4698,N_1805,N_896);
and U4699 (N_4699,N_2414,N_2476);
nor U4700 (N_4700,N_1830,N_82);
or U4701 (N_4701,N_771,N_709);
and U4702 (N_4702,N_1018,N_1881);
or U4703 (N_4703,N_1272,N_2404);
or U4704 (N_4704,N_1682,N_1764);
and U4705 (N_4705,N_509,N_199);
and U4706 (N_4706,N_50,N_234);
and U4707 (N_4707,N_251,N_37);
nand U4708 (N_4708,N_2234,N_1996);
and U4709 (N_4709,N_822,N_1315);
nor U4710 (N_4710,N_1011,N_1485);
or U4711 (N_4711,N_2091,N_1133);
nor U4712 (N_4712,N_2249,N_1057);
or U4713 (N_4713,N_1828,N_746);
nor U4714 (N_4714,N_2386,N_722);
or U4715 (N_4715,N_1395,N_1277);
nor U4716 (N_4716,N_494,N_1680);
or U4717 (N_4717,N_629,N_31);
nand U4718 (N_4718,N_402,N_1262);
nor U4719 (N_4719,N_1725,N_1926);
and U4720 (N_4720,N_2446,N_2261);
nand U4721 (N_4721,N_2342,N_2334);
or U4722 (N_4722,N_1052,N_328);
and U4723 (N_4723,N_151,N_1856);
nand U4724 (N_4724,N_177,N_1113);
nor U4725 (N_4725,N_97,N_549);
or U4726 (N_4726,N_1666,N_33);
nor U4727 (N_4727,N_244,N_448);
or U4728 (N_4728,N_741,N_1932);
nor U4729 (N_4729,N_641,N_1512);
and U4730 (N_4730,N_643,N_216);
or U4731 (N_4731,N_1167,N_2198);
or U4732 (N_4732,N_1423,N_1846);
or U4733 (N_4733,N_526,N_768);
or U4734 (N_4734,N_1882,N_235);
and U4735 (N_4735,N_1346,N_323);
or U4736 (N_4736,N_525,N_1241);
nand U4737 (N_4737,N_2165,N_83);
and U4738 (N_4738,N_1638,N_1644);
or U4739 (N_4739,N_873,N_136);
or U4740 (N_4740,N_822,N_2280);
nor U4741 (N_4741,N_261,N_520);
nand U4742 (N_4742,N_1055,N_365);
nand U4743 (N_4743,N_1075,N_2049);
or U4744 (N_4744,N_81,N_592);
and U4745 (N_4745,N_897,N_2241);
or U4746 (N_4746,N_1031,N_468);
nand U4747 (N_4747,N_138,N_428);
nor U4748 (N_4748,N_2329,N_1669);
nor U4749 (N_4749,N_150,N_2193);
nand U4750 (N_4750,N_721,N_1559);
and U4751 (N_4751,N_414,N_351);
or U4752 (N_4752,N_946,N_2427);
and U4753 (N_4753,N_1396,N_2481);
nand U4754 (N_4754,N_1352,N_2047);
nor U4755 (N_4755,N_497,N_1096);
and U4756 (N_4756,N_1318,N_1170);
nor U4757 (N_4757,N_1022,N_637);
nor U4758 (N_4758,N_2264,N_1385);
nand U4759 (N_4759,N_406,N_1845);
nand U4760 (N_4760,N_1325,N_1947);
or U4761 (N_4761,N_981,N_1669);
nor U4762 (N_4762,N_1278,N_1869);
nand U4763 (N_4763,N_597,N_811);
and U4764 (N_4764,N_2093,N_1466);
nor U4765 (N_4765,N_502,N_1606);
nand U4766 (N_4766,N_588,N_2008);
nand U4767 (N_4767,N_1166,N_566);
and U4768 (N_4768,N_31,N_1024);
and U4769 (N_4769,N_1777,N_297);
and U4770 (N_4770,N_335,N_543);
nand U4771 (N_4771,N_315,N_1007);
or U4772 (N_4772,N_639,N_1948);
nand U4773 (N_4773,N_2088,N_197);
nand U4774 (N_4774,N_888,N_2210);
and U4775 (N_4775,N_303,N_691);
nand U4776 (N_4776,N_554,N_1451);
and U4777 (N_4777,N_958,N_705);
or U4778 (N_4778,N_347,N_1524);
nand U4779 (N_4779,N_88,N_9);
nor U4780 (N_4780,N_2271,N_1360);
or U4781 (N_4781,N_1354,N_2196);
or U4782 (N_4782,N_1273,N_2341);
or U4783 (N_4783,N_1282,N_1673);
nand U4784 (N_4784,N_1715,N_1287);
or U4785 (N_4785,N_1672,N_906);
nand U4786 (N_4786,N_1959,N_413);
nor U4787 (N_4787,N_1419,N_1912);
nor U4788 (N_4788,N_1492,N_1781);
or U4789 (N_4789,N_2425,N_1676);
and U4790 (N_4790,N_1915,N_1829);
or U4791 (N_4791,N_885,N_1910);
nand U4792 (N_4792,N_564,N_2173);
or U4793 (N_4793,N_642,N_1216);
nor U4794 (N_4794,N_1036,N_2095);
nand U4795 (N_4795,N_1048,N_86);
and U4796 (N_4796,N_579,N_1013);
or U4797 (N_4797,N_1699,N_2477);
and U4798 (N_4798,N_1275,N_1140);
and U4799 (N_4799,N_1292,N_526);
nor U4800 (N_4800,N_784,N_2146);
nor U4801 (N_4801,N_1591,N_1063);
nor U4802 (N_4802,N_1328,N_1105);
or U4803 (N_4803,N_1926,N_1023);
and U4804 (N_4804,N_1032,N_182);
and U4805 (N_4805,N_615,N_519);
nor U4806 (N_4806,N_1321,N_31);
nand U4807 (N_4807,N_2168,N_1682);
nand U4808 (N_4808,N_1481,N_1431);
nand U4809 (N_4809,N_1461,N_172);
or U4810 (N_4810,N_2349,N_878);
nand U4811 (N_4811,N_2392,N_36);
or U4812 (N_4812,N_734,N_2047);
and U4813 (N_4813,N_807,N_1153);
nor U4814 (N_4814,N_1228,N_1017);
and U4815 (N_4815,N_1098,N_2496);
nor U4816 (N_4816,N_1816,N_792);
or U4817 (N_4817,N_1737,N_1376);
nor U4818 (N_4818,N_1829,N_1231);
nand U4819 (N_4819,N_504,N_242);
nor U4820 (N_4820,N_160,N_1880);
nand U4821 (N_4821,N_2298,N_522);
nand U4822 (N_4822,N_446,N_2333);
nand U4823 (N_4823,N_1086,N_21);
and U4824 (N_4824,N_766,N_1125);
nand U4825 (N_4825,N_1160,N_229);
or U4826 (N_4826,N_827,N_502);
nand U4827 (N_4827,N_296,N_1719);
or U4828 (N_4828,N_899,N_2412);
and U4829 (N_4829,N_1736,N_270);
and U4830 (N_4830,N_810,N_262);
and U4831 (N_4831,N_2467,N_394);
nor U4832 (N_4832,N_418,N_524);
or U4833 (N_4833,N_2338,N_940);
nand U4834 (N_4834,N_111,N_1156);
or U4835 (N_4835,N_270,N_1033);
nor U4836 (N_4836,N_1545,N_615);
nand U4837 (N_4837,N_2151,N_2035);
nor U4838 (N_4838,N_1754,N_511);
or U4839 (N_4839,N_1029,N_2277);
and U4840 (N_4840,N_1601,N_407);
nand U4841 (N_4841,N_386,N_353);
nand U4842 (N_4842,N_906,N_2344);
or U4843 (N_4843,N_1305,N_1447);
or U4844 (N_4844,N_897,N_1132);
and U4845 (N_4845,N_1294,N_1071);
and U4846 (N_4846,N_338,N_1540);
nand U4847 (N_4847,N_159,N_548);
nand U4848 (N_4848,N_2243,N_908);
nand U4849 (N_4849,N_2192,N_1771);
nor U4850 (N_4850,N_453,N_179);
nand U4851 (N_4851,N_1969,N_852);
and U4852 (N_4852,N_716,N_1187);
nor U4853 (N_4853,N_1773,N_1804);
nand U4854 (N_4854,N_22,N_256);
or U4855 (N_4855,N_546,N_2448);
nand U4856 (N_4856,N_145,N_987);
or U4857 (N_4857,N_152,N_1646);
or U4858 (N_4858,N_2321,N_1891);
and U4859 (N_4859,N_1599,N_2041);
nand U4860 (N_4860,N_295,N_1129);
nand U4861 (N_4861,N_221,N_678);
nor U4862 (N_4862,N_1354,N_772);
nor U4863 (N_4863,N_1502,N_1018);
nor U4864 (N_4864,N_379,N_611);
and U4865 (N_4865,N_1621,N_1927);
nor U4866 (N_4866,N_1924,N_1247);
nand U4867 (N_4867,N_1436,N_1774);
or U4868 (N_4868,N_523,N_829);
nor U4869 (N_4869,N_1265,N_1098);
nand U4870 (N_4870,N_2354,N_647);
or U4871 (N_4871,N_1616,N_256);
nand U4872 (N_4872,N_2247,N_1990);
nor U4873 (N_4873,N_341,N_1412);
nand U4874 (N_4874,N_223,N_993);
nor U4875 (N_4875,N_566,N_2362);
nand U4876 (N_4876,N_1261,N_1210);
nor U4877 (N_4877,N_304,N_1221);
nor U4878 (N_4878,N_235,N_2445);
or U4879 (N_4879,N_903,N_2438);
nand U4880 (N_4880,N_2293,N_826);
and U4881 (N_4881,N_1212,N_2079);
or U4882 (N_4882,N_913,N_351);
or U4883 (N_4883,N_2158,N_1536);
or U4884 (N_4884,N_1608,N_2002);
nor U4885 (N_4885,N_2204,N_1123);
nand U4886 (N_4886,N_501,N_265);
and U4887 (N_4887,N_2079,N_879);
or U4888 (N_4888,N_1787,N_1477);
nand U4889 (N_4889,N_210,N_308);
and U4890 (N_4890,N_1649,N_997);
nor U4891 (N_4891,N_1619,N_970);
or U4892 (N_4892,N_2403,N_2247);
nor U4893 (N_4893,N_1583,N_278);
or U4894 (N_4894,N_1580,N_1062);
nor U4895 (N_4895,N_1984,N_1402);
nor U4896 (N_4896,N_2214,N_1398);
and U4897 (N_4897,N_741,N_2390);
nor U4898 (N_4898,N_2055,N_1019);
or U4899 (N_4899,N_1565,N_2077);
and U4900 (N_4900,N_2475,N_1576);
or U4901 (N_4901,N_395,N_93);
and U4902 (N_4902,N_1672,N_705);
or U4903 (N_4903,N_695,N_247);
nor U4904 (N_4904,N_1097,N_1703);
or U4905 (N_4905,N_287,N_1776);
nand U4906 (N_4906,N_2056,N_164);
or U4907 (N_4907,N_574,N_2273);
nor U4908 (N_4908,N_1345,N_1771);
nand U4909 (N_4909,N_1795,N_132);
and U4910 (N_4910,N_1963,N_1671);
and U4911 (N_4911,N_2395,N_1366);
nor U4912 (N_4912,N_1440,N_1258);
nand U4913 (N_4913,N_26,N_873);
and U4914 (N_4914,N_897,N_743);
nand U4915 (N_4915,N_987,N_635);
or U4916 (N_4916,N_2239,N_126);
or U4917 (N_4917,N_1358,N_778);
or U4918 (N_4918,N_2002,N_1629);
or U4919 (N_4919,N_600,N_143);
xnor U4920 (N_4920,N_719,N_1273);
or U4921 (N_4921,N_152,N_1015);
and U4922 (N_4922,N_1895,N_2009);
nor U4923 (N_4923,N_1997,N_154);
nor U4924 (N_4924,N_222,N_2172);
and U4925 (N_4925,N_1647,N_178);
and U4926 (N_4926,N_1071,N_2311);
nor U4927 (N_4927,N_1759,N_397);
and U4928 (N_4928,N_299,N_809);
and U4929 (N_4929,N_987,N_830);
and U4930 (N_4930,N_29,N_1638);
or U4931 (N_4931,N_101,N_1805);
nor U4932 (N_4932,N_351,N_1192);
or U4933 (N_4933,N_592,N_1087);
nand U4934 (N_4934,N_1917,N_2276);
or U4935 (N_4935,N_539,N_1290);
and U4936 (N_4936,N_1132,N_2266);
nand U4937 (N_4937,N_44,N_848);
and U4938 (N_4938,N_458,N_876);
xnor U4939 (N_4939,N_1135,N_1107);
or U4940 (N_4940,N_2022,N_1530);
nand U4941 (N_4941,N_597,N_2082);
or U4942 (N_4942,N_2224,N_1670);
or U4943 (N_4943,N_1895,N_56);
nand U4944 (N_4944,N_2498,N_15);
nand U4945 (N_4945,N_1306,N_824);
or U4946 (N_4946,N_865,N_43);
nand U4947 (N_4947,N_2414,N_2127);
nand U4948 (N_4948,N_1732,N_1709);
nand U4949 (N_4949,N_2496,N_1688);
and U4950 (N_4950,N_1038,N_38);
nor U4951 (N_4951,N_1134,N_1120);
nand U4952 (N_4952,N_2242,N_333);
nor U4953 (N_4953,N_2086,N_642);
and U4954 (N_4954,N_179,N_934);
nor U4955 (N_4955,N_407,N_1004);
and U4956 (N_4956,N_1512,N_2204);
or U4957 (N_4957,N_349,N_2410);
or U4958 (N_4958,N_2004,N_1344);
xnor U4959 (N_4959,N_411,N_2204);
nand U4960 (N_4960,N_1851,N_1700);
or U4961 (N_4961,N_1164,N_2246);
and U4962 (N_4962,N_560,N_2020);
and U4963 (N_4963,N_376,N_622);
or U4964 (N_4964,N_1111,N_2140);
nand U4965 (N_4965,N_957,N_154);
and U4966 (N_4966,N_2187,N_963);
nand U4967 (N_4967,N_1394,N_171);
and U4968 (N_4968,N_144,N_782);
nand U4969 (N_4969,N_2327,N_82);
or U4970 (N_4970,N_1426,N_204);
nor U4971 (N_4971,N_1378,N_1839);
nor U4972 (N_4972,N_1749,N_1540);
and U4973 (N_4973,N_409,N_1876);
or U4974 (N_4974,N_1634,N_1013);
and U4975 (N_4975,N_122,N_1582);
and U4976 (N_4976,N_2459,N_1257);
nand U4977 (N_4977,N_2231,N_940);
nor U4978 (N_4978,N_1022,N_1115);
and U4979 (N_4979,N_1010,N_2350);
nor U4980 (N_4980,N_1028,N_127);
nand U4981 (N_4981,N_109,N_780);
and U4982 (N_4982,N_70,N_1614);
or U4983 (N_4983,N_2063,N_566);
or U4984 (N_4984,N_1039,N_1312);
or U4985 (N_4985,N_1951,N_835);
nand U4986 (N_4986,N_222,N_2418);
nand U4987 (N_4987,N_1023,N_509);
xnor U4988 (N_4988,N_1895,N_1256);
nor U4989 (N_4989,N_2046,N_1409);
nor U4990 (N_4990,N_2438,N_1509);
and U4991 (N_4991,N_853,N_955);
or U4992 (N_4992,N_1202,N_2198);
and U4993 (N_4993,N_55,N_1210);
nor U4994 (N_4994,N_1346,N_509);
and U4995 (N_4995,N_388,N_1594);
nor U4996 (N_4996,N_648,N_2103);
and U4997 (N_4997,N_693,N_1964);
and U4998 (N_4998,N_895,N_0);
nor U4999 (N_4999,N_1650,N_1130);
nor UO_0 (O_0,N_3767,N_4506);
nand UO_1 (O_1,N_4931,N_4496);
nor UO_2 (O_2,N_3395,N_4300);
or UO_3 (O_3,N_4198,N_2822);
and UO_4 (O_4,N_2624,N_3506);
and UO_5 (O_5,N_3037,N_4233);
nand UO_6 (O_6,N_4833,N_2987);
nor UO_7 (O_7,N_4392,N_3822);
and UO_8 (O_8,N_3363,N_4991);
or UO_9 (O_9,N_2595,N_4531);
or UO_10 (O_10,N_4159,N_3155);
nor UO_11 (O_11,N_2613,N_2729);
or UO_12 (O_12,N_4431,N_3493);
and UO_13 (O_13,N_4465,N_4718);
nand UO_14 (O_14,N_3089,N_3331);
nor UO_15 (O_15,N_4428,N_4532);
and UO_16 (O_16,N_2940,N_3518);
nor UO_17 (O_17,N_4345,N_3035);
and UO_18 (O_18,N_3367,N_2852);
nor UO_19 (O_19,N_3733,N_4761);
and UO_20 (O_20,N_2686,N_4341);
and UO_21 (O_21,N_2641,N_2976);
nor UO_22 (O_22,N_4426,N_2582);
nand UO_23 (O_23,N_4390,N_3594);
nor UO_24 (O_24,N_3620,N_3722);
nor UO_25 (O_25,N_3311,N_2887);
and UO_26 (O_26,N_3227,N_4348);
or UO_27 (O_27,N_4331,N_4443);
and UO_28 (O_28,N_3344,N_4340);
and UO_29 (O_29,N_4639,N_4652);
or UO_30 (O_30,N_4635,N_4307);
and UO_31 (O_31,N_4859,N_2732);
and UO_32 (O_32,N_2788,N_2916);
nand UO_33 (O_33,N_3102,N_3883);
and UO_34 (O_34,N_2522,N_4296);
and UO_35 (O_35,N_3081,N_4056);
nor UO_36 (O_36,N_4958,N_4544);
nor UO_37 (O_37,N_3739,N_4378);
or UO_38 (O_38,N_2751,N_3449);
and UO_39 (O_39,N_3659,N_4979);
nand UO_40 (O_40,N_4194,N_4035);
or UO_41 (O_41,N_2771,N_2651);
and UO_42 (O_42,N_4004,N_4196);
nand UO_43 (O_43,N_4369,N_4806);
or UO_44 (O_44,N_2925,N_2981);
and UO_45 (O_45,N_4642,N_2800);
or UO_46 (O_46,N_4987,N_3434);
and UO_47 (O_47,N_4608,N_3624);
or UO_48 (O_48,N_2570,N_3125);
and UO_49 (O_49,N_2529,N_4423);
or UO_50 (O_50,N_4302,N_3450);
and UO_51 (O_51,N_3663,N_3926);
xnor UO_52 (O_52,N_2539,N_3191);
nor UO_53 (O_53,N_3831,N_4155);
nand UO_54 (O_54,N_3119,N_3800);
and UO_55 (O_55,N_4411,N_3452);
and UO_56 (O_56,N_3211,N_3783);
nor UO_57 (O_57,N_2875,N_2813);
nor UO_58 (O_58,N_4006,N_2650);
nor UO_59 (O_59,N_3963,N_3480);
nor UO_60 (O_60,N_3207,N_2605);
or UO_61 (O_61,N_3684,N_3478);
or UO_62 (O_62,N_3036,N_4212);
or UO_63 (O_63,N_3007,N_2511);
or UO_64 (O_64,N_3772,N_4962);
nand UO_65 (O_65,N_4678,N_4742);
nand UO_66 (O_66,N_4589,N_3666);
nor UO_67 (O_67,N_4824,N_4151);
nand UO_68 (O_68,N_2927,N_2747);
nor UO_69 (O_69,N_4550,N_3928);
nor UO_70 (O_70,N_3676,N_4880);
or UO_71 (O_71,N_3246,N_3939);
and UO_72 (O_72,N_2520,N_3292);
or UO_73 (O_73,N_4269,N_3027);
nor UO_74 (O_74,N_3163,N_3135);
nand UO_75 (O_75,N_3188,N_3022);
and UO_76 (O_76,N_3499,N_4665);
nand UO_77 (O_77,N_3929,N_4921);
nand UO_78 (O_78,N_3203,N_3466);
nor UO_79 (O_79,N_3404,N_3534);
and UO_80 (O_80,N_4282,N_3795);
nand UO_81 (O_81,N_4590,N_3245);
nand UO_82 (O_82,N_4586,N_4808);
or UO_83 (O_83,N_3023,N_2821);
nor UO_84 (O_84,N_2778,N_2629);
and UO_85 (O_85,N_3077,N_4068);
nor UO_86 (O_86,N_2514,N_4869);
or UO_87 (O_87,N_3740,N_3540);
and UO_88 (O_88,N_3228,N_3491);
and UO_89 (O_89,N_3781,N_4516);
or UO_90 (O_90,N_3379,N_4003);
nor UO_91 (O_91,N_3157,N_4528);
and UO_92 (O_92,N_3215,N_4045);
and UO_93 (O_93,N_4055,N_3403);
nor UO_94 (O_94,N_3026,N_3849);
and UO_95 (O_95,N_3940,N_3096);
and UO_96 (O_96,N_4821,N_2691);
nand UO_97 (O_97,N_4916,N_4304);
nor UO_98 (O_98,N_2992,N_4144);
nor UO_99 (O_99,N_2979,N_4355);
nor UO_100 (O_100,N_4583,N_3786);
nor UO_101 (O_101,N_3107,N_4247);
nor UO_102 (O_102,N_4137,N_4243);
nor UO_103 (O_103,N_3932,N_3802);
and UO_104 (O_104,N_2931,N_4863);
nand UO_105 (O_105,N_2742,N_3811);
nand UO_106 (O_106,N_4146,N_3585);
nand UO_107 (O_107,N_4016,N_3523);
nor UO_108 (O_108,N_4436,N_3193);
nor UO_109 (O_109,N_4569,N_4339);
nor UO_110 (O_110,N_4103,N_3714);
nand UO_111 (O_111,N_3974,N_3583);
or UO_112 (O_112,N_4273,N_4112);
nand UO_113 (O_113,N_2572,N_4645);
nand UO_114 (O_114,N_3437,N_4142);
or UO_115 (O_115,N_4005,N_4126);
nor UO_116 (O_116,N_2921,N_3660);
nor UO_117 (O_117,N_4845,N_3182);
or UO_118 (O_118,N_4053,N_3042);
or UO_119 (O_119,N_3369,N_4083);
nor UO_120 (O_120,N_4353,N_4107);
and UO_121 (O_121,N_2560,N_2664);
nor UO_122 (O_122,N_3314,N_4794);
nor UO_123 (O_123,N_4623,N_3732);
and UO_124 (O_124,N_2748,N_2820);
and UO_125 (O_125,N_3346,N_2574);
nand UO_126 (O_126,N_2612,N_4710);
and UO_127 (O_127,N_2917,N_3580);
nor UO_128 (O_128,N_3436,N_4661);
and UO_129 (O_129,N_4322,N_3815);
and UO_130 (O_130,N_3753,N_4260);
and UO_131 (O_131,N_2885,N_3962);
and UO_132 (O_132,N_3504,N_3819);
nand UO_133 (O_133,N_3006,N_4755);
or UO_134 (O_134,N_4626,N_2886);
and UO_135 (O_135,N_3578,N_3957);
and UO_136 (O_136,N_3244,N_4701);
nand UO_137 (O_137,N_3356,N_3549);
or UO_138 (O_138,N_4250,N_3330);
nand UO_139 (O_139,N_3601,N_4604);
and UO_140 (O_140,N_4121,N_4847);
nand UO_141 (O_141,N_3003,N_2780);
nor UO_142 (O_142,N_2505,N_2578);
nand UO_143 (O_143,N_3754,N_3040);
nor UO_144 (O_144,N_4058,N_3643);
nor UO_145 (O_145,N_4326,N_3117);
or UO_146 (O_146,N_4099,N_3074);
nand UO_147 (O_147,N_4001,N_2884);
nand UO_148 (O_148,N_2654,N_3179);
nor UO_149 (O_149,N_3025,N_3969);
nand UO_150 (O_150,N_4415,N_2656);
nand UO_151 (O_151,N_3855,N_4765);
and UO_152 (O_152,N_2894,N_4416);
nand UO_153 (O_153,N_2835,N_3736);
nor UO_154 (O_154,N_2839,N_3586);
or UO_155 (O_155,N_4309,N_4807);
nor UO_156 (O_156,N_3072,N_4207);
or UO_157 (O_157,N_4796,N_3956);
and UO_158 (O_158,N_3353,N_4657);
nand UO_159 (O_159,N_4213,N_4048);
nand UO_160 (O_160,N_3977,N_3464);
nor UO_161 (O_161,N_4787,N_2846);
and UO_162 (O_162,N_2971,N_2557);
and UO_163 (O_163,N_3995,N_4454);
nand UO_164 (O_164,N_3641,N_3280);
nand UO_165 (O_165,N_4644,N_3374);
nor UO_166 (O_166,N_2934,N_4317);
nand UO_167 (O_167,N_3256,N_3275);
nand UO_168 (O_168,N_3556,N_4948);
and UO_169 (O_169,N_3285,N_3630);
and UO_170 (O_170,N_2939,N_4104);
or UO_171 (O_171,N_4747,N_4802);
nor UO_172 (O_172,N_3304,N_4980);
xor UO_173 (O_173,N_3299,N_4579);
and UO_174 (O_174,N_3655,N_4762);
nand UO_175 (O_175,N_2974,N_2907);
nand UO_176 (O_176,N_3085,N_2869);
nor UO_177 (O_177,N_3172,N_2551);
and UO_178 (O_178,N_3797,N_2982);
nor UO_179 (O_179,N_3734,N_3345);
and UO_180 (O_180,N_2502,N_3868);
or UO_181 (O_181,N_2622,N_2723);
nand UO_182 (O_182,N_3731,N_2958);
or UO_183 (O_183,N_4210,N_2797);
nand UO_184 (O_184,N_3804,N_4776);
nand UO_185 (O_185,N_3958,N_3406);
and UO_186 (O_186,N_2763,N_3692);
and UO_187 (O_187,N_4404,N_4983);
or UO_188 (O_188,N_4387,N_4556);
nor UO_189 (O_189,N_2777,N_4630);
nor UO_190 (O_190,N_3848,N_4412);
nand UO_191 (O_191,N_2893,N_3286);
nor UO_192 (O_192,N_4741,N_4929);
or UO_193 (O_193,N_3725,N_4752);
and UO_194 (O_194,N_4923,N_3834);
or UO_195 (O_195,N_4994,N_2883);
nor UO_196 (O_196,N_2781,N_3923);
nand UO_197 (O_197,N_3393,N_3278);
or UO_198 (O_198,N_4568,N_4643);
or UO_199 (O_199,N_3882,N_4649);
or UO_200 (O_200,N_4621,N_4080);
or UO_201 (O_201,N_4085,N_3837);
nor UO_202 (O_202,N_4989,N_4219);
or UO_203 (O_203,N_4344,N_4181);
nand UO_204 (O_204,N_3779,N_4864);
or UO_205 (O_205,N_3593,N_4834);
and UO_206 (O_206,N_4699,N_4704);
nor UO_207 (O_207,N_2662,N_3749);
or UO_208 (O_208,N_4777,N_3514);
or UO_209 (O_209,N_2558,N_4512);
nor UO_210 (O_210,N_3453,N_4633);
nand UO_211 (O_211,N_3381,N_2911);
nor UO_212 (O_212,N_4240,N_4203);
nand UO_213 (O_213,N_3230,N_4954);
or UO_214 (O_214,N_4206,N_4084);
nand UO_215 (O_215,N_4374,N_3495);
nand UO_216 (O_216,N_2825,N_3142);
and UO_217 (O_217,N_3571,N_4638);
nor UO_218 (O_218,N_3621,N_2997);
nand UO_219 (O_219,N_4349,N_4305);
nor UO_220 (O_220,N_3185,N_2515);
nor UO_221 (O_221,N_3647,N_3606);
nor UO_222 (O_222,N_3043,N_3844);
nand UO_223 (O_223,N_3942,N_3093);
nor UO_224 (O_224,N_3552,N_3252);
nand UO_225 (O_225,N_2577,N_3948);
and UO_226 (O_226,N_4047,N_2610);
nand UO_227 (O_227,N_3289,N_2590);
nor UO_228 (O_228,N_2644,N_2736);
or UO_229 (O_229,N_3200,N_4050);
or UO_230 (O_230,N_4095,N_4127);
nor UO_231 (O_231,N_4012,N_4458);
and UO_232 (O_232,N_3274,N_2585);
or UO_233 (O_233,N_4422,N_4848);
or UO_234 (O_234,N_4558,N_3067);
nor UO_235 (O_235,N_2961,N_2843);
or UO_236 (O_236,N_3922,N_3564);
nand UO_237 (O_237,N_4860,N_3052);
nand UO_238 (O_238,N_4354,N_2616);
nor UO_239 (O_239,N_2637,N_3156);
nor UO_240 (O_240,N_4258,N_3505);
or UO_241 (O_241,N_4238,N_2579);
nor UO_242 (O_242,N_4281,N_4602);
nand UO_243 (O_243,N_3521,N_3796);
and UO_244 (O_244,N_3116,N_3747);
nand UO_245 (O_245,N_4136,N_4907);
or UO_246 (O_246,N_2745,N_4503);
and UO_247 (O_247,N_2547,N_4509);
and UO_248 (O_248,N_4253,N_3174);
or UO_249 (O_249,N_3691,N_3303);
xnor UO_250 (O_250,N_2703,N_2943);
and UO_251 (O_251,N_2640,N_3685);
nand UO_252 (O_252,N_2532,N_4396);
nor UO_253 (O_253,N_3638,N_3937);
and UO_254 (O_254,N_2581,N_3821);
nand UO_255 (O_255,N_3924,N_4541);
or UO_256 (O_256,N_4199,N_2914);
nand UO_257 (O_257,N_2775,N_4896);
nor UO_258 (O_258,N_3129,N_4195);
or UO_259 (O_259,N_3183,N_2829);
nor UO_260 (O_260,N_2874,N_3843);
or UO_261 (O_261,N_3476,N_3916);
nand UO_262 (O_262,N_4707,N_3909);
and UO_263 (O_263,N_3675,N_3212);
and UO_264 (O_264,N_4543,N_3204);
or UO_265 (O_265,N_4469,N_4061);
nand UO_266 (O_266,N_4306,N_2833);
nand UO_267 (O_267,N_2812,N_3526);
and UO_268 (O_268,N_3765,N_4342);
and UO_269 (O_269,N_4380,N_3064);
nand UO_270 (O_270,N_3336,N_2740);
nor UO_271 (O_271,N_2692,N_4168);
and UO_272 (O_272,N_3858,N_3349);
nor UO_273 (O_273,N_3548,N_4211);
nand UO_274 (O_274,N_3118,N_4030);
nor UO_275 (O_275,N_3056,N_3799);
and UO_276 (O_276,N_4798,N_3288);
nand UO_277 (O_277,N_3972,N_3284);
and UO_278 (O_278,N_3865,N_4321);
nor UO_279 (O_279,N_3176,N_4255);
or UO_280 (O_280,N_4620,N_4793);
and UO_281 (O_281,N_3306,N_2945);
nor UO_282 (O_282,N_2752,N_4072);
nor UO_283 (O_283,N_3999,N_3435);
or UO_284 (O_284,N_3880,N_2699);
or UO_285 (O_285,N_4472,N_3904);
nor UO_286 (O_286,N_4715,N_4483);
or UO_287 (O_287,N_4116,N_4691);
or UO_288 (O_288,N_2968,N_2701);
and UO_289 (O_289,N_2550,N_3291);
or UO_290 (O_290,N_4385,N_4185);
or UO_291 (O_291,N_4890,N_4417);
and UO_292 (O_292,N_3058,N_4517);
or UO_293 (O_293,N_4031,N_3519);
and UO_294 (O_294,N_4312,N_4682);
nand UO_295 (O_295,N_2737,N_3983);
nand UO_296 (O_296,N_3399,N_3098);
or UO_297 (O_297,N_4732,N_2888);
and UO_298 (O_298,N_4425,N_3993);
and UO_299 (O_299,N_3017,N_3887);
nand UO_300 (O_300,N_2571,N_2554);
nor UO_301 (O_301,N_3508,N_2783);
nand UO_302 (O_302,N_3616,N_3354);
nor UO_303 (O_303,N_4202,N_4427);
or UO_304 (O_304,N_2678,N_2841);
nand UO_305 (O_305,N_2826,N_4365);
or UO_306 (O_306,N_2831,N_2633);
nor UO_307 (O_307,N_2635,N_2615);
or UO_308 (O_308,N_4363,N_2630);
nand UO_309 (O_309,N_3863,N_3820);
or UO_310 (O_310,N_4401,N_4837);
nor UO_311 (O_311,N_2562,N_3857);
and UO_312 (O_312,N_3300,N_4632);
nor UO_313 (O_313,N_4887,N_3699);
and UO_314 (O_314,N_4537,N_3196);
or UO_315 (O_315,N_2724,N_3944);
and UO_316 (O_316,N_4686,N_3459);
nor UO_317 (O_317,N_4395,N_3132);
and UO_318 (O_318,N_2533,N_2895);
nand UO_319 (O_319,N_4601,N_2796);
or UO_320 (O_320,N_2638,N_4235);
xnor UO_321 (O_321,N_4519,N_4337);
nand UO_322 (O_322,N_3744,N_4889);
and UO_323 (O_323,N_2568,N_4598);
nor UO_324 (O_324,N_4779,N_3808);
and UO_325 (O_325,N_3730,N_4856);
nor UO_326 (O_326,N_3968,N_4858);
nor UO_327 (O_327,N_4285,N_3010);
nand UO_328 (O_328,N_4542,N_4775);
nor UO_329 (O_329,N_3133,N_2989);
or UO_330 (O_330,N_4150,N_3294);
nand UO_331 (O_331,N_4381,N_3839);
nand UO_332 (O_332,N_2501,N_3233);
or UO_333 (O_333,N_3847,N_4578);
or UO_334 (O_334,N_3591,N_4580);
or UO_335 (O_335,N_3325,N_3386);
and UO_336 (O_336,N_3590,N_4275);
nand UO_337 (O_337,N_4640,N_4631);
and UO_338 (O_338,N_3106,N_2730);
or UO_339 (O_339,N_4504,N_4184);
nor UO_340 (O_340,N_3359,N_2566);
nand UO_341 (O_341,N_3458,N_4972);
or UO_342 (O_342,N_3422,N_2565);
nor UO_343 (O_343,N_3921,N_3716);
nand UO_344 (O_344,N_4766,N_2913);
or UO_345 (O_345,N_2779,N_3355);
nand UO_346 (O_346,N_2743,N_3342);
and UO_347 (O_347,N_3710,N_3217);
or UO_348 (O_348,N_3870,N_4036);
and UO_349 (O_349,N_3376,N_4093);
or UO_350 (O_350,N_2970,N_2591);
nand UO_351 (O_351,N_3260,N_4555);
nor UO_352 (O_352,N_3167,N_4231);
nand UO_353 (O_353,N_4825,N_2672);
or UO_354 (O_354,N_3894,N_4216);
or UO_355 (O_355,N_4904,N_4062);
nor UO_356 (O_356,N_4738,N_2768);
or UO_357 (O_357,N_4467,N_4278);
nand UO_358 (O_358,N_3712,N_3525);
and UO_359 (O_359,N_3105,N_3761);
or UO_360 (O_360,N_2891,N_2543);
nand UO_361 (O_361,N_3978,N_2504);
nand UO_362 (O_362,N_4161,N_3041);
or UO_363 (O_363,N_4624,N_3810);
nand UO_364 (O_364,N_4335,N_3757);
nor UO_365 (O_365,N_3189,N_2698);
or UO_366 (O_366,N_3689,N_3219);
nand UO_367 (O_367,N_3418,N_3907);
or UO_368 (O_368,N_3454,N_2966);
and UO_369 (O_369,N_4019,N_3210);
and UO_370 (O_370,N_3127,N_4424);
nor UO_371 (O_371,N_4810,N_2876);
nor UO_372 (O_372,N_4313,N_4187);
or UO_373 (O_373,N_4172,N_3490);
nand UO_374 (O_374,N_3618,N_3413);
nand UO_375 (O_375,N_2948,N_3014);
nor UO_376 (O_376,N_4523,N_3764);
nand UO_377 (O_377,N_4875,N_3777);
nand UO_378 (O_378,N_4057,N_3520);
nor UO_379 (O_379,N_4854,N_4754);
and UO_380 (O_380,N_3788,N_2870);
or UO_381 (O_381,N_4913,N_3087);
xnor UO_382 (O_382,N_3411,N_3720);
nand UO_383 (O_383,N_3323,N_3656);
and UO_384 (O_384,N_4986,N_4222);
and UO_385 (O_385,N_3546,N_4841);
and UO_386 (O_386,N_4595,N_4208);
and UO_387 (O_387,N_4049,N_4284);
nor UO_388 (O_388,N_4158,N_2994);
and UO_389 (O_389,N_3329,N_3134);
nor UO_390 (O_390,N_3611,N_3456);
and UO_391 (O_391,N_4367,N_2518);
and UO_392 (O_392,N_4597,N_4946);
nand UO_393 (O_393,N_4359,N_2964);
nor UO_394 (O_394,N_3442,N_3465);
and UO_395 (O_395,N_2892,N_3164);
nand UO_396 (O_396,N_3979,N_2947);
nand UO_397 (O_397,N_3131,N_4071);
and UO_398 (O_398,N_4215,N_3263);
nand UO_399 (O_399,N_3735,N_4581);
and UO_400 (O_400,N_4725,N_3084);
nor UO_401 (O_401,N_2848,N_4566);
nand UO_402 (O_402,N_4376,N_2942);
or UO_403 (O_403,N_4629,N_4486);
or UO_404 (O_404,N_2817,N_3044);
nor UO_405 (O_405,N_3619,N_4494);
nand UO_406 (O_406,N_2636,N_4835);
nor UO_407 (O_407,N_2794,N_4527);
and UO_408 (O_408,N_3139,N_4009);
nor UO_409 (O_409,N_3897,N_3690);
or UO_410 (O_410,N_3169,N_4310);
nand UO_411 (O_411,N_4485,N_4441);
and UO_412 (O_412,N_3917,N_3090);
nand UO_413 (O_413,N_4745,N_4605);
and UO_414 (O_414,N_4832,N_3852);
nor UO_415 (O_415,N_2537,N_4607);
or UO_416 (O_416,N_3239,N_4694);
or UO_417 (O_417,N_2810,N_4399);
or UO_418 (O_418,N_2584,N_2845);
nor UO_419 (O_419,N_3510,N_4939);
or UO_420 (O_420,N_4592,N_4352);
or UO_421 (O_421,N_3651,N_4830);
nand UO_422 (O_422,N_4283,N_3334);
and UO_423 (O_423,N_3662,N_2955);
nor UO_424 (O_424,N_4903,N_3768);
or UO_425 (O_425,N_2675,N_3428);
or UO_426 (O_426,N_3057,N_4702);
nand UO_427 (O_427,N_4070,N_4421);
nand UO_428 (O_428,N_4134,N_3814);
or UO_429 (O_429,N_3068,N_3190);
nor UO_430 (O_430,N_3111,N_2828);
nand UO_431 (O_431,N_2721,N_2602);
and UO_432 (O_432,N_4377,N_3080);
nand UO_433 (O_433,N_3070,N_3483);
and UO_434 (O_434,N_3533,N_2929);
or UO_435 (O_435,N_3498,N_3047);
or UO_436 (O_436,N_3512,N_4740);
nor UO_437 (O_437,N_2750,N_4239);
nand UO_438 (O_438,N_2899,N_3528);
nand UO_439 (O_439,N_4511,N_3301);
or UO_440 (O_440,N_4758,N_3216);
and UO_441 (O_441,N_4183,N_4695);
or UO_442 (O_442,N_2859,N_4968);
or UO_443 (O_443,N_3264,N_4690);
nand UO_444 (O_444,N_2623,N_4256);
nand UO_445 (O_445,N_4491,N_3824);
or UO_446 (O_446,N_4674,N_2904);
and UO_447 (O_447,N_2513,N_4462);
nand UO_448 (O_448,N_4248,N_2776);
and UO_449 (O_449,N_2712,N_3881);
or UO_450 (O_450,N_4451,N_4011);
or UO_451 (O_451,N_4291,N_2901);
and UO_452 (O_452,N_3576,N_2928);
or UO_453 (O_453,N_3845,N_4547);
and UO_454 (O_454,N_3032,N_2601);
nand UO_455 (O_455,N_3551,N_4025);
xnor UO_456 (O_456,N_4647,N_2647);
nand UO_457 (O_457,N_4364,N_4499);
nand UO_458 (O_458,N_4613,N_4906);
and UO_459 (O_459,N_3364,N_4909);
nor UO_460 (O_460,N_4998,N_3236);
or UO_461 (O_461,N_3910,N_3165);
or UO_462 (O_462,N_2707,N_3298);
nor UO_463 (O_463,N_4088,N_4379);
nand UO_464 (O_464,N_3234,N_4911);
nor UO_465 (O_465,N_3146,N_4370);
or UO_466 (O_466,N_4618,N_2842);
nor UO_467 (O_467,N_4774,N_4672);
nand UO_468 (O_468,N_4942,N_3947);
nor UO_469 (O_469,N_3703,N_3319);
nand UO_470 (O_470,N_3902,N_4188);
nor UO_471 (O_471,N_3588,N_4221);
and UO_472 (O_472,N_3108,N_4703);
nor UO_473 (O_473,N_4562,N_4915);
or UO_474 (O_474,N_4811,N_3835);
or UO_475 (O_475,N_3877,N_4298);
and UO_476 (O_476,N_4023,N_3494);
and UO_477 (O_477,N_4908,N_3574);
nor UO_478 (O_478,N_4165,N_4711);
or UO_479 (O_479,N_3809,N_4028);
or UO_480 (O_480,N_4328,N_3253);
and UO_481 (O_481,N_2738,N_3976);
xnor UO_482 (O_482,N_2983,N_4886);
and UO_483 (O_483,N_3756,N_3634);
or UO_484 (O_484,N_2774,N_4803);
or UO_485 (O_485,N_4470,N_3936);
or UO_486 (O_486,N_4816,N_4245);
and UO_487 (O_487,N_3501,N_3502);
and UO_488 (O_488,N_3864,N_3412);
nand UO_489 (O_489,N_4145,N_3097);
nand UO_490 (O_490,N_3258,N_3697);
nor UO_491 (O_491,N_4132,N_3625);
or UO_492 (O_492,N_4722,N_4726);
and UO_493 (O_493,N_4476,N_2596);
nand UO_494 (O_494,N_4201,N_3082);
xor UO_495 (O_495,N_3816,N_3572);
or UO_496 (O_496,N_2679,N_3401);
nor UO_497 (O_497,N_2922,N_4770);
or UO_498 (O_498,N_3028,N_4109);
nand UO_499 (O_499,N_2527,N_2804);
nor UO_500 (O_500,N_4997,N_4557);
or UO_501 (O_501,N_2795,N_3665);
nor UO_502 (O_502,N_3758,N_2661);
nor UO_503 (O_503,N_2705,N_4435);
nor UO_504 (O_504,N_4224,N_4254);
or UO_505 (O_505,N_3202,N_2766);
and UO_506 (O_506,N_2847,N_4820);
or UO_507 (O_507,N_2660,N_2864);
nor UO_508 (O_508,N_3516,N_3283);
nor UO_509 (O_509,N_3177,N_2592);
nand UO_510 (O_510,N_4474,N_3959);
and UO_511 (O_511,N_4829,N_4564);
nor UO_512 (O_512,N_4495,N_2681);
or UO_513 (O_513,N_3694,N_3287);
nand UO_514 (O_514,N_4677,N_3213);
or UO_515 (O_515,N_2618,N_4153);
and UO_516 (O_516,N_4280,N_3332);
nor UO_517 (O_517,N_4982,N_3024);
and UO_518 (O_518,N_2510,N_3829);
nand UO_519 (O_519,N_3051,N_3595);
nand UO_520 (O_520,N_4999,N_3950);
or UO_521 (O_521,N_3009,N_2741);
nand UO_522 (O_522,N_3417,N_2530);
or UO_523 (O_523,N_3973,N_3013);
nor UO_524 (O_524,N_3985,N_2685);
or UO_525 (O_525,N_4836,N_4698);
nor UO_526 (O_526,N_3012,N_4268);
nor UO_527 (O_527,N_2542,N_2722);
xnor UO_528 (O_528,N_4664,N_2993);
nand UO_529 (O_529,N_2995,N_3876);
nor UO_530 (O_530,N_3933,N_3095);
and UO_531 (O_531,N_4716,N_2754);
nor UO_532 (O_532,N_3751,N_4437);
nor UO_533 (O_533,N_3891,N_3075);
nor UO_534 (O_534,N_3337,N_4501);
nand UO_535 (O_535,N_4560,N_4308);
nand UO_536 (O_536,N_2844,N_4487);
nand UO_537 (O_537,N_3405,N_3099);
or UO_538 (O_538,N_3713,N_3388);
or UO_539 (O_539,N_3608,N_3841);
and UO_540 (O_540,N_2710,N_3715);
nor UO_541 (O_541,N_4293,N_2713);
nand UO_542 (O_542,N_2786,N_3539);
and UO_543 (O_543,N_4565,N_2798);
and UO_544 (O_544,N_4059,N_4670);
or UO_545 (O_545,N_3148,N_2694);
nor UO_546 (O_546,N_4898,N_4481);
nor UO_547 (O_547,N_4606,N_4043);
or UO_548 (O_548,N_4965,N_2586);
or UO_549 (O_549,N_3262,N_2523);
nand UO_550 (O_550,N_3168,N_2648);
and UO_551 (O_551,N_4038,N_3775);
nand UO_552 (O_552,N_4270,N_3402);
nor UO_553 (O_553,N_3078,N_3154);
xnor UO_554 (O_554,N_4801,N_4748);
or UO_555 (O_555,N_2603,N_3706);
or UO_556 (O_556,N_4276,N_3532);
or UO_557 (O_557,N_4819,N_3420);
or UO_558 (O_558,N_3055,N_2653);
nand UO_559 (O_559,N_3180,N_4930);
or UO_560 (O_560,N_3237,N_4933);
and UO_561 (O_561,N_2680,N_3537);
and UO_562 (O_562,N_2658,N_3729);
and UO_563 (O_563,N_4318,N_4628);
nand UO_564 (O_564,N_3711,N_3091);
nand UO_565 (O_565,N_4366,N_3687);
and UO_566 (O_566,N_2868,N_4971);
xnor UO_567 (O_567,N_4660,N_3680);
and UO_568 (O_568,N_4669,N_3535);
and UO_569 (O_569,N_3554,N_3648);
and UO_570 (O_570,N_3063,N_2854);
and UO_571 (O_571,N_2645,N_4950);
and UO_572 (O_572,N_2823,N_4037);
nor UO_573 (O_573,N_3170,N_2642);
and UO_574 (O_574,N_3986,N_4360);
and UO_575 (O_575,N_3315,N_3432);
nand UO_576 (O_576,N_3961,N_4753);
or UO_577 (O_577,N_3599,N_3240);
or UO_578 (O_578,N_3463,N_3214);
xor UO_579 (O_579,N_3147,N_4612);
nor UO_580 (O_580,N_2937,N_3243);
nand UO_581 (O_581,N_4797,N_4967);
or UO_582 (O_582,N_3582,N_4956);
and UO_583 (O_583,N_3873,N_4167);
nand UO_584 (O_584,N_4838,N_2569);
or UO_585 (O_585,N_2657,N_4683);
nand UO_586 (O_586,N_4877,N_3543);
or UO_587 (O_587,N_3197,N_2669);
or UO_588 (O_588,N_4073,N_4885);
nor UO_589 (O_589,N_3030,N_2534);
and UO_590 (O_590,N_4357,N_3793);
or UO_591 (O_591,N_4667,N_3031);
nor UO_592 (O_592,N_4163,N_3584);
or UO_593 (O_593,N_3850,N_3513);
and UO_594 (O_594,N_3991,N_2889);
nor UO_595 (O_595,N_3153,N_3198);
nor UO_596 (O_596,N_2536,N_3677);
nand UO_597 (O_597,N_2599,N_4627);
nand UO_598 (O_598,N_3536,N_4935);
and UO_599 (O_599,N_4789,N_4805);
and UO_600 (O_600,N_3340,N_2957);
nand UO_601 (O_601,N_2716,N_3555);
nand UO_602 (O_602,N_4402,N_4419);
and UO_603 (O_603,N_4782,N_3462);
and UO_604 (O_604,N_2545,N_2784);
and UO_605 (O_605,N_4242,N_4033);
and UO_606 (O_606,N_3205,N_4622);
nor UO_607 (O_607,N_3872,N_4636);
nand UO_608 (O_608,N_2726,N_3249);
nand UO_609 (O_609,N_3890,N_4572);
nor UO_610 (O_610,N_2575,N_3721);
nand UO_611 (O_611,N_4945,N_3201);
nand UO_612 (O_612,N_3199,N_3397);
and UO_613 (O_613,N_4082,N_2588);
nand UO_614 (O_614,N_4574,N_4756);
nand UO_615 (O_615,N_3104,N_2827);
nand UO_616 (O_616,N_4391,N_3527);
nor UO_617 (O_617,N_3482,N_4784);
nor UO_618 (O_618,N_4065,N_3140);
xnor UO_619 (O_619,N_4329,N_4505);
nand UO_620 (O_620,N_2573,N_4105);
nor UO_621 (O_621,N_4449,N_3447);
nor UO_622 (O_622,N_3842,N_4319);
or UO_623 (O_623,N_4540,N_4320);
nand UO_624 (O_624,N_3738,N_4717);
and UO_625 (O_625,N_2773,N_2531);
nand UO_626 (O_626,N_2512,N_4330);
or UO_627 (O_627,N_3522,N_3755);
nand UO_628 (O_628,N_3867,N_3015);
and UO_629 (O_629,N_4271,N_3664);
nor UO_630 (O_630,N_3846,N_2938);
or UO_631 (O_631,N_3679,N_4020);
and UO_632 (O_632,N_2930,N_3241);
or UO_633 (O_633,N_4135,N_3900);
nor UO_634 (O_634,N_2704,N_3339);
nand UO_635 (O_635,N_3748,N_2540);
and UO_636 (O_636,N_3497,N_4205);
or UO_637 (O_637,N_4839,N_4015);
or UO_638 (O_638,N_3238,N_2619);
nand UO_639 (O_639,N_4152,N_2863);
nor UO_640 (O_640,N_4063,N_3550);
or UO_641 (O_641,N_3511,N_4978);
or UO_642 (O_642,N_4383,N_3382);
xor UO_643 (O_643,N_3553,N_4680);
nand UO_644 (O_644,N_4910,N_4479);
nor UO_645 (O_645,N_3467,N_2598);
nand UO_646 (O_646,N_4294,N_3871);
and UO_647 (O_647,N_3784,N_3987);
and UO_648 (O_648,N_4768,N_3602);
nand UO_649 (O_649,N_3054,N_4985);
nor UO_650 (O_650,N_4791,N_4852);
or UO_651 (O_651,N_4386,N_4976);
nor UO_652 (O_652,N_3728,N_4840);
and UO_653 (O_653,N_4658,N_4008);
nor UO_654 (O_654,N_3901,N_3162);
or UO_655 (O_655,N_4535,N_3563);
nor UO_656 (O_656,N_3559,N_4066);
or UO_657 (O_657,N_4409,N_3209);
and UO_658 (O_658,N_4666,N_4881);
nor UO_659 (O_659,N_4102,N_4675);
nand UO_660 (O_660,N_4577,N_2546);
or UO_661 (O_661,N_2559,N_3869);
nor UO_662 (O_662,N_2769,N_4180);
or UO_663 (O_663,N_2728,N_4455);
or UO_664 (O_664,N_4897,N_3529);
or UO_665 (O_665,N_4123,N_4949);
nor UO_666 (O_666,N_2673,N_3076);
or UO_667 (O_667,N_4166,N_4610);
nor UO_668 (O_668,N_3138,N_4279);
nand UO_669 (O_669,N_2744,N_3614);
and UO_670 (O_670,N_4299,N_4489);
xnor UO_671 (O_671,N_2977,N_4862);
nor UO_672 (O_672,N_4778,N_4663);
nor UO_673 (O_673,N_3778,N_4178);
or UO_674 (O_674,N_4493,N_3171);
and UO_675 (O_675,N_3823,N_4162);
nand UO_676 (O_676,N_3682,N_2830);
nor UO_677 (O_677,N_4226,N_2834);
nor UO_678 (O_678,N_3235,N_4953);
and UO_679 (O_679,N_4912,N_4078);
nor UO_680 (O_680,N_4750,N_4229);
and UO_681 (O_681,N_3605,N_3309);
nand UO_682 (O_682,N_2519,N_4619);
or UO_683 (O_683,N_3653,N_3589);
nand UO_684 (O_684,N_4648,N_3470);
and UO_685 (O_685,N_3293,N_3737);
or UO_686 (O_686,N_3103,N_3965);
and UO_687 (O_687,N_4413,N_3224);
or UO_688 (O_688,N_4143,N_4125);
nand UO_689 (O_689,N_3130,N_4034);
or UO_690 (O_690,N_4400,N_3635);
and UO_691 (O_691,N_4094,N_2535);
and UO_692 (O_692,N_3431,N_2665);
and UO_693 (O_693,N_3279,N_3268);
and UO_694 (O_694,N_4044,N_4314);
or UO_695 (O_695,N_4689,N_4917);
or UO_696 (O_696,N_2882,N_2880);
and UO_697 (O_697,N_4876,N_2718);
or UO_698 (O_698,N_3048,N_3383);
nand UO_699 (O_699,N_3423,N_4027);
or UO_700 (O_700,N_4730,N_3899);
and UO_701 (O_701,N_2962,N_2715);
nor UO_702 (O_702,N_3633,N_2507);
or UO_703 (O_703,N_4723,N_3892);
or UO_704 (O_704,N_4014,N_4463);
nor UO_705 (O_705,N_3701,N_2684);
and UO_706 (O_706,N_3874,N_4585);
or UO_707 (O_707,N_3255,N_4138);
nand UO_708 (O_708,N_2700,N_4118);
and UO_709 (O_709,N_4874,N_2871);
and UO_710 (O_710,N_4287,N_4760);
nor UO_711 (O_711,N_4759,N_2801);
nand UO_712 (O_712,N_3833,N_3998);
and UO_713 (O_713,N_3908,N_3484);
nand UO_714 (O_714,N_3746,N_3251);
nor UO_715 (O_715,N_4920,N_3029);
nor UO_716 (O_716,N_4067,N_3457);
nand UO_717 (O_717,N_3092,N_2757);
nand UO_718 (O_718,N_4575,N_3137);
nor UO_719 (O_719,N_3762,N_4809);
or UO_720 (O_720,N_4518,N_4371);
and UO_721 (O_721,N_4173,N_4209);
or UO_722 (O_722,N_2789,N_4899);
or UO_723 (O_723,N_2725,N_3637);
nor UO_724 (O_724,N_3575,N_3607);
and UO_725 (O_725,N_4739,N_3400);
nor UO_726 (O_726,N_3989,N_3970);
or UO_727 (O_727,N_3187,N_4533);
nor UO_728 (O_728,N_3646,N_3375);
and UO_729 (O_729,N_4818,N_3628);
nand UO_730 (O_730,N_3250,N_4323);
nand UO_731 (O_731,N_2614,N_2548);
nand UO_732 (O_732,N_3481,N_4124);
and UO_733 (O_733,N_3062,N_2980);
nand UO_734 (O_734,N_4763,N_3851);
nor UO_735 (O_735,N_3317,N_3221);
nand UO_736 (O_736,N_3424,N_2720);
or UO_737 (O_737,N_4189,N_3538);
nor UO_738 (O_738,N_3745,N_4553);
nand UO_739 (O_739,N_4591,N_2739);
nand UO_740 (O_740,N_4884,N_2991);
nor UO_741 (O_741,N_4176,N_2861);
and UO_742 (O_742,N_3838,N_4154);
nand UO_743 (O_743,N_2996,N_3271);
or UO_744 (O_744,N_4977,N_4405);
or UO_745 (O_745,N_3570,N_3448);
nor UO_746 (O_746,N_3759,N_3971);
nand UO_747 (O_747,N_3573,N_4175);
nor UO_748 (O_748,N_2652,N_4259);
nand UO_749 (O_749,N_3530,N_2663);
and UO_750 (O_750,N_2969,N_4490);
and UO_751 (O_751,N_4720,N_4139);
nand UO_752 (O_752,N_3640,N_3088);
or UO_753 (O_753,N_4653,N_4060);
or UO_754 (O_754,N_3723,N_4656);
nor UO_755 (O_755,N_4545,N_3186);
nand UO_756 (O_756,N_4514,N_4429);
or UO_757 (O_757,N_4446,N_3297);
nor UO_758 (O_758,N_4430,N_4729);
and UO_759 (O_759,N_4459,N_3817);
nor UO_760 (O_760,N_3152,N_4696);
nor UO_761 (O_761,N_4214,N_4567);
nor UO_762 (O_762,N_4944,N_4659);
nand UO_763 (O_763,N_4932,N_3598);
nor UO_764 (O_764,N_4561,N_3039);
nor UO_765 (O_765,N_4551,N_4781);
nor UO_766 (O_766,N_2668,N_3195);
or UO_767 (O_767,N_3474,N_3654);
xnor UO_768 (O_768,N_3994,N_4684);
nand UO_769 (O_769,N_2855,N_4713);
nand UO_770 (O_770,N_3427,N_3545);
nand UO_771 (O_771,N_4074,N_3812);
nor UO_772 (O_772,N_4687,N_2561);
nor UO_773 (O_773,N_4244,N_3769);
or UO_774 (O_774,N_3708,N_2708);
nor UO_775 (O_775,N_3531,N_3489);
and UO_776 (O_776,N_2759,N_3444);
nand UO_777 (O_777,N_4927,N_3008);
nand UO_778 (O_778,N_4671,N_4995);
nor UO_779 (O_779,N_3966,N_3061);
or UO_780 (O_780,N_3446,N_2918);
and UO_781 (O_781,N_4709,N_3707);
nand UO_782 (O_782,N_4191,N_4646);
and UO_783 (O_783,N_4780,N_2950);
nor UO_784 (O_784,N_4111,N_3002);
nand UO_785 (O_785,N_4988,N_3242);
or UO_786 (O_786,N_3964,N_2959);
nor UO_787 (O_787,N_2634,N_3645);
and UO_788 (O_788,N_4098,N_3312);
and UO_789 (O_789,N_4186,N_4692);
and UO_790 (O_790,N_2919,N_4433);
nand UO_791 (O_791,N_2604,N_4744);
nor UO_792 (O_792,N_4092,N_2611);
and UO_793 (O_793,N_4228,N_3310);
nor UO_794 (O_794,N_2553,N_3524);
nand UO_795 (O_795,N_4868,N_4338);
nor UO_796 (O_796,N_4792,N_2549);
nand UO_797 (O_797,N_2593,N_2563);
nand UO_798 (O_798,N_2580,N_3652);
nand UO_799 (O_799,N_3862,N_2952);
nor UO_800 (O_800,N_3798,N_3752);
and UO_801 (O_801,N_4007,N_3113);
and UO_802 (O_802,N_4403,N_2717);
nor UO_803 (O_803,N_2506,N_4480);
nor UO_804 (O_804,N_3282,N_3350);
or UO_805 (O_805,N_3358,N_3561);
and UO_806 (O_806,N_2500,N_4614);
nor UO_807 (O_807,N_4673,N_3128);
nor UO_808 (O_808,N_2865,N_4736);
nand UO_809 (O_809,N_4343,N_3632);
nor UO_810 (O_810,N_4334,N_4879);
and UO_811 (O_811,N_2735,N_3906);
and UO_812 (O_812,N_3357,N_3144);
nor UO_813 (O_813,N_4113,N_4471);
and UO_814 (O_814,N_3912,N_3273);
and UO_815 (O_815,N_3787,N_3079);
or UO_816 (O_816,N_3579,N_3785);
nand UO_817 (O_817,N_4241,N_3160);
nand UO_818 (O_818,N_4498,N_4448);
or UO_819 (O_819,N_3477,N_2808);
or UO_820 (O_820,N_3218,N_4010);
nor UO_821 (O_821,N_3650,N_4964);
or UO_822 (O_822,N_3232,N_3141);
nor UO_823 (O_823,N_2760,N_2973);
nand UO_824 (O_824,N_4823,N_4064);
nand UO_825 (O_825,N_4200,N_4492);
nand UO_826 (O_826,N_3347,N_3384);
or UO_827 (O_827,N_3225,N_3060);
nand UO_828 (O_828,N_4131,N_3938);
and UO_829 (O_829,N_3461,N_3469);
and UO_830 (O_830,N_4955,N_4813);
nor UO_831 (O_831,N_2920,N_3486);
nand UO_832 (O_832,N_4893,N_4096);
or UO_833 (O_833,N_2898,N_3318);
or UO_834 (O_834,N_4177,N_4857);
nand UO_835 (O_835,N_4676,N_3005);
or UO_836 (O_836,N_4947,N_2627);
and UO_837 (O_837,N_2538,N_3389);
nand UO_838 (O_838,N_4957,N_2755);
and UO_839 (O_839,N_3672,N_4444);
nand UO_840 (O_840,N_4700,N_2509);
or UO_841 (O_841,N_3362,N_3394);
and UO_842 (O_842,N_2621,N_2589);
nor UO_843 (O_843,N_3980,N_2932);
nand UO_844 (O_844,N_3990,N_3488);
nor UO_845 (O_845,N_2625,N_4324);
nor UO_846 (O_846,N_3272,N_3750);
and UO_847 (O_847,N_4251,N_4831);
nor UO_848 (O_848,N_2936,N_3818);
or UO_849 (O_849,N_4922,N_3658);
nand UO_850 (O_850,N_4438,N_3370);
and UO_851 (O_851,N_3955,N_4197);
or UO_852 (O_852,N_4905,N_3338);
and UO_853 (O_853,N_3445,N_3915);
nor UO_854 (O_854,N_4693,N_3281);
or UO_855 (O_855,N_3136,N_4981);
nand UO_856 (O_856,N_2850,N_4457);
or UO_857 (O_857,N_4266,N_3678);
or UO_858 (O_858,N_4785,N_3927);
nand UO_859 (O_859,N_2819,N_4075);
nand UO_860 (O_860,N_4190,N_4861);
or UO_861 (O_861,N_3790,N_2912);
nand UO_862 (O_862,N_2985,N_2926);
or UO_863 (O_863,N_4252,N_2836);
and UO_864 (O_864,N_4051,N_3861);
nor UO_865 (O_865,N_4382,N_3905);
nand UO_866 (O_866,N_3669,N_3569);
or UO_867 (O_867,N_4225,N_3792);
nor UO_868 (O_868,N_2666,N_3702);
and UO_869 (O_869,N_3110,N_4362);
nand UO_870 (O_870,N_2516,N_4100);
nand UO_871 (O_871,N_4548,N_4609);
or UO_872 (O_872,N_3161,N_4223);
or UO_873 (O_873,N_3373,N_3276);
nor UO_874 (O_874,N_2881,N_3920);
and UO_875 (O_875,N_4616,N_4286);
and UO_876 (O_876,N_4706,N_3407);
and UO_877 (O_877,N_3409,N_4192);
nor UO_878 (O_878,N_3004,N_4129);
xor UO_879 (O_879,N_3112,N_2900);
and UO_880 (O_880,N_3231,N_2905);
and UO_881 (O_881,N_4488,N_2576);
or UO_882 (O_882,N_3261,N_4130);
nand UO_883 (O_883,N_3951,N_3943);
nand UO_884 (O_884,N_4520,N_3194);
nand UO_885 (O_885,N_3547,N_3623);
and UO_886 (O_886,N_4237,N_3184);
or UO_887 (O_887,N_2544,N_2933);
and UO_888 (O_888,N_4611,N_4358);
and UO_889 (O_889,N_3941,N_3935);
or UO_890 (O_890,N_4866,N_3175);
or UO_891 (O_891,N_2687,N_2944);
and UO_892 (O_892,N_4870,N_4393);
nor UO_893 (O_893,N_3981,N_4262);
nand UO_894 (O_894,N_3875,N_3265);
or UO_895 (O_895,N_4290,N_4257);
or UO_896 (O_896,N_3657,N_3460);
or UO_897 (O_897,N_2782,N_4963);
or UO_898 (O_898,N_4751,N_3717);
nand UO_899 (O_899,N_3509,N_2682);
or UO_900 (O_900,N_4970,N_4712);
or UO_901 (O_901,N_3914,N_3220);
nor UO_902 (O_902,N_2856,N_3604);
nor UO_903 (O_903,N_3568,N_4714);
nand UO_904 (O_904,N_4895,N_4052);
nor UO_905 (O_905,N_4539,N_3667);
and UO_906 (O_906,N_4346,N_3475);
and UO_907 (O_907,N_3996,N_4497);
nand UO_908 (O_908,N_3719,N_4389);
and UO_909 (O_909,N_4460,N_4731);
and UO_910 (O_910,N_4350,N_4466);
and UO_911 (O_911,N_2767,N_4311);
nor UO_912 (O_912,N_3763,N_4475);
and UO_913 (O_913,N_4934,N_2607);
and UO_914 (O_914,N_3949,N_3859);
nand UO_915 (O_915,N_4757,N_2858);
and UO_916 (O_916,N_3515,N_3120);
nor UO_917 (O_917,N_4418,N_3053);
nor UO_918 (O_918,N_4077,N_3742);
and UO_919 (O_919,N_3248,N_3807);
nand UO_920 (O_920,N_4156,N_4026);
nand UO_921 (O_921,N_2862,N_3390);
nor UO_922 (O_922,N_3438,N_4128);
nand UO_923 (O_923,N_2956,N_2807);
or UO_924 (O_924,N_3222,N_2818);
nand UO_925 (O_925,N_4786,N_2753);
and UO_926 (O_926,N_4473,N_3931);
nand UO_927 (O_927,N_4600,N_2879);
nor UO_928 (O_928,N_3780,N_4447);
or UO_929 (O_929,N_3360,N_2954);
nor UO_930 (O_930,N_3988,N_3704);
nand UO_931 (O_931,N_3592,N_4641);
nand UO_932 (O_932,N_3743,N_3609);
or UO_933 (O_933,N_3856,N_2689);
nand UO_934 (O_934,N_2609,N_2541);
and UO_935 (O_935,N_2521,N_4039);
and UO_936 (O_936,N_3408,N_3670);
nand UO_937 (O_937,N_2719,N_4464);
nor UO_938 (O_938,N_4546,N_4871);
nor UO_939 (O_939,N_3327,N_4685);
nor UO_940 (O_940,N_4368,N_3451);
and UO_941 (O_941,N_4795,N_3430);
or UO_942 (O_942,N_3441,N_3813);
nor UO_943 (O_943,N_3114,N_3558);
nor UO_944 (O_944,N_2924,N_2709);
nor UO_945 (O_945,N_3100,N_4993);
or UO_946 (O_946,N_2528,N_2838);
nor UO_947 (O_947,N_4888,N_4599);
and UO_948 (O_948,N_3782,N_4119);
or UO_949 (O_949,N_3507,N_3479);
nor UO_950 (O_950,N_4587,N_3320);
and UO_951 (O_951,N_3277,N_4373);
and UO_952 (O_952,N_4563,N_3305);
and UO_953 (O_953,N_4439,N_4017);
nor UO_954 (O_954,N_4408,N_2674);
or UO_955 (O_955,N_2903,N_3913);
or UO_956 (O_956,N_4990,N_3266);
or UO_957 (O_957,N_4867,N_3109);
or UO_958 (O_958,N_3414,N_3888);
nand UO_959 (O_959,N_2597,N_4737);
nor UO_960 (O_960,N_4617,N_4559);
and UO_961 (O_961,N_3496,N_3472);
nand UO_962 (O_962,N_3934,N_4783);
or UO_963 (O_963,N_3034,N_4800);
nand UO_964 (O_964,N_4406,N_3391);
nor UO_965 (O_965,N_2814,N_3351);
and UO_966 (O_966,N_4530,N_2802);
nand UO_967 (O_967,N_3794,N_3433);
nor UO_968 (O_968,N_3257,N_2902);
nor UO_969 (O_969,N_4969,N_3173);
and UO_970 (O_970,N_3854,N_3673);
and UO_971 (O_971,N_4552,N_4272);
nor UO_972 (O_972,N_4347,N_3945);
or UO_973 (O_973,N_4961,N_2999);
nor UO_974 (O_974,N_3741,N_3021);
nor UO_975 (O_975,N_4434,N_2953);
nor UO_976 (O_976,N_3700,N_4081);
or UO_977 (O_977,N_4900,N_2608);
or UO_978 (O_978,N_2832,N_3122);
nand UO_979 (O_979,N_3343,N_3975);
and UO_980 (O_980,N_4822,N_4453);
nor UO_981 (O_981,N_4507,N_3269);
nor UO_982 (O_982,N_3629,N_2631);
nand UO_983 (O_983,N_4842,N_2975);
nand UO_984 (O_984,N_2984,N_4263);
nor UO_985 (O_985,N_4232,N_2872);
and UO_986 (O_986,N_2809,N_2951);
nor UO_987 (O_987,N_4650,N_3267);
or UO_988 (O_988,N_4938,N_3372);
and UO_989 (O_989,N_3365,N_3639);
or UO_990 (O_990,N_3967,N_4032);
nor UO_991 (O_991,N_2626,N_2867);
and UO_992 (O_992,N_3398,N_2946);
and UO_993 (O_993,N_4315,N_3295);
nor UO_994 (O_994,N_3166,N_2806);
and UO_995 (O_995,N_2702,N_2639);
and UO_996 (O_996,N_3069,N_4728);
and UO_997 (O_997,N_4040,N_3542);
and UO_998 (O_998,N_4106,N_3789);
xnor UO_999 (O_999,N_2749,N_3884);
endmodule