module basic_2000_20000_2500_80_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_230,In_1010);
nor U1 (N_1,In_862,In_1350);
and U2 (N_2,In_749,In_1833);
xnor U3 (N_3,In_393,In_444);
nor U4 (N_4,In_1655,In_650);
or U5 (N_5,In_1349,In_1517);
nor U6 (N_6,In_945,In_461);
nand U7 (N_7,In_1491,In_1120);
or U8 (N_8,In_267,In_1567);
nand U9 (N_9,In_574,In_486);
and U10 (N_10,In_1379,In_928);
nand U11 (N_11,In_703,In_1217);
nand U12 (N_12,In_652,In_364);
nand U13 (N_13,In_481,In_1713);
and U14 (N_14,In_1285,In_1317);
xor U15 (N_15,In_128,In_1970);
or U16 (N_16,In_153,In_1062);
nand U17 (N_17,In_737,In_1661);
and U18 (N_18,In_156,In_398);
nor U19 (N_19,In_431,In_116);
nor U20 (N_20,In_0,In_87);
nor U21 (N_21,In_475,In_1640);
nor U22 (N_22,In_1615,In_1663);
xnor U23 (N_23,In_1590,In_1297);
nor U24 (N_24,In_1321,In_144);
and U25 (N_25,In_534,In_707);
xnor U26 (N_26,In_1277,In_458);
or U27 (N_27,In_729,In_1576);
xor U28 (N_28,In_912,In_428);
or U29 (N_29,In_1323,In_1648);
nor U30 (N_30,In_600,In_584);
or U31 (N_31,In_365,In_1084);
xor U32 (N_32,In_494,In_536);
and U33 (N_33,In_784,In_11);
nand U34 (N_34,In_257,In_66);
and U35 (N_35,In_960,In_1015);
and U36 (N_36,In_493,In_674);
nor U37 (N_37,In_1961,In_988);
and U38 (N_38,In_246,In_1080);
and U39 (N_39,In_1951,In_969);
or U40 (N_40,In_1364,In_408);
or U41 (N_41,In_1128,In_793);
and U42 (N_42,In_123,In_500);
nor U43 (N_43,In_1206,In_1465);
nand U44 (N_44,In_43,In_950);
xnor U45 (N_45,In_1522,In_605);
and U46 (N_46,In_1883,In_1733);
nand U47 (N_47,In_697,In_1985);
or U48 (N_48,In_1814,In_816);
xor U49 (N_49,In_941,In_456);
or U50 (N_50,In_795,In_339);
xor U51 (N_51,In_1371,In_345);
xnor U52 (N_52,In_228,In_358);
or U53 (N_53,In_1991,In_1275);
xnor U54 (N_54,In_555,In_1148);
and U55 (N_55,In_384,In_1469);
nand U56 (N_56,In_1542,In_303);
nand U57 (N_57,In_616,In_333);
nand U58 (N_58,In_457,In_1563);
or U59 (N_59,In_1726,In_1876);
nand U60 (N_60,In_922,In_1486);
or U61 (N_61,In_1824,In_962);
and U62 (N_62,In_1835,In_994);
nor U63 (N_63,In_1313,In_1387);
and U64 (N_64,In_632,In_1457);
nor U65 (N_65,In_1091,In_1719);
and U66 (N_66,In_1749,In_1105);
or U67 (N_67,In_453,In_1945);
nand U68 (N_68,In_1076,In_496);
xor U69 (N_69,In_846,In_1075);
nor U70 (N_70,In_328,In_682);
nand U71 (N_71,In_1644,In_427);
or U72 (N_72,In_1192,In_1758);
nand U73 (N_73,In_1827,In_1636);
nor U74 (N_74,In_1657,In_651);
or U75 (N_75,In_1798,In_680);
and U76 (N_76,In_340,In_817);
or U77 (N_77,In_1927,In_1884);
xor U78 (N_78,In_806,In_400);
xor U79 (N_79,In_971,In_69);
nand U80 (N_80,In_1841,In_1308);
and U81 (N_81,In_624,In_1548);
or U82 (N_82,In_1284,In_701);
or U83 (N_83,In_1515,In_1670);
and U84 (N_84,In_774,In_1202);
nand U85 (N_85,In_1047,In_1230);
xor U86 (N_86,In_1068,In_1740);
and U87 (N_87,In_285,In_675);
xor U88 (N_88,In_413,In_196);
nor U89 (N_89,In_1132,In_645);
and U90 (N_90,In_1152,In_1539);
nor U91 (N_91,In_756,In_1029);
or U92 (N_92,In_1595,In_1394);
nand U93 (N_93,In_582,In_1750);
and U94 (N_94,In_1435,In_242);
or U95 (N_95,In_1721,In_1169);
and U96 (N_96,In_1516,In_1107);
nor U97 (N_97,In_1845,In_1874);
and U98 (N_98,In_1240,In_1348);
and U99 (N_99,In_1543,In_149);
and U100 (N_100,In_1786,In_186);
xnor U101 (N_101,In_1931,In_522);
and U102 (N_102,In_294,In_615);
xnor U103 (N_103,In_1564,In_973);
nor U104 (N_104,In_1474,In_1906);
and U105 (N_105,In_1559,In_563);
and U106 (N_106,In_78,In_827);
or U107 (N_107,In_512,In_1188);
and U108 (N_108,In_407,In_946);
or U109 (N_109,In_1049,In_1307);
nor U110 (N_110,In_370,In_450);
nand U111 (N_111,In_526,In_306);
nand U112 (N_112,In_515,In_403);
nand U113 (N_113,In_1911,In_1079);
xnor U114 (N_114,In_1287,In_1584);
or U115 (N_115,In_872,In_1720);
and U116 (N_116,In_1825,In_552);
nor U117 (N_117,In_1801,In_1403);
nand U118 (N_118,In_1158,In_1155);
nor U119 (N_119,In_1939,In_1446);
nand U120 (N_120,In_1671,In_780);
xor U121 (N_121,In_897,In_255);
nor U122 (N_122,In_1229,In_1770);
nand U123 (N_123,In_622,In_1585);
xnor U124 (N_124,In_1051,In_1291);
nand U125 (N_125,In_264,In_934);
xor U126 (N_126,In_134,In_1019);
and U127 (N_127,In_160,In_1532);
nand U128 (N_128,In_1265,In_1214);
and U129 (N_129,In_1631,In_1470);
nand U130 (N_130,In_1889,In_1299);
or U131 (N_131,In_614,In_391);
nor U132 (N_132,In_179,In_1182);
and U133 (N_133,In_1088,In_1743);
xnor U134 (N_134,In_699,In_1060);
or U135 (N_135,In_829,In_1070);
nand U136 (N_136,In_38,In_47);
or U137 (N_137,In_942,In_1185);
nor U138 (N_138,In_42,In_250);
nor U139 (N_139,In_1099,In_1894);
and U140 (N_140,In_329,In_1968);
xnor U141 (N_141,In_1596,In_1030);
or U142 (N_142,In_845,In_1958);
nand U143 (N_143,In_418,In_1504);
nor U144 (N_144,In_227,In_711);
nor U145 (N_145,In_529,In_297);
nor U146 (N_146,In_83,In_16);
or U147 (N_147,In_1916,In_1635);
or U148 (N_148,In_910,In_1377);
nor U149 (N_149,In_320,In_1498);
and U150 (N_150,In_851,In_1565);
nand U151 (N_151,In_1157,In_1812);
nor U152 (N_152,In_1309,In_1691);
nand U153 (N_153,In_125,In_1331);
or U154 (N_154,In_1816,In_380);
or U155 (N_155,In_499,In_1557);
xnor U156 (N_156,In_1039,In_750);
nor U157 (N_157,In_1154,In_1312);
xnor U158 (N_158,In_696,In_1552);
or U159 (N_159,In_1850,In_1447);
xor U160 (N_160,In_44,In_639);
or U161 (N_161,In_234,In_1036);
or U162 (N_162,In_1804,In_1575);
or U163 (N_163,In_1043,In_1150);
or U164 (N_164,In_1395,In_871);
and U165 (N_165,In_488,In_1767);
nor U166 (N_166,In_1459,In_1855);
xnor U167 (N_167,In_68,In_1059);
xnor U168 (N_168,In_1612,In_1702);
xor U169 (N_169,In_189,In_1247);
nand U170 (N_170,In_28,In_1163);
or U171 (N_171,In_794,In_1725);
xor U172 (N_172,In_1442,In_254);
xor U173 (N_173,In_379,In_1484);
nor U174 (N_174,In_735,In_1382);
nand U175 (N_175,In_1386,In_1561);
or U176 (N_176,In_1445,In_1005);
or U177 (N_177,In_191,In_693);
nand U178 (N_178,In_80,In_1741);
xor U179 (N_179,In_288,In_550);
nor U180 (N_180,In_1058,In_820);
nand U181 (N_181,In_1257,In_1614);
or U182 (N_182,In_610,In_59);
and U183 (N_183,In_332,In_1045);
nor U184 (N_184,In_318,In_1494);
xnor U185 (N_185,In_1791,In_1956);
or U186 (N_186,In_654,In_1822);
nand U187 (N_187,In_1779,In_347);
nor U188 (N_188,In_75,In_899);
xnor U189 (N_189,In_1926,In_649);
and U190 (N_190,In_482,In_1535);
and U191 (N_191,In_107,In_1863);
or U192 (N_192,In_770,In_568);
nand U193 (N_193,In_1044,In_334);
nand U194 (N_194,In_65,In_1205);
xor U195 (N_195,In_1703,In_801);
and U196 (N_196,In_1938,In_1141);
and U197 (N_197,In_1220,In_1607);
nor U198 (N_198,In_1660,In_1864);
xor U199 (N_199,In_1625,In_1718);
or U200 (N_200,In_103,In_412);
nor U201 (N_201,In_1260,In_1338);
nor U202 (N_202,In_1930,In_1953);
and U203 (N_203,In_601,In_337);
or U204 (N_204,In_353,In_1859);
nor U205 (N_205,In_1352,In_1739);
and U206 (N_206,In_787,In_842);
nand U207 (N_207,In_302,In_856);
xor U208 (N_208,In_1149,In_1111);
nor U209 (N_209,In_1806,In_575);
xnor U210 (N_210,In_789,In_1393);
xnor U211 (N_211,In_772,In_71);
nor U212 (N_212,In_82,In_383);
and U213 (N_213,In_1024,In_175);
and U214 (N_214,In_225,In_1512);
xor U215 (N_215,In_583,In_63);
or U216 (N_216,In_1745,In_773);
nand U217 (N_217,In_197,In_507);
nor U218 (N_218,In_73,In_1977);
xnor U219 (N_219,In_1534,In_344);
xor U220 (N_220,In_1175,In_19);
or U221 (N_221,In_238,In_335);
nand U222 (N_222,In_114,In_956);
and U223 (N_223,In_866,In_671);
or U224 (N_224,In_1342,In_627);
nor U225 (N_225,In_1347,In_1238);
nand U226 (N_226,In_517,In_1658);
and U227 (N_227,In_1667,In_1065);
nand U228 (N_228,In_1608,In_677);
or U229 (N_229,In_126,In_717);
xnor U230 (N_230,In_1082,In_1983);
or U231 (N_231,In_1847,In_1586);
or U232 (N_232,In_1392,In_1279);
and U233 (N_233,In_1711,In_1137);
nand U234 (N_234,In_1156,In_448);
and U235 (N_235,In_1634,In_287);
and U236 (N_236,In_415,In_1676);
nand U237 (N_237,In_1682,In_1544);
and U238 (N_238,In_662,In_769);
nor U239 (N_239,In_768,In_535);
and U240 (N_240,In_1763,In_980);
xor U241 (N_241,In_13,In_592);
nand U242 (N_242,In_1651,In_261);
or U243 (N_243,In_991,In_1695);
nor U244 (N_244,In_1904,In_1463);
nor U245 (N_245,In_147,In_1159);
xnor U246 (N_246,In_1483,In_84);
nor U247 (N_247,In_704,In_15);
nor U248 (N_248,In_1656,In_1124);
or U249 (N_249,In_1744,In_1416);
and U250 (N_250,In_74,In_948);
xnor U251 (N_251,In_1692,In_1674);
and U252 (N_252,N_247,In_954);
xnor U253 (N_253,In_326,In_1549);
nor U254 (N_254,N_31,In_1450);
and U255 (N_255,In_105,In_1687);
or U256 (N_256,In_31,In_986);
or U257 (N_257,In_1574,In_904);
or U258 (N_258,In_1672,In_465);
or U259 (N_259,In_935,In_1980);
xor U260 (N_260,N_175,In_814);
and U261 (N_261,N_164,In_623);
nor U262 (N_262,In_1458,In_887);
nor U263 (N_263,In_7,In_1599);
or U264 (N_264,In_1139,In_1705);
or U265 (N_265,In_1629,In_163);
nor U266 (N_266,In_1908,In_1213);
xor U267 (N_267,In_1198,In_667);
and U268 (N_268,In_1899,In_1857);
nor U269 (N_269,In_542,In_1973);
or U270 (N_270,In_1121,In_1094);
and U271 (N_271,In_1208,In_859);
or U272 (N_272,In_1950,In_193);
or U273 (N_273,In_1237,In_1325);
nand U274 (N_274,In_1451,N_243);
xor U275 (N_275,In_1560,In_1852);
nand U276 (N_276,In_815,In_1322);
xnor U277 (N_277,In_1924,In_1795);
or U278 (N_278,In_1683,In_823);
and U279 (N_279,N_165,In_263);
nor U280 (N_280,In_1003,N_86);
xor U281 (N_281,In_1096,In_1501);
or U282 (N_282,N_136,In_1861);
nand U283 (N_283,In_1997,In_1730);
xor U284 (N_284,In_1410,In_420);
nand U285 (N_285,In_112,In_1174);
nand U286 (N_286,In_755,In_22);
xnor U287 (N_287,In_1306,In_736);
nand U288 (N_288,In_611,In_1722);
xnor U289 (N_289,In_1880,In_362);
and U290 (N_290,N_93,In_873);
and U291 (N_291,In_1083,In_1071);
and U292 (N_292,In_678,In_1109);
nand U293 (N_293,In_325,In_685);
nor U294 (N_294,In_30,In_1756);
and U295 (N_295,N_30,In_514);
xnor U296 (N_296,In_673,In_260);
nand U297 (N_297,In_470,In_663);
nand U298 (N_298,In_77,In_321);
and U299 (N_299,In_1955,In_541);
or U300 (N_300,In_476,N_215);
nor U301 (N_301,In_67,In_235);
nand U302 (N_302,In_599,In_1545);
nor U303 (N_303,In_9,N_44);
nor U304 (N_304,In_804,In_118);
and U305 (N_305,In_1989,In_687);
and U306 (N_306,In_1429,In_1505);
or U307 (N_307,In_399,In_1747);
nor U308 (N_308,In_174,In_848);
and U309 (N_309,In_664,In_1464);
xor U310 (N_310,In_1936,In_1396);
xor U311 (N_311,In_276,In_220);
xor U312 (N_312,In_1204,In_908);
xor U313 (N_313,In_889,In_1992);
xor U314 (N_314,In_822,In_970);
and U315 (N_315,In_58,In_12);
nor U316 (N_316,N_59,In_190);
nand U317 (N_317,In_377,In_503);
and U318 (N_318,In_274,In_1748);
or U319 (N_319,In_1456,In_1339);
or U320 (N_320,N_99,In_713);
xor U321 (N_321,In_1487,In_1568);
nor U322 (N_322,In_1689,In_39);
nand U323 (N_323,In_1489,In_1957);
nand U324 (N_324,In_1627,N_147);
xnor U325 (N_325,In_743,In_1685);
nor U326 (N_326,N_148,In_292);
or U327 (N_327,In_715,In_449);
or U328 (N_328,In_34,In_1701);
nand U329 (N_329,N_87,In_586);
xnor U330 (N_330,In_113,In_98);
nand U331 (N_331,In_524,In_1332);
nor U332 (N_332,In_1996,In_1146);
nor U333 (N_333,In_1578,In_1499);
and U334 (N_334,In_1805,In_886);
nand U335 (N_335,In_959,In_828);
or U336 (N_336,N_102,In_319);
and U337 (N_337,N_183,N_76);
xnor U338 (N_338,In_1675,In_387);
nor U339 (N_339,N_0,In_424);
nand U340 (N_340,In_1353,N_24);
xor U341 (N_341,In_372,In_1784);
nand U342 (N_342,In_949,In_1621);
nor U343 (N_343,In_1375,In_911);
and U344 (N_344,In_902,N_227);
and U345 (N_345,In_1093,In_588);
or U346 (N_346,In_1421,In_311);
nor U347 (N_347,In_4,In_625);
xor U348 (N_348,In_843,In_504);
or U349 (N_349,In_111,In_974);
nor U350 (N_350,In_1318,In_1363);
and U351 (N_351,In_1009,In_1688);
xnor U352 (N_352,In_1367,N_25);
or U353 (N_353,In_1272,In_748);
or U354 (N_354,In_1616,N_39);
and U355 (N_355,In_741,In_527);
or U356 (N_356,In_1592,In_209);
and U357 (N_357,In_930,In_240);
and U358 (N_358,N_154,In_336);
and U359 (N_359,N_149,In_436);
nor U360 (N_360,In_1063,In_1830);
xnor U361 (N_361,In_438,In_211);
and U362 (N_362,In_1488,In_1729);
nand U363 (N_363,In_700,In_1343);
nand U364 (N_364,In_1987,In_943);
nand U365 (N_365,In_612,In_1310);
or U366 (N_366,N_172,In_1751);
xnor U367 (N_367,In_630,In_1929);
nand U368 (N_368,In_477,In_1737);
nand U369 (N_369,In_577,In_441);
or U370 (N_370,In_6,In_1314);
nor U371 (N_371,In_145,N_54);
or U372 (N_372,N_235,In_587);
nand U373 (N_373,N_103,In_53);
xor U374 (N_374,In_1400,In_1604);
nor U375 (N_375,In_433,In_96);
xor U376 (N_376,In_167,In_1875);
and U377 (N_377,In_1226,In_1972);
or U378 (N_378,In_757,N_64);
or U379 (N_379,In_1370,In_1085);
nor U380 (N_380,In_879,In_17);
nor U381 (N_381,In_1654,In_1680);
xor U382 (N_382,In_1255,In_790);
nand U383 (N_383,In_1273,In_634);
nand U384 (N_384,N_221,In_422);
or U385 (N_385,N_151,In_1405);
nor U386 (N_386,In_689,N_111);
xor U387 (N_387,In_746,In_478);
nor U388 (N_388,N_153,In_1161);
and U389 (N_389,In_1669,N_191);
nand U390 (N_390,In_782,In_1301);
xor U391 (N_391,In_1362,In_1624);
xor U392 (N_392,In_1282,In_643);
nand U393 (N_393,In_1965,In_1335);
or U394 (N_394,In_861,In_1969);
xnor U395 (N_395,In_1975,In_840);
nand U396 (N_396,In_660,In_692);
nor U397 (N_397,In_1773,In_1011);
xnor U398 (N_398,N_155,In_864);
nand U399 (N_399,In_1304,In_1949);
or U400 (N_400,In_27,In_359);
or U401 (N_401,In_1383,In_1022);
nor U402 (N_402,In_309,In_501);
or U403 (N_403,In_1603,In_1577);
xnor U404 (N_404,In_25,In_1274);
nor U405 (N_405,N_237,In_944);
nand U406 (N_406,In_640,N_114);
xnor U407 (N_407,In_185,In_885);
or U408 (N_408,In_198,In_1006);
nor U409 (N_409,In_375,In_1374);
nand U410 (N_410,In_278,In_1018);
xnor U411 (N_411,In_1594,In_1241);
nor U412 (N_412,In_602,In_745);
nand U413 (N_413,In_1960,N_28);
and U414 (N_414,In_249,In_1811);
or U415 (N_415,In_1119,N_184);
and U416 (N_416,In_283,In_91);
xnor U417 (N_417,In_351,In_1320);
nand U418 (N_418,In_1253,In_936);
or U419 (N_419,In_61,In_1854);
or U420 (N_420,In_923,In_62);
or U421 (N_421,In_1935,In_1248);
nand U422 (N_422,In_49,N_159);
or U423 (N_423,In_1184,In_637);
xor U424 (N_424,In_1140,N_206);
xnor U425 (N_425,In_1340,In_925);
or U426 (N_426,N_238,In_1506);
xnor U427 (N_427,In_352,In_1513);
nor U428 (N_428,In_1984,In_1976);
and U429 (N_429,In_135,N_66);
or U430 (N_430,N_134,In_401);
or U431 (N_431,In_1978,N_48);
and U432 (N_432,N_135,In_1652);
nand U433 (N_433,In_661,In_870);
and U434 (N_434,In_1877,In_502);
nand U435 (N_435,In_1252,In_1330);
nor U436 (N_436,In_81,In_268);
and U437 (N_437,In_1920,In_1598);
nor U438 (N_438,In_683,In_1839);
nor U439 (N_439,In_533,In_1341);
or U440 (N_440,In_218,In_1519);
nand U441 (N_441,In_1160,In_1315);
or U442 (N_442,In_1872,In_1700);
nand U443 (N_443,In_1650,In_753);
or U444 (N_444,In_877,N_4);
and U445 (N_445,In_1048,In_1138);
nand U446 (N_446,In_1345,N_18);
nand U447 (N_447,In_1946,N_200);
nor U448 (N_448,In_374,In_397);
or U449 (N_449,In_388,In_839);
and U450 (N_450,N_158,In_1251);
nor U451 (N_451,In_1642,In_1990);
or U452 (N_452,In_618,In_1518);
xnor U453 (N_453,In_819,In_253);
xor U454 (N_454,In_1659,N_63);
nand U455 (N_455,In_1643,In_161);
nand U456 (N_456,In_1712,In_1476);
nor U457 (N_457,N_189,In_32);
xor U458 (N_458,In_1106,N_116);
nor U459 (N_459,In_440,In_300);
nand U460 (N_460,In_1485,N_17);
and U461 (N_461,In_199,In_1982);
and U462 (N_462,In_655,N_186);
and U463 (N_463,In_730,In_734);
xor U464 (N_464,In_1525,In_955);
nand U465 (N_465,In_1605,In_1095);
or U466 (N_466,In_591,In_1433);
nor U467 (N_467,In_392,In_1471);
and U468 (N_468,In_1694,In_993);
xor U469 (N_469,In_992,In_694);
xor U470 (N_470,N_97,In_1280);
xor U471 (N_471,In_1098,In_508);
xor U472 (N_472,N_78,In_177);
nor U473 (N_473,In_695,In_1115);
or U474 (N_474,In_324,N_29);
xor U475 (N_475,In_1041,N_140);
or U476 (N_476,In_1849,In_841);
nor U477 (N_477,In_571,In_545);
nor U478 (N_478,In_1832,In_445);
nand U479 (N_479,In_1389,In_932);
nor U480 (N_480,In_271,In_272);
xnor U481 (N_481,In_710,In_256);
and U482 (N_482,In_1886,N_138);
nor U483 (N_483,In_895,In_301);
nor U484 (N_484,In_984,N_146);
and U485 (N_485,In_231,In_811);
or U486 (N_486,In_852,In_1843);
and U487 (N_487,In_1189,In_1244);
nor U488 (N_488,In_999,In_295);
nand U489 (N_489,In_119,In_489);
xor U490 (N_490,N_10,In_1122);
nor U491 (N_491,N_190,In_759);
nor U492 (N_492,In_14,In_888);
nand U493 (N_493,In_367,In_556);
or U494 (N_494,In_1838,In_589);
or U495 (N_495,In_1922,N_161);
and U496 (N_496,In_1057,In_1061);
nand U497 (N_497,In_1461,In_1072);
or U498 (N_498,In_884,In_443);
nand U499 (N_499,In_1046,In_195);
xnor U500 (N_500,In_724,In_483);
nor U501 (N_501,In_1466,In_964);
xnor U502 (N_502,In_1449,In_99);
nand U503 (N_503,In_1042,In_1191);
xor U504 (N_504,In_224,In_1359);
and U505 (N_505,In_1896,In_1553);
xnor U506 (N_506,N_295,In_159);
or U507 (N_507,In_1180,In_1893);
and U508 (N_508,In_269,In_681);
nor U509 (N_509,In_593,In_381);
nand U510 (N_510,In_76,N_360);
or U511 (N_511,In_1263,N_358);
nand U512 (N_512,In_521,In_459);
or U513 (N_513,In_1790,In_120);
nand U514 (N_514,In_1414,N_456);
nand U515 (N_515,In_1792,N_342);
or U516 (N_516,In_117,In_1);
and U517 (N_517,In_987,In_1707);
or U518 (N_518,In_1836,In_1090);
and U519 (N_519,In_1165,In_1087);
or U520 (N_520,In_1089,N_115);
nand U521 (N_521,In_672,N_364);
nand U522 (N_522,N_198,N_196);
or U523 (N_523,In_469,In_308);
and U524 (N_524,In_1587,In_188);
or U525 (N_525,In_389,In_1034);
nand U526 (N_526,In_909,N_11);
or U527 (N_527,In_905,In_1097);
nor U528 (N_528,In_1497,N_488);
nor U529 (N_529,In_1554,In_1007);
and U530 (N_530,In_989,In_473);
or U531 (N_531,In_812,In_1329);
nor U532 (N_532,In_951,N_413);
or U533 (N_533,In_1928,In_797);
and U534 (N_534,N_344,N_317);
and U535 (N_535,In_1153,N_65);
and U536 (N_536,In_280,In_990);
and U537 (N_537,In_511,In_1591);
nand U538 (N_538,In_291,In_608);
xor U539 (N_539,In_920,N_305);
xnor U540 (N_540,In_1910,In_1626);
and U541 (N_541,In_1028,In_1221);
or U542 (N_542,In_64,N_323);
nand U543 (N_543,N_2,N_83);
and U544 (N_544,In_1215,N_19);
nand U545 (N_545,In_559,In_1135);
and U546 (N_546,In_3,In_629);
or U547 (N_547,In_860,N_280);
nand U548 (N_548,N_219,In_594);
nor U549 (N_549,In_435,In_1696);
or U550 (N_550,In_1283,In_1999);
nor U551 (N_551,In_1116,In_576);
nor U552 (N_552,In_183,In_1681);
and U553 (N_553,In_1509,N_417);
nor U554 (N_554,N_322,In_721);
nand U555 (N_555,In_151,N_6);
xor U556 (N_556,N_455,N_384);
and U557 (N_557,N_476,In_1887);
nand U558 (N_558,In_1550,In_1527);
nand U559 (N_559,In_1909,In_378);
or U560 (N_560,N_27,In_419);
or U561 (N_561,N_419,In_201);
xor U562 (N_562,In_1900,In_172);
and U563 (N_563,In_914,N_491);
nand U564 (N_564,In_1537,N_130);
nor U565 (N_565,In_314,N_283);
xor U566 (N_566,In_751,N_311);
or U567 (N_567,N_171,N_347);
and U568 (N_568,In_1819,N_210);
or U569 (N_569,In_547,In_208);
nand U570 (N_570,In_259,In_1436);
nand U571 (N_571,In_1129,In_182);
nor U572 (N_572,In_918,In_1354);
or U573 (N_573,N_192,In_1601);
or U574 (N_574,In_1738,In_1355);
and U575 (N_575,N_447,In_1647);
or U576 (N_576,In_252,In_152);
nand U577 (N_577,In_1597,N_410);
and U578 (N_578,N_363,N_156);
nand U579 (N_579,In_1579,In_233);
nand U580 (N_580,In_896,N_205);
nor U581 (N_581,N_366,In_24);
or U582 (N_582,In_1789,In_883);
nand U583 (N_583,N_234,N_20);
nand U584 (N_584,N_381,In_1197);
or U585 (N_585,N_352,In_1223);
xor U586 (N_586,In_1462,In_569);
xnor U587 (N_587,N_35,In_1211);
nand U588 (N_588,In_1050,In_1556);
nand U589 (N_589,In_638,In_853);
nand U590 (N_590,In_41,In_1546);
and U591 (N_591,In_1453,In_1580);
or U592 (N_592,N_106,In_286);
and U593 (N_593,In_1236,In_1717);
nand U594 (N_594,N_337,In_985);
or U595 (N_595,In_1468,N_353);
and U596 (N_596,N_179,In_355);
xor U597 (N_597,In_1514,In_1934);
nor U598 (N_598,In_1427,N_427);
nand U599 (N_599,In_442,In_505);
or U600 (N_600,In_26,N_374);
nor U601 (N_601,In_657,In_1170);
nor U602 (N_602,N_137,In_1757);
nor U603 (N_603,In_1858,In_1821);
or U604 (N_604,In_540,N_408);
or U605 (N_605,In_516,In_509);
nor U606 (N_606,In_110,In_1856);
nand U607 (N_607,In_1133,In_1130);
nand U608 (N_608,N_497,In_467);
nor U609 (N_609,N_436,N_367);
and U610 (N_610,In_491,In_382);
nand U611 (N_611,N_176,In_684);
xor U612 (N_612,N_383,N_89);
nand U613 (N_613,In_666,In_560);
and U614 (N_614,In_366,In_1962);
or U615 (N_615,N_433,In_425);
or U616 (N_616,In_1551,In_1008);
nand U617 (N_617,In_1617,N_94);
nor U618 (N_618,In_1302,N_401);
or U619 (N_619,N_23,N_465);
xnor U620 (N_620,In_451,N_259);
or U621 (N_621,N_22,In_1472);
nor U622 (N_622,In_1787,In_708);
or U623 (N_623,In_1117,In_1479);
nor U624 (N_624,N_12,In_1423);
nor U625 (N_625,N_438,N_228);
or U626 (N_626,In_1365,In_212);
nor U627 (N_627,In_1001,N_152);
nand U628 (N_628,In_88,In_1529);
nand U629 (N_629,In_239,In_1803);
xnor U630 (N_630,N_45,N_157);
and U631 (N_631,In_124,In_1134);
nor U632 (N_632,In_628,In_937);
nor U633 (N_633,N_480,N_294);
or U634 (N_634,In_277,In_1502);
nor U635 (N_635,In_1528,In_620);
or U636 (N_636,In_1912,N_224);
nand U637 (N_637,In_466,In_1709);
and U638 (N_638,In_764,In_368);
or U639 (N_639,In_1190,In_799);
xor U640 (N_640,N_104,In_847);
or U641 (N_641,In_850,N_392);
nor U642 (N_642,In_1074,In_1919);
xnor U643 (N_643,In_1714,N_9);
or U644 (N_644,In_631,In_169);
or U645 (N_645,N_166,N_333);
xor U646 (N_646,In_180,In_1679);
and U647 (N_647,N_426,N_463);
and U648 (N_648,In_762,In_1885);
and U649 (N_649,In_916,N_499);
or U650 (N_650,N_181,In_143);
nor U651 (N_651,N_270,In_480);
nor U652 (N_652,In_1571,In_141);
and U653 (N_653,N_478,N_483);
and U654 (N_654,In_1573,In_1524);
nand U655 (N_655,In_1998,In_157);
or U656 (N_656,N_245,In_644);
and U657 (N_657,In_155,In_162);
and U658 (N_658,In_1844,In_1200);
nor U659 (N_659,N_217,In_1337);
and U660 (N_660,N_34,In_214);
nand U661 (N_661,N_334,In_1897);
xor U662 (N_662,In_1123,In_1357);
nand U663 (N_663,In_1878,In_472);
nand U664 (N_664,In_226,In_1613);
and U665 (N_665,In_965,In_338);
nand U666 (N_666,In_1710,In_1127);
xnor U667 (N_667,In_1327,In_1862);
nand U668 (N_668,N_355,In_207);
xor U669 (N_669,In_1831,In_1637);
nor U670 (N_670,In_538,In_247);
or U671 (N_671,In_1693,N_356);
nand U672 (N_672,In_173,In_733);
xnor U673 (N_673,In_998,N_428);
and U674 (N_674,N_405,In_349);
xor U675 (N_675,In_498,In_1407);
nand U676 (N_676,N_416,In_1782);
nor U677 (N_677,In_1799,In_1760);
xnor U678 (N_678,In_1570,N_120);
xnor U679 (N_679,N_373,In_1746);
or U680 (N_680,N_430,In_1112);
nand U681 (N_681,N_255,In_1012);
nor U682 (N_682,In_1826,In_633);
and U683 (N_683,N_434,In_1728);
nand U684 (N_684,In_1031,N_16);
nand U685 (N_685,In_363,In_136);
or U686 (N_686,In_1475,In_1834);
or U687 (N_687,In_1523,N_362);
nand U688 (N_688,In_1848,In_1369);
xnor U689 (N_689,In_1428,In_1881);
or U690 (N_690,In_548,In_975);
nor U691 (N_691,In_369,In_1817);
nor U692 (N_692,In_229,In_865);
or U693 (N_693,N_421,In_411);
nor U694 (N_694,In_1940,N_460);
nand U695 (N_695,In_963,In_284);
or U696 (N_696,In_181,In_245);
or U697 (N_697,N_268,N_254);
and U698 (N_698,In_854,In_1431);
or U699 (N_699,In_1905,In_1944);
xnor U700 (N_700,In_405,In_137);
nand U701 (N_701,In_581,In_1269);
xnor U702 (N_702,In_881,N_359);
or U703 (N_703,N_298,In_1256);
nor U704 (N_704,In_1698,In_1943);
and U705 (N_705,In_1732,N_60);
and U706 (N_706,In_808,In_1533);
and U707 (N_707,In_926,In_1418);
nand U708 (N_708,N_267,N_418);
and U709 (N_709,In_564,In_251);
and U710 (N_710,N_301,N_251);
nand U711 (N_711,In_656,In_802);
nor U712 (N_712,In_1979,In_1611);
or U713 (N_713,In_298,In_553);
nand U714 (N_714,N_414,N_396);
or U715 (N_715,N_119,In_104);
or U716 (N_716,In_1196,In_1289);
xnor U717 (N_717,N_105,In_164);
xnor U718 (N_718,In_858,In_1439);
nor U719 (N_719,In_573,N_38);
and U720 (N_720,In_532,In_596);
nor U721 (N_721,In_1677,In_37);
or U722 (N_722,N_395,In_744);
or U723 (N_723,N_123,In_938);
and U724 (N_724,In_892,N_372);
and U725 (N_725,In_813,In_1723);
or U726 (N_726,In_1178,In_1290);
nand U727 (N_727,In_1020,In_421);
nor U728 (N_728,In_1495,In_1923);
and U729 (N_729,In_838,In_712);
nand U730 (N_730,N_212,In_1981);
and U731 (N_731,In_788,N_448);
or U732 (N_732,N_475,In_849);
and U733 (N_733,In_723,N_246);
nor U734 (N_734,In_1797,N_302);
nand U735 (N_735,In_953,In_868);
nor U736 (N_736,In_1002,N_47);
xnor U737 (N_737,In_995,In_184);
nor U738 (N_738,In_51,In_1628);
nor U739 (N_739,In_1227,In_1303);
or U740 (N_740,In_215,In_2);
xnor U741 (N_741,N_377,In_146);
or U742 (N_742,In_1413,N_128);
or U743 (N_743,N_209,N_141);
or U744 (N_744,N_269,In_1947);
or U745 (N_745,In_1913,In_807);
nand U746 (N_746,N_51,In_921);
or U747 (N_747,In_1915,In_1066);
and U748 (N_748,In_1641,In_423);
xor U749 (N_749,In_1638,In_1496);
and U750 (N_750,In_1520,In_726);
nand U751 (N_751,In_1823,In_1016);
xor U752 (N_752,In_1267,In_635);
and U753 (N_753,N_265,In_1530);
nor U754 (N_754,N_735,In_237);
nor U755 (N_755,In_1646,In_1668);
or U756 (N_756,In_313,In_1507);
or U757 (N_757,In_603,In_1995);
or U758 (N_758,In_1067,In_1110);
nand U759 (N_759,N_299,N_113);
or U760 (N_760,N_486,In_621);
xor U761 (N_761,In_1235,N_614);
nor U762 (N_762,N_677,In_1113);
nand U763 (N_763,N_725,In_93);
nor U764 (N_764,N_453,N_709);
xor U765 (N_765,N_324,N_230);
or U766 (N_766,In_18,In_132);
nand U767 (N_767,N_284,N_69);
nand U768 (N_768,In_1056,N_522);
nor U769 (N_769,In_394,N_738);
nand U770 (N_770,In_544,N_167);
nor U771 (N_771,In_967,N_535);
nor U772 (N_772,In_327,In_1125);
nand U773 (N_773,N_634,In_468);
nor U774 (N_774,In_171,In_1406);
xor U775 (N_775,N_110,In_244);
and U776 (N_776,N_107,In_447);
nor U777 (N_777,In_1434,In_1014);
nand U778 (N_778,N_708,N_722);
xnor U779 (N_779,In_1813,In_1891);
or U780 (N_780,N_695,In_1233);
xor U781 (N_781,In_1540,N_699);
nand U782 (N_782,In_1216,In_659);
xnor U783 (N_783,In_1785,In_1460);
nand U784 (N_784,In_1500,In_1261);
xnor U785 (N_785,In_129,N_278);
nand U786 (N_786,In_1209,In_641);
or U787 (N_787,In_1164,N_117);
or U788 (N_788,In_1917,N_489);
nand U789 (N_789,In_376,N_526);
and U790 (N_790,In_893,In_1194);
nand U791 (N_791,N_57,N_513);
nand U792 (N_792,In_54,N_551);
and U793 (N_793,N_266,In_952);
or U794 (N_794,In_924,In_1420);
and U795 (N_795,In_1086,In_1907);
xor U796 (N_796,N_681,N_679);
nand U797 (N_797,In_1481,N_654);
xnor U798 (N_798,N_611,N_244);
xor U799 (N_799,N_437,In_305);
or U800 (N_800,In_79,In_1366);
nor U801 (N_801,In_1292,N_638);
xor U802 (N_802,N_472,In_1555);
xnor U803 (N_803,In_33,In_217);
or U804 (N_804,In_1033,N_399);
nor U805 (N_805,In_1490,In_1199);
xor U806 (N_806,N_380,In_1772);
xnor U807 (N_807,In_1716,In_1145);
and U808 (N_808,N_316,In_1424);
nand U809 (N_809,In_296,N_331);
nand U810 (N_810,N_37,N_394);
xor U811 (N_811,N_55,In_1004);
and U812 (N_812,N_739,In_531);
nand U813 (N_813,N_203,In_1941);
and U814 (N_814,N_50,In_765);
xor U815 (N_815,In_1228,N_604);
nand U816 (N_816,In_139,N_688);
or U817 (N_817,In_133,In_679);
nor U818 (N_818,In_1870,In_606);
and U819 (N_819,N_400,In_1828);
and U820 (N_820,In_1173,N_602);
xnor U821 (N_821,N_36,In_519);
or U822 (N_822,N_572,N_712);
and U823 (N_823,In_1177,In_836);
and U824 (N_824,In_1538,In_1866);
nor U825 (N_825,N_188,N_81);
nor U826 (N_826,In_1100,N_271);
nand U827 (N_827,N_53,In_1136);
and U828 (N_828,In_929,In_356);
nand U829 (N_829,In_1399,N_664);
nor U830 (N_830,N_108,N_452);
or U831 (N_831,In_1092,In_342);
xnor U832 (N_832,In_719,N_594);
nor U833 (N_833,N_222,N_7);
nor U834 (N_834,N_613,In_907);
and U835 (N_835,In_1771,In_561);
or U836 (N_836,N_257,In_1622);
or U837 (N_837,N_61,In_1753);
xnor U838 (N_838,In_289,In_1017);
and U839 (N_839,In_130,In_1262);
xnor U840 (N_840,In_1810,In_776);
xor U841 (N_841,In_1794,In_127);
or U842 (N_842,In_452,N_687);
xnor U843 (N_843,In_350,N_112);
or U844 (N_844,In_1073,N_308);
or U845 (N_845,N_420,In_786);
and U846 (N_846,N_482,In_1665);
xor U847 (N_847,In_1754,N_474);
and U848 (N_848,In_1618,N_720);
xnor U849 (N_849,In_739,In_791);
xor U850 (N_850,N_501,N_213);
nand U851 (N_851,In_148,In_1918);
and U852 (N_852,In_1183,In_1879);
nand U853 (N_853,In_1473,N_689);
or U854 (N_854,In_1686,N_320);
xor U855 (N_855,N_624,N_511);
or U856 (N_856,N_208,In_1224);
or U857 (N_857,In_901,In_617);
xor U858 (N_858,N_429,In_1246);
and U859 (N_859,In_1890,N_82);
xnor U860 (N_860,In_1027,In_1402);
nand U861 (N_861,N_548,N_693);
or U862 (N_862,In_1025,N_619);
and U863 (N_863,N_502,In_410);
and U864 (N_864,In_70,In_598);
or U865 (N_865,In_894,N_332);
nand U866 (N_866,N_540,N_541);
nor U867 (N_867,In_716,In_1151);
nor U868 (N_868,In_518,In_210);
nand U869 (N_869,N_631,In_1077);
nand U870 (N_870,In_690,In_1114);
nand U871 (N_871,In_1035,N_740);
and U872 (N_872,In_439,N_14);
and U873 (N_873,N_543,In_523);
nor U874 (N_874,N_583,In_1281);
nor U875 (N_875,N_562,In_1373);
nand U876 (N_876,N_327,In_878);
nand U877 (N_877,N_258,In_1356);
nor U878 (N_878,In_1181,In_1231);
nand U879 (N_879,N_615,In_698);
xor U880 (N_880,N_517,N_635);
nand U881 (N_881,In_471,N_558);
or U882 (N_882,In_1187,N_576);
or U883 (N_883,N_143,In_558);
nor U884 (N_884,In_1868,In_417);
or U885 (N_885,In_1425,In_702);
nand U886 (N_886,In_1103,N_536);
and U887 (N_887,N_361,N_43);
xor U888 (N_888,In_1305,N_249);
xor U889 (N_889,N_412,N_385);
nor U890 (N_890,In_1172,N_461);
or U891 (N_891,N_325,In_1013);
nor U892 (N_892,N_729,N_195);
xnor U893 (N_893,In_72,N_239);
nor U894 (N_894,In_409,In_867);
nand U895 (N_895,In_983,N_591);
and U896 (N_896,In_266,In_1404);
or U897 (N_897,N_62,In_1818);
and U898 (N_898,N_406,N_534);
nor U899 (N_899,N_744,In_1632);
xor U900 (N_900,In_46,In_595);
or U901 (N_901,N_346,N_577);
or U902 (N_902,In_1254,In_279);
xnor U903 (N_903,N_500,N_330);
nor U904 (N_904,In_1480,N_132);
xnor U905 (N_905,N_126,N_552);
and U906 (N_906,N_328,N_561);
xnor U907 (N_907,In_484,In_961);
nor U908 (N_908,N_642,N_369);
and U909 (N_909,In_1678,N_74);
or U910 (N_910,In_580,In_317);
xor U911 (N_911,In_1441,N_630);
and U912 (N_912,N_595,N_160);
or U913 (N_913,In_385,N_545);
nor U914 (N_914,In_1774,In_1653);
nor U915 (N_915,In_1380,In_464);
nor U916 (N_916,N_600,In_917);
nor U917 (N_917,In_1245,N_56);
and U918 (N_918,N_529,N_525);
or U919 (N_919,N_490,N_300);
xor U920 (N_920,In_1583,N_518);
xor U921 (N_921,N_170,N_700);
or U922 (N_922,N_92,In_1316);
nor U923 (N_923,In_1412,N_713);
nor U924 (N_924,In_1298,In_100);
nor U925 (N_925,In_1055,In_1775);
or U926 (N_926,N_569,In_1793);
or U927 (N_927,In_168,In_566);
nor U928 (N_928,N_659,In_1293);
xnor U929 (N_929,In_1388,In_170);
xor U930 (N_930,In_1762,In_1384);
nand U931 (N_931,In_1360,In_543);
nand U932 (N_932,N_556,N_289);
nor U933 (N_933,In_1993,In_1921);
nor U934 (N_934,N_162,In_1319);
nand U935 (N_935,N_88,N_85);
and U936 (N_936,In_243,N_578);
nand U937 (N_937,N_341,In_55);
nor U938 (N_938,In_1895,N_546);
xnor U939 (N_939,N_589,In_236);
xor U940 (N_940,In_539,N_403);
or U941 (N_941,N_567,In_142);
nand U942 (N_942,N_504,N_451);
nand U943 (N_943,In_525,In_1783);
nand U944 (N_944,In_803,N_714);
nand U945 (N_945,In_1666,In_1593);
and U946 (N_946,In_834,N_32);
or U947 (N_947,In_474,N_603);
nor U948 (N_948,In_1225,In_1986);
nand U949 (N_949,N_470,N_13);
or U950 (N_950,N_626,In_402);
nand U951 (N_951,In_430,In_307);
and U952 (N_952,N_686,In_880);
xnor U953 (N_953,N_524,N_49);
xnor U954 (N_954,In_1266,In_1179);
nor U955 (N_955,N_557,In_1788);
and U956 (N_956,N_730,N_388);
and U957 (N_957,In_205,In_1867);
nand U958 (N_958,In_485,In_1328);
or U959 (N_959,In_1898,In_800);
or U960 (N_960,In_805,In_138);
xor U961 (N_961,In_437,In_323);
nand U962 (N_962,N_77,N_487);
xnor U963 (N_963,In_775,In_1398);
or U964 (N_964,In_1052,N_95);
xor U965 (N_965,In_315,In_857);
and U966 (N_966,N_261,In_1432);
xor U967 (N_967,In_94,In_778);
xnor U968 (N_968,In_1295,In_1966);
nor U969 (N_969,In_1336,In_1131);
nand U970 (N_970,N_178,N_272);
nor U971 (N_971,N_683,N_319);
nand U972 (N_972,N_742,In_725);
and U973 (N_973,In_1324,N_690);
or U974 (N_974,N_318,N_454);
or U975 (N_975,N_314,In_1620);
or U976 (N_976,N_606,N_98);
and U977 (N_977,In_1840,N_636);
nor U978 (N_978,N_481,In_578);
xnor U979 (N_979,N_492,N_236);
nand U980 (N_980,In_875,In_1259);
nor U981 (N_981,N_240,N_519);
nor U982 (N_982,In_939,N_671);
nor U983 (N_983,In_783,In_1764);
and U984 (N_984,In_1026,In_1351);
or U985 (N_985,N_70,In_781);
nand U986 (N_986,In_686,N_211);
and U987 (N_987,In_154,In_1358);
nand U988 (N_988,In_1925,N_559);
nand U989 (N_989,In_360,N_663);
xor U990 (N_990,In_1837,In_785);
and U991 (N_991,N_101,In_931);
xnor U992 (N_992,N_647,In_882);
xor U993 (N_993,N_335,In_766);
nand U994 (N_994,N_371,N_579);
xor U995 (N_995,In_265,N_139);
and U996 (N_996,N_637,In_216);
nand U997 (N_997,N_674,In_1808);
xnor U998 (N_998,N_262,N_233);
or U999 (N_999,In_262,N_530);
or U1000 (N_1000,N_274,N_767);
nand U1001 (N_1001,In_933,In_281);
and U1002 (N_1002,N_493,N_131);
or U1003 (N_1003,N_670,N_309);
and U1004 (N_1004,In_346,N_277);
or U1005 (N_1005,N_458,In_1344);
or U1006 (N_1006,In_429,N_962);
xnor U1007 (N_1007,In_1391,N_285);
and U1008 (N_1008,N_632,N_836);
xor U1009 (N_1009,In_809,N_898);
nor U1010 (N_1010,N_568,N_857);
nand U1011 (N_1011,N_521,In_1796);
and U1012 (N_1012,In_832,In_742);
or U1013 (N_1013,N_849,In_1882);
nor U1014 (N_1014,In_604,N_780);
nand U1015 (N_1015,N_554,N_776);
nand U1016 (N_1016,N_697,N_930);
or U1017 (N_1017,In_1376,In_1963);
xor U1018 (N_1018,N_979,In_913);
and U1019 (N_1019,In_348,In_343);
and U1020 (N_1020,N_900,In_97);
nand U1021 (N_1021,In_676,In_691);
xor U1022 (N_1022,N_640,N_644);
or U1023 (N_1023,In_1397,N_218);
or U1024 (N_1024,N_892,N_52);
xnor U1025 (N_1025,In_1201,N_538);
or U1026 (N_1026,N_779,In_1278);
nand U1027 (N_1027,In_557,In_102);
xnor U1028 (N_1028,N_425,N_880);
xor U1029 (N_1029,N_957,N_662);
nand U1030 (N_1030,N_507,N_904);
or U1031 (N_1031,N_390,N_118);
and U1032 (N_1032,N_811,In_178);
nand U1033 (N_1033,N_853,In_927);
or U1034 (N_1034,N_879,N_547);
and U1035 (N_1035,In_1234,N_174);
and U1036 (N_1036,N_891,N_980);
and U1037 (N_1037,N_498,N_875);
and U1038 (N_1038,N_617,N_908);
nand U1039 (N_1039,N_676,In_275);
xor U1040 (N_1040,N_719,N_951);
or U1041 (N_1041,N_940,In_1851);
nor U1042 (N_1042,In_23,In_855);
or U1043 (N_1043,N_984,N_370);
xnor U1044 (N_1044,N_935,In_1250);
nor U1045 (N_1045,In_222,N_555);
and U1046 (N_1046,N_760,N_468);
and U1047 (N_1047,N_340,N_718);
nor U1048 (N_1048,N_863,N_967);
or U1049 (N_1049,N_46,N_682);
or U1050 (N_1050,N_859,In_1104);
nor U1051 (N_1051,N_791,In_996);
xor U1052 (N_1052,In_1633,N_765);
nand U1053 (N_1053,In_1437,N_293);
or U1054 (N_1054,N_827,In_1562);
nand U1055 (N_1055,N_938,In_1478);
nor U1056 (N_1056,N_757,N_303);
xnor U1057 (N_1057,N_643,N_586);
nand U1058 (N_1058,N_623,N_404);
nor U1059 (N_1059,In_982,N_976);
nand U1060 (N_1060,N_607,In_1942);
or U1061 (N_1061,N_599,N_348);
or U1062 (N_1062,N_912,In_416);
nor U1063 (N_1063,N_947,In_1053);
nor U1064 (N_1064,N_816,In_176);
nand U1065 (N_1065,In_835,In_728);
nand U1066 (N_1066,In_299,N_927);
or U1067 (N_1067,N_307,In_732);
nand U1068 (N_1068,N_685,N_641);
nor U1069 (N_1069,N_226,In_979);
nand U1070 (N_1070,N_883,N_834);
nor U1071 (N_1071,N_129,N_838);
nor U1072 (N_1072,N_986,N_723);
nand U1073 (N_1073,N_622,In_1477);
and U1074 (N_1074,N_761,N_874);
xor U1075 (N_1075,In_1232,In_192);
xor U1076 (N_1076,N_970,In_131);
nor U1077 (N_1077,In_647,N_921);
and U1078 (N_1078,In_1761,N_954);
nor U1079 (N_1079,In_373,N_895);
or U1080 (N_1080,In_1959,In_165);
and U1081 (N_1081,N_920,In_506);
nor U1082 (N_1082,In_1492,N_832);
or U1083 (N_1083,In_665,N_894);
xnor U1084 (N_1084,N_509,N_40);
and U1085 (N_1085,In_900,In_221);
nor U1086 (N_1086,N_21,N_485);
nand U1087 (N_1087,In_653,In_1673);
nor U1088 (N_1088,N_902,N_783);
nand U1089 (N_1089,N_193,In_90);
nand U1090 (N_1090,N_570,N_881);
nor U1091 (N_1091,In_5,N_378);
xor U1092 (N_1092,N_746,In_8);
or U1093 (N_1093,In_718,In_727);
nand U1094 (N_1094,In_1964,N_669);
nor U1095 (N_1095,In_891,In_792);
or U1096 (N_1096,N_142,N_411);
nor U1097 (N_1097,In_95,In_158);
xnor U1098 (N_1098,In_109,N_580);
nor U1099 (N_1099,N_527,In_876);
or U1100 (N_1100,In_1526,N_916);
or U1101 (N_1101,In_390,In_1606);
nor U1102 (N_1102,N_133,In_460);
or U1103 (N_1103,N_422,In_1708);
nor U1104 (N_1104,N_873,N_590);
nor U1105 (N_1105,N_826,N_835);
or U1106 (N_1106,N_861,N_84);
nor U1107 (N_1107,In_20,In_747);
and U1108 (N_1108,N_972,In_752);
or U1109 (N_1109,N_173,In_1258);
xnor U1110 (N_1110,N_889,N_550);
nand U1111 (N_1111,N_214,In_646);
xnor U1112 (N_1112,N_924,In_1508);
nor U1113 (N_1113,In_1294,In_767);
nor U1114 (N_1114,N_560,N_982);
or U1115 (N_1115,N_42,In_187);
and U1116 (N_1116,N_726,N_310);
and U1117 (N_1117,N_809,N_665);
nand U1118 (N_1118,In_121,N_242);
and U1119 (N_1119,N_96,N_457);
xnor U1120 (N_1120,In_818,N_657);
and U1121 (N_1121,In_513,N_763);
nand U1122 (N_1122,N_913,N_715);
nor U1123 (N_1123,In_1032,In_714);
or U1124 (N_1124,In_1296,In_1390);
xnor U1125 (N_1125,N_819,In_810);
and U1126 (N_1126,In_1933,In_1218);
or U1127 (N_1127,N_858,N_817);
nand U1128 (N_1128,In_549,In_1276);
and U1129 (N_1129,In_1270,N_821);
nand U1130 (N_1130,N_639,In_1102);
nor U1131 (N_1131,N_948,In_282);
nor U1132 (N_1132,In_1649,N_282);
and U1133 (N_1133,In_1664,In_1503);
or U1134 (N_1134,In_101,N_618);
and U1135 (N_1135,N_185,N_707);
nor U1136 (N_1136,N_953,N_841);
nand U1137 (N_1137,N_252,In_626);
or U1138 (N_1138,N_721,In_10);
or U1139 (N_1139,In_1023,In_258);
nand U1140 (N_1140,In_1602,N_860);
or U1141 (N_1141,N_672,N_71);
nand U1142 (N_1142,N_528,N_985);
nand U1143 (N_1143,In_1143,N_877);
and U1144 (N_1144,N_869,N_592);
xnor U1145 (N_1145,In_636,In_658);
and U1146 (N_1146,N_656,N_609);
nor U1147 (N_1147,In_903,N_515);
nand U1148 (N_1148,In_206,N_393);
and U1149 (N_1149,N_782,In_108);
or U1150 (N_1150,N_290,N_755);
nor U1151 (N_1151,In_1249,In_273);
xor U1152 (N_1152,N_737,N_814);
or U1153 (N_1153,In_777,In_1443);
nand U1154 (N_1154,In_1902,In_1069);
nor U1155 (N_1155,N_804,In_495);
nor U1156 (N_1156,In_1203,N_431);
xnor U1157 (N_1157,N_510,In_1706);
nor U1158 (N_1158,In_1809,In_958);
xnor U1159 (N_1159,In_869,In_1372);
nand U1160 (N_1160,In_48,N_795);
or U1161 (N_1161,In_537,In_1448);
xnor U1162 (N_1162,N_596,N_965);
or U1163 (N_1163,In_1243,In_1610);
nor U1164 (N_1164,In_1144,In_976);
and U1165 (N_1165,N_825,In_331);
or U1166 (N_1166,N_402,In_1171);
and U1167 (N_1167,In_530,In_833);
or U1168 (N_1168,In_50,In_106);
xor U1169 (N_1169,N_313,N_950);
nand U1170 (N_1170,In_1776,N_585);
nand U1171 (N_1171,N_802,N_711);
nor U1172 (N_1172,In_1452,N_658);
or U1173 (N_1173,N_291,In_1914);
xnor U1174 (N_1174,N_727,N_473);
or U1175 (N_1175,In_1401,In_1581);
and U1176 (N_1176,N_605,In_232);
xor U1177 (N_1177,In_1735,N_169);
nand U1178 (N_1178,In_492,In_293);
and U1179 (N_1179,N_253,N_15);
nor U1180 (N_1180,N_999,N_990);
or U1181 (N_1181,N_747,N_616);
nor U1182 (N_1182,In_1118,In_371);
and U1183 (N_1183,N_553,N_893);
nand U1184 (N_1184,In_1892,In_554);
nand U1185 (N_1185,N_929,In_1101);
or U1186 (N_1186,In_1207,N_329);
nand U1187 (N_1187,In_1333,N_398);
or U1188 (N_1188,N_992,In_1415);
and U1189 (N_1189,In_796,N_704);
nor U1190 (N_1190,In_497,In_357);
xnor U1191 (N_1191,In_115,N_232);
nor U1192 (N_1192,In_479,In_1752);
or U1193 (N_1193,N_121,N_297);
or U1194 (N_1194,In_1037,N_306);
xnor U1195 (N_1195,In_316,N_646);
nor U1196 (N_1196,N_494,N_459);
nor U1197 (N_1197,N_542,N_759);
nand U1198 (N_1198,N_733,N_872);
or U1199 (N_1199,N_822,N_989);
nor U1200 (N_1200,In_1609,N_850);
xor U1201 (N_1201,N_287,In_1346);
nand U1202 (N_1202,N_350,N_382);
nand U1203 (N_1203,In_1699,N_512);
or U1204 (N_1204,In_1755,In_1937);
nand U1205 (N_1205,N_508,N_397);
nor U1206 (N_1206,In_1195,N_109);
xor U1207 (N_1207,In_1521,N_533);
nand U1208 (N_1208,N_775,In_1988);
nand U1209 (N_1209,N_339,In_706);
nand U1210 (N_1210,N_505,N_837);
and U1211 (N_1211,N_933,N_931);
nor U1212 (N_1212,In_446,In_720);
xnor U1213 (N_1213,N_91,In_597);
nand U1214 (N_1214,In_981,N_961);
nand U1215 (N_1215,In_354,N_903);
or U1216 (N_1216,In_1438,N_79);
or U1217 (N_1217,N_80,In_754);
or U1218 (N_1218,In_1566,N_187);
xor U1219 (N_1219,N_934,In_688);
or U1220 (N_1220,In_978,In_1444);
nor U1221 (N_1221,In_404,In_1385);
nand U1222 (N_1222,N_479,N_207);
and U1223 (N_1223,In_1454,N_906);
nor U1224 (N_1224,In_122,N_673);
and U1225 (N_1225,In_1166,N_777);
nor U1226 (N_1226,In_669,In_1081);
nor U1227 (N_1227,N_610,N_958);
and U1228 (N_1228,N_975,N_523);
or U1229 (N_1229,In_1038,In_57);
or U1230 (N_1230,N_648,In_1932);
xor U1231 (N_1231,N_987,In_312);
and U1232 (N_1232,In_434,N_983);
nor U1233 (N_1233,N_845,N_812);
nor U1234 (N_1234,N_887,N_840);
or U1235 (N_1235,N_445,N_997);
nand U1236 (N_1236,N_443,N_751);
and U1237 (N_1237,N_633,N_885);
or U1238 (N_1238,N_90,N_922);
and U1239 (N_1239,N_629,N_698);
nor U1240 (N_1240,In_705,N_564);
and U1241 (N_1241,N_321,N_145);
and U1242 (N_1242,N_520,In_1242);
nand U1243 (N_1243,N_945,N_949);
or U1244 (N_1244,N_375,N_574);
nor U1245 (N_1245,N_250,N_829);
and U1246 (N_1246,In_89,In_722);
or U1247 (N_1247,N_973,In_213);
nand U1248 (N_1248,N_928,N_338);
nand U1249 (N_1249,In_341,N_978);
nand U1250 (N_1250,N_833,N_1208);
and U1251 (N_1251,N_368,N_710);
and U1252 (N_1252,N_785,N_661);
and U1253 (N_1253,N_1057,In_1162);
nand U1254 (N_1254,N_752,In_831);
and U1255 (N_1255,N_248,In_406);
xnor U1256 (N_1256,In_1967,In_763);
nand U1257 (N_1257,N_994,N_995);
or U1258 (N_1258,N_197,N_815);
or U1259 (N_1259,N_890,N_1214);
nand U1260 (N_1260,N_514,N_296);
xor U1261 (N_1261,N_649,N_1063);
or U1262 (N_1262,N_229,N_1116);
nand U1263 (N_1263,N_1216,N_1086);
and U1264 (N_1264,N_896,N_946);
nand U1265 (N_1265,N_1171,In_1600);
xor U1266 (N_1266,N_772,In_565);
or U1267 (N_1267,In_977,N_842);
xnor U1268 (N_1268,N_588,N_587);
or U1269 (N_1269,N_598,N_304);
and U1270 (N_1270,N_766,N_537);
nor U1271 (N_1271,In_830,N_789);
nand U1272 (N_1272,N_1215,N_1127);
nand U1273 (N_1273,In_1731,In_203);
nand U1274 (N_1274,N_754,N_1061);
or U1275 (N_1275,N_532,N_379);
nand U1276 (N_1276,In_454,N_1094);
or U1277 (N_1277,In_1368,N_1074);
and U1278 (N_1278,N_273,N_1198);
nand U1279 (N_1279,N_1050,In_204);
or U1280 (N_1280,In_29,N_351);
and U1281 (N_1281,N_1067,N_977);
xnor U1282 (N_1282,N_1095,N_818);
and U1283 (N_1283,N_870,In_395);
nor U1284 (N_1284,N_1017,N_652);
or U1285 (N_1285,N_1201,N_1130);
nor U1286 (N_1286,N_584,N_144);
or U1287 (N_1287,In_1623,In_1219);
and U1288 (N_1288,N_1218,N_1203);
nor U1289 (N_1289,N_1184,N_376);
or U1290 (N_1290,N_315,N_1245);
xor U1291 (N_1291,N_923,N_1142);
or U1292 (N_1292,N_1097,N_963);
nand U1293 (N_1293,In_270,N_1042);
nor U1294 (N_1294,In_1734,N_1001);
xor U1295 (N_1295,In_1736,N_911);
nand U1296 (N_1296,N_1158,In_1021);
or U1297 (N_1297,N_1128,N_621);
xnor U1298 (N_1298,N_1124,N_1070);
xnor U1299 (N_1299,N_1143,N_750);
and U1300 (N_1300,N_312,N_471);
nor U1301 (N_1301,N_787,N_876);
nand U1302 (N_1302,N_286,N_415);
or U1303 (N_1303,N_1029,N_1038);
and U1304 (N_1304,N_1110,N_1136);
or U1305 (N_1305,N_844,N_878);
and U1306 (N_1306,N_847,N_762);
or U1307 (N_1307,N_1153,N_868);
nand U1308 (N_1308,N_778,N_1241);
nand U1309 (N_1309,In_779,N_794);
xnor U1310 (N_1310,N_202,N_1019);
and U1311 (N_1311,N_1194,In_1426);
or U1312 (N_1312,In_1176,N_1103);
and U1313 (N_1313,N_734,N_180);
or U1314 (N_1314,N_549,In_940);
and U1315 (N_1315,N_1009,N_1000);
nand U1316 (N_1316,N_1034,N_477);
or U1317 (N_1317,In_709,N_1146);
nor U1318 (N_1318,In_1054,N_784);
and U1319 (N_1319,In_590,N_854);
xnor U1320 (N_1320,In_1186,N_506);
nand U1321 (N_1321,In_906,N_1210);
nor U1322 (N_1322,N_127,N_1167);
nor U1323 (N_1323,In_619,In_1846);
nand U1324 (N_1324,In_1493,N_1052);
or U1325 (N_1325,In_45,N_279);
nand U1326 (N_1326,N_1013,N_800);
xor U1327 (N_1327,N_1150,N_1186);
xnor U1328 (N_1328,In_463,N_937);
xnor U1329 (N_1329,N_786,N_1081);
xor U1330 (N_1330,N_1147,In_1547);
xnor U1331 (N_1331,N_1140,N_1005);
and U1332 (N_1332,N_1044,N_1166);
xnor U1333 (N_1333,N_1011,N_1162);
nor U1334 (N_1334,N_1020,N_1122);
xnor U1335 (N_1335,In_1954,In_150);
and U1336 (N_1336,In_551,N_1152);
nand U1337 (N_1337,In_824,N_1154);
nor U1338 (N_1338,N_1177,N_645);
and U1339 (N_1339,In_760,In_1765);
and U1340 (N_1340,N_969,N_439);
or U1341 (N_1341,In_1334,N_625);
and U1342 (N_1342,N_1060,N_450);
nor U1343 (N_1343,In_972,N_867);
and U1344 (N_1344,N_343,N_705);
or U1345 (N_1345,N_1040,N_1048);
and U1346 (N_1346,In_562,N_667);
nand U1347 (N_1347,N_1047,In_455);
nor U1348 (N_1348,N_484,N_1155);
nand U1349 (N_1349,N_612,In_1639);
nor U1350 (N_1350,In_1948,N_231);
nor U1351 (N_1351,In_1264,N_1102);
nor U1352 (N_1352,N_220,N_68);
nor U1353 (N_1353,N_939,In_1212);
xnor U1354 (N_1354,N_797,N_843);
nand U1355 (N_1355,N_150,In_462);
nand U1356 (N_1356,N_1098,N_666);
nor U1357 (N_1357,N_1242,N_1107);
nor U1358 (N_1358,N_469,N_223);
xnor U1359 (N_1359,N_736,N_292);
and U1360 (N_1360,In_585,N_407);
xor U1361 (N_1361,In_1126,N_1120);
xnor U1362 (N_1362,In_202,N_444);
nor U1363 (N_1363,N_1062,In_36);
nor U1364 (N_1364,N_1010,N_276);
xnor U1365 (N_1365,N_955,N_168);
nor U1366 (N_1366,N_1087,In_1715);
xor U1367 (N_1367,N_466,N_901);
or U1368 (N_1368,N_125,N_336);
or U1369 (N_1369,N_684,In_1888);
nor U1370 (N_1370,In_648,N_1224);
or U1371 (N_1371,In_771,N_1049);
and U1372 (N_1372,N_539,N_899);
nand U1373 (N_1373,N_1195,N_565);
nand U1374 (N_1374,N_1219,N_345);
xnor U1375 (N_1375,N_122,In_919);
or U1376 (N_1376,N_1243,N_432);
nor U1377 (N_1377,In_1422,N_798);
xor U1378 (N_1378,In_86,N_1002);
and U1379 (N_1379,N_1223,N_770);
nor U1380 (N_1380,In_1781,N_808);
and U1381 (N_1381,N_888,N_67);
xnor U1382 (N_1382,In_731,N_907);
xnor U1383 (N_1383,N_724,In_1768);
or U1384 (N_1384,In_1000,N_563);
and U1385 (N_1385,N_391,N_716);
or U1386 (N_1386,N_974,N_1185);
and U1387 (N_1387,N_354,In_1455);
nand U1388 (N_1388,N_1156,N_1021);
nand U1389 (N_1389,N_201,N_1132);
nor U1390 (N_1390,N_799,N_884);
nor U1391 (N_1391,N_991,N_803);
nor U1392 (N_1392,N_1077,In_1222);
or U1393 (N_1393,In_613,In_1378);
xnor U1394 (N_1394,N_1229,In_758);
and U1395 (N_1395,N_566,N_544);
nand U1396 (N_1396,N_1,N_1008);
and U1397 (N_1397,N_1016,N_1036);
or U1398 (N_1398,N_1073,N_806);
nand U1399 (N_1399,N_793,N_177);
nand U1400 (N_1400,N_1033,In_567);
and U1401 (N_1401,N_952,N_442);
or U1402 (N_1402,N_1083,In_1704);
or U1403 (N_1403,In_1800,N_1206);
or U1404 (N_1404,N_608,In_1541);
and U1405 (N_1405,N_597,N_1163);
xnor U1406 (N_1406,In_1742,N_1151);
or U1407 (N_1407,N_680,N_1159);
and U1408 (N_1408,In_414,In_997);
and U1409 (N_1409,N_260,N_1004);
or U1410 (N_1410,N_830,N_1192);
or U1411 (N_1411,In_1952,N_1188);
nor U1412 (N_1412,In_1467,N_1189);
xor U1413 (N_1413,N_936,N_1030);
or U1414 (N_1414,In_520,N_959);
or U1415 (N_1415,In_52,In_1690);
xnor U1416 (N_1416,N_1231,N_1091);
xor U1417 (N_1417,In_1268,N_964);
xor U1418 (N_1418,N_1069,In_1064);
xor U1419 (N_1419,N_1024,N_788);
nor U1420 (N_1420,In_330,N_1134);
or U1421 (N_1421,N_1031,In_1271);
xnor U1422 (N_1422,In_837,In_1572);
and U1423 (N_1423,N_1032,In_1531);
xnor U1424 (N_1424,N_768,N_1199);
and U1425 (N_1425,In_140,N_703);
and U1426 (N_1426,N_1157,N_1058);
nand U1427 (N_1427,N_988,N_862);
and U1428 (N_1428,N_981,In_1300);
or U1429 (N_1429,N_943,N_968);
or U1430 (N_1430,N_1149,In_1419);
or U1431 (N_1431,N_1173,N_1041);
nand U1432 (N_1432,N_701,N_1035);
and U1433 (N_1433,N_1100,N_1064);
and U1434 (N_1434,N_182,In_844);
xnor U1435 (N_1435,N_593,N_1172);
nand U1436 (N_1436,N_1138,N_1071);
xnor U1437 (N_1437,N_971,In_1536);
or U1438 (N_1438,N_264,In_670);
and U1439 (N_1439,N_1055,N_1072);
or U1440 (N_1440,N_467,In_1778);
or U1441 (N_1441,N_905,N_281);
nand U1442 (N_1442,In_396,N_263);
or U1443 (N_1443,N_1059,N_650);
and U1444 (N_1444,N_1205,N_653);
xor U1445 (N_1445,N_696,N_753);
or U1446 (N_1446,In_821,In_1903);
xnor U1447 (N_1447,N_1232,N_1211);
xnor U1448 (N_1448,N_1119,N_1204);
xor U1449 (N_1449,In_1510,N_124);
or U1450 (N_1450,N_58,N_3);
and U1451 (N_1451,In_1239,N_993);
or U1452 (N_1452,In_60,In_798);
and U1453 (N_1453,In_1210,N_1090);
nand U1454 (N_1454,N_1114,N_852);
or U1455 (N_1455,N_1075,N_41);
xnor U1456 (N_1456,N_1236,In_1766);
and U1457 (N_1457,In_432,N_1176);
xor U1458 (N_1458,N_1139,N_1093);
nand U1459 (N_1459,N_660,N_831);
nor U1460 (N_1460,N_846,N_628);
and U1461 (N_1461,N_932,In_1630);
xnor U1462 (N_1462,N_1169,N_918);
nand U1463 (N_1463,N_1141,N_26);
and U1464 (N_1464,N_1099,N_1088);
and U1465 (N_1465,N_365,N_1018);
and U1466 (N_1466,In_92,N_1113);
and U1467 (N_1467,N_668,N_998);
nand U1468 (N_1468,N_909,N_871);
or U1469 (N_1469,N_204,In_1381);
nor U1470 (N_1470,N_446,N_440);
nor U1471 (N_1471,N_1089,In_1777);
nand U1472 (N_1472,N_516,N_1239);
nor U1473 (N_1473,N_1170,N_856);
or U1474 (N_1474,N_496,N_357);
xnor U1475 (N_1475,In_1417,In_241);
xor U1476 (N_1476,N_956,N_1164);
and U1477 (N_1477,N_771,In_1040);
or U1478 (N_1478,N_1106,In_223);
nor U1479 (N_1479,N_441,In_898);
nand U1480 (N_1480,N_1015,N_813);
or U1481 (N_1481,N_702,N_435);
nand U1482 (N_1482,In_1662,N_33);
nor U1483 (N_1483,N_1217,N_1022);
or U1484 (N_1484,N_1202,N_941);
nor U1485 (N_1485,N_627,In_219);
xnor U1486 (N_1486,N_925,N_820);
xnor U1487 (N_1487,N_1117,N_1027);
and U1488 (N_1488,N_1144,N_1037);
xor U1489 (N_1489,N_1126,In_874);
or U1490 (N_1490,In_1974,In_1684);
or U1491 (N_1491,In_826,N_1054);
nand U1492 (N_1492,N_741,N_1065);
nand U1493 (N_1493,N_1207,N_828);
or U1494 (N_1494,N_1183,In_947);
and U1495 (N_1495,In_322,N_1109);
nor U1496 (N_1496,N_1179,In_1815);
nor U1497 (N_1497,N_919,In_1971);
nand U1498 (N_1498,In_1994,N_1080);
or U1499 (N_1499,N_462,N_855);
nor U1500 (N_1500,In_528,N_1327);
nor U1501 (N_1501,N_1442,N_601);
or U1502 (N_1502,N_1264,N_790);
xnor U1503 (N_1503,In_1168,N_1486);
nand U1504 (N_1504,N_1356,N_1237);
and U1505 (N_1505,N_839,N_1404);
and U1506 (N_1506,N_651,N_1388);
nand U1507 (N_1507,N_1307,N_1397);
xor U1508 (N_1508,N_1373,N_1181);
xor U1509 (N_1509,In_304,N_1359);
and U1510 (N_1510,In_1108,N_764);
or U1511 (N_1511,In_1727,N_571);
nand U1512 (N_1512,N_389,N_1414);
nor U1513 (N_1513,N_1437,N_1482);
or U1514 (N_1514,N_1360,N_1078);
or U1515 (N_1515,N_1449,N_824);
nor U1516 (N_1516,In_490,N_1393);
or U1517 (N_1517,In_1645,N_1368);
or U1518 (N_1518,In_1759,N_1481);
and U1519 (N_1519,N_1460,N_1366);
xnor U1520 (N_1520,N_1056,N_1485);
and U1521 (N_1521,N_1455,N_886);
and U1522 (N_1522,N_1478,N_1369);
nor U1523 (N_1523,N_1253,N_1160);
nor U1524 (N_1524,In_1865,N_1274);
xnor U1525 (N_1525,In_1842,N_1007);
or U1526 (N_1526,N_1329,N_1263);
and U1527 (N_1527,N_1323,N_1240);
nand U1528 (N_1528,N_1082,N_796);
or U1529 (N_1529,N_531,N_1299);
and U1530 (N_1530,In_1901,N_1084);
nand U1531 (N_1531,N_1301,N_1330);
nand U1532 (N_1532,N_1129,N_1303);
nor U1533 (N_1533,N_1310,N_1374);
and U1534 (N_1534,N_620,N_1466);
nand U1535 (N_1535,N_1441,N_1389);
nand U1536 (N_1536,In_890,In_1167);
nand U1537 (N_1537,N_1249,N_1398);
nor U1538 (N_1538,N_1358,In_361);
xor U1539 (N_1539,N_1324,N_1465);
xnor U1540 (N_1540,N_1182,N_1079);
xor U1541 (N_1541,In_1569,N_1238);
xor U1542 (N_1542,In_487,N_1321);
or U1543 (N_1543,N_1292,N_1353);
nor U1544 (N_1544,N_1496,In_1802);
xnor U1545 (N_1545,N_1339,N_449);
and U1546 (N_1546,N_1262,N_1318);
xnor U1547 (N_1547,N_1340,N_409);
xor U1548 (N_1548,N_1252,N_1295);
or U1549 (N_1549,N_1380,N_897);
xnor U1550 (N_1550,N_728,N_756);
and U1551 (N_1551,In_290,N_1430);
or U1552 (N_1552,N_288,In_915);
nand U1553 (N_1553,N_1355,N_1428);
xor U1554 (N_1554,N_1469,In_668);
xnor U1555 (N_1555,N_1424,N_1338);
xor U1556 (N_1556,N_1385,In_1193);
or U1557 (N_1557,N_1213,N_692);
nor U1558 (N_1558,N_1480,N_1448);
and U1559 (N_1559,N_1101,N_1375);
and U1560 (N_1560,N_1335,In_1326);
nor U1561 (N_1561,In_21,N_1168);
nand U1562 (N_1562,In_1588,N_1367);
or U1563 (N_1563,N_386,N_1279);
and U1564 (N_1564,In_1873,N_1288);
and U1565 (N_1565,N_1248,N_1246);
nand U1566 (N_1566,N_910,N_1125);
nor U1567 (N_1567,N_1422,N_1121);
or U1568 (N_1568,N_1476,N_1025);
and U1569 (N_1569,N_801,N_1347);
xor U1570 (N_1570,N_1410,N_1311);
and U1571 (N_1571,N_1436,N_1402);
or U1572 (N_1572,N_1406,In_1871);
xor U1573 (N_1573,N_1439,N_807);
and U1574 (N_1574,N_1377,N_678);
and U1575 (N_1575,N_1003,N_1386);
nand U1576 (N_1576,N_1337,In_1482);
nand U1577 (N_1577,In_1511,In_1582);
xnor U1578 (N_1578,In_1558,N_1227);
or U1579 (N_1579,N_1302,In_761);
and U1580 (N_1580,In_510,N_675);
xor U1581 (N_1581,N_1419,N_1450);
and U1582 (N_1582,In_1311,N_73);
and U1583 (N_1583,In_966,In_1829);
and U1584 (N_1584,N_1470,N_1118);
nand U1585 (N_1585,N_1417,N_5);
and U1586 (N_1586,N_1443,N_1372);
and U1587 (N_1587,In_1780,N_1275);
nand U1588 (N_1588,N_781,N_1332);
nand U1589 (N_1589,N_1453,N_1461);
or U1590 (N_1590,N_805,In_1361);
and U1591 (N_1591,N_1497,In_1430);
or U1592 (N_1592,N_917,N_326);
or U1593 (N_1593,N_1278,N_865);
nand U1594 (N_1594,N_1115,In_1807);
and U1595 (N_1595,N_1255,N_1221);
nor U1596 (N_1596,N_1438,N_1379);
nor U1597 (N_1597,N_1317,N_194);
or U1598 (N_1598,N_1467,N_1413);
nor U1599 (N_1599,N_1297,N_1313);
and U1600 (N_1600,N_387,In_1147);
nor U1601 (N_1601,N_1357,N_1220);
nand U1602 (N_1602,N_1391,N_1068);
nor U1603 (N_1603,N_1350,N_1306);
nand U1604 (N_1604,In_194,N_1371);
nor U1605 (N_1605,N_1346,N_1174);
and U1606 (N_1606,N_275,N_1085);
or U1607 (N_1607,N_1468,N_758);
and U1608 (N_1608,N_1235,N_1191);
and U1609 (N_1609,In_1440,N_1344);
nor U1610 (N_1610,N_1363,N_1226);
or U1611 (N_1611,N_1309,N_1187);
xor U1612 (N_1612,N_1429,N_1490);
nor U1613 (N_1613,In_426,N_655);
xnor U1614 (N_1614,In_968,N_1014);
and U1615 (N_1615,N_1361,N_823);
or U1616 (N_1616,In_40,In_1411);
nand U1617 (N_1617,N_1270,N_1331);
nand U1618 (N_1618,N_1484,In_1820);
nor U1619 (N_1619,N_792,N_1412);
xnor U1620 (N_1620,N_1180,N_944);
xor U1621 (N_1621,N_1425,N_1294);
xnor U1622 (N_1622,N_1325,N_1390);
nand U1623 (N_1623,N_1043,N_1462);
nor U1624 (N_1624,In_572,N_1328);
nor U1625 (N_1625,N_1477,N_848);
xnor U1626 (N_1626,N_1423,N_1259);
xor U1627 (N_1627,N_691,N_1026);
xnor U1628 (N_1628,N_1105,N_1400);
nand U1629 (N_1629,N_1251,N_8);
and U1630 (N_1630,N_1315,N_1399);
or U1631 (N_1631,N_1394,N_1351);
nand U1632 (N_1632,N_1387,In_1769);
nor U1633 (N_1633,N_1108,N_1433);
or U1634 (N_1634,N_1256,N_1383);
or U1635 (N_1635,In_310,N_582);
xor U1636 (N_1636,N_1258,N_1492);
nand U1637 (N_1637,N_1305,N_1104);
and U1638 (N_1638,N_1092,N_1193);
nor U1639 (N_1639,N_1463,N_1341);
nor U1640 (N_1640,N_1348,N_1096);
nand U1641 (N_1641,N_1244,N_717);
nand U1642 (N_1642,N_1268,N_996);
nand U1643 (N_1643,N_1283,N_1434);
or U1644 (N_1644,In_1869,N_1230);
or U1645 (N_1645,N_1407,N_1234);
nor U1646 (N_1646,N_1472,In_1409);
nor U1647 (N_1647,N_1365,N_1308);
and U1648 (N_1648,N_575,N_731);
xor U1649 (N_1649,N_1261,N_1137);
and U1650 (N_1650,N_1376,N_1290);
xor U1651 (N_1651,In_1589,N_1431);
xnor U1652 (N_1652,N_1494,In_863);
and U1653 (N_1653,N_1267,N_1474);
nor U1654 (N_1654,N_1284,N_1281);
nand U1655 (N_1655,N_773,N_1479);
or U1656 (N_1656,In_386,N_1418);
or U1657 (N_1657,N_423,N_1291);
xnor U1658 (N_1658,N_1420,In_1408);
and U1659 (N_1659,N_1498,In_1619);
nor U1660 (N_1660,N_1405,N_1475);
and U1661 (N_1661,N_1370,N_1260);
and U1662 (N_1662,N_1432,N_1445);
and U1663 (N_1663,N_1271,N_1345);
or U1664 (N_1664,N_1464,N_694);
or U1665 (N_1665,N_1028,N_1415);
nand U1666 (N_1666,N_1272,N_349);
or U1667 (N_1667,N_1190,N_1196);
xor U1668 (N_1668,N_769,N_1326);
xor U1669 (N_1669,N_1403,N_810);
nand U1670 (N_1670,N_256,N_1392);
and U1671 (N_1671,N_1320,N_1225);
xnor U1672 (N_1672,N_748,In_1142);
nor U1673 (N_1673,N_1487,In_248);
or U1674 (N_1674,N_1212,In_570);
and U1675 (N_1675,N_915,N_1333);
nor U1676 (N_1676,In_200,N_1440);
and U1677 (N_1677,N_1289,N_1458);
xor U1678 (N_1678,N_1488,N_1378);
or U1679 (N_1679,In_166,N_1045);
or U1680 (N_1680,In_1724,In_1288);
and U1681 (N_1681,In_738,N_1381);
and U1682 (N_1682,N_1273,N_581);
or U1683 (N_1683,N_1499,N_1456);
and U1684 (N_1684,N_1312,N_1300);
nand U1685 (N_1685,N_199,N_1266);
or U1686 (N_1686,N_1197,N_1316);
xnor U1687 (N_1687,N_1111,N_1012);
and U1688 (N_1688,N_424,In_579);
xor U1689 (N_1689,N_1233,N_1451);
nand U1690 (N_1690,N_1265,In_609);
and U1691 (N_1691,N_1175,N_1286);
or U1692 (N_1692,N_1421,N_1200);
xor U1693 (N_1693,N_1444,N_1066);
xnor U1694 (N_1694,N_1457,N_1408);
or U1695 (N_1695,In_56,In_85);
or U1696 (N_1696,N_1352,N_1051);
nor U1697 (N_1697,N_72,N_1452);
or U1698 (N_1698,N_1416,N_1336);
nor U1699 (N_1699,N_1257,N_1495);
nand U1700 (N_1700,N_1384,N_1131);
nor U1701 (N_1701,N_1349,N_75);
and U1702 (N_1702,N_1427,N_774);
or U1703 (N_1703,N_1322,N_1411);
and U1704 (N_1704,N_1343,In_642);
nand U1705 (N_1705,In_957,N_1489);
or U1706 (N_1706,N_882,N_1023);
xnor U1707 (N_1707,N_1250,N_1277);
xor U1708 (N_1708,In_1860,N_1269);
xor U1709 (N_1709,N_1454,N_743);
or U1710 (N_1710,N_706,N_866);
and U1711 (N_1711,N_1039,N_1254);
nand U1712 (N_1712,N_732,N_216);
and U1713 (N_1713,N_1178,N_1364);
nor U1714 (N_1714,N_851,N_1409);
nand U1715 (N_1715,N_1447,N_1053);
nor U1716 (N_1716,In_35,N_1123);
xor U1717 (N_1717,N_1435,N_464);
xor U1718 (N_1718,N_1491,N_1222);
xnor U1719 (N_1719,N_1362,N_1247);
nand U1720 (N_1720,N_495,N_1287);
xor U1721 (N_1721,N_225,N_1293);
nand U1722 (N_1722,N_1276,N_1161);
nor U1723 (N_1723,N_100,N_1006);
nand U1724 (N_1724,N_966,N_1493);
or U1725 (N_1725,N_1228,N_1148);
nor U1726 (N_1726,N_1334,N_1285);
and U1727 (N_1727,N_1135,N_1298);
nor U1728 (N_1728,N_1483,N_1076);
or U1729 (N_1729,N_1446,N_864);
xnor U1730 (N_1730,In_825,N_926);
and U1731 (N_1731,N_1401,N_1426);
and U1732 (N_1732,N_745,N_241);
nand U1733 (N_1733,N_749,N_163);
or U1734 (N_1734,In_740,N_1354);
nand U1735 (N_1735,In_1853,N_1282);
nor U1736 (N_1736,In_546,N_1342);
nor U1737 (N_1737,N_1396,N_1280);
xnor U1738 (N_1738,N_1395,N_914);
xnor U1739 (N_1739,N_1296,In_1286);
and U1740 (N_1740,N_1459,N_1319);
nor U1741 (N_1741,N_503,N_1112);
and U1742 (N_1742,N_960,In_1697);
or U1743 (N_1743,N_1382,N_1473);
nand U1744 (N_1744,N_1314,In_1078);
or U1745 (N_1745,N_573,N_1133);
or U1746 (N_1746,N_1209,N_942);
or U1747 (N_1747,N_1145,N_1304);
nor U1748 (N_1748,In_607,N_1471);
and U1749 (N_1749,N_1165,N_1046);
nor U1750 (N_1750,N_1516,N_1582);
and U1751 (N_1751,N_1648,N_1689);
and U1752 (N_1752,N_1732,N_1719);
or U1753 (N_1753,N_1693,N_1527);
nor U1754 (N_1754,N_1681,N_1548);
nor U1755 (N_1755,N_1581,N_1696);
and U1756 (N_1756,N_1662,N_1700);
and U1757 (N_1757,N_1637,N_1654);
and U1758 (N_1758,N_1503,N_1640);
nand U1759 (N_1759,N_1566,N_1562);
nand U1760 (N_1760,N_1743,N_1513);
xor U1761 (N_1761,N_1567,N_1564);
nor U1762 (N_1762,N_1694,N_1603);
nor U1763 (N_1763,N_1716,N_1616);
nor U1764 (N_1764,N_1545,N_1673);
xnor U1765 (N_1765,N_1531,N_1553);
nand U1766 (N_1766,N_1680,N_1702);
or U1767 (N_1767,N_1735,N_1733);
nand U1768 (N_1768,N_1661,N_1524);
xor U1769 (N_1769,N_1738,N_1505);
or U1770 (N_1770,N_1622,N_1526);
nor U1771 (N_1771,N_1744,N_1723);
and U1772 (N_1772,N_1560,N_1515);
or U1773 (N_1773,N_1592,N_1583);
xor U1774 (N_1774,N_1659,N_1739);
nand U1775 (N_1775,N_1725,N_1520);
or U1776 (N_1776,N_1722,N_1577);
xnor U1777 (N_1777,N_1610,N_1575);
and U1778 (N_1778,N_1542,N_1502);
nor U1779 (N_1779,N_1549,N_1550);
or U1780 (N_1780,N_1574,N_1703);
or U1781 (N_1781,N_1538,N_1580);
or U1782 (N_1782,N_1593,N_1585);
xnor U1783 (N_1783,N_1709,N_1589);
and U1784 (N_1784,N_1741,N_1596);
xnor U1785 (N_1785,N_1563,N_1555);
xnor U1786 (N_1786,N_1736,N_1657);
nor U1787 (N_1787,N_1628,N_1664);
xor U1788 (N_1788,N_1539,N_1641);
xor U1789 (N_1789,N_1706,N_1587);
nand U1790 (N_1790,N_1626,N_1740);
and U1791 (N_1791,N_1636,N_1646);
and U1792 (N_1792,N_1650,N_1525);
xor U1793 (N_1793,N_1543,N_1708);
nor U1794 (N_1794,N_1670,N_1509);
nor U1795 (N_1795,N_1554,N_1615);
or U1796 (N_1796,N_1727,N_1551);
nor U1797 (N_1797,N_1695,N_1726);
or U1798 (N_1798,N_1621,N_1588);
nand U1799 (N_1799,N_1715,N_1547);
or U1800 (N_1800,N_1537,N_1688);
and U1801 (N_1801,N_1678,N_1532);
and U1802 (N_1802,N_1660,N_1675);
and U1803 (N_1803,N_1734,N_1519);
or U1804 (N_1804,N_1720,N_1748);
xnor U1805 (N_1805,N_1541,N_1728);
nand U1806 (N_1806,N_1643,N_1565);
and U1807 (N_1807,N_1528,N_1644);
and U1808 (N_1808,N_1668,N_1552);
nand U1809 (N_1809,N_1511,N_1672);
xor U1810 (N_1810,N_1590,N_1690);
and U1811 (N_1811,N_1514,N_1571);
nand U1812 (N_1812,N_1546,N_1612);
and U1813 (N_1813,N_1609,N_1620);
nor U1814 (N_1814,N_1572,N_1500);
and U1815 (N_1815,N_1512,N_1704);
nand U1816 (N_1816,N_1651,N_1721);
nand U1817 (N_1817,N_1676,N_1606);
nand U1818 (N_1818,N_1599,N_1604);
and U1819 (N_1819,N_1602,N_1578);
nand U1820 (N_1820,N_1698,N_1679);
xor U1821 (N_1821,N_1718,N_1629);
nand U1822 (N_1822,N_1559,N_1623);
xnor U1823 (N_1823,N_1665,N_1507);
or U1824 (N_1824,N_1749,N_1652);
and U1825 (N_1825,N_1501,N_1710);
nor U1826 (N_1826,N_1614,N_1663);
or U1827 (N_1827,N_1597,N_1510);
and U1828 (N_1828,N_1627,N_1687);
or U1829 (N_1829,N_1685,N_1624);
and U1830 (N_1830,N_1642,N_1529);
nor U1831 (N_1831,N_1669,N_1686);
nor U1832 (N_1832,N_1535,N_1747);
or U1833 (N_1833,N_1724,N_1534);
nand U1834 (N_1834,N_1713,N_1619);
xnor U1835 (N_1835,N_1584,N_1711);
xor U1836 (N_1836,N_1714,N_1607);
nor U1837 (N_1837,N_1717,N_1625);
or U1838 (N_1838,N_1608,N_1617);
xnor U1839 (N_1839,N_1691,N_1518);
or U1840 (N_1840,N_1558,N_1600);
xor U1841 (N_1841,N_1656,N_1645);
nor U1842 (N_1842,N_1568,N_1674);
nor U1843 (N_1843,N_1692,N_1533);
and U1844 (N_1844,N_1536,N_1638);
xnor U1845 (N_1845,N_1522,N_1540);
and U1846 (N_1846,N_1634,N_1556);
nor U1847 (N_1847,N_1729,N_1705);
xnor U1848 (N_1848,N_1666,N_1506);
xnor U1849 (N_1849,N_1517,N_1521);
xnor U1850 (N_1850,N_1569,N_1635);
or U1851 (N_1851,N_1570,N_1595);
and U1852 (N_1852,N_1649,N_1707);
nor U1853 (N_1853,N_1697,N_1586);
nor U1854 (N_1854,N_1667,N_1658);
nor U1855 (N_1855,N_1630,N_1737);
or U1856 (N_1856,N_1576,N_1653);
xnor U1857 (N_1857,N_1684,N_1639);
nor U1858 (N_1858,N_1730,N_1632);
nor U1859 (N_1859,N_1699,N_1605);
xor U1860 (N_1860,N_1647,N_1682);
nand U1861 (N_1861,N_1544,N_1508);
or U1862 (N_1862,N_1557,N_1683);
and U1863 (N_1863,N_1677,N_1561);
and U1864 (N_1864,N_1655,N_1742);
or U1865 (N_1865,N_1504,N_1591);
nand U1866 (N_1866,N_1530,N_1731);
xnor U1867 (N_1867,N_1611,N_1631);
nand U1868 (N_1868,N_1745,N_1712);
and U1869 (N_1869,N_1601,N_1701);
and U1870 (N_1870,N_1618,N_1594);
nand U1871 (N_1871,N_1746,N_1671);
nor U1872 (N_1872,N_1598,N_1633);
nand U1873 (N_1873,N_1579,N_1523);
xnor U1874 (N_1874,N_1573,N_1613);
and U1875 (N_1875,N_1642,N_1743);
xor U1876 (N_1876,N_1660,N_1591);
nor U1877 (N_1877,N_1740,N_1531);
nor U1878 (N_1878,N_1624,N_1539);
nor U1879 (N_1879,N_1704,N_1662);
nor U1880 (N_1880,N_1622,N_1640);
or U1881 (N_1881,N_1713,N_1516);
nor U1882 (N_1882,N_1722,N_1535);
and U1883 (N_1883,N_1643,N_1742);
nor U1884 (N_1884,N_1715,N_1682);
or U1885 (N_1885,N_1570,N_1707);
and U1886 (N_1886,N_1606,N_1712);
nor U1887 (N_1887,N_1645,N_1589);
or U1888 (N_1888,N_1672,N_1553);
nor U1889 (N_1889,N_1503,N_1729);
nand U1890 (N_1890,N_1501,N_1722);
or U1891 (N_1891,N_1672,N_1681);
xor U1892 (N_1892,N_1747,N_1631);
and U1893 (N_1893,N_1660,N_1635);
nor U1894 (N_1894,N_1568,N_1737);
or U1895 (N_1895,N_1645,N_1722);
xor U1896 (N_1896,N_1687,N_1594);
and U1897 (N_1897,N_1652,N_1721);
nor U1898 (N_1898,N_1673,N_1631);
xor U1899 (N_1899,N_1665,N_1515);
and U1900 (N_1900,N_1600,N_1640);
or U1901 (N_1901,N_1511,N_1610);
or U1902 (N_1902,N_1507,N_1634);
or U1903 (N_1903,N_1694,N_1658);
and U1904 (N_1904,N_1695,N_1575);
and U1905 (N_1905,N_1536,N_1589);
nor U1906 (N_1906,N_1639,N_1566);
nand U1907 (N_1907,N_1518,N_1712);
xor U1908 (N_1908,N_1644,N_1586);
nand U1909 (N_1909,N_1558,N_1721);
nand U1910 (N_1910,N_1714,N_1685);
xnor U1911 (N_1911,N_1683,N_1723);
nor U1912 (N_1912,N_1708,N_1684);
nor U1913 (N_1913,N_1658,N_1549);
and U1914 (N_1914,N_1532,N_1577);
and U1915 (N_1915,N_1590,N_1557);
and U1916 (N_1916,N_1580,N_1662);
or U1917 (N_1917,N_1608,N_1669);
or U1918 (N_1918,N_1702,N_1590);
xor U1919 (N_1919,N_1538,N_1722);
and U1920 (N_1920,N_1573,N_1615);
nand U1921 (N_1921,N_1638,N_1700);
xor U1922 (N_1922,N_1680,N_1585);
nor U1923 (N_1923,N_1528,N_1517);
nor U1924 (N_1924,N_1662,N_1654);
nor U1925 (N_1925,N_1601,N_1653);
xnor U1926 (N_1926,N_1718,N_1524);
nand U1927 (N_1927,N_1721,N_1668);
and U1928 (N_1928,N_1661,N_1704);
and U1929 (N_1929,N_1696,N_1614);
and U1930 (N_1930,N_1506,N_1635);
or U1931 (N_1931,N_1742,N_1514);
or U1932 (N_1932,N_1529,N_1608);
nand U1933 (N_1933,N_1609,N_1544);
xor U1934 (N_1934,N_1703,N_1658);
xor U1935 (N_1935,N_1748,N_1544);
nor U1936 (N_1936,N_1746,N_1699);
or U1937 (N_1937,N_1564,N_1629);
and U1938 (N_1938,N_1712,N_1508);
or U1939 (N_1939,N_1520,N_1502);
nor U1940 (N_1940,N_1673,N_1686);
xor U1941 (N_1941,N_1730,N_1649);
nand U1942 (N_1942,N_1512,N_1587);
nor U1943 (N_1943,N_1507,N_1696);
and U1944 (N_1944,N_1615,N_1627);
and U1945 (N_1945,N_1540,N_1560);
nor U1946 (N_1946,N_1699,N_1704);
nor U1947 (N_1947,N_1726,N_1583);
nor U1948 (N_1948,N_1729,N_1672);
xor U1949 (N_1949,N_1604,N_1643);
and U1950 (N_1950,N_1629,N_1549);
or U1951 (N_1951,N_1507,N_1571);
or U1952 (N_1952,N_1713,N_1549);
and U1953 (N_1953,N_1715,N_1740);
xor U1954 (N_1954,N_1655,N_1533);
xor U1955 (N_1955,N_1675,N_1677);
nor U1956 (N_1956,N_1673,N_1675);
nand U1957 (N_1957,N_1521,N_1597);
xor U1958 (N_1958,N_1505,N_1612);
nand U1959 (N_1959,N_1653,N_1670);
nand U1960 (N_1960,N_1610,N_1640);
xnor U1961 (N_1961,N_1698,N_1524);
xor U1962 (N_1962,N_1581,N_1518);
and U1963 (N_1963,N_1670,N_1503);
nand U1964 (N_1964,N_1597,N_1694);
and U1965 (N_1965,N_1644,N_1739);
nor U1966 (N_1966,N_1520,N_1631);
nand U1967 (N_1967,N_1588,N_1733);
nor U1968 (N_1968,N_1546,N_1543);
xnor U1969 (N_1969,N_1619,N_1569);
or U1970 (N_1970,N_1595,N_1546);
nand U1971 (N_1971,N_1606,N_1613);
nor U1972 (N_1972,N_1658,N_1691);
and U1973 (N_1973,N_1660,N_1588);
nor U1974 (N_1974,N_1720,N_1560);
nor U1975 (N_1975,N_1504,N_1641);
xnor U1976 (N_1976,N_1714,N_1670);
nand U1977 (N_1977,N_1722,N_1534);
nand U1978 (N_1978,N_1585,N_1683);
nand U1979 (N_1979,N_1730,N_1503);
nor U1980 (N_1980,N_1519,N_1660);
and U1981 (N_1981,N_1515,N_1525);
nor U1982 (N_1982,N_1526,N_1632);
and U1983 (N_1983,N_1621,N_1666);
nor U1984 (N_1984,N_1631,N_1698);
xor U1985 (N_1985,N_1508,N_1742);
and U1986 (N_1986,N_1663,N_1508);
nor U1987 (N_1987,N_1634,N_1582);
xor U1988 (N_1988,N_1687,N_1604);
nand U1989 (N_1989,N_1515,N_1584);
or U1990 (N_1990,N_1613,N_1557);
xnor U1991 (N_1991,N_1631,N_1540);
nor U1992 (N_1992,N_1519,N_1708);
nand U1993 (N_1993,N_1510,N_1541);
nor U1994 (N_1994,N_1586,N_1606);
nand U1995 (N_1995,N_1666,N_1512);
or U1996 (N_1996,N_1669,N_1534);
nor U1997 (N_1997,N_1637,N_1557);
xnor U1998 (N_1998,N_1522,N_1576);
nor U1999 (N_1999,N_1673,N_1560);
and U2000 (N_2000,N_1789,N_1760);
nor U2001 (N_2001,N_1781,N_1862);
or U2002 (N_2002,N_1922,N_1985);
nand U2003 (N_2003,N_1821,N_1970);
and U2004 (N_2004,N_1886,N_1990);
or U2005 (N_2005,N_1841,N_1899);
or U2006 (N_2006,N_1939,N_1795);
nand U2007 (N_2007,N_1910,N_1943);
or U2008 (N_2008,N_1796,N_1892);
nor U2009 (N_2009,N_1881,N_1914);
xnor U2010 (N_2010,N_1870,N_1843);
xnor U2011 (N_2011,N_1938,N_1890);
xor U2012 (N_2012,N_1882,N_1895);
or U2013 (N_2013,N_1949,N_1983);
nor U2014 (N_2014,N_1995,N_1942);
xor U2015 (N_2015,N_1957,N_1889);
nor U2016 (N_2016,N_1758,N_1915);
and U2017 (N_2017,N_1863,N_1997);
nor U2018 (N_2018,N_1878,N_1896);
nor U2019 (N_2019,N_1754,N_1794);
xor U2020 (N_2020,N_1903,N_1989);
or U2021 (N_2021,N_1857,N_1880);
or U2022 (N_2022,N_1973,N_1822);
nor U2023 (N_2023,N_1991,N_1996);
nand U2024 (N_2024,N_1944,N_1907);
and U2025 (N_2025,N_1993,N_1972);
nand U2026 (N_2026,N_1798,N_1877);
and U2027 (N_2027,N_1906,N_1766);
or U2028 (N_2028,N_1844,N_1848);
nor U2029 (N_2029,N_1946,N_1842);
xor U2030 (N_2030,N_1975,N_1780);
nand U2031 (N_2031,N_1787,N_1810);
and U2032 (N_2032,N_1858,N_1778);
xnor U2033 (N_2033,N_1790,N_1904);
nand U2034 (N_2034,N_1969,N_1820);
nor U2035 (N_2035,N_1759,N_1828);
nor U2036 (N_2036,N_1918,N_1998);
or U2037 (N_2037,N_1873,N_1976);
nor U2038 (N_2038,N_1913,N_1967);
or U2039 (N_2039,N_1813,N_1869);
and U2040 (N_2040,N_1901,N_1804);
nor U2041 (N_2041,N_1835,N_1819);
xor U2042 (N_2042,N_1847,N_1920);
nor U2043 (N_2043,N_1935,N_1808);
nand U2044 (N_2044,N_1802,N_1925);
and U2045 (N_2045,N_1854,N_1788);
or U2046 (N_2046,N_1897,N_1962);
nor U2047 (N_2047,N_1921,N_1966);
nor U2048 (N_2048,N_1950,N_1782);
nand U2049 (N_2049,N_1948,N_1927);
nand U2050 (N_2050,N_1887,N_1981);
or U2051 (N_2051,N_1865,N_1876);
nor U2052 (N_2052,N_1829,N_1784);
xor U2053 (N_2053,N_1814,N_1963);
nand U2054 (N_2054,N_1791,N_1987);
or U2055 (N_2055,N_1785,N_1960);
nand U2056 (N_2056,N_1752,N_1928);
or U2057 (N_2057,N_1774,N_1955);
and U2058 (N_2058,N_1786,N_1815);
and U2059 (N_2059,N_1964,N_1959);
nor U2060 (N_2060,N_1909,N_1853);
or U2061 (N_2061,N_1980,N_1974);
or U2062 (N_2062,N_1867,N_1883);
or U2063 (N_2063,N_1879,N_1768);
nand U2064 (N_2064,N_1750,N_1864);
nor U2065 (N_2065,N_1793,N_1917);
xor U2066 (N_2066,N_1958,N_1803);
xor U2067 (N_2067,N_1860,N_1941);
nor U2068 (N_2068,N_1763,N_1838);
xnor U2069 (N_2069,N_1806,N_1769);
xnor U2070 (N_2070,N_1851,N_1827);
and U2071 (N_2071,N_1805,N_1840);
nor U2072 (N_2072,N_1900,N_1850);
xor U2073 (N_2073,N_1764,N_1816);
nor U2074 (N_2074,N_1894,N_1846);
xnor U2075 (N_2075,N_1797,N_1773);
and U2076 (N_2076,N_1856,N_1994);
nand U2077 (N_2077,N_1839,N_1905);
or U2078 (N_2078,N_1872,N_1845);
or U2079 (N_2079,N_1931,N_1971);
xnor U2080 (N_2080,N_1898,N_1902);
nor U2081 (N_2081,N_1888,N_1826);
xor U2082 (N_2082,N_1751,N_1923);
nand U2083 (N_2083,N_1947,N_1837);
xor U2084 (N_2084,N_1954,N_1982);
nand U2085 (N_2085,N_1792,N_1929);
or U2086 (N_2086,N_1908,N_1823);
nand U2087 (N_2087,N_1753,N_1940);
xor U2088 (N_2088,N_1937,N_1765);
or U2089 (N_2089,N_1761,N_1932);
xor U2090 (N_2090,N_1800,N_1830);
xnor U2091 (N_2091,N_1912,N_1926);
and U2092 (N_2092,N_1783,N_1777);
nand U2093 (N_2093,N_1965,N_1911);
nand U2094 (N_2094,N_1836,N_1809);
or U2095 (N_2095,N_1916,N_1859);
or U2096 (N_2096,N_1919,N_1885);
and U2097 (N_2097,N_1945,N_1861);
and U2098 (N_2098,N_1755,N_1776);
nor U2099 (N_2099,N_1825,N_1817);
nand U2100 (N_2100,N_1855,N_1762);
and U2101 (N_2101,N_1871,N_1884);
or U2102 (N_2102,N_1866,N_1756);
nand U2103 (N_2103,N_1952,N_1951);
xor U2104 (N_2104,N_1767,N_1868);
nand U2105 (N_2105,N_1934,N_1924);
nand U2106 (N_2106,N_1961,N_1968);
or U2107 (N_2107,N_1933,N_1936);
nor U2108 (N_2108,N_1807,N_1875);
and U2109 (N_2109,N_1852,N_1893);
nor U2110 (N_2110,N_1977,N_1757);
nand U2111 (N_2111,N_1986,N_1999);
or U2112 (N_2112,N_1770,N_1833);
nand U2113 (N_2113,N_1978,N_1930);
or U2114 (N_2114,N_1818,N_1984);
or U2115 (N_2115,N_1988,N_1956);
nand U2116 (N_2116,N_1799,N_1849);
or U2117 (N_2117,N_1832,N_1771);
nor U2118 (N_2118,N_1953,N_1772);
or U2119 (N_2119,N_1831,N_1812);
or U2120 (N_2120,N_1811,N_1979);
nand U2121 (N_2121,N_1801,N_1779);
nand U2122 (N_2122,N_1992,N_1874);
and U2123 (N_2123,N_1824,N_1834);
or U2124 (N_2124,N_1775,N_1891);
nand U2125 (N_2125,N_1802,N_1789);
nand U2126 (N_2126,N_1937,N_1770);
nand U2127 (N_2127,N_1955,N_1792);
nor U2128 (N_2128,N_1866,N_1755);
and U2129 (N_2129,N_1786,N_1966);
xnor U2130 (N_2130,N_1784,N_1859);
xor U2131 (N_2131,N_1790,N_1927);
nand U2132 (N_2132,N_1980,N_1759);
or U2133 (N_2133,N_1936,N_1903);
xor U2134 (N_2134,N_1909,N_1941);
and U2135 (N_2135,N_1801,N_1803);
and U2136 (N_2136,N_1785,N_1790);
nand U2137 (N_2137,N_1839,N_1881);
or U2138 (N_2138,N_1932,N_1902);
nand U2139 (N_2139,N_1834,N_1905);
nor U2140 (N_2140,N_1992,N_1962);
nand U2141 (N_2141,N_1872,N_1750);
nand U2142 (N_2142,N_1864,N_1820);
and U2143 (N_2143,N_1781,N_1756);
xor U2144 (N_2144,N_1873,N_1824);
or U2145 (N_2145,N_1802,N_1785);
nor U2146 (N_2146,N_1899,N_1976);
nand U2147 (N_2147,N_1937,N_1923);
nand U2148 (N_2148,N_1957,N_1816);
nor U2149 (N_2149,N_1880,N_1950);
xor U2150 (N_2150,N_1981,N_1771);
nor U2151 (N_2151,N_1975,N_1883);
or U2152 (N_2152,N_1833,N_1992);
and U2153 (N_2153,N_1777,N_1799);
nor U2154 (N_2154,N_1980,N_1922);
or U2155 (N_2155,N_1874,N_1920);
and U2156 (N_2156,N_1820,N_1914);
and U2157 (N_2157,N_1884,N_1820);
and U2158 (N_2158,N_1757,N_1759);
nor U2159 (N_2159,N_1812,N_1961);
or U2160 (N_2160,N_1846,N_1942);
xor U2161 (N_2161,N_1966,N_1972);
and U2162 (N_2162,N_1894,N_1784);
and U2163 (N_2163,N_1910,N_1830);
nand U2164 (N_2164,N_1991,N_1767);
xnor U2165 (N_2165,N_1822,N_1812);
nor U2166 (N_2166,N_1757,N_1937);
xnor U2167 (N_2167,N_1951,N_1820);
and U2168 (N_2168,N_1896,N_1927);
xnor U2169 (N_2169,N_1891,N_1918);
xor U2170 (N_2170,N_1949,N_1951);
nor U2171 (N_2171,N_1953,N_1977);
nand U2172 (N_2172,N_1838,N_1765);
or U2173 (N_2173,N_1913,N_1872);
xor U2174 (N_2174,N_1752,N_1990);
nand U2175 (N_2175,N_1947,N_1879);
nor U2176 (N_2176,N_1894,N_1902);
nor U2177 (N_2177,N_1896,N_1976);
and U2178 (N_2178,N_1841,N_1940);
nand U2179 (N_2179,N_1904,N_1839);
nor U2180 (N_2180,N_1960,N_1925);
nand U2181 (N_2181,N_1785,N_1835);
xnor U2182 (N_2182,N_1855,N_1820);
and U2183 (N_2183,N_1814,N_1934);
and U2184 (N_2184,N_1795,N_1971);
and U2185 (N_2185,N_1875,N_1824);
xor U2186 (N_2186,N_1873,N_1917);
and U2187 (N_2187,N_1832,N_1935);
nand U2188 (N_2188,N_1808,N_1819);
nand U2189 (N_2189,N_1770,N_1896);
and U2190 (N_2190,N_1879,N_1761);
or U2191 (N_2191,N_1922,N_1832);
or U2192 (N_2192,N_1781,N_1951);
xor U2193 (N_2193,N_1820,N_1849);
or U2194 (N_2194,N_1889,N_1998);
or U2195 (N_2195,N_1753,N_1759);
xnor U2196 (N_2196,N_1939,N_1758);
nand U2197 (N_2197,N_1941,N_1759);
xnor U2198 (N_2198,N_1806,N_1881);
or U2199 (N_2199,N_1795,N_1828);
and U2200 (N_2200,N_1907,N_1960);
nand U2201 (N_2201,N_1773,N_1974);
nand U2202 (N_2202,N_1836,N_1996);
nor U2203 (N_2203,N_1970,N_1787);
xnor U2204 (N_2204,N_1882,N_1822);
and U2205 (N_2205,N_1986,N_1861);
nand U2206 (N_2206,N_1957,N_1762);
and U2207 (N_2207,N_1936,N_1934);
xnor U2208 (N_2208,N_1914,N_1945);
or U2209 (N_2209,N_1871,N_1877);
xnor U2210 (N_2210,N_1796,N_1776);
nor U2211 (N_2211,N_1754,N_1785);
nor U2212 (N_2212,N_1811,N_1899);
nand U2213 (N_2213,N_1906,N_1975);
nor U2214 (N_2214,N_1802,N_1943);
and U2215 (N_2215,N_1889,N_1841);
or U2216 (N_2216,N_1881,N_1882);
nand U2217 (N_2217,N_1789,N_1815);
nand U2218 (N_2218,N_1873,N_1931);
xnor U2219 (N_2219,N_1765,N_1820);
nor U2220 (N_2220,N_1785,N_1881);
and U2221 (N_2221,N_1894,N_1893);
xnor U2222 (N_2222,N_1831,N_1972);
xnor U2223 (N_2223,N_1825,N_1901);
or U2224 (N_2224,N_1931,N_1849);
or U2225 (N_2225,N_1983,N_1783);
and U2226 (N_2226,N_1998,N_1765);
nor U2227 (N_2227,N_1963,N_1944);
xor U2228 (N_2228,N_1896,N_1977);
or U2229 (N_2229,N_1871,N_1923);
xnor U2230 (N_2230,N_1901,N_1786);
nor U2231 (N_2231,N_1897,N_1919);
xor U2232 (N_2232,N_1754,N_1857);
nand U2233 (N_2233,N_1875,N_1971);
nand U2234 (N_2234,N_1976,N_1758);
nand U2235 (N_2235,N_1913,N_1758);
and U2236 (N_2236,N_1771,N_1767);
or U2237 (N_2237,N_1851,N_1955);
xnor U2238 (N_2238,N_1805,N_1827);
nor U2239 (N_2239,N_1990,N_1795);
nor U2240 (N_2240,N_1905,N_1877);
and U2241 (N_2241,N_1815,N_1891);
xnor U2242 (N_2242,N_1972,N_1905);
nor U2243 (N_2243,N_1808,N_1750);
and U2244 (N_2244,N_1962,N_1777);
and U2245 (N_2245,N_1984,N_1799);
and U2246 (N_2246,N_1807,N_1893);
and U2247 (N_2247,N_1952,N_1872);
nor U2248 (N_2248,N_1976,N_1768);
xnor U2249 (N_2249,N_1977,N_1787);
nand U2250 (N_2250,N_2230,N_2053);
and U2251 (N_2251,N_2194,N_2023);
or U2252 (N_2252,N_2037,N_2188);
nand U2253 (N_2253,N_2155,N_2096);
nand U2254 (N_2254,N_2137,N_2153);
xor U2255 (N_2255,N_2192,N_2185);
or U2256 (N_2256,N_2173,N_2209);
or U2257 (N_2257,N_2098,N_2134);
xnor U2258 (N_2258,N_2075,N_2228);
xnor U2259 (N_2259,N_2142,N_2011);
nand U2260 (N_2260,N_2108,N_2035);
nand U2261 (N_2261,N_2024,N_2206);
nor U2262 (N_2262,N_2112,N_2032);
or U2263 (N_2263,N_2141,N_2241);
nor U2264 (N_2264,N_2045,N_2130);
and U2265 (N_2265,N_2059,N_2195);
nor U2266 (N_2266,N_2086,N_2030);
nand U2267 (N_2267,N_2124,N_2058);
nand U2268 (N_2268,N_2100,N_2001);
or U2269 (N_2269,N_2160,N_2202);
xor U2270 (N_2270,N_2088,N_2213);
or U2271 (N_2271,N_2009,N_2216);
nor U2272 (N_2272,N_2013,N_2237);
nor U2273 (N_2273,N_2210,N_2022);
or U2274 (N_2274,N_2168,N_2179);
or U2275 (N_2275,N_2114,N_2070);
xor U2276 (N_2276,N_2018,N_2044);
xnor U2277 (N_2277,N_2065,N_2033);
xor U2278 (N_2278,N_2046,N_2187);
nor U2279 (N_2279,N_2060,N_2083);
nor U2280 (N_2280,N_2121,N_2102);
nand U2281 (N_2281,N_2157,N_2039);
nor U2282 (N_2282,N_2226,N_2158);
nand U2283 (N_2283,N_2150,N_2159);
xnor U2284 (N_2284,N_2235,N_2243);
and U2285 (N_2285,N_2196,N_2145);
nor U2286 (N_2286,N_2087,N_2239);
and U2287 (N_2287,N_2220,N_2020);
nor U2288 (N_2288,N_2232,N_2014);
xnor U2289 (N_2289,N_2077,N_2034);
xnor U2290 (N_2290,N_2127,N_2143);
and U2291 (N_2291,N_2218,N_2238);
xnor U2292 (N_2292,N_2122,N_2178);
or U2293 (N_2293,N_2105,N_2113);
xor U2294 (N_2294,N_2094,N_2040);
nand U2295 (N_2295,N_2169,N_2021);
nand U2296 (N_2296,N_2057,N_2138);
xor U2297 (N_2297,N_2166,N_2085);
nor U2298 (N_2298,N_2055,N_2162);
or U2299 (N_2299,N_2073,N_2131);
nor U2300 (N_2300,N_2092,N_2048);
nand U2301 (N_2301,N_2171,N_2147);
xnor U2302 (N_2302,N_2000,N_2031);
or U2303 (N_2303,N_2219,N_2082);
or U2304 (N_2304,N_2227,N_2008);
and U2305 (N_2305,N_2222,N_2090);
and U2306 (N_2306,N_2133,N_2116);
xor U2307 (N_2307,N_2139,N_2026);
and U2308 (N_2308,N_2152,N_2125);
or U2309 (N_2309,N_2107,N_2042);
nand U2310 (N_2310,N_2205,N_2076);
nand U2311 (N_2311,N_2007,N_2080);
or U2312 (N_2312,N_2191,N_2004);
or U2313 (N_2313,N_2144,N_2183);
or U2314 (N_2314,N_2248,N_2193);
xnor U2315 (N_2315,N_2167,N_2056);
xor U2316 (N_2316,N_2149,N_2089);
nor U2317 (N_2317,N_2099,N_2199);
nand U2318 (N_2318,N_2201,N_2074);
or U2319 (N_2319,N_2217,N_2180);
nand U2320 (N_2320,N_2204,N_2072);
nor U2321 (N_2321,N_2224,N_2208);
or U2322 (N_2322,N_2215,N_2132);
or U2323 (N_2323,N_2211,N_2236);
and U2324 (N_2324,N_2050,N_2063);
nor U2325 (N_2325,N_2244,N_2068);
nor U2326 (N_2326,N_2005,N_2154);
or U2327 (N_2327,N_2136,N_2229);
or U2328 (N_2328,N_2052,N_2069);
xor U2329 (N_2329,N_2110,N_2207);
nand U2330 (N_2330,N_2029,N_2214);
or U2331 (N_2331,N_2200,N_2084);
nand U2332 (N_2332,N_2181,N_2246);
xnor U2333 (N_2333,N_2109,N_2161);
nand U2334 (N_2334,N_2221,N_2120);
nor U2335 (N_2335,N_2064,N_2093);
and U2336 (N_2336,N_2016,N_2186);
and U2337 (N_2337,N_2182,N_2174);
nand U2338 (N_2338,N_2233,N_2189);
nand U2339 (N_2339,N_2197,N_2106);
nand U2340 (N_2340,N_2247,N_2165);
nand U2341 (N_2341,N_2066,N_2184);
nand U2342 (N_2342,N_2078,N_2041);
and U2343 (N_2343,N_2129,N_2027);
xor U2344 (N_2344,N_2101,N_2117);
xor U2345 (N_2345,N_2006,N_2097);
or U2346 (N_2346,N_2170,N_2119);
or U2347 (N_2347,N_2146,N_2234);
or U2348 (N_2348,N_2017,N_2225);
and U2349 (N_2349,N_2115,N_2126);
or U2350 (N_2350,N_2104,N_2240);
nor U2351 (N_2351,N_2148,N_2223);
nor U2352 (N_2352,N_2091,N_2028);
nor U2353 (N_2353,N_2123,N_2140);
nor U2354 (N_2354,N_2067,N_2015);
and U2355 (N_2355,N_2103,N_2062);
and U2356 (N_2356,N_2198,N_2212);
nand U2357 (N_2357,N_2012,N_2245);
nor U2358 (N_2358,N_2111,N_2151);
and U2359 (N_2359,N_2061,N_2051);
nand U2360 (N_2360,N_2025,N_2054);
and U2361 (N_2361,N_2043,N_2249);
nor U2362 (N_2362,N_2190,N_2242);
or U2363 (N_2363,N_2156,N_2036);
nor U2364 (N_2364,N_2164,N_2079);
and U2365 (N_2365,N_2135,N_2038);
nand U2366 (N_2366,N_2003,N_2002);
and U2367 (N_2367,N_2128,N_2177);
or U2368 (N_2368,N_2071,N_2118);
or U2369 (N_2369,N_2047,N_2019);
and U2370 (N_2370,N_2163,N_2081);
and U2371 (N_2371,N_2172,N_2203);
or U2372 (N_2372,N_2095,N_2175);
nand U2373 (N_2373,N_2049,N_2010);
or U2374 (N_2374,N_2176,N_2231);
nor U2375 (N_2375,N_2032,N_2249);
and U2376 (N_2376,N_2203,N_2023);
and U2377 (N_2377,N_2034,N_2161);
and U2378 (N_2378,N_2110,N_2010);
or U2379 (N_2379,N_2035,N_2185);
nor U2380 (N_2380,N_2001,N_2232);
xor U2381 (N_2381,N_2153,N_2003);
and U2382 (N_2382,N_2198,N_2209);
nand U2383 (N_2383,N_2178,N_2071);
and U2384 (N_2384,N_2020,N_2091);
or U2385 (N_2385,N_2115,N_2200);
and U2386 (N_2386,N_2037,N_2198);
xnor U2387 (N_2387,N_2172,N_2080);
or U2388 (N_2388,N_2243,N_2035);
and U2389 (N_2389,N_2003,N_2065);
nand U2390 (N_2390,N_2198,N_2061);
xor U2391 (N_2391,N_2222,N_2225);
or U2392 (N_2392,N_2190,N_2173);
xor U2393 (N_2393,N_2204,N_2154);
xnor U2394 (N_2394,N_2097,N_2130);
and U2395 (N_2395,N_2248,N_2221);
nand U2396 (N_2396,N_2244,N_2080);
nor U2397 (N_2397,N_2222,N_2035);
nor U2398 (N_2398,N_2162,N_2136);
xnor U2399 (N_2399,N_2230,N_2214);
nand U2400 (N_2400,N_2223,N_2034);
xor U2401 (N_2401,N_2217,N_2189);
or U2402 (N_2402,N_2129,N_2069);
or U2403 (N_2403,N_2228,N_2068);
nand U2404 (N_2404,N_2080,N_2069);
or U2405 (N_2405,N_2200,N_2089);
xnor U2406 (N_2406,N_2143,N_2028);
and U2407 (N_2407,N_2196,N_2007);
xnor U2408 (N_2408,N_2061,N_2003);
and U2409 (N_2409,N_2004,N_2136);
xnor U2410 (N_2410,N_2185,N_2015);
nor U2411 (N_2411,N_2188,N_2173);
nand U2412 (N_2412,N_2095,N_2238);
nor U2413 (N_2413,N_2010,N_2218);
or U2414 (N_2414,N_2082,N_2148);
and U2415 (N_2415,N_2153,N_2204);
nand U2416 (N_2416,N_2152,N_2249);
xor U2417 (N_2417,N_2112,N_2104);
nand U2418 (N_2418,N_2120,N_2147);
nor U2419 (N_2419,N_2078,N_2077);
or U2420 (N_2420,N_2114,N_2101);
nand U2421 (N_2421,N_2203,N_2187);
and U2422 (N_2422,N_2145,N_2143);
nand U2423 (N_2423,N_2109,N_2025);
xnor U2424 (N_2424,N_2157,N_2044);
xor U2425 (N_2425,N_2032,N_2140);
nand U2426 (N_2426,N_2008,N_2121);
and U2427 (N_2427,N_2232,N_2150);
xor U2428 (N_2428,N_2194,N_2088);
or U2429 (N_2429,N_2095,N_2096);
xor U2430 (N_2430,N_2027,N_2139);
or U2431 (N_2431,N_2102,N_2026);
xnor U2432 (N_2432,N_2062,N_2065);
or U2433 (N_2433,N_2084,N_2189);
and U2434 (N_2434,N_2128,N_2105);
and U2435 (N_2435,N_2087,N_2125);
or U2436 (N_2436,N_2132,N_2153);
nor U2437 (N_2437,N_2038,N_2115);
nor U2438 (N_2438,N_2017,N_2175);
nor U2439 (N_2439,N_2084,N_2031);
nor U2440 (N_2440,N_2217,N_2218);
and U2441 (N_2441,N_2166,N_2051);
xnor U2442 (N_2442,N_2026,N_2073);
nor U2443 (N_2443,N_2033,N_2225);
or U2444 (N_2444,N_2089,N_2132);
nor U2445 (N_2445,N_2044,N_2230);
xor U2446 (N_2446,N_2020,N_2204);
nor U2447 (N_2447,N_2223,N_2210);
or U2448 (N_2448,N_2034,N_2217);
nor U2449 (N_2449,N_2197,N_2110);
xnor U2450 (N_2450,N_2189,N_2071);
and U2451 (N_2451,N_2099,N_2047);
or U2452 (N_2452,N_2179,N_2012);
or U2453 (N_2453,N_2115,N_2119);
xnor U2454 (N_2454,N_2047,N_2133);
nand U2455 (N_2455,N_2175,N_2249);
nor U2456 (N_2456,N_2063,N_2236);
nand U2457 (N_2457,N_2158,N_2055);
or U2458 (N_2458,N_2116,N_2056);
or U2459 (N_2459,N_2062,N_2023);
nor U2460 (N_2460,N_2122,N_2166);
nand U2461 (N_2461,N_2015,N_2179);
nand U2462 (N_2462,N_2020,N_2123);
nand U2463 (N_2463,N_2034,N_2130);
nand U2464 (N_2464,N_2239,N_2053);
nand U2465 (N_2465,N_2181,N_2170);
and U2466 (N_2466,N_2093,N_2071);
or U2467 (N_2467,N_2003,N_2125);
xnor U2468 (N_2468,N_2168,N_2094);
nand U2469 (N_2469,N_2206,N_2234);
or U2470 (N_2470,N_2082,N_2232);
xnor U2471 (N_2471,N_2024,N_2118);
or U2472 (N_2472,N_2052,N_2115);
xnor U2473 (N_2473,N_2166,N_2105);
nor U2474 (N_2474,N_2070,N_2220);
xor U2475 (N_2475,N_2056,N_2145);
xnor U2476 (N_2476,N_2163,N_2138);
nor U2477 (N_2477,N_2225,N_2002);
and U2478 (N_2478,N_2104,N_2219);
and U2479 (N_2479,N_2226,N_2034);
nand U2480 (N_2480,N_2226,N_2016);
or U2481 (N_2481,N_2004,N_2058);
and U2482 (N_2482,N_2081,N_2177);
xnor U2483 (N_2483,N_2177,N_2217);
or U2484 (N_2484,N_2072,N_2216);
nand U2485 (N_2485,N_2144,N_2169);
or U2486 (N_2486,N_2061,N_2110);
or U2487 (N_2487,N_2079,N_2163);
or U2488 (N_2488,N_2231,N_2055);
and U2489 (N_2489,N_2117,N_2175);
nor U2490 (N_2490,N_2108,N_2212);
nand U2491 (N_2491,N_2240,N_2089);
or U2492 (N_2492,N_2125,N_2111);
nand U2493 (N_2493,N_2184,N_2131);
nor U2494 (N_2494,N_2086,N_2110);
nand U2495 (N_2495,N_2134,N_2151);
xor U2496 (N_2496,N_2097,N_2051);
and U2497 (N_2497,N_2135,N_2149);
nor U2498 (N_2498,N_2119,N_2201);
nand U2499 (N_2499,N_2041,N_2239);
nor U2500 (N_2500,N_2419,N_2433);
nor U2501 (N_2501,N_2448,N_2375);
nand U2502 (N_2502,N_2435,N_2454);
or U2503 (N_2503,N_2374,N_2415);
nor U2504 (N_2504,N_2377,N_2278);
and U2505 (N_2505,N_2310,N_2450);
nor U2506 (N_2506,N_2395,N_2444);
xor U2507 (N_2507,N_2460,N_2353);
xor U2508 (N_2508,N_2295,N_2269);
nand U2509 (N_2509,N_2484,N_2432);
and U2510 (N_2510,N_2262,N_2277);
nor U2511 (N_2511,N_2496,N_2421);
nor U2512 (N_2512,N_2464,N_2322);
or U2513 (N_2513,N_2253,N_2473);
and U2514 (N_2514,N_2313,N_2390);
nor U2515 (N_2515,N_2274,N_2469);
and U2516 (N_2516,N_2426,N_2294);
or U2517 (N_2517,N_2458,N_2495);
and U2518 (N_2518,N_2298,N_2346);
xnor U2519 (N_2519,N_2376,N_2416);
nand U2520 (N_2520,N_2327,N_2337);
nand U2521 (N_2521,N_2479,N_2288);
and U2522 (N_2522,N_2487,N_2431);
nor U2523 (N_2523,N_2396,N_2341);
xnor U2524 (N_2524,N_2411,N_2279);
or U2525 (N_2525,N_2489,N_2342);
nand U2526 (N_2526,N_2378,N_2345);
nor U2527 (N_2527,N_2339,N_2493);
nor U2528 (N_2528,N_2417,N_2398);
nand U2529 (N_2529,N_2358,N_2440);
nand U2530 (N_2530,N_2455,N_2486);
and U2531 (N_2531,N_2424,N_2488);
xnor U2532 (N_2532,N_2318,N_2429);
nor U2533 (N_2533,N_2474,N_2355);
nand U2534 (N_2534,N_2280,N_2323);
or U2535 (N_2535,N_2463,N_2314);
or U2536 (N_2536,N_2284,N_2401);
and U2537 (N_2537,N_2420,N_2308);
nand U2538 (N_2538,N_2364,N_2393);
and U2539 (N_2539,N_2273,N_2268);
nand U2540 (N_2540,N_2361,N_2430);
and U2541 (N_2541,N_2412,N_2438);
xor U2542 (N_2542,N_2498,N_2252);
nor U2543 (N_2543,N_2409,N_2250);
nor U2544 (N_2544,N_2351,N_2385);
and U2545 (N_2545,N_2256,N_2293);
and U2546 (N_2546,N_2399,N_2325);
nand U2547 (N_2547,N_2296,N_2297);
xnor U2548 (N_2548,N_2388,N_2367);
nand U2549 (N_2549,N_2483,N_2497);
nand U2550 (N_2550,N_2261,N_2371);
nor U2551 (N_2551,N_2373,N_2413);
xor U2552 (N_2552,N_2286,N_2457);
nand U2553 (N_2553,N_2348,N_2266);
or U2554 (N_2554,N_2456,N_2386);
nor U2555 (N_2555,N_2477,N_2272);
or U2556 (N_2556,N_2316,N_2283);
xor U2557 (N_2557,N_2303,N_2369);
and U2558 (N_2558,N_2391,N_2291);
xnor U2559 (N_2559,N_2263,N_2452);
nand U2560 (N_2560,N_2360,N_2368);
or U2561 (N_2561,N_2402,N_2257);
nor U2562 (N_2562,N_2311,N_2380);
and U2563 (N_2563,N_2405,N_2447);
nor U2564 (N_2564,N_2422,N_2251);
xor U2565 (N_2565,N_2267,N_2289);
and U2566 (N_2566,N_2326,N_2466);
nand U2567 (N_2567,N_2407,N_2425);
and U2568 (N_2568,N_2255,N_2471);
or U2569 (N_2569,N_2356,N_2389);
nand U2570 (N_2570,N_2344,N_2475);
nand U2571 (N_2571,N_2387,N_2306);
or U2572 (N_2572,N_2307,N_2352);
nor U2573 (N_2573,N_2292,N_2499);
xor U2574 (N_2574,N_2270,N_2328);
xnor U2575 (N_2575,N_2418,N_2449);
nand U2576 (N_2576,N_2258,N_2476);
and U2577 (N_2577,N_2404,N_2397);
nand U2578 (N_2578,N_2357,N_2319);
and U2579 (N_2579,N_2480,N_2461);
xnor U2580 (N_2580,N_2332,N_2372);
and U2581 (N_2581,N_2427,N_2485);
nand U2582 (N_2582,N_2264,N_2446);
nand U2583 (N_2583,N_2467,N_2414);
or U2584 (N_2584,N_2442,N_2453);
and U2585 (N_2585,N_2315,N_2276);
or U2586 (N_2586,N_2470,N_2271);
xor U2587 (N_2587,N_2320,N_2305);
and U2588 (N_2588,N_2441,N_2410);
xor U2589 (N_2589,N_2365,N_2406);
and U2590 (N_2590,N_2363,N_2312);
xnor U2591 (N_2591,N_2321,N_2381);
nor U2592 (N_2592,N_2451,N_2490);
nor U2593 (N_2593,N_2439,N_2350);
nand U2594 (N_2594,N_2478,N_2354);
nand U2595 (N_2595,N_2340,N_2382);
nor U2596 (N_2596,N_2434,N_2347);
xor U2597 (N_2597,N_2423,N_2468);
and U2598 (N_2598,N_2366,N_2285);
nor U2599 (N_2599,N_2260,N_2329);
xor U2600 (N_2600,N_2254,N_2334);
and U2601 (N_2601,N_2259,N_2301);
or U2602 (N_2602,N_2392,N_2445);
or U2603 (N_2603,N_2465,N_2403);
or U2604 (N_2604,N_2383,N_2394);
nor U2605 (N_2605,N_2370,N_2482);
or U2606 (N_2606,N_2330,N_2491);
xor U2607 (N_2607,N_2436,N_2384);
or U2608 (N_2608,N_2408,N_2324);
or U2609 (N_2609,N_2309,N_2331);
nor U2610 (N_2610,N_2317,N_2299);
nand U2611 (N_2611,N_2349,N_2265);
or U2612 (N_2612,N_2300,N_2290);
xor U2613 (N_2613,N_2362,N_2275);
nand U2614 (N_2614,N_2437,N_2481);
nand U2615 (N_2615,N_2379,N_2304);
nand U2616 (N_2616,N_2302,N_2494);
nor U2617 (N_2617,N_2282,N_2336);
and U2618 (N_2618,N_2492,N_2462);
xnor U2619 (N_2619,N_2459,N_2343);
nand U2620 (N_2620,N_2472,N_2335);
nand U2621 (N_2621,N_2281,N_2428);
nand U2622 (N_2622,N_2333,N_2359);
and U2623 (N_2623,N_2443,N_2287);
or U2624 (N_2624,N_2338,N_2400);
and U2625 (N_2625,N_2496,N_2440);
or U2626 (N_2626,N_2452,N_2391);
nand U2627 (N_2627,N_2489,N_2251);
nor U2628 (N_2628,N_2391,N_2499);
xnor U2629 (N_2629,N_2291,N_2396);
xor U2630 (N_2630,N_2412,N_2354);
nand U2631 (N_2631,N_2328,N_2291);
xnor U2632 (N_2632,N_2305,N_2435);
xnor U2633 (N_2633,N_2361,N_2350);
or U2634 (N_2634,N_2414,N_2284);
and U2635 (N_2635,N_2264,N_2360);
nand U2636 (N_2636,N_2397,N_2337);
or U2637 (N_2637,N_2415,N_2364);
and U2638 (N_2638,N_2424,N_2453);
xor U2639 (N_2639,N_2300,N_2400);
nand U2640 (N_2640,N_2363,N_2292);
xor U2641 (N_2641,N_2353,N_2336);
nand U2642 (N_2642,N_2474,N_2254);
xor U2643 (N_2643,N_2357,N_2407);
xor U2644 (N_2644,N_2437,N_2335);
nor U2645 (N_2645,N_2497,N_2250);
and U2646 (N_2646,N_2492,N_2292);
nand U2647 (N_2647,N_2277,N_2327);
nor U2648 (N_2648,N_2275,N_2314);
xor U2649 (N_2649,N_2417,N_2426);
nand U2650 (N_2650,N_2491,N_2362);
or U2651 (N_2651,N_2395,N_2462);
nor U2652 (N_2652,N_2256,N_2365);
or U2653 (N_2653,N_2333,N_2438);
and U2654 (N_2654,N_2416,N_2283);
xnor U2655 (N_2655,N_2296,N_2399);
nand U2656 (N_2656,N_2419,N_2361);
or U2657 (N_2657,N_2431,N_2259);
xnor U2658 (N_2658,N_2265,N_2465);
and U2659 (N_2659,N_2349,N_2336);
nor U2660 (N_2660,N_2420,N_2335);
and U2661 (N_2661,N_2360,N_2269);
nand U2662 (N_2662,N_2484,N_2330);
xor U2663 (N_2663,N_2486,N_2375);
nor U2664 (N_2664,N_2317,N_2414);
or U2665 (N_2665,N_2455,N_2258);
xor U2666 (N_2666,N_2274,N_2314);
or U2667 (N_2667,N_2328,N_2356);
xnor U2668 (N_2668,N_2372,N_2305);
nand U2669 (N_2669,N_2446,N_2436);
and U2670 (N_2670,N_2484,N_2362);
or U2671 (N_2671,N_2363,N_2459);
and U2672 (N_2672,N_2368,N_2307);
xnor U2673 (N_2673,N_2457,N_2384);
xor U2674 (N_2674,N_2395,N_2355);
or U2675 (N_2675,N_2443,N_2271);
nand U2676 (N_2676,N_2319,N_2370);
xor U2677 (N_2677,N_2443,N_2353);
nor U2678 (N_2678,N_2470,N_2286);
and U2679 (N_2679,N_2497,N_2307);
nor U2680 (N_2680,N_2476,N_2267);
or U2681 (N_2681,N_2302,N_2448);
nand U2682 (N_2682,N_2377,N_2400);
or U2683 (N_2683,N_2347,N_2308);
or U2684 (N_2684,N_2253,N_2376);
xor U2685 (N_2685,N_2474,N_2354);
xor U2686 (N_2686,N_2423,N_2264);
and U2687 (N_2687,N_2337,N_2444);
and U2688 (N_2688,N_2412,N_2358);
and U2689 (N_2689,N_2490,N_2274);
nand U2690 (N_2690,N_2440,N_2371);
and U2691 (N_2691,N_2420,N_2376);
and U2692 (N_2692,N_2496,N_2360);
nor U2693 (N_2693,N_2485,N_2340);
and U2694 (N_2694,N_2368,N_2337);
nand U2695 (N_2695,N_2285,N_2452);
nand U2696 (N_2696,N_2316,N_2265);
and U2697 (N_2697,N_2271,N_2403);
and U2698 (N_2698,N_2295,N_2376);
or U2699 (N_2699,N_2466,N_2480);
nor U2700 (N_2700,N_2450,N_2496);
nor U2701 (N_2701,N_2267,N_2388);
nand U2702 (N_2702,N_2270,N_2269);
or U2703 (N_2703,N_2388,N_2455);
nand U2704 (N_2704,N_2382,N_2355);
nor U2705 (N_2705,N_2397,N_2385);
or U2706 (N_2706,N_2489,N_2316);
nor U2707 (N_2707,N_2267,N_2262);
nand U2708 (N_2708,N_2442,N_2318);
xnor U2709 (N_2709,N_2289,N_2330);
nand U2710 (N_2710,N_2411,N_2300);
or U2711 (N_2711,N_2308,N_2440);
xnor U2712 (N_2712,N_2423,N_2479);
xnor U2713 (N_2713,N_2320,N_2389);
xnor U2714 (N_2714,N_2323,N_2328);
or U2715 (N_2715,N_2375,N_2379);
or U2716 (N_2716,N_2324,N_2253);
and U2717 (N_2717,N_2397,N_2333);
nor U2718 (N_2718,N_2424,N_2489);
nand U2719 (N_2719,N_2336,N_2397);
nor U2720 (N_2720,N_2345,N_2319);
and U2721 (N_2721,N_2450,N_2431);
nand U2722 (N_2722,N_2439,N_2440);
xor U2723 (N_2723,N_2443,N_2407);
and U2724 (N_2724,N_2287,N_2312);
xor U2725 (N_2725,N_2391,N_2386);
xor U2726 (N_2726,N_2336,N_2322);
and U2727 (N_2727,N_2416,N_2335);
xnor U2728 (N_2728,N_2416,N_2334);
nor U2729 (N_2729,N_2262,N_2459);
and U2730 (N_2730,N_2491,N_2481);
nand U2731 (N_2731,N_2355,N_2414);
or U2732 (N_2732,N_2486,N_2389);
nand U2733 (N_2733,N_2389,N_2394);
and U2734 (N_2734,N_2328,N_2494);
and U2735 (N_2735,N_2343,N_2326);
xor U2736 (N_2736,N_2274,N_2457);
nor U2737 (N_2737,N_2403,N_2461);
nor U2738 (N_2738,N_2340,N_2477);
nor U2739 (N_2739,N_2472,N_2337);
and U2740 (N_2740,N_2404,N_2278);
xor U2741 (N_2741,N_2252,N_2383);
nand U2742 (N_2742,N_2456,N_2359);
or U2743 (N_2743,N_2387,N_2325);
and U2744 (N_2744,N_2296,N_2430);
and U2745 (N_2745,N_2334,N_2310);
or U2746 (N_2746,N_2259,N_2364);
nand U2747 (N_2747,N_2334,N_2497);
nand U2748 (N_2748,N_2290,N_2354);
nand U2749 (N_2749,N_2311,N_2406);
nor U2750 (N_2750,N_2575,N_2737);
and U2751 (N_2751,N_2606,N_2603);
and U2752 (N_2752,N_2545,N_2646);
xor U2753 (N_2753,N_2726,N_2691);
nand U2754 (N_2754,N_2658,N_2604);
nand U2755 (N_2755,N_2611,N_2563);
nand U2756 (N_2756,N_2684,N_2679);
or U2757 (N_2757,N_2715,N_2741);
xor U2758 (N_2758,N_2521,N_2718);
nor U2759 (N_2759,N_2720,N_2742);
and U2760 (N_2760,N_2642,N_2651);
nor U2761 (N_2761,N_2697,N_2552);
xor U2762 (N_2762,N_2567,N_2556);
nand U2763 (N_2763,N_2629,N_2695);
xor U2764 (N_2764,N_2728,N_2525);
xnor U2765 (N_2765,N_2590,N_2522);
nor U2766 (N_2766,N_2625,N_2543);
nor U2767 (N_2767,N_2712,N_2580);
nand U2768 (N_2768,N_2537,N_2663);
and U2769 (N_2769,N_2595,N_2612);
nand U2770 (N_2770,N_2656,N_2548);
or U2771 (N_2771,N_2535,N_2530);
nand U2772 (N_2772,N_2633,N_2719);
or U2773 (N_2773,N_2512,N_2626);
nor U2774 (N_2774,N_2599,N_2621);
or U2775 (N_2775,N_2650,N_2637);
xnor U2776 (N_2776,N_2634,N_2581);
xor U2777 (N_2777,N_2510,N_2609);
nand U2778 (N_2778,N_2502,N_2562);
nand U2779 (N_2779,N_2618,N_2692);
and U2780 (N_2780,N_2677,N_2564);
and U2781 (N_2781,N_2733,N_2665);
or U2782 (N_2782,N_2685,N_2613);
or U2783 (N_2783,N_2743,N_2531);
xnor U2784 (N_2784,N_2542,N_2683);
nor U2785 (N_2785,N_2705,N_2717);
nor U2786 (N_2786,N_2511,N_2681);
xnor U2787 (N_2787,N_2631,N_2635);
nor U2788 (N_2788,N_2503,N_2676);
and U2789 (N_2789,N_2524,N_2598);
and U2790 (N_2790,N_2583,N_2547);
or U2791 (N_2791,N_2585,N_2690);
nand U2792 (N_2792,N_2630,N_2648);
nor U2793 (N_2793,N_2641,N_2624);
or U2794 (N_2794,N_2584,N_2528);
xnor U2795 (N_2795,N_2680,N_2571);
or U2796 (N_2796,N_2724,N_2614);
nand U2797 (N_2797,N_2597,N_2664);
and U2798 (N_2798,N_2509,N_2600);
xor U2799 (N_2799,N_2660,N_2610);
xor U2800 (N_2800,N_2501,N_2688);
nor U2801 (N_2801,N_2565,N_2632);
or U2802 (N_2802,N_2574,N_2643);
nor U2803 (N_2803,N_2572,N_2652);
xnor U2804 (N_2804,N_2670,N_2588);
and U2805 (N_2805,N_2639,N_2558);
nor U2806 (N_2806,N_2744,N_2708);
or U2807 (N_2807,N_2533,N_2532);
nor U2808 (N_2808,N_2601,N_2559);
xnor U2809 (N_2809,N_2745,N_2586);
nor U2810 (N_2810,N_2566,N_2505);
and U2811 (N_2811,N_2645,N_2546);
xor U2812 (N_2812,N_2539,N_2730);
nand U2813 (N_2813,N_2594,N_2678);
or U2814 (N_2814,N_2667,N_2638);
and U2815 (N_2815,N_2616,N_2627);
and U2816 (N_2816,N_2661,N_2689);
nor U2817 (N_2817,N_2534,N_2582);
nor U2818 (N_2818,N_2554,N_2589);
or U2819 (N_2819,N_2507,N_2504);
and U2820 (N_2820,N_2526,N_2727);
xnor U2821 (N_2821,N_2655,N_2657);
xnor U2822 (N_2822,N_2732,N_2666);
xnor U2823 (N_2823,N_2605,N_2702);
nand U2824 (N_2824,N_2662,N_2555);
or U2825 (N_2825,N_2615,N_2654);
or U2826 (N_2826,N_2696,N_2687);
and U2827 (N_2827,N_2576,N_2569);
nand U2828 (N_2828,N_2517,N_2518);
or U2829 (N_2829,N_2593,N_2536);
or U2830 (N_2830,N_2570,N_2617);
or U2831 (N_2831,N_2602,N_2608);
nor U2832 (N_2832,N_2710,N_2706);
nand U2833 (N_2833,N_2711,N_2520);
nor U2834 (N_2834,N_2746,N_2722);
nand U2835 (N_2835,N_2527,N_2682);
and U2836 (N_2836,N_2740,N_2577);
nand U2837 (N_2837,N_2694,N_2523);
nand U2838 (N_2838,N_2514,N_2591);
nand U2839 (N_2839,N_2649,N_2748);
and U2840 (N_2840,N_2636,N_2515);
xor U2841 (N_2841,N_2731,N_2736);
nor U2842 (N_2842,N_2653,N_2701);
nor U2843 (N_2843,N_2723,N_2749);
xnor U2844 (N_2844,N_2699,N_2716);
nor U2845 (N_2845,N_2561,N_2620);
nor U2846 (N_2846,N_2587,N_2541);
or U2847 (N_2847,N_2622,N_2700);
nand U2848 (N_2848,N_2686,N_2669);
and U2849 (N_2849,N_2675,N_2714);
xnor U2850 (N_2850,N_2573,N_2516);
and U2851 (N_2851,N_2519,N_2738);
nand U2852 (N_2852,N_2729,N_2713);
xnor U2853 (N_2853,N_2578,N_2747);
or U2854 (N_2854,N_2659,N_2508);
nor U2855 (N_2855,N_2628,N_2607);
nand U2856 (N_2856,N_2557,N_2513);
nand U2857 (N_2857,N_2500,N_2674);
and U2858 (N_2858,N_2647,N_2703);
xor U2859 (N_2859,N_2553,N_2693);
nand U2860 (N_2860,N_2721,N_2540);
and U2861 (N_2861,N_2709,N_2672);
nand U2862 (N_2862,N_2550,N_2725);
nor U2863 (N_2863,N_2551,N_2592);
nand U2864 (N_2864,N_2619,N_2734);
xor U2865 (N_2865,N_2538,N_2549);
nand U2866 (N_2866,N_2529,N_2596);
xor U2867 (N_2867,N_2506,N_2671);
nor U2868 (N_2868,N_2579,N_2673);
nor U2869 (N_2869,N_2623,N_2560);
and U2870 (N_2870,N_2568,N_2735);
nor U2871 (N_2871,N_2644,N_2544);
or U2872 (N_2872,N_2668,N_2707);
xor U2873 (N_2873,N_2640,N_2739);
nand U2874 (N_2874,N_2698,N_2704);
xnor U2875 (N_2875,N_2720,N_2738);
or U2876 (N_2876,N_2619,N_2581);
and U2877 (N_2877,N_2633,N_2655);
and U2878 (N_2878,N_2571,N_2690);
or U2879 (N_2879,N_2550,N_2579);
nor U2880 (N_2880,N_2679,N_2718);
or U2881 (N_2881,N_2548,N_2558);
or U2882 (N_2882,N_2638,N_2561);
xnor U2883 (N_2883,N_2560,N_2708);
nand U2884 (N_2884,N_2722,N_2613);
nand U2885 (N_2885,N_2579,N_2676);
xor U2886 (N_2886,N_2695,N_2591);
xor U2887 (N_2887,N_2633,N_2722);
and U2888 (N_2888,N_2624,N_2541);
or U2889 (N_2889,N_2643,N_2650);
nor U2890 (N_2890,N_2619,N_2741);
nand U2891 (N_2891,N_2548,N_2702);
or U2892 (N_2892,N_2573,N_2568);
xor U2893 (N_2893,N_2675,N_2680);
xor U2894 (N_2894,N_2601,N_2552);
nor U2895 (N_2895,N_2707,N_2591);
nand U2896 (N_2896,N_2539,N_2587);
nor U2897 (N_2897,N_2742,N_2737);
nor U2898 (N_2898,N_2582,N_2632);
nand U2899 (N_2899,N_2595,N_2727);
nor U2900 (N_2900,N_2510,N_2584);
nor U2901 (N_2901,N_2749,N_2581);
or U2902 (N_2902,N_2552,N_2600);
or U2903 (N_2903,N_2639,N_2601);
xnor U2904 (N_2904,N_2690,N_2520);
xnor U2905 (N_2905,N_2557,N_2590);
xor U2906 (N_2906,N_2529,N_2711);
and U2907 (N_2907,N_2649,N_2545);
or U2908 (N_2908,N_2507,N_2546);
xnor U2909 (N_2909,N_2679,N_2632);
nor U2910 (N_2910,N_2729,N_2531);
and U2911 (N_2911,N_2561,N_2502);
nor U2912 (N_2912,N_2692,N_2510);
nand U2913 (N_2913,N_2593,N_2641);
and U2914 (N_2914,N_2553,N_2522);
nor U2915 (N_2915,N_2545,N_2510);
nand U2916 (N_2916,N_2558,N_2570);
and U2917 (N_2917,N_2652,N_2701);
and U2918 (N_2918,N_2531,N_2705);
and U2919 (N_2919,N_2617,N_2502);
nor U2920 (N_2920,N_2746,N_2551);
and U2921 (N_2921,N_2689,N_2645);
nor U2922 (N_2922,N_2669,N_2620);
or U2923 (N_2923,N_2565,N_2722);
nand U2924 (N_2924,N_2548,N_2664);
nand U2925 (N_2925,N_2590,N_2583);
nor U2926 (N_2926,N_2587,N_2651);
nand U2927 (N_2927,N_2589,N_2582);
and U2928 (N_2928,N_2732,N_2702);
nor U2929 (N_2929,N_2555,N_2649);
xnor U2930 (N_2930,N_2659,N_2515);
xnor U2931 (N_2931,N_2508,N_2730);
nand U2932 (N_2932,N_2520,N_2648);
and U2933 (N_2933,N_2548,N_2711);
nand U2934 (N_2934,N_2662,N_2745);
or U2935 (N_2935,N_2558,N_2624);
and U2936 (N_2936,N_2600,N_2711);
nand U2937 (N_2937,N_2696,N_2500);
and U2938 (N_2938,N_2736,N_2561);
xnor U2939 (N_2939,N_2658,N_2659);
nand U2940 (N_2940,N_2556,N_2505);
nor U2941 (N_2941,N_2578,N_2506);
xnor U2942 (N_2942,N_2731,N_2672);
nor U2943 (N_2943,N_2627,N_2623);
nand U2944 (N_2944,N_2668,N_2685);
and U2945 (N_2945,N_2735,N_2546);
or U2946 (N_2946,N_2719,N_2552);
nand U2947 (N_2947,N_2726,N_2540);
nor U2948 (N_2948,N_2585,N_2691);
or U2949 (N_2949,N_2658,N_2687);
xnor U2950 (N_2950,N_2711,N_2608);
nand U2951 (N_2951,N_2743,N_2707);
xnor U2952 (N_2952,N_2555,N_2604);
and U2953 (N_2953,N_2630,N_2507);
or U2954 (N_2954,N_2681,N_2524);
nand U2955 (N_2955,N_2673,N_2728);
and U2956 (N_2956,N_2510,N_2575);
nand U2957 (N_2957,N_2663,N_2710);
xnor U2958 (N_2958,N_2655,N_2587);
nor U2959 (N_2959,N_2603,N_2605);
and U2960 (N_2960,N_2585,N_2728);
nand U2961 (N_2961,N_2512,N_2584);
nand U2962 (N_2962,N_2741,N_2505);
or U2963 (N_2963,N_2748,N_2606);
xor U2964 (N_2964,N_2521,N_2738);
nand U2965 (N_2965,N_2651,N_2552);
xnor U2966 (N_2966,N_2671,N_2526);
and U2967 (N_2967,N_2647,N_2564);
nor U2968 (N_2968,N_2540,N_2697);
nand U2969 (N_2969,N_2599,N_2685);
or U2970 (N_2970,N_2503,N_2537);
or U2971 (N_2971,N_2590,N_2637);
or U2972 (N_2972,N_2676,N_2663);
and U2973 (N_2973,N_2670,N_2707);
or U2974 (N_2974,N_2510,N_2681);
xor U2975 (N_2975,N_2726,N_2734);
and U2976 (N_2976,N_2579,N_2556);
or U2977 (N_2977,N_2705,N_2592);
and U2978 (N_2978,N_2549,N_2575);
xnor U2979 (N_2979,N_2561,N_2586);
xor U2980 (N_2980,N_2669,N_2690);
and U2981 (N_2981,N_2747,N_2541);
and U2982 (N_2982,N_2704,N_2514);
nor U2983 (N_2983,N_2749,N_2747);
and U2984 (N_2984,N_2522,N_2614);
nor U2985 (N_2985,N_2672,N_2742);
nand U2986 (N_2986,N_2569,N_2719);
nor U2987 (N_2987,N_2748,N_2666);
and U2988 (N_2988,N_2642,N_2604);
nand U2989 (N_2989,N_2737,N_2649);
nor U2990 (N_2990,N_2527,N_2619);
and U2991 (N_2991,N_2519,N_2656);
nand U2992 (N_2992,N_2742,N_2704);
nand U2993 (N_2993,N_2505,N_2519);
nor U2994 (N_2994,N_2524,N_2544);
xnor U2995 (N_2995,N_2578,N_2696);
xnor U2996 (N_2996,N_2542,N_2584);
and U2997 (N_2997,N_2720,N_2577);
and U2998 (N_2998,N_2549,N_2716);
xor U2999 (N_2999,N_2535,N_2617);
xnor U3000 (N_3000,N_2994,N_2833);
or U3001 (N_3001,N_2979,N_2772);
nor U3002 (N_3002,N_2767,N_2977);
and U3003 (N_3003,N_2809,N_2814);
and U3004 (N_3004,N_2806,N_2982);
or U3005 (N_3005,N_2945,N_2910);
xor U3006 (N_3006,N_2842,N_2856);
xnor U3007 (N_3007,N_2830,N_2754);
and U3008 (N_3008,N_2789,N_2850);
nor U3009 (N_3009,N_2980,N_2997);
and U3010 (N_3010,N_2916,N_2998);
xor U3011 (N_3011,N_2836,N_2808);
xor U3012 (N_3012,N_2807,N_2971);
and U3013 (N_3013,N_2987,N_2949);
and U3014 (N_3014,N_2882,N_2904);
or U3015 (N_3015,N_2775,N_2995);
nor U3016 (N_3016,N_2800,N_2975);
nand U3017 (N_3017,N_2838,N_2824);
or U3018 (N_3018,N_2947,N_2892);
and U3019 (N_3019,N_2897,N_2769);
or U3020 (N_3020,N_2907,N_2797);
nand U3021 (N_3021,N_2919,N_2844);
nand U3022 (N_3022,N_2763,N_2821);
or U3023 (N_3023,N_2954,N_2768);
nor U3024 (N_3024,N_2946,N_2942);
or U3025 (N_3025,N_2864,N_2837);
and U3026 (N_3026,N_2857,N_2788);
and U3027 (N_3027,N_2758,N_2793);
or U3028 (N_3028,N_2798,N_2981);
nor U3029 (N_3029,N_2827,N_2792);
and U3030 (N_3030,N_2866,N_2868);
or U3031 (N_3031,N_2887,N_2978);
and U3032 (N_3032,N_2848,N_2944);
or U3033 (N_3033,N_2961,N_2930);
xnor U3034 (N_3034,N_2926,N_2872);
xor U3035 (N_3035,N_2825,N_2959);
xnor U3036 (N_3036,N_2795,N_2884);
nand U3037 (N_3037,N_2770,N_2831);
nand U3038 (N_3038,N_2957,N_2900);
nor U3039 (N_3039,N_2914,N_2804);
and U3040 (N_3040,N_2828,N_2941);
or U3041 (N_3041,N_2791,N_2901);
nand U3042 (N_3042,N_2816,N_2771);
or U3043 (N_3043,N_2753,N_2822);
nand U3044 (N_3044,N_2931,N_2938);
and U3045 (N_3045,N_2880,N_2905);
xnor U3046 (N_3046,N_2801,N_2940);
xnor U3047 (N_3047,N_2921,N_2802);
xor U3048 (N_3048,N_2929,N_2948);
or U3049 (N_3049,N_2803,N_2762);
nor U3050 (N_3050,N_2765,N_2755);
nor U3051 (N_3051,N_2815,N_2786);
or U3052 (N_3052,N_2764,N_2751);
or U3053 (N_3053,N_2888,N_2932);
and U3054 (N_3054,N_2854,N_2950);
and U3055 (N_3055,N_2898,N_2790);
nand U3056 (N_3056,N_2881,N_2811);
nand U3057 (N_3057,N_2813,N_2906);
and U3058 (N_3058,N_2782,N_2925);
nand U3059 (N_3059,N_2870,N_2861);
or U3060 (N_3060,N_2976,N_2852);
xor U3061 (N_3061,N_2752,N_2962);
nand U3062 (N_3062,N_2935,N_2986);
nand U3063 (N_3063,N_2937,N_2787);
nand U3064 (N_3064,N_2779,N_2863);
or U3065 (N_3065,N_2939,N_2951);
or U3066 (N_3066,N_2909,N_2895);
and U3067 (N_3067,N_2859,N_2970);
and U3068 (N_3068,N_2777,N_2936);
or U3069 (N_3069,N_2876,N_2877);
nor U3070 (N_3070,N_2783,N_2871);
or U3071 (N_3071,N_2999,N_2760);
or U3072 (N_3072,N_2963,N_2955);
nand U3073 (N_3073,N_2989,N_2924);
xor U3074 (N_3074,N_2973,N_2851);
xnor U3075 (N_3075,N_2873,N_2757);
nor U3076 (N_3076,N_2817,N_2774);
or U3077 (N_3077,N_2883,N_2890);
nor U3078 (N_3078,N_2899,N_2820);
xor U3079 (N_3079,N_2918,N_2840);
xor U3080 (N_3080,N_2988,N_2823);
and U3081 (N_3081,N_2875,N_2927);
nand U3082 (N_3082,N_2845,N_2911);
nor U3083 (N_3083,N_2853,N_2785);
or U3084 (N_3084,N_2915,N_2839);
and U3085 (N_3085,N_2796,N_2996);
xor U3086 (N_3086,N_2794,N_2885);
or U3087 (N_3087,N_2818,N_2922);
nand U3088 (N_3088,N_2878,N_2968);
nor U3089 (N_3089,N_2913,N_2889);
and U3090 (N_3090,N_2933,N_2841);
or U3091 (N_3091,N_2849,N_2773);
or U3092 (N_3092,N_2974,N_2969);
xnor U3093 (N_3093,N_2953,N_2874);
and U3094 (N_3094,N_2964,N_2778);
xnor U3095 (N_3095,N_2826,N_2834);
or U3096 (N_3096,N_2958,N_2756);
and U3097 (N_3097,N_2819,N_2891);
nor U3098 (N_3098,N_2879,N_2862);
nand U3099 (N_3099,N_2894,N_2843);
or U3100 (N_3100,N_2923,N_2812);
or U3101 (N_3101,N_2917,N_2799);
xnor U3102 (N_3102,N_2896,N_2993);
and U3103 (N_3103,N_2983,N_2805);
nor U3104 (N_3104,N_2847,N_2886);
xor U3105 (N_3105,N_2967,N_2960);
nor U3106 (N_3106,N_2928,N_2990);
and U3107 (N_3107,N_2972,N_2965);
nor U3108 (N_3108,N_2759,N_2984);
xnor U3109 (N_3109,N_2991,N_2912);
nand U3110 (N_3110,N_2908,N_2985);
nor U3111 (N_3111,N_2810,N_2893);
nor U3112 (N_3112,N_2766,N_2966);
xnor U3113 (N_3113,N_2776,N_2943);
nor U3114 (N_3114,N_2860,N_2784);
nor U3115 (N_3115,N_2829,N_2902);
or U3116 (N_3116,N_2750,N_2846);
nand U3117 (N_3117,N_2865,N_2956);
xnor U3118 (N_3118,N_2934,N_2858);
xor U3119 (N_3119,N_2903,N_2780);
or U3120 (N_3120,N_2952,N_2867);
nor U3121 (N_3121,N_2920,N_2761);
nor U3122 (N_3122,N_2855,N_2992);
xor U3123 (N_3123,N_2835,N_2781);
and U3124 (N_3124,N_2869,N_2832);
nor U3125 (N_3125,N_2953,N_2982);
nor U3126 (N_3126,N_2887,N_2956);
xnor U3127 (N_3127,N_2815,N_2810);
nor U3128 (N_3128,N_2965,N_2762);
nand U3129 (N_3129,N_2856,N_2893);
nor U3130 (N_3130,N_2771,N_2791);
nor U3131 (N_3131,N_2763,N_2807);
xnor U3132 (N_3132,N_2986,N_2968);
nand U3133 (N_3133,N_2983,N_2874);
and U3134 (N_3134,N_2869,N_2883);
xor U3135 (N_3135,N_2833,N_2790);
xnor U3136 (N_3136,N_2901,N_2779);
or U3137 (N_3137,N_2923,N_2937);
or U3138 (N_3138,N_2977,N_2836);
nand U3139 (N_3139,N_2938,N_2988);
nand U3140 (N_3140,N_2794,N_2807);
or U3141 (N_3141,N_2970,N_2898);
xnor U3142 (N_3142,N_2778,N_2832);
or U3143 (N_3143,N_2755,N_2836);
and U3144 (N_3144,N_2844,N_2956);
xnor U3145 (N_3145,N_2761,N_2792);
nor U3146 (N_3146,N_2941,N_2759);
or U3147 (N_3147,N_2938,N_2784);
or U3148 (N_3148,N_2976,N_2826);
or U3149 (N_3149,N_2983,N_2906);
or U3150 (N_3150,N_2772,N_2860);
nand U3151 (N_3151,N_2937,N_2908);
nand U3152 (N_3152,N_2766,N_2917);
nand U3153 (N_3153,N_2912,N_2804);
or U3154 (N_3154,N_2881,N_2935);
or U3155 (N_3155,N_2808,N_2802);
and U3156 (N_3156,N_2878,N_2943);
and U3157 (N_3157,N_2756,N_2835);
and U3158 (N_3158,N_2794,N_2822);
nor U3159 (N_3159,N_2911,N_2819);
and U3160 (N_3160,N_2833,N_2897);
xnor U3161 (N_3161,N_2981,N_2892);
and U3162 (N_3162,N_2940,N_2881);
xor U3163 (N_3163,N_2862,N_2832);
or U3164 (N_3164,N_2797,N_2923);
nand U3165 (N_3165,N_2928,N_2954);
xor U3166 (N_3166,N_2948,N_2827);
nand U3167 (N_3167,N_2958,N_2834);
nor U3168 (N_3168,N_2903,N_2814);
and U3169 (N_3169,N_2919,N_2929);
or U3170 (N_3170,N_2963,N_2826);
xnor U3171 (N_3171,N_2958,N_2950);
xnor U3172 (N_3172,N_2942,N_2764);
nand U3173 (N_3173,N_2779,N_2938);
xnor U3174 (N_3174,N_2943,N_2897);
or U3175 (N_3175,N_2795,N_2980);
nor U3176 (N_3176,N_2906,N_2977);
nor U3177 (N_3177,N_2969,N_2968);
xor U3178 (N_3178,N_2967,N_2901);
nor U3179 (N_3179,N_2917,N_2895);
xor U3180 (N_3180,N_2835,N_2959);
xor U3181 (N_3181,N_2915,N_2988);
nor U3182 (N_3182,N_2844,N_2752);
or U3183 (N_3183,N_2959,N_2784);
xor U3184 (N_3184,N_2935,N_2931);
nand U3185 (N_3185,N_2871,N_2929);
nor U3186 (N_3186,N_2752,N_2795);
nor U3187 (N_3187,N_2762,N_2877);
or U3188 (N_3188,N_2975,N_2882);
or U3189 (N_3189,N_2821,N_2752);
or U3190 (N_3190,N_2756,N_2841);
and U3191 (N_3191,N_2837,N_2796);
nand U3192 (N_3192,N_2771,N_2886);
nand U3193 (N_3193,N_2954,N_2940);
nand U3194 (N_3194,N_2778,N_2985);
nand U3195 (N_3195,N_2873,N_2751);
or U3196 (N_3196,N_2825,N_2806);
or U3197 (N_3197,N_2850,N_2986);
xnor U3198 (N_3198,N_2932,N_2983);
and U3199 (N_3199,N_2798,N_2899);
xnor U3200 (N_3200,N_2820,N_2995);
and U3201 (N_3201,N_2945,N_2912);
or U3202 (N_3202,N_2989,N_2885);
or U3203 (N_3203,N_2820,N_2773);
or U3204 (N_3204,N_2960,N_2938);
and U3205 (N_3205,N_2943,N_2939);
xnor U3206 (N_3206,N_2774,N_2893);
or U3207 (N_3207,N_2990,N_2923);
nor U3208 (N_3208,N_2862,N_2859);
and U3209 (N_3209,N_2776,N_2811);
xor U3210 (N_3210,N_2874,N_2872);
nand U3211 (N_3211,N_2917,N_2913);
nor U3212 (N_3212,N_2837,N_2960);
nand U3213 (N_3213,N_2993,N_2830);
xnor U3214 (N_3214,N_2861,N_2845);
xnor U3215 (N_3215,N_2767,N_2837);
xor U3216 (N_3216,N_2903,N_2862);
xnor U3217 (N_3217,N_2978,N_2913);
xnor U3218 (N_3218,N_2777,N_2962);
or U3219 (N_3219,N_2760,N_2808);
or U3220 (N_3220,N_2968,N_2864);
nand U3221 (N_3221,N_2824,N_2811);
nor U3222 (N_3222,N_2758,N_2872);
nor U3223 (N_3223,N_2987,N_2903);
or U3224 (N_3224,N_2889,N_2988);
or U3225 (N_3225,N_2824,N_2904);
xor U3226 (N_3226,N_2757,N_2977);
xor U3227 (N_3227,N_2961,N_2837);
xnor U3228 (N_3228,N_2852,N_2768);
nor U3229 (N_3229,N_2884,N_2972);
or U3230 (N_3230,N_2781,N_2800);
xnor U3231 (N_3231,N_2978,N_2782);
xor U3232 (N_3232,N_2928,N_2875);
or U3233 (N_3233,N_2967,N_2999);
and U3234 (N_3234,N_2811,N_2856);
xnor U3235 (N_3235,N_2979,N_2923);
xor U3236 (N_3236,N_2898,N_2764);
and U3237 (N_3237,N_2762,N_2815);
nor U3238 (N_3238,N_2947,N_2890);
nor U3239 (N_3239,N_2773,N_2802);
or U3240 (N_3240,N_2939,N_2793);
or U3241 (N_3241,N_2834,N_2955);
nand U3242 (N_3242,N_2883,N_2785);
xor U3243 (N_3243,N_2769,N_2778);
or U3244 (N_3244,N_2840,N_2916);
nand U3245 (N_3245,N_2953,N_2768);
or U3246 (N_3246,N_2997,N_2808);
nand U3247 (N_3247,N_2818,N_2967);
and U3248 (N_3248,N_2765,N_2953);
nor U3249 (N_3249,N_2800,N_2877);
xnor U3250 (N_3250,N_3217,N_3103);
or U3251 (N_3251,N_3008,N_3171);
nor U3252 (N_3252,N_3028,N_3180);
nand U3253 (N_3253,N_3106,N_3042);
xor U3254 (N_3254,N_3036,N_3170);
and U3255 (N_3255,N_3117,N_3218);
or U3256 (N_3256,N_3099,N_3179);
xor U3257 (N_3257,N_3080,N_3239);
or U3258 (N_3258,N_3110,N_3158);
or U3259 (N_3259,N_3151,N_3005);
and U3260 (N_3260,N_3160,N_3115);
nand U3261 (N_3261,N_3119,N_3069);
nand U3262 (N_3262,N_3079,N_3035);
xnor U3263 (N_3263,N_3240,N_3195);
nand U3264 (N_3264,N_3202,N_3121);
or U3265 (N_3265,N_3082,N_3232);
or U3266 (N_3266,N_3033,N_3246);
nand U3267 (N_3267,N_3113,N_3237);
nand U3268 (N_3268,N_3162,N_3203);
and U3269 (N_3269,N_3006,N_3076);
nor U3270 (N_3270,N_3017,N_3127);
and U3271 (N_3271,N_3230,N_3175);
nand U3272 (N_3272,N_3015,N_3053);
nand U3273 (N_3273,N_3215,N_3126);
xor U3274 (N_3274,N_3147,N_3224);
xnor U3275 (N_3275,N_3128,N_3020);
or U3276 (N_3276,N_3013,N_3130);
nor U3277 (N_3277,N_3152,N_3227);
nor U3278 (N_3278,N_3137,N_3124);
nand U3279 (N_3279,N_3003,N_3025);
or U3280 (N_3280,N_3049,N_3140);
nor U3281 (N_3281,N_3112,N_3067);
nand U3282 (N_3282,N_3010,N_3201);
or U3283 (N_3283,N_3241,N_3223);
nor U3284 (N_3284,N_3046,N_3186);
and U3285 (N_3285,N_3167,N_3163);
xnor U3286 (N_3286,N_3122,N_3037);
nand U3287 (N_3287,N_3138,N_3136);
and U3288 (N_3288,N_3095,N_3166);
or U3289 (N_3289,N_3145,N_3062);
nand U3290 (N_3290,N_3032,N_3084);
nor U3291 (N_3291,N_3209,N_3159);
nand U3292 (N_3292,N_3078,N_3018);
nand U3293 (N_3293,N_3043,N_3189);
or U3294 (N_3294,N_3029,N_3083);
xnor U3295 (N_3295,N_3088,N_3229);
xor U3296 (N_3296,N_3014,N_3068);
nand U3297 (N_3297,N_3093,N_3114);
or U3298 (N_3298,N_3208,N_3231);
and U3299 (N_3299,N_3098,N_3011);
nor U3300 (N_3300,N_3101,N_3222);
nand U3301 (N_3301,N_3055,N_3057);
nor U3302 (N_3302,N_3176,N_3225);
and U3303 (N_3303,N_3031,N_3236);
xnor U3304 (N_3304,N_3123,N_3219);
and U3305 (N_3305,N_3086,N_3199);
nor U3306 (N_3306,N_3107,N_3047);
and U3307 (N_3307,N_3038,N_3154);
xor U3308 (N_3308,N_3161,N_3148);
nor U3309 (N_3309,N_3194,N_3207);
xnor U3310 (N_3310,N_3149,N_3039);
or U3311 (N_3311,N_3129,N_3064);
nor U3312 (N_3312,N_3023,N_3181);
nor U3313 (N_3313,N_3156,N_3000);
xnor U3314 (N_3314,N_3073,N_3021);
and U3315 (N_3315,N_3234,N_3007);
nor U3316 (N_3316,N_3030,N_3193);
xnor U3317 (N_3317,N_3172,N_3085);
nor U3318 (N_3318,N_3157,N_3188);
xnor U3319 (N_3319,N_3004,N_3102);
nand U3320 (N_3320,N_3090,N_3109);
nand U3321 (N_3321,N_3089,N_3216);
and U3322 (N_3322,N_3060,N_3104);
nand U3323 (N_3323,N_3196,N_3116);
xor U3324 (N_3324,N_3168,N_3135);
or U3325 (N_3325,N_3205,N_3244);
and U3326 (N_3326,N_3243,N_3187);
nand U3327 (N_3327,N_3132,N_3174);
and U3328 (N_3328,N_3050,N_3108);
nor U3329 (N_3329,N_3092,N_3210);
or U3330 (N_3330,N_3185,N_3024);
or U3331 (N_3331,N_3146,N_3065);
and U3332 (N_3332,N_3245,N_3063);
xnor U3333 (N_3333,N_3075,N_3204);
nor U3334 (N_3334,N_3220,N_3134);
and U3335 (N_3335,N_3051,N_3077);
or U3336 (N_3336,N_3087,N_3200);
nand U3337 (N_3337,N_3183,N_3097);
nand U3338 (N_3338,N_3249,N_3071);
and U3339 (N_3339,N_3233,N_3094);
and U3340 (N_3340,N_3198,N_3058);
xnor U3341 (N_3341,N_3091,N_3081);
or U3342 (N_3342,N_3169,N_3153);
nand U3343 (N_3343,N_3143,N_3178);
nand U3344 (N_3344,N_3012,N_3206);
nand U3345 (N_3345,N_3150,N_3061);
nand U3346 (N_3346,N_3056,N_3131);
or U3347 (N_3347,N_3155,N_3173);
nand U3348 (N_3348,N_3120,N_3022);
nor U3349 (N_3349,N_3212,N_3221);
nand U3350 (N_3350,N_3184,N_3242);
and U3351 (N_3351,N_3228,N_3190);
or U3352 (N_3352,N_3027,N_3096);
or U3353 (N_3353,N_3072,N_3001);
and U3354 (N_3354,N_3070,N_3016);
xnor U3355 (N_3355,N_3111,N_3191);
xnor U3356 (N_3356,N_3045,N_3066);
xnor U3357 (N_3357,N_3177,N_3034);
nand U3358 (N_3358,N_3105,N_3182);
xor U3359 (N_3359,N_3165,N_3139);
xnor U3360 (N_3360,N_3026,N_3235);
nor U3361 (N_3361,N_3197,N_3059);
nor U3362 (N_3362,N_3164,N_3074);
xor U3363 (N_3363,N_3040,N_3041);
and U3364 (N_3364,N_3133,N_3214);
nor U3365 (N_3365,N_3226,N_3142);
and U3366 (N_3366,N_3100,N_3054);
nor U3367 (N_3367,N_3144,N_3125);
and U3368 (N_3368,N_3247,N_3192);
or U3369 (N_3369,N_3238,N_3141);
and U3370 (N_3370,N_3211,N_3019);
and U3371 (N_3371,N_3048,N_3044);
and U3372 (N_3372,N_3002,N_3213);
or U3373 (N_3373,N_3248,N_3009);
or U3374 (N_3374,N_3052,N_3118);
or U3375 (N_3375,N_3004,N_3139);
nor U3376 (N_3376,N_3233,N_3081);
or U3377 (N_3377,N_3201,N_3206);
or U3378 (N_3378,N_3042,N_3111);
nor U3379 (N_3379,N_3073,N_3097);
and U3380 (N_3380,N_3125,N_3151);
or U3381 (N_3381,N_3030,N_3248);
and U3382 (N_3382,N_3064,N_3124);
nor U3383 (N_3383,N_3162,N_3126);
or U3384 (N_3384,N_3022,N_3080);
nor U3385 (N_3385,N_3157,N_3166);
xnor U3386 (N_3386,N_3114,N_3085);
nor U3387 (N_3387,N_3037,N_3140);
or U3388 (N_3388,N_3192,N_3008);
nor U3389 (N_3389,N_3041,N_3151);
and U3390 (N_3390,N_3064,N_3158);
and U3391 (N_3391,N_3005,N_3158);
nand U3392 (N_3392,N_3219,N_3008);
nor U3393 (N_3393,N_3041,N_3076);
xor U3394 (N_3394,N_3228,N_3098);
nor U3395 (N_3395,N_3027,N_3245);
or U3396 (N_3396,N_3017,N_3223);
nor U3397 (N_3397,N_3152,N_3029);
or U3398 (N_3398,N_3010,N_3084);
and U3399 (N_3399,N_3117,N_3001);
or U3400 (N_3400,N_3002,N_3236);
or U3401 (N_3401,N_3006,N_3080);
nand U3402 (N_3402,N_3129,N_3110);
and U3403 (N_3403,N_3218,N_3043);
nand U3404 (N_3404,N_3051,N_3229);
or U3405 (N_3405,N_3190,N_3162);
nor U3406 (N_3406,N_3164,N_3055);
and U3407 (N_3407,N_3167,N_3135);
and U3408 (N_3408,N_3126,N_3145);
nand U3409 (N_3409,N_3003,N_3181);
xnor U3410 (N_3410,N_3115,N_3031);
xor U3411 (N_3411,N_3220,N_3037);
and U3412 (N_3412,N_3058,N_3201);
xnor U3413 (N_3413,N_3190,N_3030);
xnor U3414 (N_3414,N_3067,N_3200);
or U3415 (N_3415,N_3043,N_3209);
nor U3416 (N_3416,N_3223,N_3007);
xor U3417 (N_3417,N_3229,N_3023);
nand U3418 (N_3418,N_3206,N_3211);
nor U3419 (N_3419,N_3027,N_3139);
nor U3420 (N_3420,N_3012,N_3219);
xor U3421 (N_3421,N_3013,N_3212);
nor U3422 (N_3422,N_3163,N_3021);
nand U3423 (N_3423,N_3224,N_3220);
nand U3424 (N_3424,N_3218,N_3096);
and U3425 (N_3425,N_3016,N_3186);
or U3426 (N_3426,N_3196,N_3195);
nor U3427 (N_3427,N_3202,N_3135);
or U3428 (N_3428,N_3221,N_3053);
nor U3429 (N_3429,N_3187,N_3039);
nor U3430 (N_3430,N_3046,N_3057);
xor U3431 (N_3431,N_3234,N_3220);
and U3432 (N_3432,N_3174,N_3091);
nand U3433 (N_3433,N_3212,N_3075);
or U3434 (N_3434,N_3025,N_3190);
xor U3435 (N_3435,N_3091,N_3033);
and U3436 (N_3436,N_3040,N_3198);
nand U3437 (N_3437,N_3209,N_3099);
xor U3438 (N_3438,N_3238,N_3044);
xor U3439 (N_3439,N_3197,N_3070);
or U3440 (N_3440,N_3140,N_3176);
nor U3441 (N_3441,N_3201,N_3241);
nand U3442 (N_3442,N_3209,N_3182);
or U3443 (N_3443,N_3151,N_3032);
or U3444 (N_3444,N_3233,N_3207);
nor U3445 (N_3445,N_3203,N_3085);
or U3446 (N_3446,N_3052,N_3113);
xor U3447 (N_3447,N_3106,N_3185);
xnor U3448 (N_3448,N_3016,N_3102);
nor U3449 (N_3449,N_3130,N_3073);
nand U3450 (N_3450,N_3121,N_3040);
nand U3451 (N_3451,N_3056,N_3029);
nor U3452 (N_3452,N_3233,N_3225);
nand U3453 (N_3453,N_3175,N_3171);
nor U3454 (N_3454,N_3021,N_3043);
or U3455 (N_3455,N_3237,N_3092);
or U3456 (N_3456,N_3115,N_3100);
and U3457 (N_3457,N_3214,N_3181);
and U3458 (N_3458,N_3238,N_3247);
or U3459 (N_3459,N_3196,N_3027);
nand U3460 (N_3460,N_3090,N_3202);
xor U3461 (N_3461,N_3172,N_3003);
nor U3462 (N_3462,N_3066,N_3108);
nor U3463 (N_3463,N_3112,N_3126);
and U3464 (N_3464,N_3202,N_3200);
or U3465 (N_3465,N_3244,N_3164);
nand U3466 (N_3466,N_3105,N_3054);
nor U3467 (N_3467,N_3164,N_3123);
xor U3468 (N_3468,N_3194,N_3210);
nor U3469 (N_3469,N_3049,N_3036);
and U3470 (N_3470,N_3139,N_3112);
nor U3471 (N_3471,N_3021,N_3010);
nor U3472 (N_3472,N_3147,N_3171);
xor U3473 (N_3473,N_3001,N_3050);
or U3474 (N_3474,N_3104,N_3198);
or U3475 (N_3475,N_3153,N_3228);
or U3476 (N_3476,N_3113,N_3018);
nand U3477 (N_3477,N_3032,N_3062);
or U3478 (N_3478,N_3067,N_3113);
nor U3479 (N_3479,N_3091,N_3242);
nor U3480 (N_3480,N_3145,N_3142);
xor U3481 (N_3481,N_3213,N_3062);
and U3482 (N_3482,N_3246,N_3160);
nor U3483 (N_3483,N_3068,N_3049);
nand U3484 (N_3484,N_3039,N_3150);
xor U3485 (N_3485,N_3156,N_3044);
nor U3486 (N_3486,N_3143,N_3123);
or U3487 (N_3487,N_3033,N_3058);
and U3488 (N_3488,N_3065,N_3106);
or U3489 (N_3489,N_3070,N_3043);
and U3490 (N_3490,N_3205,N_3033);
xnor U3491 (N_3491,N_3186,N_3011);
xor U3492 (N_3492,N_3012,N_3003);
nor U3493 (N_3493,N_3240,N_3045);
and U3494 (N_3494,N_3109,N_3081);
or U3495 (N_3495,N_3058,N_3221);
xnor U3496 (N_3496,N_3051,N_3075);
nand U3497 (N_3497,N_3212,N_3116);
xnor U3498 (N_3498,N_3173,N_3162);
and U3499 (N_3499,N_3143,N_3106);
nor U3500 (N_3500,N_3487,N_3280);
xor U3501 (N_3501,N_3335,N_3349);
xnor U3502 (N_3502,N_3459,N_3479);
nand U3503 (N_3503,N_3347,N_3252);
xor U3504 (N_3504,N_3442,N_3320);
nand U3505 (N_3505,N_3283,N_3463);
and U3506 (N_3506,N_3375,N_3438);
nor U3507 (N_3507,N_3289,N_3414);
and U3508 (N_3508,N_3425,N_3431);
and U3509 (N_3509,N_3476,N_3398);
nand U3510 (N_3510,N_3344,N_3358);
xnor U3511 (N_3511,N_3295,N_3357);
nand U3512 (N_3512,N_3382,N_3352);
and U3513 (N_3513,N_3466,N_3361);
or U3514 (N_3514,N_3415,N_3269);
and U3515 (N_3515,N_3498,N_3403);
nor U3516 (N_3516,N_3406,N_3342);
xnor U3517 (N_3517,N_3462,N_3400);
and U3518 (N_3518,N_3376,N_3418);
nor U3519 (N_3519,N_3278,N_3381);
xnor U3520 (N_3520,N_3451,N_3399);
or U3521 (N_3521,N_3273,N_3363);
nor U3522 (N_3522,N_3341,N_3338);
nor U3523 (N_3523,N_3493,N_3259);
and U3524 (N_3524,N_3480,N_3276);
or U3525 (N_3525,N_3460,N_3397);
xnor U3526 (N_3526,N_3380,N_3478);
or U3527 (N_3527,N_3383,N_3263);
xnor U3528 (N_3528,N_3410,N_3465);
xnor U3529 (N_3529,N_3299,N_3481);
or U3530 (N_3530,N_3390,N_3339);
nand U3531 (N_3531,N_3433,N_3319);
and U3532 (N_3532,N_3251,N_3346);
or U3533 (N_3533,N_3302,N_3270);
xor U3534 (N_3534,N_3353,N_3440);
and U3535 (N_3535,N_3362,N_3387);
xnor U3536 (N_3536,N_3419,N_3405);
xnor U3537 (N_3537,N_3277,N_3354);
and U3538 (N_3538,N_3321,N_3391);
xnor U3539 (N_3539,N_3429,N_3483);
and U3540 (N_3540,N_3286,N_3298);
xnor U3541 (N_3541,N_3492,N_3271);
nor U3542 (N_3542,N_3309,N_3413);
and U3543 (N_3543,N_3450,N_3407);
or U3544 (N_3544,N_3448,N_3323);
nor U3545 (N_3545,N_3261,N_3472);
nand U3546 (N_3546,N_3423,N_3422);
or U3547 (N_3547,N_3260,N_3337);
xnor U3548 (N_3548,N_3444,N_3435);
or U3549 (N_3549,N_3365,N_3436);
and U3550 (N_3550,N_3474,N_3386);
and U3551 (N_3551,N_3475,N_3432);
nor U3552 (N_3552,N_3256,N_3412);
and U3553 (N_3553,N_3470,N_3464);
nor U3554 (N_3554,N_3409,N_3421);
and U3555 (N_3555,N_3351,N_3332);
or U3556 (N_3556,N_3402,N_3385);
nand U3557 (N_3557,N_3439,N_3424);
xor U3558 (N_3558,N_3284,N_3427);
nand U3559 (N_3559,N_3485,N_3411);
xor U3560 (N_3560,N_3486,N_3304);
and U3561 (N_3561,N_3404,N_3275);
nor U3562 (N_3562,N_3279,N_3272);
nor U3563 (N_3563,N_3258,N_3288);
or U3564 (N_3564,N_3325,N_3262);
nor U3565 (N_3565,N_3453,N_3452);
and U3566 (N_3566,N_3310,N_3489);
or U3567 (N_3567,N_3458,N_3447);
nand U3568 (N_3568,N_3360,N_3328);
nand U3569 (N_3569,N_3308,N_3355);
nor U3570 (N_3570,N_3467,N_3292);
or U3571 (N_3571,N_3408,N_3281);
nor U3572 (N_3572,N_3446,N_3266);
xnor U3573 (N_3573,N_3428,N_3255);
nand U3574 (N_3574,N_3396,N_3377);
xnor U3575 (N_3575,N_3454,N_3265);
xnor U3576 (N_3576,N_3374,N_3471);
nand U3577 (N_3577,N_3426,N_3291);
nor U3578 (N_3578,N_3268,N_3401);
nand U3579 (N_3579,N_3322,N_3333);
xnor U3580 (N_3580,N_3345,N_3364);
or U3581 (N_3581,N_3297,N_3379);
or U3582 (N_3582,N_3469,N_3378);
nor U3583 (N_3583,N_3324,N_3494);
nand U3584 (N_3584,N_3334,N_3370);
or U3585 (N_3585,N_3497,N_3372);
nand U3586 (N_3586,N_3416,N_3317);
or U3587 (N_3587,N_3343,N_3253);
nand U3588 (N_3588,N_3490,N_3457);
and U3589 (N_3589,N_3484,N_3434);
xor U3590 (N_3590,N_3392,N_3395);
or U3591 (N_3591,N_3449,N_3257);
or U3592 (N_3592,N_3488,N_3312);
xnor U3593 (N_3593,N_3430,N_3293);
or U3594 (N_3594,N_3329,N_3499);
and U3595 (N_3595,N_3441,N_3282);
and U3596 (N_3596,N_3294,N_3473);
or U3597 (N_3597,N_3371,N_3356);
nor U3598 (N_3598,N_3327,N_3330);
nand U3599 (N_3599,N_3326,N_3331);
or U3600 (N_3600,N_3443,N_3316);
and U3601 (N_3601,N_3496,N_3373);
xor U3602 (N_3602,N_3274,N_3388);
nand U3603 (N_3603,N_3340,N_3287);
nand U3604 (N_3604,N_3359,N_3314);
nand U3605 (N_3605,N_3384,N_3420);
or U3606 (N_3606,N_3394,N_3267);
nor U3607 (N_3607,N_3368,N_3468);
and U3608 (N_3608,N_3348,N_3336);
xor U3609 (N_3609,N_3437,N_3306);
or U3610 (N_3610,N_3300,N_3495);
and U3611 (N_3611,N_3250,N_3254);
nand U3612 (N_3612,N_3445,N_3315);
xor U3613 (N_3613,N_3313,N_3366);
xor U3614 (N_3614,N_3301,N_3455);
nand U3615 (N_3615,N_3311,N_3307);
nand U3616 (N_3616,N_3482,N_3318);
and U3617 (N_3617,N_3369,N_3305);
xnor U3618 (N_3618,N_3264,N_3367);
nand U3619 (N_3619,N_3296,N_3393);
nor U3620 (N_3620,N_3303,N_3477);
nand U3621 (N_3621,N_3389,N_3417);
and U3622 (N_3622,N_3456,N_3285);
nand U3623 (N_3623,N_3290,N_3461);
or U3624 (N_3624,N_3491,N_3350);
and U3625 (N_3625,N_3365,N_3286);
xnor U3626 (N_3626,N_3295,N_3454);
xnor U3627 (N_3627,N_3388,N_3370);
and U3628 (N_3628,N_3262,N_3456);
xnor U3629 (N_3629,N_3468,N_3319);
nor U3630 (N_3630,N_3255,N_3389);
nor U3631 (N_3631,N_3428,N_3368);
nand U3632 (N_3632,N_3343,N_3251);
or U3633 (N_3633,N_3319,N_3465);
nor U3634 (N_3634,N_3347,N_3259);
xor U3635 (N_3635,N_3460,N_3426);
and U3636 (N_3636,N_3368,N_3392);
nand U3637 (N_3637,N_3429,N_3409);
or U3638 (N_3638,N_3457,N_3458);
and U3639 (N_3639,N_3496,N_3439);
xor U3640 (N_3640,N_3348,N_3310);
nor U3641 (N_3641,N_3459,N_3315);
and U3642 (N_3642,N_3258,N_3359);
nand U3643 (N_3643,N_3333,N_3466);
xor U3644 (N_3644,N_3386,N_3291);
xnor U3645 (N_3645,N_3483,N_3329);
xor U3646 (N_3646,N_3384,N_3312);
xnor U3647 (N_3647,N_3384,N_3293);
xnor U3648 (N_3648,N_3494,N_3443);
nor U3649 (N_3649,N_3489,N_3393);
nor U3650 (N_3650,N_3273,N_3486);
nor U3651 (N_3651,N_3455,N_3498);
nand U3652 (N_3652,N_3497,N_3297);
and U3653 (N_3653,N_3279,N_3439);
or U3654 (N_3654,N_3464,N_3461);
nor U3655 (N_3655,N_3495,N_3281);
xor U3656 (N_3656,N_3429,N_3261);
nor U3657 (N_3657,N_3375,N_3390);
and U3658 (N_3658,N_3327,N_3408);
xnor U3659 (N_3659,N_3253,N_3447);
nor U3660 (N_3660,N_3467,N_3372);
and U3661 (N_3661,N_3322,N_3365);
xnor U3662 (N_3662,N_3300,N_3276);
and U3663 (N_3663,N_3375,N_3329);
nand U3664 (N_3664,N_3439,N_3475);
and U3665 (N_3665,N_3261,N_3446);
nor U3666 (N_3666,N_3316,N_3404);
xnor U3667 (N_3667,N_3438,N_3429);
xnor U3668 (N_3668,N_3437,N_3433);
and U3669 (N_3669,N_3418,N_3385);
and U3670 (N_3670,N_3275,N_3484);
or U3671 (N_3671,N_3414,N_3290);
and U3672 (N_3672,N_3421,N_3366);
nor U3673 (N_3673,N_3418,N_3494);
xnor U3674 (N_3674,N_3466,N_3396);
nor U3675 (N_3675,N_3423,N_3485);
and U3676 (N_3676,N_3394,N_3351);
and U3677 (N_3677,N_3363,N_3277);
and U3678 (N_3678,N_3463,N_3266);
xor U3679 (N_3679,N_3419,N_3332);
or U3680 (N_3680,N_3326,N_3433);
or U3681 (N_3681,N_3450,N_3352);
nand U3682 (N_3682,N_3314,N_3459);
nand U3683 (N_3683,N_3389,N_3394);
nand U3684 (N_3684,N_3310,N_3473);
xnor U3685 (N_3685,N_3450,N_3354);
nand U3686 (N_3686,N_3368,N_3284);
nand U3687 (N_3687,N_3301,N_3424);
or U3688 (N_3688,N_3355,N_3345);
xnor U3689 (N_3689,N_3411,N_3314);
or U3690 (N_3690,N_3327,N_3313);
and U3691 (N_3691,N_3450,N_3348);
nand U3692 (N_3692,N_3459,N_3451);
nand U3693 (N_3693,N_3401,N_3294);
nand U3694 (N_3694,N_3346,N_3305);
and U3695 (N_3695,N_3292,N_3347);
nor U3696 (N_3696,N_3324,N_3414);
nand U3697 (N_3697,N_3347,N_3417);
and U3698 (N_3698,N_3334,N_3477);
xor U3699 (N_3699,N_3358,N_3490);
or U3700 (N_3700,N_3386,N_3358);
xnor U3701 (N_3701,N_3472,N_3310);
and U3702 (N_3702,N_3300,N_3354);
or U3703 (N_3703,N_3260,N_3344);
and U3704 (N_3704,N_3409,N_3392);
nor U3705 (N_3705,N_3377,N_3436);
xor U3706 (N_3706,N_3407,N_3436);
and U3707 (N_3707,N_3281,N_3318);
xnor U3708 (N_3708,N_3309,N_3369);
xnor U3709 (N_3709,N_3422,N_3491);
or U3710 (N_3710,N_3423,N_3438);
nand U3711 (N_3711,N_3399,N_3336);
nor U3712 (N_3712,N_3490,N_3458);
and U3713 (N_3713,N_3269,N_3449);
nor U3714 (N_3714,N_3461,N_3469);
xor U3715 (N_3715,N_3318,N_3433);
and U3716 (N_3716,N_3291,N_3341);
nor U3717 (N_3717,N_3339,N_3452);
or U3718 (N_3718,N_3267,N_3264);
or U3719 (N_3719,N_3467,N_3450);
nor U3720 (N_3720,N_3480,N_3360);
and U3721 (N_3721,N_3278,N_3347);
or U3722 (N_3722,N_3411,N_3361);
nand U3723 (N_3723,N_3375,N_3429);
nor U3724 (N_3724,N_3487,N_3337);
and U3725 (N_3725,N_3318,N_3473);
nor U3726 (N_3726,N_3384,N_3354);
xnor U3727 (N_3727,N_3326,N_3277);
nor U3728 (N_3728,N_3274,N_3383);
nor U3729 (N_3729,N_3403,N_3437);
nand U3730 (N_3730,N_3450,N_3280);
and U3731 (N_3731,N_3422,N_3430);
xnor U3732 (N_3732,N_3350,N_3250);
and U3733 (N_3733,N_3357,N_3314);
or U3734 (N_3734,N_3266,N_3418);
or U3735 (N_3735,N_3257,N_3354);
nor U3736 (N_3736,N_3495,N_3320);
nor U3737 (N_3737,N_3442,N_3472);
or U3738 (N_3738,N_3326,N_3383);
xor U3739 (N_3739,N_3434,N_3327);
xor U3740 (N_3740,N_3298,N_3315);
and U3741 (N_3741,N_3305,N_3429);
or U3742 (N_3742,N_3404,N_3337);
or U3743 (N_3743,N_3259,N_3335);
and U3744 (N_3744,N_3262,N_3495);
nand U3745 (N_3745,N_3416,N_3463);
nor U3746 (N_3746,N_3404,N_3345);
xor U3747 (N_3747,N_3458,N_3397);
or U3748 (N_3748,N_3391,N_3384);
and U3749 (N_3749,N_3379,N_3388);
xnor U3750 (N_3750,N_3635,N_3629);
and U3751 (N_3751,N_3634,N_3605);
or U3752 (N_3752,N_3707,N_3595);
nor U3753 (N_3753,N_3659,N_3661);
or U3754 (N_3754,N_3719,N_3645);
or U3755 (N_3755,N_3510,N_3601);
xnor U3756 (N_3756,N_3523,N_3552);
or U3757 (N_3757,N_3647,N_3614);
nor U3758 (N_3758,N_3714,N_3585);
xor U3759 (N_3759,N_3651,N_3726);
nand U3760 (N_3760,N_3607,N_3620);
or U3761 (N_3761,N_3644,N_3716);
nor U3762 (N_3762,N_3710,N_3658);
xor U3763 (N_3763,N_3618,N_3590);
or U3764 (N_3764,N_3638,N_3627);
nor U3765 (N_3765,N_3515,N_3741);
or U3766 (N_3766,N_3666,N_3583);
nor U3767 (N_3767,N_3554,N_3739);
nor U3768 (N_3768,N_3597,N_3530);
nand U3769 (N_3769,N_3631,N_3591);
nand U3770 (N_3770,N_3720,N_3536);
or U3771 (N_3771,N_3551,N_3587);
nand U3772 (N_3772,N_3640,N_3520);
and U3773 (N_3773,N_3503,N_3539);
or U3774 (N_3774,N_3692,N_3722);
nand U3775 (N_3775,N_3660,N_3600);
nand U3776 (N_3776,N_3648,N_3745);
or U3777 (N_3777,N_3502,N_3636);
and U3778 (N_3778,N_3557,N_3513);
nand U3779 (N_3779,N_3748,N_3695);
nand U3780 (N_3780,N_3561,N_3671);
or U3781 (N_3781,N_3681,N_3623);
xnor U3782 (N_3782,N_3559,N_3519);
nand U3783 (N_3783,N_3596,N_3628);
nor U3784 (N_3784,N_3594,N_3678);
nand U3785 (N_3785,N_3565,N_3746);
xor U3786 (N_3786,N_3579,N_3641);
and U3787 (N_3787,N_3679,N_3526);
xnor U3788 (N_3788,N_3700,N_3732);
xor U3789 (N_3789,N_3699,N_3609);
or U3790 (N_3790,N_3571,N_3549);
and U3791 (N_3791,N_3673,N_3735);
and U3792 (N_3792,N_3617,N_3599);
nand U3793 (N_3793,N_3672,N_3637);
nor U3794 (N_3794,N_3507,N_3667);
xor U3795 (N_3795,N_3553,N_3740);
xnor U3796 (N_3796,N_3567,N_3531);
nand U3797 (N_3797,N_3569,N_3577);
nand U3798 (N_3798,N_3603,N_3548);
and U3799 (N_3799,N_3622,N_3527);
or U3800 (N_3800,N_3731,N_3742);
nor U3801 (N_3801,N_3506,N_3537);
or U3802 (N_3802,N_3524,N_3540);
or U3803 (N_3803,N_3509,N_3542);
nor U3804 (N_3804,N_3602,N_3684);
nand U3805 (N_3805,N_3690,N_3514);
nand U3806 (N_3806,N_3535,N_3687);
nor U3807 (N_3807,N_3576,N_3677);
nand U3808 (N_3808,N_3717,N_3642);
nand U3809 (N_3809,N_3639,N_3703);
or U3810 (N_3810,N_3737,N_3697);
and U3811 (N_3811,N_3630,N_3545);
and U3812 (N_3812,N_3500,N_3625);
or U3813 (N_3813,N_3566,N_3501);
nand U3814 (N_3814,N_3610,N_3749);
and U3815 (N_3815,N_3588,N_3615);
or U3816 (N_3816,N_3619,N_3706);
nand U3817 (N_3817,N_3543,N_3680);
xor U3818 (N_3818,N_3532,N_3705);
nand U3819 (N_3819,N_3611,N_3516);
nand U3820 (N_3820,N_3547,N_3698);
or U3821 (N_3821,N_3562,N_3612);
xor U3822 (N_3822,N_3743,N_3589);
nor U3823 (N_3823,N_3708,N_3721);
nor U3824 (N_3824,N_3581,N_3688);
nor U3825 (N_3825,N_3655,N_3682);
and U3826 (N_3826,N_3693,N_3546);
or U3827 (N_3827,N_3694,N_3723);
and U3828 (N_3828,N_3649,N_3729);
or U3829 (N_3829,N_3675,N_3534);
or U3830 (N_3830,N_3712,N_3616);
and U3831 (N_3831,N_3522,N_3517);
nor U3832 (N_3832,N_3696,N_3633);
or U3833 (N_3833,N_3704,N_3715);
or U3834 (N_3834,N_3727,N_3574);
nor U3835 (N_3835,N_3730,N_3738);
nor U3836 (N_3836,N_3580,N_3573);
nor U3837 (N_3837,N_3643,N_3701);
or U3838 (N_3838,N_3568,N_3654);
and U3839 (N_3839,N_3572,N_3550);
or U3840 (N_3840,N_3686,N_3511);
or U3841 (N_3841,N_3593,N_3725);
nor U3842 (N_3842,N_3747,N_3670);
xor U3843 (N_3843,N_3663,N_3560);
xnor U3844 (N_3844,N_3683,N_3504);
nand U3845 (N_3845,N_3653,N_3613);
or U3846 (N_3846,N_3578,N_3584);
xor U3847 (N_3847,N_3505,N_3656);
or U3848 (N_3848,N_3652,N_3529);
or U3849 (N_3849,N_3702,N_3512);
or U3850 (N_3850,N_3736,N_3668);
or U3851 (N_3851,N_3713,N_3563);
nor U3852 (N_3852,N_3621,N_3604);
nor U3853 (N_3853,N_3624,N_3662);
nand U3854 (N_3854,N_3592,N_3538);
nor U3855 (N_3855,N_3674,N_3669);
and U3856 (N_3856,N_3508,N_3709);
or U3857 (N_3857,N_3676,N_3606);
nor U3858 (N_3858,N_3711,N_3734);
and U3859 (N_3859,N_3575,N_3570);
or U3860 (N_3860,N_3586,N_3528);
or U3861 (N_3861,N_3646,N_3608);
nand U3862 (N_3862,N_3744,N_3521);
and U3863 (N_3863,N_3598,N_3733);
xor U3864 (N_3864,N_3533,N_3582);
nor U3865 (N_3865,N_3541,N_3555);
nand U3866 (N_3866,N_3626,N_3728);
xor U3867 (N_3867,N_3544,N_3518);
nand U3868 (N_3868,N_3657,N_3650);
xnor U3869 (N_3869,N_3664,N_3632);
and U3870 (N_3870,N_3724,N_3525);
and U3871 (N_3871,N_3556,N_3564);
xor U3872 (N_3872,N_3691,N_3718);
or U3873 (N_3873,N_3665,N_3558);
and U3874 (N_3874,N_3689,N_3685);
nor U3875 (N_3875,N_3588,N_3651);
xor U3876 (N_3876,N_3529,N_3734);
xor U3877 (N_3877,N_3524,N_3545);
xor U3878 (N_3878,N_3686,N_3587);
and U3879 (N_3879,N_3709,N_3603);
xnor U3880 (N_3880,N_3613,N_3592);
nor U3881 (N_3881,N_3503,N_3683);
xnor U3882 (N_3882,N_3524,N_3705);
nor U3883 (N_3883,N_3688,N_3707);
xnor U3884 (N_3884,N_3658,N_3501);
or U3885 (N_3885,N_3652,N_3619);
nor U3886 (N_3886,N_3597,N_3578);
xor U3887 (N_3887,N_3537,N_3659);
xor U3888 (N_3888,N_3714,N_3670);
and U3889 (N_3889,N_3736,N_3604);
or U3890 (N_3890,N_3709,N_3716);
xnor U3891 (N_3891,N_3515,N_3564);
or U3892 (N_3892,N_3612,N_3671);
nor U3893 (N_3893,N_3700,N_3524);
xor U3894 (N_3894,N_3510,N_3681);
and U3895 (N_3895,N_3686,N_3603);
and U3896 (N_3896,N_3526,N_3692);
or U3897 (N_3897,N_3519,N_3605);
xnor U3898 (N_3898,N_3591,N_3639);
xnor U3899 (N_3899,N_3636,N_3655);
nand U3900 (N_3900,N_3546,N_3685);
or U3901 (N_3901,N_3581,N_3682);
xor U3902 (N_3902,N_3528,N_3660);
xnor U3903 (N_3903,N_3637,N_3632);
nor U3904 (N_3904,N_3554,N_3700);
xnor U3905 (N_3905,N_3600,N_3619);
or U3906 (N_3906,N_3694,N_3658);
nand U3907 (N_3907,N_3743,N_3520);
and U3908 (N_3908,N_3567,N_3659);
or U3909 (N_3909,N_3681,N_3688);
nand U3910 (N_3910,N_3650,N_3515);
and U3911 (N_3911,N_3673,N_3573);
or U3912 (N_3912,N_3584,N_3526);
nand U3913 (N_3913,N_3698,N_3689);
nand U3914 (N_3914,N_3687,N_3744);
or U3915 (N_3915,N_3590,N_3539);
or U3916 (N_3916,N_3693,N_3682);
and U3917 (N_3917,N_3652,N_3744);
or U3918 (N_3918,N_3541,N_3697);
xnor U3919 (N_3919,N_3648,N_3583);
nand U3920 (N_3920,N_3644,N_3562);
nor U3921 (N_3921,N_3725,N_3686);
nand U3922 (N_3922,N_3611,N_3667);
nor U3923 (N_3923,N_3734,N_3610);
and U3924 (N_3924,N_3573,N_3735);
xnor U3925 (N_3925,N_3569,N_3603);
xor U3926 (N_3926,N_3669,N_3613);
or U3927 (N_3927,N_3697,N_3675);
xor U3928 (N_3928,N_3722,N_3723);
xnor U3929 (N_3929,N_3583,N_3748);
xnor U3930 (N_3930,N_3529,N_3735);
and U3931 (N_3931,N_3506,N_3646);
and U3932 (N_3932,N_3559,N_3500);
nand U3933 (N_3933,N_3642,N_3500);
nand U3934 (N_3934,N_3725,N_3534);
and U3935 (N_3935,N_3525,N_3656);
xor U3936 (N_3936,N_3512,N_3532);
and U3937 (N_3937,N_3675,N_3722);
and U3938 (N_3938,N_3666,N_3527);
and U3939 (N_3939,N_3671,N_3656);
nand U3940 (N_3940,N_3731,N_3718);
nor U3941 (N_3941,N_3678,N_3735);
xnor U3942 (N_3942,N_3603,N_3657);
or U3943 (N_3943,N_3641,N_3541);
nor U3944 (N_3944,N_3600,N_3605);
nor U3945 (N_3945,N_3606,N_3646);
nor U3946 (N_3946,N_3557,N_3702);
nand U3947 (N_3947,N_3642,N_3737);
nor U3948 (N_3948,N_3525,N_3635);
xnor U3949 (N_3949,N_3582,N_3720);
and U3950 (N_3950,N_3529,N_3554);
or U3951 (N_3951,N_3736,N_3571);
and U3952 (N_3952,N_3615,N_3731);
nor U3953 (N_3953,N_3568,N_3577);
xnor U3954 (N_3954,N_3545,N_3571);
nand U3955 (N_3955,N_3695,N_3621);
nor U3956 (N_3956,N_3631,N_3608);
nand U3957 (N_3957,N_3637,N_3556);
xnor U3958 (N_3958,N_3727,N_3505);
and U3959 (N_3959,N_3626,N_3660);
nor U3960 (N_3960,N_3521,N_3668);
xnor U3961 (N_3961,N_3715,N_3718);
xnor U3962 (N_3962,N_3620,N_3646);
and U3963 (N_3963,N_3604,N_3575);
and U3964 (N_3964,N_3724,N_3691);
xor U3965 (N_3965,N_3593,N_3599);
or U3966 (N_3966,N_3584,N_3510);
nand U3967 (N_3967,N_3713,N_3670);
nand U3968 (N_3968,N_3719,N_3529);
and U3969 (N_3969,N_3690,N_3711);
or U3970 (N_3970,N_3593,N_3701);
nand U3971 (N_3971,N_3554,N_3524);
and U3972 (N_3972,N_3726,N_3527);
nand U3973 (N_3973,N_3624,N_3565);
nor U3974 (N_3974,N_3530,N_3695);
and U3975 (N_3975,N_3642,N_3610);
nand U3976 (N_3976,N_3716,N_3605);
or U3977 (N_3977,N_3715,N_3682);
and U3978 (N_3978,N_3583,N_3543);
nand U3979 (N_3979,N_3733,N_3730);
xor U3980 (N_3980,N_3571,N_3657);
nand U3981 (N_3981,N_3673,N_3564);
or U3982 (N_3982,N_3654,N_3554);
nand U3983 (N_3983,N_3617,N_3592);
nor U3984 (N_3984,N_3637,N_3720);
nor U3985 (N_3985,N_3500,N_3724);
and U3986 (N_3986,N_3704,N_3598);
nor U3987 (N_3987,N_3516,N_3662);
xnor U3988 (N_3988,N_3607,N_3584);
or U3989 (N_3989,N_3700,N_3629);
nand U3990 (N_3990,N_3649,N_3733);
nand U3991 (N_3991,N_3733,N_3677);
nor U3992 (N_3992,N_3612,N_3738);
xnor U3993 (N_3993,N_3646,N_3650);
and U3994 (N_3994,N_3749,N_3665);
nand U3995 (N_3995,N_3746,N_3511);
or U3996 (N_3996,N_3556,N_3700);
nor U3997 (N_3997,N_3698,N_3735);
or U3998 (N_3998,N_3580,N_3746);
xnor U3999 (N_3999,N_3599,N_3669);
xor U4000 (N_4000,N_3855,N_3750);
or U4001 (N_4001,N_3790,N_3769);
and U4002 (N_4002,N_3977,N_3998);
or U4003 (N_4003,N_3800,N_3816);
xnor U4004 (N_4004,N_3797,N_3980);
and U4005 (N_4005,N_3793,N_3883);
nor U4006 (N_4006,N_3838,N_3831);
xnor U4007 (N_4007,N_3969,N_3988);
or U4008 (N_4008,N_3906,N_3939);
nand U4009 (N_4009,N_3914,N_3785);
or U4010 (N_4010,N_3928,N_3801);
nor U4011 (N_4011,N_3865,N_3956);
xor U4012 (N_4012,N_3994,N_3978);
or U4013 (N_4013,N_3965,N_3915);
and U4014 (N_4014,N_3751,N_3856);
and U4015 (N_4015,N_3817,N_3786);
xor U4016 (N_4016,N_3889,N_3820);
or U4017 (N_4017,N_3905,N_3760);
nand U4018 (N_4018,N_3992,N_3904);
and U4019 (N_4019,N_3806,N_3868);
and U4020 (N_4020,N_3850,N_3986);
nand U4021 (N_4021,N_3964,N_3772);
xnor U4022 (N_4022,N_3809,N_3872);
xor U4023 (N_4023,N_3822,N_3810);
nand U4024 (N_4024,N_3877,N_3869);
or U4025 (N_4025,N_3794,N_3918);
nand U4026 (N_4026,N_3803,N_3879);
or U4027 (N_4027,N_3972,N_3976);
nand U4028 (N_4028,N_3917,N_3788);
or U4029 (N_4029,N_3871,N_3922);
nor U4030 (N_4030,N_3840,N_3948);
nand U4031 (N_4031,N_3919,N_3759);
nor U4032 (N_4032,N_3848,N_3881);
xnor U4033 (N_4033,N_3947,N_3863);
and U4034 (N_4034,N_3824,N_3890);
nand U4035 (N_4035,N_3973,N_3970);
and U4036 (N_4036,N_3814,N_3934);
nand U4037 (N_4037,N_3908,N_3841);
and U4038 (N_4038,N_3828,N_3784);
nand U4039 (N_4039,N_3950,N_3954);
xnor U4040 (N_4040,N_3953,N_3882);
and U4041 (N_4041,N_3787,N_3993);
xnor U4042 (N_4042,N_3896,N_3899);
nand U4043 (N_4043,N_3911,N_3995);
xnor U4044 (N_4044,N_3913,N_3932);
xnor U4045 (N_4045,N_3952,N_3791);
nor U4046 (N_4046,N_3891,N_3756);
nand U4047 (N_4047,N_3999,N_3780);
nor U4048 (N_4048,N_3781,N_3862);
nor U4049 (N_4049,N_3762,N_3900);
and U4050 (N_4050,N_3808,N_3774);
nor U4051 (N_4051,N_3961,N_3929);
nand U4052 (N_4052,N_3847,N_3842);
and U4053 (N_4053,N_3955,N_3778);
and U4054 (N_4054,N_3893,N_3827);
nor U4055 (N_4055,N_3851,N_3974);
or U4056 (N_4056,N_3798,N_3894);
and U4057 (N_4057,N_3942,N_3935);
or U4058 (N_4058,N_3864,N_3873);
and U4059 (N_4059,N_3898,N_3807);
xor U4060 (N_4060,N_3990,N_3799);
nor U4061 (N_4061,N_3936,N_3958);
or U4062 (N_4062,N_3897,N_3779);
and U4063 (N_4063,N_3860,N_3804);
nor U4064 (N_4064,N_3776,N_3854);
and U4065 (N_4065,N_3792,N_3996);
nor U4066 (N_4066,N_3885,N_3796);
or U4067 (N_4067,N_3773,N_3761);
nand U4068 (N_4068,N_3819,N_3921);
and U4069 (N_4069,N_3937,N_3823);
xor U4070 (N_4070,N_3920,N_3907);
nand U4071 (N_4071,N_3775,N_3979);
and U4072 (N_4072,N_3924,N_3834);
nand U4073 (N_4073,N_3984,N_3811);
nand U4074 (N_4074,N_3876,N_3870);
nor U4075 (N_4075,N_3821,N_3857);
xor U4076 (N_4076,N_3829,N_3933);
nand U4077 (N_4077,N_3782,N_3962);
nor U4078 (N_4078,N_3812,N_3960);
and U4079 (N_4079,N_3757,N_3795);
nor U4080 (N_4080,N_3789,N_3763);
or U4081 (N_4081,N_3943,N_3892);
and U4082 (N_4082,N_3989,N_3887);
or U4083 (N_4083,N_3944,N_3815);
nor U4084 (N_4084,N_3783,N_3818);
or U4085 (N_4085,N_3813,N_3941);
and U4086 (N_4086,N_3987,N_3846);
xnor U4087 (N_4087,N_3771,N_3923);
or U4088 (N_4088,N_3981,N_3967);
and U4089 (N_4089,N_3888,N_3839);
nor U4090 (N_4090,N_3758,N_3858);
nand U4091 (N_4091,N_3752,N_3874);
or U4092 (N_4092,N_3764,N_3849);
xor U4093 (N_4093,N_3853,N_3959);
nor U4094 (N_4094,N_3826,N_3938);
nand U4095 (N_4095,N_3844,N_3884);
nor U4096 (N_4096,N_3845,N_3930);
xnor U4097 (N_4097,N_3766,N_3886);
nand U4098 (N_4098,N_3880,N_3901);
or U4099 (N_4099,N_3805,N_3765);
nor U4100 (N_4100,N_3832,N_3866);
nand U4101 (N_4101,N_3755,N_3878);
xnor U4102 (N_4102,N_3957,N_3997);
nor U4103 (N_4103,N_3859,N_3983);
nor U4104 (N_4104,N_3895,N_3903);
or U4105 (N_4105,N_3833,N_3940);
and U4106 (N_4106,N_3946,N_3837);
and U4107 (N_4107,N_3912,N_3835);
nor U4108 (N_4108,N_3767,N_3830);
and U4109 (N_4109,N_3836,N_3843);
and U4110 (N_4110,N_3754,N_3768);
xor U4111 (N_4111,N_3975,N_3991);
and U4112 (N_4112,N_3852,N_3968);
and U4113 (N_4113,N_3982,N_3966);
or U4114 (N_4114,N_3926,N_3963);
and U4115 (N_4115,N_3971,N_3985);
nor U4116 (N_4116,N_3931,N_3825);
or U4117 (N_4117,N_3777,N_3902);
or U4118 (N_4118,N_3770,N_3910);
xnor U4119 (N_4119,N_3945,N_3949);
or U4120 (N_4120,N_3802,N_3951);
xor U4121 (N_4121,N_3861,N_3875);
or U4122 (N_4122,N_3925,N_3909);
xor U4123 (N_4123,N_3927,N_3916);
nand U4124 (N_4124,N_3753,N_3867);
nor U4125 (N_4125,N_3806,N_3986);
or U4126 (N_4126,N_3886,N_3945);
xor U4127 (N_4127,N_3985,N_3811);
xnor U4128 (N_4128,N_3823,N_3780);
or U4129 (N_4129,N_3775,N_3843);
nand U4130 (N_4130,N_3874,N_3852);
nand U4131 (N_4131,N_3885,N_3798);
or U4132 (N_4132,N_3999,N_3952);
and U4133 (N_4133,N_3812,N_3770);
nor U4134 (N_4134,N_3934,N_3917);
and U4135 (N_4135,N_3962,N_3986);
nand U4136 (N_4136,N_3797,N_3898);
xnor U4137 (N_4137,N_3973,N_3925);
nand U4138 (N_4138,N_3793,N_3897);
and U4139 (N_4139,N_3868,N_3970);
and U4140 (N_4140,N_3816,N_3999);
and U4141 (N_4141,N_3893,N_3822);
nor U4142 (N_4142,N_3889,N_3969);
or U4143 (N_4143,N_3835,N_3910);
or U4144 (N_4144,N_3889,N_3893);
or U4145 (N_4145,N_3835,N_3802);
and U4146 (N_4146,N_3764,N_3797);
nor U4147 (N_4147,N_3839,N_3822);
nor U4148 (N_4148,N_3890,N_3760);
xor U4149 (N_4149,N_3814,N_3763);
xnor U4150 (N_4150,N_3774,N_3824);
or U4151 (N_4151,N_3787,N_3891);
and U4152 (N_4152,N_3765,N_3999);
xnor U4153 (N_4153,N_3998,N_3886);
and U4154 (N_4154,N_3998,N_3925);
nand U4155 (N_4155,N_3942,N_3980);
or U4156 (N_4156,N_3750,N_3811);
or U4157 (N_4157,N_3909,N_3962);
or U4158 (N_4158,N_3916,N_3995);
and U4159 (N_4159,N_3894,N_3791);
and U4160 (N_4160,N_3830,N_3955);
and U4161 (N_4161,N_3916,N_3810);
or U4162 (N_4162,N_3801,N_3983);
nand U4163 (N_4163,N_3859,N_3927);
xnor U4164 (N_4164,N_3752,N_3953);
nor U4165 (N_4165,N_3769,N_3761);
nand U4166 (N_4166,N_3943,N_3995);
nand U4167 (N_4167,N_3977,N_3826);
nand U4168 (N_4168,N_3923,N_3764);
and U4169 (N_4169,N_3810,N_3801);
nor U4170 (N_4170,N_3786,N_3792);
xor U4171 (N_4171,N_3758,N_3951);
or U4172 (N_4172,N_3764,N_3759);
nor U4173 (N_4173,N_3920,N_3951);
xnor U4174 (N_4174,N_3855,N_3986);
nand U4175 (N_4175,N_3930,N_3995);
nor U4176 (N_4176,N_3992,N_3789);
nor U4177 (N_4177,N_3766,N_3838);
or U4178 (N_4178,N_3935,N_3906);
nand U4179 (N_4179,N_3926,N_3989);
and U4180 (N_4180,N_3861,N_3908);
xnor U4181 (N_4181,N_3857,N_3836);
nand U4182 (N_4182,N_3846,N_3810);
xor U4183 (N_4183,N_3923,N_3922);
xnor U4184 (N_4184,N_3985,N_3795);
or U4185 (N_4185,N_3958,N_3822);
xnor U4186 (N_4186,N_3911,N_3968);
xnor U4187 (N_4187,N_3882,N_3964);
or U4188 (N_4188,N_3953,N_3954);
nor U4189 (N_4189,N_3972,N_3783);
nand U4190 (N_4190,N_3778,N_3795);
nand U4191 (N_4191,N_3825,N_3862);
xnor U4192 (N_4192,N_3968,N_3945);
and U4193 (N_4193,N_3879,N_3935);
xnor U4194 (N_4194,N_3840,N_3809);
or U4195 (N_4195,N_3984,N_3834);
nor U4196 (N_4196,N_3944,N_3910);
and U4197 (N_4197,N_3783,N_3854);
and U4198 (N_4198,N_3838,N_3865);
or U4199 (N_4199,N_3833,N_3861);
and U4200 (N_4200,N_3760,N_3819);
or U4201 (N_4201,N_3989,N_3993);
xor U4202 (N_4202,N_3888,N_3809);
and U4203 (N_4203,N_3957,N_3771);
and U4204 (N_4204,N_3959,N_3813);
nor U4205 (N_4205,N_3950,N_3767);
nand U4206 (N_4206,N_3817,N_3879);
nand U4207 (N_4207,N_3859,N_3900);
xnor U4208 (N_4208,N_3785,N_3764);
nor U4209 (N_4209,N_3986,N_3960);
xor U4210 (N_4210,N_3770,N_3793);
nand U4211 (N_4211,N_3967,N_3945);
nor U4212 (N_4212,N_3857,N_3870);
xor U4213 (N_4213,N_3803,N_3849);
nor U4214 (N_4214,N_3897,N_3964);
xor U4215 (N_4215,N_3899,N_3757);
or U4216 (N_4216,N_3939,N_3812);
or U4217 (N_4217,N_3781,N_3984);
or U4218 (N_4218,N_3941,N_3863);
nor U4219 (N_4219,N_3765,N_3919);
nor U4220 (N_4220,N_3998,N_3895);
or U4221 (N_4221,N_3820,N_3934);
or U4222 (N_4222,N_3918,N_3958);
nand U4223 (N_4223,N_3917,N_3827);
or U4224 (N_4224,N_3843,N_3996);
nand U4225 (N_4225,N_3857,N_3804);
xnor U4226 (N_4226,N_3835,N_3804);
nor U4227 (N_4227,N_3925,N_3912);
nand U4228 (N_4228,N_3923,N_3867);
nand U4229 (N_4229,N_3902,N_3947);
and U4230 (N_4230,N_3919,N_3917);
xnor U4231 (N_4231,N_3787,N_3947);
nor U4232 (N_4232,N_3798,N_3970);
nand U4233 (N_4233,N_3815,N_3779);
and U4234 (N_4234,N_3872,N_3762);
nand U4235 (N_4235,N_3925,N_3954);
nor U4236 (N_4236,N_3831,N_3842);
xor U4237 (N_4237,N_3893,N_3899);
xor U4238 (N_4238,N_3826,N_3945);
xnor U4239 (N_4239,N_3983,N_3912);
and U4240 (N_4240,N_3920,N_3808);
xor U4241 (N_4241,N_3750,N_3988);
and U4242 (N_4242,N_3789,N_3926);
nand U4243 (N_4243,N_3769,N_3886);
nand U4244 (N_4244,N_3861,N_3877);
or U4245 (N_4245,N_3757,N_3814);
nand U4246 (N_4246,N_3941,N_3750);
nand U4247 (N_4247,N_3897,N_3903);
or U4248 (N_4248,N_3947,N_3755);
or U4249 (N_4249,N_3766,N_3919);
or U4250 (N_4250,N_4040,N_4010);
xnor U4251 (N_4251,N_4129,N_4210);
nor U4252 (N_4252,N_4008,N_4224);
or U4253 (N_4253,N_4054,N_4045);
and U4254 (N_4254,N_4028,N_4220);
nor U4255 (N_4255,N_4149,N_4241);
xor U4256 (N_4256,N_4061,N_4070);
nor U4257 (N_4257,N_4099,N_4094);
and U4258 (N_4258,N_4147,N_4193);
xnor U4259 (N_4259,N_4090,N_4237);
nand U4260 (N_4260,N_4156,N_4022);
and U4261 (N_4261,N_4135,N_4113);
nor U4262 (N_4262,N_4198,N_4199);
and U4263 (N_4263,N_4244,N_4080);
nand U4264 (N_4264,N_4053,N_4180);
xnor U4265 (N_4265,N_4165,N_4043);
or U4266 (N_4266,N_4005,N_4068);
nor U4267 (N_4267,N_4013,N_4071);
and U4268 (N_4268,N_4153,N_4195);
nor U4269 (N_4269,N_4222,N_4118);
xor U4270 (N_4270,N_4171,N_4213);
xnor U4271 (N_4271,N_4027,N_4229);
or U4272 (N_4272,N_4228,N_4137);
nor U4273 (N_4273,N_4182,N_4212);
nand U4274 (N_4274,N_4217,N_4073);
or U4275 (N_4275,N_4009,N_4203);
nor U4276 (N_4276,N_4082,N_4218);
nor U4277 (N_4277,N_4230,N_4020);
xor U4278 (N_4278,N_4015,N_4187);
and U4279 (N_4279,N_4100,N_4109);
xnor U4280 (N_4280,N_4007,N_4000);
xnor U4281 (N_4281,N_4246,N_4078);
or U4282 (N_4282,N_4160,N_4112);
xnor U4283 (N_4283,N_4023,N_4108);
and U4284 (N_4284,N_4125,N_4041);
xor U4285 (N_4285,N_4170,N_4235);
nor U4286 (N_4286,N_4231,N_4056);
or U4287 (N_4287,N_4039,N_4117);
nand U4288 (N_4288,N_4166,N_4225);
and U4289 (N_4289,N_4163,N_4106);
nand U4290 (N_4290,N_4038,N_4092);
or U4291 (N_4291,N_4243,N_4131);
nor U4292 (N_4292,N_4001,N_4143);
nor U4293 (N_4293,N_4204,N_4034);
xor U4294 (N_4294,N_4223,N_4173);
or U4295 (N_4295,N_4191,N_4064);
nand U4296 (N_4296,N_4240,N_4035);
xnor U4297 (N_4297,N_4029,N_4002);
nor U4298 (N_4298,N_4144,N_4055);
nor U4299 (N_4299,N_4037,N_4105);
nor U4300 (N_4300,N_4164,N_4026);
and U4301 (N_4301,N_4172,N_4036);
and U4302 (N_4302,N_4159,N_4024);
nor U4303 (N_4303,N_4111,N_4183);
xor U4304 (N_4304,N_4091,N_4248);
and U4305 (N_4305,N_4067,N_4018);
nor U4306 (N_4306,N_4192,N_4057);
nand U4307 (N_4307,N_4233,N_4221);
nor U4308 (N_4308,N_4211,N_4148);
and U4309 (N_4309,N_4059,N_4161);
xnor U4310 (N_4310,N_4033,N_4088);
nor U4311 (N_4311,N_4158,N_4044);
xor U4312 (N_4312,N_4104,N_4145);
or U4313 (N_4313,N_4123,N_4115);
nand U4314 (N_4314,N_4150,N_4048);
xnor U4315 (N_4315,N_4077,N_4107);
xnor U4316 (N_4316,N_4157,N_4152);
and U4317 (N_4317,N_4179,N_4176);
xor U4318 (N_4318,N_4174,N_4087);
nand U4319 (N_4319,N_4114,N_4049);
and U4320 (N_4320,N_4184,N_4169);
or U4321 (N_4321,N_4216,N_4134);
and U4322 (N_4322,N_4102,N_4019);
nand U4323 (N_4323,N_4226,N_4011);
and U4324 (N_4324,N_4079,N_4101);
xnor U4325 (N_4325,N_4074,N_4093);
nor U4326 (N_4326,N_4188,N_4146);
xor U4327 (N_4327,N_4081,N_4052);
and U4328 (N_4328,N_4083,N_4050);
xnor U4329 (N_4329,N_4249,N_4234);
nor U4330 (N_4330,N_4089,N_4168);
or U4331 (N_4331,N_4215,N_4151);
nor U4332 (N_4332,N_4051,N_4116);
nand U4333 (N_4333,N_4096,N_4095);
xor U4334 (N_4334,N_4245,N_4127);
and U4335 (N_4335,N_4030,N_4058);
nand U4336 (N_4336,N_4232,N_4194);
or U4337 (N_4337,N_4136,N_4017);
or U4338 (N_4338,N_4097,N_4242);
nor U4339 (N_4339,N_4196,N_4181);
and U4340 (N_4340,N_4167,N_4130);
or U4341 (N_4341,N_4065,N_4025);
or U4342 (N_4342,N_4206,N_4086);
nor U4343 (N_4343,N_4205,N_4154);
xor U4344 (N_4344,N_4060,N_4006);
or U4345 (N_4345,N_4124,N_4012);
xnor U4346 (N_4346,N_4247,N_4128);
and U4347 (N_4347,N_4133,N_4139);
nor U4348 (N_4348,N_4142,N_4084);
xnor U4349 (N_4349,N_4076,N_4103);
nor U4350 (N_4350,N_4072,N_4214);
xnor U4351 (N_4351,N_4200,N_4162);
and U4352 (N_4352,N_4069,N_4032);
nand U4353 (N_4353,N_4236,N_4021);
nand U4354 (N_4354,N_4042,N_4140);
and U4355 (N_4355,N_4178,N_4132);
or U4356 (N_4356,N_4141,N_4122);
nand U4357 (N_4357,N_4201,N_4075);
nor U4358 (N_4358,N_4177,N_4085);
or U4359 (N_4359,N_4126,N_4155);
nand U4360 (N_4360,N_4031,N_4003);
xnor U4361 (N_4361,N_4138,N_4016);
and U4362 (N_4362,N_4066,N_4098);
nor U4363 (N_4363,N_4227,N_4046);
xnor U4364 (N_4364,N_4189,N_4110);
xnor U4365 (N_4365,N_4185,N_4239);
xnor U4366 (N_4366,N_4119,N_4186);
or U4367 (N_4367,N_4238,N_4121);
nor U4368 (N_4368,N_4063,N_4202);
xnor U4369 (N_4369,N_4219,N_4209);
nor U4370 (N_4370,N_4207,N_4004);
nand U4371 (N_4371,N_4062,N_4014);
and U4372 (N_4372,N_4190,N_4197);
and U4373 (N_4373,N_4047,N_4175);
and U4374 (N_4374,N_4120,N_4208);
or U4375 (N_4375,N_4027,N_4043);
xnor U4376 (N_4376,N_4222,N_4201);
and U4377 (N_4377,N_4213,N_4055);
or U4378 (N_4378,N_4134,N_4071);
and U4379 (N_4379,N_4187,N_4083);
or U4380 (N_4380,N_4161,N_4155);
or U4381 (N_4381,N_4123,N_4236);
nor U4382 (N_4382,N_4176,N_4172);
and U4383 (N_4383,N_4161,N_4197);
or U4384 (N_4384,N_4140,N_4127);
xor U4385 (N_4385,N_4141,N_4174);
nor U4386 (N_4386,N_4064,N_4215);
xnor U4387 (N_4387,N_4058,N_4150);
xor U4388 (N_4388,N_4119,N_4242);
xnor U4389 (N_4389,N_4057,N_4000);
xor U4390 (N_4390,N_4073,N_4046);
or U4391 (N_4391,N_4238,N_4175);
and U4392 (N_4392,N_4024,N_4030);
xnor U4393 (N_4393,N_4093,N_4002);
nor U4394 (N_4394,N_4071,N_4103);
xor U4395 (N_4395,N_4245,N_4208);
nor U4396 (N_4396,N_4128,N_4214);
nor U4397 (N_4397,N_4144,N_4008);
nor U4398 (N_4398,N_4167,N_4218);
nand U4399 (N_4399,N_4198,N_4228);
nor U4400 (N_4400,N_4041,N_4069);
nand U4401 (N_4401,N_4159,N_4226);
xor U4402 (N_4402,N_4167,N_4017);
nand U4403 (N_4403,N_4092,N_4110);
or U4404 (N_4404,N_4185,N_4170);
nand U4405 (N_4405,N_4235,N_4030);
and U4406 (N_4406,N_4226,N_4126);
xor U4407 (N_4407,N_4083,N_4220);
nand U4408 (N_4408,N_4189,N_4197);
nor U4409 (N_4409,N_4211,N_4048);
and U4410 (N_4410,N_4024,N_4057);
and U4411 (N_4411,N_4024,N_4098);
or U4412 (N_4412,N_4185,N_4207);
or U4413 (N_4413,N_4068,N_4201);
xor U4414 (N_4414,N_4156,N_4098);
nand U4415 (N_4415,N_4075,N_4094);
or U4416 (N_4416,N_4055,N_4238);
or U4417 (N_4417,N_4022,N_4240);
or U4418 (N_4418,N_4080,N_4099);
nor U4419 (N_4419,N_4226,N_4070);
or U4420 (N_4420,N_4120,N_4154);
nor U4421 (N_4421,N_4104,N_4135);
nand U4422 (N_4422,N_4203,N_4218);
or U4423 (N_4423,N_4128,N_4145);
xor U4424 (N_4424,N_4076,N_4048);
nor U4425 (N_4425,N_4201,N_4007);
xor U4426 (N_4426,N_4068,N_4138);
and U4427 (N_4427,N_4196,N_4122);
and U4428 (N_4428,N_4016,N_4092);
nor U4429 (N_4429,N_4202,N_4164);
nand U4430 (N_4430,N_4118,N_4142);
xor U4431 (N_4431,N_4225,N_4092);
or U4432 (N_4432,N_4138,N_4184);
nand U4433 (N_4433,N_4173,N_4236);
xnor U4434 (N_4434,N_4232,N_4104);
nor U4435 (N_4435,N_4160,N_4085);
or U4436 (N_4436,N_4118,N_4214);
nor U4437 (N_4437,N_4076,N_4204);
nand U4438 (N_4438,N_4127,N_4191);
nor U4439 (N_4439,N_4061,N_4130);
nand U4440 (N_4440,N_4161,N_4095);
and U4441 (N_4441,N_4021,N_4031);
and U4442 (N_4442,N_4014,N_4079);
nor U4443 (N_4443,N_4110,N_4100);
or U4444 (N_4444,N_4120,N_4219);
xor U4445 (N_4445,N_4083,N_4079);
nor U4446 (N_4446,N_4231,N_4057);
nor U4447 (N_4447,N_4023,N_4185);
nor U4448 (N_4448,N_4179,N_4215);
or U4449 (N_4449,N_4053,N_4070);
xor U4450 (N_4450,N_4211,N_4030);
xnor U4451 (N_4451,N_4030,N_4206);
nand U4452 (N_4452,N_4166,N_4057);
or U4453 (N_4453,N_4068,N_4008);
and U4454 (N_4454,N_4146,N_4147);
and U4455 (N_4455,N_4080,N_4157);
xor U4456 (N_4456,N_4134,N_4057);
xnor U4457 (N_4457,N_4194,N_4119);
nor U4458 (N_4458,N_4008,N_4221);
xor U4459 (N_4459,N_4234,N_4165);
nor U4460 (N_4460,N_4235,N_4075);
nor U4461 (N_4461,N_4234,N_4128);
or U4462 (N_4462,N_4212,N_4028);
nand U4463 (N_4463,N_4093,N_4212);
and U4464 (N_4464,N_4135,N_4221);
nand U4465 (N_4465,N_4202,N_4207);
or U4466 (N_4466,N_4128,N_4115);
and U4467 (N_4467,N_4057,N_4033);
and U4468 (N_4468,N_4190,N_4224);
nand U4469 (N_4469,N_4211,N_4107);
xnor U4470 (N_4470,N_4019,N_4169);
or U4471 (N_4471,N_4022,N_4160);
nand U4472 (N_4472,N_4081,N_4223);
nand U4473 (N_4473,N_4095,N_4166);
xor U4474 (N_4474,N_4110,N_4059);
or U4475 (N_4475,N_4246,N_4127);
xnor U4476 (N_4476,N_4237,N_4157);
xnor U4477 (N_4477,N_4086,N_4228);
xor U4478 (N_4478,N_4188,N_4189);
nor U4479 (N_4479,N_4202,N_4009);
xnor U4480 (N_4480,N_4106,N_4111);
and U4481 (N_4481,N_4082,N_4048);
xnor U4482 (N_4482,N_4034,N_4217);
xor U4483 (N_4483,N_4118,N_4098);
nand U4484 (N_4484,N_4198,N_4033);
nor U4485 (N_4485,N_4062,N_4227);
or U4486 (N_4486,N_4235,N_4139);
xor U4487 (N_4487,N_4054,N_4090);
xor U4488 (N_4488,N_4221,N_4239);
nor U4489 (N_4489,N_4173,N_4129);
nor U4490 (N_4490,N_4092,N_4099);
nor U4491 (N_4491,N_4047,N_4153);
or U4492 (N_4492,N_4153,N_4220);
xor U4493 (N_4493,N_4056,N_4141);
or U4494 (N_4494,N_4102,N_4096);
or U4495 (N_4495,N_4056,N_4022);
and U4496 (N_4496,N_4201,N_4096);
xnor U4497 (N_4497,N_4164,N_4065);
nor U4498 (N_4498,N_4247,N_4189);
or U4499 (N_4499,N_4046,N_4044);
nor U4500 (N_4500,N_4416,N_4282);
nand U4501 (N_4501,N_4346,N_4273);
nand U4502 (N_4502,N_4414,N_4478);
nand U4503 (N_4503,N_4355,N_4340);
and U4504 (N_4504,N_4314,N_4260);
xor U4505 (N_4505,N_4253,N_4426);
xor U4506 (N_4506,N_4250,N_4387);
xnor U4507 (N_4507,N_4358,N_4392);
xnor U4508 (N_4508,N_4263,N_4373);
or U4509 (N_4509,N_4278,N_4337);
xnor U4510 (N_4510,N_4378,N_4393);
and U4511 (N_4511,N_4388,N_4305);
xor U4512 (N_4512,N_4413,N_4298);
xor U4513 (N_4513,N_4476,N_4284);
nand U4514 (N_4514,N_4364,N_4334);
nand U4515 (N_4515,N_4315,N_4394);
or U4516 (N_4516,N_4446,N_4437);
or U4517 (N_4517,N_4385,N_4348);
nand U4518 (N_4518,N_4482,N_4408);
nor U4519 (N_4519,N_4429,N_4491);
xor U4520 (N_4520,N_4493,N_4331);
and U4521 (N_4521,N_4397,N_4275);
and U4522 (N_4522,N_4400,N_4359);
nor U4523 (N_4523,N_4494,N_4308);
and U4524 (N_4524,N_4262,N_4329);
xnor U4525 (N_4525,N_4288,N_4422);
xor U4526 (N_4526,N_4454,N_4440);
or U4527 (N_4527,N_4402,N_4318);
and U4528 (N_4528,N_4445,N_4498);
and U4529 (N_4529,N_4432,N_4285);
nor U4530 (N_4530,N_4450,N_4370);
nand U4531 (N_4531,N_4291,N_4431);
nor U4532 (N_4532,N_4274,N_4424);
nand U4533 (N_4533,N_4404,N_4295);
and U4534 (N_4534,N_4490,N_4276);
xor U4535 (N_4535,N_4347,N_4470);
or U4536 (N_4536,N_4419,N_4286);
and U4537 (N_4537,N_4354,N_4384);
nor U4538 (N_4538,N_4409,N_4495);
xnor U4539 (N_4539,N_4390,N_4254);
or U4540 (N_4540,N_4336,N_4433);
nor U4541 (N_4541,N_4366,N_4327);
nor U4542 (N_4542,N_4447,N_4303);
nor U4543 (N_4543,N_4463,N_4255);
and U4544 (N_4544,N_4441,N_4391);
nor U4545 (N_4545,N_4398,N_4389);
nand U4546 (N_4546,N_4386,N_4496);
and U4547 (N_4547,N_4466,N_4427);
or U4548 (N_4548,N_4425,N_4335);
and U4549 (N_4549,N_4372,N_4434);
or U4550 (N_4550,N_4452,N_4383);
nor U4551 (N_4551,N_4451,N_4328);
or U4552 (N_4552,N_4251,N_4479);
xnor U4553 (N_4553,N_4266,N_4483);
and U4554 (N_4554,N_4380,N_4277);
xnor U4555 (N_4555,N_4339,N_4345);
nand U4556 (N_4556,N_4330,N_4369);
nand U4557 (N_4557,N_4350,N_4297);
or U4558 (N_4558,N_4306,N_4343);
xnor U4559 (N_4559,N_4455,N_4472);
or U4560 (N_4560,N_4351,N_4267);
nor U4561 (N_4561,N_4468,N_4459);
xor U4562 (N_4562,N_4406,N_4293);
nor U4563 (N_4563,N_4417,N_4368);
nor U4564 (N_4564,N_4428,N_4499);
nand U4565 (N_4565,N_4280,N_4311);
or U4566 (N_4566,N_4279,N_4294);
xor U4567 (N_4567,N_4289,N_4471);
nor U4568 (N_4568,N_4264,N_4377);
xor U4569 (N_4569,N_4310,N_4415);
nor U4570 (N_4570,N_4489,N_4460);
nor U4571 (N_4571,N_4480,N_4321);
nor U4572 (N_4572,N_4258,N_4395);
nor U4573 (N_4573,N_4362,N_4283);
or U4574 (N_4574,N_4448,N_4497);
nor U4575 (N_4575,N_4265,N_4312);
xor U4576 (N_4576,N_4486,N_4271);
or U4577 (N_4577,N_4325,N_4317);
and U4578 (N_4578,N_4256,N_4443);
nor U4579 (N_4579,N_4374,N_4412);
nand U4580 (N_4580,N_4464,N_4323);
or U4581 (N_4581,N_4473,N_4461);
or U4582 (N_4582,N_4367,N_4469);
xor U4583 (N_4583,N_4444,N_4281);
and U4584 (N_4584,N_4488,N_4322);
xor U4585 (N_4585,N_4423,N_4300);
nor U4586 (N_4586,N_4487,N_4467);
xor U4587 (N_4587,N_4379,N_4403);
xnor U4588 (N_4588,N_4360,N_4357);
nor U4589 (N_4589,N_4309,N_4349);
or U4590 (N_4590,N_4361,N_4257);
xnor U4591 (N_4591,N_4338,N_4333);
nand U4592 (N_4592,N_4324,N_4439);
nor U4593 (N_4593,N_4405,N_4287);
nor U4594 (N_4594,N_4481,N_4363);
xor U4595 (N_4595,N_4352,N_4457);
and U4596 (N_4596,N_4353,N_4465);
and U4597 (N_4597,N_4484,N_4420);
xnor U4598 (N_4598,N_4319,N_4401);
and U4599 (N_4599,N_4410,N_4301);
nor U4600 (N_4600,N_4399,N_4302);
nand U4601 (N_4601,N_4252,N_4332);
or U4602 (N_4602,N_4299,N_4269);
nand U4603 (N_4603,N_4304,N_4436);
nor U4604 (N_4604,N_4296,N_4356);
or U4605 (N_4605,N_4365,N_4326);
and U4606 (N_4606,N_4259,N_4442);
xor U4607 (N_4607,N_4492,N_4477);
and U4608 (N_4608,N_4292,N_4396);
xor U4609 (N_4609,N_4435,N_4270);
nor U4610 (N_4610,N_4456,N_4313);
xnor U4611 (N_4611,N_4342,N_4316);
and U4612 (N_4612,N_4449,N_4407);
nand U4613 (N_4613,N_4268,N_4418);
and U4614 (N_4614,N_4290,N_4376);
or U4615 (N_4615,N_4462,N_4411);
nand U4616 (N_4616,N_4382,N_4261);
nand U4617 (N_4617,N_4272,N_4430);
or U4618 (N_4618,N_4438,N_4421);
nand U4619 (N_4619,N_4458,N_4485);
xnor U4620 (N_4620,N_4375,N_4341);
and U4621 (N_4621,N_4474,N_4307);
xnor U4622 (N_4622,N_4381,N_4453);
nor U4623 (N_4623,N_4320,N_4371);
nand U4624 (N_4624,N_4475,N_4344);
or U4625 (N_4625,N_4472,N_4343);
and U4626 (N_4626,N_4353,N_4410);
or U4627 (N_4627,N_4432,N_4287);
xnor U4628 (N_4628,N_4460,N_4307);
xor U4629 (N_4629,N_4379,N_4274);
or U4630 (N_4630,N_4409,N_4340);
nand U4631 (N_4631,N_4351,N_4337);
xor U4632 (N_4632,N_4285,N_4450);
nand U4633 (N_4633,N_4380,N_4285);
nor U4634 (N_4634,N_4462,N_4331);
or U4635 (N_4635,N_4384,N_4360);
nor U4636 (N_4636,N_4484,N_4488);
or U4637 (N_4637,N_4447,N_4483);
or U4638 (N_4638,N_4491,N_4316);
or U4639 (N_4639,N_4263,N_4349);
nor U4640 (N_4640,N_4473,N_4460);
or U4641 (N_4641,N_4318,N_4322);
xnor U4642 (N_4642,N_4267,N_4405);
xor U4643 (N_4643,N_4443,N_4497);
xnor U4644 (N_4644,N_4434,N_4404);
nand U4645 (N_4645,N_4293,N_4278);
and U4646 (N_4646,N_4405,N_4473);
and U4647 (N_4647,N_4317,N_4405);
and U4648 (N_4648,N_4259,N_4303);
nor U4649 (N_4649,N_4456,N_4453);
xor U4650 (N_4650,N_4386,N_4419);
or U4651 (N_4651,N_4277,N_4306);
nand U4652 (N_4652,N_4394,N_4366);
and U4653 (N_4653,N_4277,N_4299);
nand U4654 (N_4654,N_4311,N_4386);
nand U4655 (N_4655,N_4492,N_4330);
nor U4656 (N_4656,N_4419,N_4495);
nand U4657 (N_4657,N_4349,N_4405);
and U4658 (N_4658,N_4354,N_4476);
nand U4659 (N_4659,N_4491,N_4394);
or U4660 (N_4660,N_4306,N_4370);
nor U4661 (N_4661,N_4404,N_4472);
nor U4662 (N_4662,N_4298,N_4418);
and U4663 (N_4663,N_4478,N_4320);
xnor U4664 (N_4664,N_4414,N_4374);
or U4665 (N_4665,N_4270,N_4309);
and U4666 (N_4666,N_4472,N_4325);
nand U4667 (N_4667,N_4368,N_4273);
nor U4668 (N_4668,N_4436,N_4496);
xor U4669 (N_4669,N_4462,N_4421);
nor U4670 (N_4670,N_4368,N_4405);
or U4671 (N_4671,N_4305,N_4335);
or U4672 (N_4672,N_4480,N_4415);
xor U4673 (N_4673,N_4436,N_4307);
nand U4674 (N_4674,N_4262,N_4393);
nand U4675 (N_4675,N_4285,N_4358);
nand U4676 (N_4676,N_4457,N_4362);
xor U4677 (N_4677,N_4411,N_4340);
nor U4678 (N_4678,N_4405,N_4378);
and U4679 (N_4679,N_4419,N_4474);
or U4680 (N_4680,N_4438,N_4487);
xor U4681 (N_4681,N_4499,N_4436);
nor U4682 (N_4682,N_4276,N_4333);
nor U4683 (N_4683,N_4380,N_4341);
nand U4684 (N_4684,N_4315,N_4471);
nor U4685 (N_4685,N_4424,N_4402);
and U4686 (N_4686,N_4493,N_4349);
nor U4687 (N_4687,N_4271,N_4479);
or U4688 (N_4688,N_4412,N_4465);
nor U4689 (N_4689,N_4403,N_4365);
xnor U4690 (N_4690,N_4352,N_4344);
nor U4691 (N_4691,N_4308,N_4261);
nand U4692 (N_4692,N_4264,N_4382);
or U4693 (N_4693,N_4350,N_4395);
nand U4694 (N_4694,N_4395,N_4308);
and U4695 (N_4695,N_4444,N_4337);
or U4696 (N_4696,N_4287,N_4378);
nand U4697 (N_4697,N_4320,N_4414);
and U4698 (N_4698,N_4303,N_4398);
nor U4699 (N_4699,N_4305,N_4339);
and U4700 (N_4700,N_4413,N_4338);
nand U4701 (N_4701,N_4396,N_4451);
nor U4702 (N_4702,N_4444,N_4493);
or U4703 (N_4703,N_4423,N_4310);
and U4704 (N_4704,N_4356,N_4438);
and U4705 (N_4705,N_4339,N_4344);
nor U4706 (N_4706,N_4496,N_4465);
and U4707 (N_4707,N_4486,N_4335);
nand U4708 (N_4708,N_4451,N_4437);
or U4709 (N_4709,N_4420,N_4482);
nand U4710 (N_4710,N_4426,N_4413);
and U4711 (N_4711,N_4425,N_4413);
and U4712 (N_4712,N_4427,N_4330);
nor U4713 (N_4713,N_4405,N_4347);
xnor U4714 (N_4714,N_4457,N_4285);
nor U4715 (N_4715,N_4465,N_4345);
nor U4716 (N_4716,N_4347,N_4300);
and U4717 (N_4717,N_4287,N_4465);
xnor U4718 (N_4718,N_4424,N_4450);
xnor U4719 (N_4719,N_4255,N_4471);
or U4720 (N_4720,N_4338,N_4271);
nand U4721 (N_4721,N_4257,N_4377);
nor U4722 (N_4722,N_4294,N_4328);
xor U4723 (N_4723,N_4333,N_4450);
or U4724 (N_4724,N_4262,N_4274);
nand U4725 (N_4725,N_4370,N_4452);
nor U4726 (N_4726,N_4334,N_4363);
and U4727 (N_4727,N_4403,N_4482);
nor U4728 (N_4728,N_4341,N_4289);
and U4729 (N_4729,N_4256,N_4301);
and U4730 (N_4730,N_4330,N_4253);
nor U4731 (N_4731,N_4282,N_4347);
xnor U4732 (N_4732,N_4393,N_4358);
and U4733 (N_4733,N_4385,N_4497);
and U4734 (N_4734,N_4489,N_4476);
xor U4735 (N_4735,N_4327,N_4411);
or U4736 (N_4736,N_4455,N_4449);
or U4737 (N_4737,N_4405,N_4357);
and U4738 (N_4738,N_4393,N_4426);
nand U4739 (N_4739,N_4375,N_4317);
nor U4740 (N_4740,N_4461,N_4440);
and U4741 (N_4741,N_4364,N_4269);
or U4742 (N_4742,N_4278,N_4327);
xor U4743 (N_4743,N_4320,N_4285);
xor U4744 (N_4744,N_4373,N_4295);
nand U4745 (N_4745,N_4486,N_4438);
or U4746 (N_4746,N_4431,N_4387);
and U4747 (N_4747,N_4486,N_4326);
or U4748 (N_4748,N_4456,N_4250);
and U4749 (N_4749,N_4480,N_4345);
xnor U4750 (N_4750,N_4736,N_4590);
xnor U4751 (N_4751,N_4749,N_4582);
xnor U4752 (N_4752,N_4622,N_4666);
and U4753 (N_4753,N_4686,N_4656);
and U4754 (N_4754,N_4525,N_4579);
nor U4755 (N_4755,N_4522,N_4673);
or U4756 (N_4756,N_4671,N_4681);
nor U4757 (N_4757,N_4532,N_4564);
or U4758 (N_4758,N_4511,N_4628);
nor U4759 (N_4759,N_4706,N_4743);
xnor U4760 (N_4760,N_4589,N_4549);
nand U4761 (N_4761,N_4542,N_4573);
nor U4762 (N_4762,N_4696,N_4591);
or U4763 (N_4763,N_4701,N_4655);
nand U4764 (N_4764,N_4615,N_4596);
xor U4765 (N_4765,N_4558,N_4657);
nand U4766 (N_4766,N_4592,N_4692);
nor U4767 (N_4767,N_4740,N_4560);
xnor U4768 (N_4768,N_4715,N_4719);
xnor U4769 (N_4769,N_4555,N_4621);
nor U4770 (N_4770,N_4593,N_4746);
xor U4771 (N_4771,N_4711,N_4738);
or U4772 (N_4772,N_4714,N_4517);
nand U4773 (N_4773,N_4665,N_4705);
and U4774 (N_4774,N_4712,N_4587);
xor U4775 (N_4775,N_4627,N_4651);
and U4776 (N_4776,N_4739,N_4570);
xnor U4777 (N_4777,N_4732,N_4648);
xor U4778 (N_4778,N_4562,N_4724);
and U4779 (N_4779,N_4637,N_4616);
or U4780 (N_4780,N_4684,N_4745);
nand U4781 (N_4781,N_4718,N_4513);
nor U4782 (N_4782,N_4641,N_4682);
nand U4783 (N_4783,N_4728,N_4578);
or U4784 (N_4784,N_4584,N_4586);
nor U4785 (N_4785,N_4594,N_4546);
xor U4786 (N_4786,N_4610,N_4623);
nand U4787 (N_4787,N_4703,N_4625);
and U4788 (N_4788,N_4547,N_4672);
or U4789 (N_4789,N_4509,N_4512);
or U4790 (N_4790,N_4653,N_4550);
or U4791 (N_4791,N_4537,N_4722);
nor U4792 (N_4792,N_4548,N_4742);
and U4793 (N_4793,N_4565,N_4646);
nor U4794 (N_4794,N_4519,N_4664);
xor U4795 (N_4795,N_4630,N_4678);
xnor U4796 (N_4796,N_4510,N_4611);
nor U4797 (N_4797,N_4580,N_4563);
nor U4798 (N_4798,N_4620,N_4588);
or U4799 (N_4799,N_4601,N_4649);
and U4800 (N_4800,N_4551,N_4516);
nor U4801 (N_4801,N_4608,N_4571);
nand U4802 (N_4802,N_4605,N_4663);
nand U4803 (N_4803,N_4561,N_4668);
or U4804 (N_4804,N_4635,N_4693);
and U4805 (N_4805,N_4647,N_4652);
xor U4806 (N_4806,N_4502,N_4735);
xnor U4807 (N_4807,N_4528,N_4687);
nand U4808 (N_4808,N_4734,N_4661);
nand U4809 (N_4809,N_4741,N_4520);
or U4810 (N_4810,N_4574,N_4670);
or U4811 (N_4811,N_4527,N_4639);
nor U4812 (N_4812,N_4631,N_4634);
and U4813 (N_4813,N_4675,N_4606);
nor U4814 (N_4814,N_4729,N_4723);
nand U4815 (N_4815,N_4534,N_4521);
nor U4816 (N_4816,N_4538,N_4710);
nand U4817 (N_4817,N_4618,N_4514);
nor U4818 (N_4818,N_4515,N_4748);
and U4819 (N_4819,N_4662,N_4683);
or U4820 (N_4820,N_4613,N_4691);
xor U4821 (N_4821,N_4576,N_4698);
nand U4822 (N_4822,N_4543,N_4599);
or U4823 (N_4823,N_4737,N_4541);
nor U4824 (N_4824,N_4677,N_4626);
and U4825 (N_4825,N_4603,N_4642);
nand U4826 (N_4826,N_4524,N_4636);
nand U4827 (N_4827,N_4733,N_4569);
and U4828 (N_4828,N_4747,N_4685);
or U4829 (N_4829,N_4654,N_4552);
xor U4830 (N_4830,N_4539,N_4650);
nand U4831 (N_4831,N_4544,N_4572);
xor U4832 (N_4832,N_4600,N_4717);
xnor U4833 (N_4833,N_4645,N_4583);
nand U4834 (N_4834,N_4597,N_4531);
xor U4835 (N_4835,N_4501,N_4633);
or U4836 (N_4836,N_4695,N_4533);
nor U4837 (N_4837,N_4730,N_4504);
xnor U4838 (N_4838,N_4659,N_4614);
nand U4839 (N_4839,N_4640,N_4617);
xor U4840 (N_4840,N_4535,N_4523);
nand U4841 (N_4841,N_4667,N_4629);
nor U4842 (N_4842,N_4554,N_4689);
nand U4843 (N_4843,N_4674,N_4721);
xnor U4844 (N_4844,N_4506,N_4553);
nand U4845 (N_4845,N_4720,N_4676);
nor U4846 (N_4846,N_4704,N_4575);
xnor U4847 (N_4847,N_4612,N_4568);
xor U4848 (N_4848,N_4556,N_4503);
nor U4849 (N_4849,N_4581,N_4518);
xnor U4850 (N_4850,N_4660,N_4702);
and U4851 (N_4851,N_4577,N_4744);
xor U4852 (N_4852,N_4540,N_4526);
xor U4853 (N_4853,N_4679,N_4507);
and U4854 (N_4854,N_4658,N_4536);
or U4855 (N_4855,N_4709,N_4725);
xnor U4856 (N_4856,N_4609,N_4713);
xor U4857 (N_4857,N_4731,N_4529);
and U4858 (N_4858,N_4557,N_4566);
xnor U4859 (N_4859,N_4624,N_4595);
and U4860 (N_4860,N_4602,N_4680);
nor U4861 (N_4861,N_4690,N_4559);
nand U4862 (N_4862,N_4726,N_4669);
nor U4863 (N_4863,N_4707,N_4619);
nor U4864 (N_4864,N_4500,N_4643);
or U4865 (N_4865,N_4727,N_4688);
and U4866 (N_4866,N_4697,N_4716);
and U4867 (N_4867,N_4508,N_4604);
nand U4868 (N_4868,N_4530,N_4598);
nor U4869 (N_4869,N_4700,N_4585);
nor U4870 (N_4870,N_4699,N_4567);
and U4871 (N_4871,N_4644,N_4694);
xor U4872 (N_4872,N_4632,N_4638);
and U4873 (N_4873,N_4545,N_4607);
nand U4874 (N_4874,N_4708,N_4505);
nor U4875 (N_4875,N_4672,N_4648);
xor U4876 (N_4876,N_4594,N_4662);
or U4877 (N_4877,N_4698,N_4713);
or U4878 (N_4878,N_4636,N_4713);
nor U4879 (N_4879,N_4584,N_4665);
or U4880 (N_4880,N_4504,N_4523);
nand U4881 (N_4881,N_4600,N_4731);
xnor U4882 (N_4882,N_4581,N_4641);
xor U4883 (N_4883,N_4509,N_4598);
or U4884 (N_4884,N_4733,N_4503);
and U4885 (N_4885,N_4642,N_4607);
nor U4886 (N_4886,N_4723,N_4608);
nand U4887 (N_4887,N_4699,N_4730);
xnor U4888 (N_4888,N_4731,N_4564);
nand U4889 (N_4889,N_4626,N_4548);
xnor U4890 (N_4890,N_4519,N_4564);
nor U4891 (N_4891,N_4584,N_4729);
and U4892 (N_4892,N_4509,N_4734);
and U4893 (N_4893,N_4644,N_4634);
nor U4894 (N_4894,N_4543,N_4630);
nor U4895 (N_4895,N_4645,N_4687);
and U4896 (N_4896,N_4645,N_4740);
xor U4897 (N_4897,N_4700,N_4545);
nand U4898 (N_4898,N_4516,N_4692);
nand U4899 (N_4899,N_4721,N_4706);
nor U4900 (N_4900,N_4737,N_4705);
nand U4901 (N_4901,N_4574,N_4565);
nand U4902 (N_4902,N_4629,N_4704);
nor U4903 (N_4903,N_4604,N_4723);
nand U4904 (N_4904,N_4557,N_4655);
nand U4905 (N_4905,N_4641,N_4738);
nand U4906 (N_4906,N_4630,N_4642);
xnor U4907 (N_4907,N_4721,N_4562);
or U4908 (N_4908,N_4577,N_4670);
or U4909 (N_4909,N_4630,N_4550);
nor U4910 (N_4910,N_4505,N_4715);
nor U4911 (N_4911,N_4721,N_4588);
xor U4912 (N_4912,N_4744,N_4667);
xor U4913 (N_4913,N_4623,N_4594);
xnor U4914 (N_4914,N_4722,N_4682);
xor U4915 (N_4915,N_4708,N_4565);
or U4916 (N_4916,N_4690,N_4552);
and U4917 (N_4917,N_4553,N_4581);
nor U4918 (N_4918,N_4695,N_4666);
nor U4919 (N_4919,N_4552,N_4641);
nand U4920 (N_4920,N_4663,N_4706);
or U4921 (N_4921,N_4734,N_4624);
and U4922 (N_4922,N_4636,N_4548);
or U4923 (N_4923,N_4609,N_4727);
xor U4924 (N_4924,N_4583,N_4517);
and U4925 (N_4925,N_4604,N_4548);
nand U4926 (N_4926,N_4522,N_4510);
and U4927 (N_4927,N_4730,N_4644);
and U4928 (N_4928,N_4669,N_4539);
and U4929 (N_4929,N_4648,N_4736);
nand U4930 (N_4930,N_4689,N_4575);
and U4931 (N_4931,N_4707,N_4582);
xnor U4932 (N_4932,N_4676,N_4574);
nand U4933 (N_4933,N_4704,N_4749);
and U4934 (N_4934,N_4678,N_4590);
nand U4935 (N_4935,N_4713,N_4727);
xnor U4936 (N_4936,N_4523,N_4565);
nor U4937 (N_4937,N_4582,N_4577);
or U4938 (N_4938,N_4509,N_4565);
nor U4939 (N_4939,N_4630,N_4692);
nor U4940 (N_4940,N_4537,N_4598);
nand U4941 (N_4941,N_4686,N_4595);
and U4942 (N_4942,N_4699,N_4643);
or U4943 (N_4943,N_4571,N_4683);
or U4944 (N_4944,N_4668,N_4671);
nor U4945 (N_4945,N_4749,N_4731);
xor U4946 (N_4946,N_4532,N_4606);
nand U4947 (N_4947,N_4652,N_4569);
or U4948 (N_4948,N_4550,N_4508);
and U4949 (N_4949,N_4518,N_4573);
nand U4950 (N_4950,N_4652,N_4702);
nor U4951 (N_4951,N_4712,N_4695);
or U4952 (N_4952,N_4547,N_4600);
or U4953 (N_4953,N_4573,N_4709);
xor U4954 (N_4954,N_4512,N_4735);
or U4955 (N_4955,N_4640,N_4709);
nand U4956 (N_4956,N_4726,N_4705);
or U4957 (N_4957,N_4730,N_4628);
nor U4958 (N_4958,N_4568,N_4566);
nand U4959 (N_4959,N_4594,N_4729);
and U4960 (N_4960,N_4672,N_4581);
or U4961 (N_4961,N_4542,N_4749);
nand U4962 (N_4962,N_4618,N_4672);
xnor U4963 (N_4963,N_4589,N_4632);
or U4964 (N_4964,N_4680,N_4515);
nand U4965 (N_4965,N_4580,N_4643);
or U4966 (N_4966,N_4632,N_4564);
and U4967 (N_4967,N_4510,N_4683);
or U4968 (N_4968,N_4593,N_4731);
and U4969 (N_4969,N_4678,N_4639);
nor U4970 (N_4970,N_4589,N_4717);
nor U4971 (N_4971,N_4574,N_4655);
and U4972 (N_4972,N_4694,N_4584);
and U4973 (N_4973,N_4541,N_4520);
nand U4974 (N_4974,N_4631,N_4668);
and U4975 (N_4975,N_4707,N_4736);
or U4976 (N_4976,N_4663,N_4689);
nor U4977 (N_4977,N_4641,N_4517);
nor U4978 (N_4978,N_4603,N_4554);
xor U4979 (N_4979,N_4523,N_4567);
xnor U4980 (N_4980,N_4539,N_4630);
xnor U4981 (N_4981,N_4546,N_4561);
or U4982 (N_4982,N_4543,N_4617);
or U4983 (N_4983,N_4733,N_4553);
and U4984 (N_4984,N_4587,N_4518);
or U4985 (N_4985,N_4687,N_4509);
or U4986 (N_4986,N_4691,N_4554);
nand U4987 (N_4987,N_4720,N_4633);
xor U4988 (N_4988,N_4614,N_4512);
or U4989 (N_4989,N_4527,N_4712);
or U4990 (N_4990,N_4745,N_4597);
nor U4991 (N_4991,N_4630,N_4693);
nor U4992 (N_4992,N_4620,N_4722);
and U4993 (N_4993,N_4634,N_4601);
nand U4994 (N_4994,N_4657,N_4533);
nor U4995 (N_4995,N_4535,N_4563);
xnor U4996 (N_4996,N_4621,N_4506);
xor U4997 (N_4997,N_4613,N_4672);
nand U4998 (N_4998,N_4597,N_4615);
and U4999 (N_4999,N_4580,N_4628);
xor U5000 (N_5000,N_4818,N_4887);
and U5001 (N_5001,N_4944,N_4976);
or U5002 (N_5002,N_4935,N_4776);
nor U5003 (N_5003,N_4845,N_4751);
nand U5004 (N_5004,N_4847,N_4852);
nand U5005 (N_5005,N_4820,N_4995);
or U5006 (N_5006,N_4987,N_4871);
or U5007 (N_5007,N_4966,N_4898);
and U5008 (N_5008,N_4991,N_4848);
and U5009 (N_5009,N_4901,N_4836);
nand U5010 (N_5010,N_4822,N_4839);
xor U5011 (N_5011,N_4977,N_4816);
nand U5012 (N_5012,N_4921,N_4959);
nor U5013 (N_5013,N_4905,N_4856);
or U5014 (N_5014,N_4910,N_4828);
nor U5015 (N_5015,N_4876,N_4814);
nand U5016 (N_5016,N_4796,N_4780);
nand U5017 (N_5017,N_4834,N_4967);
xor U5018 (N_5018,N_4764,N_4767);
or U5019 (N_5019,N_4992,N_4924);
nand U5020 (N_5020,N_4941,N_4753);
or U5021 (N_5021,N_4855,N_4833);
nor U5022 (N_5022,N_4841,N_4953);
nand U5023 (N_5023,N_4791,N_4934);
xnor U5024 (N_5024,N_4785,N_4909);
xnor U5025 (N_5025,N_4875,N_4908);
nand U5026 (N_5026,N_4774,N_4919);
or U5027 (N_5027,N_4769,N_4893);
and U5028 (N_5028,N_4789,N_4755);
or U5029 (N_5029,N_4807,N_4870);
or U5030 (N_5030,N_4787,N_4958);
and U5031 (N_5031,N_4851,N_4911);
nor U5032 (N_5032,N_4765,N_4752);
nor U5033 (N_5033,N_4808,N_4894);
nand U5034 (N_5034,N_4784,N_4920);
nor U5035 (N_5035,N_4990,N_4929);
or U5036 (N_5036,N_4813,N_4943);
nand U5037 (N_5037,N_4849,N_4823);
xor U5038 (N_5038,N_4927,N_4951);
xnor U5039 (N_5039,N_4954,N_4904);
nand U5040 (N_5040,N_4989,N_4915);
nor U5041 (N_5041,N_4859,N_4773);
or U5042 (N_5042,N_4946,N_4975);
nor U5043 (N_5043,N_4970,N_4979);
nor U5044 (N_5044,N_4864,N_4799);
xor U5045 (N_5045,N_4937,N_4838);
or U5046 (N_5046,N_4805,N_4949);
nor U5047 (N_5047,N_4968,N_4998);
nand U5048 (N_5048,N_4926,N_4783);
or U5049 (N_5049,N_4984,N_4819);
nand U5050 (N_5050,N_4829,N_4997);
or U5051 (N_5051,N_4940,N_4854);
nand U5052 (N_5052,N_4883,N_4768);
or U5053 (N_5053,N_4928,N_4810);
nor U5054 (N_5054,N_4772,N_4971);
xnor U5055 (N_5055,N_4775,N_4884);
and U5056 (N_5056,N_4891,N_4840);
and U5057 (N_5057,N_4857,N_4917);
nor U5058 (N_5058,N_4801,N_4936);
or U5059 (N_5059,N_4914,N_4962);
xnor U5060 (N_5060,N_4881,N_4939);
nor U5061 (N_5061,N_4860,N_4868);
xor U5062 (N_5062,N_4996,N_4757);
nor U5063 (N_5063,N_4931,N_4877);
nand U5064 (N_5064,N_4826,N_4932);
nor U5065 (N_5065,N_4797,N_4812);
or U5066 (N_5066,N_4957,N_4892);
xnor U5067 (N_5067,N_4982,N_4873);
xnor U5068 (N_5068,N_4882,N_4897);
xor U5069 (N_5069,N_4974,N_4872);
or U5070 (N_5070,N_4835,N_4798);
xor U5071 (N_5071,N_4961,N_4777);
xnor U5072 (N_5072,N_4889,N_4942);
nand U5073 (N_5073,N_4771,N_4809);
nand U5074 (N_5074,N_4916,N_4913);
xor U5075 (N_5075,N_4782,N_4985);
or U5076 (N_5076,N_4779,N_4888);
and U5077 (N_5077,N_4906,N_4861);
or U5078 (N_5078,N_4862,N_4879);
and U5079 (N_5079,N_4790,N_4763);
nand U5080 (N_5080,N_4761,N_4903);
xor U5081 (N_5081,N_4788,N_4885);
or U5082 (N_5082,N_4912,N_4886);
nand U5083 (N_5083,N_4950,N_4844);
nor U5084 (N_5084,N_4978,N_4955);
or U5085 (N_5085,N_4918,N_4762);
nand U5086 (N_5086,N_4825,N_4933);
nor U5087 (N_5087,N_4811,N_4874);
and U5088 (N_5088,N_4750,N_4945);
xnor U5089 (N_5089,N_4754,N_4969);
nor U5090 (N_5090,N_4999,N_4952);
or U5091 (N_5091,N_4900,N_4793);
nor U5092 (N_5092,N_4922,N_4832);
nor U5093 (N_5093,N_4842,N_4981);
nand U5094 (N_5094,N_4907,N_4923);
xor U5095 (N_5095,N_4964,N_4880);
nand U5096 (N_5096,N_4824,N_4831);
nand U5097 (N_5097,N_4846,N_4786);
and U5098 (N_5098,N_4827,N_4792);
nand U5099 (N_5099,N_4986,N_4766);
nor U5100 (N_5100,N_4993,N_4865);
nand U5101 (N_5101,N_4869,N_4756);
nor U5102 (N_5102,N_4778,N_4858);
and U5103 (N_5103,N_4947,N_4803);
nor U5104 (N_5104,N_4837,N_4804);
or U5105 (N_5105,N_4994,N_4965);
and U5106 (N_5106,N_4806,N_4821);
xor U5107 (N_5107,N_4770,N_4758);
or U5108 (N_5108,N_4843,N_4973);
or U5109 (N_5109,N_4815,N_4850);
or U5110 (N_5110,N_4890,N_4878);
and U5111 (N_5111,N_4948,N_4972);
and U5112 (N_5112,N_4802,N_4866);
nor U5113 (N_5113,N_4794,N_4988);
xor U5114 (N_5114,N_4760,N_4980);
xnor U5115 (N_5115,N_4938,N_4930);
and U5116 (N_5116,N_4830,N_4863);
xnor U5117 (N_5117,N_4800,N_4896);
and U5118 (N_5118,N_4960,N_4902);
xor U5119 (N_5119,N_4963,N_4853);
nor U5120 (N_5120,N_4759,N_4899);
nor U5121 (N_5121,N_4817,N_4895);
xor U5122 (N_5122,N_4956,N_4867);
nor U5123 (N_5123,N_4925,N_4781);
nor U5124 (N_5124,N_4983,N_4795);
and U5125 (N_5125,N_4924,N_4772);
or U5126 (N_5126,N_4980,N_4921);
nand U5127 (N_5127,N_4788,N_4839);
xor U5128 (N_5128,N_4970,N_4921);
xor U5129 (N_5129,N_4982,N_4979);
or U5130 (N_5130,N_4943,N_4897);
and U5131 (N_5131,N_4987,N_4813);
xor U5132 (N_5132,N_4874,N_4773);
nand U5133 (N_5133,N_4960,N_4994);
and U5134 (N_5134,N_4983,N_4875);
and U5135 (N_5135,N_4832,N_4995);
or U5136 (N_5136,N_4932,N_4971);
xor U5137 (N_5137,N_4756,N_4798);
nand U5138 (N_5138,N_4809,N_4756);
xor U5139 (N_5139,N_4887,N_4820);
nand U5140 (N_5140,N_4900,N_4838);
and U5141 (N_5141,N_4989,N_4793);
or U5142 (N_5142,N_4806,N_4954);
and U5143 (N_5143,N_4911,N_4949);
xnor U5144 (N_5144,N_4868,N_4889);
and U5145 (N_5145,N_4985,N_4937);
xor U5146 (N_5146,N_4821,N_4953);
xnor U5147 (N_5147,N_4942,N_4953);
nand U5148 (N_5148,N_4774,N_4816);
or U5149 (N_5149,N_4937,N_4833);
nand U5150 (N_5150,N_4861,N_4752);
and U5151 (N_5151,N_4793,N_4878);
and U5152 (N_5152,N_4846,N_4764);
nand U5153 (N_5153,N_4928,N_4920);
nor U5154 (N_5154,N_4828,N_4781);
or U5155 (N_5155,N_4763,N_4829);
and U5156 (N_5156,N_4934,N_4978);
or U5157 (N_5157,N_4868,N_4855);
or U5158 (N_5158,N_4887,N_4964);
and U5159 (N_5159,N_4917,N_4864);
nor U5160 (N_5160,N_4916,N_4857);
or U5161 (N_5161,N_4935,N_4826);
nand U5162 (N_5162,N_4933,N_4993);
nand U5163 (N_5163,N_4924,N_4771);
and U5164 (N_5164,N_4805,N_4758);
nor U5165 (N_5165,N_4899,N_4828);
nand U5166 (N_5166,N_4880,N_4990);
and U5167 (N_5167,N_4974,N_4811);
or U5168 (N_5168,N_4796,N_4935);
xnor U5169 (N_5169,N_4788,N_4967);
or U5170 (N_5170,N_4940,N_4879);
and U5171 (N_5171,N_4807,N_4971);
and U5172 (N_5172,N_4886,N_4960);
nand U5173 (N_5173,N_4936,N_4823);
or U5174 (N_5174,N_4859,N_4929);
xor U5175 (N_5175,N_4959,N_4938);
or U5176 (N_5176,N_4962,N_4765);
xnor U5177 (N_5177,N_4793,N_4824);
and U5178 (N_5178,N_4970,N_4969);
or U5179 (N_5179,N_4817,N_4826);
xnor U5180 (N_5180,N_4959,N_4849);
and U5181 (N_5181,N_4772,N_4896);
and U5182 (N_5182,N_4883,N_4843);
xnor U5183 (N_5183,N_4903,N_4888);
or U5184 (N_5184,N_4957,N_4913);
xnor U5185 (N_5185,N_4855,N_4990);
or U5186 (N_5186,N_4889,N_4911);
or U5187 (N_5187,N_4875,N_4984);
xnor U5188 (N_5188,N_4813,N_4807);
and U5189 (N_5189,N_4983,N_4920);
and U5190 (N_5190,N_4827,N_4777);
or U5191 (N_5191,N_4754,N_4893);
nand U5192 (N_5192,N_4839,N_4897);
nand U5193 (N_5193,N_4885,N_4810);
xnor U5194 (N_5194,N_4916,N_4824);
and U5195 (N_5195,N_4987,N_4850);
or U5196 (N_5196,N_4921,N_4974);
and U5197 (N_5197,N_4809,N_4792);
nor U5198 (N_5198,N_4767,N_4968);
xnor U5199 (N_5199,N_4818,N_4837);
and U5200 (N_5200,N_4875,N_4798);
xnor U5201 (N_5201,N_4999,N_4981);
nand U5202 (N_5202,N_4999,N_4820);
xor U5203 (N_5203,N_4936,N_4867);
xnor U5204 (N_5204,N_4778,N_4771);
nand U5205 (N_5205,N_4834,N_4873);
and U5206 (N_5206,N_4881,N_4805);
xnor U5207 (N_5207,N_4930,N_4995);
nand U5208 (N_5208,N_4796,N_4820);
or U5209 (N_5209,N_4754,N_4967);
nand U5210 (N_5210,N_4769,N_4870);
and U5211 (N_5211,N_4993,N_4885);
xor U5212 (N_5212,N_4905,N_4898);
xor U5213 (N_5213,N_4944,N_4822);
or U5214 (N_5214,N_4999,N_4768);
nor U5215 (N_5215,N_4771,N_4893);
and U5216 (N_5216,N_4997,N_4782);
xnor U5217 (N_5217,N_4770,N_4973);
nand U5218 (N_5218,N_4871,N_4845);
or U5219 (N_5219,N_4934,N_4886);
nand U5220 (N_5220,N_4842,N_4882);
or U5221 (N_5221,N_4799,N_4946);
nand U5222 (N_5222,N_4944,N_4885);
xnor U5223 (N_5223,N_4814,N_4993);
nand U5224 (N_5224,N_4971,N_4917);
xnor U5225 (N_5225,N_4914,N_4828);
xnor U5226 (N_5226,N_4811,N_4916);
and U5227 (N_5227,N_4757,N_4760);
nand U5228 (N_5228,N_4866,N_4959);
nand U5229 (N_5229,N_4817,N_4861);
xnor U5230 (N_5230,N_4899,N_4988);
xnor U5231 (N_5231,N_4974,N_4864);
xnor U5232 (N_5232,N_4900,N_4962);
and U5233 (N_5233,N_4893,N_4960);
nand U5234 (N_5234,N_4993,N_4970);
xor U5235 (N_5235,N_4996,N_4943);
nor U5236 (N_5236,N_4924,N_4831);
nor U5237 (N_5237,N_4970,N_4750);
nand U5238 (N_5238,N_4913,N_4879);
and U5239 (N_5239,N_4914,N_4889);
and U5240 (N_5240,N_4763,N_4923);
and U5241 (N_5241,N_4921,N_4998);
nor U5242 (N_5242,N_4831,N_4798);
nor U5243 (N_5243,N_4942,N_4919);
and U5244 (N_5244,N_4882,N_4778);
or U5245 (N_5245,N_4874,N_4865);
and U5246 (N_5246,N_4842,N_4973);
xor U5247 (N_5247,N_4909,N_4976);
or U5248 (N_5248,N_4878,N_4860);
nor U5249 (N_5249,N_4750,N_4872);
nor U5250 (N_5250,N_5171,N_5243);
nand U5251 (N_5251,N_5066,N_5044);
nand U5252 (N_5252,N_5120,N_5089);
nor U5253 (N_5253,N_5148,N_5144);
xor U5254 (N_5254,N_5127,N_5074);
nand U5255 (N_5255,N_5049,N_5134);
nand U5256 (N_5256,N_5205,N_5226);
xnor U5257 (N_5257,N_5113,N_5121);
nand U5258 (N_5258,N_5235,N_5024);
or U5259 (N_5259,N_5093,N_5136);
or U5260 (N_5260,N_5197,N_5220);
or U5261 (N_5261,N_5234,N_5155);
nand U5262 (N_5262,N_5130,N_5137);
nand U5263 (N_5263,N_5064,N_5102);
or U5264 (N_5264,N_5142,N_5214);
or U5265 (N_5265,N_5018,N_5054);
nand U5266 (N_5266,N_5019,N_5182);
and U5267 (N_5267,N_5020,N_5218);
xor U5268 (N_5268,N_5005,N_5163);
nand U5269 (N_5269,N_5114,N_5047);
xnor U5270 (N_5270,N_5085,N_5170);
nor U5271 (N_5271,N_5068,N_5147);
or U5272 (N_5272,N_5132,N_5126);
and U5273 (N_5273,N_5225,N_5196);
and U5274 (N_5274,N_5037,N_5149);
nor U5275 (N_5275,N_5061,N_5108);
and U5276 (N_5276,N_5216,N_5029);
nor U5277 (N_5277,N_5026,N_5161);
xor U5278 (N_5278,N_5115,N_5014);
and U5279 (N_5279,N_5128,N_5200);
nor U5280 (N_5280,N_5236,N_5143);
nand U5281 (N_5281,N_5230,N_5201);
nand U5282 (N_5282,N_5215,N_5055);
or U5283 (N_5283,N_5237,N_5183);
and U5284 (N_5284,N_5246,N_5125);
and U5285 (N_5285,N_5194,N_5103);
xnor U5286 (N_5286,N_5112,N_5206);
and U5287 (N_5287,N_5199,N_5123);
and U5288 (N_5288,N_5139,N_5135);
nor U5289 (N_5289,N_5110,N_5077);
or U5290 (N_5290,N_5092,N_5013);
nand U5291 (N_5291,N_5084,N_5032);
xor U5292 (N_5292,N_5070,N_5208);
and U5293 (N_5293,N_5079,N_5030);
xnor U5294 (N_5294,N_5238,N_5184);
nand U5295 (N_5295,N_5229,N_5154);
or U5296 (N_5296,N_5033,N_5035);
nand U5297 (N_5297,N_5189,N_5025);
and U5298 (N_5298,N_5232,N_5164);
nor U5299 (N_5299,N_5247,N_5156);
nand U5300 (N_5300,N_5105,N_5198);
xor U5301 (N_5301,N_5192,N_5187);
xor U5302 (N_5302,N_5086,N_5094);
nand U5303 (N_5303,N_5076,N_5056);
and U5304 (N_5304,N_5111,N_5219);
or U5305 (N_5305,N_5221,N_5099);
and U5306 (N_5306,N_5138,N_5028);
nand U5307 (N_5307,N_5248,N_5117);
nand U5308 (N_5308,N_5087,N_5202);
nand U5309 (N_5309,N_5078,N_5146);
and U5310 (N_5310,N_5165,N_5193);
and U5311 (N_5311,N_5222,N_5186);
xnor U5312 (N_5312,N_5012,N_5001);
or U5313 (N_5313,N_5158,N_5195);
and U5314 (N_5314,N_5104,N_5041);
xor U5315 (N_5315,N_5015,N_5071);
and U5316 (N_5316,N_5129,N_5209);
nand U5317 (N_5317,N_5212,N_5053);
xnor U5318 (N_5318,N_5242,N_5168);
and U5319 (N_5319,N_5177,N_5075);
and U5320 (N_5320,N_5207,N_5191);
nand U5321 (N_5321,N_5059,N_5040);
nor U5322 (N_5322,N_5160,N_5042);
or U5323 (N_5323,N_5095,N_5181);
or U5324 (N_5324,N_5213,N_5003);
xnor U5325 (N_5325,N_5211,N_5073);
nor U5326 (N_5326,N_5052,N_5091);
nor U5327 (N_5327,N_5060,N_5048);
or U5328 (N_5328,N_5167,N_5006);
and U5329 (N_5329,N_5017,N_5245);
nand U5330 (N_5330,N_5016,N_5227);
or U5331 (N_5331,N_5036,N_5097);
xor U5332 (N_5332,N_5151,N_5228);
or U5333 (N_5333,N_5180,N_5249);
xnor U5334 (N_5334,N_5010,N_5133);
nor U5335 (N_5335,N_5162,N_5116);
or U5336 (N_5336,N_5080,N_5058);
and U5337 (N_5337,N_5172,N_5027);
nand U5338 (N_5338,N_5153,N_5224);
or U5339 (N_5339,N_5081,N_5023);
or U5340 (N_5340,N_5090,N_5004);
xnor U5341 (N_5341,N_5223,N_5009);
nand U5342 (N_5342,N_5150,N_5000);
nor U5343 (N_5343,N_5022,N_5100);
nor U5344 (N_5344,N_5141,N_5157);
nand U5345 (N_5345,N_5179,N_5007);
or U5346 (N_5346,N_5185,N_5188);
nand U5347 (N_5347,N_5175,N_5031);
nand U5348 (N_5348,N_5106,N_5008);
nand U5349 (N_5349,N_5169,N_5145);
nand U5350 (N_5350,N_5231,N_5045);
or U5351 (N_5351,N_5065,N_5176);
and U5352 (N_5352,N_5166,N_5109);
and U5353 (N_5353,N_5203,N_5210);
or U5354 (N_5354,N_5107,N_5131);
and U5355 (N_5355,N_5159,N_5002);
nand U5356 (N_5356,N_5096,N_5051);
xnor U5357 (N_5357,N_5057,N_5152);
nand U5358 (N_5358,N_5240,N_5082);
and U5359 (N_5359,N_5043,N_5069);
and U5360 (N_5360,N_5118,N_5072);
nor U5361 (N_5361,N_5122,N_5204);
nand U5362 (N_5362,N_5039,N_5173);
nand U5363 (N_5363,N_5217,N_5174);
or U5364 (N_5364,N_5067,N_5011);
xor U5365 (N_5365,N_5124,N_5178);
xor U5366 (N_5366,N_5050,N_5119);
or U5367 (N_5367,N_5190,N_5046);
or U5368 (N_5368,N_5101,N_5140);
nor U5369 (N_5369,N_5098,N_5021);
or U5370 (N_5370,N_5244,N_5038);
xnor U5371 (N_5371,N_5083,N_5088);
xnor U5372 (N_5372,N_5063,N_5233);
nand U5373 (N_5373,N_5239,N_5241);
xnor U5374 (N_5374,N_5034,N_5062);
or U5375 (N_5375,N_5243,N_5217);
or U5376 (N_5376,N_5097,N_5213);
nor U5377 (N_5377,N_5082,N_5090);
nand U5378 (N_5378,N_5023,N_5241);
xnor U5379 (N_5379,N_5015,N_5115);
and U5380 (N_5380,N_5080,N_5239);
xor U5381 (N_5381,N_5217,N_5147);
and U5382 (N_5382,N_5231,N_5062);
xnor U5383 (N_5383,N_5247,N_5172);
and U5384 (N_5384,N_5217,N_5171);
or U5385 (N_5385,N_5126,N_5017);
xor U5386 (N_5386,N_5040,N_5222);
xnor U5387 (N_5387,N_5169,N_5022);
nand U5388 (N_5388,N_5055,N_5021);
xnor U5389 (N_5389,N_5113,N_5042);
or U5390 (N_5390,N_5232,N_5124);
nand U5391 (N_5391,N_5142,N_5240);
and U5392 (N_5392,N_5132,N_5106);
and U5393 (N_5393,N_5099,N_5158);
and U5394 (N_5394,N_5104,N_5064);
or U5395 (N_5395,N_5171,N_5057);
nand U5396 (N_5396,N_5069,N_5194);
or U5397 (N_5397,N_5245,N_5136);
xnor U5398 (N_5398,N_5056,N_5070);
xor U5399 (N_5399,N_5135,N_5184);
nor U5400 (N_5400,N_5209,N_5135);
or U5401 (N_5401,N_5201,N_5140);
xnor U5402 (N_5402,N_5244,N_5149);
and U5403 (N_5403,N_5088,N_5080);
nand U5404 (N_5404,N_5184,N_5116);
and U5405 (N_5405,N_5210,N_5144);
nor U5406 (N_5406,N_5169,N_5063);
xnor U5407 (N_5407,N_5165,N_5129);
and U5408 (N_5408,N_5132,N_5226);
nor U5409 (N_5409,N_5109,N_5197);
nor U5410 (N_5410,N_5059,N_5161);
nor U5411 (N_5411,N_5197,N_5118);
nand U5412 (N_5412,N_5054,N_5176);
or U5413 (N_5413,N_5239,N_5170);
nor U5414 (N_5414,N_5236,N_5156);
or U5415 (N_5415,N_5151,N_5044);
or U5416 (N_5416,N_5190,N_5223);
or U5417 (N_5417,N_5227,N_5055);
nor U5418 (N_5418,N_5104,N_5151);
nand U5419 (N_5419,N_5020,N_5049);
or U5420 (N_5420,N_5245,N_5226);
nand U5421 (N_5421,N_5179,N_5201);
or U5422 (N_5422,N_5123,N_5168);
and U5423 (N_5423,N_5072,N_5043);
or U5424 (N_5424,N_5053,N_5113);
or U5425 (N_5425,N_5149,N_5158);
and U5426 (N_5426,N_5030,N_5087);
nor U5427 (N_5427,N_5155,N_5044);
and U5428 (N_5428,N_5148,N_5104);
and U5429 (N_5429,N_5078,N_5242);
nor U5430 (N_5430,N_5226,N_5109);
xor U5431 (N_5431,N_5055,N_5009);
and U5432 (N_5432,N_5113,N_5213);
xnor U5433 (N_5433,N_5199,N_5127);
or U5434 (N_5434,N_5169,N_5163);
xor U5435 (N_5435,N_5183,N_5062);
xnor U5436 (N_5436,N_5193,N_5029);
nand U5437 (N_5437,N_5166,N_5080);
and U5438 (N_5438,N_5169,N_5241);
or U5439 (N_5439,N_5229,N_5128);
xnor U5440 (N_5440,N_5190,N_5246);
or U5441 (N_5441,N_5017,N_5059);
or U5442 (N_5442,N_5035,N_5204);
xnor U5443 (N_5443,N_5094,N_5158);
nand U5444 (N_5444,N_5001,N_5056);
xnor U5445 (N_5445,N_5200,N_5044);
nor U5446 (N_5446,N_5092,N_5051);
or U5447 (N_5447,N_5244,N_5063);
xnor U5448 (N_5448,N_5181,N_5203);
or U5449 (N_5449,N_5236,N_5072);
nand U5450 (N_5450,N_5003,N_5059);
and U5451 (N_5451,N_5189,N_5106);
and U5452 (N_5452,N_5215,N_5026);
or U5453 (N_5453,N_5155,N_5185);
nand U5454 (N_5454,N_5200,N_5085);
xnor U5455 (N_5455,N_5238,N_5075);
xor U5456 (N_5456,N_5027,N_5119);
nor U5457 (N_5457,N_5203,N_5015);
nor U5458 (N_5458,N_5184,N_5165);
or U5459 (N_5459,N_5040,N_5071);
nand U5460 (N_5460,N_5206,N_5080);
xnor U5461 (N_5461,N_5089,N_5036);
and U5462 (N_5462,N_5169,N_5019);
or U5463 (N_5463,N_5213,N_5107);
or U5464 (N_5464,N_5148,N_5014);
xor U5465 (N_5465,N_5182,N_5209);
nand U5466 (N_5466,N_5212,N_5086);
nor U5467 (N_5467,N_5232,N_5213);
nor U5468 (N_5468,N_5196,N_5071);
and U5469 (N_5469,N_5233,N_5242);
nor U5470 (N_5470,N_5017,N_5129);
xnor U5471 (N_5471,N_5164,N_5179);
nand U5472 (N_5472,N_5209,N_5073);
nor U5473 (N_5473,N_5114,N_5131);
and U5474 (N_5474,N_5219,N_5168);
and U5475 (N_5475,N_5148,N_5133);
nor U5476 (N_5476,N_5093,N_5114);
and U5477 (N_5477,N_5095,N_5003);
xor U5478 (N_5478,N_5108,N_5204);
xnor U5479 (N_5479,N_5049,N_5100);
nor U5480 (N_5480,N_5065,N_5089);
nand U5481 (N_5481,N_5126,N_5226);
xor U5482 (N_5482,N_5043,N_5110);
xnor U5483 (N_5483,N_5093,N_5165);
xor U5484 (N_5484,N_5031,N_5165);
nor U5485 (N_5485,N_5179,N_5207);
nor U5486 (N_5486,N_5159,N_5150);
xor U5487 (N_5487,N_5063,N_5061);
xnor U5488 (N_5488,N_5129,N_5091);
nor U5489 (N_5489,N_5100,N_5059);
or U5490 (N_5490,N_5181,N_5073);
or U5491 (N_5491,N_5067,N_5059);
xor U5492 (N_5492,N_5097,N_5237);
nor U5493 (N_5493,N_5146,N_5087);
and U5494 (N_5494,N_5160,N_5041);
and U5495 (N_5495,N_5012,N_5190);
and U5496 (N_5496,N_5174,N_5133);
xor U5497 (N_5497,N_5164,N_5069);
and U5498 (N_5498,N_5075,N_5241);
nand U5499 (N_5499,N_5214,N_5057);
xnor U5500 (N_5500,N_5260,N_5335);
xnor U5501 (N_5501,N_5256,N_5327);
nand U5502 (N_5502,N_5287,N_5396);
or U5503 (N_5503,N_5254,N_5434);
and U5504 (N_5504,N_5405,N_5401);
xnor U5505 (N_5505,N_5473,N_5252);
or U5506 (N_5506,N_5407,N_5420);
xnor U5507 (N_5507,N_5492,N_5317);
or U5508 (N_5508,N_5482,N_5476);
nor U5509 (N_5509,N_5378,N_5293);
nand U5510 (N_5510,N_5422,N_5448);
nand U5511 (N_5511,N_5319,N_5341);
nor U5512 (N_5512,N_5379,N_5373);
nor U5513 (N_5513,N_5475,N_5450);
xor U5514 (N_5514,N_5261,N_5390);
and U5515 (N_5515,N_5384,N_5343);
or U5516 (N_5516,N_5302,N_5483);
nor U5517 (N_5517,N_5380,N_5470);
nor U5518 (N_5518,N_5352,N_5445);
and U5519 (N_5519,N_5326,N_5342);
xor U5520 (N_5520,N_5251,N_5312);
xnor U5521 (N_5521,N_5354,N_5348);
nand U5522 (N_5522,N_5403,N_5416);
nand U5523 (N_5523,N_5376,N_5338);
and U5524 (N_5524,N_5438,N_5320);
nor U5525 (N_5525,N_5439,N_5307);
xor U5526 (N_5526,N_5368,N_5477);
nor U5527 (N_5527,N_5421,N_5441);
and U5528 (N_5528,N_5406,N_5290);
and U5529 (N_5529,N_5485,N_5336);
or U5530 (N_5530,N_5364,N_5316);
xnor U5531 (N_5531,N_5334,N_5299);
nand U5532 (N_5532,N_5346,N_5276);
nand U5533 (N_5533,N_5369,N_5488);
xnor U5534 (N_5534,N_5387,N_5271);
or U5535 (N_5535,N_5371,N_5493);
xor U5536 (N_5536,N_5321,N_5350);
nor U5537 (N_5537,N_5402,N_5363);
xor U5538 (N_5538,N_5463,N_5392);
and U5539 (N_5539,N_5372,N_5412);
or U5540 (N_5540,N_5433,N_5386);
nor U5541 (N_5541,N_5385,N_5487);
nor U5542 (N_5542,N_5353,N_5471);
and U5543 (N_5543,N_5451,N_5272);
nor U5544 (N_5544,N_5367,N_5255);
xnor U5545 (N_5545,N_5355,N_5417);
nand U5546 (N_5546,N_5397,N_5395);
nand U5547 (N_5547,N_5262,N_5486);
nor U5548 (N_5548,N_5258,N_5329);
xor U5549 (N_5549,N_5310,N_5359);
nand U5550 (N_5550,N_5452,N_5468);
nor U5551 (N_5551,N_5459,N_5311);
or U5552 (N_5552,N_5298,N_5496);
or U5553 (N_5553,N_5361,N_5305);
and U5554 (N_5554,N_5300,N_5456);
or U5555 (N_5555,N_5408,N_5288);
xor U5556 (N_5556,N_5279,N_5399);
nor U5557 (N_5557,N_5495,N_5388);
xor U5558 (N_5558,N_5425,N_5351);
nand U5559 (N_5559,N_5398,N_5362);
nand U5560 (N_5560,N_5337,N_5484);
or U5561 (N_5561,N_5436,N_5285);
xor U5562 (N_5562,N_5332,N_5466);
or U5563 (N_5563,N_5275,N_5499);
nand U5564 (N_5564,N_5446,N_5318);
nor U5565 (N_5565,N_5479,N_5462);
nor U5566 (N_5566,N_5419,N_5283);
nor U5567 (N_5567,N_5382,N_5366);
xor U5568 (N_5568,N_5423,N_5404);
xor U5569 (N_5569,N_5280,N_5347);
xor U5570 (N_5570,N_5328,N_5340);
xnor U5571 (N_5571,N_5357,N_5391);
and U5572 (N_5572,N_5315,N_5264);
or U5573 (N_5573,N_5281,N_5297);
nor U5574 (N_5574,N_5410,N_5274);
nand U5575 (N_5575,N_5447,N_5374);
or U5576 (N_5576,N_5427,N_5432);
or U5577 (N_5577,N_5467,N_5306);
and U5578 (N_5578,N_5429,N_5322);
and U5579 (N_5579,N_5472,N_5313);
xnor U5580 (N_5580,N_5469,N_5286);
or U5581 (N_5581,N_5303,N_5444);
xnor U5582 (N_5582,N_5413,N_5291);
and U5583 (N_5583,N_5377,N_5418);
nor U5584 (N_5584,N_5284,N_5282);
nand U5585 (N_5585,N_5424,N_5344);
nor U5586 (N_5586,N_5497,N_5259);
and U5587 (N_5587,N_5269,N_5333);
nor U5588 (N_5588,N_5266,N_5325);
or U5589 (N_5589,N_5430,N_5461);
nor U5590 (N_5590,N_5381,N_5465);
nor U5591 (N_5591,N_5331,N_5440);
xor U5592 (N_5592,N_5292,N_5383);
nor U5593 (N_5593,N_5370,N_5265);
xnor U5594 (N_5594,N_5414,N_5435);
or U5595 (N_5595,N_5494,N_5449);
or U5596 (N_5596,N_5314,N_5394);
nand U5597 (N_5597,N_5454,N_5457);
nor U5598 (N_5598,N_5443,N_5323);
nor U5599 (N_5599,N_5428,N_5481);
xnor U5600 (N_5600,N_5455,N_5442);
nand U5601 (N_5601,N_5409,N_5278);
xor U5602 (N_5602,N_5273,N_5268);
xnor U5603 (N_5603,N_5358,N_5375);
nor U5604 (N_5604,N_5478,N_5289);
or U5605 (N_5605,N_5296,N_5309);
nand U5606 (N_5606,N_5257,N_5277);
nor U5607 (N_5607,N_5330,N_5349);
nand U5608 (N_5608,N_5360,N_5389);
nor U5609 (N_5609,N_5415,N_5324);
nor U5610 (N_5610,N_5267,N_5250);
and U5611 (N_5611,N_5460,N_5437);
or U5612 (N_5612,N_5480,N_5431);
and U5613 (N_5613,N_5253,N_5498);
nand U5614 (N_5614,N_5453,N_5489);
xor U5615 (N_5615,N_5411,N_5345);
and U5616 (N_5616,N_5491,N_5270);
nor U5617 (N_5617,N_5490,N_5426);
and U5618 (N_5618,N_5304,N_5393);
or U5619 (N_5619,N_5400,N_5464);
xnor U5620 (N_5620,N_5356,N_5458);
xor U5621 (N_5621,N_5301,N_5263);
nand U5622 (N_5622,N_5294,N_5308);
or U5623 (N_5623,N_5365,N_5339);
and U5624 (N_5624,N_5474,N_5295);
and U5625 (N_5625,N_5386,N_5374);
or U5626 (N_5626,N_5261,N_5363);
nand U5627 (N_5627,N_5368,N_5497);
nor U5628 (N_5628,N_5472,N_5425);
or U5629 (N_5629,N_5304,N_5418);
and U5630 (N_5630,N_5469,N_5316);
nor U5631 (N_5631,N_5284,N_5452);
and U5632 (N_5632,N_5398,N_5491);
nor U5633 (N_5633,N_5371,N_5424);
nand U5634 (N_5634,N_5342,N_5312);
or U5635 (N_5635,N_5412,N_5397);
or U5636 (N_5636,N_5362,N_5350);
nand U5637 (N_5637,N_5499,N_5262);
and U5638 (N_5638,N_5337,N_5250);
and U5639 (N_5639,N_5432,N_5419);
or U5640 (N_5640,N_5258,N_5454);
xnor U5641 (N_5641,N_5250,N_5377);
and U5642 (N_5642,N_5384,N_5317);
and U5643 (N_5643,N_5465,N_5467);
xor U5644 (N_5644,N_5485,N_5397);
or U5645 (N_5645,N_5307,N_5310);
xnor U5646 (N_5646,N_5432,N_5485);
nor U5647 (N_5647,N_5400,N_5296);
or U5648 (N_5648,N_5404,N_5342);
and U5649 (N_5649,N_5401,N_5383);
xor U5650 (N_5650,N_5363,N_5296);
nor U5651 (N_5651,N_5303,N_5255);
or U5652 (N_5652,N_5387,N_5470);
or U5653 (N_5653,N_5444,N_5364);
xor U5654 (N_5654,N_5407,N_5319);
nand U5655 (N_5655,N_5459,N_5388);
and U5656 (N_5656,N_5332,N_5451);
and U5657 (N_5657,N_5452,N_5478);
nand U5658 (N_5658,N_5263,N_5450);
and U5659 (N_5659,N_5282,N_5340);
or U5660 (N_5660,N_5457,N_5405);
nor U5661 (N_5661,N_5468,N_5456);
or U5662 (N_5662,N_5485,N_5434);
and U5663 (N_5663,N_5479,N_5380);
nand U5664 (N_5664,N_5316,N_5380);
nor U5665 (N_5665,N_5445,N_5448);
nor U5666 (N_5666,N_5265,N_5267);
nor U5667 (N_5667,N_5423,N_5409);
or U5668 (N_5668,N_5390,N_5307);
or U5669 (N_5669,N_5463,N_5466);
nand U5670 (N_5670,N_5257,N_5316);
and U5671 (N_5671,N_5400,N_5355);
xnor U5672 (N_5672,N_5470,N_5336);
xor U5673 (N_5673,N_5285,N_5350);
or U5674 (N_5674,N_5267,N_5355);
or U5675 (N_5675,N_5285,N_5302);
nand U5676 (N_5676,N_5455,N_5359);
or U5677 (N_5677,N_5272,N_5432);
xnor U5678 (N_5678,N_5431,N_5250);
xnor U5679 (N_5679,N_5481,N_5445);
nand U5680 (N_5680,N_5460,N_5267);
xor U5681 (N_5681,N_5412,N_5424);
and U5682 (N_5682,N_5270,N_5489);
nand U5683 (N_5683,N_5346,N_5345);
nand U5684 (N_5684,N_5421,N_5352);
nand U5685 (N_5685,N_5388,N_5462);
xnor U5686 (N_5686,N_5272,N_5422);
and U5687 (N_5687,N_5250,N_5327);
nor U5688 (N_5688,N_5472,N_5316);
nor U5689 (N_5689,N_5488,N_5366);
or U5690 (N_5690,N_5257,N_5290);
nor U5691 (N_5691,N_5339,N_5402);
or U5692 (N_5692,N_5360,N_5408);
or U5693 (N_5693,N_5337,N_5322);
or U5694 (N_5694,N_5425,N_5268);
xnor U5695 (N_5695,N_5275,N_5324);
xor U5696 (N_5696,N_5437,N_5454);
nor U5697 (N_5697,N_5365,N_5402);
nor U5698 (N_5698,N_5297,N_5476);
xnor U5699 (N_5699,N_5410,N_5381);
nand U5700 (N_5700,N_5406,N_5307);
or U5701 (N_5701,N_5278,N_5297);
or U5702 (N_5702,N_5258,N_5327);
xor U5703 (N_5703,N_5401,N_5445);
xor U5704 (N_5704,N_5367,N_5384);
nand U5705 (N_5705,N_5336,N_5331);
or U5706 (N_5706,N_5410,N_5349);
or U5707 (N_5707,N_5410,N_5255);
or U5708 (N_5708,N_5322,N_5473);
xor U5709 (N_5709,N_5284,N_5270);
or U5710 (N_5710,N_5408,N_5450);
and U5711 (N_5711,N_5478,N_5480);
xnor U5712 (N_5712,N_5322,N_5499);
or U5713 (N_5713,N_5449,N_5466);
or U5714 (N_5714,N_5337,N_5435);
nand U5715 (N_5715,N_5403,N_5363);
xor U5716 (N_5716,N_5385,N_5340);
and U5717 (N_5717,N_5457,N_5470);
nand U5718 (N_5718,N_5266,N_5488);
or U5719 (N_5719,N_5439,N_5461);
xor U5720 (N_5720,N_5311,N_5452);
nor U5721 (N_5721,N_5370,N_5400);
nand U5722 (N_5722,N_5437,N_5449);
and U5723 (N_5723,N_5338,N_5331);
nor U5724 (N_5724,N_5290,N_5306);
and U5725 (N_5725,N_5335,N_5483);
and U5726 (N_5726,N_5416,N_5462);
xnor U5727 (N_5727,N_5285,N_5420);
nor U5728 (N_5728,N_5436,N_5394);
nand U5729 (N_5729,N_5352,N_5277);
nor U5730 (N_5730,N_5322,N_5377);
xnor U5731 (N_5731,N_5252,N_5372);
and U5732 (N_5732,N_5258,N_5339);
or U5733 (N_5733,N_5333,N_5375);
and U5734 (N_5734,N_5328,N_5325);
nand U5735 (N_5735,N_5375,N_5340);
or U5736 (N_5736,N_5498,N_5304);
xor U5737 (N_5737,N_5253,N_5464);
nor U5738 (N_5738,N_5267,N_5341);
xnor U5739 (N_5739,N_5287,N_5354);
nand U5740 (N_5740,N_5417,N_5305);
nand U5741 (N_5741,N_5434,N_5293);
xor U5742 (N_5742,N_5332,N_5256);
or U5743 (N_5743,N_5310,N_5423);
and U5744 (N_5744,N_5494,N_5314);
nor U5745 (N_5745,N_5319,N_5367);
nand U5746 (N_5746,N_5433,N_5392);
nand U5747 (N_5747,N_5332,N_5432);
and U5748 (N_5748,N_5480,N_5300);
xnor U5749 (N_5749,N_5462,N_5465);
xor U5750 (N_5750,N_5655,N_5621);
and U5751 (N_5751,N_5589,N_5578);
or U5752 (N_5752,N_5748,N_5568);
nor U5753 (N_5753,N_5741,N_5582);
xnor U5754 (N_5754,N_5673,N_5500);
xor U5755 (N_5755,N_5606,N_5711);
nand U5756 (N_5756,N_5556,N_5574);
or U5757 (N_5757,N_5543,N_5648);
xnor U5758 (N_5758,N_5581,N_5680);
and U5759 (N_5759,N_5546,N_5623);
nand U5760 (N_5760,N_5514,N_5722);
or U5761 (N_5761,N_5615,N_5629);
nor U5762 (N_5762,N_5735,N_5674);
or U5763 (N_5763,N_5745,N_5704);
xnor U5764 (N_5764,N_5517,N_5594);
and U5765 (N_5765,N_5566,N_5573);
or U5766 (N_5766,N_5605,N_5620);
and U5767 (N_5767,N_5631,N_5628);
and U5768 (N_5768,N_5625,N_5636);
nand U5769 (N_5769,N_5721,N_5522);
and U5770 (N_5770,N_5511,N_5718);
or U5771 (N_5771,N_5603,N_5508);
nand U5772 (N_5772,N_5697,N_5627);
xor U5773 (N_5773,N_5563,N_5665);
or U5774 (N_5774,N_5521,N_5667);
nand U5775 (N_5775,N_5576,N_5687);
nor U5776 (N_5776,N_5746,N_5661);
nand U5777 (N_5777,N_5541,N_5707);
or U5778 (N_5778,N_5678,N_5698);
nand U5779 (N_5779,N_5717,N_5702);
and U5780 (N_5780,N_5658,N_5656);
and U5781 (N_5781,N_5677,N_5690);
xor U5782 (N_5782,N_5641,N_5539);
xnor U5783 (N_5783,N_5577,N_5531);
xor U5784 (N_5784,N_5557,N_5716);
xor U5785 (N_5785,N_5545,N_5599);
xnor U5786 (N_5786,N_5709,N_5713);
xnor U5787 (N_5787,N_5724,N_5561);
nand U5788 (N_5788,N_5725,N_5688);
or U5789 (N_5789,N_5512,N_5670);
or U5790 (N_5790,N_5731,N_5579);
nand U5791 (N_5791,N_5564,N_5518);
and U5792 (N_5792,N_5558,N_5684);
nand U5793 (N_5793,N_5715,N_5683);
nand U5794 (N_5794,N_5747,N_5657);
or U5795 (N_5795,N_5602,N_5618);
xnor U5796 (N_5796,N_5727,N_5696);
or U5797 (N_5797,N_5549,N_5572);
nor U5798 (N_5798,N_5634,N_5570);
nor U5799 (N_5799,N_5613,N_5614);
nand U5800 (N_5800,N_5525,N_5530);
and U5801 (N_5801,N_5528,N_5749);
nand U5802 (N_5802,N_5699,N_5672);
nand U5803 (N_5803,N_5509,N_5538);
nand U5804 (N_5804,N_5555,N_5583);
xor U5805 (N_5805,N_5700,N_5565);
or U5806 (N_5806,N_5624,N_5560);
and U5807 (N_5807,N_5596,N_5652);
or U5808 (N_5808,N_5710,N_5647);
nor U5809 (N_5809,N_5681,N_5626);
nor U5810 (N_5810,N_5616,N_5501);
nor U5811 (N_5811,N_5695,N_5679);
nor U5812 (N_5812,N_5744,N_5692);
or U5813 (N_5813,N_5600,N_5736);
or U5814 (N_5814,N_5633,N_5617);
xnor U5815 (N_5815,N_5686,N_5732);
xor U5816 (N_5816,N_5723,N_5671);
xor U5817 (N_5817,N_5593,N_5638);
nand U5818 (N_5818,N_5646,N_5554);
nor U5819 (N_5819,N_5575,N_5654);
and U5820 (N_5820,N_5571,N_5653);
nor U5821 (N_5821,N_5726,N_5585);
nand U5822 (N_5822,N_5693,N_5701);
nand U5823 (N_5823,N_5743,N_5642);
or U5824 (N_5824,N_5567,N_5740);
nand U5825 (N_5825,N_5608,N_5590);
xnor U5826 (N_5826,N_5551,N_5635);
nand U5827 (N_5827,N_5552,N_5529);
xor U5828 (N_5828,N_5535,N_5675);
and U5829 (N_5829,N_5651,N_5506);
or U5830 (N_5830,N_5685,N_5728);
xnor U5831 (N_5831,N_5664,N_5534);
or U5832 (N_5832,N_5662,N_5720);
xnor U5833 (N_5833,N_5729,N_5586);
xnor U5834 (N_5834,N_5588,N_5640);
nor U5835 (N_5835,N_5540,N_5519);
or U5836 (N_5836,N_5659,N_5604);
or U5837 (N_5837,N_5595,N_5553);
nand U5838 (N_5838,N_5520,N_5513);
or U5839 (N_5839,N_5502,N_5533);
and U5840 (N_5840,N_5632,N_5547);
and U5841 (N_5841,N_5691,N_5607);
nand U5842 (N_5842,N_5562,N_5510);
nand U5843 (N_5843,N_5649,N_5592);
nor U5844 (N_5844,N_5612,N_5703);
or U5845 (N_5845,N_5584,N_5619);
nor U5846 (N_5846,N_5597,N_5705);
and U5847 (N_5847,N_5550,N_5503);
nor U5848 (N_5848,N_5598,N_5610);
xnor U5849 (N_5849,N_5676,N_5548);
nor U5850 (N_5850,N_5708,N_5668);
and U5851 (N_5851,N_5719,N_5515);
nand U5852 (N_5852,N_5587,N_5730);
xor U5853 (N_5853,N_5569,N_5714);
nand U5854 (N_5854,N_5516,N_5622);
or U5855 (N_5855,N_5601,N_5666);
or U5856 (N_5856,N_5643,N_5630);
or U5857 (N_5857,N_5526,N_5544);
nor U5858 (N_5858,N_5712,N_5532);
nor U5859 (N_5859,N_5507,N_5536);
or U5860 (N_5860,N_5689,N_5738);
xor U5861 (N_5861,N_5537,N_5639);
xnor U5862 (N_5862,N_5737,N_5644);
xnor U5863 (N_5863,N_5650,N_5734);
and U5864 (N_5864,N_5523,N_5733);
nor U5865 (N_5865,N_5669,N_5542);
nor U5866 (N_5866,N_5706,N_5742);
nor U5867 (N_5867,N_5694,N_5611);
nand U5868 (N_5868,N_5609,N_5663);
nor U5869 (N_5869,N_5645,N_5591);
and U5870 (N_5870,N_5504,N_5527);
xnor U5871 (N_5871,N_5524,N_5637);
and U5872 (N_5872,N_5682,N_5505);
xnor U5873 (N_5873,N_5559,N_5660);
or U5874 (N_5874,N_5739,N_5580);
xor U5875 (N_5875,N_5683,N_5717);
nor U5876 (N_5876,N_5555,N_5524);
nand U5877 (N_5877,N_5651,N_5676);
nand U5878 (N_5878,N_5512,N_5697);
nor U5879 (N_5879,N_5605,N_5561);
or U5880 (N_5880,N_5746,N_5623);
nor U5881 (N_5881,N_5589,N_5649);
nand U5882 (N_5882,N_5654,N_5706);
nor U5883 (N_5883,N_5715,N_5590);
and U5884 (N_5884,N_5543,N_5643);
nor U5885 (N_5885,N_5732,N_5552);
and U5886 (N_5886,N_5559,N_5709);
xnor U5887 (N_5887,N_5678,N_5637);
nor U5888 (N_5888,N_5694,N_5607);
nor U5889 (N_5889,N_5719,N_5616);
or U5890 (N_5890,N_5672,N_5665);
or U5891 (N_5891,N_5567,N_5619);
xnor U5892 (N_5892,N_5529,N_5662);
xor U5893 (N_5893,N_5608,N_5531);
or U5894 (N_5894,N_5569,N_5605);
or U5895 (N_5895,N_5701,N_5615);
xnor U5896 (N_5896,N_5722,N_5683);
or U5897 (N_5897,N_5638,N_5642);
or U5898 (N_5898,N_5506,N_5633);
nor U5899 (N_5899,N_5661,N_5693);
nor U5900 (N_5900,N_5559,N_5519);
and U5901 (N_5901,N_5642,N_5683);
nor U5902 (N_5902,N_5643,N_5540);
nor U5903 (N_5903,N_5734,N_5597);
nand U5904 (N_5904,N_5537,N_5748);
nand U5905 (N_5905,N_5565,N_5665);
nor U5906 (N_5906,N_5636,N_5532);
xnor U5907 (N_5907,N_5519,N_5695);
or U5908 (N_5908,N_5554,N_5727);
or U5909 (N_5909,N_5635,N_5614);
xnor U5910 (N_5910,N_5716,N_5559);
nor U5911 (N_5911,N_5612,N_5742);
nand U5912 (N_5912,N_5600,N_5543);
and U5913 (N_5913,N_5578,N_5568);
nor U5914 (N_5914,N_5509,N_5717);
and U5915 (N_5915,N_5539,N_5725);
nor U5916 (N_5916,N_5712,N_5652);
and U5917 (N_5917,N_5618,N_5643);
or U5918 (N_5918,N_5501,N_5673);
and U5919 (N_5919,N_5526,N_5718);
nor U5920 (N_5920,N_5528,N_5520);
or U5921 (N_5921,N_5531,N_5586);
nor U5922 (N_5922,N_5678,N_5581);
and U5923 (N_5923,N_5594,N_5747);
nor U5924 (N_5924,N_5516,N_5604);
nor U5925 (N_5925,N_5565,N_5704);
xnor U5926 (N_5926,N_5628,N_5651);
and U5927 (N_5927,N_5721,N_5729);
or U5928 (N_5928,N_5583,N_5616);
or U5929 (N_5929,N_5737,N_5507);
nand U5930 (N_5930,N_5737,N_5587);
nand U5931 (N_5931,N_5684,N_5567);
nor U5932 (N_5932,N_5735,N_5653);
xnor U5933 (N_5933,N_5548,N_5668);
nor U5934 (N_5934,N_5565,N_5671);
nand U5935 (N_5935,N_5502,N_5557);
nand U5936 (N_5936,N_5530,N_5702);
nand U5937 (N_5937,N_5550,N_5736);
xnor U5938 (N_5938,N_5508,N_5665);
or U5939 (N_5939,N_5552,N_5588);
and U5940 (N_5940,N_5699,N_5538);
nor U5941 (N_5941,N_5525,N_5554);
nand U5942 (N_5942,N_5749,N_5683);
nor U5943 (N_5943,N_5541,N_5651);
nand U5944 (N_5944,N_5552,N_5555);
or U5945 (N_5945,N_5612,N_5652);
and U5946 (N_5946,N_5627,N_5701);
and U5947 (N_5947,N_5669,N_5616);
xor U5948 (N_5948,N_5647,N_5620);
and U5949 (N_5949,N_5619,N_5576);
xnor U5950 (N_5950,N_5668,N_5569);
or U5951 (N_5951,N_5647,N_5560);
and U5952 (N_5952,N_5696,N_5693);
nand U5953 (N_5953,N_5515,N_5520);
and U5954 (N_5954,N_5502,N_5705);
or U5955 (N_5955,N_5652,N_5644);
nor U5956 (N_5956,N_5638,N_5536);
nor U5957 (N_5957,N_5665,N_5603);
and U5958 (N_5958,N_5501,N_5517);
nand U5959 (N_5959,N_5555,N_5638);
xor U5960 (N_5960,N_5630,N_5504);
nand U5961 (N_5961,N_5593,N_5581);
or U5962 (N_5962,N_5616,N_5545);
nor U5963 (N_5963,N_5577,N_5623);
nand U5964 (N_5964,N_5675,N_5586);
and U5965 (N_5965,N_5641,N_5600);
xor U5966 (N_5966,N_5704,N_5520);
nor U5967 (N_5967,N_5737,N_5512);
nand U5968 (N_5968,N_5683,N_5548);
or U5969 (N_5969,N_5702,N_5561);
nand U5970 (N_5970,N_5743,N_5530);
or U5971 (N_5971,N_5560,N_5604);
nor U5972 (N_5972,N_5646,N_5687);
and U5973 (N_5973,N_5501,N_5694);
or U5974 (N_5974,N_5721,N_5581);
nand U5975 (N_5975,N_5660,N_5615);
nor U5976 (N_5976,N_5734,N_5503);
or U5977 (N_5977,N_5672,N_5703);
and U5978 (N_5978,N_5649,N_5736);
nor U5979 (N_5979,N_5530,N_5656);
xor U5980 (N_5980,N_5594,N_5616);
or U5981 (N_5981,N_5715,N_5687);
xor U5982 (N_5982,N_5638,N_5572);
and U5983 (N_5983,N_5642,N_5700);
nand U5984 (N_5984,N_5741,N_5600);
or U5985 (N_5985,N_5579,N_5708);
xnor U5986 (N_5986,N_5724,N_5745);
nand U5987 (N_5987,N_5543,N_5707);
and U5988 (N_5988,N_5735,N_5723);
xnor U5989 (N_5989,N_5553,N_5633);
nand U5990 (N_5990,N_5574,N_5516);
and U5991 (N_5991,N_5679,N_5625);
or U5992 (N_5992,N_5733,N_5710);
and U5993 (N_5993,N_5584,N_5651);
and U5994 (N_5994,N_5616,N_5578);
and U5995 (N_5995,N_5625,N_5711);
xor U5996 (N_5996,N_5723,N_5616);
and U5997 (N_5997,N_5511,N_5534);
nand U5998 (N_5998,N_5591,N_5692);
and U5999 (N_5999,N_5514,N_5709);
and U6000 (N_6000,N_5886,N_5786);
nand U6001 (N_6001,N_5806,N_5803);
nand U6002 (N_6002,N_5938,N_5773);
and U6003 (N_6003,N_5812,N_5889);
nor U6004 (N_6004,N_5999,N_5972);
nand U6005 (N_6005,N_5960,N_5827);
and U6006 (N_6006,N_5768,N_5922);
and U6007 (N_6007,N_5897,N_5967);
or U6008 (N_6008,N_5787,N_5893);
or U6009 (N_6009,N_5823,N_5840);
or U6010 (N_6010,N_5920,N_5849);
nand U6011 (N_6011,N_5791,N_5944);
or U6012 (N_6012,N_5924,N_5935);
and U6013 (N_6013,N_5921,N_5801);
xnor U6014 (N_6014,N_5814,N_5983);
nor U6015 (N_6015,N_5951,N_5809);
xor U6016 (N_6016,N_5813,N_5961);
nor U6017 (N_6017,N_5928,N_5973);
xor U6018 (N_6018,N_5887,N_5871);
nand U6019 (N_6019,N_5923,N_5764);
nand U6020 (N_6020,N_5978,N_5866);
nand U6021 (N_6021,N_5877,N_5789);
and U6022 (N_6022,N_5971,N_5891);
or U6023 (N_6023,N_5955,N_5766);
or U6024 (N_6024,N_5908,N_5865);
nor U6025 (N_6025,N_5947,N_5900);
nand U6026 (N_6026,N_5868,N_5847);
nor U6027 (N_6027,N_5784,N_5909);
xor U6028 (N_6028,N_5850,N_5800);
xor U6029 (N_6029,N_5763,N_5846);
or U6030 (N_6030,N_5883,N_5892);
nor U6031 (N_6031,N_5986,N_5838);
nor U6032 (N_6032,N_5862,N_5925);
and U6033 (N_6033,N_5761,N_5844);
nand U6034 (N_6034,N_5918,N_5941);
nor U6035 (N_6035,N_5762,N_5911);
xnor U6036 (N_6036,N_5952,N_5811);
or U6037 (N_6037,N_5832,N_5851);
nand U6038 (N_6038,N_5959,N_5898);
or U6039 (N_6039,N_5818,N_5817);
and U6040 (N_6040,N_5962,N_5772);
nor U6041 (N_6041,N_5853,N_5807);
or U6042 (N_6042,N_5836,N_5993);
xor U6043 (N_6043,N_5954,N_5808);
xnor U6044 (N_6044,N_5802,N_5859);
or U6045 (N_6045,N_5948,N_5881);
or U6046 (N_6046,N_5899,N_5816);
nor U6047 (N_6047,N_5781,N_5869);
and U6048 (N_6048,N_5863,N_5839);
or U6049 (N_6049,N_5906,N_5828);
nand U6050 (N_6050,N_5820,N_5867);
nand U6051 (N_6051,N_5917,N_5966);
and U6052 (N_6052,N_5824,N_5919);
and U6053 (N_6053,N_5884,N_5970);
or U6054 (N_6054,N_5937,N_5785);
or U6055 (N_6055,N_5930,N_5907);
or U6056 (N_6056,N_5984,N_5777);
xnor U6057 (N_6057,N_5751,N_5934);
nand U6058 (N_6058,N_5979,N_5914);
or U6059 (N_6059,N_5950,N_5957);
or U6060 (N_6060,N_5991,N_5878);
xnor U6061 (N_6061,N_5830,N_5780);
or U6062 (N_6062,N_5890,N_5776);
xor U6063 (N_6063,N_5874,N_5754);
nor U6064 (N_6064,N_5974,N_5858);
xor U6065 (N_6065,N_5775,N_5799);
nor U6066 (N_6066,N_5942,N_5805);
or U6067 (N_6067,N_5852,N_5931);
nor U6068 (N_6068,N_5804,N_5835);
xor U6069 (N_6069,N_5992,N_5760);
xor U6070 (N_6070,N_5879,N_5774);
or U6071 (N_6071,N_5753,N_5940);
nand U6072 (N_6072,N_5755,N_5997);
and U6073 (N_6073,N_5793,N_5896);
or U6074 (N_6074,N_5821,N_5829);
or U6075 (N_6075,N_5790,N_5756);
nand U6076 (N_6076,N_5822,N_5913);
xnor U6077 (N_6077,N_5904,N_5943);
nor U6078 (N_6078,N_5965,N_5825);
xnor U6079 (N_6079,N_5949,N_5982);
or U6080 (N_6080,N_5988,N_5985);
xor U6081 (N_6081,N_5998,N_5882);
and U6082 (N_6082,N_5953,N_5765);
xnor U6083 (N_6083,N_5870,N_5946);
nor U6084 (N_6084,N_5905,N_5956);
or U6085 (N_6085,N_5770,N_5758);
or U6086 (N_6086,N_5927,N_5842);
and U6087 (N_6087,N_5888,N_5903);
nand U6088 (N_6088,N_5788,N_5980);
nand U6089 (N_6089,N_5994,N_5861);
xor U6090 (N_6090,N_5932,N_5769);
nor U6091 (N_6091,N_5841,N_5834);
xnor U6092 (N_6092,N_5860,N_5778);
nor U6093 (N_6093,N_5855,N_5963);
xor U6094 (N_6094,N_5767,N_5771);
xnor U6095 (N_6095,N_5873,N_5936);
xor U6096 (N_6096,N_5990,N_5783);
nand U6097 (N_6097,N_5996,N_5857);
xnor U6098 (N_6098,N_5989,N_5782);
and U6099 (N_6099,N_5969,N_5964);
or U6100 (N_6100,N_5958,N_5926);
nand U6101 (N_6101,N_5915,N_5976);
nand U6102 (N_6102,N_5779,N_5872);
nand U6103 (N_6103,N_5981,N_5752);
xnor U6104 (N_6104,N_5875,N_5880);
or U6105 (N_6105,N_5831,N_5819);
nor U6106 (N_6106,N_5810,N_5876);
nand U6107 (N_6107,N_5902,N_5895);
xor U6108 (N_6108,N_5833,N_5916);
nor U6109 (N_6109,N_5794,N_5796);
xor U6110 (N_6110,N_5856,N_5848);
nor U6111 (N_6111,N_5995,N_5933);
nor U6112 (N_6112,N_5759,N_5987);
or U6113 (N_6113,N_5843,N_5977);
nand U6114 (N_6114,N_5910,N_5968);
or U6115 (N_6115,N_5864,N_5885);
xnor U6116 (N_6116,N_5854,N_5826);
xor U6117 (N_6117,N_5975,N_5795);
nand U6118 (N_6118,N_5945,N_5792);
nor U6119 (N_6119,N_5815,N_5901);
nand U6120 (N_6120,N_5750,N_5757);
and U6121 (N_6121,N_5939,N_5912);
nor U6122 (N_6122,N_5894,N_5929);
and U6123 (N_6123,N_5837,N_5845);
nand U6124 (N_6124,N_5797,N_5798);
xor U6125 (N_6125,N_5967,N_5835);
or U6126 (N_6126,N_5780,N_5988);
nand U6127 (N_6127,N_5924,N_5867);
and U6128 (N_6128,N_5920,N_5952);
xnor U6129 (N_6129,N_5762,N_5961);
nand U6130 (N_6130,N_5832,N_5807);
xor U6131 (N_6131,N_5920,N_5901);
xor U6132 (N_6132,N_5789,N_5826);
and U6133 (N_6133,N_5928,N_5819);
and U6134 (N_6134,N_5855,N_5773);
nand U6135 (N_6135,N_5927,N_5987);
or U6136 (N_6136,N_5911,N_5898);
nor U6137 (N_6137,N_5993,N_5899);
nand U6138 (N_6138,N_5924,N_5997);
nor U6139 (N_6139,N_5769,N_5777);
and U6140 (N_6140,N_5989,N_5896);
nor U6141 (N_6141,N_5853,N_5886);
and U6142 (N_6142,N_5752,N_5911);
nand U6143 (N_6143,N_5784,N_5932);
nand U6144 (N_6144,N_5925,N_5905);
nand U6145 (N_6145,N_5988,N_5752);
nor U6146 (N_6146,N_5787,N_5926);
or U6147 (N_6147,N_5791,N_5794);
xnor U6148 (N_6148,N_5951,N_5767);
nor U6149 (N_6149,N_5945,N_5972);
nand U6150 (N_6150,N_5998,N_5878);
nor U6151 (N_6151,N_5832,N_5978);
nand U6152 (N_6152,N_5869,N_5810);
or U6153 (N_6153,N_5950,N_5903);
or U6154 (N_6154,N_5851,N_5880);
nor U6155 (N_6155,N_5790,N_5780);
xnor U6156 (N_6156,N_5930,N_5946);
nand U6157 (N_6157,N_5803,N_5775);
and U6158 (N_6158,N_5983,N_5939);
and U6159 (N_6159,N_5976,N_5804);
nor U6160 (N_6160,N_5851,N_5775);
and U6161 (N_6161,N_5963,N_5913);
and U6162 (N_6162,N_5771,N_5840);
or U6163 (N_6163,N_5851,N_5763);
and U6164 (N_6164,N_5814,N_5789);
and U6165 (N_6165,N_5914,N_5967);
or U6166 (N_6166,N_5810,N_5757);
or U6167 (N_6167,N_5982,N_5993);
xor U6168 (N_6168,N_5867,N_5970);
nand U6169 (N_6169,N_5776,N_5955);
xnor U6170 (N_6170,N_5829,N_5803);
xor U6171 (N_6171,N_5788,N_5835);
or U6172 (N_6172,N_5865,N_5994);
nor U6173 (N_6173,N_5783,N_5931);
and U6174 (N_6174,N_5895,N_5871);
nor U6175 (N_6175,N_5844,N_5914);
xnor U6176 (N_6176,N_5932,N_5855);
nand U6177 (N_6177,N_5851,N_5850);
xnor U6178 (N_6178,N_5868,N_5844);
nor U6179 (N_6179,N_5937,N_5769);
or U6180 (N_6180,N_5813,N_5817);
and U6181 (N_6181,N_5971,N_5932);
and U6182 (N_6182,N_5999,N_5918);
nand U6183 (N_6183,N_5893,N_5793);
and U6184 (N_6184,N_5758,N_5884);
and U6185 (N_6185,N_5992,N_5793);
nand U6186 (N_6186,N_5852,N_5939);
nand U6187 (N_6187,N_5795,N_5853);
and U6188 (N_6188,N_5964,N_5847);
xor U6189 (N_6189,N_5862,N_5843);
and U6190 (N_6190,N_5857,N_5760);
and U6191 (N_6191,N_5896,N_5919);
xnor U6192 (N_6192,N_5975,N_5964);
xnor U6193 (N_6193,N_5779,N_5863);
and U6194 (N_6194,N_5910,N_5772);
nor U6195 (N_6195,N_5906,N_5895);
nor U6196 (N_6196,N_5761,N_5960);
or U6197 (N_6197,N_5828,N_5990);
and U6198 (N_6198,N_5812,N_5940);
nor U6199 (N_6199,N_5996,N_5850);
or U6200 (N_6200,N_5817,N_5901);
xor U6201 (N_6201,N_5989,N_5919);
or U6202 (N_6202,N_5978,N_5802);
or U6203 (N_6203,N_5814,N_5816);
xnor U6204 (N_6204,N_5994,N_5807);
or U6205 (N_6205,N_5939,N_5943);
and U6206 (N_6206,N_5992,N_5984);
xor U6207 (N_6207,N_5819,N_5800);
xnor U6208 (N_6208,N_5773,N_5834);
xor U6209 (N_6209,N_5892,N_5866);
or U6210 (N_6210,N_5893,N_5780);
xnor U6211 (N_6211,N_5878,N_5978);
xnor U6212 (N_6212,N_5893,N_5956);
and U6213 (N_6213,N_5887,N_5851);
or U6214 (N_6214,N_5967,N_5768);
or U6215 (N_6215,N_5853,N_5969);
nor U6216 (N_6216,N_5839,N_5938);
or U6217 (N_6217,N_5814,N_5910);
and U6218 (N_6218,N_5809,N_5980);
or U6219 (N_6219,N_5859,N_5983);
xor U6220 (N_6220,N_5829,N_5801);
xnor U6221 (N_6221,N_5880,N_5966);
xor U6222 (N_6222,N_5897,N_5753);
nand U6223 (N_6223,N_5929,N_5944);
xnor U6224 (N_6224,N_5940,N_5981);
nor U6225 (N_6225,N_5819,N_5769);
nand U6226 (N_6226,N_5992,N_5824);
and U6227 (N_6227,N_5877,N_5926);
or U6228 (N_6228,N_5840,N_5847);
xnor U6229 (N_6229,N_5965,N_5997);
nand U6230 (N_6230,N_5750,N_5888);
or U6231 (N_6231,N_5750,N_5890);
or U6232 (N_6232,N_5991,N_5837);
xnor U6233 (N_6233,N_5892,N_5943);
xnor U6234 (N_6234,N_5750,N_5782);
or U6235 (N_6235,N_5976,N_5774);
or U6236 (N_6236,N_5834,N_5873);
nand U6237 (N_6237,N_5816,N_5900);
or U6238 (N_6238,N_5946,N_5791);
nand U6239 (N_6239,N_5819,N_5840);
nor U6240 (N_6240,N_5824,N_5875);
and U6241 (N_6241,N_5979,N_5893);
xor U6242 (N_6242,N_5757,N_5828);
nand U6243 (N_6243,N_5919,N_5878);
or U6244 (N_6244,N_5763,N_5986);
nor U6245 (N_6245,N_5776,N_5923);
nor U6246 (N_6246,N_5937,N_5971);
nor U6247 (N_6247,N_5876,N_5893);
and U6248 (N_6248,N_5810,N_5916);
xnor U6249 (N_6249,N_5893,N_5781);
or U6250 (N_6250,N_6199,N_6220);
xnor U6251 (N_6251,N_6024,N_6080);
xor U6252 (N_6252,N_6202,N_6093);
nand U6253 (N_6253,N_6246,N_6168);
or U6254 (N_6254,N_6060,N_6205);
nor U6255 (N_6255,N_6057,N_6111);
and U6256 (N_6256,N_6137,N_6065);
nor U6257 (N_6257,N_6023,N_6110);
and U6258 (N_6258,N_6094,N_6142);
or U6259 (N_6259,N_6006,N_6163);
and U6260 (N_6260,N_6003,N_6236);
or U6261 (N_6261,N_6122,N_6095);
and U6262 (N_6262,N_6174,N_6155);
or U6263 (N_6263,N_6054,N_6182);
nor U6264 (N_6264,N_6209,N_6156);
nor U6265 (N_6265,N_6154,N_6249);
xnor U6266 (N_6266,N_6063,N_6153);
xor U6267 (N_6267,N_6086,N_6184);
and U6268 (N_6268,N_6067,N_6196);
and U6269 (N_6269,N_6071,N_6005);
xnor U6270 (N_6270,N_6096,N_6077);
nand U6271 (N_6271,N_6058,N_6218);
and U6272 (N_6272,N_6195,N_6130);
and U6273 (N_6273,N_6239,N_6053);
and U6274 (N_6274,N_6243,N_6066);
xor U6275 (N_6275,N_6172,N_6132);
and U6276 (N_6276,N_6148,N_6121);
nand U6277 (N_6277,N_6138,N_6007);
nor U6278 (N_6278,N_6244,N_6165);
and U6279 (N_6279,N_6192,N_6079);
nor U6280 (N_6280,N_6028,N_6129);
xor U6281 (N_6281,N_6048,N_6151);
or U6282 (N_6282,N_6046,N_6045);
and U6283 (N_6283,N_6128,N_6189);
or U6284 (N_6284,N_6108,N_6204);
xnor U6285 (N_6285,N_6139,N_6029);
and U6286 (N_6286,N_6207,N_6185);
nor U6287 (N_6287,N_6113,N_6214);
or U6288 (N_6288,N_6087,N_6090);
or U6289 (N_6289,N_6149,N_6124);
nand U6290 (N_6290,N_6183,N_6242);
or U6291 (N_6291,N_6186,N_6241);
nand U6292 (N_6292,N_6098,N_6061);
or U6293 (N_6293,N_6064,N_6198);
and U6294 (N_6294,N_6038,N_6103);
nor U6295 (N_6295,N_6041,N_6167);
and U6296 (N_6296,N_6009,N_6247);
or U6297 (N_6297,N_6179,N_6008);
nand U6298 (N_6298,N_6015,N_6216);
and U6299 (N_6299,N_6131,N_6112);
and U6300 (N_6300,N_6092,N_6193);
nor U6301 (N_6301,N_6194,N_6187);
nor U6302 (N_6302,N_6225,N_6208);
and U6303 (N_6303,N_6200,N_6070);
and U6304 (N_6304,N_6245,N_6085);
nor U6305 (N_6305,N_6089,N_6036);
nor U6306 (N_6306,N_6176,N_6178);
nand U6307 (N_6307,N_6030,N_6211);
xnor U6308 (N_6308,N_6217,N_6160);
nand U6309 (N_6309,N_6232,N_6221);
xor U6310 (N_6310,N_6206,N_6016);
and U6311 (N_6311,N_6115,N_6039);
xnor U6312 (N_6312,N_6072,N_6091);
nor U6313 (N_6313,N_6099,N_6040);
xnor U6314 (N_6314,N_6147,N_6228);
or U6315 (N_6315,N_6177,N_6224);
xnor U6316 (N_6316,N_6166,N_6049);
nand U6317 (N_6317,N_6031,N_6120);
nor U6318 (N_6318,N_6222,N_6173);
nor U6319 (N_6319,N_6034,N_6033);
and U6320 (N_6320,N_6068,N_6170);
nand U6321 (N_6321,N_6237,N_6180);
or U6322 (N_6322,N_6078,N_6227);
or U6323 (N_6323,N_6106,N_6226);
xnor U6324 (N_6324,N_6162,N_6010);
xor U6325 (N_6325,N_6000,N_6025);
and U6326 (N_6326,N_6125,N_6169);
nand U6327 (N_6327,N_6083,N_6141);
and U6328 (N_6328,N_6118,N_6074);
nand U6329 (N_6329,N_6215,N_6104);
xnor U6330 (N_6330,N_6212,N_6026);
or U6331 (N_6331,N_6145,N_6144);
xnor U6332 (N_6332,N_6002,N_6011);
xor U6333 (N_6333,N_6001,N_6088);
nand U6334 (N_6334,N_6117,N_6157);
or U6335 (N_6335,N_6059,N_6107);
xnor U6336 (N_6336,N_6219,N_6234);
nand U6337 (N_6337,N_6019,N_6159);
xnor U6338 (N_6338,N_6126,N_6109);
or U6339 (N_6339,N_6047,N_6235);
xor U6340 (N_6340,N_6100,N_6081);
xor U6341 (N_6341,N_6062,N_6014);
or U6342 (N_6342,N_6230,N_6140);
or U6343 (N_6343,N_6055,N_6032);
xor U6344 (N_6344,N_6119,N_6134);
nand U6345 (N_6345,N_6056,N_6136);
nor U6346 (N_6346,N_6042,N_6020);
nand U6347 (N_6347,N_6229,N_6210);
nand U6348 (N_6348,N_6158,N_6013);
nor U6349 (N_6349,N_6043,N_6123);
or U6350 (N_6350,N_6181,N_6191);
nand U6351 (N_6351,N_6175,N_6052);
and U6352 (N_6352,N_6150,N_6051);
nor U6353 (N_6353,N_6197,N_6116);
nor U6354 (N_6354,N_6240,N_6233);
xnor U6355 (N_6355,N_6143,N_6133);
and U6356 (N_6356,N_6084,N_6073);
nand U6357 (N_6357,N_6018,N_6188);
nand U6358 (N_6358,N_6105,N_6135);
or U6359 (N_6359,N_6161,N_6213);
xor U6360 (N_6360,N_6044,N_6201);
nand U6361 (N_6361,N_6127,N_6203);
nand U6362 (N_6362,N_6004,N_6238);
or U6363 (N_6363,N_6248,N_6069);
nor U6364 (N_6364,N_6101,N_6146);
nor U6365 (N_6365,N_6102,N_6190);
and U6366 (N_6366,N_6223,N_6075);
and U6367 (N_6367,N_6164,N_6012);
and U6368 (N_6368,N_6027,N_6076);
nand U6369 (N_6369,N_6037,N_6097);
and U6370 (N_6370,N_6114,N_6171);
nor U6371 (N_6371,N_6152,N_6050);
nor U6372 (N_6372,N_6022,N_6017);
or U6373 (N_6373,N_6231,N_6082);
nor U6374 (N_6374,N_6035,N_6021);
nand U6375 (N_6375,N_6217,N_6181);
xnor U6376 (N_6376,N_6085,N_6019);
or U6377 (N_6377,N_6155,N_6040);
nand U6378 (N_6378,N_6161,N_6166);
nand U6379 (N_6379,N_6171,N_6145);
nand U6380 (N_6380,N_6089,N_6072);
or U6381 (N_6381,N_6094,N_6026);
and U6382 (N_6382,N_6041,N_6080);
nor U6383 (N_6383,N_6172,N_6023);
or U6384 (N_6384,N_6223,N_6100);
or U6385 (N_6385,N_6172,N_6011);
nand U6386 (N_6386,N_6201,N_6239);
or U6387 (N_6387,N_6241,N_6026);
nand U6388 (N_6388,N_6048,N_6081);
and U6389 (N_6389,N_6214,N_6194);
xor U6390 (N_6390,N_6236,N_6070);
xor U6391 (N_6391,N_6111,N_6155);
nor U6392 (N_6392,N_6046,N_6021);
nor U6393 (N_6393,N_6136,N_6025);
or U6394 (N_6394,N_6101,N_6106);
xnor U6395 (N_6395,N_6106,N_6222);
and U6396 (N_6396,N_6163,N_6241);
nor U6397 (N_6397,N_6090,N_6198);
nor U6398 (N_6398,N_6238,N_6228);
nand U6399 (N_6399,N_6054,N_6088);
and U6400 (N_6400,N_6220,N_6189);
and U6401 (N_6401,N_6076,N_6016);
and U6402 (N_6402,N_6126,N_6143);
and U6403 (N_6403,N_6185,N_6117);
nand U6404 (N_6404,N_6231,N_6227);
nor U6405 (N_6405,N_6194,N_6059);
nor U6406 (N_6406,N_6061,N_6145);
xnor U6407 (N_6407,N_6189,N_6152);
xnor U6408 (N_6408,N_6008,N_6027);
nand U6409 (N_6409,N_6024,N_6084);
or U6410 (N_6410,N_6121,N_6149);
or U6411 (N_6411,N_6035,N_6141);
nor U6412 (N_6412,N_6197,N_6158);
nand U6413 (N_6413,N_6212,N_6130);
and U6414 (N_6414,N_6012,N_6025);
xnor U6415 (N_6415,N_6051,N_6184);
nor U6416 (N_6416,N_6103,N_6170);
nor U6417 (N_6417,N_6200,N_6017);
xnor U6418 (N_6418,N_6126,N_6015);
or U6419 (N_6419,N_6241,N_6071);
or U6420 (N_6420,N_6155,N_6102);
xor U6421 (N_6421,N_6008,N_6089);
nand U6422 (N_6422,N_6219,N_6032);
nor U6423 (N_6423,N_6128,N_6076);
or U6424 (N_6424,N_6237,N_6227);
nor U6425 (N_6425,N_6219,N_6158);
nand U6426 (N_6426,N_6005,N_6148);
xnor U6427 (N_6427,N_6025,N_6210);
nand U6428 (N_6428,N_6067,N_6118);
nand U6429 (N_6429,N_6113,N_6111);
and U6430 (N_6430,N_6056,N_6133);
or U6431 (N_6431,N_6211,N_6226);
xnor U6432 (N_6432,N_6248,N_6165);
nand U6433 (N_6433,N_6124,N_6206);
nor U6434 (N_6434,N_6180,N_6201);
xor U6435 (N_6435,N_6083,N_6066);
xor U6436 (N_6436,N_6093,N_6094);
xnor U6437 (N_6437,N_6244,N_6167);
and U6438 (N_6438,N_6230,N_6094);
or U6439 (N_6439,N_6134,N_6218);
or U6440 (N_6440,N_6187,N_6220);
or U6441 (N_6441,N_6098,N_6020);
xor U6442 (N_6442,N_6173,N_6108);
nor U6443 (N_6443,N_6014,N_6039);
xor U6444 (N_6444,N_6067,N_6061);
and U6445 (N_6445,N_6213,N_6226);
and U6446 (N_6446,N_6175,N_6011);
and U6447 (N_6447,N_6231,N_6124);
xnor U6448 (N_6448,N_6108,N_6066);
nor U6449 (N_6449,N_6124,N_6177);
xor U6450 (N_6450,N_6172,N_6070);
xnor U6451 (N_6451,N_6121,N_6200);
nor U6452 (N_6452,N_6209,N_6123);
nand U6453 (N_6453,N_6073,N_6180);
or U6454 (N_6454,N_6091,N_6163);
or U6455 (N_6455,N_6116,N_6075);
or U6456 (N_6456,N_6004,N_6217);
xnor U6457 (N_6457,N_6033,N_6213);
or U6458 (N_6458,N_6222,N_6087);
nand U6459 (N_6459,N_6199,N_6072);
nor U6460 (N_6460,N_6101,N_6076);
and U6461 (N_6461,N_6054,N_6147);
nand U6462 (N_6462,N_6055,N_6196);
or U6463 (N_6463,N_6020,N_6192);
and U6464 (N_6464,N_6064,N_6170);
nand U6465 (N_6465,N_6167,N_6011);
nor U6466 (N_6466,N_6189,N_6215);
or U6467 (N_6467,N_6166,N_6177);
and U6468 (N_6468,N_6130,N_6245);
and U6469 (N_6469,N_6044,N_6121);
xor U6470 (N_6470,N_6029,N_6158);
or U6471 (N_6471,N_6159,N_6018);
or U6472 (N_6472,N_6015,N_6050);
xor U6473 (N_6473,N_6241,N_6200);
and U6474 (N_6474,N_6110,N_6009);
or U6475 (N_6475,N_6189,N_6065);
and U6476 (N_6476,N_6103,N_6175);
and U6477 (N_6477,N_6172,N_6092);
nor U6478 (N_6478,N_6066,N_6105);
xor U6479 (N_6479,N_6112,N_6123);
or U6480 (N_6480,N_6102,N_6175);
or U6481 (N_6481,N_6007,N_6235);
xnor U6482 (N_6482,N_6113,N_6229);
or U6483 (N_6483,N_6238,N_6061);
and U6484 (N_6484,N_6041,N_6170);
nand U6485 (N_6485,N_6086,N_6158);
xor U6486 (N_6486,N_6238,N_6138);
and U6487 (N_6487,N_6126,N_6100);
nand U6488 (N_6488,N_6052,N_6042);
xnor U6489 (N_6489,N_6238,N_6043);
xnor U6490 (N_6490,N_6094,N_6132);
nand U6491 (N_6491,N_6230,N_6145);
nor U6492 (N_6492,N_6221,N_6057);
xnor U6493 (N_6493,N_6179,N_6228);
or U6494 (N_6494,N_6089,N_6065);
or U6495 (N_6495,N_6190,N_6012);
nand U6496 (N_6496,N_6249,N_6113);
nor U6497 (N_6497,N_6005,N_6174);
nor U6498 (N_6498,N_6112,N_6001);
or U6499 (N_6499,N_6108,N_6062);
or U6500 (N_6500,N_6367,N_6336);
xor U6501 (N_6501,N_6423,N_6374);
and U6502 (N_6502,N_6252,N_6340);
or U6503 (N_6503,N_6314,N_6344);
or U6504 (N_6504,N_6315,N_6408);
nor U6505 (N_6505,N_6273,N_6468);
xnor U6506 (N_6506,N_6381,N_6259);
xor U6507 (N_6507,N_6432,N_6452);
xor U6508 (N_6508,N_6473,N_6339);
nand U6509 (N_6509,N_6390,N_6364);
and U6510 (N_6510,N_6430,N_6475);
and U6511 (N_6511,N_6351,N_6316);
nand U6512 (N_6512,N_6376,N_6328);
and U6513 (N_6513,N_6458,N_6282);
xor U6514 (N_6514,N_6288,N_6426);
nand U6515 (N_6515,N_6378,N_6298);
or U6516 (N_6516,N_6299,N_6280);
xor U6517 (N_6517,N_6379,N_6386);
or U6518 (N_6518,N_6313,N_6312);
xor U6519 (N_6519,N_6361,N_6333);
and U6520 (N_6520,N_6261,N_6391);
or U6521 (N_6521,N_6493,N_6255);
and U6522 (N_6522,N_6472,N_6420);
nand U6523 (N_6523,N_6264,N_6384);
nor U6524 (N_6524,N_6284,N_6440);
nor U6525 (N_6525,N_6331,N_6485);
nand U6526 (N_6526,N_6251,N_6360);
xnor U6527 (N_6527,N_6466,N_6429);
and U6528 (N_6528,N_6478,N_6303);
nand U6529 (N_6529,N_6447,N_6395);
xor U6530 (N_6530,N_6304,N_6460);
nand U6531 (N_6531,N_6488,N_6349);
xor U6532 (N_6532,N_6301,N_6355);
nor U6533 (N_6533,N_6276,N_6393);
xor U6534 (N_6534,N_6383,N_6289);
nand U6535 (N_6535,N_6467,N_6327);
xnor U6536 (N_6536,N_6256,N_6266);
and U6537 (N_6537,N_6342,N_6375);
nor U6538 (N_6538,N_6490,N_6291);
and U6539 (N_6539,N_6491,N_6498);
nand U6540 (N_6540,N_6449,N_6250);
nor U6541 (N_6541,N_6320,N_6334);
or U6542 (N_6542,N_6428,N_6437);
or U6543 (N_6543,N_6330,N_6354);
nand U6544 (N_6544,N_6456,N_6418);
nand U6545 (N_6545,N_6396,N_6308);
and U6546 (N_6546,N_6325,N_6403);
nand U6547 (N_6547,N_6380,N_6495);
nand U6548 (N_6548,N_6319,N_6404);
or U6549 (N_6549,N_6335,N_6450);
xor U6550 (N_6550,N_6347,N_6425);
or U6551 (N_6551,N_6494,N_6496);
nand U6552 (N_6552,N_6463,N_6269);
nor U6553 (N_6553,N_6388,N_6372);
or U6554 (N_6554,N_6323,N_6353);
or U6555 (N_6555,N_6332,N_6476);
nor U6556 (N_6556,N_6318,N_6369);
or U6557 (N_6557,N_6497,N_6435);
xnor U6558 (N_6558,N_6302,N_6482);
or U6559 (N_6559,N_6471,N_6457);
nand U6560 (N_6560,N_6442,N_6492);
xnor U6561 (N_6561,N_6479,N_6281);
and U6562 (N_6562,N_6489,N_6270);
xor U6563 (N_6563,N_6343,N_6401);
or U6564 (N_6564,N_6477,N_6277);
or U6565 (N_6565,N_6398,N_6337);
nor U6566 (N_6566,N_6368,N_6346);
nor U6567 (N_6567,N_6263,N_6499);
or U6568 (N_6568,N_6394,N_6387);
and U6569 (N_6569,N_6417,N_6412);
or U6570 (N_6570,N_6271,N_6258);
and U6571 (N_6571,N_6300,N_6462);
and U6572 (N_6572,N_6406,N_6309);
nand U6573 (N_6573,N_6483,N_6373);
nand U6574 (N_6574,N_6285,N_6464);
xnor U6575 (N_6575,N_6416,N_6371);
xnor U6576 (N_6576,N_6307,N_6257);
nor U6577 (N_6577,N_6451,N_6326);
and U6578 (N_6578,N_6441,N_6274);
nor U6579 (N_6579,N_6287,N_6366);
xor U6580 (N_6580,N_6352,N_6292);
xor U6581 (N_6581,N_6310,N_6350);
or U6582 (N_6582,N_6415,N_6348);
nand U6583 (N_6583,N_6317,N_6265);
xnor U6584 (N_6584,N_6283,N_6290);
and U6585 (N_6585,N_6392,N_6311);
nand U6586 (N_6586,N_6296,N_6419);
nor U6587 (N_6587,N_6487,N_6357);
nor U6588 (N_6588,N_6443,N_6422);
xnor U6589 (N_6589,N_6329,N_6397);
or U6590 (N_6590,N_6409,N_6286);
nor U6591 (N_6591,N_6474,N_6321);
and U6592 (N_6592,N_6481,N_6254);
nor U6593 (N_6593,N_6262,N_6446);
nand U6594 (N_6594,N_6434,N_6445);
and U6595 (N_6595,N_6453,N_6358);
xnor U6596 (N_6596,N_6444,N_6370);
or U6597 (N_6597,N_6278,N_6385);
nor U6598 (N_6598,N_6433,N_6253);
xor U6599 (N_6599,N_6469,N_6427);
nand U6600 (N_6600,N_6407,N_6338);
nand U6601 (N_6601,N_6402,N_6341);
nor U6602 (N_6602,N_6297,N_6356);
xnor U6603 (N_6603,N_6414,N_6324);
nand U6604 (N_6604,N_6470,N_6382);
nor U6605 (N_6605,N_6454,N_6399);
and U6606 (N_6606,N_6459,N_6365);
nor U6607 (N_6607,N_6438,N_6322);
or U6608 (N_6608,N_6480,N_6424);
xor U6609 (N_6609,N_6306,N_6279);
xnor U6610 (N_6610,N_6421,N_6484);
and U6611 (N_6611,N_6405,N_6400);
or U6612 (N_6612,N_6448,N_6486);
nand U6613 (N_6613,N_6389,N_6436);
nor U6614 (N_6614,N_6305,N_6294);
xnor U6615 (N_6615,N_6377,N_6410);
and U6616 (N_6616,N_6268,N_6431);
nor U6617 (N_6617,N_6295,N_6363);
nand U6618 (N_6618,N_6260,N_6455);
nor U6619 (N_6619,N_6465,N_6267);
nor U6620 (N_6620,N_6413,N_6345);
or U6621 (N_6621,N_6272,N_6362);
nand U6622 (N_6622,N_6359,N_6461);
or U6623 (N_6623,N_6411,N_6293);
or U6624 (N_6624,N_6439,N_6275);
xnor U6625 (N_6625,N_6460,N_6281);
or U6626 (N_6626,N_6426,N_6466);
xor U6627 (N_6627,N_6314,N_6450);
and U6628 (N_6628,N_6374,N_6329);
or U6629 (N_6629,N_6357,N_6421);
nand U6630 (N_6630,N_6375,N_6311);
or U6631 (N_6631,N_6489,N_6308);
or U6632 (N_6632,N_6284,N_6335);
nand U6633 (N_6633,N_6361,N_6369);
nor U6634 (N_6634,N_6272,N_6281);
nor U6635 (N_6635,N_6482,N_6295);
nand U6636 (N_6636,N_6314,N_6271);
or U6637 (N_6637,N_6266,N_6297);
and U6638 (N_6638,N_6464,N_6459);
nor U6639 (N_6639,N_6363,N_6482);
and U6640 (N_6640,N_6266,N_6377);
nor U6641 (N_6641,N_6464,N_6460);
xor U6642 (N_6642,N_6268,N_6444);
and U6643 (N_6643,N_6346,N_6311);
or U6644 (N_6644,N_6278,N_6426);
and U6645 (N_6645,N_6473,N_6303);
nand U6646 (N_6646,N_6311,N_6283);
nor U6647 (N_6647,N_6397,N_6339);
nand U6648 (N_6648,N_6340,N_6496);
nand U6649 (N_6649,N_6324,N_6408);
xor U6650 (N_6650,N_6440,N_6334);
or U6651 (N_6651,N_6279,N_6269);
nand U6652 (N_6652,N_6483,N_6347);
nor U6653 (N_6653,N_6481,N_6397);
and U6654 (N_6654,N_6463,N_6351);
or U6655 (N_6655,N_6376,N_6492);
nor U6656 (N_6656,N_6453,N_6360);
nor U6657 (N_6657,N_6271,N_6430);
and U6658 (N_6658,N_6314,N_6474);
and U6659 (N_6659,N_6402,N_6322);
and U6660 (N_6660,N_6280,N_6346);
nor U6661 (N_6661,N_6413,N_6273);
nor U6662 (N_6662,N_6366,N_6484);
nor U6663 (N_6663,N_6422,N_6456);
nand U6664 (N_6664,N_6332,N_6324);
and U6665 (N_6665,N_6322,N_6413);
xor U6666 (N_6666,N_6338,N_6253);
nand U6667 (N_6667,N_6326,N_6313);
and U6668 (N_6668,N_6409,N_6313);
nor U6669 (N_6669,N_6296,N_6455);
or U6670 (N_6670,N_6254,N_6333);
and U6671 (N_6671,N_6324,N_6377);
or U6672 (N_6672,N_6483,N_6339);
xnor U6673 (N_6673,N_6438,N_6475);
nand U6674 (N_6674,N_6473,N_6265);
nor U6675 (N_6675,N_6265,N_6359);
xnor U6676 (N_6676,N_6461,N_6370);
and U6677 (N_6677,N_6453,N_6316);
nor U6678 (N_6678,N_6375,N_6309);
xor U6679 (N_6679,N_6414,N_6499);
nor U6680 (N_6680,N_6274,N_6320);
or U6681 (N_6681,N_6276,N_6432);
nor U6682 (N_6682,N_6296,N_6362);
nand U6683 (N_6683,N_6295,N_6373);
nor U6684 (N_6684,N_6362,N_6289);
nor U6685 (N_6685,N_6417,N_6360);
nand U6686 (N_6686,N_6359,N_6432);
nand U6687 (N_6687,N_6341,N_6330);
nand U6688 (N_6688,N_6303,N_6298);
nor U6689 (N_6689,N_6283,N_6346);
nand U6690 (N_6690,N_6333,N_6391);
and U6691 (N_6691,N_6349,N_6419);
nand U6692 (N_6692,N_6351,N_6286);
nor U6693 (N_6693,N_6256,N_6444);
nand U6694 (N_6694,N_6298,N_6485);
and U6695 (N_6695,N_6305,N_6298);
nand U6696 (N_6696,N_6315,N_6394);
nand U6697 (N_6697,N_6321,N_6264);
nand U6698 (N_6698,N_6312,N_6480);
nand U6699 (N_6699,N_6437,N_6392);
xor U6700 (N_6700,N_6466,N_6342);
or U6701 (N_6701,N_6470,N_6421);
nor U6702 (N_6702,N_6275,N_6462);
nor U6703 (N_6703,N_6302,N_6272);
xor U6704 (N_6704,N_6488,N_6327);
nand U6705 (N_6705,N_6399,N_6321);
and U6706 (N_6706,N_6321,N_6499);
or U6707 (N_6707,N_6336,N_6253);
nand U6708 (N_6708,N_6255,N_6444);
and U6709 (N_6709,N_6279,N_6442);
nor U6710 (N_6710,N_6447,N_6377);
nand U6711 (N_6711,N_6299,N_6294);
nor U6712 (N_6712,N_6291,N_6416);
or U6713 (N_6713,N_6335,N_6499);
or U6714 (N_6714,N_6322,N_6275);
nand U6715 (N_6715,N_6296,N_6376);
nand U6716 (N_6716,N_6481,N_6439);
or U6717 (N_6717,N_6476,N_6491);
and U6718 (N_6718,N_6411,N_6433);
or U6719 (N_6719,N_6439,N_6435);
or U6720 (N_6720,N_6298,N_6344);
nand U6721 (N_6721,N_6432,N_6461);
nand U6722 (N_6722,N_6318,N_6394);
and U6723 (N_6723,N_6351,N_6288);
nor U6724 (N_6724,N_6358,N_6430);
nor U6725 (N_6725,N_6372,N_6349);
nand U6726 (N_6726,N_6387,N_6433);
xor U6727 (N_6727,N_6327,N_6446);
xnor U6728 (N_6728,N_6478,N_6287);
or U6729 (N_6729,N_6337,N_6378);
xnor U6730 (N_6730,N_6306,N_6431);
and U6731 (N_6731,N_6259,N_6282);
or U6732 (N_6732,N_6423,N_6404);
nor U6733 (N_6733,N_6334,N_6324);
xnor U6734 (N_6734,N_6489,N_6374);
xnor U6735 (N_6735,N_6356,N_6454);
xor U6736 (N_6736,N_6284,N_6414);
nor U6737 (N_6737,N_6320,N_6253);
nand U6738 (N_6738,N_6386,N_6267);
or U6739 (N_6739,N_6372,N_6366);
nand U6740 (N_6740,N_6395,N_6489);
nand U6741 (N_6741,N_6266,N_6313);
nand U6742 (N_6742,N_6404,N_6306);
nand U6743 (N_6743,N_6379,N_6338);
nand U6744 (N_6744,N_6284,N_6460);
nor U6745 (N_6745,N_6419,N_6311);
or U6746 (N_6746,N_6391,N_6343);
xnor U6747 (N_6747,N_6459,N_6452);
nor U6748 (N_6748,N_6454,N_6449);
or U6749 (N_6749,N_6289,N_6283);
xor U6750 (N_6750,N_6724,N_6689);
nand U6751 (N_6751,N_6686,N_6595);
or U6752 (N_6752,N_6588,N_6570);
nand U6753 (N_6753,N_6690,N_6551);
and U6754 (N_6754,N_6587,N_6628);
xnor U6755 (N_6755,N_6531,N_6541);
and U6756 (N_6756,N_6731,N_6610);
or U6757 (N_6757,N_6533,N_6563);
or U6758 (N_6758,N_6516,N_6675);
and U6759 (N_6759,N_6692,N_6561);
and U6760 (N_6760,N_6621,N_6511);
or U6761 (N_6761,N_6627,N_6733);
xor U6762 (N_6762,N_6558,N_6529);
nor U6763 (N_6763,N_6674,N_6723);
nand U6764 (N_6764,N_6712,N_6709);
nand U6765 (N_6765,N_6634,N_6727);
nand U6766 (N_6766,N_6722,N_6737);
and U6767 (N_6767,N_6693,N_6503);
or U6768 (N_6768,N_6636,N_6644);
or U6769 (N_6769,N_6642,N_6713);
and U6770 (N_6770,N_6580,N_6565);
or U6771 (N_6771,N_6645,N_6545);
nor U6772 (N_6772,N_6515,N_6677);
or U6773 (N_6773,N_6547,N_6615);
nand U6774 (N_6774,N_6747,N_6653);
nor U6775 (N_6775,N_6619,N_6654);
nand U6776 (N_6776,N_6743,N_6659);
or U6777 (N_6777,N_6643,N_6656);
nand U6778 (N_6778,N_6520,N_6593);
nand U6779 (N_6779,N_6523,N_6519);
xnor U6780 (N_6780,N_6652,N_6745);
or U6781 (N_6781,N_6602,N_6576);
nor U6782 (N_6782,N_6734,N_6539);
nor U6783 (N_6783,N_6632,N_6666);
or U6784 (N_6784,N_6599,N_6537);
and U6785 (N_6785,N_6566,N_6728);
nand U6786 (N_6786,N_6660,N_6746);
nor U6787 (N_6787,N_6608,N_6741);
xnor U6788 (N_6788,N_6556,N_6742);
xor U6789 (N_6789,N_6639,N_6564);
xor U6790 (N_6790,N_6577,N_6585);
nand U6791 (N_6791,N_6601,N_6646);
xnor U6792 (N_6792,N_6510,N_6518);
nand U6793 (N_6793,N_6597,N_6683);
or U6794 (N_6794,N_6716,N_6504);
or U6795 (N_6795,N_6600,N_6530);
nand U6796 (N_6796,N_6502,N_6676);
xnor U6797 (N_6797,N_6662,N_6586);
nor U6798 (N_6798,N_6552,N_6721);
nor U6799 (N_6799,N_6719,N_6637);
xor U6800 (N_6800,N_6670,N_6631);
nor U6801 (N_6801,N_6679,N_6700);
or U6802 (N_6802,N_6506,N_6657);
and U6803 (N_6803,N_6567,N_6740);
nor U6804 (N_6804,N_6623,N_6549);
nand U6805 (N_6805,N_6574,N_6651);
or U6806 (N_6806,N_6594,N_6612);
and U6807 (N_6807,N_6649,N_6617);
nor U6808 (N_6808,N_6604,N_6698);
nand U6809 (N_6809,N_6535,N_6614);
or U6810 (N_6810,N_6616,N_6629);
nand U6811 (N_6811,N_6553,N_6544);
nor U6812 (N_6812,N_6680,N_6596);
and U6813 (N_6813,N_6702,N_6715);
or U6814 (N_6814,N_6581,N_6592);
nand U6815 (N_6815,N_6582,N_6748);
nor U6816 (N_6816,N_6732,N_6710);
xor U6817 (N_6817,N_6572,N_6671);
and U6818 (N_6818,N_6528,N_6667);
or U6819 (N_6819,N_6684,N_6507);
nor U6820 (N_6820,N_6681,N_6718);
nor U6821 (N_6821,N_6625,N_6707);
or U6822 (N_6822,N_6749,N_6514);
xor U6823 (N_6823,N_6606,N_6687);
xor U6824 (N_6824,N_6609,N_6678);
nor U6825 (N_6825,N_6611,N_6560);
and U6826 (N_6826,N_6682,N_6613);
nor U6827 (N_6827,N_6543,N_6590);
nand U6828 (N_6828,N_6534,N_6501);
nor U6829 (N_6829,N_6697,N_6708);
nand U6830 (N_6830,N_6701,N_6641);
or U6831 (N_6831,N_6550,N_6729);
nor U6832 (N_6832,N_6694,N_6583);
xor U6833 (N_6833,N_6717,N_6532);
and U6834 (N_6834,N_6536,N_6521);
nand U6835 (N_6835,N_6573,N_6562);
or U6836 (N_6836,N_6578,N_6633);
or U6837 (N_6837,N_6735,N_6524);
or U6838 (N_6838,N_6526,N_6720);
nor U6839 (N_6839,N_6665,N_6669);
or U6840 (N_6840,N_6673,N_6569);
and U6841 (N_6841,N_6591,N_6685);
nor U6842 (N_6842,N_6726,N_6618);
xor U6843 (N_6843,N_6704,N_6517);
xor U6844 (N_6844,N_6688,N_6699);
xor U6845 (N_6845,N_6672,N_6658);
nor U6846 (N_6846,N_6647,N_6512);
and U6847 (N_6847,N_6705,N_6661);
and U6848 (N_6848,N_6546,N_6542);
or U6849 (N_6849,N_6714,N_6571);
and U6850 (N_6850,N_6725,N_6635);
or U6851 (N_6851,N_6711,N_6738);
nor U6852 (N_6852,N_6500,N_6527);
xnor U6853 (N_6853,N_6626,N_6736);
and U6854 (N_6854,N_6607,N_6555);
nor U6855 (N_6855,N_6744,N_6554);
nor U6856 (N_6856,N_6540,N_6703);
or U6857 (N_6857,N_6640,N_6730);
or U6858 (N_6858,N_6589,N_6650);
and U6859 (N_6859,N_6598,N_6706);
nand U6860 (N_6860,N_6691,N_6664);
nand U6861 (N_6861,N_6739,N_6548);
and U6862 (N_6862,N_6695,N_6648);
xnor U6863 (N_6863,N_6696,N_6557);
and U6864 (N_6864,N_6505,N_6525);
nor U6865 (N_6865,N_6568,N_6509);
nor U6866 (N_6866,N_6513,N_6579);
and U6867 (N_6867,N_6538,N_6663);
nor U6868 (N_6868,N_6584,N_6559);
nor U6869 (N_6869,N_6575,N_6630);
and U6870 (N_6870,N_6622,N_6605);
nor U6871 (N_6871,N_6508,N_6603);
and U6872 (N_6872,N_6522,N_6620);
or U6873 (N_6873,N_6624,N_6655);
and U6874 (N_6874,N_6638,N_6668);
or U6875 (N_6875,N_6503,N_6734);
or U6876 (N_6876,N_6683,N_6735);
nor U6877 (N_6877,N_6656,N_6708);
nand U6878 (N_6878,N_6706,N_6735);
nand U6879 (N_6879,N_6731,N_6676);
and U6880 (N_6880,N_6539,N_6580);
nand U6881 (N_6881,N_6711,N_6531);
xor U6882 (N_6882,N_6559,N_6684);
nand U6883 (N_6883,N_6564,N_6585);
or U6884 (N_6884,N_6723,N_6542);
nand U6885 (N_6885,N_6671,N_6646);
xor U6886 (N_6886,N_6631,N_6581);
xnor U6887 (N_6887,N_6545,N_6567);
and U6888 (N_6888,N_6710,N_6706);
nand U6889 (N_6889,N_6660,N_6638);
and U6890 (N_6890,N_6576,N_6688);
nor U6891 (N_6891,N_6531,N_6690);
and U6892 (N_6892,N_6747,N_6531);
nand U6893 (N_6893,N_6690,N_6617);
nand U6894 (N_6894,N_6692,N_6641);
xor U6895 (N_6895,N_6666,N_6595);
nand U6896 (N_6896,N_6665,N_6505);
nand U6897 (N_6897,N_6504,N_6654);
or U6898 (N_6898,N_6728,N_6592);
or U6899 (N_6899,N_6542,N_6510);
xor U6900 (N_6900,N_6533,N_6690);
nor U6901 (N_6901,N_6748,N_6683);
and U6902 (N_6902,N_6688,N_6545);
and U6903 (N_6903,N_6632,N_6671);
nand U6904 (N_6904,N_6730,N_6661);
xnor U6905 (N_6905,N_6560,N_6664);
nor U6906 (N_6906,N_6696,N_6509);
or U6907 (N_6907,N_6563,N_6511);
and U6908 (N_6908,N_6662,N_6504);
or U6909 (N_6909,N_6504,N_6606);
and U6910 (N_6910,N_6697,N_6508);
nand U6911 (N_6911,N_6729,N_6652);
nor U6912 (N_6912,N_6627,N_6594);
nand U6913 (N_6913,N_6551,N_6669);
or U6914 (N_6914,N_6746,N_6549);
xnor U6915 (N_6915,N_6614,N_6565);
xor U6916 (N_6916,N_6633,N_6508);
or U6917 (N_6917,N_6607,N_6601);
or U6918 (N_6918,N_6728,N_6674);
and U6919 (N_6919,N_6600,N_6661);
xor U6920 (N_6920,N_6690,N_6661);
nand U6921 (N_6921,N_6601,N_6571);
xnor U6922 (N_6922,N_6550,N_6595);
xnor U6923 (N_6923,N_6715,N_6517);
nor U6924 (N_6924,N_6573,N_6696);
nand U6925 (N_6925,N_6692,N_6595);
nand U6926 (N_6926,N_6650,N_6643);
nor U6927 (N_6927,N_6654,N_6639);
xor U6928 (N_6928,N_6641,N_6590);
nand U6929 (N_6929,N_6577,N_6651);
nor U6930 (N_6930,N_6725,N_6713);
xor U6931 (N_6931,N_6524,N_6530);
nor U6932 (N_6932,N_6540,N_6697);
nand U6933 (N_6933,N_6590,N_6730);
or U6934 (N_6934,N_6605,N_6612);
nand U6935 (N_6935,N_6628,N_6716);
and U6936 (N_6936,N_6518,N_6733);
xnor U6937 (N_6937,N_6642,N_6677);
nor U6938 (N_6938,N_6696,N_6744);
nor U6939 (N_6939,N_6683,N_6556);
or U6940 (N_6940,N_6627,N_6695);
and U6941 (N_6941,N_6620,N_6716);
or U6942 (N_6942,N_6618,N_6633);
or U6943 (N_6943,N_6604,N_6552);
or U6944 (N_6944,N_6611,N_6605);
or U6945 (N_6945,N_6591,N_6633);
or U6946 (N_6946,N_6570,N_6721);
xnor U6947 (N_6947,N_6742,N_6546);
nand U6948 (N_6948,N_6631,N_6616);
or U6949 (N_6949,N_6683,N_6563);
and U6950 (N_6950,N_6732,N_6738);
or U6951 (N_6951,N_6605,N_6718);
xnor U6952 (N_6952,N_6583,N_6614);
nand U6953 (N_6953,N_6593,N_6621);
and U6954 (N_6954,N_6673,N_6622);
and U6955 (N_6955,N_6722,N_6532);
nor U6956 (N_6956,N_6643,N_6618);
xor U6957 (N_6957,N_6696,N_6680);
xor U6958 (N_6958,N_6540,N_6637);
xnor U6959 (N_6959,N_6693,N_6749);
xnor U6960 (N_6960,N_6576,N_6696);
xnor U6961 (N_6961,N_6557,N_6667);
and U6962 (N_6962,N_6659,N_6607);
xor U6963 (N_6963,N_6658,N_6712);
and U6964 (N_6964,N_6676,N_6574);
and U6965 (N_6965,N_6622,N_6737);
or U6966 (N_6966,N_6608,N_6536);
nor U6967 (N_6967,N_6637,N_6506);
and U6968 (N_6968,N_6628,N_6679);
xnor U6969 (N_6969,N_6706,N_6609);
and U6970 (N_6970,N_6587,N_6639);
xnor U6971 (N_6971,N_6577,N_6647);
or U6972 (N_6972,N_6642,N_6539);
or U6973 (N_6973,N_6630,N_6581);
or U6974 (N_6974,N_6633,N_6738);
and U6975 (N_6975,N_6727,N_6691);
and U6976 (N_6976,N_6628,N_6701);
nor U6977 (N_6977,N_6540,N_6660);
and U6978 (N_6978,N_6662,N_6510);
and U6979 (N_6979,N_6661,N_6587);
xor U6980 (N_6980,N_6747,N_6718);
nand U6981 (N_6981,N_6674,N_6574);
or U6982 (N_6982,N_6634,N_6596);
nor U6983 (N_6983,N_6591,N_6520);
xor U6984 (N_6984,N_6676,N_6623);
nand U6985 (N_6985,N_6590,N_6548);
nor U6986 (N_6986,N_6651,N_6552);
nor U6987 (N_6987,N_6688,N_6513);
or U6988 (N_6988,N_6704,N_6716);
or U6989 (N_6989,N_6576,N_6680);
and U6990 (N_6990,N_6592,N_6663);
xor U6991 (N_6991,N_6738,N_6534);
nor U6992 (N_6992,N_6649,N_6702);
and U6993 (N_6993,N_6577,N_6628);
or U6994 (N_6994,N_6711,N_6603);
xor U6995 (N_6995,N_6512,N_6595);
nand U6996 (N_6996,N_6602,N_6661);
nand U6997 (N_6997,N_6533,N_6735);
xor U6998 (N_6998,N_6695,N_6623);
nand U6999 (N_6999,N_6664,N_6598);
nor U7000 (N_7000,N_6938,N_6968);
nand U7001 (N_7001,N_6953,N_6802);
nor U7002 (N_7002,N_6793,N_6757);
nand U7003 (N_7003,N_6995,N_6919);
nand U7004 (N_7004,N_6814,N_6801);
and U7005 (N_7005,N_6976,N_6884);
nor U7006 (N_7006,N_6855,N_6779);
xor U7007 (N_7007,N_6877,N_6911);
nor U7008 (N_7008,N_6846,N_6851);
or U7009 (N_7009,N_6903,N_6901);
and U7010 (N_7010,N_6992,N_6822);
nor U7011 (N_7011,N_6896,N_6962);
nand U7012 (N_7012,N_6894,N_6811);
and U7013 (N_7013,N_6983,N_6831);
nor U7014 (N_7014,N_6778,N_6907);
or U7015 (N_7015,N_6763,N_6817);
xnor U7016 (N_7016,N_6967,N_6952);
nand U7017 (N_7017,N_6838,N_6806);
xnor U7018 (N_7018,N_6860,N_6957);
xor U7019 (N_7019,N_6932,N_6834);
and U7020 (N_7020,N_6808,N_6782);
xor U7021 (N_7021,N_6959,N_6942);
nor U7022 (N_7022,N_6833,N_6818);
nor U7023 (N_7023,N_6856,N_6853);
or U7024 (N_7024,N_6984,N_6956);
nor U7025 (N_7025,N_6985,N_6898);
or U7026 (N_7026,N_6905,N_6866);
and U7027 (N_7027,N_6914,N_6918);
and U7028 (N_7028,N_6832,N_6789);
nand U7029 (N_7029,N_6844,N_6913);
or U7030 (N_7030,N_6797,N_6847);
xor U7031 (N_7031,N_6977,N_6764);
xor U7032 (N_7032,N_6929,N_6785);
or U7033 (N_7033,N_6787,N_6840);
nand U7034 (N_7034,N_6777,N_6863);
or U7035 (N_7035,N_6839,N_6949);
or U7036 (N_7036,N_6972,N_6998);
nand U7037 (N_7037,N_6842,N_6836);
nor U7038 (N_7038,N_6876,N_6925);
or U7039 (N_7039,N_6788,N_6939);
nand U7040 (N_7040,N_6935,N_6902);
nand U7041 (N_7041,N_6857,N_6991);
nand U7042 (N_7042,N_6889,N_6899);
or U7043 (N_7043,N_6994,N_6852);
nand U7044 (N_7044,N_6859,N_6774);
nor U7045 (N_7045,N_6878,N_6762);
nand U7046 (N_7046,N_6837,N_6845);
and U7047 (N_7047,N_6882,N_6965);
nor U7048 (N_7048,N_6750,N_6820);
nor U7049 (N_7049,N_6821,N_6804);
xor U7050 (N_7050,N_6987,N_6854);
xnor U7051 (N_7051,N_6828,N_6997);
nand U7052 (N_7052,N_6941,N_6924);
or U7053 (N_7053,N_6955,N_6966);
nor U7054 (N_7054,N_6969,N_6880);
or U7055 (N_7055,N_6993,N_6819);
nand U7056 (N_7056,N_6861,N_6883);
nor U7057 (N_7057,N_6867,N_6803);
xnor U7058 (N_7058,N_6825,N_6843);
or U7059 (N_7059,N_6928,N_6761);
xor U7060 (N_7060,N_6879,N_6973);
nor U7061 (N_7061,N_6810,N_6970);
xor U7062 (N_7062,N_6865,N_6862);
xor U7063 (N_7063,N_6940,N_6873);
xnor U7064 (N_7064,N_6826,N_6963);
or U7065 (N_7065,N_6892,N_6950);
and U7066 (N_7066,N_6891,N_6781);
xnor U7067 (N_7067,N_6947,N_6786);
or U7068 (N_7068,N_6944,N_6943);
xor U7069 (N_7069,N_6835,N_6796);
and U7070 (N_7070,N_6981,N_6791);
and U7071 (N_7071,N_6794,N_6827);
nand U7072 (N_7072,N_6800,N_6980);
nand U7073 (N_7073,N_6986,N_6915);
xor U7074 (N_7074,N_6922,N_6875);
nand U7075 (N_7075,N_6760,N_6758);
or U7076 (N_7076,N_6869,N_6978);
nor U7077 (N_7077,N_6982,N_6799);
and U7078 (N_7078,N_6885,N_6769);
nor U7079 (N_7079,N_6868,N_6824);
xnor U7080 (N_7080,N_6999,N_6795);
nand U7081 (N_7081,N_6809,N_6767);
nor U7082 (N_7082,N_6816,N_6900);
and U7083 (N_7083,N_6921,N_6829);
or U7084 (N_7084,N_6979,N_6906);
nand U7085 (N_7085,N_6807,N_6945);
xnor U7086 (N_7086,N_6926,N_6961);
or U7087 (N_7087,N_6766,N_6784);
nor U7088 (N_7088,N_6916,N_6773);
or U7089 (N_7089,N_6920,N_6870);
xnor U7090 (N_7090,N_6752,N_6770);
nand U7091 (N_7091,N_6872,N_6908);
nor U7092 (N_7092,N_6815,N_6904);
nand U7093 (N_7093,N_6849,N_6813);
and U7094 (N_7094,N_6996,N_6772);
and U7095 (N_7095,N_6858,N_6792);
or U7096 (N_7096,N_6812,N_6895);
nor U7097 (N_7097,N_6912,N_6753);
xnor U7098 (N_7098,N_6848,N_6910);
xnor U7099 (N_7099,N_6805,N_6931);
nand U7100 (N_7100,N_6933,N_6964);
nand U7101 (N_7101,N_6755,N_6887);
nor U7102 (N_7102,N_6990,N_6881);
nor U7103 (N_7103,N_6909,N_6886);
or U7104 (N_7104,N_6989,N_6830);
or U7105 (N_7105,N_6850,N_6988);
or U7106 (N_7106,N_6798,N_6974);
nor U7107 (N_7107,N_6917,N_6754);
xnor U7108 (N_7108,N_6951,N_6971);
or U7109 (N_7109,N_6937,N_6768);
nand U7110 (N_7110,N_6888,N_6934);
and U7111 (N_7111,N_6871,N_6775);
nand U7112 (N_7112,N_6930,N_6841);
or U7113 (N_7113,N_6958,N_6893);
or U7114 (N_7114,N_6783,N_6936);
and U7115 (N_7115,N_6954,N_6897);
nand U7116 (N_7116,N_6864,N_6765);
xor U7117 (N_7117,N_6946,N_6927);
or U7118 (N_7118,N_6948,N_6874);
or U7119 (N_7119,N_6759,N_6890);
or U7120 (N_7120,N_6771,N_6751);
and U7121 (N_7121,N_6780,N_6960);
and U7122 (N_7122,N_6790,N_6823);
xor U7123 (N_7123,N_6776,N_6975);
nand U7124 (N_7124,N_6923,N_6756);
xor U7125 (N_7125,N_6781,N_6946);
nand U7126 (N_7126,N_6883,N_6918);
nand U7127 (N_7127,N_6949,N_6796);
nand U7128 (N_7128,N_6867,N_6881);
nand U7129 (N_7129,N_6935,N_6783);
xor U7130 (N_7130,N_6914,N_6795);
or U7131 (N_7131,N_6813,N_6907);
and U7132 (N_7132,N_6878,N_6892);
nor U7133 (N_7133,N_6976,N_6820);
xnor U7134 (N_7134,N_6920,N_6783);
xor U7135 (N_7135,N_6766,N_6918);
nor U7136 (N_7136,N_6843,N_6848);
or U7137 (N_7137,N_6764,N_6973);
or U7138 (N_7138,N_6828,N_6784);
nand U7139 (N_7139,N_6901,N_6855);
nand U7140 (N_7140,N_6844,N_6862);
nand U7141 (N_7141,N_6844,N_6956);
or U7142 (N_7142,N_6923,N_6796);
or U7143 (N_7143,N_6923,N_6978);
xor U7144 (N_7144,N_6839,N_6887);
nor U7145 (N_7145,N_6831,N_6885);
nor U7146 (N_7146,N_6780,N_6768);
and U7147 (N_7147,N_6811,N_6891);
nand U7148 (N_7148,N_6933,N_6776);
xor U7149 (N_7149,N_6841,N_6894);
xnor U7150 (N_7150,N_6840,N_6845);
nor U7151 (N_7151,N_6990,N_6843);
nor U7152 (N_7152,N_6819,N_6944);
and U7153 (N_7153,N_6976,N_6824);
and U7154 (N_7154,N_6916,N_6986);
nor U7155 (N_7155,N_6760,N_6854);
and U7156 (N_7156,N_6819,N_6862);
and U7157 (N_7157,N_6886,N_6821);
nand U7158 (N_7158,N_6914,N_6911);
nand U7159 (N_7159,N_6946,N_6963);
nand U7160 (N_7160,N_6837,N_6836);
or U7161 (N_7161,N_6969,N_6846);
xor U7162 (N_7162,N_6900,N_6984);
or U7163 (N_7163,N_6980,N_6781);
nand U7164 (N_7164,N_6848,N_6835);
nor U7165 (N_7165,N_6948,N_6904);
nand U7166 (N_7166,N_6999,N_6823);
nor U7167 (N_7167,N_6789,N_6750);
or U7168 (N_7168,N_6989,N_6906);
or U7169 (N_7169,N_6848,N_6924);
or U7170 (N_7170,N_6954,N_6982);
or U7171 (N_7171,N_6967,N_6860);
xor U7172 (N_7172,N_6973,N_6941);
or U7173 (N_7173,N_6968,N_6989);
nor U7174 (N_7174,N_6900,N_6848);
or U7175 (N_7175,N_6771,N_6776);
nor U7176 (N_7176,N_6807,N_6858);
xor U7177 (N_7177,N_6824,N_6784);
xor U7178 (N_7178,N_6801,N_6976);
nor U7179 (N_7179,N_6959,N_6766);
nor U7180 (N_7180,N_6772,N_6884);
nand U7181 (N_7181,N_6992,N_6906);
nand U7182 (N_7182,N_6867,N_6889);
and U7183 (N_7183,N_6869,N_6971);
and U7184 (N_7184,N_6839,N_6801);
xor U7185 (N_7185,N_6982,N_6791);
nor U7186 (N_7186,N_6992,N_6866);
and U7187 (N_7187,N_6821,N_6753);
or U7188 (N_7188,N_6870,N_6771);
nor U7189 (N_7189,N_6908,N_6763);
nor U7190 (N_7190,N_6769,N_6759);
and U7191 (N_7191,N_6907,N_6802);
nor U7192 (N_7192,N_6775,N_6911);
and U7193 (N_7193,N_6840,N_6782);
nand U7194 (N_7194,N_6914,N_6820);
nor U7195 (N_7195,N_6874,N_6923);
or U7196 (N_7196,N_6896,N_6796);
nor U7197 (N_7197,N_6755,N_6774);
nor U7198 (N_7198,N_6840,N_6940);
nor U7199 (N_7199,N_6865,N_6761);
and U7200 (N_7200,N_6751,N_6845);
nor U7201 (N_7201,N_6797,N_6827);
xnor U7202 (N_7202,N_6804,N_6861);
nand U7203 (N_7203,N_6796,N_6845);
and U7204 (N_7204,N_6867,N_6835);
xor U7205 (N_7205,N_6864,N_6971);
nand U7206 (N_7206,N_6858,N_6920);
nor U7207 (N_7207,N_6827,N_6921);
nand U7208 (N_7208,N_6965,N_6960);
xnor U7209 (N_7209,N_6973,N_6958);
xnor U7210 (N_7210,N_6962,N_6978);
or U7211 (N_7211,N_6890,N_6906);
xnor U7212 (N_7212,N_6759,N_6958);
xnor U7213 (N_7213,N_6863,N_6918);
or U7214 (N_7214,N_6959,N_6866);
nand U7215 (N_7215,N_6871,N_6948);
nor U7216 (N_7216,N_6978,N_6966);
nor U7217 (N_7217,N_6922,N_6896);
nand U7218 (N_7218,N_6810,N_6886);
nor U7219 (N_7219,N_6895,N_6940);
nand U7220 (N_7220,N_6892,N_6904);
or U7221 (N_7221,N_6830,N_6752);
and U7222 (N_7222,N_6895,N_6778);
xnor U7223 (N_7223,N_6989,N_6949);
and U7224 (N_7224,N_6898,N_6797);
or U7225 (N_7225,N_6787,N_6811);
nor U7226 (N_7226,N_6912,N_6989);
and U7227 (N_7227,N_6870,N_6906);
or U7228 (N_7228,N_6824,N_6787);
xnor U7229 (N_7229,N_6897,N_6763);
xnor U7230 (N_7230,N_6880,N_6994);
nand U7231 (N_7231,N_6782,N_6794);
and U7232 (N_7232,N_6769,N_6972);
and U7233 (N_7233,N_6992,N_6936);
nor U7234 (N_7234,N_6873,N_6920);
and U7235 (N_7235,N_6801,N_6955);
nor U7236 (N_7236,N_6903,N_6966);
and U7237 (N_7237,N_6809,N_6959);
or U7238 (N_7238,N_6809,N_6906);
nand U7239 (N_7239,N_6940,N_6770);
and U7240 (N_7240,N_6751,N_6852);
or U7241 (N_7241,N_6890,N_6856);
and U7242 (N_7242,N_6930,N_6762);
nand U7243 (N_7243,N_6860,N_6925);
xnor U7244 (N_7244,N_6789,N_6949);
and U7245 (N_7245,N_6777,N_6933);
or U7246 (N_7246,N_6963,N_6909);
and U7247 (N_7247,N_6788,N_6885);
and U7248 (N_7248,N_6786,N_6830);
nand U7249 (N_7249,N_6958,N_6880);
and U7250 (N_7250,N_7080,N_7088);
nand U7251 (N_7251,N_7190,N_7206);
nor U7252 (N_7252,N_7132,N_7180);
nor U7253 (N_7253,N_7071,N_7143);
or U7254 (N_7254,N_7053,N_7100);
nor U7255 (N_7255,N_7097,N_7136);
nor U7256 (N_7256,N_7072,N_7240);
xor U7257 (N_7257,N_7042,N_7197);
nand U7258 (N_7258,N_7068,N_7173);
xor U7259 (N_7259,N_7020,N_7022);
xnor U7260 (N_7260,N_7064,N_7189);
xnor U7261 (N_7261,N_7035,N_7224);
and U7262 (N_7262,N_7041,N_7203);
xnor U7263 (N_7263,N_7138,N_7044);
xnor U7264 (N_7264,N_7060,N_7109);
nor U7265 (N_7265,N_7156,N_7193);
or U7266 (N_7266,N_7168,N_7013);
and U7267 (N_7267,N_7162,N_7188);
and U7268 (N_7268,N_7147,N_7220);
or U7269 (N_7269,N_7200,N_7104);
nand U7270 (N_7270,N_7055,N_7078);
nor U7271 (N_7271,N_7122,N_7063);
or U7272 (N_7272,N_7117,N_7087);
nor U7273 (N_7273,N_7076,N_7187);
and U7274 (N_7274,N_7232,N_7134);
nor U7275 (N_7275,N_7141,N_7026);
or U7276 (N_7276,N_7149,N_7073);
and U7277 (N_7277,N_7107,N_7160);
xnor U7278 (N_7278,N_7079,N_7165);
and U7279 (N_7279,N_7059,N_7219);
and U7280 (N_7280,N_7050,N_7177);
xor U7281 (N_7281,N_7181,N_7030);
xor U7282 (N_7282,N_7084,N_7212);
or U7283 (N_7283,N_7011,N_7052);
nor U7284 (N_7284,N_7176,N_7093);
xor U7285 (N_7285,N_7008,N_7046);
nor U7286 (N_7286,N_7236,N_7032);
nand U7287 (N_7287,N_7056,N_7161);
nand U7288 (N_7288,N_7194,N_7112);
and U7289 (N_7289,N_7159,N_7094);
or U7290 (N_7290,N_7021,N_7144);
or U7291 (N_7291,N_7126,N_7028);
or U7292 (N_7292,N_7205,N_7127);
nor U7293 (N_7293,N_7047,N_7137);
or U7294 (N_7294,N_7214,N_7036);
or U7295 (N_7295,N_7183,N_7249);
and U7296 (N_7296,N_7024,N_7045);
xnor U7297 (N_7297,N_7043,N_7216);
or U7298 (N_7298,N_7081,N_7103);
nand U7299 (N_7299,N_7110,N_7179);
and U7300 (N_7300,N_7015,N_7199);
xnor U7301 (N_7301,N_7098,N_7146);
nor U7302 (N_7302,N_7034,N_7234);
or U7303 (N_7303,N_7211,N_7051);
nor U7304 (N_7304,N_7054,N_7151);
and U7305 (N_7305,N_7130,N_7226);
nor U7306 (N_7306,N_7196,N_7089);
and U7307 (N_7307,N_7012,N_7017);
nand U7308 (N_7308,N_7065,N_7208);
or U7309 (N_7309,N_7092,N_7006);
nor U7310 (N_7310,N_7185,N_7154);
and U7311 (N_7311,N_7119,N_7075);
nand U7312 (N_7312,N_7067,N_7218);
or U7313 (N_7313,N_7003,N_7010);
nor U7314 (N_7314,N_7111,N_7246);
and U7315 (N_7315,N_7031,N_7039);
nand U7316 (N_7316,N_7131,N_7082);
xnor U7317 (N_7317,N_7201,N_7191);
nor U7318 (N_7318,N_7228,N_7115);
nor U7319 (N_7319,N_7145,N_7086);
and U7320 (N_7320,N_7049,N_7106);
nor U7321 (N_7321,N_7023,N_7114);
xnor U7322 (N_7322,N_7155,N_7248);
nand U7323 (N_7323,N_7120,N_7038);
or U7324 (N_7324,N_7237,N_7231);
nor U7325 (N_7325,N_7192,N_7007);
nand U7326 (N_7326,N_7095,N_7005);
xnor U7327 (N_7327,N_7016,N_7004);
and U7328 (N_7328,N_7221,N_7217);
xnor U7329 (N_7329,N_7101,N_7166);
xor U7330 (N_7330,N_7062,N_7083);
and U7331 (N_7331,N_7215,N_7040);
xnor U7332 (N_7332,N_7230,N_7009);
nor U7333 (N_7333,N_7125,N_7202);
nor U7334 (N_7334,N_7163,N_7148);
xnor U7335 (N_7335,N_7241,N_7066);
and U7336 (N_7336,N_7002,N_7069);
nand U7337 (N_7337,N_7169,N_7121);
xor U7338 (N_7338,N_7245,N_7061);
and U7339 (N_7339,N_7129,N_7239);
and U7340 (N_7340,N_7142,N_7077);
or U7341 (N_7341,N_7198,N_7223);
xnor U7342 (N_7342,N_7242,N_7000);
nand U7343 (N_7343,N_7070,N_7157);
nand U7344 (N_7344,N_7027,N_7150);
nor U7345 (N_7345,N_7235,N_7184);
or U7346 (N_7346,N_7172,N_7133);
xor U7347 (N_7347,N_7118,N_7171);
or U7348 (N_7348,N_7116,N_7222);
nor U7349 (N_7349,N_7074,N_7029);
and U7350 (N_7350,N_7213,N_7113);
nand U7351 (N_7351,N_7014,N_7037);
and U7352 (N_7352,N_7128,N_7135);
xor U7353 (N_7353,N_7057,N_7167);
nor U7354 (N_7354,N_7090,N_7091);
or U7355 (N_7355,N_7227,N_7158);
nand U7356 (N_7356,N_7105,N_7225);
nor U7357 (N_7357,N_7140,N_7058);
xnor U7358 (N_7358,N_7033,N_7102);
xor U7359 (N_7359,N_7186,N_7244);
nand U7360 (N_7360,N_7108,N_7178);
nand U7361 (N_7361,N_7247,N_7229);
or U7362 (N_7362,N_7019,N_7182);
and U7363 (N_7363,N_7099,N_7025);
nand U7364 (N_7364,N_7139,N_7048);
and U7365 (N_7365,N_7238,N_7209);
nor U7366 (N_7366,N_7085,N_7170);
and U7367 (N_7367,N_7243,N_7207);
or U7368 (N_7368,N_7153,N_7175);
nor U7369 (N_7369,N_7124,N_7018);
or U7370 (N_7370,N_7001,N_7152);
xor U7371 (N_7371,N_7210,N_7233);
or U7372 (N_7372,N_7174,N_7164);
nand U7373 (N_7373,N_7096,N_7204);
nand U7374 (N_7374,N_7123,N_7195);
xnor U7375 (N_7375,N_7020,N_7171);
or U7376 (N_7376,N_7090,N_7182);
nor U7377 (N_7377,N_7143,N_7205);
and U7378 (N_7378,N_7132,N_7028);
or U7379 (N_7379,N_7188,N_7247);
or U7380 (N_7380,N_7097,N_7126);
nor U7381 (N_7381,N_7005,N_7045);
and U7382 (N_7382,N_7085,N_7067);
or U7383 (N_7383,N_7113,N_7027);
or U7384 (N_7384,N_7027,N_7235);
or U7385 (N_7385,N_7200,N_7049);
nand U7386 (N_7386,N_7051,N_7077);
or U7387 (N_7387,N_7180,N_7100);
xnor U7388 (N_7388,N_7128,N_7106);
nand U7389 (N_7389,N_7073,N_7229);
nand U7390 (N_7390,N_7008,N_7074);
or U7391 (N_7391,N_7205,N_7165);
nor U7392 (N_7392,N_7172,N_7001);
nor U7393 (N_7393,N_7146,N_7232);
nor U7394 (N_7394,N_7052,N_7217);
nand U7395 (N_7395,N_7244,N_7126);
or U7396 (N_7396,N_7051,N_7196);
nand U7397 (N_7397,N_7029,N_7046);
nor U7398 (N_7398,N_7219,N_7091);
nand U7399 (N_7399,N_7012,N_7189);
nor U7400 (N_7400,N_7087,N_7017);
xnor U7401 (N_7401,N_7183,N_7170);
or U7402 (N_7402,N_7153,N_7164);
or U7403 (N_7403,N_7173,N_7009);
nor U7404 (N_7404,N_7043,N_7018);
nor U7405 (N_7405,N_7121,N_7097);
xnor U7406 (N_7406,N_7056,N_7163);
or U7407 (N_7407,N_7245,N_7194);
and U7408 (N_7408,N_7070,N_7190);
nor U7409 (N_7409,N_7162,N_7042);
and U7410 (N_7410,N_7110,N_7081);
xor U7411 (N_7411,N_7045,N_7068);
nor U7412 (N_7412,N_7192,N_7146);
or U7413 (N_7413,N_7143,N_7082);
nand U7414 (N_7414,N_7242,N_7126);
or U7415 (N_7415,N_7049,N_7096);
nand U7416 (N_7416,N_7175,N_7009);
and U7417 (N_7417,N_7106,N_7069);
nor U7418 (N_7418,N_7038,N_7050);
xor U7419 (N_7419,N_7214,N_7092);
or U7420 (N_7420,N_7237,N_7025);
or U7421 (N_7421,N_7223,N_7030);
and U7422 (N_7422,N_7230,N_7202);
xor U7423 (N_7423,N_7054,N_7062);
or U7424 (N_7424,N_7098,N_7228);
xnor U7425 (N_7425,N_7187,N_7050);
nor U7426 (N_7426,N_7170,N_7199);
xor U7427 (N_7427,N_7227,N_7095);
nand U7428 (N_7428,N_7054,N_7072);
xnor U7429 (N_7429,N_7028,N_7096);
nor U7430 (N_7430,N_7011,N_7085);
and U7431 (N_7431,N_7100,N_7179);
nor U7432 (N_7432,N_7118,N_7170);
nor U7433 (N_7433,N_7091,N_7048);
and U7434 (N_7434,N_7134,N_7118);
xnor U7435 (N_7435,N_7174,N_7030);
or U7436 (N_7436,N_7136,N_7167);
and U7437 (N_7437,N_7121,N_7094);
nand U7438 (N_7438,N_7241,N_7007);
nand U7439 (N_7439,N_7086,N_7193);
and U7440 (N_7440,N_7114,N_7174);
xor U7441 (N_7441,N_7125,N_7050);
or U7442 (N_7442,N_7226,N_7194);
and U7443 (N_7443,N_7129,N_7249);
xor U7444 (N_7444,N_7081,N_7093);
or U7445 (N_7445,N_7090,N_7106);
or U7446 (N_7446,N_7174,N_7170);
nor U7447 (N_7447,N_7084,N_7161);
and U7448 (N_7448,N_7018,N_7058);
nand U7449 (N_7449,N_7004,N_7120);
or U7450 (N_7450,N_7163,N_7236);
nand U7451 (N_7451,N_7001,N_7202);
nor U7452 (N_7452,N_7217,N_7060);
and U7453 (N_7453,N_7086,N_7236);
and U7454 (N_7454,N_7213,N_7172);
or U7455 (N_7455,N_7138,N_7247);
xor U7456 (N_7456,N_7003,N_7236);
or U7457 (N_7457,N_7118,N_7023);
xnor U7458 (N_7458,N_7135,N_7140);
or U7459 (N_7459,N_7239,N_7035);
xor U7460 (N_7460,N_7222,N_7207);
or U7461 (N_7461,N_7219,N_7117);
nand U7462 (N_7462,N_7186,N_7151);
xor U7463 (N_7463,N_7138,N_7246);
nand U7464 (N_7464,N_7063,N_7108);
nor U7465 (N_7465,N_7120,N_7231);
or U7466 (N_7466,N_7195,N_7209);
nand U7467 (N_7467,N_7090,N_7238);
nand U7468 (N_7468,N_7185,N_7039);
or U7469 (N_7469,N_7163,N_7000);
nor U7470 (N_7470,N_7243,N_7162);
xor U7471 (N_7471,N_7225,N_7062);
nand U7472 (N_7472,N_7098,N_7112);
and U7473 (N_7473,N_7069,N_7056);
xor U7474 (N_7474,N_7237,N_7083);
xnor U7475 (N_7475,N_7217,N_7190);
and U7476 (N_7476,N_7100,N_7064);
and U7477 (N_7477,N_7235,N_7248);
nor U7478 (N_7478,N_7181,N_7101);
nand U7479 (N_7479,N_7130,N_7063);
and U7480 (N_7480,N_7078,N_7147);
or U7481 (N_7481,N_7099,N_7158);
nor U7482 (N_7482,N_7172,N_7026);
or U7483 (N_7483,N_7078,N_7059);
and U7484 (N_7484,N_7006,N_7131);
or U7485 (N_7485,N_7230,N_7019);
nand U7486 (N_7486,N_7149,N_7061);
nor U7487 (N_7487,N_7042,N_7026);
and U7488 (N_7488,N_7077,N_7248);
xnor U7489 (N_7489,N_7147,N_7131);
and U7490 (N_7490,N_7152,N_7165);
and U7491 (N_7491,N_7130,N_7083);
nand U7492 (N_7492,N_7023,N_7241);
nor U7493 (N_7493,N_7104,N_7117);
nand U7494 (N_7494,N_7141,N_7107);
nand U7495 (N_7495,N_7034,N_7202);
nand U7496 (N_7496,N_7040,N_7229);
xor U7497 (N_7497,N_7189,N_7013);
nor U7498 (N_7498,N_7091,N_7212);
and U7499 (N_7499,N_7159,N_7178);
or U7500 (N_7500,N_7335,N_7478);
nand U7501 (N_7501,N_7289,N_7447);
and U7502 (N_7502,N_7389,N_7407);
xor U7503 (N_7503,N_7326,N_7384);
or U7504 (N_7504,N_7424,N_7324);
and U7505 (N_7505,N_7339,N_7340);
and U7506 (N_7506,N_7349,N_7329);
or U7507 (N_7507,N_7322,N_7325);
nor U7508 (N_7508,N_7401,N_7367);
or U7509 (N_7509,N_7438,N_7465);
and U7510 (N_7510,N_7254,N_7468);
or U7511 (N_7511,N_7261,N_7319);
or U7512 (N_7512,N_7290,N_7444);
or U7513 (N_7513,N_7453,N_7347);
or U7514 (N_7514,N_7355,N_7291);
nand U7515 (N_7515,N_7459,N_7286);
nand U7516 (N_7516,N_7393,N_7271);
or U7517 (N_7517,N_7442,N_7299);
nor U7518 (N_7518,N_7433,N_7492);
or U7519 (N_7519,N_7440,N_7486);
nor U7520 (N_7520,N_7262,N_7451);
nand U7521 (N_7521,N_7489,N_7275);
nor U7522 (N_7522,N_7422,N_7314);
or U7523 (N_7523,N_7348,N_7304);
and U7524 (N_7524,N_7467,N_7400);
and U7525 (N_7525,N_7449,N_7318);
and U7526 (N_7526,N_7456,N_7398);
and U7527 (N_7527,N_7315,N_7491);
nand U7528 (N_7528,N_7352,N_7374);
xor U7529 (N_7529,N_7338,N_7321);
or U7530 (N_7530,N_7327,N_7266);
nand U7531 (N_7531,N_7448,N_7446);
or U7532 (N_7532,N_7375,N_7431);
xnor U7533 (N_7533,N_7333,N_7488);
nand U7534 (N_7534,N_7414,N_7403);
nand U7535 (N_7535,N_7471,N_7436);
nor U7536 (N_7536,N_7421,N_7293);
and U7537 (N_7537,N_7463,N_7455);
xnor U7538 (N_7538,N_7300,N_7425);
nand U7539 (N_7539,N_7399,N_7493);
nand U7540 (N_7540,N_7415,N_7269);
nand U7541 (N_7541,N_7281,N_7420);
xor U7542 (N_7542,N_7409,N_7294);
nand U7543 (N_7543,N_7474,N_7377);
nor U7544 (N_7544,N_7426,N_7292);
or U7545 (N_7545,N_7280,N_7371);
nand U7546 (N_7546,N_7270,N_7361);
xor U7547 (N_7547,N_7383,N_7481);
or U7548 (N_7548,N_7341,N_7419);
and U7549 (N_7549,N_7317,N_7250);
nand U7550 (N_7550,N_7285,N_7255);
nor U7551 (N_7551,N_7394,N_7387);
or U7552 (N_7552,N_7330,N_7258);
nand U7553 (N_7553,N_7365,N_7282);
or U7554 (N_7554,N_7476,N_7469);
xor U7555 (N_7555,N_7303,N_7411);
nor U7556 (N_7556,N_7482,N_7429);
xor U7557 (N_7557,N_7434,N_7410);
xnor U7558 (N_7558,N_7360,N_7391);
or U7559 (N_7559,N_7395,N_7356);
nand U7560 (N_7560,N_7274,N_7379);
or U7561 (N_7561,N_7350,N_7336);
and U7562 (N_7562,N_7323,N_7268);
nor U7563 (N_7563,N_7364,N_7278);
or U7564 (N_7564,N_7477,N_7288);
xnor U7565 (N_7565,N_7480,N_7316);
nor U7566 (N_7566,N_7260,N_7272);
or U7567 (N_7567,N_7345,N_7344);
nor U7568 (N_7568,N_7351,N_7450);
nor U7569 (N_7569,N_7382,N_7405);
nor U7570 (N_7570,N_7334,N_7435);
or U7571 (N_7571,N_7416,N_7257);
and U7572 (N_7572,N_7494,N_7466);
xor U7573 (N_7573,N_7284,N_7483);
nor U7574 (N_7574,N_7497,N_7259);
nor U7575 (N_7575,N_7283,N_7311);
nand U7576 (N_7576,N_7308,N_7253);
and U7577 (N_7577,N_7445,N_7484);
nor U7578 (N_7578,N_7328,N_7462);
xnor U7579 (N_7579,N_7392,N_7404);
xor U7580 (N_7580,N_7287,N_7313);
nand U7581 (N_7581,N_7475,N_7373);
and U7582 (N_7582,N_7252,N_7297);
xnor U7583 (N_7583,N_7363,N_7331);
nand U7584 (N_7584,N_7457,N_7470);
nor U7585 (N_7585,N_7385,N_7452);
or U7586 (N_7586,N_7485,N_7498);
nor U7587 (N_7587,N_7376,N_7490);
and U7588 (N_7588,N_7427,N_7310);
and U7589 (N_7589,N_7305,N_7265);
nand U7590 (N_7590,N_7309,N_7413);
nand U7591 (N_7591,N_7332,N_7402);
or U7592 (N_7592,N_7378,N_7251);
nor U7593 (N_7593,N_7381,N_7472);
nand U7594 (N_7594,N_7337,N_7437);
and U7595 (N_7595,N_7366,N_7354);
nand U7596 (N_7596,N_7487,N_7296);
and U7597 (N_7597,N_7256,N_7353);
nand U7598 (N_7598,N_7390,N_7273);
xor U7599 (N_7599,N_7495,N_7359);
xor U7600 (N_7600,N_7423,N_7368);
xnor U7601 (N_7601,N_7479,N_7432);
nor U7602 (N_7602,N_7454,N_7277);
nor U7603 (N_7603,N_7408,N_7388);
nand U7604 (N_7604,N_7380,N_7267);
and U7605 (N_7605,N_7386,N_7441);
xnor U7606 (N_7606,N_7342,N_7362);
or U7607 (N_7607,N_7396,N_7295);
xnor U7608 (N_7608,N_7430,N_7496);
or U7609 (N_7609,N_7264,N_7460);
nand U7610 (N_7610,N_7406,N_7279);
nor U7611 (N_7611,N_7397,N_7443);
xnor U7612 (N_7612,N_7370,N_7263);
xnor U7613 (N_7613,N_7346,N_7464);
and U7614 (N_7614,N_7307,N_7320);
or U7615 (N_7615,N_7369,N_7301);
or U7616 (N_7616,N_7343,N_7312);
nor U7617 (N_7617,N_7473,N_7358);
nor U7618 (N_7618,N_7276,N_7439);
nand U7619 (N_7619,N_7306,N_7372);
xnor U7620 (N_7620,N_7428,N_7499);
and U7621 (N_7621,N_7302,N_7461);
or U7622 (N_7622,N_7417,N_7412);
nor U7623 (N_7623,N_7298,N_7357);
xor U7624 (N_7624,N_7458,N_7418);
or U7625 (N_7625,N_7390,N_7494);
and U7626 (N_7626,N_7385,N_7394);
and U7627 (N_7627,N_7321,N_7350);
nor U7628 (N_7628,N_7297,N_7341);
or U7629 (N_7629,N_7428,N_7419);
nor U7630 (N_7630,N_7451,N_7485);
or U7631 (N_7631,N_7398,N_7462);
xor U7632 (N_7632,N_7274,N_7344);
xnor U7633 (N_7633,N_7373,N_7296);
xor U7634 (N_7634,N_7418,N_7439);
nor U7635 (N_7635,N_7478,N_7407);
nand U7636 (N_7636,N_7468,N_7312);
and U7637 (N_7637,N_7411,N_7466);
xnor U7638 (N_7638,N_7337,N_7405);
xnor U7639 (N_7639,N_7305,N_7424);
nand U7640 (N_7640,N_7466,N_7479);
nor U7641 (N_7641,N_7440,N_7464);
and U7642 (N_7642,N_7429,N_7468);
nor U7643 (N_7643,N_7438,N_7480);
xor U7644 (N_7644,N_7400,N_7470);
nor U7645 (N_7645,N_7470,N_7311);
and U7646 (N_7646,N_7252,N_7349);
nor U7647 (N_7647,N_7406,N_7408);
xnor U7648 (N_7648,N_7384,N_7453);
or U7649 (N_7649,N_7448,N_7343);
xnor U7650 (N_7650,N_7273,N_7481);
and U7651 (N_7651,N_7323,N_7272);
xor U7652 (N_7652,N_7343,N_7394);
and U7653 (N_7653,N_7485,N_7406);
or U7654 (N_7654,N_7388,N_7477);
nand U7655 (N_7655,N_7287,N_7393);
nor U7656 (N_7656,N_7404,N_7299);
nand U7657 (N_7657,N_7254,N_7346);
nand U7658 (N_7658,N_7488,N_7435);
xnor U7659 (N_7659,N_7372,N_7322);
or U7660 (N_7660,N_7343,N_7254);
xnor U7661 (N_7661,N_7303,N_7429);
or U7662 (N_7662,N_7275,N_7464);
or U7663 (N_7663,N_7326,N_7411);
nand U7664 (N_7664,N_7365,N_7490);
nor U7665 (N_7665,N_7327,N_7457);
and U7666 (N_7666,N_7389,N_7457);
and U7667 (N_7667,N_7257,N_7330);
nor U7668 (N_7668,N_7397,N_7367);
xnor U7669 (N_7669,N_7348,N_7339);
or U7670 (N_7670,N_7292,N_7440);
nand U7671 (N_7671,N_7435,N_7459);
and U7672 (N_7672,N_7321,N_7348);
or U7673 (N_7673,N_7345,N_7319);
xnor U7674 (N_7674,N_7337,N_7408);
xnor U7675 (N_7675,N_7413,N_7362);
xnor U7676 (N_7676,N_7387,N_7415);
and U7677 (N_7677,N_7430,N_7302);
or U7678 (N_7678,N_7257,N_7289);
nor U7679 (N_7679,N_7444,N_7445);
nor U7680 (N_7680,N_7418,N_7284);
nor U7681 (N_7681,N_7406,N_7282);
xor U7682 (N_7682,N_7310,N_7400);
or U7683 (N_7683,N_7457,N_7418);
nand U7684 (N_7684,N_7279,N_7276);
or U7685 (N_7685,N_7437,N_7466);
and U7686 (N_7686,N_7492,N_7498);
and U7687 (N_7687,N_7386,N_7336);
and U7688 (N_7688,N_7323,N_7346);
nand U7689 (N_7689,N_7467,N_7341);
nand U7690 (N_7690,N_7388,N_7456);
or U7691 (N_7691,N_7319,N_7326);
and U7692 (N_7692,N_7258,N_7254);
nand U7693 (N_7693,N_7287,N_7423);
and U7694 (N_7694,N_7350,N_7462);
nand U7695 (N_7695,N_7461,N_7267);
xnor U7696 (N_7696,N_7338,N_7272);
xnor U7697 (N_7697,N_7450,N_7312);
nand U7698 (N_7698,N_7447,N_7480);
and U7699 (N_7699,N_7325,N_7345);
or U7700 (N_7700,N_7463,N_7449);
nor U7701 (N_7701,N_7483,N_7367);
nand U7702 (N_7702,N_7482,N_7434);
or U7703 (N_7703,N_7273,N_7402);
and U7704 (N_7704,N_7392,N_7441);
or U7705 (N_7705,N_7298,N_7375);
nor U7706 (N_7706,N_7443,N_7476);
nor U7707 (N_7707,N_7462,N_7432);
nand U7708 (N_7708,N_7356,N_7455);
xnor U7709 (N_7709,N_7330,N_7431);
or U7710 (N_7710,N_7402,N_7456);
xnor U7711 (N_7711,N_7388,N_7451);
and U7712 (N_7712,N_7321,N_7364);
xor U7713 (N_7713,N_7444,N_7491);
and U7714 (N_7714,N_7277,N_7353);
xor U7715 (N_7715,N_7309,N_7324);
nor U7716 (N_7716,N_7492,N_7360);
xnor U7717 (N_7717,N_7365,N_7339);
or U7718 (N_7718,N_7360,N_7280);
nor U7719 (N_7719,N_7341,N_7455);
or U7720 (N_7720,N_7363,N_7372);
nand U7721 (N_7721,N_7387,N_7407);
nor U7722 (N_7722,N_7335,N_7367);
nor U7723 (N_7723,N_7260,N_7493);
nand U7724 (N_7724,N_7276,N_7360);
xnor U7725 (N_7725,N_7259,N_7356);
or U7726 (N_7726,N_7444,N_7373);
or U7727 (N_7727,N_7462,N_7472);
nor U7728 (N_7728,N_7391,N_7405);
nor U7729 (N_7729,N_7383,N_7299);
nor U7730 (N_7730,N_7396,N_7485);
or U7731 (N_7731,N_7336,N_7293);
xnor U7732 (N_7732,N_7294,N_7464);
xor U7733 (N_7733,N_7298,N_7464);
or U7734 (N_7734,N_7273,N_7290);
and U7735 (N_7735,N_7460,N_7485);
nor U7736 (N_7736,N_7467,N_7332);
or U7737 (N_7737,N_7331,N_7254);
nor U7738 (N_7738,N_7425,N_7372);
and U7739 (N_7739,N_7462,N_7260);
xnor U7740 (N_7740,N_7315,N_7269);
nor U7741 (N_7741,N_7452,N_7352);
xor U7742 (N_7742,N_7420,N_7469);
nand U7743 (N_7743,N_7472,N_7385);
or U7744 (N_7744,N_7495,N_7342);
nor U7745 (N_7745,N_7317,N_7285);
nor U7746 (N_7746,N_7426,N_7396);
xor U7747 (N_7747,N_7256,N_7453);
xnor U7748 (N_7748,N_7423,N_7450);
and U7749 (N_7749,N_7384,N_7461);
and U7750 (N_7750,N_7670,N_7611);
or U7751 (N_7751,N_7626,N_7582);
xnor U7752 (N_7752,N_7716,N_7725);
nor U7753 (N_7753,N_7657,N_7647);
nand U7754 (N_7754,N_7588,N_7649);
nand U7755 (N_7755,N_7513,N_7684);
or U7756 (N_7756,N_7604,N_7742);
nor U7757 (N_7757,N_7656,N_7636);
and U7758 (N_7758,N_7594,N_7708);
and U7759 (N_7759,N_7517,N_7702);
xnor U7760 (N_7760,N_7525,N_7516);
nand U7761 (N_7761,N_7538,N_7722);
nor U7762 (N_7762,N_7614,N_7562);
nor U7763 (N_7763,N_7704,N_7741);
or U7764 (N_7764,N_7613,N_7584);
nand U7765 (N_7765,N_7527,N_7712);
and U7766 (N_7766,N_7601,N_7624);
and U7767 (N_7767,N_7532,N_7509);
or U7768 (N_7768,N_7526,N_7537);
or U7769 (N_7769,N_7633,N_7746);
and U7770 (N_7770,N_7747,N_7618);
nand U7771 (N_7771,N_7703,N_7678);
nand U7772 (N_7772,N_7677,N_7603);
nand U7773 (N_7773,N_7502,N_7609);
and U7774 (N_7774,N_7713,N_7570);
or U7775 (N_7775,N_7616,N_7694);
or U7776 (N_7776,N_7720,N_7607);
and U7777 (N_7777,N_7659,N_7697);
or U7778 (N_7778,N_7736,N_7683);
nand U7779 (N_7779,N_7507,N_7638);
nand U7780 (N_7780,N_7520,N_7530);
nor U7781 (N_7781,N_7714,N_7691);
xor U7782 (N_7782,N_7685,N_7731);
xor U7783 (N_7783,N_7709,N_7695);
and U7784 (N_7784,N_7675,N_7682);
nand U7785 (N_7785,N_7654,N_7748);
nor U7786 (N_7786,N_7580,N_7625);
nor U7787 (N_7787,N_7514,N_7730);
xor U7788 (N_7788,N_7553,N_7566);
nand U7789 (N_7789,N_7653,N_7558);
or U7790 (N_7790,N_7599,N_7700);
nor U7791 (N_7791,N_7512,N_7669);
xor U7792 (N_7792,N_7658,N_7710);
and U7793 (N_7793,N_7726,N_7504);
nor U7794 (N_7794,N_7533,N_7590);
nor U7795 (N_7795,N_7667,N_7688);
xor U7796 (N_7796,N_7606,N_7506);
nand U7797 (N_7797,N_7587,N_7648);
or U7798 (N_7798,N_7620,N_7738);
nor U7799 (N_7799,N_7508,N_7642);
nor U7800 (N_7800,N_7529,N_7552);
nor U7801 (N_7801,N_7510,N_7701);
and U7802 (N_7802,N_7575,N_7727);
xor U7803 (N_7803,N_7643,N_7621);
xnor U7804 (N_7804,N_7598,N_7576);
or U7805 (N_7805,N_7548,N_7541);
xnor U7806 (N_7806,N_7545,N_7577);
nor U7807 (N_7807,N_7744,N_7534);
or U7808 (N_7808,N_7503,N_7637);
or U7809 (N_7809,N_7559,N_7585);
xor U7810 (N_7810,N_7557,N_7554);
and U7811 (N_7811,N_7630,N_7500);
or U7812 (N_7812,N_7539,N_7573);
nor U7813 (N_7813,N_7672,N_7628);
and U7814 (N_7814,N_7662,N_7743);
xnor U7815 (N_7815,N_7634,N_7693);
xor U7816 (N_7816,N_7724,N_7673);
or U7817 (N_7817,N_7592,N_7623);
xnor U7818 (N_7818,N_7661,N_7615);
nor U7819 (N_7819,N_7597,N_7668);
xnor U7820 (N_7820,N_7536,N_7687);
nand U7821 (N_7821,N_7589,N_7728);
and U7822 (N_7822,N_7698,N_7681);
or U7823 (N_7823,N_7549,N_7602);
nor U7824 (N_7824,N_7629,N_7522);
and U7825 (N_7825,N_7567,N_7515);
nor U7826 (N_7826,N_7671,N_7505);
and U7827 (N_7827,N_7627,N_7739);
and U7828 (N_7828,N_7610,N_7640);
xor U7829 (N_7829,N_7561,N_7535);
nand U7830 (N_7830,N_7655,N_7521);
nor U7831 (N_7831,N_7528,N_7718);
xnor U7832 (N_7832,N_7531,N_7680);
and U7833 (N_7833,N_7569,N_7674);
xor U7834 (N_7834,N_7737,N_7711);
nand U7835 (N_7835,N_7581,N_7565);
or U7836 (N_7836,N_7556,N_7519);
and U7837 (N_7837,N_7735,N_7689);
and U7838 (N_7838,N_7555,N_7740);
or U7839 (N_7839,N_7563,N_7664);
or U7840 (N_7840,N_7717,N_7600);
or U7841 (N_7841,N_7733,N_7651);
or U7842 (N_7842,N_7608,N_7696);
and U7843 (N_7843,N_7571,N_7666);
or U7844 (N_7844,N_7622,N_7749);
nand U7845 (N_7845,N_7560,N_7501);
nand U7846 (N_7846,N_7734,N_7542);
or U7847 (N_7847,N_7635,N_7690);
xor U7848 (N_7848,N_7572,N_7705);
xnor U7849 (N_7849,N_7676,N_7650);
xnor U7850 (N_7850,N_7605,N_7692);
or U7851 (N_7851,N_7518,N_7596);
nand U7852 (N_7852,N_7551,N_7564);
or U7853 (N_7853,N_7699,N_7745);
nor U7854 (N_7854,N_7686,N_7644);
and U7855 (N_7855,N_7639,N_7574);
nand U7856 (N_7856,N_7715,N_7591);
and U7857 (N_7857,N_7547,N_7619);
nor U7858 (N_7858,N_7568,N_7550);
and U7859 (N_7859,N_7524,N_7612);
nand U7860 (N_7860,N_7645,N_7583);
nand U7861 (N_7861,N_7729,N_7578);
or U7862 (N_7862,N_7540,N_7707);
and U7863 (N_7863,N_7721,N_7732);
nor U7864 (N_7864,N_7652,N_7586);
or U7865 (N_7865,N_7679,N_7723);
xnor U7866 (N_7866,N_7719,N_7632);
or U7867 (N_7867,N_7523,N_7663);
and U7868 (N_7868,N_7546,N_7579);
nand U7869 (N_7869,N_7511,N_7595);
or U7870 (N_7870,N_7660,N_7641);
xnor U7871 (N_7871,N_7631,N_7593);
and U7872 (N_7872,N_7646,N_7706);
and U7873 (N_7873,N_7665,N_7617);
nand U7874 (N_7874,N_7543,N_7544);
nand U7875 (N_7875,N_7642,N_7729);
and U7876 (N_7876,N_7572,N_7724);
and U7877 (N_7877,N_7672,N_7588);
xnor U7878 (N_7878,N_7584,N_7506);
or U7879 (N_7879,N_7607,N_7671);
or U7880 (N_7880,N_7735,N_7716);
nor U7881 (N_7881,N_7553,N_7695);
and U7882 (N_7882,N_7525,N_7679);
xnor U7883 (N_7883,N_7663,N_7650);
and U7884 (N_7884,N_7583,N_7604);
xor U7885 (N_7885,N_7732,N_7690);
xor U7886 (N_7886,N_7628,N_7725);
nor U7887 (N_7887,N_7502,N_7633);
nor U7888 (N_7888,N_7598,N_7560);
nor U7889 (N_7889,N_7600,N_7629);
and U7890 (N_7890,N_7529,N_7647);
xor U7891 (N_7891,N_7506,N_7691);
or U7892 (N_7892,N_7574,N_7692);
or U7893 (N_7893,N_7639,N_7648);
and U7894 (N_7894,N_7569,N_7670);
nand U7895 (N_7895,N_7544,N_7527);
nand U7896 (N_7896,N_7551,N_7623);
nand U7897 (N_7897,N_7539,N_7564);
xor U7898 (N_7898,N_7700,N_7691);
or U7899 (N_7899,N_7645,N_7553);
and U7900 (N_7900,N_7589,N_7574);
nor U7901 (N_7901,N_7641,N_7649);
nand U7902 (N_7902,N_7744,N_7509);
nand U7903 (N_7903,N_7521,N_7661);
nand U7904 (N_7904,N_7679,N_7686);
nand U7905 (N_7905,N_7682,N_7655);
nor U7906 (N_7906,N_7671,N_7557);
and U7907 (N_7907,N_7566,N_7514);
xor U7908 (N_7908,N_7533,N_7718);
and U7909 (N_7909,N_7555,N_7643);
nand U7910 (N_7910,N_7734,N_7717);
or U7911 (N_7911,N_7546,N_7501);
xnor U7912 (N_7912,N_7633,N_7516);
and U7913 (N_7913,N_7638,N_7522);
or U7914 (N_7914,N_7622,N_7560);
nor U7915 (N_7915,N_7680,N_7597);
and U7916 (N_7916,N_7688,N_7744);
nand U7917 (N_7917,N_7661,N_7563);
nand U7918 (N_7918,N_7532,N_7667);
or U7919 (N_7919,N_7720,N_7732);
nor U7920 (N_7920,N_7689,N_7557);
xor U7921 (N_7921,N_7732,N_7653);
or U7922 (N_7922,N_7577,N_7626);
or U7923 (N_7923,N_7731,N_7575);
xor U7924 (N_7924,N_7688,N_7531);
and U7925 (N_7925,N_7729,N_7611);
xor U7926 (N_7926,N_7582,N_7552);
nor U7927 (N_7927,N_7562,N_7523);
xor U7928 (N_7928,N_7662,N_7747);
xnor U7929 (N_7929,N_7712,N_7599);
and U7930 (N_7930,N_7683,N_7570);
xnor U7931 (N_7931,N_7511,N_7691);
nand U7932 (N_7932,N_7598,N_7566);
nand U7933 (N_7933,N_7653,N_7623);
nor U7934 (N_7934,N_7642,N_7638);
nand U7935 (N_7935,N_7528,N_7601);
and U7936 (N_7936,N_7593,N_7620);
nor U7937 (N_7937,N_7704,N_7622);
xnor U7938 (N_7938,N_7707,N_7580);
nor U7939 (N_7939,N_7677,N_7531);
and U7940 (N_7940,N_7601,N_7745);
nor U7941 (N_7941,N_7680,N_7543);
nor U7942 (N_7942,N_7539,N_7594);
nand U7943 (N_7943,N_7707,N_7658);
and U7944 (N_7944,N_7592,N_7631);
nor U7945 (N_7945,N_7571,N_7658);
or U7946 (N_7946,N_7700,N_7502);
or U7947 (N_7947,N_7636,N_7539);
and U7948 (N_7948,N_7671,N_7586);
and U7949 (N_7949,N_7744,N_7524);
or U7950 (N_7950,N_7575,N_7701);
nand U7951 (N_7951,N_7703,N_7705);
or U7952 (N_7952,N_7569,N_7693);
and U7953 (N_7953,N_7545,N_7622);
or U7954 (N_7954,N_7703,N_7553);
nor U7955 (N_7955,N_7528,N_7515);
nand U7956 (N_7956,N_7604,N_7703);
and U7957 (N_7957,N_7738,N_7713);
or U7958 (N_7958,N_7584,N_7683);
nand U7959 (N_7959,N_7644,N_7703);
xor U7960 (N_7960,N_7713,N_7587);
nand U7961 (N_7961,N_7603,N_7715);
nand U7962 (N_7962,N_7665,N_7698);
nand U7963 (N_7963,N_7531,N_7721);
xor U7964 (N_7964,N_7725,N_7560);
and U7965 (N_7965,N_7518,N_7603);
nand U7966 (N_7966,N_7539,N_7714);
xor U7967 (N_7967,N_7578,N_7746);
or U7968 (N_7968,N_7684,N_7569);
or U7969 (N_7969,N_7738,N_7640);
xor U7970 (N_7970,N_7549,N_7510);
or U7971 (N_7971,N_7551,N_7535);
nor U7972 (N_7972,N_7684,N_7542);
xor U7973 (N_7973,N_7519,N_7701);
nand U7974 (N_7974,N_7683,N_7705);
or U7975 (N_7975,N_7714,N_7616);
or U7976 (N_7976,N_7654,N_7659);
and U7977 (N_7977,N_7608,N_7626);
nand U7978 (N_7978,N_7735,N_7585);
and U7979 (N_7979,N_7510,N_7519);
or U7980 (N_7980,N_7685,N_7713);
xnor U7981 (N_7981,N_7500,N_7660);
xnor U7982 (N_7982,N_7528,N_7727);
xnor U7983 (N_7983,N_7585,N_7679);
and U7984 (N_7984,N_7549,N_7737);
nand U7985 (N_7985,N_7560,N_7515);
or U7986 (N_7986,N_7557,N_7586);
or U7987 (N_7987,N_7643,N_7577);
nor U7988 (N_7988,N_7705,N_7543);
or U7989 (N_7989,N_7727,N_7587);
nor U7990 (N_7990,N_7630,N_7621);
nand U7991 (N_7991,N_7685,N_7730);
and U7992 (N_7992,N_7592,N_7711);
nor U7993 (N_7993,N_7628,N_7636);
or U7994 (N_7994,N_7565,N_7621);
xnor U7995 (N_7995,N_7638,N_7631);
or U7996 (N_7996,N_7731,N_7743);
nor U7997 (N_7997,N_7720,N_7583);
nor U7998 (N_7998,N_7680,N_7689);
xor U7999 (N_7999,N_7617,N_7533);
or U8000 (N_8000,N_7865,N_7881);
xor U8001 (N_8001,N_7960,N_7959);
and U8002 (N_8002,N_7769,N_7891);
nand U8003 (N_8003,N_7793,N_7836);
nand U8004 (N_8004,N_7958,N_7977);
nand U8005 (N_8005,N_7906,N_7874);
nand U8006 (N_8006,N_7777,N_7939);
or U8007 (N_8007,N_7817,N_7890);
or U8008 (N_8008,N_7967,N_7846);
or U8009 (N_8009,N_7822,N_7909);
xnor U8010 (N_8010,N_7968,N_7912);
or U8011 (N_8011,N_7987,N_7843);
and U8012 (N_8012,N_7823,N_7767);
and U8013 (N_8013,N_7762,N_7980);
and U8014 (N_8014,N_7857,N_7768);
nor U8015 (N_8015,N_7872,N_7933);
xnor U8016 (N_8016,N_7819,N_7898);
nand U8017 (N_8017,N_7760,N_7855);
xor U8018 (N_8018,N_7908,N_7814);
xor U8019 (N_8019,N_7896,N_7991);
and U8020 (N_8020,N_7884,N_7785);
xnor U8021 (N_8021,N_7950,N_7880);
and U8022 (N_8022,N_7985,N_7752);
nand U8023 (N_8023,N_7876,N_7918);
xnor U8024 (N_8024,N_7799,N_7756);
xnor U8025 (N_8025,N_7816,N_7835);
nor U8026 (N_8026,N_7784,N_7791);
and U8027 (N_8027,N_7910,N_7834);
xnor U8028 (N_8028,N_7928,N_7911);
or U8029 (N_8029,N_7848,N_7839);
or U8030 (N_8030,N_7921,N_7922);
or U8031 (N_8031,N_7947,N_7753);
nor U8032 (N_8032,N_7946,N_7829);
xor U8033 (N_8033,N_7774,N_7997);
xnor U8034 (N_8034,N_7783,N_7900);
xnor U8035 (N_8035,N_7955,N_7897);
or U8036 (N_8036,N_7779,N_7901);
nand U8037 (N_8037,N_7929,N_7869);
xnor U8038 (N_8038,N_7805,N_7969);
xnor U8039 (N_8039,N_7943,N_7917);
xor U8040 (N_8040,N_7919,N_7804);
nor U8041 (N_8041,N_7830,N_7831);
xor U8042 (N_8042,N_7871,N_7966);
nand U8043 (N_8043,N_7931,N_7889);
and U8044 (N_8044,N_7993,N_7974);
nand U8045 (N_8045,N_7838,N_7941);
nand U8046 (N_8046,N_7851,N_7965);
and U8047 (N_8047,N_7826,N_7860);
or U8048 (N_8048,N_7853,N_7759);
and U8049 (N_8049,N_7914,N_7798);
xor U8050 (N_8050,N_7766,N_7988);
nand U8051 (N_8051,N_7878,N_7961);
and U8052 (N_8052,N_7953,N_7778);
xor U8053 (N_8053,N_7780,N_7757);
and U8054 (N_8054,N_7932,N_7875);
or U8055 (N_8055,N_7786,N_7776);
xor U8056 (N_8056,N_7802,N_7975);
or U8057 (N_8057,N_7982,N_7934);
nor U8058 (N_8058,N_7821,N_7925);
xnor U8059 (N_8059,N_7942,N_7755);
xor U8060 (N_8060,N_7847,N_7809);
xor U8061 (N_8061,N_7894,N_7832);
xor U8062 (N_8062,N_7840,N_7818);
nand U8063 (N_8063,N_7984,N_7842);
nor U8064 (N_8064,N_7983,N_7949);
nand U8065 (N_8065,N_7770,N_7892);
and U8066 (N_8066,N_7820,N_7913);
nor U8067 (N_8067,N_7926,N_7996);
xnor U8068 (N_8068,N_7761,N_7915);
nor U8069 (N_8069,N_7886,N_7981);
nor U8070 (N_8070,N_7999,N_7879);
nand U8071 (N_8071,N_7994,N_7899);
nand U8072 (N_8072,N_7751,N_7863);
or U8073 (N_8073,N_7864,N_7870);
nor U8074 (N_8074,N_7877,N_7893);
xor U8075 (N_8075,N_7807,N_7989);
nand U8076 (N_8076,N_7775,N_7963);
xnor U8077 (N_8077,N_7923,N_7945);
nor U8078 (N_8078,N_7765,N_7808);
nor U8079 (N_8079,N_7992,N_7764);
nand U8080 (N_8080,N_7986,N_7868);
or U8081 (N_8081,N_7858,N_7976);
nand U8082 (N_8082,N_7979,N_7907);
or U8083 (N_8083,N_7773,N_7781);
xnor U8084 (N_8084,N_7971,N_7867);
nand U8085 (N_8085,N_7973,N_7935);
xnor U8086 (N_8086,N_7957,N_7970);
and U8087 (N_8087,N_7990,N_7803);
nor U8088 (N_8088,N_7978,N_7888);
xnor U8089 (N_8089,N_7861,N_7924);
nand U8090 (N_8090,N_7854,N_7902);
and U8091 (N_8091,N_7948,N_7862);
or U8092 (N_8092,N_7885,N_7782);
xnor U8093 (N_8093,N_7859,N_7952);
and U8094 (N_8094,N_7873,N_7824);
nand U8095 (N_8095,N_7937,N_7837);
nor U8096 (N_8096,N_7811,N_7962);
xnor U8097 (N_8097,N_7795,N_7972);
xor U8098 (N_8098,N_7828,N_7845);
nor U8099 (N_8099,N_7936,N_7882);
nand U8100 (N_8100,N_7849,N_7850);
nor U8101 (N_8101,N_7763,N_7800);
nand U8102 (N_8102,N_7788,N_7792);
xor U8103 (N_8103,N_7787,N_7954);
or U8104 (N_8104,N_7940,N_7951);
nand U8105 (N_8105,N_7927,N_7806);
and U8106 (N_8106,N_7813,N_7772);
nand U8107 (N_8107,N_7797,N_7789);
nor U8108 (N_8108,N_7758,N_7930);
xor U8109 (N_8109,N_7916,N_7844);
or U8110 (N_8110,N_7903,N_7841);
nor U8111 (N_8111,N_7771,N_7956);
nor U8112 (N_8112,N_7883,N_7796);
or U8113 (N_8113,N_7852,N_7825);
nand U8114 (N_8114,N_7920,N_7754);
and U8115 (N_8115,N_7810,N_7964);
and U8116 (N_8116,N_7866,N_7944);
and U8117 (N_8117,N_7938,N_7998);
xor U8118 (N_8118,N_7833,N_7827);
and U8119 (N_8119,N_7815,N_7856);
nand U8120 (N_8120,N_7895,N_7812);
or U8121 (N_8121,N_7790,N_7801);
nor U8122 (N_8122,N_7995,N_7750);
nor U8123 (N_8123,N_7905,N_7904);
nand U8124 (N_8124,N_7887,N_7794);
xnor U8125 (N_8125,N_7806,N_7864);
and U8126 (N_8126,N_7910,N_7857);
or U8127 (N_8127,N_7773,N_7872);
nand U8128 (N_8128,N_7825,N_7811);
or U8129 (N_8129,N_7928,N_7934);
xnor U8130 (N_8130,N_7875,N_7862);
nand U8131 (N_8131,N_7759,N_7824);
nand U8132 (N_8132,N_7832,N_7937);
nor U8133 (N_8133,N_7845,N_7858);
nor U8134 (N_8134,N_7859,N_7953);
nor U8135 (N_8135,N_7994,N_7904);
nand U8136 (N_8136,N_7990,N_7753);
nand U8137 (N_8137,N_7792,N_7859);
xnor U8138 (N_8138,N_7924,N_7998);
xor U8139 (N_8139,N_7907,N_7767);
nor U8140 (N_8140,N_7896,N_7881);
nor U8141 (N_8141,N_7778,N_7929);
and U8142 (N_8142,N_7901,N_7781);
and U8143 (N_8143,N_7812,N_7863);
nor U8144 (N_8144,N_7917,N_7982);
xnor U8145 (N_8145,N_7961,N_7912);
nand U8146 (N_8146,N_7914,N_7882);
or U8147 (N_8147,N_7910,N_7904);
xnor U8148 (N_8148,N_7938,N_7882);
nor U8149 (N_8149,N_7901,N_7840);
xor U8150 (N_8150,N_7929,N_7777);
nand U8151 (N_8151,N_7853,N_7856);
or U8152 (N_8152,N_7873,N_7970);
and U8153 (N_8153,N_7882,N_7869);
or U8154 (N_8154,N_7972,N_7988);
nand U8155 (N_8155,N_7770,N_7763);
nand U8156 (N_8156,N_7951,N_7993);
nand U8157 (N_8157,N_7836,N_7849);
and U8158 (N_8158,N_7818,N_7995);
and U8159 (N_8159,N_7771,N_7819);
or U8160 (N_8160,N_7827,N_7957);
xor U8161 (N_8161,N_7977,N_7910);
or U8162 (N_8162,N_7811,N_7862);
xor U8163 (N_8163,N_7762,N_7955);
xor U8164 (N_8164,N_7894,N_7986);
and U8165 (N_8165,N_7806,N_7940);
xor U8166 (N_8166,N_7973,N_7771);
nor U8167 (N_8167,N_7752,N_7883);
and U8168 (N_8168,N_7887,N_7888);
and U8169 (N_8169,N_7853,N_7836);
nand U8170 (N_8170,N_7870,N_7829);
or U8171 (N_8171,N_7958,N_7786);
nand U8172 (N_8172,N_7921,N_7908);
and U8173 (N_8173,N_7799,N_7827);
nor U8174 (N_8174,N_7783,N_7808);
or U8175 (N_8175,N_7989,N_7915);
nor U8176 (N_8176,N_7874,N_7845);
or U8177 (N_8177,N_7912,N_7948);
or U8178 (N_8178,N_7965,N_7989);
nand U8179 (N_8179,N_7877,N_7803);
nor U8180 (N_8180,N_7756,N_7901);
and U8181 (N_8181,N_7814,N_7776);
nand U8182 (N_8182,N_7816,N_7938);
and U8183 (N_8183,N_7921,N_7818);
xor U8184 (N_8184,N_7924,N_7917);
and U8185 (N_8185,N_7890,N_7810);
and U8186 (N_8186,N_7926,N_7866);
and U8187 (N_8187,N_7751,N_7825);
xnor U8188 (N_8188,N_7836,N_7896);
xor U8189 (N_8189,N_7877,N_7772);
nor U8190 (N_8190,N_7867,N_7917);
nor U8191 (N_8191,N_7787,N_7826);
xor U8192 (N_8192,N_7945,N_7858);
or U8193 (N_8193,N_7867,N_7946);
xor U8194 (N_8194,N_7953,N_7878);
or U8195 (N_8195,N_7904,N_7854);
nor U8196 (N_8196,N_7768,N_7781);
nand U8197 (N_8197,N_7859,N_7969);
and U8198 (N_8198,N_7850,N_7861);
or U8199 (N_8199,N_7805,N_7795);
or U8200 (N_8200,N_7929,N_7764);
xnor U8201 (N_8201,N_7780,N_7777);
xnor U8202 (N_8202,N_7944,N_7975);
nor U8203 (N_8203,N_7801,N_7841);
nor U8204 (N_8204,N_7827,N_7951);
nor U8205 (N_8205,N_7978,N_7923);
nor U8206 (N_8206,N_7830,N_7885);
nand U8207 (N_8207,N_7995,N_7874);
nand U8208 (N_8208,N_7857,N_7752);
xor U8209 (N_8209,N_7825,N_7913);
xor U8210 (N_8210,N_7932,N_7893);
and U8211 (N_8211,N_7869,N_7876);
nor U8212 (N_8212,N_7846,N_7855);
or U8213 (N_8213,N_7858,N_7846);
nand U8214 (N_8214,N_7956,N_7810);
xnor U8215 (N_8215,N_7890,N_7771);
or U8216 (N_8216,N_7788,N_7893);
or U8217 (N_8217,N_7971,N_7801);
xor U8218 (N_8218,N_7931,N_7777);
and U8219 (N_8219,N_7783,N_7837);
nor U8220 (N_8220,N_7842,N_7866);
nand U8221 (N_8221,N_7779,N_7948);
nand U8222 (N_8222,N_7873,N_7909);
nor U8223 (N_8223,N_7919,N_7906);
and U8224 (N_8224,N_7786,N_7890);
or U8225 (N_8225,N_7967,N_7761);
or U8226 (N_8226,N_7897,N_7962);
or U8227 (N_8227,N_7972,N_7904);
or U8228 (N_8228,N_7755,N_7821);
xnor U8229 (N_8229,N_7843,N_7952);
nand U8230 (N_8230,N_7798,N_7857);
nand U8231 (N_8231,N_7894,N_7870);
nand U8232 (N_8232,N_7975,N_7928);
nor U8233 (N_8233,N_7964,N_7780);
nor U8234 (N_8234,N_7880,N_7948);
nand U8235 (N_8235,N_7919,N_7898);
nand U8236 (N_8236,N_7902,N_7990);
nor U8237 (N_8237,N_7797,N_7829);
xnor U8238 (N_8238,N_7783,N_7980);
and U8239 (N_8239,N_7937,N_7826);
xor U8240 (N_8240,N_7856,N_7763);
nor U8241 (N_8241,N_7788,N_7877);
nand U8242 (N_8242,N_7885,N_7905);
or U8243 (N_8243,N_7763,N_7772);
xor U8244 (N_8244,N_7787,N_7818);
or U8245 (N_8245,N_7989,N_7963);
nand U8246 (N_8246,N_7894,N_7919);
xnor U8247 (N_8247,N_7759,N_7750);
nand U8248 (N_8248,N_7983,N_7811);
nand U8249 (N_8249,N_7991,N_7944);
and U8250 (N_8250,N_8162,N_8115);
and U8251 (N_8251,N_8224,N_8113);
and U8252 (N_8252,N_8069,N_8022);
or U8253 (N_8253,N_8174,N_8144);
or U8254 (N_8254,N_8193,N_8038);
nor U8255 (N_8255,N_8017,N_8195);
xnor U8256 (N_8256,N_8083,N_8192);
or U8257 (N_8257,N_8033,N_8056);
or U8258 (N_8258,N_8212,N_8152);
and U8259 (N_8259,N_8126,N_8078);
and U8260 (N_8260,N_8114,N_8238);
nand U8261 (N_8261,N_8156,N_8211);
nand U8262 (N_8262,N_8042,N_8041);
nand U8263 (N_8263,N_8050,N_8019);
xor U8264 (N_8264,N_8004,N_8121);
nand U8265 (N_8265,N_8061,N_8150);
xor U8266 (N_8266,N_8124,N_8007);
or U8267 (N_8267,N_8190,N_8170);
xnor U8268 (N_8268,N_8220,N_8165);
nor U8269 (N_8269,N_8117,N_8024);
xnor U8270 (N_8270,N_8227,N_8160);
nand U8271 (N_8271,N_8099,N_8134);
nor U8272 (N_8272,N_8239,N_8157);
xor U8273 (N_8273,N_8025,N_8008);
nand U8274 (N_8274,N_8182,N_8068);
nor U8275 (N_8275,N_8085,N_8035);
xnor U8276 (N_8276,N_8032,N_8149);
and U8277 (N_8277,N_8072,N_8058);
xnor U8278 (N_8278,N_8073,N_8055);
xnor U8279 (N_8279,N_8111,N_8026);
and U8280 (N_8280,N_8218,N_8013);
xnor U8281 (N_8281,N_8234,N_8060);
or U8282 (N_8282,N_8082,N_8015);
nand U8283 (N_8283,N_8161,N_8005);
or U8284 (N_8284,N_8120,N_8003);
nor U8285 (N_8285,N_8171,N_8226);
nor U8286 (N_8286,N_8028,N_8009);
or U8287 (N_8287,N_8070,N_8228);
and U8288 (N_8288,N_8065,N_8048);
and U8289 (N_8289,N_8179,N_8040);
and U8290 (N_8290,N_8000,N_8016);
nor U8291 (N_8291,N_8147,N_8063);
and U8292 (N_8292,N_8027,N_8184);
or U8293 (N_8293,N_8046,N_8047);
xnor U8294 (N_8294,N_8225,N_8062);
nor U8295 (N_8295,N_8189,N_8088);
and U8296 (N_8296,N_8232,N_8103);
xnor U8297 (N_8297,N_8104,N_8107);
or U8298 (N_8298,N_8079,N_8138);
xnor U8299 (N_8299,N_8209,N_8136);
xor U8300 (N_8300,N_8213,N_8164);
nand U8301 (N_8301,N_8178,N_8173);
nand U8302 (N_8302,N_8119,N_8202);
nand U8303 (N_8303,N_8175,N_8148);
or U8304 (N_8304,N_8181,N_8044);
and U8305 (N_8305,N_8131,N_8118);
nand U8306 (N_8306,N_8166,N_8177);
nor U8307 (N_8307,N_8203,N_8030);
and U8308 (N_8308,N_8123,N_8154);
nor U8309 (N_8309,N_8219,N_8102);
or U8310 (N_8310,N_8122,N_8116);
nand U8311 (N_8311,N_8172,N_8045);
or U8312 (N_8312,N_8110,N_8183);
xnor U8313 (N_8313,N_8106,N_8043);
and U8314 (N_8314,N_8034,N_8204);
and U8315 (N_8315,N_8018,N_8101);
xor U8316 (N_8316,N_8249,N_8021);
xnor U8317 (N_8317,N_8080,N_8037);
nand U8318 (N_8318,N_8067,N_8094);
nand U8319 (N_8319,N_8205,N_8247);
xnor U8320 (N_8320,N_8053,N_8127);
or U8321 (N_8321,N_8141,N_8071);
nor U8322 (N_8322,N_8095,N_8243);
and U8323 (N_8323,N_8169,N_8155);
or U8324 (N_8324,N_8105,N_8158);
and U8325 (N_8325,N_8133,N_8167);
xnor U8326 (N_8326,N_8198,N_8240);
or U8327 (N_8327,N_8229,N_8130);
or U8328 (N_8328,N_8143,N_8200);
and U8329 (N_8329,N_8207,N_8168);
nor U8330 (N_8330,N_8153,N_8074);
or U8331 (N_8331,N_8146,N_8129);
nor U8332 (N_8332,N_8230,N_8010);
xnor U8333 (N_8333,N_8093,N_8235);
xor U8334 (N_8334,N_8020,N_8180);
nor U8335 (N_8335,N_8215,N_8151);
and U8336 (N_8336,N_8187,N_8197);
nand U8337 (N_8337,N_8011,N_8191);
nor U8338 (N_8338,N_8208,N_8039);
nand U8339 (N_8339,N_8236,N_8201);
xor U8340 (N_8340,N_8223,N_8217);
and U8341 (N_8341,N_8241,N_8242);
or U8342 (N_8342,N_8214,N_8096);
xnor U8343 (N_8343,N_8087,N_8098);
and U8344 (N_8344,N_8051,N_8145);
and U8345 (N_8345,N_8091,N_8128);
or U8346 (N_8346,N_8075,N_8066);
or U8347 (N_8347,N_8139,N_8142);
nand U8348 (N_8348,N_8132,N_8108);
xor U8349 (N_8349,N_8206,N_8186);
and U8350 (N_8350,N_8163,N_8216);
nand U8351 (N_8351,N_8248,N_8244);
nand U8352 (N_8352,N_8237,N_8023);
and U8353 (N_8353,N_8222,N_8233);
nor U8354 (N_8354,N_8006,N_8185);
xor U8355 (N_8355,N_8064,N_8002);
nor U8356 (N_8356,N_8092,N_8081);
nor U8357 (N_8357,N_8176,N_8196);
nand U8358 (N_8358,N_8001,N_8090);
nand U8359 (N_8359,N_8012,N_8245);
nand U8360 (N_8360,N_8031,N_8086);
or U8361 (N_8361,N_8231,N_8057);
xor U8362 (N_8362,N_8059,N_8077);
or U8363 (N_8363,N_8221,N_8159);
nor U8364 (N_8364,N_8135,N_8109);
nand U8365 (N_8365,N_8188,N_8029);
nand U8366 (N_8366,N_8049,N_8137);
and U8367 (N_8367,N_8199,N_8246);
and U8368 (N_8368,N_8097,N_8052);
or U8369 (N_8369,N_8076,N_8014);
nor U8370 (N_8370,N_8054,N_8100);
xnor U8371 (N_8371,N_8112,N_8036);
and U8372 (N_8372,N_8140,N_8194);
or U8373 (N_8373,N_8125,N_8210);
xnor U8374 (N_8374,N_8084,N_8089);
and U8375 (N_8375,N_8183,N_8108);
nand U8376 (N_8376,N_8200,N_8024);
or U8377 (N_8377,N_8037,N_8151);
and U8378 (N_8378,N_8137,N_8153);
nor U8379 (N_8379,N_8145,N_8244);
nand U8380 (N_8380,N_8157,N_8014);
or U8381 (N_8381,N_8009,N_8066);
or U8382 (N_8382,N_8152,N_8241);
nor U8383 (N_8383,N_8119,N_8139);
xnor U8384 (N_8384,N_8197,N_8087);
xnor U8385 (N_8385,N_8045,N_8137);
and U8386 (N_8386,N_8023,N_8218);
nand U8387 (N_8387,N_8170,N_8065);
nor U8388 (N_8388,N_8151,N_8213);
and U8389 (N_8389,N_8000,N_8120);
xor U8390 (N_8390,N_8202,N_8067);
nand U8391 (N_8391,N_8115,N_8136);
nand U8392 (N_8392,N_8100,N_8178);
and U8393 (N_8393,N_8246,N_8132);
or U8394 (N_8394,N_8182,N_8053);
and U8395 (N_8395,N_8030,N_8220);
nand U8396 (N_8396,N_8238,N_8117);
and U8397 (N_8397,N_8108,N_8028);
xor U8398 (N_8398,N_8226,N_8072);
xor U8399 (N_8399,N_8059,N_8121);
nand U8400 (N_8400,N_8132,N_8045);
and U8401 (N_8401,N_8198,N_8010);
nand U8402 (N_8402,N_8048,N_8014);
or U8403 (N_8403,N_8076,N_8185);
nor U8404 (N_8404,N_8075,N_8121);
nand U8405 (N_8405,N_8213,N_8142);
nand U8406 (N_8406,N_8090,N_8149);
xnor U8407 (N_8407,N_8153,N_8128);
xnor U8408 (N_8408,N_8187,N_8202);
or U8409 (N_8409,N_8003,N_8090);
xor U8410 (N_8410,N_8004,N_8199);
and U8411 (N_8411,N_8234,N_8010);
and U8412 (N_8412,N_8138,N_8015);
nand U8413 (N_8413,N_8181,N_8213);
nand U8414 (N_8414,N_8074,N_8035);
nand U8415 (N_8415,N_8117,N_8049);
nor U8416 (N_8416,N_8033,N_8232);
or U8417 (N_8417,N_8224,N_8019);
and U8418 (N_8418,N_8099,N_8011);
or U8419 (N_8419,N_8173,N_8007);
or U8420 (N_8420,N_8053,N_8010);
nand U8421 (N_8421,N_8100,N_8109);
nand U8422 (N_8422,N_8006,N_8149);
or U8423 (N_8423,N_8022,N_8233);
nor U8424 (N_8424,N_8064,N_8069);
or U8425 (N_8425,N_8106,N_8072);
or U8426 (N_8426,N_8064,N_8232);
nor U8427 (N_8427,N_8083,N_8233);
nor U8428 (N_8428,N_8234,N_8147);
and U8429 (N_8429,N_8112,N_8029);
xor U8430 (N_8430,N_8188,N_8079);
and U8431 (N_8431,N_8224,N_8043);
and U8432 (N_8432,N_8150,N_8146);
or U8433 (N_8433,N_8055,N_8115);
xor U8434 (N_8434,N_8095,N_8067);
nand U8435 (N_8435,N_8055,N_8158);
xnor U8436 (N_8436,N_8009,N_8180);
or U8437 (N_8437,N_8078,N_8220);
nand U8438 (N_8438,N_8150,N_8051);
and U8439 (N_8439,N_8189,N_8194);
or U8440 (N_8440,N_8161,N_8118);
xnor U8441 (N_8441,N_8013,N_8066);
nor U8442 (N_8442,N_8177,N_8069);
nand U8443 (N_8443,N_8146,N_8126);
xnor U8444 (N_8444,N_8165,N_8002);
nand U8445 (N_8445,N_8200,N_8035);
nor U8446 (N_8446,N_8106,N_8234);
xor U8447 (N_8447,N_8072,N_8046);
nand U8448 (N_8448,N_8105,N_8032);
nand U8449 (N_8449,N_8125,N_8134);
xor U8450 (N_8450,N_8172,N_8090);
and U8451 (N_8451,N_8048,N_8170);
xor U8452 (N_8452,N_8022,N_8079);
and U8453 (N_8453,N_8151,N_8089);
or U8454 (N_8454,N_8060,N_8048);
nand U8455 (N_8455,N_8120,N_8149);
nor U8456 (N_8456,N_8050,N_8021);
nor U8457 (N_8457,N_8065,N_8082);
xor U8458 (N_8458,N_8116,N_8008);
xnor U8459 (N_8459,N_8183,N_8098);
xor U8460 (N_8460,N_8042,N_8161);
or U8461 (N_8461,N_8052,N_8235);
xnor U8462 (N_8462,N_8098,N_8029);
or U8463 (N_8463,N_8116,N_8208);
or U8464 (N_8464,N_8024,N_8207);
nand U8465 (N_8465,N_8030,N_8053);
or U8466 (N_8466,N_8116,N_8135);
nor U8467 (N_8467,N_8038,N_8022);
nand U8468 (N_8468,N_8104,N_8244);
or U8469 (N_8469,N_8145,N_8224);
or U8470 (N_8470,N_8051,N_8213);
xor U8471 (N_8471,N_8221,N_8078);
nand U8472 (N_8472,N_8077,N_8115);
nor U8473 (N_8473,N_8055,N_8239);
nor U8474 (N_8474,N_8081,N_8220);
nor U8475 (N_8475,N_8011,N_8228);
nand U8476 (N_8476,N_8172,N_8088);
nor U8477 (N_8477,N_8004,N_8042);
and U8478 (N_8478,N_8116,N_8037);
nand U8479 (N_8479,N_8140,N_8063);
or U8480 (N_8480,N_8023,N_8102);
nand U8481 (N_8481,N_8013,N_8024);
and U8482 (N_8482,N_8057,N_8139);
nor U8483 (N_8483,N_8248,N_8242);
nand U8484 (N_8484,N_8046,N_8035);
xnor U8485 (N_8485,N_8096,N_8105);
or U8486 (N_8486,N_8156,N_8129);
or U8487 (N_8487,N_8149,N_8072);
nand U8488 (N_8488,N_8094,N_8168);
nand U8489 (N_8489,N_8190,N_8090);
nor U8490 (N_8490,N_8044,N_8248);
xnor U8491 (N_8491,N_8093,N_8167);
or U8492 (N_8492,N_8048,N_8112);
and U8493 (N_8493,N_8065,N_8197);
or U8494 (N_8494,N_8151,N_8123);
nand U8495 (N_8495,N_8066,N_8111);
xnor U8496 (N_8496,N_8123,N_8218);
nor U8497 (N_8497,N_8172,N_8157);
nor U8498 (N_8498,N_8247,N_8017);
xnor U8499 (N_8499,N_8114,N_8142);
and U8500 (N_8500,N_8462,N_8330);
or U8501 (N_8501,N_8386,N_8398);
xor U8502 (N_8502,N_8451,N_8434);
and U8503 (N_8503,N_8322,N_8353);
nor U8504 (N_8504,N_8362,N_8358);
and U8505 (N_8505,N_8418,N_8277);
and U8506 (N_8506,N_8493,N_8416);
xor U8507 (N_8507,N_8412,N_8389);
nor U8508 (N_8508,N_8490,N_8421);
or U8509 (N_8509,N_8297,N_8305);
nand U8510 (N_8510,N_8361,N_8365);
nand U8511 (N_8511,N_8474,N_8431);
nand U8512 (N_8512,N_8308,N_8454);
xor U8513 (N_8513,N_8479,N_8435);
or U8514 (N_8514,N_8400,N_8376);
nor U8515 (N_8515,N_8284,N_8312);
and U8516 (N_8516,N_8496,N_8494);
and U8517 (N_8517,N_8366,N_8269);
or U8518 (N_8518,N_8430,N_8285);
and U8519 (N_8519,N_8280,N_8283);
xor U8520 (N_8520,N_8360,N_8293);
and U8521 (N_8521,N_8448,N_8380);
or U8522 (N_8522,N_8304,N_8393);
nor U8523 (N_8523,N_8488,N_8267);
nand U8524 (N_8524,N_8388,N_8282);
nand U8525 (N_8525,N_8429,N_8492);
nor U8526 (N_8526,N_8368,N_8455);
and U8527 (N_8527,N_8468,N_8327);
xor U8528 (N_8528,N_8343,N_8445);
nor U8529 (N_8529,N_8325,N_8346);
or U8530 (N_8530,N_8423,N_8347);
xnor U8531 (N_8531,N_8495,N_8254);
and U8532 (N_8532,N_8310,N_8324);
nand U8533 (N_8533,N_8291,N_8279);
nand U8534 (N_8534,N_8301,N_8344);
nand U8535 (N_8535,N_8482,N_8475);
and U8536 (N_8536,N_8403,N_8485);
xnor U8537 (N_8537,N_8471,N_8384);
nor U8538 (N_8538,N_8261,N_8401);
nand U8539 (N_8539,N_8436,N_8422);
nor U8540 (N_8540,N_8300,N_8369);
xor U8541 (N_8541,N_8337,N_8395);
nand U8542 (N_8542,N_8316,N_8409);
xor U8543 (N_8543,N_8264,N_8491);
nor U8544 (N_8544,N_8320,N_8356);
xor U8545 (N_8545,N_8457,N_8394);
nor U8546 (N_8546,N_8273,N_8306);
or U8547 (N_8547,N_8397,N_8498);
xor U8548 (N_8548,N_8458,N_8499);
nand U8549 (N_8549,N_8303,N_8456);
nand U8550 (N_8550,N_8335,N_8315);
or U8551 (N_8551,N_8323,N_8417);
nand U8552 (N_8552,N_8378,N_8363);
nor U8553 (N_8553,N_8294,N_8481);
or U8554 (N_8554,N_8274,N_8486);
nand U8555 (N_8555,N_8326,N_8396);
and U8556 (N_8556,N_8357,N_8390);
or U8557 (N_8557,N_8450,N_8428);
nor U8558 (N_8558,N_8253,N_8317);
or U8559 (N_8559,N_8404,N_8460);
nand U8560 (N_8560,N_8387,N_8374);
and U8561 (N_8561,N_8392,N_8379);
xor U8562 (N_8562,N_8381,N_8426);
nand U8563 (N_8563,N_8408,N_8453);
nor U8564 (N_8564,N_8497,N_8487);
nor U8565 (N_8565,N_8255,N_8336);
or U8566 (N_8566,N_8351,N_8465);
nand U8567 (N_8567,N_8333,N_8250);
nor U8568 (N_8568,N_8367,N_8260);
nand U8569 (N_8569,N_8289,N_8359);
and U8570 (N_8570,N_8287,N_8463);
nor U8571 (N_8571,N_8372,N_8473);
xnor U8572 (N_8572,N_8257,N_8470);
or U8573 (N_8573,N_8272,N_8447);
nand U8574 (N_8574,N_8268,N_8349);
nor U8575 (N_8575,N_8484,N_8371);
nand U8576 (N_8576,N_8328,N_8410);
or U8577 (N_8577,N_8437,N_8307);
nand U8578 (N_8578,N_8442,N_8318);
and U8579 (N_8579,N_8278,N_8443);
and U8580 (N_8580,N_8399,N_8414);
xnor U8581 (N_8581,N_8281,N_8413);
xor U8582 (N_8582,N_8266,N_8252);
and U8583 (N_8583,N_8292,N_8433);
nand U8584 (N_8584,N_8461,N_8407);
or U8585 (N_8585,N_8298,N_8377);
xnor U8586 (N_8586,N_8352,N_8342);
and U8587 (N_8587,N_8329,N_8364);
nand U8588 (N_8588,N_8478,N_8286);
xnor U8589 (N_8589,N_8424,N_8469);
nor U8590 (N_8590,N_8313,N_8391);
and U8591 (N_8591,N_8348,N_8340);
and U8592 (N_8592,N_8476,N_8402);
or U8593 (N_8593,N_8405,N_8373);
or U8594 (N_8594,N_8472,N_8262);
and U8595 (N_8595,N_8295,N_8275);
xor U8596 (N_8596,N_8263,N_8420);
xnor U8597 (N_8597,N_8444,N_8258);
nor U8598 (N_8598,N_8467,N_8332);
or U8599 (N_8599,N_8382,N_8383);
and U8600 (N_8600,N_8350,N_8319);
xnor U8601 (N_8601,N_8464,N_8341);
or U8602 (N_8602,N_8321,N_8276);
nor U8603 (N_8603,N_8425,N_8345);
nand U8604 (N_8604,N_8489,N_8370);
nor U8605 (N_8605,N_8375,N_8338);
and U8606 (N_8606,N_8339,N_8256);
nand U8607 (N_8607,N_8480,N_8432);
and U8608 (N_8608,N_8296,N_8415);
nor U8609 (N_8609,N_8411,N_8251);
nand U8610 (N_8610,N_8299,N_8452);
nor U8611 (N_8611,N_8441,N_8314);
and U8612 (N_8612,N_8290,N_8302);
nand U8613 (N_8613,N_8259,N_8311);
xor U8614 (N_8614,N_8483,N_8354);
or U8615 (N_8615,N_8406,N_8309);
and U8616 (N_8616,N_8427,N_8355);
nand U8617 (N_8617,N_8440,N_8265);
nor U8618 (N_8618,N_8466,N_8439);
or U8619 (N_8619,N_8288,N_8449);
nor U8620 (N_8620,N_8270,N_8334);
nor U8621 (N_8621,N_8459,N_8446);
or U8622 (N_8622,N_8477,N_8438);
nor U8623 (N_8623,N_8385,N_8331);
and U8624 (N_8624,N_8271,N_8419);
or U8625 (N_8625,N_8422,N_8277);
nor U8626 (N_8626,N_8499,N_8496);
or U8627 (N_8627,N_8450,N_8318);
xor U8628 (N_8628,N_8357,N_8277);
and U8629 (N_8629,N_8386,N_8406);
nor U8630 (N_8630,N_8313,N_8327);
nand U8631 (N_8631,N_8398,N_8252);
nand U8632 (N_8632,N_8454,N_8466);
nor U8633 (N_8633,N_8405,N_8425);
xnor U8634 (N_8634,N_8315,N_8383);
or U8635 (N_8635,N_8385,N_8323);
and U8636 (N_8636,N_8469,N_8357);
or U8637 (N_8637,N_8367,N_8372);
or U8638 (N_8638,N_8399,N_8351);
xor U8639 (N_8639,N_8254,N_8465);
and U8640 (N_8640,N_8447,N_8470);
nand U8641 (N_8641,N_8422,N_8493);
xor U8642 (N_8642,N_8323,N_8357);
nand U8643 (N_8643,N_8250,N_8499);
nand U8644 (N_8644,N_8275,N_8447);
and U8645 (N_8645,N_8346,N_8479);
or U8646 (N_8646,N_8464,N_8390);
nor U8647 (N_8647,N_8454,N_8403);
nand U8648 (N_8648,N_8318,N_8281);
or U8649 (N_8649,N_8429,N_8363);
nor U8650 (N_8650,N_8343,N_8334);
nand U8651 (N_8651,N_8326,N_8415);
nand U8652 (N_8652,N_8335,N_8297);
or U8653 (N_8653,N_8408,N_8435);
or U8654 (N_8654,N_8322,N_8313);
or U8655 (N_8655,N_8334,N_8308);
xor U8656 (N_8656,N_8411,N_8334);
and U8657 (N_8657,N_8326,N_8257);
and U8658 (N_8658,N_8272,N_8313);
nand U8659 (N_8659,N_8440,N_8266);
nand U8660 (N_8660,N_8499,N_8311);
and U8661 (N_8661,N_8294,N_8311);
xor U8662 (N_8662,N_8499,N_8397);
or U8663 (N_8663,N_8418,N_8485);
nor U8664 (N_8664,N_8317,N_8364);
xor U8665 (N_8665,N_8318,N_8353);
nand U8666 (N_8666,N_8301,N_8327);
xor U8667 (N_8667,N_8470,N_8314);
nor U8668 (N_8668,N_8259,N_8280);
and U8669 (N_8669,N_8471,N_8390);
and U8670 (N_8670,N_8294,N_8391);
or U8671 (N_8671,N_8421,N_8489);
xor U8672 (N_8672,N_8394,N_8274);
and U8673 (N_8673,N_8454,N_8413);
or U8674 (N_8674,N_8354,N_8325);
nor U8675 (N_8675,N_8334,N_8395);
and U8676 (N_8676,N_8400,N_8279);
and U8677 (N_8677,N_8281,N_8338);
or U8678 (N_8678,N_8271,N_8496);
xor U8679 (N_8679,N_8381,N_8344);
xnor U8680 (N_8680,N_8468,N_8442);
or U8681 (N_8681,N_8363,N_8276);
or U8682 (N_8682,N_8312,N_8296);
nand U8683 (N_8683,N_8465,N_8461);
xor U8684 (N_8684,N_8456,N_8396);
nand U8685 (N_8685,N_8405,N_8358);
xnor U8686 (N_8686,N_8292,N_8380);
xnor U8687 (N_8687,N_8456,N_8364);
nor U8688 (N_8688,N_8415,N_8392);
xnor U8689 (N_8689,N_8270,N_8329);
or U8690 (N_8690,N_8340,N_8401);
nand U8691 (N_8691,N_8390,N_8421);
nor U8692 (N_8692,N_8391,N_8380);
nor U8693 (N_8693,N_8442,N_8422);
nor U8694 (N_8694,N_8260,N_8464);
and U8695 (N_8695,N_8330,N_8347);
nand U8696 (N_8696,N_8419,N_8381);
xnor U8697 (N_8697,N_8449,N_8376);
nand U8698 (N_8698,N_8357,N_8495);
and U8699 (N_8699,N_8461,N_8428);
nor U8700 (N_8700,N_8270,N_8465);
nand U8701 (N_8701,N_8342,N_8455);
nand U8702 (N_8702,N_8413,N_8269);
nand U8703 (N_8703,N_8378,N_8310);
nor U8704 (N_8704,N_8294,N_8288);
or U8705 (N_8705,N_8463,N_8455);
xnor U8706 (N_8706,N_8293,N_8472);
xor U8707 (N_8707,N_8338,N_8376);
xor U8708 (N_8708,N_8448,N_8440);
nor U8709 (N_8709,N_8366,N_8399);
nor U8710 (N_8710,N_8479,N_8387);
nand U8711 (N_8711,N_8363,N_8332);
xnor U8712 (N_8712,N_8430,N_8363);
nor U8713 (N_8713,N_8359,N_8290);
xnor U8714 (N_8714,N_8496,N_8336);
or U8715 (N_8715,N_8343,N_8285);
and U8716 (N_8716,N_8298,N_8433);
or U8717 (N_8717,N_8361,N_8360);
or U8718 (N_8718,N_8391,N_8298);
and U8719 (N_8719,N_8478,N_8445);
nand U8720 (N_8720,N_8491,N_8396);
nor U8721 (N_8721,N_8497,N_8284);
or U8722 (N_8722,N_8463,N_8397);
xnor U8723 (N_8723,N_8484,N_8346);
and U8724 (N_8724,N_8379,N_8498);
xor U8725 (N_8725,N_8397,N_8491);
nor U8726 (N_8726,N_8388,N_8393);
or U8727 (N_8727,N_8448,N_8314);
nand U8728 (N_8728,N_8477,N_8309);
or U8729 (N_8729,N_8313,N_8368);
and U8730 (N_8730,N_8439,N_8277);
xnor U8731 (N_8731,N_8434,N_8340);
nor U8732 (N_8732,N_8314,N_8335);
or U8733 (N_8733,N_8478,N_8256);
and U8734 (N_8734,N_8287,N_8269);
nand U8735 (N_8735,N_8262,N_8473);
xor U8736 (N_8736,N_8308,N_8290);
nand U8737 (N_8737,N_8369,N_8322);
nand U8738 (N_8738,N_8295,N_8320);
xor U8739 (N_8739,N_8308,N_8387);
nand U8740 (N_8740,N_8408,N_8457);
and U8741 (N_8741,N_8378,N_8441);
or U8742 (N_8742,N_8461,N_8357);
and U8743 (N_8743,N_8360,N_8338);
nand U8744 (N_8744,N_8363,N_8420);
xnor U8745 (N_8745,N_8290,N_8259);
xnor U8746 (N_8746,N_8392,N_8461);
nand U8747 (N_8747,N_8394,N_8310);
xor U8748 (N_8748,N_8455,N_8471);
and U8749 (N_8749,N_8317,N_8341);
nor U8750 (N_8750,N_8649,N_8734);
xor U8751 (N_8751,N_8619,N_8676);
and U8752 (N_8752,N_8632,N_8665);
nand U8753 (N_8753,N_8741,N_8587);
and U8754 (N_8754,N_8535,N_8728);
or U8755 (N_8755,N_8575,N_8512);
and U8756 (N_8756,N_8723,N_8545);
nand U8757 (N_8757,N_8605,N_8613);
xnor U8758 (N_8758,N_8722,N_8530);
nand U8759 (N_8759,N_8670,N_8509);
xnor U8760 (N_8760,N_8745,N_8547);
nand U8761 (N_8761,N_8655,N_8663);
or U8762 (N_8762,N_8636,N_8556);
and U8763 (N_8763,N_8646,N_8560);
or U8764 (N_8764,N_8581,N_8580);
xnor U8765 (N_8765,N_8507,N_8710);
nand U8766 (N_8766,N_8682,N_8715);
nand U8767 (N_8767,N_8612,N_8548);
nor U8768 (N_8768,N_8572,N_8673);
or U8769 (N_8769,N_8600,N_8518);
or U8770 (N_8770,N_8533,N_8737);
xnor U8771 (N_8771,N_8594,N_8539);
nor U8772 (N_8772,N_8573,N_8576);
nand U8773 (N_8773,N_8521,N_8617);
or U8774 (N_8774,N_8569,N_8644);
xnor U8775 (N_8775,N_8583,N_8564);
nand U8776 (N_8776,N_8528,N_8584);
nor U8777 (N_8777,N_8510,N_8519);
nor U8778 (N_8778,N_8540,N_8597);
and U8779 (N_8779,N_8658,N_8708);
and U8780 (N_8780,N_8595,N_8546);
nor U8781 (N_8781,N_8659,N_8561);
xnor U8782 (N_8782,N_8668,N_8608);
and U8783 (N_8783,N_8610,N_8630);
nand U8784 (N_8784,N_8680,N_8589);
nand U8785 (N_8785,N_8701,N_8681);
or U8786 (N_8786,N_8622,N_8724);
nor U8787 (N_8787,N_8506,N_8667);
and U8788 (N_8788,N_8664,N_8558);
nand U8789 (N_8789,N_8672,N_8689);
xor U8790 (N_8790,N_8690,N_8542);
nand U8791 (N_8791,N_8679,N_8743);
nor U8792 (N_8792,N_8517,N_8567);
nand U8793 (N_8793,N_8727,N_8529);
nor U8794 (N_8794,N_8652,N_8603);
and U8795 (N_8795,N_8543,N_8733);
and U8796 (N_8796,N_8642,N_8643);
xnor U8797 (N_8797,N_8718,N_8588);
nand U8798 (N_8798,N_8691,N_8502);
nor U8799 (N_8799,N_8744,N_8515);
xor U8800 (N_8800,N_8732,N_8685);
nand U8801 (N_8801,N_8598,N_8639);
nor U8802 (N_8802,N_8522,N_8696);
and U8803 (N_8803,N_8505,N_8541);
nand U8804 (N_8804,N_8574,N_8514);
or U8805 (N_8805,N_8604,N_8503);
xnor U8806 (N_8806,N_8614,N_8633);
nor U8807 (N_8807,N_8693,N_8648);
xor U8808 (N_8808,N_8544,N_8531);
nor U8809 (N_8809,N_8534,N_8578);
or U8810 (N_8810,N_8730,N_8538);
nor U8811 (N_8811,N_8585,N_8717);
or U8812 (N_8812,N_8566,N_8686);
xnor U8813 (N_8813,N_8704,N_8735);
nor U8814 (N_8814,N_8635,N_8516);
nor U8815 (N_8815,N_8525,N_8562);
xnor U8816 (N_8816,N_8621,N_8638);
nor U8817 (N_8817,N_8592,N_8695);
and U8818 (N_8818,N_8713,N_8707);
nor U8819 (N_8819,N_8500,N_8729);
and U8820 (N_8820,N_8662,N_8523);
nand U8821 (N_8821,N_8669,N_8747);
nor U8822 (N_8822,N_8654,N_8563);
and U8823 (N_8823,N_8641,N_8684);
nor U8824 (N_8824,N_8615,N_8624);
nor U8825 (N_8825,N_8570,N_8629);
nand U8826 (N_8826,N_8565,N_8553);
and U8827 (N_8827,N_8602,N_8623);
nand U8828 (N_8828,N_8666,N_8552);
xnor U8829 (N_8829,N_8627,N_8705);
or U8830 (N_8830,N_8590,N_8716);
or U8831 (N_8831,N_8628,N_8596);
xnor U8832 (N_8832,N_8720,N_8508);
nand U8833 (N_8833,N_8601,N_8513);
xnor U8834 (N_8834,N_8609,N_8618);
nand U8835 (N_8835,N_8748,N_8714);
nand U8836 (N_8836,N_8599,N_8694);
or U8837 (N_8837,N_8551,N_8520);
xor U8838 (N_8838,N_8625,N_8721);
or U8839 (N_8839,N_8550,N_8645);
xnor U8840 (N_8840,N_8524,N_8749);
nor U8841 (N_8841,N_8593,N_8586);
and U8842 (N_8842,N_8711,N_8719);
or U8843 (N_8843,N_8536,N_8626);
nor U8844 (N_8844,N_8660,N_8697);
nand U8845 (N_8845,N_8537,N_8631);
or U8846 (N_8846,N_8571,N_8554);
nor U8847 (N_8847,N_8582,N_8504);
nand U8848 (N_8848,N_8634,N_8640);
xor U8849 (N_8849,N_8650,N_8739);
xnor U8850 (N_8850,N_8616,N_8577);
nor U8851 (N_8851,N_8532,N_8526);
and U8852 (N_8852,N_8637,N_8738);
xor U8853 (N_8853,N_8555,N_8740);
nand U8854 (N_8854,N_8678,N_8661);
xnor U8855 (N_8855,N_8656,N_8675);
or U8856 (N_8856,N_8726,N_8549);
xnor U8857 (N_8857,N_8692,N_8674);
nand U8858 (N_8858,N_8731,N_8742);
xor U8859 (N_8859,N_8706,N_8671);
or U8860 (N_8860,N_8700,N_8559);
or U8861 (N_8861,N_8527,N_8709);
nand U8862 (N_8862,N_8703,N_8687);
or U8863 (N_8863,N_8677,N_8606);
nor U8864 (N_8864,N_8579,N_8611);
and U8865 (N_8865,N_8688,N_8683);
nand U8866 (N_8866,N_8620,N_8557);
and U8867 (N_8867,N_8725,N_8698);
nor U8868 (N_8868,N_8702,N_8712);
or U8869 (N_8869,N_8651,N_8591);
or U8870 (N_8870,N_8653,N_8699);
nor U8871 (N_8871,N_8746,N_8657);
and U8872 (N_8872,N_8607,N_8736);
nand U8873 (N_8873,N_8501,N_8647);
or U8874 (N_8874,N_8568,N_8511);
and U8875 (N_8875,N_8593,N_8600);
and U8876 (N_8876,N_8545,N_8557);
nand U8877 (N_8877,N_8709,N_8689);
and U8878 (N_8878,N_8574,N_8520);
or U8879 (N_8879,N_8661,N_8602);
nor U8880 (N_8880,N_8619,N_8524);
or U8881 (N_8881,N_8605,N_8548);
xnor U8882 (N_8882,N_8580,N_8662);
and U8883 (N_8883,N_8721,N_8671);
xor U8884 (N_8884,N_8516,N_8623);
nor U8885 (N_8885,N_8703,N_8516);
or U8886 (N_8886,N_8558,N_8734);
or U8887 (N_8887,N_8577,N_8738);
nand U8888 (N_8888,N_8641,N_8517);
nand U8889 (N_8889,N_8725,N_8582);
nand U8890 (N_8890,N_8526,N_8651);
xnor U8891 (N_8891,N_8692,N_8546);
and U8892 (N_8892,N_8567,N_8573);
nand U8893 (N_8893,N_8593,N_8626);
or U8894 (N_8894,N_8611,N_8657);
nor U8895 (N_8895,N_8705,N_8658);
xor U8896 (N_8896,N_8501,N_8634);
or U8897 (N_8897,N_8657,N_8620);
and U8898 (N_8898,N_8581,N_8724);
nand U8899 (N_8899,N_8712,N_8708);
and U8900 (N_8900,N_8679,N_8714);
and U8901 (N_8901,N_8621,N_8741);
and U8902 (N_8902,N_8536,N_8585);
and U8903 (N_8903,N_8574,N_8595);
xnor U8904 (N_8904,N_8737,N_8635);
xnor U8905 (N_8905,N_8724,N_8623);
nor U8906 (N_8906,N_8717,N_8582);
nand U8907 (N_8907,N_8504,N_8587);
and U8908 (N_8908,N_8679,N_8651);
and U8909 (N_8909,N_8672,N_8507);
nor U8910 (N_8910,N_8592,N_8607);
nand U8911 (N_8911,N_8727,N_8736);
nor U8912 (N_8912,N_8597,N_8739);
nor U8913 (N_8913,N_8500,N_8728);
nand U8914 (N_8914,N_8662,N_8592);
xnor U8915 (N_8915,N_8694,N_8528);
nand U8916 (N_8916,N_8647,N_8744);
nand U8917 (N_8917,N_8654,N_8734);
or U8918 (N_8918,N_8671,N_8613);
xor U8919 (N_8919,N_8725,N_8531);
nor U8920 (N_8920,N_8560,N_8681);
nand U8921 (N_8921,N_8646,N_8631);
nand U8922 (N_8922,N_8647,N_8642);
nand U8923 (N_8923,N_8519,N_8704);
xnor U8924 (N_8924,N_8676,N_8578);
nor U8925 (N_8925,N_8659,N_8716);
or U8926 (N_8926,N_8509,N_8556);
xor U8927 (N_8927,N_8725,N_8701);
or U8928 (N_8928,N_8685,N_8708);
nand U8929 (N_8929,N_8708,N_8590);
nand U8930 (N_8930,N_8736,N_8713);
or U8931 (N_8931,N_8518,N_8739);
or U8932 (N_8932,N_8647,N_8609);
nand U8933 (N_8933,N_8703,N_8695);
nor U8934 (N_8934,N_8644,N_8656);
nor U8935 (N_8935,N_8708,N_8743);
nor U8936 (N_8936,N_8579,N_8641);
xnor U8937 (N_8937,N_8645,N_8737);
and U8938 (N_8938,N_8508,N_8627);
xor U8939 (N_8939,N_8671,N_8631);
or U8940 (N_8940,N_8654,N_8636);
nor U8941 (N_8941,N_8519,N_8746);
and U8942 (N_8942,N_8683,N_8749);
nor U8943 (N_8943,N_8745,N_8523);
xnor U8944 (N_8944,N_8618,N_8525);
xnor U8945 (N_8945,N_8631,N_8649);
xor U8946 (N_8946,N_8604,N_8697);
nand U8947 (N_8947,N_8723,N_8595);
nor U8948 (N_8948,N_8680,N_8536);
or U8949 (N_8949,N_8628,N_8517);
xor U8950 (N_8950,N_8643,N_8596);
nor U8951 (N_8951,N_8749,N_8748);
nand U8952 (N_8952,N_8528,N_8613);
nand U8953 (N_8953,N_8652,N_8663);
nor U8954 (N_8954,N_8666,N_8661);
xnor U8955 (N_8955,N_8570,N_8684);
and U8956 (N_8956,N_8566,N_8573);
nor U8957 (N_8957,N_8506,N_8564);
or U8958 (N_8958,N_8574,N_8745);
xnor U8959 (N_8959,N_8736,N_8527);
xor U8960 (N_8960,N_8586,N_8543);
nand U8961 (N_8961,N_8505,N_8578);
or U8962 (N_8962,N_8505,N_8728);
nand U8963 (N_8963,N_8621,N_8505);
xor U8964 (N_8964,N_8584,N_8661);
xor U8965 (N_8965,N_8629,N_8709);
and U8966 (N_8966,N_8746,N_8625);
xnor U8967 (N_8967,N_8698,N_8595);
nor U8968 (N_8968,N_8564,N_8740);
nand U8969 (N_8969,N_8746,N_8681);
and U8970 (N_8970,N_8528,N_8670);
or U8971 (N_8971,N_8664,N_8673);
and U8972 (N_8972,N_8652,N_8634);
and U8973 (N_8973,N_8589,N_8578);
and U8974 (N_8974,N_8576,N_8602);
nor U8975 (N_8975,N_8671,N_8503);
xnor U8976 (N_8976,N_8731,N_8682);
and U8977 (N_8977,N_8540,N_8569);
xnor U8978 (N_8978,N_8648,N_8603);
nand U8979 (N_8979,N_8555,N_8699);
and U8980 (N_8980,N_8702,N_8695);
and U8981 (N_8981,N_8500,N_8567);
or U8982 (N_8982,N_8529,N_8682);
and U8983 (N_8983,N_8705,N_8544);
nor U8984 (N_8984,N_8548,N_8561);
nor U8985 (N_8985,N_8504,N_8609);
and U8986 (N_8986,N_8512,N_8523);
nor U8987 (N_8987,N_8605,N_8551);
nor U8988 (N_8988,N_8688,N_8691);
nor U8989 (N_8989,N_8669,N_8745);
nor U8990 (N_8990,N_8575,N_8719);
nand U8991 (N_8991,N_8654,N_8678);
xnor U8992 (N_8992,N_8654,N_8550);
nor U8993 (N_8993,N_8740,N_8714);
or U8994 (N_8994,N_8592,N_8689);
and U8995 (N_8995,N_8746,N_8626);
xnor U8996 (N_8996,N_8694,N_8548);
nand U8997 (N_8997,N_8585,N_8628);
and U8998 (N_8998,N_8693,N_8587);
nand U8999 (N_8999,N_8668,N_8660);
nor U9000 (N_9000,N_8984,N_8784);
and U9001 (N_9001,N_8862,N_8897);
and U9002 (N_9002,N_8907,N_8750);
nor U9003 (N_9003,N_8911,N_8978);
or U9004 (N_9004,N_8752,N_8900);
nand U9005 (N_9005,N_8792,N_8910);
and U9006 (N_9006,N_8974,N_8780);
xnor U9007 (N_9007,N_8965,N_8990);
nor U9008 (N_9008,N_8946,N_8966);
nor U9009 (N_9009,N_8989,N_8806);
nand U9010 (N_9010,N_8918,N_8759);
and U9011 (N_9011,N_8781,N_8980);
and U9012 (N_9012,N_8985,N_8793);
and U9013 (N_9013,N_8800,N_8765);
xor U9014 (N_9014,N_8901,N_8832);
nand U9015 (N_9015,N_8875,N_8882);
xor U9016 (N_9016,N_8828,N_8856);
or U9017 (N_9017,N_8790,N_8767);
and U9018 (N_9018,N_8973,N_8843);
xnor U9019 (N_9019,N_8887,N_8755);
and U9020 (N_9020,N_8997,N_8820);
and U9021 (N_9021,N_8947,N_8952);
nor U9022 (N_9022,N_8977,N_8787);
and U9023 (N_9023,N_8905,N_8867);
nand U9024 (N_9024,N_8883,N_8925);
nand U9025 (N_9025,N_8857,N_8945);
nor U9026 (N_9026,N_8927,N_8913);
or U9027 (N_9027,N_8836,N_8889);
nor U9028 (N_9028,N_8881,N_8801);
nor U9029 (N_9029,N_8812,N_8786);
xor U9030 (N_9030,N_8877,N_8924);
nor U9031 (N_9031,N_8768,N_8824);
or U9032 (N_9032,N_8931,N_8854);
or U9033 (N_9033,N_8773,N_8930);
xnor U9034 (N_9034,N_8842,N_8860);
and U9035 (N_9035,N_8811,N_8975);
nand U9036 (N_9036,N_8845,N_8833);
nand U9037 (N_9037,N_8822,N_8783);
and U9038 (N_9038,N_8933,N_8823);
xor U9039 (N_9039,N_8782,N_8868);
xnor U9040 (N_9040,N_8953,N_8878);
nand U9041 (N_9041,N_8858,N_8864);
nand U9042 (N_9042,N_8758,N_8915);
or U9043 (N_9043,N_8816,N_8825);
nand U9044 (N_9044,N_8969,N_8892);
nor U9045 (N_9045,N_8950,N_8839);
and U9046 (N_9046,N_8993,N_8899);
xor U9047 (N_9047,N_8754,N_8869);
and U9048 (N_9048,N_8919,N_8834);
xor U9049 (N_9049,N_8796,N_8779);
and U9050 (N_9050,N_8830,N_8971);
or U9051 (N_9051,N_8995,N_8872);
nand U9052 (N_9052,N_8753,N_8770);
nand U9053 (N_9053,N_8943,N_8916);
nor U9054 (N_9054,N_8805,N_8769);
and U9055 (N_9055,N_8976,N_8791);
or U9056 (N_9056,N_8983,N_8934);
nor U9057 (N_9057,N_8936,N_8807);
or U9058 (N_9058,N_8939,N_8988);
and U9059 (N_9059,N_8837,N_8999);
nor U9060 (N_9060,N_8855,N_8859);
nand U9061 (N_9061,N_8844,N_8849);
nand U9062 (N_9062,N_8831,N_8847);
nand U9063 (N_9063,N_8871,N_8917);
or U9064 (N_9064,N_8902,N_8829);
or U9065 (N_9065,N_8895,N_8914);
nand U9066 (N_9066,N_8766,N_8826);
or U9067 (N_9067,N_8891,N_8874);
nand U9068 (N_9068,N_8760,N_8870);
and U9069 (N_9069,N_8850,N_8876);
or U9070 (N_9070,N_8957,N_8951);
nor U9071 (N_9071,N_8838,N_8798);
xnor U9072 (N_9072,N_8873,N_8958);
and U9073 (N_9073,N_8795,N_8851);
xnor U9074 (N_9074,N_8863,N_8762);
xnor U9075 (N_9075,N_8785,N_8763);
nor U9076 (N_9076,N_8813,N_8948);
nand U9077 (N_9077,N_8757,N_8967);
nand U9078 (N_9078,N_8986,N_8802);
or U9079 (N_9079,N_8960,N_8888);
nor U9080 (N_9080,N_8848,N_8810);
xnor U9081 (N_9081,N_8865,N_8809);
or U9082 (N_9082,N_8932,N_8761);
nor U9083 (N_9083,N_8909,N_8774);
nand U9084 (N_9084,N_8776,N_8938);
nand U9085 (N_9085,N_8817,N_8880);
and U9086 (N_9086,N_8808,N_8998);
and U9087 (N_9087,N_8898,N_8789);
nor U9088 (N_9088,N_8852,N_8970);
xnor U9089 (N_9089,N_8968,N_8890);
nand U9090 (N_9090,N_8937,N_8799);
xor U9091 (N_9091,N_8908,N_8949);
nor U9092 (N_9092,N_8987,N_8827);
or U9093 (N_9093,N_8981,N_8835);
or U9094 (N_9094,N_8912,N_8942);
xor U9095 (N_9095,N_8972,N_8804);
and U9096 (N_9096,N_8885,N_8771);
nand U9097 (N_9097,N_8982,N_8803);
nand U9098 (N_9098,N_8788,N_8935);
or U9099 (N_9099,N_8955,N_8959);
nor U9100 (N_9100,N_8879,N_8991);
and U9101 (N_9101,N_8846,N_8814);
nor U9102 (N_9102,N_8819,N_8923);
nand U9103 (N_9103,N_8821,N_8961);
and U9104 (N_9104,N_8896,N_8841);
and U9105 (N_9105,N_8884,N_8956);
or U9106 (N_9106,N_8992,N_8922);
nor U9107 (N_9107,N_8979,N_8940);
nand U9108 (N_9108,N_8772,N_8775);
and U9109 (N_9109,N_8944,N_8962);
and U9110 (N_9110,N_8906,N_8921);
nand U9111 (N_9111,N_8751,N_8866);
xnor U9112 (N_9112,N_8996,N_8954);
and U9113 (N_9113,N_8861,N_8994);
or U9114 (N_9114,N_8777,N_8840);
xnor U9115 (N_9115,N_8894,N_8928);
nand U9116 (N_9116,N_8794,N_8778);
and U9117 (N_9117,N_8853,N_8903);
and U9118 (N_9118,N_8815,N_8764);
or U9119 (N_9119,N_8797,N_8963);
xnor U9120 (N_9120,N_8818,N_8941);
and U9121 (N_9121,N_8886,N_8756);
xor U9122 (N_9122,N_8904,N_8926);
xnor U9123 (N_9123,N_8893,N_8920);
nand U9124 (N_9124,N_8964,N_8929);
and U9125 (N_9125,N_8994,N_8804);
and U9126 (N_9126,N_8783,N_8844);
and U9127 (N_9127,N_8854,N_8903);
or U9128 (N_9128,N_8829,N_8926);
xnor U9129 (N_9129,N_8934,N_8873);
nor U9130 (N_9130,N_8767,N_8807);
nand U9131 (N_9131,N_8769,N_8858);
xnor U9132 (N_9132,N_8822,N_8798);
xnor U9133 (N_9133,N_8964,N_8818);
or U9134 (N_9134,N_8985,N_8867);
nor U9135 (N_9135,N_8867,N_8982);
xor U9136 (N_9136,N_8806,N_8869);
nand U9137 (N_9137,N_8977,N_8795);
xor U9138 (N_9138,N_8975,N_8957);
xnor U9139 (N_9139,N_8902,N_8867);
nor U9140 (N_9140,N_8804,N_8973);
and U9141 (N_9141,N_8870,N_8873);
nor U9142 (N_9142,N_8762,N_8788);
nor U9143 (N_9143,N_8858,N_8750);
or U9144 (N_9144,N_8969,N_8854);
nor U9145 (N_9145,N_8986,N_8960);
nand U9146 (N_9146,N_8916,N_8869);
nand U9147 (N_9147,N_8918,N_8917);
nand U9148 (N_9148,N_8855,N_8998);
or U9149 (N_9149,N_8993,N_8780);
or U9150 (N_9150,N_8867,N_8771);
xnor U9151 (N_9151,N_8920,N_8898);
nor U9152 (N_9152,N_8762,N_8948);
or U9153 (N_9153,N_8833,N_8849);
xnor U9154 (N_9154,N_8884,N_8816);
nor U9155 (N_9155,N_8751,N_8949);
nand U9156 (N_9156,N_8976,N_8788);
xor U9157 (N_9157,N_8935,N_8893);
and U9158 (N_9158,N_8914,N_8857);
nand U9159 (N_9159,N_8924,N_8959);
and U9160 (N_9160,N_8871,N_8854);
nand U9161 (N_9161,N_8982,N_8962);
or U9162 (N_9162,N_8821,N_8933);
nand U9163 (N_9163,N_8931,N_8828);
or U9164 (N_9164,N_8960,N_8957);
nand U9165 (N_9165,N_8957,N_8792);
or U9166 (N_9166,N_8994,N_8972);
xnor U9167 (N_9167,N_8771,N_8996);
nor U9168 (N_9168,N_8815,N_8967);
nand U9169 (N_9169,N_8972,N_8933);
xnor U9170 (N_9170,N_8867,N_8812);
nor U9171 (N_9171,N_8871,N_8940);
xor U9172 (N_9172,N_8938,N_8948);
or U9173 (N_9173,N_8853,N_8828);
nand U9174 (N_9174,N_8909,N_8951);
xor U9175 (N_9175,N_8918,N_8798);
xor U9176 (N_9176,N_8832,N_8993);
or U9177 (N_9177,N_8862,N_8975);
or U9178 (N_9178,N_8825,N_8814);
nand U9179 (N_9179,N_8802,N_8768);
and U9180 (N_9180,N_8998,N_8967);
or U9181 (N_9181,N_8760,N_8912);
and U9182 (N_9182,N_8813,N_8982);
or U9183 (N_9183,N_8783,N_8856);
and U9184 (N_9184,N_8961,N_8764);
and U9185 (N_9185,N_8806,N_8893);
and U9186 (N_9186,N_8773,N_8843);
and U9187 (N_9187,N_8815,N_8969);
or U9188 (N_9188,N_8927,N_8871);
and U9189 (N_9189,N_8838,N_8906);
and U9190 (N_9190,N_8948,N_8808);
nand U9191 (N_9191,N_8761,N_8971);
or U9192 (N_9192,N_8782,N_8816);
nor U9193 (N_9193,N_8858,N_8926);
nor U9194 (N_9194,N_8973,N_8842);
nor U9195 (N_9195,N_8995,N_8796);
and U9196 (N_9196,N_8831,N_8986);
nor U9197 (N_9197,N_8900,N_8964);
nand U9198 (N_9198,N_8952,N_8927);
or U9199 (N_9199,N_8991,N_8844);
nor U9200 (N_9200,N_8968,N_8761);
nand U9201 (N_9201,N_8806,N_8888);
nor U9202 (N_9202,N_8832,N_8905);
nor U9203 (N_9203,N_8756,N_8877);
nor U9204 (N_9204,N_8762,N_8936);
nand U9205 (N_9205,N_8888,N_8962);
xor U9206 (N_9206,N_8801,N_8856);
or U9207 (N_9207,N_8798,N_8759);
nor U9208 (N_9208,N_8797,N_8988);
nand U9209 (N_9209,N_8982,N_8968);
nand U9210 (N_9210,N_8797,N_8885);
xor U9211 (N_9211,N_8824,N_8798);
and U9212 (N_9212,N_8975,N_8781);
or U9213 (N_9213,N_8955,N_8997);
nand U9214 (N_9214,N_8893,N_8967);
and U9215 (N_9215,N_8979,N_8858);
nand U9216 (N_9216,N_8758,N_8769);
or U9217 (N_9217,N_8831,N_8942);
nand U9218 (N_9218,N_8751,N_8946);
or U9219 (N_9219,N_8942,N_8968);
xor U9220 (N_9220,N_8896,N_8903);
nor U9221 (N_9221,N_8899,N_8918);
or U9222 (N_9222,N_8929,N_8799);
xor U9223 (N_9223,N_8952,N_8896);
xor U9224 (N_9224,N_8793,N_8764);
or U9225 (N_9225,N_8777,N_8925);
and U9226 (N_9226,N_8778,N_8796);
nand U9227 (N_9227,N_8917,N_8899);
and U9228 (N_9228,N_8788,N_8872);
nand U9229 (N_9229,N_8941,N_8888);
nand U9230 (N_9230,N_8996,N_8972);
xnor U9231 (N_9231,N_8923,N_8804);
xnor U9232 (N_9232,N_8844,N_8782);
and U9233 (N_9233,N_8906,N_8983);
nor U9234 (N_9234,N_8765,N_8901);
nand U9235 (N_9235,N_8862,N_8875);
or U9236 (N_9236,N_8762,N_8945);
and U9237 (N_9237,N_8825,N_8953);
nand U9238 (N_9238,N_8805,N_8873);
or U9239 (N_9239,N_8815,N_8864);
or U9240 (N_9240,N_8826,N_8858);
or U9241 (N_9241,N_8902,N_8761);
nand U9242 (N_9242,N_8795,N_8894);
and U9243 (N_9243,N_8977,N_8819);
or U9244 (N_9244,N_8987,N_8933);
nand U9245 (N_9245,N_8932,N_8931);
or U9246 (N_9246,N_8768,N_8856);
nand U9247 (N_9247,N_8890,N_8900);
nand U9248 (N_9248,N_8800,N_8805);
and U9249 (N_9249,N_8824,N_8754);
and U9250 (N_9250,N_9164,N_9238);
nand U9251 (N_9251,N_9095,N_9121);
or U9252 (N_9252,N_9142,N_9216);
nand U9253 (N_9253,N_9237,N_9102);
or U9254 (N_9254,N_9171,N_9040);
xor U9255 (N_9255,N_9062,N_9036);
and U9256 (N_9256,N_9103,N_9090);
and U9257 (N_9257,N_9220,N_9014);
or U9258 (N_9258,N_9246,N_9154);
and U9259 (N_9259,N_9181,N_9074);
or U9260 (N_9260,N_9055,N_9041);
and U9261 (N_9261,N_9063,N_9033);
nand U9262 (N_9262,N_9003,N_9155);
nor U9263 (N_9263,N_9110,N_9198);
nor U9264 (N_9264,N_9099,N_9166);
nand U9265 (N_9265,N_9089,N_9059);
or U9266 (N_9266,N_9066,N_9039);
xnor U9267 (N_9267,N_9162,N_9179);
and U9268 (N_9268,N_9168,N_9038);
and U9269 (N_9269,N_9030,N_9128);
or U9270 (N_9270,N_9150,N_9097);
xor U9271 (N_9271,N_9084,N_9035);
nand U9272 (N_9272,N_9115,N_9165);
nand U9273 (N_9273,N_9034,N_9206);
nand U9274 (N_9274,N_9050,N_9088);
nor U9275 (N_9275,N_9138,N_9159);
nand U9276 (N_9276,N_9054,N_9013);
or U9277 (N_9277,N_9113,N_9126);
and U9278 (N_9278,N_9133,N_9208);
and U9279 (N_9279,N_9131,N_9104);
nand U9280 (N_9280,N_9079,N_9184);
xor U9281 (N_9281,N_9200,N_9195);
xor U9282 (N_9282,N_9144,N_9147);
and U9283 (N_9283,N_9057,N_9178);
or U9284 (N_9284,N_9217,N_9002);
or U9285 (N_9285,N_9046,N_9082);
nor U9286 (N_9286,N_9176,N_9191);
nand U9287 (N_9287,N_9085,N_9210);
xnor U9288 (N_9288,N_9174,N_9146);
nor U9289 (N_9289,N_9072,N_9249);
nand U9290 (N_9290,N_9111,N_9228);
and U9291 (N_9291,N_9005,N_9173);
xor U9292 (N_9292,N_9167,N_9242);
and U9293 (N_9293,N_9073,N_9199);
and U9294 (N_9294,N_9248,N_9230);
nand U9295 (N_9295,N_9009,N_9105);
xor U9296 (N_9296,N_9020,N_9053);
nand U9297 (N_9297,N_9027,N_9067);
xnor U9298 (N_9298,N_9145,N_9207);
or U9299 (N_9299,N_9119,N_9170);
nand U9300 (N_9300,N_9172,N_9117);
nand U9301 (N_9301,N_9160,N_9158);
xnor U9302 (N_9302,N_9149,N_9243);
xor U9303 (N_9303,N_9087,N_9045);
or U9304 (N_9304,N_9225,N_9008);
and U9305 (N_9305,N_9136,N_9094);
nand U9306 (N_9306,N_9222,N_9204);
xor U9307 (N_9307,N_9161,N_9051);
nand U9308 (N_9308,N_9049,N_9240);
or U9309 (N_9309,N_9157,N_9213);
or U9310 (N_9310,N_9132,N_9232);
nand U9311 (N_9311,N_9052,N_9007);
xnor U9312 (N_9312,N_9185,N_9018);
nor U9313 (N_9313,N_9188,N_9196);
xnor U9314 (N_9314,N_9148,N_9192);
and U9315 (N_9315,N_9010,N_9015);
nand U9316 (N_9316,N_9071,N_9042);
nor U9317 (N_9317,N_9024,N_9244);
nand U9318 (N_9318,N_9135,N_9233);
nor U9319 (N_9319,N_9109,N_9177);
nor U9320 (N_9320,N_9022,N_9189);
and U9321 (N_9321,N_9224,N_9006);
nand U9322 (N_9322,N_9065,N_9202);
nand U9323 (N_9323,N_9226,N_9236);
nand U9324 (N_9324,N_9026,N_9075);
xnor U9325 (N_9325,N_9182,N_9205);
nand U9326 (N_9326,N_9151,N_9156);
xnor U9327 (N_9327,N_9058,N_9069);
or U9328 (N_9328,N_9078,N_9068);
nand U9329 (N_9329,N_9227,N_9029);
or U9330 (N_9330,N_9193,N_9197);
or U9331 (N_9331,N_9223,N_9234);
or U9332 (N_9332,N_9076,N_9048);
and U9333 (N_9333,N_9194,N_9056);
xor U9334 (N_9334,N_9175,N_9060);
and U9335 (N_9335,N_9219,N_9061);
xor U9336 (N_9336,N_9134,N_9016);
xnor U9337 (N_9337,N_9247,N_9092);
or U9338 (N_9338,N_9209,N_9077);
and U9339 (N_9339,N_9031,N_9187);
and U9340 (N_9340,N_9120,N_9043);
nor U9341 (N_9341,N_9143,N_9153);
nand U9342 (N_9342,N_9239,N_9139);
nand U9343 (N_9343,N_9245,N_9093);
nor U9344 (N_9344,N_9116,N_9186);
nand U9345 (N_9345,N_9130,N_9070);
xor U9346 (N_9346,N_9218,N_9083);
xnor U9347 (N_9347,N_9221,N_9203);
xor U9348 (N_9348,N_9047,N_9037);
and U9349 (N_9349,N_9129,N_9023);
xnor U9350 (N_9350,N_9212,N_9169);
and U9351 (N_9351,N_9235,N_9107);
nand U9352 (N_9352,N_9001,N_9017);
or U9353 (N_9353,N_9137,N_9011);
nor U9354 (N_9354,N_9183,N_9231);
nor U9355 (N_9355,N_9127,N_9163);
or U9356 (N_9356,N_9241,N_9229);
nor U9357 (N_9357,N_9080,N_9112);
nand U9358 (N_9358,N_9096,N_9012);
xnor U9359 (N_9359,N_9098,N_9214);
or U9360 (N_9360,N_9100,N_9125);
nor U9361 (N_9361,N_9152,N_9124);
xor U9362 (N_9362,N_9101,N_9122);
nand U9363 (N_9363,N_9140,N_9025);
nor U9364 (N_9364,N_9086,N_9000);
xnor U9365 (N_9365,N_9201,N_9021);
nand U9366 (N_9366,N_9081,N_9114);
or U9367 (N_9367,N_9019,N_9091);
nor U9368 (N_9368,N_9028,N_9064);
or U9369 (N_9369,N_9141,N_9032);
nor U9370 (N_9370,N_9123,N_9118);
nand U9371 (N_9371,N_9190,N_9004);
nor U9372 (N_9372,N_9106,N_9108);
nor U9373 (N_9373,N_9180,N_9044);
or U9374 (N_9374,N_9211,N_9215);
or U9375 (N_9375,N_9063,N_9138);
and U9376 (N_9376,N_9189,N_9051);
or U9377 (N_9377,N_9102,N_9057);
nand U9378 (N_9378,N_9105,N_9225);
nor U9379 (N_9379,N_9130,N_9082);
nor U9380 (N_9380,N_9110,N_9095);
nor U9381 (N_9381,N_9215,N_9060);
nor U9382 (N_9382,N_9009,N_9043);
nand U9383 (N_9383,N_9243,N_9041);
nand U9384 (N_9384,N_9232,N_9142);
xor U9385 (N_9385,N_9167,N_9067);
xnor U9386 (N_9386,N_9087,N_9012);
xnor U9387 (N_9387,N_9071,N_9053);
nand U9388 (N_9388,N_9182,N_9070);
and U9389 (N_9389,N_9042,N_9082);
nor U9390 (N_9390,N_9226,N_9181);
and U9391 (N_9391,N_9147,N_9158);
xnor U9392 (N_9392,N_9054,N_9092);
xor U9393 (N_9393,N_9056,N_9069);
xnor U9394 (N_9394,N_9174,N_9057);
nand U9395 (N_9395,N_9143,N_9120);
xnor U9396 (N_9396,N_9231,N_9199);
and U9397 (N_9397,N_9148,N_9191);
nand U9398 (N_9398,N_9073,N_9230);
nor U9399 (N_9399,N_9011,N_9027);
or U9400 (N_9400,N_9154,N_9138);
nand U9401 (N_9401,N_9126,N_9159);
and U9402 (N_9402,N_9054,N_9114);
or U9403 (N_9403,N_9039,N_9086);
nand U9404 (N_9404,N_9172,N_9042);
nor U9405 (N_9405,N_9151,N_9170);
or U9406 (N_9406,N_9202,N_9167);
and U9407 (N_9407,N_9065,N_9160);
and U9408 (N_9408,N_9159,N_9136);
xor U9409 (N_9409,N_9120,N_9082);
nand U9410 (N_9410,N_9024,N_9103);
or U9411 (N_9411,N_9017,N_9236);
and U9412 (N_9412,N_9123,N_9241);
xor U9413 (N_9413,N_9195,N_9131);
or U9414 (N_9414,N_9062,N_9248);
nor U9415 (N_9415,N_9160,N_9094);
nor U9416 (N_9416,N_9118,N_9081);
xor U9417 (N_9417,N_9225,N_9218);
and U9418 (N_9418,N_9152,N_9069);
and U9419 (N_9419,N_9184,N_9181);
nand U9420 (N_9420,N_9125,N_9141);
and U9421 (N_9421,N_9247,N_9035);
nand U9422 (N_9422,N_9026,N_9035);
nand U9423 (N_9423,N_9242,N_9150);
nor U9424 (N_9424,N_9168,N_9104);
nand U9425 (N_9425,N_9092,N_9115);
nand U9426 (N_9426,N_9143,N_9176);
and U9427 (N_9427,N_9176,N_9230);
xor U9428 (N_9428,N_9056,N_9215);
xor U9429 (N_9429,N_9080,N_9202);
and U9430 (N_9430,N_9185,N_9056);
nand U9431 (N_9431,N_9193,N_9043);
nand U9432 (N_9432,N_9224,N_9092);
nor U9433 (N_9433,N_9005,N_9211);
or U9434 (N_9434,N_9114,N_9180);
xnor U9435 (N_9435,N_9122,N_9008);
or U9436 (N_9436,N_9174,N_9050);
or U9437 (N_9437,N_9043,N_9001);
nand U9438 (N_9438,N_9167,N_9099);
xor U9439 (N_9439,N_9123,N_9012);
nor U9440 (N_9440,N_9148,N_9037);
or U9441 (N_9441,N_9219,N_9049);
and U9442 (N_9442,N_9027,N_9110);
nand U9443 (N_9443,N_9210,N_9105);
and U9444 (N_9444,N_9109,N_9101);
or U9445 (N_9445,N_9095,N_9080);
nand U9446 (N_9446,N_9142,N_9144);
and U9447 (N_9447,N_9244,N_9110);
xnor U9448 (N_9448,N_9082,N_9246);
and U9449 (N_9449,N_9087,N_9072);
xnor U9450 (N_9450,N_9022,N_9069);
or U9451 (N_9451,N_9055,N_9144);
nor U9452 (N_9452,N_9168,N_9246);
nor U9453 (N_9453,N_9121,N_9080);
xnor U9454 (N_9454,N_9000,N_9157);
nor U9455 (N_9455,N_9230,N_9098);
or U9456 (N_9456,N_9027,N_9025);
and U9457 (N_9457,N_9061,N_9116);
xnor U9458 (N_9458,N_9144,N_9236);
or U9459 (N_9459,N_9022,N_9198);
nor U9460 (N_9460,N_9037,N_9115);
nor U9461 (N_9461,N_9023,N_9192);
and U9462 (N_9462,N_9164,N_9067);
xnor U9463 (N_9463,N_9132,N_9093);
nor U9464 (N_9464,N_9198,N_9164);
nand U9465 (N_9465,N_9147,N_9022);
or U9466 (N_9466,N_9210,N_9078);
or U9467 (N_9467,N_9119,N_9031);
nor U9468 (N_9468,N_9035,N_9242);
nor U9469 (N_9469,N_9028,N_9086);
and U9470 (N_9470,N_9120,N_9155);
nand U9471 (N_9471,N_9203,N_9179);
and U9472 (N_9472,N_9108,N_9005);
or U9473 (N_9473,N_9095,N_9204);
or U9474 (N_9474,N_9008,N_9120);
nand U9475 (N_9475,N_9010,N_9002);
xor U9476 (N_9476,N_9179,N_9224);
or U9477 (N_9477,N_9209,N_9248);
or U9478 (N_9478,N_9107,N_9045);
xnor U9479 (N_9479,N_9062,N_9037);
nand U9480 (N_9480,N_9014,N_9206);
and U9481 (N_9481,N_9171,N_9176);
or U9482 (N_9482,N_9038,N_9011);
nand U9483 (N_9483,N_9131,N_9229);
and U9484 (N_9484,N_9133,N_9201);
nor U9485 (N_9485,N_9174,N_9114);
and U9486 (N_9486,N_9083,N_9150);
nor U9487 (N_9487,N_9219,N_9234);
or U9488 (N_9488,N_9159,N_9113);
or U9489 (N_9489,N_9077,N_9220);
nor U9490 (N_9490,N_9248,N_9065);
and U9491 (N_9491,N_9188,N_9231);
nand U9492 (N_9492,N_9143,N_9011);
or U9493 (N_9493,N_9019,N_9034);
nor U9494 (N_9494,N_9223,N_9066);
xor U9495 (N_9495,N_9105,N_9217);
nand U9496 (N_9496,N_9189,N_9059);
xor U9497 (N_9497,N_9191,N_9071);
xnor U9498 (N_9498,N_9201,N_9017);
or U9499 (N_9499,N_9204,N_9033);
xnor U9500 (N_9500,N_9302,N_9315);
and U9501 (N_9501,N_9377,N_9469);
or U9502 (N_9502,N_9351,N_9486);
nor U9503 (N_9503,N_9250,N_9254);
nand U9504 (N_9504,N_9323,N_9400);
nor U9505 (N_9505,N_9256,N_9482);
xnor U9506 (N_9506,N_9262,N_9496);
or U9507 (N_9507,N_9405,N_9494);
xor U9508 (N_9508,N_9467,N_9415);
nand U9509 (N_9509,N_9450,N_9460);
nor U9510 (N_9510,N_9295,N_9436);
and U9511 (N_9511,N_9454,N_9352);
nand U9512 (N_9512,N_9423,N_9350);
nor U9513 (N_9513,N_9458,N_9392);
or U9514 (N_9514,N_9406,N_9327);
nor U9515 (N_9515,N_9286,N_9252);
and U9516 (N_9516,N_9338,N_9471);
nor U9517 (N_9517,N_9408,N_9331);
or U9518 (N_9518,N_9253,N_9297);
nor U9519 (N_9519,N_9489,N_9288);
or U9520 (N_9520,N_9270,N_9306);
nand U9521 (N_9521,N_9346,N_9407);
nand U9522 (N_9522,N_9485,N_9434);
and U9523 (N_9523,N_9381,N_9470);
and U9524 (N_9524,N_9422,N_9363);
and U9525 (N_9525,N_9308,N_9364);
nor U9526 (N_9526,N_9361,N_9399);
nand U9527 (N_9527,N_9367,N_9280);
nand U9528 (N_9528,N_9292,N_9257);
nor U9529 (N_9529,N_9487,N_9276);
and U9530 (N_9530,N_9445,N_9261);
nor U9531 (N_9531,N_9376,N_9359);
and U9532 (N_9532,N_9424,N_9401);
xnor U9533 (N_9533,N_9437,N_9264);
nor U9534 (N_9534,N_9390,N_9457);
xnor U9535 (N_9535,N_9490,N_9465);
nor U9536 (N_9536,N_9272,N_9274);
xnor U9537 (N_9537,N_9427,N_9289);
and U9538 (N_9538,N_9317,N_9296);
nor U9539 (N_9539,N_9410,N_9355);
or U9540 (N_9540,N_9481,N_9329);
nor U9541 (N_9541,N_9451,N_9301);
xor U9542 (N_9542,N_9340,N_9389);
and U9543 (N_9543,N_9268,N_9371);
or U9544 (N_9544,N_9365,N_9275);
xnor U9545 (N_9545,N_9319,N_9342);
or U9546 (N_9546,N_9335,N_9412);
xor U9547 (N_9547,N_9466,N_9440);
nor U9548 (N_9548,N_9375,N_9391);
nor U9549 (N_9549,N_9337,N_9345);
xor U9550 (N_9550,N_9429,N_9314);
xor U9551 (N_9551,N_9271,N_9368);
or U9552 (N_9552,N_9298,N_9349);
xnor U9553 (N_9553,N_9475,N_9397);
nor U9554 (N_9554,N_9320,N_9366);
nand U9555 (N_9555,N_9476,N_9294);
or U9556 (N_9556,N_9369,N_9461);
and U9557 (N_9557,N_9267,N_9384);
nand U9558 (N_9558,N_9398,N_9318);
nand U9559 (N_9559,N_9348,N_9499);
nand U9560 (N_9560,N_9388,N_9446);
nand U9561 (N_9561,N_9343,N_9484);
nor U9562 (N_9562,N_9326,N_9452);
and U9563 (N_9563,N_9497,N_9324);
nor U9564 (N_9564,N_9263,N_9425);
and U9565 (N_9565,N_9421,N_9431);
nand U9566 (N_9566,N_9339,N_9277);
xor U9567 (N_9567,N_9447,N_9307);
and U9568 (N_9568,N_9341,N_9449);
nand U9569 (N_9569,N_9353,N_9479);
and U9570 (N_9570,N_9443,N_9378);
nand U9571 (N_9571,N_9334,N_9304);
or U9572 (N_9572,N_9394,N_9409);
xor U9573 (N_9573,N_9332,N_9459);
or U9574 (N_9574,N_9333,N_9300);
xnor U9575 (N_9575,N_9258,N_9305);
nand U9576 (N_9576,N_9285,N_9453);
xnor U9577 (N_9577,N_9251,N_9372);
or U9578 (N_9578,N_9311,N_9416);
xor U9579 (N_9579,N_9448,N_9291);
nor U9580 (N_9580,N_9395,N_9266);
xor U9581 (N_9581,N_9385,N_9419);
and U9582 (N_9582,N_9309,N_9473);
nand U9583 (N_9583,N_9498,N_9358);
nand U9584 (N_9584,N_9303,N_9462);
nand U9585 (N_9585,N_9354,N_9483);
nand U9586 (N_9586,N_9370,N_9379);
nor U9587 (N_9587,N_9347,N_9413);
or U9588 (N_9588,N_9330,N_9477);
xor U9589 (N_9589,N_9468,N_9492);
and U9590 (N_9590,N_9310,N_9290);
nor U9591 (N_9591,N_9441,N_9420);
nor U9592 (N_9592,N_9360,N_9491);
xnor U9593 (N_9593,N_9356,N_9278);
nand U9594 (N_9594,N_9322,N_9428);
nand U9595 (N_9595,N_9417,N_9382);
xor U9596 (N_9596,N_9287,N_9488);
nor U9597 (N_9597,N_9373,N_9444);
xor U9598 (N_9598,N_9299,N_9442);
nand U9599 (N_9599,N_9411,N_9312);
xor U9600 (N_9600,N_9336,N_9402);
nor U9601 (N_9601,N_9282,N_9255);
xor U9602 (N_9602,N_9478,N_9493);
or U9603 (N_9603,N_9432,N_9321);
nand U9604 (N_9604,N_9259,N_9273);
and U9605 (N_9605,N_9269,N_9313);
nand U9606 (N_9606,N_9344,N_9279);
nand U9607 (N_9607,N_9430,N_9383);
nand U9608 (N_9608,N_9463,N_9386);
xnor U9609 (N_9609,N_9433,N_9325);
nand U9610 (N_9610,N_9393,N_9380);
nor U9611 (N_9611,N_9404,N_9456);
xnor U9612 (N_9612,N_9374,N_9265);
nand U9613 (N_9613,N_9464,N_9357);
nand U9614 (N_9614,N_9495,N_9455);
nor U9615 (N_9615,N_9426,N_9474);
nor U9616 (N_9616,N_9260,N_9439);
nand U9617 (N_9617,N_9414,N_9293);
xnor U9618 (N_9618,N_9284,N_9362);
or U9619 (N_9619,N_9387,N_9418);
and U9620 (N_9620,N_9480,N_9283);
or U9621 (N_9621,N_9472,N_9328);
nand U9622 (N_9622,N_9281,N_9396);
nor U9623 (N_9623,N_9435,N_9438);
nand U9624 (N_9624,N_9403,N_9316);
and U9625 (N_9625,N_9346,N_9459);
nand U9626 (N_9626,N_9344,N_9498);
or U9627 (N_9627,N_9282,N_9273);
xnor U9628 (N_9628,N_9311,N_9487);
and U9629 (N_9629,N_9452,N_9424);
or U9630 (N_9630,N_9289,N_9356);
nand U9631 (N_9631,N_9294,N_9445);
xor U9632 (N_9632,N_9416,N_9322);
and U9633 (N_9633,N_9400,N_9349);
and U9634 (N_9634,N_9290,N_9473);
nor U9635 (N_9635,N_9490,N_9251);
xor U9636 (N_9636,N_9327,N_9281);
xnor U9637 (N_9637,N_9486,N_9319);
nand U9638 (N_9638,N_9484,N_9331);
nand U9639 (N_9639,N_9482,N_9415);
or U9640 (N_9640,N_9274,N_9414);
nor U9641 (N_9641,N_9369,N_9304);
and U9642 (N_9642,N_9377,N_9381);
and U9643 (N_9643,N_9350,N_9421);
nor U9644 (N_9644,N_9364,N_9279);
nand U9645 (N_9645,N_9498,N_9338);
xor U9646 (N_9646,N_9475,N_9353);
or U9647 (N_9647,N_9479,N_9333);
or U9648 (N_9648,N_9489,N_9278);
nor U9649 (N_9649,N_9261,N_9359);
nor U9650 (N_9650,N_9268,N_9357);
or U9651 (N_9651,N_9458,N_9335);
or U9652 (N_9652,N_9408,N_9301);
or U9653 (N_9653,N_9345,N_9427);
or U9654 (N_9654,N_9398,N_9420);
nand U9655 (N_9655,N_9480,N_9470);
nor U9656 (N_9656,N_9331,N_9416);
or U9657 (N_9657,N_9482,N_9275);
or U9658 (N_9658,N_9263,N_9364);
nand U9659 (N_9659,N_9364,N_9327);
or U9660 (N_9660,N_9363,N_9437);
or U9661 (N_9661,N_9414,N_9372);
and U9662 (N_9662,N_9495,N_9450);
nor U9663 (N_9663,N_9320,N_9471);
or U9664 (N_9664,N_9371,N_9317);
or U9665 (N_9665,N_9470,N_9255);
nand U9666 (N_9666,N_9427,N_9450);
and U9667 (N_9667,N_9319,N_9397);
nand U9668 (N_9668,N_9383,N_9349);
xor U9669 (N_9669,N_9383,N_9474);
and U9670 (N_9670,N_9341,N_9298);
or U9671 (N_9671,N_9275,N_9357);
xnor U9672 (N_9672,N_9445,N_9389);
nand U9673 (N_9673,N_9422,N_9293);
nand U9674 (N_9674,N_9358,N_9378);
xnor U9675 (N_9675,N_9299,N_9318);
or U9676 (N_9676,N_9372,N_9410);
nor U9677 (N_9677,N_9333,N_9348);
or U9678 (N_9678,N_9317,N_9354);
and U9679 (N_9679,N_9383,N_9437);
nand U9680 (N_9680,N_9436,N_9460);
nor U9681 (N_9681,N_9272,N_9335);
xor U9682 (N_9682,N_9338,N_9391);
xor U9683 (N_9683,N_9388,N_9488);
nor U9684 (N_9684,N_9294,N_9376);
and U9685 (N_9685,N_9337,N_9439);
nand U9686 (N_9686,N_9475,N_9318);
or U9687 (N_9687,N_9369,N_9366);
nor U9688 (N_9688,N_9450,N_9468);
nand U9689 (N_9689,N_9356,N_9355);
xnor U9690 (N_9690,N_9288,N_9304);
nand U9691 (N_9691,N_9395,N_9359);
and U9692 (N_9692,N_9383,N_9340);
or U9693 (N_9693,N_9300,N_9400);
nand U9694 (N_9694,N_9333,N_9424);
xnor U9695 (N_9695,N_9279,N_9417);
nand U9696 (N_9696,N_9438,N_9470);
xnor U9697 (N_9697,N_9351,N_9414);
nand U9698 (N_9698,N_9359,N_9416);
and U9699 (N_9699,N_9356,N_9304);
nand U9700 (N_9700,N_9496,N_9374);
nand U9701 (N_9701,N_9281,N_9416);
and U9702 (N_9702,N_9421,N_9427);
nand U9703 (N_9703,N_9466,N_9318);
or U9704 (N_9704,N_9280,N_9314);
and U9705 (N_9705,N_9266,N_9347);
nand U9706 (N_9706,N_9396,N_9251);
and U9707 (N_9707,N_9455,N_9339);
nor U9708 (N_9708,N_9307,N_9260);
nand U9709 (N_9709,N_9361,N_9257);
and U9710 (N_9710,N_9461,N_9305);
nor U9711 (N_9711,N_9285,N_9434);
nor U9712 (N_9712,N_9293,N_9424);
and U9713 (N_9713,N_9374,N_9471);
nor U9714 (N_9714,N_9321,N_9349);
nand U9715 (N_9715,N_9291,N_9304);
nor U9716 (N_9716,N_9412,N_9312);
xnor U9717 (N_9717,N_9290,N_9437);
nor U9718 (N_9718,N_9319,N_9494);
and U9719 (N_9719,N_9319,N_9365);
nand U9720 (N_9720,N_9297,N_9339);
nand U9721 (N_9721,N_9413,N_9462);
and U9722 (N_9722,N_9427,N_9337);
or U9723 (N_9723,N_9322,N_9306);
xnor U9724 (N_9724,N_9287,N_9265);
xor U9725 (N_9725,N_9456,N_9479);
and U9726 (N_9726,N_9437,N_9310);
xnor U9727 (N_9727,N_9348,N_9258);
or U9728 (N_9728,N_9322,N_9457);
nor U9729 (N_9729,N_9495,N_9465);
and U9730 (N_9730,N_9337,N_9357);
nand U9731 (N_9731,N_9412,N_9365);
and U9732 (N_9732,N_9429,N_9330);
nor U9733 (N_9733,N_9399,N_9435);
or U9734 (N_9734,N_9344,N_9473);
or U9735 (N_9735,N_9390,N_9324);
or U9736 (N_9736,N_9341,N_9330);
and U9737 (N_9737,N_9273,N_9431);
xnor U9738 (N_9738,N_9301,N_9386);
xnor U9739 (N_9739,N_9298,N_9432);
nor U9740 (N_9740,N_9311,N_9280);
nand U9741 (N_9741,N_9341,N_9445);
xor U9742 (N_9742,N_9259,N_9355);
nor U9743 (N_9743,N_9384,N_9315);
or U9744 (N_9744,N_9449,N_9452);
or U9745 (N_9745,N_9310,N_9382);
and U9746 (N_9746,N_9392,N_9360);
or U9747 (N_9747,N_9279,N_9255);
nand U9748 (N_9748,N_9478,N_9325);
nor U9749 (N_9749,N_9441,N_9406);
xor U9750 (N_9750,N_9603,N_9616);
and U9751 (N_9751,N_9540,N_9619);
nand U9752 (N_9752,N_9669,N_9517);
xnor U9753 (N_9753,N_9732,N_9601);
nor U9754 (N_9754,N_9743,N_9746);
or U9755 (N_9755,N_9585,N_9519);
nor U9756 (N_9756,N_9509,N_9582);
xnor U9757 (N_9757,N_9648,N_9524);
nor U9758 (N_9758,N_9573,N_9738);
nor U9759 (N_9759,N_9660,N_9566);
or U9760 (N_9760,N_9640,N_9745);
nor U9761 (N_9761,N_9633,N_9578);
or U9762 (N_9762,N_9598,N_9689);
or U9763 (N_9763,N_9708,N_9500);
nor U9764 (N_9764,N_9718,N_9703);
nor U9765 (N_9765,N_9705,N_9602);
nor U9766 (N_9766,N_9664,N_9711);
and U9767 (N_9767,N_9688,N_9674);
nand U9768 (N_9768,N_9695,N_9522);
nand U9769 (N_9769,N_9503,N_9505);
nor U9770 (N_9770,N_9696,N_9572);
xor U9771 (N_9771,N_9506,N_9672);
or U9772 (N_9772,N_9597,N_9610);
xnor U9773 (N_9773,N_9581,N_9733);
nor U9774 (N_9774,N_9704,N_9706);
nand U9775 (N_9775,N_9560,N_9516);
xnor U9776 (N_9776,N_9707,N_9681);
xnor U9777 (N_9777,N_9550,N_9568);
xor U9778 (N_9778,N_9624,N_9694);
or U9779 (N_9779,N_9556,N_9561);
nor U9780 (N_9780,N_9538,N_9700);
and U9781 (N_9781,N_9571,N_9565);
nor U9782 (N_9782,N_9641,N_9722);
nand U9783 (N_9783,N_9562,N_9629);
xor U9784 (N_9784,N_9611,N_9589);
and U9785 (N_9785,N_9595,N_9668);
nand U9786 (N_9786,N_9606,N_9567);
nor U9787 (N_9787,N_9512,N_9510);
xor U9788 (N_9788,N_9584,N_9529);
xnor U9789 (N_9789,N_9592,N_9559);
xnor U9790 (N_9790,N_9740,N_9713);
xnor U9791 (N_9791,N_9587,N_9580);
nand U9792 (N_9792,N_9575,N_9545);
nor U9793 (N_9793,N_9749,N_9638);
xor U9794 (N_9794,N_9627,N_9650);
nand U9795 (N_9795,N_9670,N_9590);
nor U9796 (N_9796,N_9644,N_9715);
or U9797 (N_9797,N_9645,N_9729);
or U9798 (N_9798,N_9662,N_9655);
nor U9799 (N_9799,N_9748,N_9637);
nand U9800 (N_9800,N_9731,N_9551);
xor U9801 (N_9801,N_9532,N_9613);
and U9802 (N_9802,N_9557,N_9667);
nor U9803 (N_9803,N_9631,N_9690);
nand U9804 (N_9804,N_9625,N_9537);
and U9805 (N_9805,N_9628,N_9725);
nand U9806 (N_9806,N_9596,N_9721);
nor U9807 (N_9807,N_9521,N_9594);
or U9808 (N_9808,N_9717,N_9724);
nor U9809 (N_9809,N_9663,N_9739);
nand U9810 (N_9810,N_9563,N_9554);
xnor U9811 (N_9811,N_9723,N_9656);
nor U9812 (N_9812,N_9621,N_9525);
xnor U9813 (N_9813,N_9514,N_9548);
or U9814 (N_9814,N_9747,N_9515);
nand U9815 (N_9815,N_9552,N_9617);
and U9816 (N_9816,N_9586,N_9574);
nand U9817 (N_9817,N_9744,N_9685);
nor U9818 (N_9818,N_9736,N_9697);
or U9819 (N_9819,N_9511,N_9651);
or U9820 (N_9820,N_9683,N_9634);
xnor U9821 (N_9821,N_9675,N_9702);
xnor U9822 (N_9822,N_9530,N_9534);
nor U9823 (N_9823,N_9659,N_9599);
nand U9824 (N_9824,N_9665,N_9543);
or U9825 (N_9825,N_9646,N_9647);
nor U9826 (N_9826,N_9693,N_9553);
xor U9827 (N_9827,N_9501,N_9642);
and U9828 (N_9828,N_9671,N_9654);
and U9829 (N_9829,N_9653,N_9709);
xnor U9830 (N_9830,N_9536,N_9555);
and U9831 (N_9831,N_9679,N_9547);
nand U9832 (N_9832,N_9684,N_9735);
and U9833 (N_9833,N_9504,N_9569);
or U9834 (N_9834,N_9570,N_9701);
and U9835 (N_9835,N_9591,N_9535);
nand U9836 (N_9836,N_9686,N_9608);
nor U9837 (N_9837,N_9636,N_9622);
nand U9838 (N_9838,N_9520,N_9558);
xor U9839 (N_9839,N_9579,N_9712);
xnor U9840 (N_9840,N_9716,N_9691);
nor U9841 (N_9841,N_9523,N_9605);
or U9842 (N_9842,N_9680,N_9742);
and U9843 (N_9843,N_9682,N_9658);
or U9844 (N_9844,N_9614,N_9528);
nand U9845 (N_9845,N_9698,N_9507);
and U9846 (N_9846,N_9615,N_9518);
and U9847 (N_9847,N_9583,N_9657);
and U9848 (N_9848,N_9541,N_9577);
or U9849 (N_9849,N_9728,N_9593);
or U9850 (N_9850,N_9687,N_9720);
xnor U9851 (N_9851,N_9677,N_9531);
nor U9852 (N_9852,N_9730,N_9609);
nand U9853 (N_9853,N_9604,N_9737);
nand U9854 (N_9854,N_9600,N_9533);
nand U9855 (N_9855,N_9666,N_9564);
and U9856 (N_9856,N_9527,N_9741);
and U9857 (N_9857,N_9661,N_9673);
xor U9858 (N_9858,N_9635,N_9643);
xnor U9859 (N_9859,N_9526,N_9630);
nand U9860 (N_9860,N_9549,N_9714);
or U9861 (N_9861,N_9710,N_9639);
nor U9862 (N_9862,N_9652,N_9588);
xnor U9863 (N_9863,N_9678,N_9542);
nor U9864 (N_9864,N_9612,N_9726);
nand U9865 (N_9865,N_9546,N_9623);
nor U9866 (N_9866,N_9626,N_9576);
nand U9867 (N_9867,N_9699,N_9618);
nor U9868 (N_9868,N_9649,N_9692);
nor U9869 (N_9869,N_9502,N_9632);
and U9870 (N_9870,N_9539,N_9719);
nor U9871 (N_9871,N_9676,N_9734);
and U9872 (N_9872,N_9620,N_9607);
nand U9873 (N_9873,N_9727,N_9544);
nor U9874 (N_9874,N_9508,N_9513);
or U9875 (N_9875,N_9673,N_9614);
nand U9876 (N_9876,N_9702,N_9739);
nor U9877 (N_9877,N_9611,N_9627);
xor U9878 (N_9878,N_9637,N_9537);
and U9879 (N_9879,N_9601,N_9675);
nand U9880 (N_9880,N_9685,N_9674);
and U9881 (N_9881,N_9500,N_9601);
nand U9882 (N_9882,N_9730,N_9694);
or U9883 (N_9883,N_9645,N_9590);
and U9884 (N_9884,N_9739,N_9641);
and U9885 (N_9885,N_9639,N_9546);
xor U9886 (N_9886,N_9553,N_9555);
or U9887 (N_9887,N_9521,N_9681);
and U9888 (N_9888,N_9705,N_9736);
nand U9889 (N_9889,N_9574,N_9626);
nor U9890 (N_9890,N_9744,N_9690);
or U9891 (N_9891,N_9525,N_9734);
nor U9892 (N_9892,N_9742,N_9557);
or U9893 (N_9893,N_9697,N_9596);
xor U9894 (N_9894,N_9643,N_9726);
nand U9895 (N_9895,N_9730,N_9636);
nor U9896 (N_9896,N_9704,N_9654);
and U9897 (N_9897,N_9516,N_9562);
and U9898 (N_9898,N_9507,N_9548);
xnor U9899 (N_9899,N_9714,N_9681);
xnor U9900 (N_9900,N_9547,N_9606);
nand U9901 (N_9901,N_9560,N_9538);
xor U9902 (N_9902,N_9743,N_9720);
and U9903 (N_9903,N_9734,N_9509);
xnor U9904 (N_9904,N_9551,N_9682);
xor U9905 (N_9905,N_9748,N_9679);
xnor U9906 (N_9906,N_9726,N_9521);
xnor U9907 (N_9907,N_9587,N_9583);
nor U9908 (N_9908,N_9651,N_9668);
nor U9909 (N_9909,N_9574,N_9593);
nor U9910 (N_9910,N_9559,N_9543);
xnor U9911 (N_9911,N_9592,N_9644);
and U9912 (N_9912,N_9724,N_9626);
nor U9913 (N_9913,N_9535,N_9631);
nor U9914 (N_9914,N_9514,N_9516);
or U9915 (N_9915,N_9706,N_9594);
nand U9916 (N_9916,N_9748,N_9698);
or U9917 (N_9917,N_9685,N_9646);
nor U9918 (N_9918,N_9674,N_9747);
or U9919 (N_9919,N_9717,N_9695);
or U9920 (N_9920,N_9535,N_9506);
or U9921 (N_9921,N_9529,N_9610);
xnor U9922 (N_9922,N_9509,N_9568);
or U9923 (N_9923,N_9589,N_9511);
nand U9924 (N_9924,N_9658,N_9618);
nand U9925 (N_9925,N_9576,N_9596);
and U9926 (N_9926,N_9502,N_9551);
or U9927 (N_9927,N_9538,N_9615);
or U9928 (N_9928,N_9749,N_9570);
nand U9929 (N_9929,N_9674,N_9556);
xor U9930 (N_9930,N_9675,N_9650);
xor U9931 (N_9931,N_9560,N_9537);
nor U9932 (N_9932,N_9547,N_9527);
xor U9933 (N_9933,N_9712,N_9578);
xor U9934 (N_9934,N_9506,N_9521);
nor U9935 (N_9935,N_9640,N_9723);
and U9936 (N_9936,N_9579,N_9683);
or U9937 (N_9937,N_9560,N_9688);
and U9938 (N_9938,N_9729,N_9629);
nor U9939 (N_9939,N_9551,N_9639);
xor U9940 (N_9940,N_9531,N_9641);
nor U9941 (N_9941,N_9663,N_9534);
or U9942 (N_9942,N_9690,N_9548);
nand U9943 (N_9943,N_9623,N_9505);
or U9944 (N_9944,N_9709,N_9681);
xnor U9945 (N_9945,N_9553,N_9716);
or U9946 (N_9946,N_9595,N_9620);
and U9947 (N_9947,N_9676,N_9551);
nand U9948 (N_9948,N_9706,N_9688);
xnor U9949 (N_9949,N_9654,N_9720);
nor U9950 (N_9950,N_9658,N_9720);
nand U9951 (N_9951,N_9718,N_9532);
and U9952 (N_9952,N_9739,N_9565);
nor U9953 (N_9953,N_9691,N_9581);
xor U9954 (N_9954,N_9693,N_9636);
xnor U9955 (N_9955,N_9574,N_9613);
xnor U9956 (N_9956,N_9582,N_9558);
nor U9957 (N_9957,N_9541,N_9709);
or U9958 (N_9958,N_9730,N_9740);
nand U9959 (N_9959,N_9663,N_9610);
nor U9960 (N_9960,N_9626,N_9712);
nand U9961 (N_9961,N_9571,N_9673);
and U9962 (N_9962,N_9706,N_9670);
nand U9963 (N_9963,N_9511,N_9555);
nor U9964 (N_9964,N_9603,N_9529);
xnor U9965 (N_9965,N_9747,N_9602);
nand U9966 (N_9966,N_9503,N_9658);
and U9967 (N_9967,N_9687,N_9645);
nand U9968 (N_9968,N_9658,N_9552);
xnor U9969 (N_9969,N_9584,N_9555);
or U9970 (N_9970,N_9590,N_9587);
or U9971 (N_9971,N_9570,N_9724);
nor U9972 (N_9972,N_9635,N_9730);
and U9973 (N_9973,N_9667,N_9609);
and U9974 (N_9974,N_9522,N_9531);
xnor U9975 (N_9975,N_9694,N_9692);
nand U9976 (N_9976,N_9621,N_9640);
or U9977 (N_9977,N_9601,N_9618);
and U9978 (N_9978,N_9749,N_9717);
nand U9979 (N_9979,N_9701,N_9634);
xor U9980 (N_9980,N_9671,N_9633);
nand U9981 (N_9981,N_9572,N_9536);
and U9982 (N_9982,N_9599,N_9676);
nand U9983 (N_9983,N_9646,N_9724);
nand U9984 (N_9984,N_9513,N_9583);
xnor U9985 (N_9985,N_9511,N_9572);
xnor U9986 (N_9986,N_9664,N_9578);
or U9987 (N_9987,N_9747,N_9591);
or U9988 (N_9988,N_9594,N_9650);
and U9989 (N_9989,N_9550,N_9662);
or U9990 (N_9990,N_9578,N_9579);
and U9991 (N_9991,N_9644,N_9502);
xnor U9992 (N_9992,N_9663,N_9674);
and U9993 (N_9993,N_9611,N_9573);
and U9994 (N_9994,N_9733,N_9613);
xor U9995 (N_9995,N_9529,N_9502);
nand U9996 (N_9996,N_9568,N_9687);
xnor U9997 (N_9997,N_9570,N_9545);
xor U9998 (N_9998,N_9635,N_9674);
or U9999 (N_9999,N_9508,N_9577);
xnor U10000 (N_10000,N_9762,N_9908);
xnor U10001 (N_10001,N_9931,N_9811);
xor U10002 (N_10002,N_9778,N_9873);
or U10003 (N_10003,N_9957,N_9767);
xnor U10004 (N_10004,N_9951,N_9855);
nor U10005 (N_10005,N_9876,N_9964);
or U10006 (N_10006,N_9754,N_9925);
and U10007 (N_10007,N_9832,N_9850);
or U10008 (N_10008,N_9787,N_9766);
xor U10009 (N_10009,N_9985,N_9882);
nand U10010 (N_10010,N_9889,N_9835);
and U10011 (N_10011,N_9904,N_9831);
nor U10012 (N_10012,N_9768,N_9907);
and U10013 (N_10013,N_9948,N_9939);
nand U10014 (N_10014,N_9955,N_9804);
xor U10015 (N_10015,N_9929,N_9937);
or U10016 (N_10016,N_9828,N_9868);
or U10017 (N_10017,N_9847,N_9865);
and U10018 (N_10018,N_9901,N_9842);
nor U10019 (N_10019,N_9848,N_9887);
xnor U10020 (N_10020,N_9986,N_9896);
nand U10021 (N_10021,N_9892,N_9814);
and U10022 (N_10022,N_9914,N_9779);
or U10023 (N_10023,N_9796,N_9859);
nor U10024 (N_10024,N_9755,N_9952);
nor U10025 (N_10025,N_9954,N_9823);
or U10026 (N_10026,N_9756,N_9979);
xor U10027 (N_10027,N_9940,N_9810);
xor U10028 (N_10028,N_9959,N_9906);
xor U10029 (N_10029,N_9813,N_9818);
nor U10030 (N_10030,N_9763,N_9982);
nor U10031 (N_10031,N_9841,N_9820);
xor U10032 (N_10032,N_9911,N_9885);
nand U10033 (N_10033,N_9932,N_9984);
nor U10034 (N_10034,N_9783,N_9830);
or U10035 (N_10035,N_9854,N_9960);
nand U10036 (N_10036,N_9874,N_9785);
nor U10037 (N_10037,N_9843,N_9983);
and U10038 (N_10038,N_9805,N_9998);
nand U10039 (N_10039,N_9794,N_9819);
nor U10040 (N_10040,N_9938,N_9981);
nand U10041 (N_10041,N_9836,N_9870);
or U10042 (N_10042,N_9757,N_9967);
and U10043 (N_10043,N_9872,N_9950);
nand U10044 (N_10044,N_9879,N_9913);
or U10045 (N_10045,N_9944,N_9991);
xnor U10046 (N_10046,N_9788,N_9976);
nor U10047 (N_10047,N_9912,N_9958);
and U10048 (N_10048,N_9797,N_9936);
nor U10049 (N_10049,N_9933,N_9962);
or U10050 (N_10050,N_9884,N_9917);
and U10051 (N_10051,N_9878,N_9845);
nor U10052 (N_10052,N_9922,N_9776);
nor U10053 (N_10053,N_9930,N_9775);
xnor U10054 (N_10054,N_9765,N_9822);
or U10055 (N_10055,N_9934,N_9774);
xnor U10056 (N_10056,N_9849,N_9894);
and U10057 (N_10057,N_9803,N_9942);
nand U10058 (N_10058,N_9992,N_9866);
xnor U10059 (N_10059,N_9903,N_9807);
nor U10060 (N_10060,N_9902,N_9916);
and U10061 (N_10061,N_9996,N_9927);
nand U10062 (N_10062,N_9971,N_9978);
and U10063 (N_10063,N_9900,N_9881);
or U10064 (N_10064,N_9846,N_9946);
xor U10065 (N_10065,N_9844,N_9915);
and U10066 (N_10066,N_9837,N_9863);
and U10067 (N_10067,N_9824,N_9821);
or U10068 (N_10068,N_9840,N_9816);
nor U10069 (N_10069,N_9781,N_9759);
nand U10070 (N_10070,N_9806,N_9851);
and U10071 (N_10071,N_9947,N_9926);
and U10072 (N_10072,N_9888,N_9815);
nand U10073 (N_10073,N_9993,N_9780);
or U10074 (N_10074,N_9980,N_9970);
xnor U10075 (N_10075,N_9969,N_9753);
or U10076 (N_10076,N_9989,N_9793);
nand U10077 (N_10077,N_9994,N_9924);
xnor U10078 (N_10078,N_9829,N_9858);
and U10079 (N_10079,N_9956,N_9790);
nand U10080 (N_10080,N_9860,N_9891);
or U10081 (N_10081,N_9751,N_9875);
xor U10082 (N_10082,N_9784,N_9941);
xnor U10083 (N_10083,N_9909,N_9801);
and U10084 (N_10084,N_9999,N_9867);
or U10085 (N_10085,N_9852,N_9973);
and U10086 (N_10086,N_9990,N_9921);
or U10087 (N_10087,N_9923,N_9883);
nand U10088 (N_10088,N_9817,N_9825);
and U10089 (N_10089,N_9897,N_9995);
nand U10090 (N_10090,N_9965,N_9795);
xnor U10091 (N_10091,N_9802,N_9974);
or U10092 (N_10092,N_9750,N_9880);
xnor U10093 (N_10093,N_9910,N_9792);
xor U10094 (N_10094,N_9943,N_9782);
nor U10095 (N_10095,N_9862,N_9853);
or U10096 (N_10096,N_9786,N_9895);
nand U10097 (N_10097,N_9773,N_9752);
nor U10098 (N_10098,N_9758,N_9791);
and U10099 (N_10099,N_9856,N_9953);
and U10100 (N_10100,N_9949,N_9769);
nor U10101 (N_10101,N_9877,N_9988);
and U10102 (N_10102,N_9833,N_9771);
nor U10103 (N_10103,N_9945,N_9764);
nand U10104 (N_10104,N_9864,N_9772);
and U10105 (N_10105,N_9809,N_9857);
nor U10106 (N_10106,N_9770,N_9918);
nand U10107 (N_10107,N_9905,N_9920);
nor U10108 (N_10108,N_9760,N_9838);
nor U10109 (N_10109,N_9961,N_9977);
and U10110 (N_10110,N_9972,N_9834);
and U10111 (N_10111,N_9827,N_9997);
xor U10112 (N_10112,N_9826,N_9800);
xnor U10113 (N_10113,N_9886,N_9869);
nor U10114 (N_10114,N_9761,N_9935);
nand U10115 (N_10115,N_9893,N_9871);
nor U10116 (N_10116,N_9899,N_9808);
nor U10117 (N_10117,N_9839,N_9928);
nand U10118 (N_10118,N_9798,N_9968);
nor U10119 (N_10119,N_9777,N_9987);
or U10120 (N_10120,N_9975,N_9966);
xor U10121 (N_10121,N_9890,N_9789);
nand U10122 (N_10122,N_9963,N_9812);
nor U10123 (N_10123,N_9799,N_9919);
xor U10124 (N_10124,N_9898,N_9861);
nand U10125 (N_10125,N_9909,N_9887);
nor U10126 (N_10126,N_9900,N_9996);
xor U10127 (N_10127,N_9953,N_9798);
nand U10128 (N_10128,N_9938,N_9971);
xor U10129 (N_10129,N_9923,N_9986);
nor U10130 (N_10130,N_9793,N_9960);
xor U10131 (N_10131,N_9885,N_9759);
nand U10132 (N_10132,N_9920,N_9993);
xnor U10133 (N_10133,N_9839,N_9929);
xor U10134 (N_10134,N_9826,N_9955);
nand U10135 (N_10135,N_9956,N_9861);
or U10136 (N_10136,N_9868,N_9917);
nor U10137 (N_10137,N_9772,N_9852);
or U10138 (N_10138,N_9931,N_9915);
or U10139 (N_10139,N_9966,N_9751);
or U10140 (N_10140,N_9959,N_9789);
and U10141 (N_10141,N_9859,N_9917);
nor U10142 (N_10142,N_9830,N_9771);
nor U10143 (N_10143,N_9989,N_9817);
or U10144 (N_10144,N_9895,N_9966);
and U10145 (N_10145,N_9894,N_9966);
nand U10146 (N_10146,N_9915,N_9930);
nor U10147 (N_10147,N_9802,N_9933);
nand U10148 (N_10148,N_9888,N_9774);
and U10149 (N_10149,N_9879,N_9803);
nand U10150 (N_10150,N_9860,N_9963);
and U10151 (N_10151,N_9753,N_9953);
nor U10152 (N_10152,N_9979,N_9906);
and U10153 (N_10153,N_9982,N_9953);
and U10154 (N_10154,N_9920,N_9848);
xor U10155 (N_10155,N_9813,N_9795);
nor U10156 (N_10156,N_9817,N_9782);
and U10157 (N_10157,N_9981,N_9801);
and U10158 (N_10158,N_9923,N_9800);
nand U10159 (N_10159,N_9917,N_9768);
xnor U10160 (N_10160,N_9933,N_9839);
and U10161 (N_10161,N_9939,N_9989);
xor U10162 (N_10162,N_9779,N_9896);
nand U10163 (N_10163,N_9833,N_9960);
xnor U10164 (N_10164,N_9857,N_9960);
or U10165 (N_10165,N_9917,N_9830);
and U10166 (N_10166,N_9906,N_9901);
and U10167 (N_10167,N_9861,N_9851);
or U10168 (N_10168,N_9961,N_9975);
nor U10169 (N_10169,N_9961,N_9786);
xnor U10170 (N_10170,N_9850,N_9826);
or U10171 (N_10171,N_9949,N_9788);
or U10172 (N_10172,N_9967,N_9868);
nand U10173 (N_10173,N_9838,N_9871);
nor U10174 (N_10174,N_9998,N_9972);
or U10175 (N_10175,N_9854,N_9912);
xor U10176 (N_10176,N_9948,N_9929);
nor U10177 (N_10177,N_9877,N_9847);
or U10178 (N_10178,N_9873,N_9989);
nor U10179 (N_10179,N_9794,N_9896);
nand U10180 (N_10180,N_9915,N_9810);
nand U10181 (N_10181,N_9918,N_9841);
or U10182 (N_10182,N_9932,N_9998);
or U10183 (N_10183,N_9798,N_9991);
nand U10184 (N_10184,N_9764,N_9883);
nor U10185 (N_10185,N_9977,N_9905);
and U10186 (N_10186,N_9791,N_9946);
nand U10187 (N_10187,N_9834,N_9987);
and U10188 (N_10188,N_9954,N_9784);
nor U10189 (N_10189,N_9895,N_9986);
nor U10190 (N_10190,N_9797,N_9894);
or U10191 (N_10191,N_9770,N_9867);
nand U10192 (N_10192,N_9855,N_9961);
nand U10193 (N_10193,N_9846,N_9879);
or U10194 (N_10194,N_9798,N_9799);
nand U10195 (N_10195,N_9809,N_9910);
xor U10196 (N_10196,N_9959,N_9771);
nand U10197 (N_10197,N_9750,N_9951);
nand U10198 (N_10198,N_9998,N_9901);
or U10199 (N_10199,N_9961,N_9831);
or U10200 (N_10200,N_9936,N_9935);
nor U10201 (N_10201,N_9847,N_9776);
and U10202 (N_10202,N_9939,N_9950);
or U10203 (N_10203,N_9833,N_9826);
nor U10204 (N_10204,N_9847,N_9828);
or U10205 (N_10205,N_9980,N_9924);
and U10206 (N_10206,N_9814,N_9965);
or U10207 (N_10207,N_9939,N_9971);
nand U10208 (N_10208,N_9793,N_9841);
nand U10209 (N_10209,N_9819,N_9778);
nor U10210 (N_10210,N_9898,N_9987);
xnor U10211 (N_10211,N_9807,N_9942);
nor U10212 (N_10212,N_9995,N_9994);
and U10213 (N_10213,N_9798,N_9823);
or U10214 (N_10214,N_9893,N_9892);
xnor U10215 (N_10215,N_9873,N_9840);
nor U10216 (N_10216,N_9756,N_9856);
xor U10217 (N_10217,N_9801,N_9830);
xnor U10218 (N_10218,N_9945,N_9882);
nor U10219 (N_10219,N_9971,N_9983);
nor U10220 (N_10220,N_9823,N_9895);
xnor U10221 (N_10221,N_9823,N_9820);
and U10222 (N_10222,N_9754,N_9955);
and U10223 (N_10223,N_9938,N_9801);
xnor U10224 (N_10224,N_9921,N_9783);
nor U10225 (N_10225,N_9937,N_9861);
xor U10226 (N_10226,N_9856,N_9813);
nand U10227 (N_10227,N_9934,N_9832);
nor U10228 (N_10228,N_9761,N_9859);
nor U10229 (N_10229,N_9988,N_9890);
and U10230 (N_10230,N_9986,N_9921);
or U10231 (N_10231,N_9935,N_9782);
xor U10232 (N_10232,N_9853,N_9761);
and U10233 (N_10233,N_9980,N_9793);
nand U10234 (N_10234,N_9966,N_9977);
or U10235 (N_10235,N_9808,N_9760);
nor U10236 (N_10236,N_9977,N_9893);
nor U10237 (N_10237,N_9910,N_9922);
xor U10238 (N_10238,N_9933,N_9815);
nand U10239 (N_10239,N_9756,N_9880);
nand U10240 (N_10240,N_9857,N_9800);
nor U10241 (N_10241,N_9830,N_9752);
nand U10242 (N_10242,N_9785,N_9782);
nor U10243 (N_10243,N_9821,N_9872);
nor U10244 (N_10244,N_9953,N_9824);
nand U10245 (N_10245,N_9997,N_9905);
nor U10246 (N_10246,N_9985,N_9824);
and U10247 (N_10247,N_9840,N_9804);
or U10248 (N_10248,N_9939,N_9785);
nor U10249 (N_10249,N_9846,N_9894);
and U10250 (N_10250,N_10184,N_10080);
nor U10251 (N_10251,N_10144,N_10194);
nand U10252 (N_10252,N_10173,N_10009);
nand U10253 (N_10253,N_10198,N_10070);
and U10254 (N_10254,N_10245,N_10005);
nor U10255 (N_10255,N_10044,N_10149);
xnor U10256 (N_10256,N_10189,N_10195);
or U10257 (N_10257,N_10153,N_10137);
or U10258 (N_10258,N_10180,N_10082);
nor U10259 (N_10259,N_10102,N_10056);
or U10260 (N_10260,N_10246,N_10227);
nor U10261 (N_10261,N_10028,N_10064);
and U10262 (N_10262,N_10143,N_10096);
and U10263 (N_10263,N_10230,N_10172);
and U10264 (N_10264,N_10065,N_10190);
nand U10265 (N_10265,N_10163,N_10222);
or U10266 (N_10266,N_10016,N_10213);
nand U10267 (N_10267,N_10147,N_10103);
and U10268 (N_10268,N_10117,N_10032);
nor U10269 (N_10269,N_10212,N_10226);
and U10270 (N_10270,N_10146,N_10128);
nand U10271 (N_10271,N_10175,N_10017);
xor U10272 (N_10272,N_10012,N_10097);
and U10273 (N_10273,N_10066,N_10238);
nor U10274 (N_10274,N_10109,N_10191);
and U10275 (N_10275,N_10186,N_10068);
or U10276 (N_10276,N_10014,N_10131);
nand U10277 (N_10277,N_10161,N_10036);
or U10278 (N_10278,N_10239,N_10072);
nand U10279 (N_10279,N_10202,N_10225);
xnor U10280 (N_10280,N_10214,N_10145);
nand U10281 (N_10281,N_10063,N_10140);
nor U10282 (N_10282,N_10092,N_10188);
and U10283 (N_10283,N_10248,N_10001);
or U10284 (N_10284,N_10129,N_10156);
or U10285 (N_10285,N_10174,N_10023);
or U10286 (N_10286,N_10240,N_10168);
or U10287 (N_10287,N_10133,N_10077);
and U10288 (N_10288,N_10229,N_10224);
nor U10289 (N_10289,N_10209,N_10197);
nand U10290 (N_10290,N_10166,N_10039);
nand U10291 (N_10291,N_10236,N_10125);
xnor U10292 (N_10292,N_10199,N_10217);
nand U10293 (N_10293,N_10169,N_10167);
nand U10294 (N_10294,N_10182,N_10019);
or U10295 (N_10295,N_10081,N_10094);
and U10296 (N_10296,N_10207,N_10051);
and U10297 (N_10297,N_10142,N_10004);
or U10298 (N_10298,N_10078,N_10135);
or U10299 (N_10299,N_10013,N_10008);
nand U10300 (N_10300,N_10216,N_10221);
xnor U10301 (N_10301,N_10151,N_10218);
or U10302 (N_10302,N_10057,N_10244);
and U10303 (N_10303,N_10046,N_10231);
nand U10304 (N_10304,N_10134,N_10114);
xnor U10305 (N_10305,N_10215,N_10148);
or U10306 (N_10306,N_10090,N_10141);
xnor U10307 (N_10307,N_10124,N_10024);
or U10308 (N_10308,N_10034,N_10223);
xor U10309 (N_10309,N_10108,N_10037);
xor U10310 (N_10310,N_10206,N_10185);
nand U10311 (N_10311,N_10073,N_10157);
or U10312 (N_10312,N_10091,N_10062);
nor U10313 (N_10313,N_10021,N_10043);
and U10314 (N_10314,N_10000,N_10093);
xor U10315 (N_10315,N_10241,N_10079);
and U10316 (N_10316,N_10177,N_10119);
and U10317 (N_10317,N_10113,N_10232);
nor U10318 (N_10318,N_10127,N_10165);
nand U10319 (N_10319,N_10130,N_10006);
nand U10320 (N_10320,N_10035,N_10058);
or U10321 (N_10321,N_10041,N_10192);
nand U10322 (N_10322,N_10203,N_10042);
nor U10323 (N_10323,N_10181,N_10170);
nand U10324 (N_10324,N_10155,N_10158);
nand U10325 (N_10325,N_10183,N_10139);
and U10326 (N_10326,N_10187,N_10200);
nor U10327 (N_10327,N_10122,N_10045);
and U10328 (N_10328,N_10069,N_10228);
and U10329 (N_10329,N_10115,N_10107);
xor U10330 (N_10330,N_10049,N_10136);
nor U10331 (N_10331,N_10022,N_10138);
or U10332 (N_10332,N_10054,N_10061);
and U10333 (N_10333,N_10018,N_10249);
nor U10334 (N_10334,N_10003,N_10031);
and U10335 (N_10335,N_10193,N_10110);
nor U10336 (N_10336,N_10060,N_10152);
nor U10337 (N_10337,N_10204,N_10120);
or U10338 (N_10338,N_10086,N_10087);
nand U10339 (N_10339,N_10020,N_10038);
nor U10340 (N_10340,N_10116,N_10029);
nor U10341 (N_10341,N_10075,N_10076);
xor U10342 (N_10342,N_10112,N_10105);
and U10343 (N_10343,N_10040,N_10201);
xor U10344 (N_10344,N_10067,N_10111);
xnor U10345 (N_10345,N_10196,N_10098);
xnor U10346 (N_10346,N_10007,N_10088);
nand U10347 (N_10347,N_10208,N_10101);
or U10348 (N_10348,N_10074,N_10234);
nor U10349 (N_10349,N_10084,N_10176);
nand U10350 (N_10350,N_10164,N_10150);
xnor U10351 (N_10351,N_10154,N_10015);
and U10352 (N_10352,N_10052,N_10053);
xor U10353 (N_10353,N_10159,N_10100);
nand U10354 (N_10354,N_10050,N_10048);
nor U10355 (N_10355,N_10099,N_10121);
nand U10356 (N_10356,N_10055,N_10162);
and U10357 (N_10357,N_10089,N_10027);
nor U10358 (N_10358,N_10132,N_10205);
or U10359 (N_10359,N_10219,N_10010);
and U10360 (N_10360,N_10025,N_10247);
and U10361 (N_10361,N_10243,N_10104);
nor U10362 (N_10362,N_10047,N_10033);
or U10363 (N_10363,N_10083,N_10095);
xnor U10364 (N_10364,N_10235,N_10106);
nor U10365 (N_10365,N_10123,N_10059);
xor U10366 (N_10366,N_10126,N_10118);
nand U10367 (N_10367,N_10211,N_10233);
nand U10368 (N_10368,N_10242,N_10179);
and U10369 (N_10369,N_10171,N_10071);
xor U10370 (N_10370,N_10026,N_10178);
and U10371 (N_10371,N_10011,N_10160);
nand U10372 (N_10372,N_10002,N_10210);
xnor U10373 (N_10373,N_10237,N_10220);
xor U10374 (N_10374,N_10085,N_10030);
nand U10375 (N_10375,N_10148,N_10086);
and U10376 (N_10376,N_10215,N_10183);
nand U10377 (N_10377,N_10093,N_10076);
nor U10378 (N_10378,N_10189,N_10017);
or U10379 (N_10379,N_10194,N_10249);
nor U10380 (N_10380,N_10078,N_10070);
or U10381 (N_10381,N_10142,N_10195);
xor U10382 (N_10382,N_10007,N_10076);
or U10383 (N_10383,N_10134,N_10104);
nor U10384 (N_10384,N_10061,N_10224);
or U10385 (N_10385,N_10086,N_10154);
nor U10386 (N_10386,N_10063,N_10237);
and U10387 (N_10387,N_10027,N_10022);
nand U10388 (N_10388,N_10007,N_10175);
nor U10389 (N_10389,N_10177,N_10165);
and U10390 (N_10390,N_10094,N_10107);
and U10391 (N_10391,N_10124,N_10249);
or U10392 (N_10392,N_10184,N_10113);
or U10393 (N_10393,N_10049,N_10111);
nand U10394 (N_10394,N_10184,N_10153);
or U10395 (N_10395,N_10091,N_10051);
and U10396 (N_10396,N_10117,N_10005);
nand U10397 (N_10397,N_10188,N_10082);
xor U10398 (N_10398,N_10037,N_10015);
xor U10399 (N_10399,N_10205,N_10047);
or U10400 (N_10400,N_10132,N_10037);
xor U10401 (N_10401,N_10188,N_10208);
or U10402 (N_10402,N_10023,N_10105);
nand U10403 (N_10403,N_10150,N_10111);
and U10404 (N_10404,N_10126,N_10210);
nor U10405 (N_10405,N_10222,N_10156);
xnor U10406 (N_10406,N_10055,N_10056);
and U10407 (N_10407,N_10168,N_10176);
nor U10408 (N_10408,N_10172,N_10126);
nor U10409 (N_10409,N_10170,N_10098);
or U10410 (N_10410,N_10070,N_10159);
xnor U10411 (N_10411,N_10214,N_10144);
nand U10412 (N_10412,N_10055,N_10027);
and U10413 (N_10413,N_10083,N_10055);
nor U10414 (N_10414,N_10067,N_10021);
or U10415 (N_10415,N_10018,N_10006);
and U10416 (N_10416,N_10037,N_10225);
or U10417 (N_10417,N_10141,N_10155);
and U10418 (N_10418,N_10125,N_10247);
nor U10419 (N_10419,N_10003,N_10083);
nor U10420 (N_10420,N_10239,N_10026);
or U10421 (N_10421,N_10032,N_10245);
or U10422 (N_10422,N_10221,N_10101);
and U10423 (N_10423,N_10189,N_10034);
and U10424 (N_10424,N_10079,N_10247);
nor U10425 (N_10425,N_10031,N_10036);
xnor U10426 (N_10426,N_10088,N_10123);
nand U10427 (N_10427,N_10218,N_10163);
and U10428 (N_10428,N_10003,N_10135);
xor U10429 (N_10429,N_10055,N_10206);
nand U10430 (N_10430,N_10123,N_10094);
or U10431 (N_10431,N_10054,N_10183);
nor U10432 (N_10432,N_10208,N_10112);
and U10433 (N_10433,N_10179,N_10201);
xnor U10434 (N_10434,N_10157,N_10054);
nor U10435 (N_10435,N_10138,N_10197);
nand U10436 (N_10436,N_10064,N_10194);
or U10437 (N_10437,N_10062,N_10152);
or U10438 (N_10438,N_10103,N_10030);
xor U10439 (N_10439,N_10121,N_10006);
nor U10440 (N_10440,N_10145,N_10135);
and U10441 (N_10441,N_10054,N_10242);
nor U10442 (N_10442,N_10226,N_10063);
nor U10443 (N_10443,N_10068,N_10160);
and U10444 (N_10444,N_10172,N_10224);
nor U10445 (N_10445,N_10174,N_10225);
nand U10446 (N_10446,N_10067,N_10048);
nor U10447 (N_10447,N_10009,N_10069);
xor U10448 (N_10448,N_10155,N_10016);
nor U10449 (N_10449,N_10240,N_10020);
nand U10450 (N_10450,N_10023,N_10159);
xor U10451 (N_10451,N_10206,N_10021);
and U10452 (N_10452,N_10067,N_10238);
or U10453 (N_10453,N_10036,N_10094);
xor U10454 (N_10454,N_10075,N_10176);
nor U10455 (N_10455,N_10061,N_10180);
or U10456 (N_10456,N_10197,N_10038);
nand U10457 (N_10457,N_10049,N_10121);
or U10458 (N_10458,N_10229,N_10101);
xnor U10459 (N_10459,N_10017,N_10211);
nor U10460 (N_10460,N_10062,N_10164);
xnor U10461 (N_10461,N_10104,N_10128);
nand U10462 (N_10462,N_10223,N_10109);
and U10463 (N_10463,N_10141,N_10087);
or U10464 (N_10464,N_10018,N_10098);
and U10465 (N_10465,N_10027,N_10212);
or U10466 (N_10466,N_10121,N_10066);
xnor U10467 (N_10467,N_10077,N_10002);
and U10468 (N_10468,N_10147,N_10143);
nand U10469 (N_10469,N_10169,N_10116);
xor U10470 (N_10470,N_10121,N_10171);
or U10471 (N_10471,N_10195,N_10058);
and U10472 (N_10472,N_10071,N_10018);
and U10473 (N_10473,N_10059,N_10109);
and U10474 (N_10474,N_10063,N_10248);
or U10475 (N_10475,N_10199,N_10206);
and U10476 (N_10476,N_10209,N_10092);
nor U10477 (N_10477,N_10184,N_10055);
nand U10478 (N_10478,N_10156,N_10002);
nor U10479 (N_10479,N_10177,N_10179);
nor U10480 (N_10480,N_10117,N_10081);
nor U10481 (N_10481,N_10054,N_10079);
and U10482 (N_10482,N_10202,N_10106);
xor U10483 (N_10483,N_10211,N_10098);
and U10484 (N_10484,N_10041,N_10132);
or U10485 (N_10485,N_10172,N_10144);
or U10486 (N_10486,N_10188,N_10145);
nand U10487 (N_10487,N_10074,N_10039);
nand U10488 (N_10488,N_10066,N_10164);
nor U10489 (N_10489,N_10041,N_10115);
nand U10490 (N_10490,N_10202,N_10072);
and U10491 (N_10491,N_10247,N_10120);
nand U10492 (N_10492,N_10114,N_10216);
xor U10493 (N_10493,N_10014,N_10240);
nand U10494 (N_10494,N_10035,N_10071);
xnor U10495 (N_10495,N_10216,N_10200);
and U10496 (N_10496,N_10240,N_10169);
nor U10497 (N_10497,N_10198,N_10161);
or U10498 (N_10498,N_10082,N_10177);
and U10499 (N_10499,N_10204,N_10028);
nand U10500 (N_10500,N_10431,N_10270);
xor U10501 (N_10501,N_10322,N_10430);
or U10502 (N_10502,N_10301,N_10439);
nand U10503 (N_10503,N_10398,N_10260);
nand U10504 (N_10504,N_10469,N_10420);
nor U10505 (N_10505,N_10458,N_10449);
or U10506 (N_10506,N_10372,N_10323);
nor U10507 (N_10507,N_10298,N_10484);
xnor U10508 (N_10508,N_10394,N_10489);
nor U10509 (N_10509,N_10391,N_10411);
nor U10510 (N_10510,N_10286,N_10274);
xor U10511 (N_10511,N_10284,N_10360);
xnor U10512 (N_10512,N_10253,N_10349);
xnor U10513 (N_10513,N_10328,N_10313);
nor U10514 (N_10514,N_10272,N_10319);
nand U10515 (N_10515,N_10318,N_10281);
nor U10516 (N_10516,N_10412,N_10424);
and U10517 (N_10517,N_10289,N_10258);
or U10518 (N_10518,N_10354,N_10340);
xnor U10519 (N_10519,N_10355,N_10392);
nand U10520 (N_10520,N_10396,N_10265);
and U10521 (N_10521,N_10475,N_10345);
nor U10522 (N_10522,N_10423,N_10324);
nand U10523 (N_10523,N_10380,N_10481);
or U10524 (N_10524,N_10436,N_10418);
xor U10525 (N_10525,N_10432,N_10419);
nor U10526 (N_10526,N_10496,N_10462);
nand U10527 (N_10527,N_10337,N_10421);
xor U10528 (N_10528,N_10405,N_10454);
or U10529 (N_10529,N_10485,N_10402);
nor U10530 (N_10530,N_10478,N_10305);
or U10531 (N_10531,N_10275,N_10288);
nor U10532 (N_10532,N_10291,N_10387);
nor U10533 (N_10533,N_10314,N_10262);
xnor U10534 (N_10534,N_10498,N_10366);
xor U10535 (N_10535,N_10342,N_10304);
xor U10536 (N_10536,N_10447,N_10339);
nand U10537 (N_10537,N_10351,N_10254);
xnor U10538 (N_10538,N_10369,N_10297);
and U10539 (N_10539,N_10317,N_10331);
nor U10540 (N_10540,N_10327,N_10480);
xnor U10541 (N_10541,N_10473,N_10279);
nand U10542 (N_10542,N_10310,N_10385);
nor U10543 (N_10543,N_10311,N_10470);
nand U10544 (N_10544,N_10467,N_10371);
or U10545 (N_10545,N_10368,N_10290);
and U10546 (N_10546,N_10472,N_10381);
xnor U10547 (N_10547,N_10388,N_10476);
xor U10548 (N_10548,N_10451,N_10296);
and U10549 (N_10549,N_10433,N_10408);
and U10550 (N_10550,N_10383,N_10400);
xor U10551 (N_10551,N_10403,N_10378);
or U10552 (N_10552,N_10488,N_10440);
or U10553 (N_10553,N_10429,N_10344);
xor U10554 (N_10554,N_10268,N_10350);
and U10555 (N_10555,N_10259,N_10346);
nor U10556 (N_10556,N_10477,N_10307);
nand U10557 (N_10557,N_10329,N_10266);
xnor U10558 (N_10558,N_10401,N_10308);
and U10559 (N_10559,N_10428,N_10468);
and U10560 (N_10560,N_10263,N_10490);
or U10561 (N_10561,N_10374,N_10409);
and U10562 (N_10562,N_10399,N_10395);
and U10563 (N_10563,N_10267,N_10493);
xor U10564 (N_10564,N_10413,N_10356);
nand U10565 (N_10565,N_10358,N_10278);
or U10566 (N_10566,N_10309,N_10334);
nand U10567 (N_10567,N_10287,N_10359);
or U10568 (N_10568,N_10257,N_10406);
nand U10569 (N_10569,N_10416,N_10251);
nor U10570 (N_10570,N_10495,N_10415);
nor U10571 (N_10571,N_10295,N_10492);
and U10572 (N_10572,N_10370,N_10497);
xor U10573 (N_10573,N_10277,N_10269);
xor U10574 (N_10574,N_10474,N_10250);
or U10575 (N_10575,N_10273,N_10362);
and U10576 (N_10576,N_10414,N_10283);
and U10577 (N_10577,N_10361,N_10325);
and U10578 (N_10578,N_10443,N_10384);
nand U10579 (N_10579,N_10292,N_10382);
xor U10580 (N_10580,N_10410,N_10446);
nor U10581 (N_10581,N_10255,N_10459);
and U10582 (N_10582,N_10457,N_10336);
nor U10583 (N_10583,N_10312,N_10452);
and U10584 (N_10584,N_10343,N_10352);
nor U10585 (N_10585,N_10445,N_10326);
and U10586 (N_10586,N_10364,N_10363);
nor U10587 (N_10587,N_10455,N_10365);
nor U10588 (N_10588,N_10422,N_10464);
nor U10589 (N_10589,N_10453,N_10456);
or U10590 (N_10590,N_10303,N_10448);
nand U10591 (N_10591,N_10315,N_10494);
nor U10592 (N_10592,N_10407,N_10425);
xnor U10593 (N_10593,N_10377,N_10330);
nand U10594 (N_10594,N_10379,N_10357);
nand U10595 (N_10595,N_10280,N_10487);
xnor U10596 (N_10596,N_10499,N_10461);
nor U10597 (N_10597,N_10483,N_10276);
nor U10598 (N_10598,N_10300,N_10367);
xnor U10599 (N_10599,N_10426,N_10335);
nor U10600 (N_10600,N_10390,N_10332);
nand U10601 (N_10601,N_10338,N_10321);
or U10602 (N_10602,N_10376,N_10282);
xnor U10603 (N_10603,N_10466,N_10450);
xor U10604 (N_10604,N_10438,N_10482);
nor U10605 (N_10605,N_10348,N_10306);
nor U10606 (N_10606,N_10299,N_10271);
or U10607 (N_10607,N_10404,N_10316);
nand U10608 (N_10608,N_10293,N_10471);
and U10609 (N_10609,N_10435,N_10373);
and U10610 (N_10610,N_10353,N_10463);
xor U10611 (N_10611,N_10434,N_10389);
and U10612 (N_10612,N_10486,N_10444);
nor U10613 (N_10613,N_10264,N_10375);
and U10614 (N_10614,N_10417,N_10460);
and U10615 (N_10615,N_10479,N_10347);
or U10616 (N_10616,N_10427,N_10397);
xnor U10617 (N_10617,N_10285,N_10256);
nand U10618 (N_10618,N_10252,N_10386);
and U10619 (N_10619,N_10333,N_10442);
or U10620 (N_10620,N_10491,N_10320);
xor U10621 (N_10621,N_10302,N_10437);
or U10622 (N_10622,N_10393,N_10294);
xnor U10623 (N_10623,N_10261,N_10441);
nand U10624 (N_10624,N_10341,N_10465);
and U10625 (N_10625,N_10432,N_10280);
and U10626 (N_10626,N_10290,N_10466);
or U10627 (N_10627,N_10448,N_10447);
or U10628 (N_10628,N_10282,N_10382);
nand U10629 (N_10629,N_10273,N_10313);
nor U10630 (N_10630,N_10331,N_10250);
xor U10631 (N_10631,N_10377,N_10480);
or U10632 (N_10632,N_10440,N_10447);
and U10633 (N_10633,N_10331,N_10385);
or U10634 (N_10634,N_10348,N_10419);
and U10635 (N_10635,N_10471,N_10488);
nand U10636 (N_10636,N_10272,N_10405);
or U10637 (N_10637,N_10492,N_10280);
or U10638 (N_10638,N_10310,N_10407);
xnor U10639 (N_10639,N_10461,N_10321);
nor U10640 (N_10640,N_10468,N_10404);
nand U10641 (N_10641,N_10337,N_10463);
xnor U10642 (N_10642,N_10352,N_10402);
or U10643 (N_10643,N_10332,N_10480);
and U10644 (N_10644,N_10353,N_10338);
and U10645 (N_10645,N_10427,N_10384);
and U10646 (N_10646,N_10395,N_10360);
and U10647 (N_10647,N_10376,N_10373);
or U10648 (N_10648,N_10437,N_10271);
xnor U10649 (N_10649,N_10287,N_10314);
xor U10650 (N_10650,N_10390,N_10472);
nand U10651 (N_10651,N_10426,N_10307);
and U10652 (N_10652,N_10399,N_10414);
nor U10653 (N_10653,N_10362,N_10494);
xor U10654 (N_10654,N_10272,N_10293);
and U10655 (N_10655,N_10461,N_10420);
or U10656 (N_10656,N_10290,N_10367);
or U10657 (N_10657,N_10461,N_10256);
xnor U10658 (N_10658,N_10302,N_10482);
xor U10659 (N_10659,N_10427,N_10293);
nor U10660 (N_10660,N_10330,N_10470);
and U10661 (N_10661,N_10316,N_10282);
nor U10662 (N_10662,N_10463,N_10396);
and U10663 (N_10663,N_10431,N_10277);
nand U10664 (N_10664,N_10377,N_10491);
xor U10665 (N_10665,N_10338,N_10447);
nand U10666 (N_10666,N_10412,N_10360);
nand U10667 (N_10667,N_10392,N_10336);
nor U10668 (N_10668,N_10306,N_10489);
nand U10669 (N_10669,N_10436,N_10385);
nand U10670 (N_10670,N_10256,N_10386);
nor U10671 (N_10671,N_10494,N_10359);
or U10672 (N_10672,N_10427,N_10420);
xnor U10673 (N_10673,N_10261,N_10252);
xor U10674 (N_10674,N_10416,N_10456);
nand U10675 (N_10675,N_10322,N_10432);
xor U10676 (N_10676,N_10371,N_10251);
nor U10677 (N_10677,N_10425,N_10323);
xor U10678 (N_10678,N_10370,N_10366);
nor U10679 (N_10679,N_10469,N_10260);
nand U10680 (N_10680,N_10435,N_10356);
nor U10681 (N_10681,N_10303,N_10447);
nor U10682 (N_10682,N_10463,N_10419);
xor U10683 (N_10683,N_10364,N_10348);
nor U10684 (N_10684,N_10316,N_10252);
and U10685 (N_10685,N_10360,N_10393);
xnor U10686 (N_10686,N_10337,N_10393);
and U10687 (N_10687,N_10442,N_10253);
or U10688 (N_10688,N_10344,N_10354);
nand U10689 (N_10689,N_10461,N_10375);
nand U10690 (N_10690,N_10449,N_10439);
xor U10691 (N_10691,N_10421,N_10266);
nor U10692 (N_10692,N_10441,N_10321);
nand U10693 (N_10693,N_10326,N_10411);
nand U10694 (N_10694,N_10343,N_10418);
or U10695 (N_10695,N_10352,N_10405);
nor U10696 (N_10696,N_10489,N_10385);
nand U10697 (N_10697,N_10289,N_10271);
nand U10698 (N_10698,N_10283,N_10374);
and U10699 (N_10699,N_10436,N_10393);
and U10700 (N_10700,N_10439,N_10454);
xnor U10701 (N_10701,N_10472,N_10491);
nand U10702 (N_10702,N_10379,N_10397);
and U10703 (N_10703,N_10391,N_10315);
nor U10704 (N_10704,N_10291,N_10475);
nand U10705 (N_10705,N_10403,N_10284);
and U10706 (N_10706,N_10307,N_10395);
or U10707 (N_10707,N_10398,N_10335);
nand U10708 (N_10708,N_10295,N_10446);
xor U10709 (N_10709,N_10406,N_10382);
or U10710 (N_10710,N_10406,N_10369);
and U10711 (N_10711,N_10278,N_10374);
or U10712 (N_10712,N_10483,N_10397);
nor U10713 (N_10713,N_10406,N_10287);
nor U10714 (N_10714,N_10448,N_10252);
and U10715 (N_10715,N_10258,N_10460);
nor U10716 (N_10716,N_10263,N_10292);
xor U10717 (N_10717,N_10250,N_10344);
nor U10718 (N_10718,N_10317,N_10384);
xor U10719 (N_10719,N_10476,N_10261);
xor U10720 (N_10720,N_10327,N_10493);
and U10721 (N_10721,N_10327,N_10329);
xnor U10722 (N_10722,N_10444,N_10285);
and U10723 (N_10723,N_10469,N_10475);
or U10724 (N_10724,N_10329,N_10391);
nand U10725 (N_10725,N_10405,N_10416);
nand U10726 (N_10726,N_10287,N_10385);
or U10727 (N_10727,N_10481,N_10394);
xor U10728 (N_10728,N_10294,N_10255);
nand U10729 (N_10729,N_10259,N_10390);
and U10730 (N_10730,N_10295,N_10450);
nor U10731 (N_10731,N_10283,N_10295);
or U10732 (N_10732,N_10304,N_10375);
xor U10733 (N_10733,N_10306,N_10369);
xor U10734 (N_10734,N_10481,N_10430);
or U10735 (N_10735,N_10461,N_10313);
or U10736 (N_10736,N_10353,N_10380);
or U10737 (N_10737,N_10417,N_10475);
nor U10738 (N_10738,N_10440,N_10263);
nand U10739 (N_10739,N_10380,N_10460);
or U10740 (N_10740,N_10418,N_10305);
xnor U10741 (N_10741,N_10416,N_10273);
xnor U10742 (N_10742,N_10268,N_10355);
nor U10743 (N_10743,N_10427,N_10460);
nand U10744 (N_10744,N_10345,N_10383);
nand U10745 (N_10745,N_10344,N_10406);
and U10746 (N_10746,N_10441,N_10316);
and U10747 (N_10747,N_10383,N_10444);
nor U10748 (N_10748,N_10478,N_10366);
or U10749 (N_10749,N_10368,N_10432);
and U10750 (N_10750,N_10680,N_10588);
nor U10751 (N_10751,N_10596,N_10747);
nor U10752 (N_10752,N_10713,N_10547);
xor U10753 (N_10753,N_10624,N_10659);
and U10754 (N_10754,N_10562,N_10669);
nand U10755 (N_10755,N_10571,N_10687);
nor U10756 (N_10756,N_10725,N_10568);
xor U10757 (N_10757,N_10678,N_10663);
or U10758 (N_10758,N_10619,N_10598);
nand U10759 (N_10759,N_10548,N_10511);
and U10760 (N_10760,N_10664,N_10708);
nand U10761 (N_10761,N_10650,N_10580);
and U10762 (N_10762,N_10572,N_10696);
and U10763 (N_10763,N_10577,N_10600);
nor U10764 (N_10764,N_10576,N_10656);
and U10765 (N_10765,N_10585,N_10605);
nor U10766 (N_10766,N_10666,N_10734);
and U10767 (N_10767,N_10639,N_10525);
nand U10768 (N_10768,N_10565,N_10699);
nand U10769 (N_10769,N_10646,N_10712);
nand U10770 (N_10770,N_10684,N_10643);
nor U10771 (N_10771,N_10567,N_10545);
and U10772 (N_10772,N_10535,N_10675);
nand U10773 (N_10773,N_10508,N_10622);
or U10774 (N_10774,N_10590,N_10717);
xor U10775 (N_10775,N_10737,N_10701);
xor U10776 (N_10776,N_10569,N_10595);
xor U10777 (N_10777,N_10673,N_10514);
xnor U10778 (N_10778,N_10703,N_10670);
xnor U10779 (N_10779,N_10632,N_10745);
nor U10780 (N_10780,N_10536,N_10587);
and U10781 (N_10781,N_10606,N_10665);
and U10782 (N_10782,N_10733,N_10630);
or U10783 (N_10783,N_10652,N_10607);
or U10784 (N_10784,N_10540,N_10515);
or U10785 (N_10785,N_10529,N_10566);
xnor U10786 (N_10786,N_10517,N_10724);
xnor U10787 (N_10787,N_10718,N_10671);
nor U10788 (N_10788,N_10532,N_10629);
and U10789 (N_10789,N_10626,N_10504);
nand U10790 (N_10790,N_10557,N_10592);
xor U10791 (N_10791,N_10520,N_10731);
nor U10792 (N_10792,N_10561,N_10645);
and U10793 (N_10793,N_10640,N_10594);
nor U10794 (N_10794,N_10519,N_10705);
or U10795 (N_10795,N_10593,N_10710);
and U10796 (N_10796,N_10716,N_10608);
nor U10797 (N_10797,N_10621,N_10702);
xor U10798 (N_10798,N_10554,N_10628);
xor U10799 (N_10799,N_10558,N_10611);
nand U10800 (N_10800,N_10527,N_10615);
and U10801 (N_10801,N_10677,N_10722);
and U10802 (N_10802,N_10563,N_10732);
nand U10803 (N_10803,N_10638,N_10668);
nand U10804 (N_10804,N_10522,N_10573);
nor U10805 (N_10805,N_10648,N_10721);
and U10806 (N_10806,N_10667,N_10521);
and U10807 (N_10807,N_10686,N_10604);
xnor U10808 (N_10808,N_10586,N_10609);
or U10809 (N_10809,N_10637,N_10591);
xnor U10810 (N_10810,N_10583,N_10662);
or U10811 (N_10811,N_10743,N_10575);
or U10812 (N_10812,N_10534,N_10556);
or U10813 (N_10813,N_10570,N_10582);
and U10814 (N_10814,N_10502,N_10706);
nor U10815 (N_10815,N_10660,N_10505);
or U10816 (N_10816,N_10711,N_10616);
xor U10817 (N_10817,N_10681,N_10719);
nand U10818 (N_10818,N_10651,N_10542);
nor U10819 (N_10819,N_10507,N_10693);
or U10820 (N_10820,N_10523,N_10715);
and U10821 (N_10821,N_10612,N_10676);
nand U10822 (N_10822,N_10501,N_10634);
or U10823 (N_10823,N_10738,N_10528);
nor U10824 (N_10824,N_10533,N_10655);
xor U10825 (N_10825,N_10530,N_10692);
nand U10826 (N_10826,N_10506,N_10682);
nor U10827 (N_10827,N_10579,N_10553);
and U10828 (N_10828,N_10574,N_10516);
nand U10829 (N_10829,N_10647,N_10589);
nand U10830 (N_10830,N_10564,N_10672);
or U10831 (N_10831,N_10661,N_10538);
and U10832 (N_10832,N_10642,N_10625);
nor U10833 (N_10833,N_10513,N_10539);
or U10834 (N_10834,N_10510,N_10623);
nand U10835 (N_10835,N_10658,N_10500);
and U10836 (N_10836,N_10578,N_10729);
and U10837 (N_10837,N_10700,N_10739);
or U10838 (N_10838,N_10620,N_10560);
nand U10839 (N_10839,N_10730,N_10653);
nand U10840 (N_10840,N_10531,N_10741);
and U10841 (N_10841,N_10631,N_10726);
or U10842 (N_10842,N_10627,N_10654);
or U10843 (N_10843,N_10691,N_10742);
nand U10844 (N_10844,N_10636,N_10551);
or U10845 (N_10845,N_10617,N_10601);
and U10846 (N_10846,N_10748,N_10688);
or U10847 (N_10847,N_10599,N_10559);
nand U10848 (N_10848,N_10550,N_10690);
nor U10849 (N_10849,N_10714,N_10707);
and U10850 (N_10850,N_10503,N_10704);
nand U10851 (N_10851,N_10735,N_10610);
nor U10852 (N_10852,N_10657,N_10685);
and U10853 (N_10853,N_10543,N_10633);
and U10854 (N_10854,N_10537,N_10644);
nor U10855 (N_10855,N_10727,N_10584);
or U10856 (N_10856,N_10744,N_10512);
nand U10857 (N_10857,N_10603,N_10683);
or U10858 (N_10858,N_10698,N_10544);
nor U10859 (N_10859,N_10613,N_10740);
xor U10860 (N_10860,N_10746,N_10736);
nand U10861 (N_10861,N_10546,N_10695);
nand U10862 (N_10862,N_10674,N_10541);
xnor U10863 (N_10863,N_10618,N_10614);
or U10864 (N_10864,N_10518,N_10526);
and U10865 (N_10865,N_10552,N_10728);
nand U10866 (N_10866,N_10649,N_10749);
nor U10867 (N_10867,N_10689,N_10720);
xnor U10868 (N_10868,N_10723,N_10679);
and U10869 (N_10869,N_10549,N_10581);
or U10870 (N_10870,N_10635,N_10524);
nor U10871 (N_10871,N_10641,N_10709);
nor U10872 (N_10872,N_10555,N_10602);
nand U10873 (N_10873,N_10694,N_10697);
xor U10874 (N_10874,N_10509,N_10597);
and U10875 (N_10875,N_10660,N_10543);
and U10876 (N_10876,N_10591,N_10732);
and U10877 (N_10877,N_10559,N_10509);
and U10878 (N_10878,N_10552,N_10562);
or U10879 (N_10879,N_10661,N_10648);
nor U10880 (N_10880,N_10594,N_10592);
xor U10881 (N_10881,N_10607,N_10720);
xnor U10882 (N_10882,N_10716,N_10739);
or U10883 (N_10883,N_10684,N_10625);
nand U10884 (N_10884,N_10745,N_10681);
nand U10885 (N_10885,N_10525,N_10533);
and U10886 (N_10886,N_10664,N_10653);
nand U10887 (N_10887,N_10553,N_10660);
nand U10888 (N_10888,N_10583,N_10666);
or U10889 (N_10889,N_10651,N_10742);
xnor U10890 (N_10890,N_10544,N_10567);
and U10891 (N_10891,N_10505,N_10665);
nand U10892 (N_10892,N_10612,N_10637);
or U10893 (N_10893,N_10529,N_10527);
nor U10894 (N_10894,N_10650,N_10607);
or U10895 (N_10895,N_10641,N_10727);
or U10896 (N_10896,N_10535,N_10620);
and U10897 (N_10897,N_10618,N_10674);
xnor U10898 (N_10898,N_10592,N_10683);
nor U10899 (N_10899,N_10536,N_10528);
nor U10900 (N_10900,N_10626,N_10704);
nor U10901 (N_10901,N_10689,N_10620);
and U10902 (N_10902,N_10677,N_10612);
nor U10903 (N_10903,N_10568,N_10549);
nor U10904 (N_10904,N_10719,N_10534);
nor U10905 (N_10905,N_10683,N_10557);
xnor U10906 (N_10906,N_10649,N_10657);
and U10907 (N_10907,N_10661,N_10555);
or U10908 (N_10908,N_10657,N_10684);
xor U10909 (N_10909,N_10716,N_10591);
and U10910 (N_10910,N_10590,N_10589);
nand U10911 (N_10911,N_10704,N_10516);
xor U10912 (N_10912,N_10567,N_10643);
nor U10913 (N_10913,N_10712,N_10716);
nor U10914 (N_10914,N_10734,N_10583);
and U10915 (N_10915,N_10630,N_10632);
nor U10916 (N_10916,N_10684,N_10700);
nor U10917 (N_10917,N_10625,N_10639);
nor U10918 (N_10918,N_10706,N_10557);
or U10919 (N_10919,N_10626,N_10723);
nand U10920 (N_10920,N_10691,N_10560);
nor U10921 (N_10921,N_10605,N_10637);
or U10922 (N_10922,N_10625,N_10670);
or U10923 (N_10923,N_10560,N_10748);
nand U10924 (N_10924,N_10540,N_10664);
xor U10925 (N_10925,N_10591,N_10633);
nand U10926 (N_10926,N_10505,N_10546);
and U10927 (N_10927,N_10685,N_10698);
nor U10928 (N_10928,N_10657,N_10614);
or U10929 (N_10929,N_10625,N_10692);
nor U10930 (N_10930,N_10535,N_10593);
xnor U10931 (N_10931,N_10644,N_10621);
or U10932 (N_10932,N_10746,N_10581);
or U10933 (N_10933,N_10575,N_10579);
xor U10934 (N_10934,N_10520,N_10672);
or U10935 (N_10935,N_10702,N_10544);
nor U10936 (N_10936,N_10575,N_10654);
nand U10937 (N_10937,N_10680,N_10731);
or U10938 (N_10938,N_10514,N_10742);
nand U10939 (N_10939,N_10525,N_10570);
nor U10940 (N_10940,N_10744,N_10647);
xnor U10941 (N_10941,N_10524,N_10715);
or U10942 (N_10942,N_10554,N_10518);
xnor U10943 (N_10943,N_10664,N_10524);
or U10944 (N_10944,N_10656,N_10524);
nor U10945 (N_10945,N_10672,N_10707);
nand U10946 (N_10946,N_10728,N_10507);
and U10947 (N_10947,N_10594,N_10610);
xor U10948 (N_10948,N_10615,N_10537);
or U10949 (N_10949,N_10684,N_10594);
and U10950 (N_10950,N_10539,N_10528);
xor U10951 (N_10951,N_10585,N_10669);
xnor U10952 (N_10952,N_10699,N_10596);
xor U10953 (N_10953,N_10572,N_10672);
nand U10954 (N_10954,N_10676,N_10716);
nand U10955 (N_10955,N_10701,N_10564);
and U10956 (N_10956,N_10631,N_10508);
nor U10957 (N_10957,N_10559,N_10715);
or U10958 (N_10958,N_10530,N_10715);
and U10959 (N_10959,N_10678,N_10606);
or U10960 (N_10960,N_10507,N_10656);
and U10961 (N_10961,N_10556,N_10537);
or U10962 (N_10962,N_10553,N_10566);
and U10963 (N_10963,N_10517,N_10520);
xnor U10964 (N_10964,N_10647,N_10635);
nand U10965 (N_10965,N_10718,N_10519);
or U10966 (N_10966,N_10740,N_10530);
or U10967 (N_10967,N_10715,N_10727);
nand U10968 (N_10968,N_10638,N_10706);
nor U10969 (N_10969,N_10518,N_10569);
xnor U10970 (N_10970,N_10744,N_10589);
nand U10971 (N_10971,N_10504,N_10650);
nand U10972 (N_10972,N_10551,N_10671);
nand U10973 (N_10973,N_10601,N_10692);
or U10974 (N_10974,N_10688,N_10638);
nor U10975 (N_10975,N_10657,N_10526);
or U10976 (N_10976,N_10657,N_10575);
nor U10977 (N_10977,N_10726,N_10640);
nand U10978 (N_10978,N_10537,N_10663);
nor U10979 (N_10979,N_10505,N_10554);
or U10980 (N_10980,N_10647,N_10747);
nand U10981 (N_10981,N_10646,N_10603);
nand U10982 (N_10982,N_10631,N_10507);
nand U10983 (N_10983,N_10556,N_10749);
nor U10984 (N_10984,N_10708,N_10632);
and U10985 (N_10985,N_10622,N_10637);
nand U10986 (N_10986,N_10527,N_10575);
xor U10987 (N_10987,N_10709,N_10683);
nand U10988 (N_10988,N_10556,N_10576);
xor U10989 (N_10989,N_10746,N_10694);
nor U10990 (N_10990,N_10706,N_10563);
or U10991 (N_10991,N_10694,N_10739);
nand U10992 (N_10992,N_10650,N_10725);
or U10993 (N_10993,N_10709,N_10593);
nand U10994 (N_10994,N_10641,N_10609);
and U10995 (N_10995,N_10636,N_10708);
nor U10996 (N_10996,N_10672,N_10562);
and U10997 (N_10997,N_10616,N_10602);
nor U10998 (N_10998,N_10724,N_10645);
nand U10999 (N_10999,N_10607,N_10749);
nand U11000 (N_11000,N_10969,N_10778);
or U11001 (N_11001,N_10774,N_10810);
xnor U11002 (N_11002,N_10933,N_10889);
and U11003 (N_11003,N_10826,N_10761);
and U11004 (N_11004,N_10956,N_10907);
xor U11005 (N_11005,N_10823,N_10800);
and U11006 (N_11006,N_10948,N_10968);
or U11007 (N_11007,N_10755,N_10875);
xnor U11008 (N_11008,N_10811,N_10750);
nand U11009 (N_11009,N_10777,N_10920);
xnor U11010 (N_11010,N_10849,N_10851);
and U11011 (N_11011,N_10841,N_10939);
and U11012 (N_11012,N_10883,N_10971);
nand U11013 (N_11013,N_10817,N_10863);
or U11014 (N_11014,N_10877,N_10819);
xnor U11015 (N_11015,N_10832,N_10768);
nand U11016 (N_11016,N_10775,N_10977);
or U11017 (N_11017,N_10813,N_10882);
nand U11018 (N_11018,N_10902,N_10936);
nand U11019 (N_11019,N_10890,N_10859);
nand U11020 (N_11020,N_10873,N_10757);
and U11021 (N_11021,N_10850,N_10862);
nor U11022 (N_11022,N_10974,N_10988);
xnor U11023 (N_11023,N_10764,N_10967);
nor U11024 (N_11024,N_10952,N_10912);
and U11025 (N_11025,N_10833,N_10904);
and U11026 (N_11026,N_10847,N_10756);
or U11027 (N_11027,N_10991,N_10994);
and U11028 (N_11028,N_10916,N_10887);
or U11029 (N_11029,N_10843,N_10760);
nand U11030 (N_11030,N_10866,N_10987);
or U11031 (N_11031,N_10802,N_10781);
or U11032 (N_11032,N_10923,N_10752);
nor U11033 (N_11033,N_10997,N_10790);
and U11034 (N_11034,N_10783,N_10930);
nor U11035 (N_11035,N_10938,N_10905);
nand U11036 (N_11036,N_10769,N_10865);
nor U11037 (N_11037,N_10899,N_10792);
and U11038 (N_11038,N_10979,N_10780);
or U11039 (N_11039,N_10796,N_10824);
or U11040 (N_11040,N_10942,N_10945);
nand U11041 (N_11041,N_10839,N_10835);
xnor U11042 (N_11042,N_10919,N_10753);
nand U11043 (N_11043,N_10922,N_10791);
and U11044 (N_11044,N_10868,N_10857);
and U11045 (N_11045,N_10888,N_10989);
or U11046 (N_11046,N_10763,N_10874);
xor U11047 (N_11047,N_10871,N_10898);
or U11048 (N_11048,N_10869,N_10954);
or U11049 (N_11049,N_10966,N_10815);
nor U11050 (N_11050,N_10840,N_10758);
nor U11051 (N_11051,N_10953,N_10829);
nor U11052 (N_11052,N_10911,N_10998);
nor U11053 (N_11053,N_10897,N_10986);
nor U11054 (N_11054,N_10807,N_10947);
or U11055 (N_11055,N_10965,N_10771);
nand U11056 (N_11056,N_10921,N_10981);
nor U11057 (N_11057,N_10838,N_10894);
nor U11058 (N_11058,N_10782,N_10928);
nor U11059 (N_11059,N_10961,N_10992);
xor U11060 (N_11060,N_10949,N_10805);
or U11061 (N_11061,N_10821,N_10766);
nor U11062 (N_11062,N_10809,N_10957);
xnor U11063 (N_11063,N_10804,N_10931);
or U11064 (N_11064,N_10880,N_10937);
or U11065 (N_11065,N_10825,N_10795);
or U11066 (N_11066,N_10858,N_10844);
xor U11067 (N_11067,N_10785,N_10754);
nor U11068 (N_11068,N_10915,N_10798);
and U11069 (N_11069,N_10935,N_10959);
nor U11070 (N_11070,N_10765,N_10980);
nand U11071 (N_11071,N_10794,N_10845);
or U11072 (N_11072,N_10946,N_10926);
nor U11073 (N_11073,N_10895,N_10940);
and U11074 (N_11074,N_10993,N_10941);
nand U11075 (N_11075,N_10878,N_10834);
or U11076 (N_11076,N_10784,N_10908);
nor U11077 (N_11077,N_10881,N_10884);
or U11078 (N_11078,N_10818,N_10836);
nor U11079 (N_11079,N_10885,N_10886);
nand U11080 (N_11080,N_10892,N_10831);
nor U11081 (N_11081,N_10879,N_10978);
xor U11082 (N_11082,N_10893,N_10853);
and U11083 (N_11083,N_10779,N_10906);
and U11084 (N_11084,N_10972,N_10996);
xor U11085 (N_11085,N_10909,N_10918);
nand U11086 (N_11086,N_10896,N_10995);
xnor U11087 (N_11087,N_10861,N_10799);
xor U11088 (N_11088,N_10934,N_10901);
or U11089 (N_11089,N_10773,N_10820);
and U11090 (N_11090,N_10951,N_10990);
nand U11091 (N_11091,N_10958,N_10856);
and U11092 (N_11092,N_10914,N_10924);
and U11093 (N_11093,N_10822,N_10950);
nor U11094 (N_11094,N_10854,N_10797);
and U11095 (N_11095,N_10842,N_10943);
or U11096 (N_11096,N_10976,N_10929);
or U11097 (N_11097,N_10770,N_10910);
xor U11098 (N_11098,N_10787,N_10860);
xnor U11099 (N_11099,N_10876,N_10944);
or U11100 (N_11100,N_10759,N_10827);
nand U11101 (N_11101,N_10867,N_10872);
nor U11102 (N_11102,N_10793,N_10806);
nand U11103 (N_11103,N_10975,N_10983);
nor U11104 (N_11104,N_10828,N_10808);
nand U11105 (N_11105,N_10762,N_10788);
xor U11106 (N_11106,N_10962,N_10927);
xnor U11107 (N_11107,N_10985,N_10870);
and U11108 (N_11108,N_10814,N_10751);
xnor U11109 (N_11109,N_10891,N_10970);
and U11110 (N_11110,N_10801,N_10776);
nor U11111 (N_11111,N_10812,N_10932);
or U11112 (N_11112,N_10903,N_10964);
and U11113 (N_11113,N_10955,N_10925);
nand U11114 (N_11114,N_10816,N_10864);
nor U11115 (N_11115,N_10837,N_10900);
xor U11116 (N_11116,N_10772,N_10789);
xor U11117 (N_11117,N_10786,N_10984);
xnor U11118 (N_11118,N_10963,N_10803);
xnor U11119 (N_11119,N_10846,N_10852);
or U11120 (N_11120,N_10913,N_10848);
nor U11121 (N_11121,N_10982,N_10999);
and U11122 (N_11122,N_10830,N_10917);
nand U11123 (N_11123,N_10973,N_10767);
nand U11124 (N_11124,N_10855,N_10960);
nor U11125 (N_11125,N_10832,N_10825);
xnor U11126 (N_11126,N_10967,N_10775);
nand U11127 (N_11127,N_10791,N_10850);
nor U11128 (N_11128,N_10775,N_10832);
or U11129 (N_11129,N_10843,N_10803);
nor U11130 (N_11130,N_10851,N_10991);
nor U11131 (N_11131,N_10924,N_10750);
nor U11132 (N_11132,N_10795,N_10983);
xor U11133 (N_11133,N_10858,N_10882);
and U11134 (N_11134,N_10900,N_10968);
and U11135 (N_11135,N_10984,N_10930);
xnor U11136 (N_11136,N_10886,N_10770);
or U11137 (N_11137,N_10809,N_10932);
nor U11138 (N_11138,N_10934,N_10808);
nor U11139 (N_11139,N_10858,N_10820);
and U11140 (N_11140,N_10877,N_10796);
and U11141 (N_11141,N_10983,N_10979);
xnor U11142 (N_11142,N_10916,N_10921);
or U11143 (N_11143,N_10938,N_10925);
and U11144 (N_11144,N_10972,N_10951);
or U11145 (N_11145,N_10961,N_10918);
and U11146 (N_11146,N_10860,N_10830);
xnor U11147 (N_11147,N_10782,N_10845);
or U11148 (N_11148,N_10938,N_10950);
nor U11149 (N_11149,N_10888,N_10856);
nand U11150 (N_11150,N_10800,N_10910);
nor U11151 (N_11151,N_10846,N_10882);
nor U11152 (N_11152,N_10799,N_10803);
xor U11153 (N_11153,N_10803,N_10778);
or U11154 (N_11154,N_10871,N_10860);
or U11155 (N_11155,N_10934,N_10858);
or U11156 (N_11156,N_10940,N_10846);
nor U11157 (N_11157,N_10790,N_10968);
nor U11158 (N_11158,N_10920,N_10804);
nand U11159 (N_11159,N_10987,N_10975);
nand U11160 (N_11160,N_10792,N_10893);
xnor U11161 (N_11161,N_10986,N_10837);
or U11162 (N_11162,N_10914,N_10823);
xnor U11163 (N_11163,N_10762,N_10961);
and U11164 (N_11164,N_10756,N_10881);
xor U11165 (N_11165,N_10810,N_10816);
xor U11166 (N_11166,N_10932,N_10820);
nand U11167 (N_11167,N_10807,N_10864);
xnor U11168 (N_11168,N_10964,N_10826);
or U11169 (N_11169,N_10996,N_10953);
and U11170 (N_11170,N_10948,N_10793);
nand U11171 (N_11171,N_10998,N_10754);
nand U11172 (N_11172,N_10913,N_10979);
xor U11173 (N_11173,N_10766,N_10853);
nand U11174 (N_11174,N_10862,N_10917);
or U11175 (N_11175,N_10952,N_10965);
and U11176 (N_11176,N_10813,N_10867);
nor U11177 (N_11177,N_10875,N_10857);
xor U11178 (N_11178,N_10879,N_10976);
xnor U11179 (N_11179,N_10995,N_10908);
and U11180 (N_11180,N_10894,N_10820);
nand U11181 (N_11181,N_10887,N_10880);
and U11182 (N_11182,N_10935,N_10914);
or U11183 (N_11183,N_10864,N_10899);
xnor U11184 (N_11184,N_10806,N_10812);
nand U11185 (N_11185,N_10809,N_10911);
nor U11186 (N_11186,N_10935,N_10987);
or U11187 (N_11187,N_10965,N_10928);
and U11188 (N_11188,N_10830,N_10935);
xnor U11189 (N_11189,N_10787,N_10833);
or U11190 (N_11190,N_10782,N_10989);
and U11191 (N_11191,N_10835,N_10771);
and U11192 (N_11192,N_10910,N_10872);
nand U11193 (N_11193,N_10757,N_10786);
nand U11194 (N_11194,N_10976,N_10817);
nand U11195 (N_11195,N_10977,N_10843);
nand U11196 (N_11196,N_10936,N_10751);
and U11197 (N_11197,N_10995,N_10952);
nand U11198 (N_11198,N_10985,N_10974);
nand U11199 (N_11199,N_10972,N_10794);
or U11200 (N_11200,N_10927,N_10807);
or U11201 (N_11201,N_10802,N_10862);
and U11202 (N_11202,N_10822,N_10974);
nand U11203 (N_11203,N_10793,N_10820);
or U11204 (N_11204,N_10887,N_10835);
and U11205 (N_11205,N_10857,N_10809);
and U11206 (N_11206,N_10975,N_10873);
and U11207 (N_11207,N_10759,N_10810);
xor U11208 (N_11208,N_10876,N_10774);
and U11209 (N_11209,N_10862,N_10869);
xnor U11210 (N_11210,N_10920,N_10796);
or U11211 (N_11211,N_10780,N_10918);
nor U11212 (N_11212,N_10882,N_10965);
xor U11213 (N_11213,N_10989,N_10771);
or U11214 (N_11214,N_10888,N_10944);
or U11215 (N_11215,N_10900,N_10910);
and U11216 (N_11216,N_10947,N_10945);
nand U11217 (N_11217,N_10834,N_10954);
and U11218 (N_11218,N_10955,N_10892);
nor U11219 (N_11219,N_10903,N_10798);
and U11220 (N_11220,N_10876,N_10770);
or U11221 (N_11221,N_10782,N_10816);
and U11222 (N_11222,N_10868,N_10750);
nand U11223 (N_11223,N_10994,N_10894);
nor U11224 (N_11224,N_10845,N_10802);
nand U11225 (N_11225,N_10940,N_10978);
xor U11226 (N_11226,N_10941,N_10996);
nand U11227 (N_11227,N_10768,N_10896);
and U11228 (N_11228,N_10902,N_10893);
nor U11229 (N_11229,N_10818,N_10857);
or U11230 (N_11230,N_10942,N_10857);
nor U11231 (N_11231,N_10989,N_10968);
nand U11232 (N_11232,N_10904,N_10905);
nor U11233 (N_11233,N_10850,N_10833);
nor U11234 (N_11234,N_10964,N_10918);
nand U11235 (N_11235,N_10857,N_10908);
and U11236 (N_11236,N_10861,N_10865);
and U11237 (N_11237,N_10839,N_10966);
xnor U11238 (N_11238,N_10798,N_10762);
nor U11239 (N_11239,N_10932,N_10896);
or U11240 (N_11240,N_10971,N_10867);
or U11241 (N_11241,N_10861,N_10817);
or U11242 (N_11242,N_10876,N_10802);
xnor U11243 (N_11243,N_10943,N_10783);
and U11244 (N_11244,N_10956,N_10911);
or U11245 (N_11245,N_10939,N_10977);
xor U11246 (N_11246,N_10829,N_10757);
nor U11247 (N_11247,N_10844,N_10963);
and U11248 (N_11248,N_10941,N_10854);
and U11249 (N_11249,N_10794,N_10941);
and U11250 (N_11250,N_11059,N_11172);
and U11251 (N_11251,N_11164,N_11070);
nor U11252 (N_11252,N_11103,N_11010);
or U11253 (N_11253,N_11209,N_11182);
and U11254 (N_11254,N_11248,N_11204);
nor U11255 (N_11255,N_11023,N_11246);
nor U11256 (N_11256,N_11210,N_11086);
or U11257 (N_11257,N_11180,N_11161);
xnor U11258 (N_11258,N_11163,N_11237);
nor U11259 (N_11259,N_11061,N_11045);
and U11260 (N_11260,N_11082,N_11242);
or U11261 (N_11261,N_11033,N_11102);
or U11262 (N_11262,N_11247,N_11143);
nand U11263 (N_11263,N_11175,N_11094);
nor U11264 (N_11264,N_11193,N_11043);
or U11265 (N_11265,N_11171,N_11063);
nand U11266 (N_11266,N_11200,N_11190);
nor U11267 (N_11267,N_11145,N_11092);
and U11268 (N_11268,N_11126,N_11024);
xor U11269 (N_11269,N_11220,N_11060);
xor U11270 (N_11270,N_11212,N_11104);
xor U11271 (N_11271,N_11123,N_11158);
and U11272 (N_11272,N_11199,N_11111);
xor U11273 (N_11273,N_11122,N_11165);
xnor U11274 (N_11274,N_11095,N_11150);
or U11275 (N_11275,N_11176,N_11062);
and U11276 (N_11276,N_11013,N_11219);
or U11277 (N_11277,N_11213,N_11167);
xnor U11278 (N_11278,N_11117,N_11072);
and U11279 (N_11279,N_11148,N_11008);
and U11280 (N_11280,N_11053,N_11106);
nand U11281 (N_11281,N_11173,N_11138);
and U11282 (N_11282,N_11157,N_11196);
nand U11283 (N_11283,N_11056,N_11118);
xnor U11284 (N_11284,N_11216,N_11130);
and U11285 (N_11285,N_11127,N_11064);
nor U11286 (N_11286,N_11132,N_11168);
nand U11287 (N_11287,N_11189,N_11039);
xor U11288 (N_11288,N_11003,N_11227);
or U11289 (N_11289,N_11113,N_11006);
and U11290 (N_11290,N_11208,N_11218);
xor U11291 (N_11291,N_11194,N_11048);
nand U11292 (N_11292,N_11203,N_11207);
nor U11293 (N_11293,N_11169,N_11239);
xnor U11294 (N_11294,N_11088,N_11046);
nand U11295 (N_11295,N_11058,N_11001);
xnor U11296 (N_11296,N_11037,N_11038);
nor U11297 (N_11297,N_11015,N_11052);
or U11298 (N_11298,N_11068,N_11151);
or U11299 (N_11299,N_11174,N_11206);
or U11300 (N_11300,N_11085,N_11134);
and U11301 (N_11301,N_11012,N_11125);
nand U11302 (N_11302,N_11146,N_11074);
or U11303 (N_11303,N_11186,N_11087);
nor U11304 (N_11304,N_11002,N_11119);
nand U11305 (N_11305,N_11071,N_11027);
nand U11306 (N_11306,N_11028,N_11110);
or U11307 (N_11307,N_11178,N_11047);
and U11308 (N_11308,N_11017,N_11042);
nand U11309 (N_11309,N_11223,N_11249);
or U11310 (N_11310,N_11044,N_11098);
xor U11311 (N_11311,N_11155,N_11244);
nor U11312 (N_11312,N_11066,N_11166);
nor U11313 (N_11313,N_11097,N_11049);
nor U11314 (N_11314,N_11004,N_11029);
xor U11315 (N_11315,N_11035,N_11211);
xnor U11316 (N_11316,N_11089,N_11141);
and U11317 (N_11317,N_11078,N_11234);
nand U11318 (N_11318,N_11214,N_11099);
or U11319 (N_11319,N_11065,N_11222);
nor U11320 (N_11320,N_11075,N_11225);
nor U11321 (N_11321,N_11187,N_11069);
and U11322 (N_11322,N_11215,N_11055);
nor U11323 (N_11323,N_11091,N_11217);
or U11324 (N_11324,N_11019,N_11235);
nand U11325 (N_11325,N_11073,N_11243);
xnor U11326 (N_11326,N_11057,N_11129);
and U11327 (N_11327,N_11205,N_11188);
xor U11328 (N_11328,N_11112,N_11241);
nand U11329 (N_11329,N_11133,N_11152);
xnor U11330 (N_11330,N_11018,N_11009);
and U11331 (N_11331,N_11226,N_11139);
nor U11332 (N_11332,N_11154,N_11128);
xor U11333 (N_11333,N_11121,N_11170);
xor U11334 (N_11334,N_11156,N_11080);
nor U11335 (N_11335,N_11108,N_11016);
or U11336 (N_11336,N_11021,N_11031);
nand U11337 (N_11337,N_11005,N_11153);
xnor U11338 (N_11338,N_11109,N_11084);
and U11339 (N_11339,N_11177,N_11184);
nand U11340 (N_11340,N_11115,N_11124);
or U11341 (N_11341,N_11032,N_11198);
xor U11342 (N_11342,N_11135,N_11179);
nand U11343 (N_11343,N_11240,N_11159);
or U11344 (N_11344,N_11181,N_11233);
and U11345 (N_11345,N_11034,N_11051);
or U11346 (N_11346,N_11195,N_11011);
nor U11347 (N_11347,N_11191,N_11185);
nand U11348 (N_11348,N_11036,N_11224);
and U11349 (N_11349,N_11120,N_11081);
xnor U11350 (N_11350,N_11020,N_11202);
and U11351 (N_11351,N_11077,N_11232);
nor U11352 (N_11352,N_11100,N_11192);
or U11353 (N_11353,N_11221,N_11114);
nor U11354 (N_11354,N_11183,N_11144);
nor U11355 (N_11355,N_11245,N_11041);
or U11356 (N_11356,N_11083,N_11067);
and U11357 (N_11357,N_11228,N_11142);
nor U11358 (N_11358,N_11136,N_11054);
xor U11359 (N_11359,N_11140,N_11236);
and U11360 (N_11360,N_11197,N_11116);
xor U11361 (N_11361,N_11090,N_11131);
nand U11362 (N_11362,N_11093,N_11050);
xnor U11363 (N_11363,N_11230,N_11201);
xnor U11364 (N_11364,N_11030,N_11014);
nor U11365 (N_11365,N_11147,N_11238);
or U11366 (N_11366,N_11231,N_11149);
nor U11367 (N_11367,N_11105,N_11000);
xnor U11368 (N_11368,N_11162,N_11040);
or U11369 (N_11369,N_11025,N_11079);
or U11370 (N_11370,N_11026,N_11137);
nor U11371 (N_11371,N_11007,N_11160);
or U11372 (N_11372,N_11101,N_11096);
or U11373 (N_11373,N_11076,N_11229);
or U11374 (N_11374,N_11107,N_11022);
nor U11375 (N_11375,N_11184,N_11243);
nor U11376 (N_11376,N_11050,N_11062);
nand U11377 (N_11377,N_11188,N_11008);
and U11378 (N_11378,N_11199,N_11110);
or U11379 (N_11379,N_11024,N_11205);
xnor U11380 (N_11380,N_11041,N_11149);
nor U11381 (N_11381,N_11157,N_11207);
and U11382 (N_11382,N_11169,N_11009);
nor U11383 (N_11383,N_11192,N_11141);
nand U11384 (N_11384,N_11077,N_11200);
and U11385 (N_11385,N_11209,N_11220);
or U11386 (N_11386,N_11067,N_11026);
xor U11387 (N_11387,N_11183,N_11232);
xor U11388 (N_11388,N_11174,N_11043);
and U11389 (N_11389,N_11105,N_11015);
nor U11390 (N_11390,N_11040,N_11166);
nor U11391 (N_11391,N_11067,N_11133);
and U11392 (N_11392,N_11233,N_11232);
or U11393 (N_11393,N_11175,N_11236);
or U11394 (N_11394,N_11024,N_11177);
nor U11395 (N_11395,N_11193,N_11057);
xor U11396 (N_11396,N_11008,N_11120);
xnor U11397 (N_11397,N_11030,N_11048);
xor U11398 (N_11398,N_11228,N_11238);
nor U11399 (N_11399,N_11044,N_11207);
nor U11400 (N_11400,N_11021,N_11152);
nand U11401 (N_11401,N_11034,N_11227);
nand U11402 (N_11402,N_11021,N_11137);
nand U11403 (N_11403,N_11017,N_11209);
nor U11404 (N_11404,N_11116,N_11134);
nand U11405 (N_11405,N_11027,N_11224);
nor U11406 (N_11406,N_11129,N_11156);
xnor U11407 (N_11407,N_11132,N_11079);
and U11408 (N_11408,N_11120,N_11073);
or U11409 (N_11409,N_11143,N_11153);
and U11410 (N_11410,N_11119,N_11062);
and U11411 (N_11411,N_11197,N_11109);
nor U11412 (N_11412,N_11201,N_11146);
nand U11413 (N_11413,N_11232,N_11085);
or U11414 (N_11414,N_11081,N_11211);
and U11415 (N_11415,N_11072,N_11002);
and U11416 (N_11416,N_11162,N_11195);
or U11417 (N_11417,N_11163,N_11138);
or U11418 (N_11418,N_11087,N_11217);
or U11419 (N_11419,N_11109,N_11025);
nand U11420 (N_11420,N_11071,N_11191);
xnor U11421 (N_11421,N_11192,N_11224);
or U11422 (N_11422,N_11141,N_11180);
or U11423 (N_11423,N_11183,N_11102);
nand U11424 (N_11424,N_11081,N_11233);
xor U11425 (N_11425,N_11098,N_11119);
xor U11426 (N_11426,N_11086,N_11150);
nand U11427 (N_11427,N_11236,N_11049);
or U11428 (N_11428,N_11124,N_11106);
or U11429 (N_11429,N_11230,N_11064);
and U11430 (N_11430,N_11204,N_11142);
xor U11431 (N_11431,N_11098,N_11015);
xor U11432 (N_11432,N_11053,N_11017);
nand U11433 (N_11433,N_11012,N_11152);
and U11434 (N_11434,N_11168,N_11126);
and U11435 (N_11435,N_11140,N_11104);
nor U11436 (N_11436,N_11211,N_11180);
nand U11437 (N_11437,N_11032,N_11139);
nand U11438 (N_11438,N_11071,N_11037);
or U11439 (N_11439,N_11130,N_11214);
xor U11440 (N_11440,N_11203,N_11046);
or U11441 (N_11441,N_11221,N_11174);
nand U11442 (N_11442,N_11184,N_11220);
and U11443 (N_11443,N_11174,N_11012);
nand U11444 (N_11444,N_11043,N_11162);
nor U11445 (N_11445,N_11050,N_11111);
nor U11446 (N_11446,N_11017,N_11124);
and U11447 (N_11447,N_11231,N_11007);
nor U11448 (N_11448,N_11055,N_11075);
xor U11449 (N_11449,N_11109,N_11062);
and U11450 (N_11450,N_11148,N_11086);
xnor U11451 (N_11451,N_11204,N_11086);
and U11452 (N_11452,N_11030,N_11145);
and U11453 (N_11453,N_11154,N_11049);
nor U11454 (N_11454,N_11016,N_11128);
nand U11455 (N_11455,N_11180,N_11184);
nor U11456 (N_11456,N_11001,N_11132);
or U11457 (N_11457,N_11006,N_11001);
and U11458 (N_11458,N_11133,N_11079);
nand U11459 (N_11459,N_11017,N_11242);
nor U11460 (N_11460,N_11067,N_11079);
nand U11461 (N_11461,N_11103,N_11177);
nand U11462 (N_11462,N_11130,N_11114);
xor U11463 (N_11463,N_11084,N_11179);
or U11464 (N_11464,N_11130,N_11141);
and U11465 (N_11465,N_11196,N_11194);
xnor U11466 (N_11466,N_11067,N_11238);
xnor U11467 (N_11467,N_11060,N_11041);
nor U11468 (N_11468,N_11111,N_11124);
nand U11469 (N_11469,N_11149,N_11119);
nand U11470 (N_11470,N_11212,N_11029);
nor U11471 (N_11471,N_11082,N_11196);
nor U11472 (N_11472,N_11247,N_11044);
nor U11473 (N_11473,N_11175,N_11006);
nand U11474 (N_11474,N_11011,N_11121);
xnor U11475 (N_11475,N_11191,N_11148);
nand U11476 (N_11476,N_11030,N_11211);
and U11477 (N_11477,N_11126,N_11119);
nor U11478 (N_11478,N_11060,N_11058);
nor U11479 (N_11479,N_11123,N_11107);
and U11480 (N_11480,N_11202,N_11026);
nand U11481 (N_11481,N_11241,N_11177);
xor U11482 (N_11482,N_11218,N_11164);
nor U11483 (N_11483,N_11184,N_11004);
and U11484 (N_11484,N_11178,N_11056);
nor U11485 (N_11485,N_11063,N_11055);
nand U11486 (N_11486,N_11139,N_11012);
and U11487 (N_11487,N_11193,N_11063);
or U11488 (N_11488,N_11015,N_11181);
nor U11489 (N_11489,N_11124,N_11021);
nand U11490 (N_11490,N_11161,N_11147);
or U11491 (N_11491,N_11245,N_11205);
and U11492 (N_11492,N_11211,N_11134);
or U11493 (N_11493,N_11035,N_11023);
or U11494 (N_11494,N_11159,N_11126);
or U11495 (N_11495,N_11144,N_11122);
xor U11496 (N_11496,N_11146,N_11034);
and U11497 (N_11497,N_11027,N_11187);
nand U11498 (N_11498,N_11154,N_11063);
nor U11499 (N_11499,N_11056,N_11141);
nor U11500 (N_11500,N_11481,N_11402);
or U11501 (N_11501,N_11443,N_11298);
nand U11502 (N_11502,N_11454,N_11318);
nand U11503 (N_11503,N_11476,N_11490);
xor U11504 (N_11504,N_11302,N_11282);
nor U11505 (N_11505,N_11472,N_11280);
or U11506 (N_11506,N_11449,N_11459);
or U11507 (N_11507,N_11495,N_11419);
or U11508 (N_11508,N_11285,N_11266);
xnor U11509 (N_11509,N_11373,N_11300);
and U11510 (N_11510,N_11406,N_11331);
or U11511 (N_11511,N_11347,N_11294);
nor U11512 (N_11512,N_11283,N_11417);
nand U11513 (N_11513,N_11326,N_11336);
nand U11514 (N_11514,N_11332,N_11363);
nor U11515 (N_11515,N_11440,N_11252);
nor U11516 (N_11516,N_11457,N_11384);
or U11517 (N_11517,N_11311,N_11425);
xnor U11518 (N_11518,N_11342,N_11256);
xor U11519 (N_11519,N_11376,N_11381);
and U11520 (N_11520,N_11405,N_11491);
nand U11521 (N_11521,N_11355,N_11487);
and U11522 (N_11522,N_11484,N_11343);
or U11523 (N_11523,N_11387,N_11414);
or U11524 (N_11524,N_11360,N_11400);
or U11525 (N_11525,N_11354,N_11250);
xor U11526 (N_11526,N_11409,N_11377);
and U11527 (N_11527,N_11492,N_11262);
or U11528 (N_11528,N_11295,N_11442);
and U11529 (N_11529,N_11396,N_11321);
xor U11530 (N_11530,N_11327,N_11395);
and U11531 (N_11531,N_11309,N_11392);
xnor U11532 (N_11532,N_11310,N_11398);
and U11533 (N_11533,N_11374,N_11483);
and U11534 (N_11534,N_11437,N_11279);
nand U11535 (N_11535,N_11290,N_11272);
or U11536 (N_11536,N_11452,N_11438);
xor U11537 (N_11537,N_11370,N_11284);
or U11538 (N_11538,N_11307,N_11352);
xor U11539 (N_11539,N_11391,N_11359);
or U11540 (N_11540,N_11386,N_11447);
and U11541 (N_11541,N_11274,N_11338);
or U11542 (N_11542,N_11308,N_11435);
xor U11543 (N_11543,N_11351,N_11275);
and U11544 (N_11544,N_11413,N_11305);
and U11545 (N_11545,N_11312,N_11340);
or U11546 (N_11546,N_11314,N_11291);
nor U11547 (N_11547,N_11463,N_11410);
xor U11548 (N_11548,N_11477,N_11334);
nor U11549 (N_11549,N_11431,N_11407);
nand U11550 (N_11550,N_11493,N_11324);
nor U11551 (N_11551,N_11255,N_11479);
or U11552 (N_11552,N_11323,N_11404);
xnor U11553 (N_11553,N_11445,N_11416);
xor U11554 (N_11554,N_11267,N_11315);
and U11555 (N_11555,N_11403,N_11270);
nor U11556 (N_11556,N_11455,N_11380);
or U11557 (N_11557,N_11488,N_11469);
nor U11558 (N_11558,N_11337,N_11464);
or U11559 (N_11559,N_11458,N_11480);
nand U11560 (N_11560,N_11357,N_11401);
and U11561 (N_11561,N_11433,N_11286);
and U11562 (N_11562,N_11341,N_11394);
or U11563 (N_11563,N_11273,N_11303);
and U11564 (N_11564,N_11426,N_11329);
xnor U11565 (N_11565,N_11299,N_11371);
nor U11566 (N_11566,N_11288,N_11497);
xor U11567 (N_11567,N_11325,N_11482);
and U11568 (N_11568,N_11261,N_11254);
or U11569 (N_11569,N_11368,N_11264);
and U11570 (N_11570,N_11268,N_11421);
nor U11571 (N_11571,N_11257,N_11260);
nand U11572 (N_11572,N_11420,N_11486);
nand U11573 (N_11573,N_11429,N_11375);
nor U11574 (N_11574,N_11385,N_11320);
or U11575 (N_11575,N_11446,N_11448);
nand U11576 (N_11576,N_11301,N_11453);
xnor U11577 (N_11577,N_11361,N_11296);
nor U11578 (N_11578,N_11263,N_11485);
nor U11579 (N_11579,N_11471,N_11430);
or U11580 (N_11580,N_11258,N_11439);
xnor U11581 (N_11581,N_11271,N_11292);
nor U11582 (N_11582,N_11478,N_11276);
xor U11583 (N_11583,N_11427,N_11397);
nand U11584 (N_11584,N_11378,N_11399);
nand U11585 (N_11585,N_11349,N_11415);
or U11586 (N_11586,N_11278,N_11251);
nor U11587 (N_11587,N_11322,N_11335);
xor U11588 (N_11588,N_11441,N_11259);
nand U11589 (N_11589,N_11328,N_11408);
nor U11590 (N_11590,N_11372,N_11316);
or U11591 (N_11591,N_11350,N_11393);
nand U11592 (N_11592,N_11346,N_11383);
nor U11593 (N_11593,N_11313,N_11277);
and U11594 (N_11594,N_11494,N_11319);
nor U11595 (N_11595,N_11356,N_11411);
or U11596 (N_11596,N_11297,N_11367);
and U11597 (N_11597,N_11382,N_11498);
nor U11598 (N_11598,N_11358,N_11475);
and U11599 (N_11599,N_11281,N_11287);
and U11600 (N_11600,N_11450,N_11436);
xor U11601 (N_11601,N_11473,N_11345);
xnor U11602 (N_11602,N_11366,N_11362);
xor U11603 (N_11603,N_11462,N_11388);
nor U11604 (N_11604,N_11474,N_11317);
xnor U11605 (N_11605,N_11496,N_11424);
nand U11606 (N_11606,N_11333,N_11465);
nor U11607 (N_11607,N_11466,N_11390);
nor U11608 (N_11608,N_11499,N_11304);
or U11609 (N_11609,N_11293,N_11253);
nand U11610 (N_11610,N_11369,N_11265);
and U11611 (N_11611,N_11348,N_11489);
and U11612 (N_11612,N_11353,N_11379);
xnor U11613 (N_11613,N_11389,N_11339);
nor U11614 (N_11614,N_11422,N_11365);
nor U11615 (N_11615,N_11467,N_11444);
and U11616 (N_11616,N_11269,N_11460);
nor U11617 (N_11617,N_11330,N_11456);
and U11618 (N_11618,N_11461,N_11434);
nor U11619 (N_11619,N_11306,N_11364);
and U11620 (N_11620,N_11344,N_11432);
nand U11621 (N_11621,N_11289,N_11451);
nor U11622 (N_11622,N_11468,N_11470);
nor U11623 (N_11623,N_11423,N_11428);
or U11624 (N_11624,N_11412,N_11418);
xor U11625 (N_11625,N_11285,N_11422);
xor U11626 (N_11626,N_11479,N_11457);
and U11627 (N_11627,N_11253,N_11254);
nor U11628 (N_11628,N_11450,N_11446);
nor U11629 (N_11629,N_11261,N_11392);
and U11630 (N_11630,N_11359,N_11331);
nand U11631 (N_11631,N_11368,N_11493);
nand U11632 (N_11632,N_11345,N_11272);
nand U11633 (N_11633,N_11393,N_11414);
nand U11634 (N_11634,N_11292,N_11263);
or U11635 (N_11635,N_11319,N_11382);
nand U11636 (N_11636,N_11438,N_11329);
nand U11637 (N_11637,N_11397,N_11364);
and U11638 (N_11638,N_11283,N_11252);
xnor U11639 (N_11639,N_11324,N_11297);
or U11640 (N_11640,N_11491,N_11453);
nand U11641 (N_11641,N_11335,N_11487);
nand U11642 (N_11642,N_11251,N_11339);
nor U11643 (N_11643,N_11467,N_11454);
nor U11644 (N_11644,N_11398,N_11314);
nand U11645 (N_11645,N_11371,N_11441);
nand U11646 (N_11646,N_11478,N_11413);
or U11647 (N_11647,N_11250,N_11455);
and U11648 (N_11648,N_11478,N_11341);
nor U11649 (N_11649,N_11345,N_11428);
nand U11650 (N_11650,N_11490,N_11294);
and U11651 (N_11651,N_11292,N_11353);
nor U11652 (N_11652,N_11338,N_11438);
and U11653 (N_11653,N_11438,N_11273);
xor U11654 (N_11654,N_11456,N_11449);
and U11655 (N_11655,N_11364,N_11344);
xor U11656 (N_11656,N_11268,N_11255);
nand U11657 (N_11657,N_11408,N_11487);
or U11658 (N_11658,N_11459,N_11305);
or U11659 (N_11659,N_11419,N_11315);
nand U11660 (N_11660,N_11402,N_11447);
nor U11661 (N_11661,N_11376,N_11325);
xor U11662 (N_11662,N_11314,N_11396);
and U11663 (N_11663,N_11482,N_11268);
xnor U11664 (N_11664,N_11460,N_11448);
xor U11665 (N_11665,N_11406,N_11411);
xor U11666 (N_11666,N_11386,N_11481);
nand U11667 (N_11667,N_11388,N_11411);
nor U11668 (N_11668,N_11306,N_11499);
xnor U11669 (N_11669,N_11255,N_11433);
nor U11670 (N_11670,N_11428,N_11457);
xor U11671 (N_11671,N_11359,N_11476);
nand U11672 (N_11672,N_11310,N_11461);
nand U11673 (N_11673,N_11303,N_11403);
and U11674 (N_11674,N_11268,N_11401);
nor U11675 (N_11675,N_11346,N_11397);
and U11676 (N_11676,N_11492,N_11360);
and U11677 (N_11677,N_11318,N_11386);
and U11678 (N_11678,N_11418,N_11339);
or U11679 (N_11679,N_11431,N_11455);
nand U11680 (N_11680,N_11257,N_11344);
or U11681 (N_11681,N_11357,N_11354);
nor U11682 (N_11682,N_11439,N_11426);
nor U11683 (N_11683,N_11351,N_11459);
nor U11684 (N_11684,N_11436,N_11460);
and U11685 (N_11685,N_11320,N_11455);
and U11686 (N_11686,N_11351,N_11377);
nand U11687 (N_11687,N_11371,N_11392);
and U11688 (N_11688,N_11294,N_11340);
nand U11689 (N_11689,N_11424,N_11439);
or U11690 (N_11690,N_11296,N_11318);
xor U11691 (N_11691,N_11280,N_11471);
xnor U11692 (N_11692,N_11324,N_11472);
xor U11693 (N_11693,N_11341,N_11342);
and U11694 (N_11694,N_11344,N_11420);
nand U11695 (N_11695,N_11391,N_11383);
xor U11696 (N_11696,N_11317,N_11466);
nor U11697 (N_11697,N_11284,N_11366);
xnor U11698 (N_11698,N_11429,N_11319);
nand U11699 (N_11699,N_11452,N_11381);
xor U11700 (N_11700,N_11418,N_11320);
and U11701 (N_11701,N_11409,N_11293);
or U11702 (N_11702,N_11396,N_11388);
nand U11703 (N_11703,N_11481,N_11446);
nor U11704 (N_11704,N_11431,N_11443);
nor U11705 (N_11705,N_11336,N_11353);
xnor U11706 (N_11706,N_11290,N_11405);
and U11707 (N_11707,N_11310,N_11488);
nand U11708 (N_11708,N_11352,N_11427);
nand U11709 (N_11709,N_11440,N_11494);
xor U11710 (N_11710,N_11288,N_11271);
nand U11711 (N_11711,N_11462,N_11406);
and U11712 (N_11712,N_11338,N_11417);
nor U11713 (N_11713,N_11373,N_11334);
nor U11714 (N_11714,N_11436,N_11338);
and U11715 (N_11715,N_11423,N_11266);
xnor U11716 (N_11716,N_11266,N_11378);
or U11717 (N_11717,N_11287,N_11267);
nor U11718 (N_11718,N_11308,N_11283);
nor U11719 (N_11719,N_11339,N_11456);
nand U11720 (N_11720,N_11279,N_11370);
or U11721 (N_11721,N_11307,N_11388);
and U11722 (N_11722,N_11492,N_11477);
nor U11723 (N_11723,N_11337,N_11402);
nor U11724 (N_11724,N_11384,N_11494);
nor U11725 (N_11725,N_11299,N_11458);
nor U11726 (N_11726,N_11488,N_11273);
xnor U11727 (N_11727,N_11461,N_11395);
and U11728 (N_11728,N_11463,N_11440);
or U11729 (N_11729,N_11396,N_11455);
nand U11730 (N_11730,N_11261,N_11256);
or U11731 (N_11731,N_11284,N_11367);
xnor U11732 (N_11732,N_11316,N_11478);
or U11733 (N_11733,N_11456,N_11328);
or U11734 (N_11734,N_11252,N_11492);
or U11735 (N_11735,N_11342,N_11289);
and U11736 (N_11736,N_11484,N_11364);
nand U11737 (N_11737,N_11375,N_11348);
nor U11738 (N_11738,N_11333,N_11348);
or U11739 (N_11739,N_11309,N_11489);
and U11740 (N_11740,N_11341,N_11275);
nor U11741 (N_11741,N_11483,N_11477);
nand U11742 (N_11742,N_11436,N_11305);
nor U11743 (N_11743,N_11426,N_11478);
or U11744 (N_11744,N_11273,N_11376);
nand U11745 (N_11745,N_11382,N_11413);
or U11746 (N_11746,N_11470,N_11392);
or U11747 (N_11747,N_11427,N_11444);
nor U11748 (N_11748,N_11497,N_11494);
nand U11749 (N_11749,N_11414,N_11325);
and U11750 (N_11750,N_11562,N_11747);
nor U11751 (N_11751,N_11737,N_11576);
nand U11752 (N_11752,N_11678,N_11508);
nand U11753 (N_11753,N_11500,N_11661);
nand U11754 (N_11754,N_11506,N_11592);
and U11755 (N_11755,N_11726,N_11668);
xor U11756 (N_11756,N_11510,N_11734);
and U11757 (N_11757,N_11691,N_11638);
nor U11758 (N_11758,N_11512,N_11641);
and U11759 (N_11759,N_11679,N_11743);
nor U11760 (N_11760,N_11527,N_11602);
nor U11761 (N_11761,N_11636,N_11736);
nand U11762 (N_11762,N_11507,N_11700);
nor U11763 (N_11763,N_11572,N_11728);
nand U11764 (N_11764,N_11684,N_11702);
nor U11765 (N_11765,N_11729,N_11598);
nand U11766 (N_11766,N_11669,N_11676);
nand U11767 (N_11767,N_11509,N_11695);
or U11768 (N_11768,N_11670,N_11682);
and U11769 (N_11769,N_11630,N_11586);
xor U11770 (N_11770,N_11651,N_11658);
xnor U11771 (N_11771,N_11687,N_11521);
nor U11772 (N_11772,N_11574,N_11735);
nor U11773 (N_11773,N_11525,N_11552);
nand U11774 (N_11774,N_11530,N_11650);
nand U11775 (N_11775,N_11551,N_11704);
xnor U11776 (N_11776,N_11631,N_11637);
xnor U11777 (N_11777,N_11643,N_11706);
xor U11778 (N_11778,N_11590,N_11714);
and U11779 (N_11779,N_11642,N_11712);
xnor U11780 (N_11780,N_11600,N_11513);
or U11781 (N_11781,N_11559,N_11730);
and U11782 (N_11782,N_11742,N_11555);
and U11783 (N_11783,N_11583,N_11564);
xnor U11784 (N_11784,N_11522,N_11585);
nor U11785 (N_11785,N_11733,N_11595);
xor U11786 (N_11786,N_11724,N_11698);
nand U11787 (N_11787,N_11718,N_11674);
nand U11788 (N_11788,N_11705,N_11579);
xor U11789 (N_11789,N_11685,N_11648);
and U11790 (N_11790,N_11701,N_11554);
nor U11791 (N_11791,N_11548,N_11688);
nand U11792 (N_11792,N_11556,N_11645);
and U11793 (N_11793,N_11709,N_11605);
and U11794 (N_11794,N_11671,N_11569);
xnor U11795 (N_11795,N_11514,N_11596);
nand U11796 (N_11796,N_11649,N_11511);
or U11797 (N_11797,N_11640,N_11597);
nor U11798 (N_11798,N_11609,N_11577);
nand U11799 (N_11799,N_11553,N_11738);
or U11800 (N_11800,N_11599,N_11571);
nor U11801 (N_11801,N_11731,N_11518);
and U11802 (N_11802,N_11719,N_11673);
and U11803 (N_11803,N_11567,N_11607);
nor U11804 (N_11804,N_11581,N_11550);
nor U11805 (N_11805,N_11722,N_11620);
nand U11806 (N_11806,N_11739,N_11666);
and U11807 (N_11807,N_11613,N_11502);
or U11808 (N_11808,N_11561,N_11715);
and U11809 (N_11809,N_11626,N_11524);
nand U11810 (N_11810,N_11717,N_11618);
or U11811 (N_11811,N_11711,N_11660);
nand U11812 (N_11812,N_11611,N_11603);
and U11813 (N_11813,N_11628,N_11624);
and U11814 (N_11814,N_11665,N_11653);
nor U11815 (N_11815,N_11681,N_11710);
and U11816 (N_11816,N_11732,N_11632);
and U11817 (N_11817,N_11617,N_11619);
xnor U11818 (N_11818,N_11543,N_11633);
xor U11819 (N_11819,N_11708,N_11625);
or U11820 (N_11820,N_11634,N_11520);
xor U11821 (N_11821,N_11699,N_11713);
and U11822 (N_11822,N_11504,N_11565);
nor U11823 (N_11823,N_11557,N_11534);
and U11824 (N_11824,N_11696,N_11544);
xor U11825 (N_11825,N_11541,N_11536);
nand U11826 (N_11826,N_11588,N_11621);
xor U11827 (N_11827,N_11531,N_11558);
or U11828 (N_11828,N_11537,N_11675);
nor U11829 (N_11829,N_11654,N_11538);
nor U11830 (N_11830,N_11519,N_11582);
xor U11831 (N_11831,N_11601,N_11655);
xor U11832 (N_11832,N_11573,N_11545);
or U11833 (N_11833,N_11677,N_11694);
nand U11834 (N_11834,N_11746,N_11664);
xnor U11835 (N_11835,N_11744,N_11516);
or U11836 (N_11836,N_11741,N_11535);
nand U11837 (N_11837,N_11680,N_11547);
or U11838 (N_11838,N_11690,N_11652);
nor U11839 (N_11839,N_11515,N_11697);
or U11840 (N_11840,N_11542,N_11644);
and U11841 (N_11841,N_11594,N_11659);
or U11842 (N_11842,N_11627,N_11612);
nor U11843 (N_11843,N_11657,N_11745);
nor U11844 (N_11844,N_11689,N_11748);
or U11845 (N_11845,N_11686,N_11589);
and U11846 (N_11846,N_11578,N_11528);
nor U11847 (N_11847,N_11740,N_11692);
and U11848 (N_11848,N_11533,N_11584);
nand U11849 (N_11849,N_11503,N_11610);
nand U11850 (N_11850,N_11667,N_11749);
nand U11851 (N_11851,N_11635,N_11526);
or U11852 (N_11852,N_11639,N_11591);
or U11853 (N_11853,N_11656,N_11532);
nand U11854 (N_11854,N_11614,N_11560);
xnor U11855 (N_11855,N_11716,N_11549);
nand U11856 (N_11856,N_11725,N_11616);
nor U11857 (N_11857,N_11517,N_11546);
or U11858 (N_11858,N_11662,N_11563);
and U11859 (N_11859,N_11629,N_11580);
or U11860 (N_11860,N_11568,N_11505);
and U11861 (N_11861,N_11540,N_11615);
xnor U11862 (N_11862,N_11647,N_11721);
and U11863 (N_11863,N_11593,N_11672);
xnor U11864 (N_11864,N_11575,N_11646);
nand U11865 (N_11865,N_11523,N_11683);
xor U11866 (N_11866,N_11663,N_11720);
and U11867 (N_11867,N_11707,N_11604);
and U11868 (N_11868,N_11570,N_11539);
and U11869 (N_11869,N_11566,N_11727);
nor U11870 (N_11870,N_11623,N_11501);
and U11871 (N_11871,N_11606,N_11622);
nor U11872 (N_11872,N_11723,N_11693);
nor U11873 (N_11873,N_11703,N_11529);
and U11874 (N_11874,N_11608,N_11587);
xnor U11875 (N_11875,N_11573,N_11609);
and U11876 (N_11876,N_11550,N_11703);
nand U11877 (N_11877,N_11579,N_11563);
nor U11878 (N_11878,N_11737,N_11740);
or U11879 (N_11879,N_11578,N_11500);
nor U11880 (N_11880,N_11580,N_11634);
nor U11881 (N_11881,N_11519,N_11657);
and U11882 (N_11882,N_11538,N_11589);
or U11883 (N_11883,N_11698,N_11556);
xor U11884 (N_11884,N_11569,N_11532);
and U11885 (N_11885,N_11716,N_11712);
or U11886 (N_11886,N_11722,N_11697);
xor U11887 (N_11887,N_11737,N_11745);
nor U11888 (N_11888,N_11672,N_11537);
or U11889 (N_11889,N_11605,N_11628);
and U11890 (N_11890,N_11613,N_11747);
or U11891 (N_11891,N_11556,N_11737);
or U11892 (N_11892,N_11639,N_11505);
nor U11893 (N_11893,N_11692,N_11749);
nand U11894 (N_11894,N_11557,N_11525);
or U11895 (N_11895,N_11692,N_11652);
or U11896 (N_11896,N_11525,N_11633);
or U11897 (N_11897,N_11666,N_11506);
nor U11898 (N_11898,N_11685,N_11509);
xnor U11899 (N_11899,N_11518,N_11665);
xor U11900 (N_11900,N_11543,N_11566);
or U11901 (N_11901,N_11512,N_11613);
xnor U11902 (N_11902,N_11707,N_11729);
nand U11903 (N_11903,N_11656,N_11699);
nor U11904 (N_11904,N_11615,N_11569);
or U11905 (N_11905,N_11509,N_11614);
nand U11906 (N_11906,N_11684,N_11738);
nand U11907 (N_11907,N_11585,N_11573);
or U11908 (N_11908,N_11706,N_11673);
or U11909 (N_11909,N_11699,N_11727);
xnor U11910 (N_11910,N_11572,N_11603);
xnor U11911 (N_11911,N_11683,N_11567);
xor U11912 (N_11912,N_11528,N_11560);
or U11913 (N_11913,N_11590,N_11689);
xor U11914 (N_11914,N_11560,N_11537);
or U11915 (N_11915,N_11660,N_11596);
and U11916 (N_11916,N_11647,N_11642);
and U11917 (N_11917,N_11708,N_11703);
nor U11918 (N_11918,N_11595,N_11718);
or U11919 (N_11919,N_11675,N_11520);
nand U11920 (N_11920,N_11665,N_11695);
nand U11921 (N_11921,N_11643,N_11524);
xnor U11922 (N_11922,N_11525,N_11651);
xor U11923 (N_11923,N_11643,N_11563);
nand U11924 (N_11924,N_11648,N_11524);
nor U11925 (N_11925,N_11702,N_11712);
or U11926 (N_11926,N_11529,N_11596);
nor U11927 (N_11927,N_11694,N_11704);
and U11928 (N_11928,N_11701,N_11574);
nand U11929 (N_11929,N_11510,N_11610);
nor U11930 (N_11930,N_11565,N_11725);
nand U11931 (N_11931,N_11706,N_11667);
nand U11932 (N_11932,N_11665,N_11610);
nand U11933 (N_11933,N_11535,N_11587);
xor U11934 (N_11934,N_11589,N_11600);
and U11935 (N_11935,N_11741,N_11633);
and U11936 (N_11936,N_11691,N_11674);
and U11937 (N_11937,N_11584,N_11534);
and U11938 (N_11938,N_11677,N_11549);
or U11939 (N_11939,N_11570,N_11659);
xnor U11940 (N_11940,N_11596,N_11707);
nor U11941 (N_11941,N_11724,N_11718);
or U11942 (N_11942,N_11582,N_11564);
and U11943 (N_11943,N_11508,N_11621);
or U11944 (N_11944,N_11618,N_11651);
and U11945 (N_11945,N_11699,N_11523);
and U11946 (N_11946,N_11737,N_11525);
nor U11947 (N_11947,N_11719,N_11597);
nand U11948 (N_11948,N_11672,N_11614);
or U11949 (N_11949,N_11502,N_11614);
or U11950 (N_11950,N_11706,N_11540);
or U11951 (N_11951,N_11700,N_11709);
nor U11952 (N_11952,N_11716,N_11568);
nor U11953 (N_11953,N_11548,N_11657);
nor U11954 (N_11954,N_11513,N_11706);
and U11955 (N_11955,N_11636,N_11613);
nand U11956 (N_11956,N_11575,N_11713);
or U11957 (N_11957,N_11597,N_11601);
nor U11958 (N_11958,N_11512,N_11637);
nand U11959 (N_11959,N_11575,N_11686);
nand U11960 (N_11960,N_11523,N_11557);
or U11961 (N_11961,N_11724,N_11645);
nor U11962 (N_11962,N_11696,N_11713);
nor U11963 (N_11963,N_11650,N_11639);
and U11964 (N_11964,N_11553,N_11689);
and U11965 (N_11965,N_11700,N_11554);
nor U11966 (N_11966,N_11707,N_11711);
nor U11967 (N_11967,N_11585,N_11730);
xor U11968 (N_11968,N_11566,N_11608);
xnor U11969 (N_11969,N_11692,N_11727);
xnor U11970 (N_11970,N_11501,N_11619);
xor U11971 (N_11971,N_11664,N_11586);
or U11972 (N_11972,N_11610,N_11738);
nand U11973 (N_11973,N_11682,N_11731);
nand U11974 (N_11974,N_11665,N_11555);
nand U11975 (N_11975,N_11711,N_11604);
xnor U11976 (N_11976,N_11581,N_11628);
xor U11977 (N_11977,N_11727,N_11688);
xnor U11978 (N_11978,N_11703,N_11634);
nor U11979 (N_11979,N_11575,N_11550);
xor U11980 (N_11980,N_11659,N_11633);
xor U11981 (N_11981,N_11564,N_11529);
nor U11982 (N_11982,N_11514,N_11679);
and U11983 (N_11983,N_11502,N_11648);
and U11984 (N_11984,N_11720,N_11530);
nand U11985 (N_11985,N_11596,N_11748);
or U11986 (N_11986,N_11616,N_11738);
nand U11987 (N_11987,N_11571,N_11587);
and U11988 (N_11988,N_11562,N_11631);
or U11989 (N_11989,N_11738,N_11565);
and U11990 (N_11990,N_11548,N_11571);
nand U11991 (N_11991,N_11609,N_11706);
or U11992 (N_11992,N_11644,N_11747);
nor U11993 (N_11993,N_11559,N_11538);
nor U11994 (N_11994,N_11736,N_11648);
and U11995 (N_11995,N_11726,N_11734);
and U11996 (N_11996,N_11682,N_11582);
nor U11997 (N_11997,N_11566,N_11519);
xnor U11998 (N_11998,N_11647,N_11551);
nand U11999 (N_11999,N_11533,N_11717);
and U12000 (N_12000,N_11885,N_11944);
nand U12001 (N_12001,N_11849,N_11994);
nor U12002 (N_12002,N_11955,N_11813);
nor U12003 (N_12003,N_11870,N_11788);
nor U12004 (N_12004,N_11847,N_11804);
and U12005 (N_12005,N_11898,N_11838);
or U12006 (N_12006,N_11853,N_11786);
and U12007 (N_12007,N_11881,N_11910);
and U12008 (N_12008,N_11753,N_11795);
xnor U12009 (N_12009,N_11907,N_11775);
or U12010 (N_12010,N_11999,N_11829);
nor U12011 (N_12011,N_11904,N_11946);
and U12012 (N_12012,N_11997,N_11842);
xnor U12013 (N_12013,N_11941,N_11961);
and U12014 (N_12014,N_11972,N_11943);
or U12015 (N_12015,N_11934,N_11773);
or U12016 (N_12016,N_11759,N_11960);
nor U12017 (N_12017,N_11976,N_11968);
xnor U12018 (N_12018,N_11835,N_11852);
nor U12019 (N_12019,N_11792,N_11769);
and U12020 (N_12020,N_11952,N_11858);
nor U12021 (N_12021,N_11823,N_11861);
and U12022 (N_12022,N_11958,N_11901);
nand U12023 (N_12023,N_11876,N_11906);
nand U12024 (N_12024,N_11819,N_11988);
and U12025 (N_12025,N_11974,N_11883);
nand U12026 (N_12026,N_11796,N_11756);
or U12027 (N_12027,N_11887,N_11772);
and U12028 (N_12028,N_11929,N_11755);
nand U12029 (N_12029,N_11874,N_11766);
xnor U12030 (N_12030,N_11857,N_11873);
or U12031 (N_12031,N_11806,N_11800);
and U12032 (N_12032,N_11754,N_11875);
or U12033 (N_12033,N_11758,N_11866);
nor U12034 (N_12034,N_11893,N_11820);
and U12035 (N_12035,N_11980,N_11880);
and U12036 (N_12036,N_11937,N_11799);
nor U12037 (N_12037,N_11839,N_11942);
nor U12038 (N_12038,N_11809,N_11831);
nor U12039 (N_12039,N_11751,N_11895);
nor U12040 (N_12040,N_11841,N_11768);
xnor U12041 (N_12041,N_11815,N_11783);
xnor U12042 (N_12042,N_11990,N_11844);
xnor U12043 (N_12043,N_11791,N_11939);
nor U12044 (N_12044,N_11957,N_11965);
and U12045 (N_12045,N_11856,N_11816);
nand U12046 (N_12046,N_11973,N_11948);
or U12047 (N_12047,N_11771,N_11921);
and U12048 (N_12048,N_11900,N_11811);
and U12049 (N_12049,N_11925,N_11863);
and U12050 (N_12050,N_11851,N_11827);
xnor U12051 (N_12051,N_11808,N_11989);
and U12052 (N_12052,N_11889,N_11764);
xor U12053 (N_12053,N_11949,N_11987);
and U12054 (N_12054,N_11963,N_11912);
or U12055 (N_12055,N_11966,N_11777);
nor U12056 (N_12056,N_11935,N_11828);
nor U12057 (N_12057,N_11862,N_11762);
nand U12058 (N_12058,N_11830,N_11860);
nor U12059 (N_12059,N_11978,N_11812);
and U12060 (N_12060,N_11867,N_11964);
and U12061 (N_12061,N_11911,N_11750);
nor U12062 (N_12062,N_11918,N_11781);
xnor U12063 (N_12063,N_11959,N_11846);
or U12064 (N_12064,N_11803,N_11878);
or U12065 (N_12065,N_11882,N_11969);
and U12066 (N_12066,N_11779,N_11919);
nor U12067 (N_12067,N_11761,N_11832);
xnor U12068 (N_12068,N_11940,N_11985);
xor U12069 (N_12069,N_11774,N_11825);
and U12070 (N_12070,N_11810,N_11932);
and U12071 (N_12071,N_11903,N_11854);
xor U12072 (N_12072,N_11787,N_11891);
and U12073 (N_12073,N_11986,N_11837);
nor U12074 (N_12074,N_11909,N_11822);
xor U12075 (N_12075,N_11938,N_11877);
nand U12076 (N_12076,N_11840,N_11872);
or U12077 (N_12077,N_11782,N_11814);
and U12078 (N_12078,N_11834,N_11767);
and U12079 (N_12079,N_11884,N_11890);
xor U12080 (N_12080,N_11996,N_11992);
nand U12081 (N_12081,N_11780,N_11776);
nand U12082 (N_12082,N_11982,N_11864);
nand U12083 (N_12083,N_11802,N_11798);
and U12084 (N_12084,N_11926,N_11850);
nor U12085 (N_12085,N_11924,N_11896);
and U12086 (N_12086,N_11905,N_11848);
nand U12087 (N_12087,N_11894,N_11833);
or U12088 (N_12088,N_11923,N_11855);
nand U12089 (N_12089,N_11778,N_11975);
nor U12090 (N_12090,N_11865,N_11908);
or U12091 (N_12091,N_11826,N_11981);
or U12092 (N_12092,N_11836,N_11763);
xor U12093 (N_12093,N_11794,N_11953);
nand U12094 (N_12094,N_11869,N_11995);
nand U12095 (N_12095,N_11807,N_11821);
nand U12096 (N_12096,N_11993,N_11817);
nand U12097 (N_12097,N_11962,N_11752);
or U12098 (N_12098,N_11984,N_11845);
nand U12099 (N_12099,N_11971,N_11914);
nor U12100 (N_12100,N_11897,N_11805);
xor U12101 (N_12101,N_11868,N_11928);
and U12102 (N_12102,N_11760,N_11917);
xor U12103 (N_12103,N_11991,N_11859);
and U12104 (N_12104,N_11801,N_11902);
and U12105 (N_12105,N_11797,N_11931);
or U12106 (N_12106,N_11979,N_11983);
nand U12107 (N_12107,N_11793,N_11977);
nor U12108 (N_12108,N_11954,N_11930);
nand U12109 (N_12109,N_11947,N_11945);
nand U12110 (N_12110,N_11770,N_11790);
xnor U12111 (N_12111,N_11956,N_11888);
xnor U12112 (N_12112,N_11892,N_11998);
nor U12113 (N_12113,N_11922,N_11933);
nor U12114 (N_12114,N_11765,N_11879);
nand U12115 (N_12115,N_11784,N_11913);
xnor U12116 (N_12116,N_11967,N_11936);
and U12117 (N_12117,N_11950,N_11915);
or U12118 (N_12118,N_11970,N_11757);
or U12119 (N_12119,N_11824,N_11916);
nor U12120 (N_12120,N_11927,N_11899);
xor U12121 (N_12121,N_11789,N_11843);
nand U12122 (N_12122,N_11920,N_11886);
or U12123 (N_12123,N_11818,N_11785);
and U12124 (N_12124,N_11871,N_11951);
and U12125 (N_12125,N_11845,N_11797);
nor U12126 (N_12126,N_11842,N_11951);
or U12127 (N_12127,N_11751,N_11987);
xor U12128 (N_12128,N_11779,N_11847);
xor U12129 (N_12129,N_11751,N_11859);
or U12130 (N_12130,N_11835,N_11780);
xor U12131 (N_12131,N_11868,N_11937);
nor U12132 (N_12132,N_11755,N_11826);
nand U12133 (N_12133,N_11996,N_11893);
xnor U12134 (N_12134,N_11991,N_11806);
xnor U12135 (N_12135,N_11853,N_11947);
nand U12136 (N_12136,N_11895,N_11843);
and U12137 (N_12137,N_11977,N_11936);
xor U12138 (N_12138,N_11810,N_11895);
and U12139 (N_12139,N_11962,N_11926);
nor U12140 (N_12140,N_11918,N_11990);
or U12141 (N_12141,N_11927,N_11906);
or U12142 (N_12142,N_11976,N_11792);
and U12143 (N_12143,N_11866,N_11977);
and U12144 (N_12144,N_11944,N_11890);
nor U12145 (N_12145,N_11785,N_11867);
nand U12146 (N_12146,N_11786,N_11921);
nand U12147 (N_12147,N_11753,N_11866);
and U12148 (N_12148,N_11778,N_11981);
and U12149 (N_12149,N_11993,N_11938);
or U12150 (N_12150,N_11998,N_11962);
nor U12151 (N_12151,N_11874,N_11850);
nand U12152 (N_12152,N_11792,N_11761);
nor U12153 (N_12153,N_11817,N_11946);
nand U12154 (N_12154,N_11924,N_11819);
or U12155 (N_12155,N_11857,N_11877);
nand U12156 (N_12156,N_11926,N_11973);
nor U12157 (N_12157,N_11930,N_11819);
nor U12158 (N_12158,N_11930,N_11886);
xor U12159 (N_12159,N_11952,N_11824);
and U12160 (N_12160,N_11819,N_11865);
nor U12161 (N_12161,N_11911,N_11899);
nand U12162 (N_12162,N_11887,N_11981);
xor U12163 (N_12163,N_11954,N_11894);
or U12164 (N_12164,N_11986,N_11783);
or U12165 (N_12165,N_11830,N_11912);
and U12166 (N_12166,N_11925,N_11883);
xnor U12167 (N_12167,N_11978,N_11979);
or U12168 (N_12168,N_11973,N_11887);
or U12169 (N_12169,N_11954,N_11837);
or U12170 (N_12170,N_11883,N_11773);
and U12171 (N_12171,N_11784,N_11994);
nor U12172 (N_12172,N_11876,N_11891);
xnor U12173 (N_12173,N_11877,N_11774);
nor U12174 (N_12174,N_11952,N_11975);
or U12175 (N_12175,N_11788,N_11898);
and U12176 (N_12176,N_11903,N_11806);
and U12177 (N_12177,N_11900,N_11877);
nand U12178 (N_12178,N_11869,N_11831);
or U12179 (N_12179,N_11932,N_11835);
nor U12180 (N_12180,N_11772,N_11771);
nand U12181 (N_12181,N_11770,N_11754);
nor U12182 (N_12182,N_11904,N_11771);
nor U12183 (N_12183,N_11809,N_11932);
xor U12184 (N_12184,N_11790,N_11951);
or U12185 (N_12185,N_11830,N_11858);
and U12186 (N_12186,N_11783,N_11889);
xnor U12187 (N_12187,N_11779,N_11921);
nand U12188 (N_12188,N_11810,N_11811);
or U12189 (N_12189,N_11811,N_11827);
or U12190 (N_12190,N_11938,N_11900);
xor U12191 (N_12191,N_11882,N_11757);
and U12192 (N_12192,N_11979,N_11925);
and U12193 (N_12193,N_11777,N_11820);
and U12194 (N_12194,N_11983,N_11894);
and U12195 (N_12195,N_11858,N_11995);
and U12196 (N_12196,N_11984,N_11959);
or U12197 (N_12197,N_11909,N_11847);
xor U12198 (N_12198,N_11779,N_11977);
and U12199 (N_12199,N_11766,N_11962);
xnor U12200 (N_12200,N_11764,N_11766);
xor U12201 (N_12201,N_11848,N_11961);
nand U12202 (N_12202,N_11857,N_11810);
or U12203 (N_12203,N_11771,N_11943);
xor U12204 (N_12204,N_11937,N_11801);
xnor U12205 (N_12205,N_11786,N_11957);
nand U12206 (N_12206,N_11826,N_11874);
or U12207 (N_12207,N_11984,N_11975);
xnor U12208 (N_12208,N_11929,N_11765);
xor U12209 (N_12209,N_11894,N_11969);
and U12210 (N_12210,N_11942,N_11785);
nor U12211 (N_12211,N_11842,N_11775);
nor U12212 (N_12212,N_11817,N_11955);
nor U12213 (N_12213,N_11929,N_11845);
and U12214 (N_12214,N_11780,N_11909);
and U12215 (N_12215,N_11861,N_11878);
and U12216 (N_12216,N_11782,N_11881);
xnor U12217 (N_12217,N_11960,N_11815);
nor U12218 (N_12218,N_11860,N_11907);
xor U12219 (N_12219,N_11894,N_11985);
xor U12220 (N_12220,N_11913,N_11855);
or U12221 (N_12221,N_11873,N_11770);
or U12222 (N_12222,N_11866,N_11867);
and U12223 (N_12223,N_11836,N_11949);
nand U12224 (N_12224,N_11811,N_11844);
and U12225 (N_12225,N_11922,N_11877);
nor U12226 (N_12226,N_11990,N_11927);
xnor U12227 (N_12227,N_11790,N_11935);
xor U12228 (N_12228,N_11940,N_11846);
xnor U12229 (N_12229,N_11936,N_11859);
nand U12230 (N_12230,N_11792,N_11891);
nand U12231 (N_12231,N_11804,N_11819);
nor U12232 (N_12232,N_11782,N_11950);
and U12233 (N_12233,N_11994,N_11775);
nor U12234 (N_12234,N_11891,N_11861);
nor U12235 (N_12235,N_11841,N_11972);
nor U12236 (N_12236,N_11833,N_11872);
nand U12237 (N_12237,N_11959,N_11914);
nand U12238 (N_12238,N_11978,N_11843);
and U12239 (N_12239,N_11844,N_11788);
nor U12240 (N_12240,N_11944,N_11791);
or U12241 (N_12241,N_11839,N_11951);
nor U12242 (N_12242,N_11864,N_11876);
nand U12243 (N_12243,N_11876,N_11981);
nand U12244 (N_12244,N_11975,N_11965);
xnor U12245 (N_12245,N_11960,N_11854);
nor U12246 (N_12246,N_11826,N_11966);
or U12247 (N_12247,N_11911,N_11883);
and U12248 (N_12248,N_11958,N_11862);
nand U12249 (N_12249,N_11946,N_11801);
nand U12250 (N_12250,N_12019,N_12207);
nand U12251 (N_12251,N_12031,N_12092);
or U12252 (N_12252,N_12076,N_12221);
and U12253 (N_12253,N_12114,N_12223);
and U12254 (N_12254,N_12184,N_12150);
nor U12255 (N_12255,N_12053,N_12090);
or U12256 (N_12256,N_12145,N_12132);
and U12257 (N_12257,N_12008,N_12035);
xor U12258 (N_12258,N_12119,N_12083);
xor U12259 (N_12259,N_12183,N_12203);
nor U12260 (N_12260,N_12111,N_12208);
xnor U12261 (N_12261,N_12056,N_12196);
and U12262 (N_12262,N_12023,N_12147);
nor U12263 (N_12263,N_12153,N_12093);
nand U12264 (N_12264,N_12185,N_12170);
nand U12265 (N_12265,N_12206,N_12245);
nor U12266 (N_12266,N_12131,N_12099);
or U12267 (N_12267,N_12158,N_12188);
nor U12268 (N_12268,N_12074,N_12211);
nand U12269 (N_12269,N_12108,N_12159);
or U12270 (N_12270,N_12059,N_12015);
nand U12271 (N_12271,N_12115,N_12103);
and U12272 (N_12272,N_12167,N_12040);
xor U12273 (N_12273,N_12061,N_12126);
or U12274 (N_12274,N_12200,N_12064);
xnor U12275 (N_12275,N_12179,N_12052);
or U12276 (N_12276,N_12045,N_12144);
nand U12277 (N_12277,N_12063,N_12229);
nor U12278 (N_12278,N_12189,N_12146);
xnor U12279 (N_12279,N_12133,N_12072);
nor U12280 (N_12280,N_12033,N_12138);
nor U12281 (N_12281,N_12181,N_12065);
and U12282 (N_12282,N_12136,N_12050);
xor U12283 (N_12283,N_12148,N_12178);
xnor U12284 (N_12284,N_12001,N_12006);
and U12285 (N_12285,N_12247,N_12209);
xor U12286 (N_12286,N_12112,N_12215);
xor U12287 (N_12287,N_12149,N_12244);
xnor U12288 (N_12288,N_12192,N_12029);
nor U12289 (N_12289,N_12000,N_12172);
or U12290 (N_12290,N_12041,N_12037);
xnor U12291 (N_12291,N_12141,N_12049);
or U12292 (N_12292,N_12080,N_12177);
nand U12293 (N_12293,N_12113,N_12225);
nor U12294 (N_12294,N_12171,N_12060);
and U12295 (N_12295,N_12154,N_12216);
and U12296 (N_12296,N_12166,N_12084);
nand U12297 (N_12297,N_12106,N_12193);
xnor U12298 (N_12298,N_12066,N_12213);
or U12299 (N_12299,N_12165,N_12226);
nand U12300 (N_12300,N_12249,N_12231);
and U12301 (N_12301,N_12034,N_12068);
xnor U12302 (N_12302,N_12224,N_12143);
nor U12303 (N_12303,N_12004,N_12218);
or U12304 (N_12304,N_12161,N_12139);
and U12305 (N_12305,N_12051,N_12246);
nor U12306 (N_12306,N_12077,N_12030);
or U12307 (N_12307,N_12107,N_12152);
or U12308 (N_12308,N_12122,N_12009);
nor U12309 (N_12309,N_12240,N_12238);
or U12310 (N_12310,N_12239,N_12021);
nor U12311 (N_12311,N_12017,N_12058);
nor U12312 (N_12312,N_12094,N_12130);
nor U12313 (N_12313,N_12027,N_12191);
or U12314 (N_12314,N_12101,N_12222);
or U12315 (N_12315,N_12014,N_12214);
nor U12316 (N_12316,N_12012,N_12228);
nand U12317 (N_12317,N_12095,N_12118);
xor U12318 (N_12318,N_12085,N_12007);
nand U12319 (N_12319,N_12024,N_12142);
and U12320 (N_12320,N_12232,N_12109);
and U12321 (N_12321,N_12135,N_12176);
and U12322 (N_12322,N_12087,N_12174);
nand U12323 (N_12323,N_12018,N_12230);
nor U12324 (N_12324,N_12089,N_12005);
nor U12325 (N_12325,N_12233,N_12079);
nand U12326 (N_12326,N_12102,N_12204);
and U12327 (N_12327,N_12182,N_12201);
and U12328 (N_12328,N_12104,N_12157);
and U12329 (N_12329,N_12198,N_12160);
xnor U12330 (N_12330,N_12235,N_12243);
nand U12331 (N_12331,N_12124,N_12036);
nor U12332 (N_12332,N_12010,N_12129);
nand U12333 (N_12333,N_12241,N_12190);
xnor U12334 (N_12334,N_12237,N_12162);
nor U12335 (N_12335,N_12180,N_12151);
xor U12336 (N_12336,N_12038,N_12047);
and U12337 (N_12337,N_12046,N_12199);
nand U12338 (N_12338,N_12073,N_12120);
nand U12339 (N_12339,N_12210,N_12123);
or U12340 (N_12340,N_12098,N_12082);
nor U12341 (N_12341,N_12219,N_12140);
or U12342 (N_12342,N_12054,N_12220);
nand U12343 (N_12343,N_12013,N_12091);
and U12344 (N_12344,N_12197,N_12105);
or U12345 (N_12345,N_12128,N_12202);
or U12346 (N_12346,N_12227,N_12088);
nand U12347 (N_12347,N_12003,N_12057);
nand U12348 (N_12348,N_12086,N_12062);
nand U12349 (N_12349,N_12097,N_12195);
nor U12350 (N_12350,N_12134,N_12028);
xnor U12351 (N_12351,N_12187,N_12164);
nor U12352 (N_12352,N_12067,N_12039);
and U12353 (N_12353,N_12169,N_12055);
and U12354 (N_12354,N_12070,N_12026);
nand U12355 (N_12355,N_12194,N_12069);
nor U12356 (N_12356,N_12156,N_12081);
and U12357 (N_12357,N_12186,N_12096);
xnor U12358 (N_12358,N_12075,N_12100);
xor U12359 (N_12359,N_12242,N_12234);
nor U12360 (N_12360,N_12110,N_12125);
nor U12361 (N_12361,N_12020,N_12236);
nand U12362 (N_12362,N_12048,N_12116);
or U12363 (N_12363,N_12155,N_12212);
or U12364 (N_12364,N_12205,N_12022);
xnor U12365 (N_12365,N_12025,N_12173);
or U12366 (N_12366,N_12002,N_12016);
or U12367 (N_12367,N_12137,N_12127);
or U12368 (N_12368,N_12168,N_12117);
xnor U12369 (N_12369,N_12071,N_12217);
nand U12370 (N_12370,N_12175,N_12248);
or U12371 (N_12371,N_12121,N_12044);
nor U12372 (N_12372,N_12011,N_12078);
nand U12373 (N_12373,N_12042,N_12163);
or U12374 (N_12374,N_12032,N_12043);
and U12375 (N_12375,N_12085,N_12143);
nand U12376 (N_12376,N_12055,N_12097);
xor U12377 (N_12377,N_12212,N_12209);
xnor U12378 (N_12378,N_12224,N_12174);
nor U12379 (N_12379,N_12071,N_12122);
xor U12380 (N_12380,N_12072,N_12179);
nand U12381 (N_12381,N_12246,N_12091);
nor U12382 (N_12382,N_12231,N_12214);
xor U12383 (N_12383,N_12170,N_12071);
xor U12384 (N_12384,N_12222,N_12148);
xor U12385 (N_12385,N_12034,N_12097);
xor U12386 (N_12386,N_12177,N_12227);
nand U12387 (N_12387,N_12233,N_12019);
or U12388 (N_12388,N_12077,N_12001);
and U12389 (N_12389,N_12028,N_12191);
nand U12390 (N_12390,N_12218,N_12156);
xnor U12391 (N_12391,N_12185,N_12068);
or U12392 (N_12392,N_12048,N_12078);
xnor U12393 (N_12393,N_12083,N_12009);
nor U12394 (N_12394,N_12022,N_12047);
or U12395 (N_12395,N_12188,N_12180);
or U12396 (N_12396,N_12179,N_12217);
and U12397 (N_12397,N_12193,N_12206);
nand U12398 (N_12398,N_12213,N_12225);
and U12399 (N_12399,N_12088,N_12131);
or U12400 (N_12400,N_12204,N_12225);
and U12401 (N_12401,N_12156,N_12064);
nor U12402 (N_12402,N_12206,N_12054);
and U12403 (N_12403,N_12102,N_12162);
nor U12404 (N_12404,N_12071,N_12236);
xor U12405 (N_12405,N_12033,N_12166);
and U12406 (N_12406,N_12052,N_12006);
nand U12407 (N_12407,N_12241,N_12055);
nor U12408 (N_12408,N_12235,N_12000);
nand U12409 (N_12409,N_12070,N_12039);
and U12410 (N_12410,N_12241,N_12185);
xor U12411 (N_12411,N_12224,N_12021);
nor U12412 (N_12412,N_12019,N_12037);
xnor U12413 (N_12413,N_12111,N_12057);
and U12414 (N_12414,N_12035,N_12032);
and U12415 (N_12415,N_12161,N_12086);
and U12416 (N_12416,N_12058,N_12011);
nor U12417 (N_12417,N_12181,N_12120);
or U12418 (N_12418,N_12114,N_12175);
and U12419 (N_12419,N_12008,N_12011);
and U12420 (N_12420,N_12075,N_12151);
nand U12421 (N_12421,N_12006,N_12099);
xnor U12422 (N_12422,N_12228,N_12158);
or U12423 (N_12423,N_12018,N_12178);
xor U12424 (N_12424,N_12206,N_12026);
or U12425 (N_12425,N_12201,N_12124);
nand U12426 (N_12426,N_12025,N_12133);
xnor U12427 (N_12427,N_12089,N_12153);
or U12428 (N_12428,N_12178,N_12130);
and U12429 (N_12429,N_12117,N_12175);
nand U12430 (N_12430,N_12105,N_12123);
xnor U12431 (N_12431,N_12092,N_12125);
nor U12432 (N_12432,N_12228,N_12039);
nor U12433 (N_12433,N_12048,N_12074);
nand U12434 (N_12434,N_12131,N_12136);
nor U12435 (N_12435,N_12054,N_12157);
and U12436 (N_12436,N_12104,N_12125);
and U12437 (N_12437,N_12078,N_12038);
nand U12438 (N_12438,N_12095,N_12222);
or U12439 (N_12439,N_12037,N_12130);
or U12440 (N_12440,N_12230,N_12078);
nand U12441 (N_12441,N_12175,N_12160);
and U12442 (N_12442,N_12093,N_12041);
xnor U12443 (N_12443,N_12127,N_12041);
nand U12444 (N_12444,N_12030,N_12043);
xor U12445 (N_12445,N_12170,N_12070);
nor U12446 (N_12446,N_12167,N_12226);
or U12447 (N_12447,N_12098,N_12247);
nor U12448 (N_12448,N_12101,N_12168);
or U12449 (N_12449,N_12080,N_12185);
or U12450 (N_12450,N_12051,N_12129);
or U12451 (N_12451,N_12139,N_12236);
or U12452 (N_12452,N_12219,N_12045);
or U12453 (N_12453,N_12055,N_12213);
nand U12454 (N_12454,N_12100,N_12116);
nor U12455 (N_12455,N_12037,N_12206);
xor U12456 (N_12456,N_12005,N_12116);
xor U12457 (N_12457,N_12045,N_12137);
nand U12458 (N_12458,N_12121,N_12055);
or U12459 (N_12459,N_12014,N_12067);
or U12460 (N_12460,N_12125,N_12216);
and U12461 (N_12461,N_12151,N_12239);
xnor U12462 (N_12462,N_12150,N_12145);
and U12463 (N_12463,N_12223,N_12160);
and U12464 (N_12464,N_12047,N_12009);
nand U12465 (N_12465,N_12070,N_12108);
nand U12466 (N_12466,N_12021,N_12079);
and U12467 (N_12467,N_12201,N_12087);
xnor U12468 (N_12468,N_12171,N_12156);
or U12469 (N_12469,N_12156,N_12005);
nand U12470 (N_12470,N_12016,N_12126);
or U12471 (N_12471,N_12085,N_12111);
and U12472 (N_12472,N_12199,N_12201);
xnor U12473 (N_12473,N_12068,N_12165);
nor U12474 (N_12474,N_12133,N_12248);
and U12475 (N_12475,N_12049,N_12080);
and U12476 (N_12476,N_12054,N_12216);
or U12477 (N_12477,N_12004,N_12162);
xnor U12478 (N_12478,N_12017,N_12042);
or U12479 (N_12479,N_12106,N_12068);
nand U12480 (N_12480,N_12238,N_12227);
and U12481 (N_12481,N_12005,N_12249);
and U12482 (N_12482,N_12113,N_12064);
and U12483 (N_12483,N_12207,N_12120);
or U12484 (N_12484,N_12035,N_12125);
nor U12485 (N_12485,N_12020,N_12048);
xnor U12486 (N_12486,N_12092,N_12085);
or U12487 (N_12487,N_12042,N_12125);
and U12488 (N_12488,N_12104,N_12184);
xor U12489 (N_12489,N_12211,N_12003);
or U12490 (N_12490,N_12233,N_12039);
nor U12491 (N_12491,N_12037,N_12167);
nor U12492 (N_12492,N_12249,N_12190);
nand U12493 (N_12493,N_12120,N_12074);
and U12494 (N_12494,N_12213,N_12038);
and U12495 (N_12495,N_12147,N_12135);
and U12496 (N_12496,N_12099,N_12153);
and U12497 (N_12497,N_12071,N_12040);
or U12498 (N_12498,N_12168,N_12249);
or U12499 (N_12499,N_12130,N_12066);
xor U12500 (N_12500,N_12252,N_12447);
and U12501 (N_12501,N_12493,N_12456);
nand U12502 (N_12502,N_12475,N_12414);
xor U12503 (N_12503,N_12365,N_12441);
nand U12504 (N_12504,N_12410,N_12304);
nand U12505 (N_12505,N_12359,N_12257);
or U12506 (N_12506,N_12490,N_12299);
and U12507 (N_12507,N_12318,N_12491);
nand U12508 (N_12508,N_12273,N_12339);
nor U12509 (N_12509,N_12377,N_12366);
or U12510 (N_12510,N_12262,N_12483);
and U12511 (N_12511,N_12401,N_12451);
nand U12512 (N_12512,N_12425,N_12400);
nand U12513 (N_12513,N_12322,N_12361);
nor U12514 (N_12514,N_12353,N_12297);
xnor U12515 (N_12515,N_12427,N_12474);
xnor U12516 (N_12516,N_12268,N_12415);
or U12517 (N_12517,N_12409,N_12394);
nor U12518 (N_12518,N_12323,N_12423);
and U12519 (N_12519,N_12419,N_12298);
nor U12520 (N_12520,N_12387,N_12476);
nor U12521 (N_12521,N_12312,N_12358);
nand U12522 (N_12522,N_12471,N_12311);
and U12523 (N_12523,N_12424,N_12272);
and U12524 (N_12524,N_12284,N_12346);
xor U12525 (N_12525,N_12464,N_12340);
nand U12526 (N_12526,N_12363,N_12412);
nor U12527 (N_12527,N_12496,N_12289);
or U12528 (N_12528,N_12319,N_12329);
and U12529 (N_12529,N_12397,N_12437);
nor U12530 (N_12530,N_12482,N_12351);
xor U12531 (N_12531,N_12477,N_12270);
nor U12532 (N_12532,N_12416,N_12458);
nand U12533 (N_12533,N_12435,N_12372);
and U12534 (N_12534,N_12269,N_12436);
nand U12535 (N_12535,N_12281,N_12385);
xor U12536 (N_12536,N_12306,N_12497);
nor U12537 (N_12537,N_12379,N_12429);
nand U12538 (N_12538,N_12278,N_12440);
or U12539 (N_12539,N_12328,N_12466);
nor U12540 (N_12540,N_12388,N_12448);
and U12541 (N_12541,N_12454,N_12347);
or U12542 (N_12542,N_12367,N_12399);
and U12543 (N_12543,N_12384,N_12260);
nor U12544 (N_12544,N_12364,N_12258);
and U12545 (N_12545,N_12489,N_12283);
nand U12546 (N_12546,N_12277,N_12295);
and U12547 (N_12547,N_12398,N_12468);
xnor U12548 (N_12548,N_12461,N_12368);
and U12549 (N_12549,N_12370,N_12444);
xnor U12550 (N_12550,N_12354,N_12293);
nand U12551 (N_12551,N_12263,N_12287);
nand U12552 (N_12552,N_12313,N_12405);
and U12553 (N_12553,N_12264,N_12335);
xor U12554 (N_12554,N_12487,N_12465);
xor U12555 (N_12555,N_12406,N_12307);
and U12556 (N_12556,N_12422,N_12479);
xor U12557 (N_12557,N_12314,N_12256);
and U12558 (N_12558,N_12325,N_12395);
and U12559 (N_12559,N_12420,N_12334);
nor U12560 (N_12560,N_12426,N_12430);
or U12561 (N_12561,N_12338,N_12250);
nor U12562 (N_12562,N_12373,N_12499);
or U12563 (N_12563,N_12342,N_12467);
and U12564 (N_12564,N_12291,N_12402);
and U12565 (N_12565,N_12371,N_12492);
xnor U12566 (N_12566,N_12376,N_12431);
nor U12567 (N_12567,N_12341,N_12393);
and U12568 (N_12568,N_12383,N_12472);
xnor U12569 (N_12569,N_12326,N_12271);
xnor U12570 (N_12570,N_12288,N_12421);
and U12571 (N_12571,N_12438,N_12344);
xnor U12572 (N_12572,N_12362,N_12469);
or U12573 (N_12573,N_12337,N_12348);
or U12574 (N_12574,N_12254,N_12375);
and U12575 (N_12575,N_12434,N_12290);
nand U12576 (N_12576,N_12350,N_12349);
or U12577 (N_12577,N_12336,N_12411);
or U12578 (N_12578,N_12305,N_12282);
and U12579 (N_12579,N_12428,N_12478);
nor U12580 (N_12580,N_12452,N_12386);
nor U12581 (N_12581,N_12494,N_12296);
nand U12582 (N_12582,N_12484,N_12463);
nand U12583 (N_12583,N_12408,N_12392);
nand U12584 (N_12584,N_12450,N_12374);
or U12585 (N_12585,N_12253,N_12321);
or U12586 (N_12586,N_12396,N_12470);
xor U12587 (N_12587,N_12378,N_12407);
xnor U12588 (N_12588,N_12433,N_12275);
nand U12589 (N_12589,N_12389,N_12455);
or U12590 (N_12590,N_12259,N_12357);
or U12591 (N_12591,N_12360,N_12315);
nor U12592 (N_12592,N_12418,N_12330);
nand U12593 (N_12593,N_12453,N_12301);
nand U12594 (N_12594,N_12279,N_12300);
nor U12595 (N_12595,N_12324,N_12443);
or U12596 (N_12596,N_12309,N_12286);
nor U12597 (N_12597,N_12473,N_12462);
or U12598 (N_12598,N_12345,N_12403);
or U12599 (N_12599,N_12486,N_12310);
xnor U12600 (N_12600,N_12303,N_12261);
nor U12601 (N_12601,N_12308,N_12317);
nor U12602 (N_12602,N_12356,N_12343);
xnor U12603 (N_12603,N_12457,N_12413);
nand U12604 (N_12604,N_12276,N_12380);
or U12605 (N_12605,N_12274,N_12495);
and U12606 (N_12606,N_12391,N_12332);
xnor U12607 (N_12607,N_12352,N_12302);
or U12608 (N_12608,N_12449,N_12266);
nor U12609 (N_12609,N_12316,N_12285);
nand U12610 (N_12610,N_12480,N_12381);
xnor U12611 (N_12611,N_12481,N_12432);
nand U12612 (N_12612,N_12439,N_12251);
xor U12613 (N_12613,N_12404,N_12446);
and U12614 (N_12614,N_12327,N_12369);
and U12615 (N_12615,N_12382,N_12355);
xor U12616 (N_12616,N_12280,N_12417);
or U12617 (N_12617,N_12498,N_12488);
nor U12618 (N_12618,N_12292,N_12333);
or U12619 (N_12619,N_12265,N_12445);
nor U12620 (N_12620,N_12267,N_12442);
nor U12621 (N_12621,N_12320,N_12255);
xor U12622 (N_12622,N_12485,N_12294);
xor U12623 (N_12623,N_12331,N_12390);
xor U12624 (N_12624,N_12460,N_12459);
or U12625 (N_12625,N_12375,N_12252);
nor U12626 (N_12626,N_12270,N_12271);
nor U12627 (N_12627,N_12457,N_12462);
and U12628 (N_12628,N_12263,N_12315);
and U12629 (N_12629,N_12330,N_12443);
nand U12630 (N_12630,N_12369,N_12308);
nor U12631 (N_12631,N_12382,N_12404);
or U12632 (N_12632,N_12424,N_12285);
nor U12633 (N_12633,N_12454,N_12498);
and U12634 (N_12634,N_12358,N_12431);
or U12635 (N_12635,N_12305,N_12475);
and U12636 (N_12636,N_12370,N_12465);
xor U12637 (N_12637,N_12254,N_12363);
and U12638 (N_12638,N_12332,N_12333);
and U12639 (N_12639,N_12255,N_12464);
nand U12640 (N_12640,N_12397,N_12434);
or U12641 (N_12641,N_12432,N_12409);
or U12642 (N_12642,N_12441,N_12424);
nand U12643 (N_12643,N_12358,N_12311);
nor U12644 (N_12644,N_12340,N_12253);
or U12645 (N_12645,N_12498,N_12410);
nand U12646 (N_12646,N_12286,N_12323);
nor U12647 (N_12647,N_12454,N_12449);
or U12648 (N_12648,N_12261,N_12381);
nand U12649 (N_12649,N_12256,N_12391);
nor U12650 (N_12650,N_12353,N_12377);
or U12651 (N_12651,N_12323,N_12420);
or U12652 (N_12652,N_12404,N_12285);
and U12653 (N_12653,N_12415,N_12294);
nor U12654 (N_12654,N_12395,N_12413);
xnor U12655 (N_12655,N_12293,N_12251);
xor U12656 (N_12656,N_12336,N_12344);
and U12657 (N_12657,N_12303,N_12476);
or U12658 (N_12658,N_12303,N_12485);
xor U12659 (N_12659,N_12404,N_12411);
or U12660 (N_12660,N_12381,N_12368);
nor U12661 (N_12661,N_12453,N_12331);
xnor U12662 (N_12662,N_12443,N_12480);
nor U12663 (N_12663,N_12482,N_12321);
and U12664 (N_12664,N_12379,N_12365);
nand U12665 (N_12665,N_12442,N_12438);
xnor U12666 (N_12666,N_12358,N_12413);
or U12667 (N_12667,N_12325,N_12364);
nor U12668 (N_12668,N_12382,N_12477);
or U12669 (N_12669,N_12394,N_12484);
nand U12670 (N_12670,N_12373,N_12359);
nand U12671 (N_12671,N_12352,N_12457);
nor U12672 (N_12672,N_12254,N_12311);
xnor U12673 (N_12673,N_12430,N_12397);
nand U12674 (N_12674,N_12312,N_12268);
and U12675 (N_12675,N_12485,N_12468);
nor U12676 (N_12676,N_12476,N_12378);
and U12677 (N_12677,N_12459,N_12309);
and U12678 (N_12678,N_12379,N_12271);
and U12679 (N_12679,N_12252,N_12475);
and U12680 (N_12680,N_12341,N_12385);
nand U12681 (N_12681,N_12349,N_12353);
and U12682 (N_12682,N_12309,N_12448);
and U12683 (N_12683,N_12250,N_12323);
xnor U12684 (N_12684,N_12390,N_12351);
or U12685 (N_12685,N_12387,N_12335);
and U12686 (N_12686,N_12339,N_12445);
nor U12687 (N_12687,N_12291,N_12464);
xor U12688 (N_12688,N_12483,N_12346);
nor U12689 (N_12689,N_12284,N_12494);
nor U12690 (N_12690,N_12312,N_12446);
xnor U12691 (N_12691,N_12347,N_12430);
xnor U12692 (N_12692,N_12440,N_12451);
or U12693 (N_12693,N_12251,N_12398);
and U12694 (N_12694,N_12297,N_12250);
or U12695 (N_12695,N_12363,N_12481);
or U12696 (N_12696,N_12346,N_12430);
nor U12697 (N_12697,N_12307,N_12262);
nand U12698 (N_12698,N_12368,N_12350);
and U12699 (N_12699,N_12456,N_12282);
or U12700 (N_12700,N_12258,N_12458);
xnor U12701 (N_12701,N_12382,N_12428);
xnor U12702 (N_12702,N_12468,N_12445);
nor U12703 (N_12703,N_12437,N_12283);
or U12704 (N_12704,N_12304,N_12324);
nor U12705 (N_12705,N_12291,N_12445);
xnor U12706 (N_12706,N_12479,N_12352);
or U12707 (N_12707,N_12473,N_12388);
and U12708 (N_12708,N_12392,N_12352);
nand U12709 (N_12709,N_12480,N_12258);
nand U12710 (N_12710,N_12434,N_12377);
and U12711 (N_12711,N_12463,N_12407);
xor U12712 (N_12712,N_12461,N_12399);
nand U12713 (N_12713,N_12257,N_12486);
nand U12714 (N_12714,N_12303,N_12304);
and U12715 (N_12715,N_12355,N_12284);
and U12716 (N_12716,N_12293,N_12494);
xnor U12717 (N_12717,N_12296,N_12465);
and U12718 (N_12718,N_12483,N_12272);
or U12719 (N_12719,N_12386,N_12489);
nand U12720 (N_12720,N_12497,N_12473);
nor U12721 (N_12721,N_12494,N_12266);
nand U12722 (N_12722,N_12453,N_12271);
nor U12723 (N_12723,N_12268,N_12486);
xor U12724 (N_12724,N_12418,N_12408);
and U12725 (N_12725,N_12406,N_12498);
nor U12726 (N_12726,N_12384,N_12475);
or U12727 (N_12727,N_12348,N_12442);
xor U12728 (N_12728,N_12437,N_12347);
or U12729 (N_12729,N_12334,N_12283);
and U12730 (N_12730,N_12433,N_12303);
nand U12731 (N_12731,N_12448,N_12338);
nand U12732 (N_12732,N_12256,N_12264);
xnor U12733 (N_12733,N_12311,N_12420);
xnor U12734 (N_12734,N_12435,N_12253);
or U12735 (N_12735,N_12390,N_12342);
and U12736 (N_12736,N_12322,N_12328);
and U12737 (N_12737,N_12459,N_12267);
xor U12738 (N_12738,N_12303,N_12357);
or U12739 (N_12739,N_12493,N_12310);
xor U12740 (N_12740,N_12420,N_12489);
nor U12741 (N_12741,N_12467,N_12297);
nand U12742 (N_12742,N_12314,N_12399);
and U12743 (N_12743,N_12283,N_12291);
nor U12744 (N_12744,N_12348,N_12422);
nor U12745 (N_12745,N_12428,N_12451);
xor U12746 (N_12746,N_12335,N_12409);
and U12747 (N_12747,N_12346,N_12260);
xnor U12748 (N_12748,N_12313,N_12493);
or U12749 (N_12749,N_12328,N_12446);
xnor U12750 (N_12750,N_12676,N_12687);
and U12751 (N_12751,N_12598,N_12626);
nand U12752 (N_12752,N_12670,N_12613);
nor U12753 (N_12753,N_12673,N_12570);
nand U12754 (N_12754,N_12719,N_12678);
or U12755 (N_12755,N_12520,N_12715);
nand U12756 (N_12756,N_12631,N_12500);
and U12757 (N_12757,N_12659,N_12674);
or U12758 (N_12758,N_12623,N_12664);
xnor U12759 (N_12759,N_12711,N_12616);
xor U12760 (N_12760,N_12541,N_12528);
nor U12761 (N_12761,N_12727,N_12524);
and U12762 (N_12762,N_12635,N_12648);
and U12763 (N_12763,N_12621,N_12696);
and U12764 (N_12764,N_12606,N_12557);
nor U12765 (N_12765,N_12505,N_12547);
nand U12766 (N_12766,N_12747,N_12587);
or U12767 (N_12767,N_12698,N_12543);
nand U12768 (N_12768,N_12633,N_12539);
nor U12769 (N_12769,N_12605,N_12739);
nand U12770 (N_12770,N_12681,N_12562);
and U12771 (N_12771,N_12749,N_12634);
xnor U12772 (N_12772,N_12572,N_12685);
nand U12773 (N_12773,N_12584,N_12502);
and U12774 (N_12774,N_12590,N_12571);
xnor U12775 (N_12775,N_12545,N_12740);
nor U12776 (N_12776,N_12675,N_12551);
xor U12777 (N_12777,N_12736,N_12503);
and U12778 (N_12778,N_12684,N_12732);
and U12779 (N_12779,N_12507,N_12531);
nand U12780 (N_12780,N_12511,N_12733);
nor U12781 (N_12781,N_12591,N_12576);
nand U12782 (N_12782,N_12529,N_12712);
xor U12783 (N_12783,N_12692,N_12512);
xor U12784 (N_12784,N_12699,N_12513);
nand U12785 (N_12785,N_12730,N_12700);
and U12786 (N_12786,N_12628,N_12564);
or U12787 (N_12787,N_12627,N_12560);
nor U12788 (N_12788,N_12637,N_12565);
xor U12789 (N_12789,N_12599,N_12672);
nand U12790 (N_12790,N_12552,N_12629);
and U12791 (N_12791,N_12726,N_12636);
and U12792 (N_12792,N_12604,N_12706);
nand U12793 (N_12793,N_12583,N_12538);
nor U12794 (N_12794,N_12669,N_12640);
nor U12795 (N_12795,N_12581,N_12718);
xnor U12796 (N_12796,N_12555,N_12745);
or U12797 (N_12797,N_12653,N_12592);
xnor U12798 (N_12798,N_12559,N_12625);
and U12799 (N_12799,N_12519,N_12533);
or U12800 (N_12800,N_12611,N_12721);
and U12801 (N_12801,N_12716,N_12697);
xor U12802 (N_12802,N_12647,N_12680);
or U12803 (N_12803,N_12738,N_12723);
nor U12804 (N_12804,N_12509,N_12523);
and U12805 (N_12805,N_12683,N_12608);
or U12806 (N_12806,N_12580,N_12556);
nor U12807 (N_12807,N_12662,N_12702);
nor U12808 (N_12808,N_12667,N_12663);
or U12809 (N_12809,N_12582,N_12546);
nand U12810 (N_12810,N_12731,N_12708);
nor U12811 (N_12811,N_12530,N_12563);
xor U12812 (N_12812,N_12554,N_12518);
nand U12813 (N_12813,N_12639,N_12506);
and U12814 (N_12814,N_12722,N_12594);
and U12815 (N_12815,N_12661,N_12713);
nand U12816 (N_12816,N_12666,N_12578);
nand U12817 (N_12817,N_12561,N_12588);
nand U12818 (N_12818,N_12532,N_12642);
and U12819 (N_12819,N_12612,N_12746);
xnor U12820 (N_12820,N_12579,N_12501);
xnor U12821 (N_12821,N_12617,N_12682);
nand U12822 (N_12822,N_12693,N_12744);
or U12823 (N_12823,N_12724,N_12595);
nor U12824 (N_12824,N_12568,N_12553);
nand U12825 (N_12825,N_12743,N_12650);
and U12826 (N_12826,N_12707,N_12609);
xnor U12827 (N_12827,N_12655,N_12527);
nor U12828 (N_12828,N_12610,N_12549);
and U12829 (N_12829,N_12624,N_12607);
or U12830 (N_12830,N_12548,N_12589);
xnor U12831 (N_12831,N_12646,N_12710);
and U12832 (N_12832,N_12689,N_12622);
xnor U12833 (N_12833,N_12603,N_12586);
or U12834 (N_12834,N_12656,N_12615);
nor U12835 (N_12835,N_12614,N_12645);
and U12836 (N_12836,N_12695,N_12654);
or U12837 (N_12837,N_12575,N_12686);
or U12838 (N_12838,N_12665,N_12735);
and U12839 (N_12839,N_12644,N_12522);
nand U12840 (N_12840,N_12597,N_12585);
and U12841 (N_12841,N_12643,N_12688);
xnor U12842 (N_12842,N_12558,N_12671);
nor U12843 (N_12843,N_12652,N_12714);
xnor U12844 (N_12844,N_12510,N_12737);
nand U12845 (N_12845,N_12630,N_12540);
nand U12846 (N_12846,N_12720,N_12573);
nand U12847 (N_12847,N_12704,N_12668);
nor U12848 (N_12848,N_12638,N_12658);
and U12849 (N_12849,N_12729,N_12728);
and U12850 (N_12850,N_12517,N_12618);
nand U12851 (N_12851,N_12550,N_12593);
or U12852 (N_12852,N_12537,N_12725);
and U12853 (N_12853,N_12632,N_12734);
or U12854 (N_12854,N_12709,N_12619);
or U12855 (N_12855,N_12651,N_12742);
nand U12856 (N_12856,N_12748,N_12515);
and U12857 (N_12857,N_12504,N_12521);
nor U12858 (N_12858,N_12703,N_12536);
or U12859 (N_12859,N_12717,N_12535);
and U12860 (N_12860,N_12567,N_12600);
nand U12861 (N_12861,N_12690,N_12660);
nor U12862 (N_12862,N_12574,N_12514);
xor U12863 (N_12863,N_12566,N_12596);
or U12864 (N_12864,N_12542,N_12516);
and U12865 (N_12865,N_12701,N_12569);
nand U12866 (N_12866,N_12544,N_12534);
xor U12867 (N_12867,N_12601,N_12525);
nand U12868 (N_12868,N_12705,N_12602);
and U12869 (N_12869,N_12526,N_12691);
and U12870 (N_12870,N_12677,N_12741);
nand U12871 (N_12871,N_12620,N_12679);
or U12872 (N_12872,N_12649,N_12694);
nand U12873 (N_12873,N_12508,N_12641);
xor U12874 (N_12874,N_12657,N_12577);
and U12875 (N_12875,N_12548,N_12508);
nand U12876 (N_12876,N_12626,N_12592);
and U12877 (N_12877,N_12726,N_12599);
or U12878 (N_12878,N_12528,N_12590);
nor U12879 (N_12879,N_12562,N_12650);
xor U12880 (N_12880,N_12579,N_12525);
xnor U12881 (N_12881,N_12683,N_12623);
or U12882 (N_12882,N_12668,N_12592);
xnor U12883 (N_12883,N_12665,N_12597);
and U12884 (N_12884,N_12649,N_12722);
or U12885 (N_12885,N_12647,N_12656);
or U12886 (N_12886,N_12518,N_12645);
nor U12887 (N_12887,N_12731,N_12632);
or U12888 (N_12888,N_12652,N_12639);
nor U12889 (N_12889,N_12536,N_12552);
nand U12890 (N_12890,N_12654,N_12674);
xnor U12891 (N_12891,N_12617,N_12659);
nand U12892 (N_12892,N_12738,N_12560);
nand U12893 (N_12893,N_12737,N_12622);
nand U12894 (N_12894,N_12671,N_12580);
xor U12895 (N_12895,N_12520,N_12527);
and U12896 (N_12896,N_12598,N_12580);
and U12897 (N_12897,N_12729,N_12569);
nand U12898 (N_12898,N_12570,N_12528);
xor U12899 (N_12899,N_12637,N_12730);
or U12900 (N_12900,N_12575,N_12608);
nand U12901 (N_12901,N_12681,N_12649);
or U12902 (N_12902,N_12696,N_12597);
xor U12903 (N_12903,N_12509,N_12571);
nand U12904 (N_12904,N_12661,N_12613);
or U12905 (N_12905,N_12559,N_12525);
and U12906 (N_12906,N_12512,N_12573);
nor U12907 (N_12907,N_12540,N_12638);
or U12908 (N_12908,N_12656,N_12718);
and U12909 (N_12909,N_12590,N_12706);
xnor U12910 (N_12910,N_12573,N_12679);
xor U12911 (N_12911,N_12669,N_12510);
xor U12912 (N_12912,N_12617,N_12688);
nand U12913 (N_12913,N_12618,N_12544);
nand U12914 (N_12914,N_12543,N_12504);
or U12915 (N_12915,N_12612,N_12565);
and U12916 (N_12916,N_12516,N_12529);
nand U12917 (N_12917,N_12707,N_12562);
and U12918 (N_12918,N_12662,N_12653);
or U12919 (N_12919,N_12589,N_12649);
or U12920 (N_12920,N_12525,N_12605);
or U12921 (N_12921,N_12735,N_12588);
and U12922 (N_12922,N_12519,N_12637);
nand U12923 (N_12923,N_12545,N_12529);
nand U12924 (N_12924,N_12615,N_12729);
nand U12925 (N_12925,N_12706,N_12609);
or U12926 (N_12926,N_12618,N_12554);
and U12927 (N_12927,N_12617,N_12558);
xnor U12928 (N_12928,N_12699,N_12597);
nor U12929 (N_12929,N_12658,N_12632);
nand U12930 (N_12930,N_12602,N_12506);
and U12931 (N_12931,N_12536,N_12578);
nor U12932 (N_12932,N_12656,N_12596);
nor U12933 (N_12933,N_12749,N_12508);
or U12934 (N_12934,N_12636,N_12671);
nor U12935 (N_12935,N_12515,N_12604);
nand U12936 (N_12936,N_12507,N_12691);
or U12937 (N_12937,N_12723,N_12531);
or U12938 (N_12938,N_12730,N_12630);
nand U12939 (N_12939,N_12741,N_12502);
xor U12940 (N_12940,N_12523,N_12562);
nand U12941 (N_12941,N_12521,N_12578);
xnor U12942 (N_12942,N_12688,N_12700);
and U12943 (N_12943,N_12597,N_12725);
nand U12944 (N_12944,N_12508,N_12659);
nand U12945 (N_12945,N_12525,N_12626);
or U12946 (N_12946,N_12748,N_12535);
nor U12947 (N_12947,N_12548,N_12526);
and U12948 (N_12948,N_12731,N_12605);
and U12949 (N_12949,N_12685,N_12510);
or U12950 (N_12950,N_12512,N_12660);
xor U12951 (N_12951,N_12689,N_12655);
nand U12952 (N_12952,N_12633,N_12598);
xor U12953 (N_12953,N_12519,N_12616);
nor U12954 (N_12954,N_12585,N_12535);
and U12955 (N_12955,N_12532,N_12547);
and U12956 (N_12956,N_12692,N_12597);
xor U12957 (N_12957,N_12712,N_12576);
nand U12958 (N_12958,N_12654,N_12635);
nand U12959 (N_12959,N_12748,N_12739);
or U12960 (N_12960,N_12747,N_12657);
or U12961 (N_12961,N_12562,N_12661);
nand U12962 (N_12962,N_12543,N_12744);
and U12963 (N_12963,N_12578,N_12619);
or U12964 (N_12964,N_12659,N_12536);
or U12965 (N_12965,N_12523,N_12617);
or U12966 (N_12966,N_12582,N_12654);
and U12967 (N_12967,N_12503,N_12518);
and U12968 (N_12968,N_12573,N_12653);
or U12969 (N_12969,N_12675,N_12701);
xnor U12970 (N_12970,N_12575,N_12536);
nor U12971 (N_12971,N_12720,N_12585);
nand U12972 (N_12972,N_12507,N_12535);
nand U12973 (N_12973,N_12568,N_12629);
and U12974 (N_12974,N_12715,N_12638);
nor U12975 (N_12975,N_12687,N_12654);
and U12976 (N_12976,N_12506,N_12680);
nor U12977 (N_12977,N_12603,N_12679);
and U12978 (N_12978,N_12553,N_12563);
xor U12979 (N_12979,N_12700,N_12548);
nor U12980 (N_12980,N_12726,N_12666);
nor U12981 (N_12981,N_12503,N_12538);
and U12982 (N_12982,N_12571,N_12691);
nand U12983 (N_12983,N_12748,N_12620);
nor U12984 (N_12984,N_12621,N_12626);
xnor U12985 (N_12985,N_12745,N_12720);
or U12986 (N_12986,N_12633,N_12715);
xor U12987 (N_12987,N_12653,N_12689);
or U12988 (N_12988,N_12555,N_12561);
and U12989 (N_12989,N_12701,N_12533);
and U12990 (N_12990,N_12514,N_12551);
and U12991 (N_12991,N_12635,N_12542);
nor U12992 (N_12992,N_12565,N_12583);
and U12993 (N_12993,N_12645,N_12551);
xor U12994 (N_12994,N_12686,N_12608);
or U12995 (N_12995,N_12560,N_12639);
nand U12996 (N_12996,N_12720,N_12522);
xor U12997 (N_12997,N_12641,N_12747);
nand U12998 (N_12998,N_12566,N_12684);
nor U12999 (N_12999,N_12542,N_12556);
or U13000 (N_13000,N_12935,N_12947);
or U13001 (N_13001,N_12827,N_12834);
or U13002 (N_13002,N_12898,N_12972);
and U13003 (N_13003,N_12760,N_12755);
or U13004 (N_13004,N_12783,N_12857);
nand U13005 (N_13005,N_12881,N_12767);
xnor U13006 (N_13006,N_12911,N_12975);
or U13007 (N_13007,N_12756,N_12776);
or U13008 (N_13008,N_12766,N_12978);
xnor U13009 (N_13009,N_12893,N_12835);
nand U13010 (N_13010,N_12809,N_12877);
nor U13011 (N_13011,N_12851,N_12949);
nand U13012 (N_13012,N_12904,N_12885);
xnor U13013 (N_13013,N_12837,N_12791);
nand U13014 (N_13014,N_12995,N_12805);
nor U13015 (N_13015,N_12982,N_12894);
xnor U13016 (N_13016,N_12924,N_12757);
nand U13017 (N_13017,N_12840,N_12925);
nand U13018 (N_13018,N_12933,N_12994);
nand U13019 (N_13019,N_12909,N_12774);
and U13020 (N_13020,N_12944,N_12957);
or U13021 (N_13021,N_12966,N_12931);
or U13022 (N_13022,N_12872,N_12792);
nand U13023 (N_13023,N_12770,N_12910);
nor U13024 (N_13024,N_12915,N_12960);
xor U13025 (N_13025,N_12919,N_12846);
nand U13026 (N_13026,N_12812,N_12977);
and U13027 (N_13027,N_12815,N_12901);
xor U13028 (N_13028,N_12779,N_12876);
or U13029 (N_13029,N_12921,N_12914);
or U13030 (N_13030,N_12956,N_12789);
xnor U13031 (N_13031,N_12917,N_12762);
and U13032 (N_13032,N_12985,N_12942);
or U13033 (N_13033,N_12861,N_12821);
xor U13034 (N_13034,N_12764,N_12996);
or U13035 (N_13035,N_12855,N_12831);
nand U13036 (N_13036,N_12973,N_12858);
nor U13037 (N_13037,N_12988,N_12822);
or U13038 (N_13038,N_12899,N_12871);
xnor U13039 (N_13039,N_12900,N_12806);
and U13040 (N_13040,N_12912,N_12907);
nand U13041 (N_13041,N_12884,N_12948);
nand U13042 (N_13042,N_12984,N_12986);
and U13043 (N_13043,N_12974,N_12759);
or U13044 (N_13044,N_12798,N_12813);
xnor U13045 (N_13045,N_12775,N_12926);
or U13046 (N_13046,N_12810,N_12784);
xor U13047 (N_13047,N_12879,N_12790);
and U13048 (N_13048,N_12889,N_12826);
nor U13049 (N_13049,N_12954,N_12820);
nand U13050 (N_13050,N_12838,N_12953);
or U13051 (N_13051,N_12916,N_12895);
and U13052 (N_13052,N_12869,N_12753);
and U13053 (N_13053,N_12998,N_12941);
nand U13054 (N_13054,N_12788,N_12999);
and U13055 (N_13055,N_12839,N_12906);
and U13056 (N_13056,N_12829,N_12795);
nand U13057 (N_13057,N_12945,N_12955);
nor U13058 (N_13058,N_12754,N_12856);
and U13059 (N_13059,N_12797,N_12842);
and U13060 (N_13060,N_12801,N_12825);
xnor U13061 (N_13061,N_12865,N_12993);
or U13062 (N_13062,N_12934,N_12800);
nand U13063 (N_13063,N_12782,N_12940);
or U13064 (N_13064,N_12905,N_12892);
nor U13065 (N_13065,N_12841,N_12918);
and U13066 (N_13066,N_12991,N_12823);
and U13067 (N_13067,N_12878,N_12781);
nor U13068 (N_13068,N_12751,N_12969);
or U13069 (N_13069,N_12963,N_12853);
xor U13070 (N_13070,N_12794,N_12785);
xor U13071 (N_13071,N_12828,N_12964);
nand U13072 (N_13072,N_12952,N_12943);
and U13073 (N_13073,N_12928,N_12890);
and U13074 (N_13074,N_12843,N_12807);
xor U13075 (N_13075,N_12814,N_12780);
xor U13076 (N_13076,N_12971,N_12833);
xnor U13077 (N_13077,N_12946,N_12987);
nand U13078 (N_13078,N_12970,N_12875);
nand U13079 (N_13079,N_12886,N_12818);
nand U13080 (N_13080,N_12832,N_12824);
nor U13081 (N_13081,N_12854,N_12950);
xor U13082 (N_13082,N_12967,N_12938);
nand U13083 (N_13083,N_12903,N_12796);
xnor U13084 (N_13084,N_12777,N_12787);
nand U13085 (N_13085,N_12868,N_12896);
nand U13086 (N_13086,N_12852,N_12962);
nor U13087 (N_13087,N_12836,N_12930);
and U13088 (N_13088,N_12761,N_12765);
or U13089 (N_13089,N_12864,N_12873);
nor U13090 (N_13090,N_12819,N_12990);
nor U13091 (N_13091,N_12763,N_12768);
or U13092 (N_13092,N_12908,N_12887);
nand U13093 (N_13093,N_12750,N_12965);
nand U13094 (N_13094,N_12830,N_12803);
and U13095 (N_13095,N_12923,N_12927);
nand U13096 (N_13096,N_12773,N_12811);
xor U13097 (N_13097,N_12920,N_12983);
and U13098 (N_13098,N_12844,N_12808);
and U13099 (N_13099,N_12867,N_12932);
nand U13100 (N_13100,N_12981,N_12848);
or U13101 (N_13101,N_12997,N_12888);
xor U13102 (N_13102,N_12793,N_12863);
and U13103 (N_13103,N_12913,N_12870);
or U13104 (N_13104,N_12936,N_12771);
and U13105 (N_13105,N_12980,N_12786);
or U13106 (N_13106,N_12976,N_12860);
and U13107 (N_13107,N_12847,N_12897);
nor U13108 (N_13108,N_12850,N_12937);
and U13109 (N_13109,N_12859,N_12845);
xor U13110 (N_13110,N_12802,N_12758);
nor U13111 (N_13111,N_12880,N_12939);
and U13112 (N_13112,N_12817,N_12922);
or U13113 (N_13113,N_12979,N_12874);
and U13114 (N_13114,N_12769,N_12799);
or U13115 (N_13115,N_12816,N_12968);
nor U13116 (N_13116,N_12891,N_12902);
and U13117 (N_13117,N_12883,N_12849);
nor U13118 (N_13118,N_12862,N_12959);
xnor U13119 (N_13119,N_12772,N_12804);
nand U13120 (N_13120,N_12958,N_12882);
nand U13121 (N_13121,N_12866,N_12992);
nand U13122 (N_13122,N_12778,N_12951);
nor U13123 (N_13123,N_12929,N_12989);
or U13124 (N_13124,N_12752,N_12961);
xnor U13125 (N_13125,N_12937,N_12830);
xnor U13126 (N_13126,N_12977,N_12864);
xor U13127 (N_13127,N_12891,N_12878);
or U13128 (N_13128,N_12806,N_12878);
xnor U13129 (N_13129,N_12803,N_12908);
or U13130 (N_13130,N_12863,N_12755);
xnor U13131 (N_13131,N_12992,N_12900);
xor U13132 (N_13132,N_12769,N_12937);
nor U13133 (N_13133,N_12800,N_12912);
or U13134 (N_13134,N_12972,N_12788);
and U13135 (N_13135,N_12765,N_12796);
nor U13136 (N_13136,N_12868,N_12764);
or U13137 (N_13137,N_12827,N_12794);
nand U13138 (N_13138,N_12948,N_12927);
and U13139 (N_13139,N_12884,N_12786);
or U13140 (N_13140,N_12901,N_12828);
nor U13141 (N_13141,N_12950,N_12755);
or U13142 (N_13142,N_12764,N_12843);
or U13143 (N_13143,N_12872,N_12791);
and U13144 (N_13144,N_12776,N_12897);
nand U13145 (N_13145,N_12907,N_12831);
or U13146 (N_13146,N_12969,N_12974);
or U13147 (N_13147,N_12928,N_12832);
xnor U13148 (N_13148,N_12770,N_12943);
xor U13149 (N_13149,N_12839,N_12751);
nand U13150 (N_13150,N_12812,N_12814);
nor U13151 (N_13151,N_12786,N_12848);
xor U13152 (N_13152,N_12796,N_12984);
xor U13153 (N_13153,N_12937,N_12853);
and U13154 (N_13154,N_12794,N_12952);
and U13155 (N_13155,N_12991,N_12801);
xnor U13156 (N_13156,N_12832,N_12920);
nor U13157 (N_13157,N_12816,N_12984);
or U13158 (N_13158,N_12937,N_12969);
xor U13159 (N_13159,N_12821,N_12936);
or U13160 (N_13160,N_12792,N_12826);
xnor U13161 (N_13161,N_12906,N_12925);
nand U13162 (N_13162,N_12796,N_12959);
or U13163 (N_13163,N_12862,N_12807);
nand U13164 (N_13164,N_12873,N_12792);
or U13165 (N_13165,N_12807,N_12887);
or U13166 (N_13166,N_12776,N_12774);
and U13167 (N_13167,N_12863,N_12915);
nand U13168 (N_13168,N_12857,N_12959);
xnor U13169 (N_13169,N_12768,N_12914);
xnor U13170 (N_13170,N_12980,N_12890);
xor U13171 (N_13171,N_12886,N_12982);
nor U13172 (N_13172,N_12848,N_12756);
and U13173 (N_13173,N_12849,N_12808);
nand U13174 (N_13174,N_12761,N_12767);
xor U13175 (N_13175,N_12938,N_12863);
or U13176 (N_13176,N_12997,N_12921);
nand U13177 (N_13177,N_12846,N_12962);
and U13178 (N_13178,N_12833,N_12885);
or U13179 (N_13179,N_12988,N_12865);
xor U13180 (N_13180,N_12999,N_12925);
nor U13181 (N_13181,N_12843,N_12766);
nor U13182 (N_13182,N_12925,N_12824);
nand U13183 (N_13183,N_12900,N_12865);
nor U13184 (N_13184,N_12755,N_12908);
xnor U13185 (N_13185,N_12858,N_12763);
and U13186 (N_13186,N_12842,N_12762);
xor U13187 (N_13187,N_12963,N_12884);
or U13188 (N_13188,N_12902,N_12774);
or U13189 (N_13189,N_12904,N_12957);
and U13190 (N_13190,N_12866,N_12851);
nor U13191 (N_13191,N_12982,N_12996);
xor U13192 (N_13192,N_12921,N_12947);
and U13193 (N_13193,N_12806,N_12890);
or U13194 (N_13194,N_12818,N_12899);
xnor U13195 (N_13195,N_12854,N_12843);
nand U13196 (N_13196,N_12771,N_12758);
and U13197 (N_13197,N_12918,N_12857);
nand U13198 (N_13198,N_12816,N_12898);
xnor U13199 (N_13199,N_12760,N_12781);
xor U13200 (N_13200,N_12901,N_12845);
nand U13201 (N_13201,N_12852,N_12920);
and U13202 (N_13202,N_12866,N_12915);
nand U13203 (N_13203,N_12790,N_12821);
nor U13204 (N_13204,N_12833,N_12987);
nor U13205 (N_13205,N_12873,N_12978);
or U13206 (N_13206,N_12922,N_12923);
xnor U13207 (N_13207,N_12940,N_12796);
nand U13208 (N_13208,N_12864,N_12997);
or U13209 (N_13209,N_12973,N_12917);
and U13210 (N_13210,N_12786,N_12769);
xor U13211 (N_13211,N_12912,N_12808);
nand U13212 (N_13212,N_12777,N_12901);
and U13213 (N_13213,N_12903,N_12849);
xnor U13214 (N_13214,N_12904,N_12888);
nand U13215 (N_13215,N_12945,N_12939);
nand U13216 (N_13216,N_12901,N_12816);
nor U13217 (N_13217,N_12969,N_12842);
or U13218 (N_13218,N_12886,N_12783);
nand U13219 (N_13219,N_12761,N_12816);
and U13220 (N_13220,N_12977,N_12833);
nand U13221 (N_13221,N_12910,N_12781);
and U13222 (N_13222,N_12954,N_12962);
nor U13223 (N_13223,N_12934,N_12942);
xnor U13224 (N_13224,N_12832,N_12913);
or U13225 (N_13225,N_12796,N_12999);
or U13226 (N_13226,N_12994,N_12974);
nand U13227 (N_13227,N_12964,N_12786);
xor U13228 (N_13228,N_12984,N_12880);
or U13229 (N_13229,N_12758,N_12989);
and U13230 (N_13230,N_12750,N_12839);
xor U13231 (N_13231,N_12824,N_12953);
or U13232 (N_13232,N_12994,N_12834);
xnor U13233 (N_13233,N_12751,N_12871);
or U13234 (N_13234,N_12861,N_12794);
and U13235 (N_13235,N_12855,N_12851);
nand U13236 (N_13236,N_12928,N_12996);
and U13237 (N_13237,N_12937,N_12807);
nor U13238 (N_13238,N_12916,N_12790);
nor U13239 (N_13239,N_12798,N_12812);
or U13240 (N_13240,N_12751,N_12892);
nor U13241 (N_13241,N_12820,N_12997);
nor U13242 (N_13242,N_12953,N_12814);
nand U13243 (N_13243,N_12983,N_12804);
and U13244 (N_13244,N_12958,N_12835);
nand U13245 (N_13245,N_12904,N_12890);
xor U13246 (N_13246,N_12812,N_12875);
nand U13247 (N_13247,N_12852,N_12921);
and U13248 (N_13248,N_12825,N_12765);
nand U13249 (N_13249,N_12994,N_12815);
and U13250 (N_13250,N_13106,N_13191);
nand U13251 (N_13251,N_13245,N_13158);
and U13252 (N_13252,N_13115,N_13196);
or U13253 (N_13253,N_13183,N_13070);
or U13254 (N_13254,N_13119,N_13021);
and U13255 (N_13255,N_13233,N_13152);
nand U13256 (N_13256,N_13068,N_13050);
nand U13257 (N_13257,N_13081,N_13084);
and U13258 (N_13258,N_13020,N_13229);
and U13259 (N_13259,N_13127,N_13022);
nor U13260 (N_13260,N_13006,N_13142);
nand U13261 (N_13261,N_13216,N_13109);
nor U13262 (N_13262,N_13019,N_13210);
nand U13263 (N_13263,N_13248,N_13143);
nor U13264 (N_13264,N_13061,N_13237);
xnor U13265 (N_13265,N_13150,N_13141);
nand U13266 (N_13266,N_13186,N_13113);
or U13267 (N_13267,N_13015,N_13121);
nor U13268 (N_13268,N_13016,N_13002);
or U13269 (N_13269,N_13181,N_13165);
xnor U13270 (N_13270,N_13195,N_13083);
nand U13271 (N_13271,N_13041,N_13073);
nor U13272 (N_13272,N_13148,N_13146);
nand U13273 (N_13273,N_13036,N_13174);
nor U13274 (N_13274,N_13235,N_13076);
and U13275 (N_13275,N_13105,N_13096);
nor U13276 (N_13276,N_13088,N_13133);
nand U13277 (N_13277,N_13046,N_13167);
nand U13278 (N_13278,N_13197,N_13093);
and U13279 (N_13279,N_13193,N_13043);
and U13280 (N_13280,N_13102,N_13219);
and U13281 (N_13281,N_13222,N_13187);
and U13282 (N_13282,N_13204,N_13063);
nand U13283 (N_13283,N_13010,N_13014);
xnor U13284 (N_13284,N_13045,N_13030);
nand U13285 (N_13285,N_13129,N_13018);
nand U13286 (N_13286,N_13042,N_13132);
xnor U13287 (N_13287,N_13031,N_13244);
and U13288 (N_13288,N_13124,N_13051);
or U13289 (N_13289,N_13069,N_13159);
and U13290 (N_13290,N_13053,N_13185);
nor U13291 (N_13291,N_13044,N_13205);
nand U13292 (N_13292,N_13139,N_13226);
and U13293 (N_13293,N_13240,N_13224);
and U13294 (N_13294,N_13049,N_13190);
nor U13295 (N_13295,N_13220,N_13039);
or U13296 (N_13296,N_13172,N_13035);
or U13297 (N_13297,N_13247,N_13151);
nand U13298 (N_13298,N_13156,N_13200);
nand U13299 (N_13299,N_13178,N_13242);
and U13300 (N_13300,N_13163,N_13128);
nand U13301 (N_13301,N_13080,N_13095);
nand U13302 (N_13302,N_13176,N_13192);
nor U13303 (N_13303,N_13231,N_13234);
nor U13304 (N_13304,N_13147,N_13241);
nor U13305 (N_13305,N_13103,N_13203);
and U13306 (N_13306,N_13059,N_13225);
and U13307 (N_13307,N_13125,N_13078);
xor U13308 (N_13308,N_13120,N_13025);
xnor U13309 (N_13309,N_13038,N_13209);
nand U13310 (N_13310,N_13208,N_13004);
nor U13311 (N_13311,N_13162,N_13098);
or U13312 (N_13312,N_13087,N_13201);
or U13313 (N_13313,N_13028,N_13211);
nand U13314 (N_13314,N_13228,N_13107);
xnor U13315 (N_13315,N_13173,N_13072);
or U13316 (N_13316,N_13013,N_13111);
and U13317 (N_13317,N_13189,N_13243);
and U13318 (N_13318,N_13137,N_13180);
or U13319 (N_13319,N_13136,N_13144);
and U13320 (N_13320,N_13218,N_13024);
xor U13321 (N_13321,N_13091,N_13086);
xnor U13322 (N_13322,N_13122,N_13246);
xnor U13323 (N_13323,N_13062,N_13145);
xnor U13324 (N_13324,N_13232,N_13198);
and U13325 (N_13325,N_13037,N_13227);
and U13326 (N_13326,N_13026,N_13135);
nand U13327 (N_13327,N_13157,N_13074);
nor U13328 (N_13328,N_13118,N_13108);
nand U13329 (N_13329,N_13206,N_13090);
nand U13330 (N_13330,N_13011,N_13160);
or U13331 (N_13331,N_13239,N_13012);
nor U13332 (N_13332,N_13194,N_13065);
or U13333 (N_13333,N_13164,N_13184);
nand U13334 (N_13334,N_13008,N_13140);
nor U13335 (N_13335,N_13055,N_13238);
or U13336 (N_13336,N_13131,N_13005);
nand U13337 (N_13337,N_13077,N_13202);
nand U13338 (N_13338,N_13134,N_13123);
nor U13339 (N_13339,N_13126,N_13064);
or U13340 (N_13340,N_13213,N_13230);
xor U13341 (N_13341,N_13000,N_13215);
or U13342 (N_13342,N_13236,N_13027);
nand U13343 (N_13343,N_13168,N_13177);
nand U13344 (N_13344,N_13040,N_13085);
xor U13345 (N_13345,N_13170,N_13199);
or U13346 (N_13346,N_13112,N_13217);
or U13347 (N_13347,N_13138,N_13182);
xor U13348 (N_13348,N_13249,N_13089);
or U13349 (N_13349,N_13104,N_13188);
and U13350 (N_13350,N_13221,N_13169);
xor U13351 (N_13351,N_13056,N_13114);
and U13352 (N_13352,N_13033,N_13054);
nand U13353 (N_13353,N_13057,N_13082);
xor U13354 (N_13354,N_13101,N_13166);
or U13355 (N_13355,N_13097,N_13047);
nor U13356 (N_13356,N_13003,N_13034);
nand U13357 (N_13357,N_13116,N_13079);
nor U13358 (N_13358,N_13171,N_13075);
nand U13359 (N_13359,N_13032,N_13066);
or U13360 (N_13360,N_13110,N_13179);
nor U13361 (N_13361,N_13023,N_13212);
and U13362 (N_13362,N_13130,N_13099);
nand U13363 (N_13363,N_13058,N_13154);
or U13364 (N_13364,N_13223,N_13100);
or U13365 (N_13365,N_13175,N_13117);
or U13366 (N_13366,N_13007,N_13017);
nand U13367 (N_13367,N_13009,N_13161);
or U13368 (N_13368,N_13071,N_13029);
nand U13369 (N_13369,N_13155,N_13001);
or U13370 (N_13370,N_13052,N_13207);
or U13371 (N_13371,N_13214,N_13153);
and U13372 (N_13372,N_13092,N_13149);
nand U13373 (N_13373,N_13060,N_13094);
nand U13374 (N_13374,N_13048,N_13067);
xor U13375 (N_13375,N_13129,N_13137);
and U13376 (N_13376,N_13233,N_13232);
nor U13377 (N_13377,N_13210,N_13116);
nor U13378 (N_13378,N_13190,N_13215);
and U13379 (N_13379,N_13140,N_13069);
xor U13380 (N_13380,N_13066,N_13013);
or U13381 (N_13381,N_13192,N_13020);
nor U13382 (N_13382,N_13176,N_13179);
and U13383 (N_13383,N_13216,N_13201);
xnor U13384 (N_13384,N_13084,N_13171);
nand U13385 (N_13385,N_13005,N_13248);
and U13386 (N_13386,N_13067,N_13214);
xnor U13387 (N_13387,N_13175,N_13024);
nand U13388 (N_13388,N_13219,N_13004);
nor U13389 (N_13389,N_13041,N_13240);
nor U13390 (N_13390,N_13010,N_13024);
and U13391 (N_13391,N_13126,N_13108);
and U13392 (N_13392,N_13169,N_13228);
or U13393 (N_13393,N_13093,N_13220);
xnor U13394 (N_13394,N_13163,N_13122);
nor U13395 (N_13395,N_13135,N_13138);
nor U13396 (N_13396,N_13140,N_13216);
xor U13397 (N_13397,N_13064,N_13109);
and U13398 (N_13398,N_13236,N_13193);
xor U13399 (N_13399,N_13106,N_13075);
nor U13400 (N_13400,N_13046,N_13244);
nand U13401 (N_13401,N_13053,N_13193);
xnor U13402 (N_13402,N_13198,N_13215);
or U13403 (N_13403,N_13100,N_13132);
xnor U13404 (N_13404,N_13093,N_13219);
nand U13405 (N_13405,N_13201,N_13238);
and U13406 (N_13406,N_13238,N_13101);
xor U13407 (N_13407,N_13045,N_13001);
or U13408 (N_13408,N_13179,N_13057);
nor U13409 (N_13409,N_13134,N_13226);
or U13410 (N_13410,N_13136,N_13182);
or U13411 (N_13411,N_13209,N_13078);
nand U13412 (N_13412,N_13150,N_13076);
nand U13413 (N_13413,N_13070,N_13137);
nand U13414 (N_13414,N_13209,N_13133);
and U13415 (N_13415,N_13215,N_13007);
nand U13416 (N_13416,N_13193,N_13107);
xnor U13417 (N_13417,N_13234,N_13057);
or U13418 (N_13418,N_13200,N_13035);
xnor U13419 (N_13419,N_13239,N_13073);
xnor U13420 (N_13420,N_13238,N_13196);
and U13421 (N_13421,N_13129,N_13180);
nand U13422 (N_13422,N_13009,N_13098);
and U13423 (N_13423,N_13163,N_13235);
xnor U13424 (N_13424,N_13053,N_13141);
nor U13425 (N_13425,N_13018,N_13017);
xor U13426 (N_13426,N_13153,N_13135);
or U13427 (N_13427,N_13137,N_13241);
or U13428 (N_13428,N_13221,N_13132);
nand U13429 (N_13429,N_13043,N_13007);
and U13430 (N_13430,N_13090,N_13162);
or U13431 (N_13431,N_13247,N_13112);
xnor U13432 (N_13432,N_13011,N_13042);
xor U13433 (N_13433,N_13033,N_13003);
nor U13434 (N_13434,N_13226,N_13168);
or U13435 (N_13435,N_13200,N_13237);
xor U13436 (N_13436,N_13219,N_13106);
nand U13437 (N_13437,N_13213,N_13059);
nand U13438 (N_13438,N_13131,N_13100);
nor U13439 (N_13439,N_13171,N_13231);
xor U13440 (N_13440,N_13166,N_13214);
nand U13441 (N_13441,N_13001,N_13218);
xnor U13442 (N_13442,N_13002,N_13099);
nor U13443 (N_13443,N_13238,N_13046);
xnor U13444 (N_13444,N_13032,N_13043);
nor U13445 (N_13445,N_13048,N_13063);
xor U13446 (N_13446,N_13020,N_13054);
xnor U13447 (N_13447,N_13121,N_13102);
nor U13448 (N_13448,N_13061,N_13105);
and U13449 (N_13449,N_13150,N_13237);
xor U13450 (N_13450,N_13212,N_13051);
or U13451 (N_13451,N_13189,N_13030);
nor U13452 (N_13452,N_13215,N_13023);
xor U13453 (N_13453,N_13068,N_13117);
nor U13454 (N_13454,N_13225,N_13014);
and U13455 (N_13455,N_13184,N_13079);
and U13456 (N_13456,N_13007,N_13014);
or U13457 (N_13457,N_13120,N_13204);
and U13458 (N_13458,N_13186,N_13212);
or U13459 (N_13459,N_13081,N_13035);
and U13460 (N_13460,N_13139,N_13121);
xnor U13461 (N_13461,N_13128,N_13193);
nand U13462 (N_13462,N_13117,N_13238);
or U13463 (N_13463,N_13244,N_13212);
or U13464 (N_13464,N_13217,N_13229);
xnor U13465 (N_13465,N_13158,N_13196);
nor U13466 (N_13466,N_13089,N_13141);
nand U13467 (N_13467,N_13154,N_13107);
xnor U13468 (N_13468,N_13200,N_13000);
nand U13469 (N_13469,N_13181,N_13077);
xor U13470 (N_13470,N_13183,N_13093);
and U13471 (N_13471,N_13239,N_13023);
or U13472 (N_13472,N_13028,N_13245);
nor U13473 (N_13473,N_13065,N_13079);
nor U13474 (N_13474,N_13172,N_13153);
nand U13475 (N_13475,N_13179,N_13031);
or U13476 (N_13476,N_13142,N_13140);
nor U13477 (N_13477,N_13140,N_13070);
or U13478 (N_13478,N_13075,N_13210);
nor U13479 (N_13479,N_13107,N_13058);
nor U13480 (N_13480,N_13098,N_13002);
nor U13481 (N_13481,N_13053,N_13085);
and U13482 (N_13482,N_13191,N_13055);
and U13483 (N_13483,N_13229,N_13238);
xor U13484 (N_13484,N_13235,N_13002);
or U13485 (N_13485,N_13004,N_13181);
nor U13486 (N_13486,N_13165,N_13185);
and U13487 (N_13487,N_13092,N_13147);
and U13488 (N_13488,N_13112,N_13098);
nand U13489 (N_13489,N_13037,N_13066);
and U13490 (N_13490,N_13101,N_13007);
nor U13491 (N_13491,N_13089,N_13169);
nor U13492 (N_13492,N_13083,N_13244);
xnor U13493 (N_13493,N_13168,N_13144);
and U13494 (N_13494,N_13141,N_13028);
and U13495 (N_13495,N_13188,N_13133);
nor U13496 (N_13496,N_13017,N_13126);
nand U13497 (N_13497,N_13049,N_13003);
or U13498 (N_13498,N_13216,N_13193);
or U13499 (N_13499,N_13131,N_13237);
xor U13500 (N_13500,N_13255,N_13302);
nor U13501 (N_13501,N_13458,N_13283);
nor U13502 (N_13502,N_13471,N_13385);
xnor U13503 (N_13503,N_13331,N_13474);
or U13504 (N_13504,N_13390,N_13407);
or U13505 (N_13505,N_13461,N_13335);
nand U13506 (N_13506,N_13381,N_13483);
nand U13507 (N_13507,N_13279,N_13480);
nand U13508 (N_13508,N_13484,N_13443);
nand U13509 (N_13509,N_13432,N_13475);
or U13510 (N_13510,N_13430,N_13391);
or U13511 (N_13511,N_13415,N_13456);
and U13512 (N_13512,N_13256,N_13460);
nand U13513 (N_13513,N_13413,N_13379);
xor U13514 (N_13514,N_13463,N_13312);
nand U13515 (N_13515,N_13298,N_13394);
nand U13516 (N_13516,N_13343,N_13462);
and U13517 (N_13517,N_13285,N_13276);
and U13518 (N_13518,N_13265,N_13448);
xor U13519 (N_13519,N_13490,N_13498);
or U13520 (N_13520,N_13376,N_13465);
xor U13521 (N_13521,N_13497,N_13327);
xnor U13522 (N_13522,N_13295,N_13401);
nor U13523 (N_13523,N_13307,N_13478);
or U13524 (N_13524,N_13397,N_13297);
and U13525 (N_13525,N_13324,N_13356);
or U13526 (N_13526,N_13429,N_13425);
and U13527 (N_13527,N_13319,N_13344);
and U13528 (N_13528,N_13308,N_13272);
and U13529 (N_13529,N_13380,N_13486);
and U13530 (N_13530,N_13280,N_13291);
or U13531 (N_13531,N_13436,N_13491);
xor U13532 (N_13532,N_13284,N_13253);
or U13533 (N_13533,N_13301,N_13426);
nor U13534 (N_13534,N_13469,N_13314);
nor U13535 (N_13535,N_13468,N_13330);
xnor U13536 (N_13536,N_13420,N_13410);
nor U13537 (N_13537,N_13277,N_13346);
nand U13538 (N_13538,N_13336,N_13322);
or U13539 (N_13539,N_13325,N_13287);
or U13540 (N_13540,N_13311,N_13384);
nor U13541 (N_13541,N_13366,N_13288);
nor U13542 (N_13542,N_13364,N_13453);
or U13543 (N_13543,N_13489,N_13338);
and U13544 (N_13544,N_13306,N_13328);
or U13545 (N_13545,N_13477,N_13290);
and U13546 (N_13546,N_13270,N_13438);
nor U13547 (N_13547,N_13303,N_13359);
xor U13548 (N_13548,N_13329,N_13442);
or U13549 (N_13549,N_13423,N_13360);
nand U13550 (N_13550,N_13398,N_13345);
nand U13551 (N_13551,N_13309,N_13414);
and U13552 (N_13552,N_13485,N_13267);
nor U13553 (N_13553,N_13446,N_13395);
nand U13554 (N_13554,N_13383,N_13332);
nor U13555 (N_13555,N_13386,N_13431);
nand U13556 (N_13556,N_13358,N_13493);
nor U13557 (N_13557,N_13388,N_13282);
nand U13558 (N_13558,N_13403,N_13370);
xor U13559 (N_13559,N_13355,N_13450);
or U13560 (N_13560,N_13274,N_13447);
and U13561 (N_13561,N_13402,N_13399);
xor U13562 (N_13562,N_13252,N_13317);
and U13563 (N_13563,N_13348,N_13339);
nor U13564 (N_13564,N_13352,N_13451);
nor U13565 (N_13565,N_13393,N_13310);
xor U13566 (N_13566,N_13315,N_13496);
nand U13567 (N_13567,N_13363,N_13340);
nor U13568 (N_13568,N_13320,N_13289);
nor U13569 (N_13569,N_13378,N_13264);
nand U13570 (N_13570,N_13408,N_13300);
or U13571 (N_13571,N_13374,N_13492);
xnor U13572 (N_13572,N_13412,N_13440);
nor U13573 (N_13573,N_13495,N_13278);
nand U13574 (N_13574,N_13472,N_13433);
nand U13575 (N_13575,N_13457,N_13254);
nand U13576 (N_13576,N_13481,N_13494);
xnor U13577 (N_13577,N_13441,N_13392);
and U13578 (N_13578,N_13444,N_13350);
nor U13579 (N_13579,N_13313,N_13464);
nand U13580 (N_13580,N_13445,N_13417);
or U13581 (N_13581,N_13437,N_13353);
xnor U13582 (N_13582,N_13361,N_13449);
nand U13583 (N_13583,N_13373,N_13467);
and U13584 (N_13584,N_13422,N_13258);
and U13585 (N_13585,N_13326,N_13418);
or U13586 (N_13586,N_13427,N_13260);
nand U13587 (N_13587,N_13405,N_13263);
xor U13588 (N_13588,N_13294,N_13455);
or U13589 (N_13589,N_13488,N_13342);
and U13590 (N_13590,N_13259,N_13286);
and U13591 (N_13591,N_13337,N_13268);
or U13592 (N_13592,N_13434,N_13375);
or U13593 (N_13593,N_13357,N_13473);
xnor U13594 (N_13594,N_13305,N_13281);
or U13595 (N_13595,N_13296,N_13368);
nand U13596 (N_13596,N_13349,N_13424);
nor U13597 (N_13597,N_13257,N_13416);
xor U13598 (N_13598,N_13250,N_13251);
nand U13599 (N_13599,N_13476,N_13459);
nand U13600 (N_13600,N_13318,N_13428);
and U13601 (N_13601,N_13316,N_13411);
or U13602 (N_13602,N_13365,N_13435);
nor U13603 (N_13603,N_13499,N_13269);
and U13604 (N_13604,N_13354,N_13334);
nor U13605 (N_13605,N_13275,N_13304);
nor U13606 (N_13606,N_13369,N_13466);
and U13607 (N_13607,N_13452,N_13347);
and U13608 (N_13608,N_13273,N_13409);
nor U13609 (N_13609,N_13271,N_13293);
nor U13610 (N_13610,N_13419,N_13421);
nor U13611 (N_13611,N_13382,N_13292);
nor U13612 (N_13612,N_13404,N_13377);
xor U13613 (N_13613,N_13299,N_13479);
or U13614 (N_13614,N_13341,N_13321);
or U13615 (N_13615,N_13371,N_13454);
nor U13616 (N_13616,N_13487,N_13333);
nand U13617 (N_13617,N_13372,N_13323);
nand U13618 (N_13618,N_13396,N_13400);
or U13619 (N_13619,N_13470,N_13351);
or U13620 (N_13620,N_13266,N_13482);
nand U13621 (N_13621,N_13387,N_13439);
and U13622 (N_13622,N_13362,N_13367);
xor U13623 (N_13623,N_13389,N_13262);
nor U13624 (N_13624,N_13406,N_13261);
nand U13625 (N_13625,N_13399,N_13254);
nor U13626 (N_13626,N_13444,N_13417);
or U13627 (N_13627,N_13471,N_13383);
or U13628 (N_13628,N_13429,N_13449);
nand U13629 (N_13629,N_13392,N_13315);
and U13630 (N_13630,N_13491,N_13426);
and U13631 (N_13631,N_13268,N_13267);
and U13632 (N_13632,N_13335,N_13275);
nor U13633 (N_13633,N_13294,N_13357);
xor U13634 (N_13634,N_13463,N_13280);
nor U13635 (N_13635,N_13404,N_13320);
nand U13636 (N_13636,N_13255,N_13489);
and U13637 (N_13637,N_13433,N_13399);
or U13638 (N_13638,N_13444,N_13471);
nor U13639 (N_13639,N_13451,N_13449);
and U13640 (N_13640,N_13406,N_13430);
nand U13641 (N_13641,N_13326,N_13306);
nand U13642 (N_13642,N_13305,N_13323);
and U13643 (N_13643,N_13266,N_13282);
nor U13644 (N_13644,N_13450,N_13458);
or U13645 (N_13645,N_13382,N_13273);
or U13646 (N_13646,N_13401,N_13337);
nand U13647 (N_13647,N_13497,N_13432);
nand U13648 (N_13648,N_13336,N_13434);
nand U13649 (N_13649,N_13264,N_13268);
and U13650 (N_13650,N_13365,N_13296);
or U13651 (N_13651,N_13293,N_13291);
nand U13652 (N_13652,N_13368,N_13414);
nand U13653 (N_13653,N_13391,N_13459);
and U13654 (N_13654,N_13376,N_13483);
and U13655 (N_13655,N_13310,N_13446);
nand U13656 (N_13656,N_13454,N_13299);
nand U13657 (N_13657,N_13274,N_13298);
and U13658 (N_13658,N_13303,N_13461);
xnor U13659 (N_13659,N_13349,N_13288);
and U13660 (N_13660,N_13323,N_13368);
or U13661 (N_13661,N_13344,N_13262);
xor U13662 (N_13662,N_13272,N_13258);
or U13663 (N_13663,N_13373,N_13256);
or U13664 (N_13664,N_13419,N_13414);
xnor U13665 (N_13665,N_13429,N_13412);
xnor U13666 (N_13666,N_13440,N_13481);
and U13667 (N_13667,N_13400,N_13447);
xor U13668 (N_13668,N_13288,N_13352);
or U13669 (N_13669,N_13416,N_13489);
nor U13670 (N_13670,N_13377,N_13337);
and U13671 (N_13671,N_13407,N_13439);
nor U13672 (N_13672,N_13307,N_13272);
or U13673 (N_13673,N_13273,N_13264);
xnor U13674 (N_13674,N_13402,N_13423);
or U13675 (N_13675,N_13307,N_13255);
nand U13676 (N_13676,N_13341,N_13497);
nand U13677 (N_13677,N_13402,N_13484);
nor U13678 (N_13678,N_13383,N_13389);
or U13679 (N_13679,N_13436,N_13283);
nand U13680 (N_13680,N_13416,N_13364);
xnor U13681 (N_13681,N_13261,N_13485);
nor U13682 (N_13682,N_13364,N_13271);
nand U13683 (N_13683,N_13330,N_13425);
and U13684 (N_13684,N_13402,N_13392);
nor U13685 (N_13685,N_13378,N_13313);
and U13686 (N_13686,N_13491,N_13260);
nand U13687 (N_13687,N_13423,N_13315);
and U13688 (N_13688,N_13338,N_13479);
xnor U13689 (N_13689,N_13284,N_13296);
xor U13690 (N_13690,N_13483,N_13407);
and U13691 (N_13691,N_13482,N_13291);
xor U13692 (N_13692,N_13361,N_13438);
xor U13693 (N_13693,N_13278,N_13303);
and U13694 (N_13694,N_13486,N_13485);
and U13695 (N_13695,N_13483,N_13426);
nor U13696 (N_13696,N_13489,N_13341);
nor U13697 (N_13697,N_13449,N_13370);
nor U13698 (N_13698,N_13264,N_13335);
or U13699 (N_13699,N_13486,N_13499);
or U13700 (N_13700,N_13288,N_13312);
nand U13701 (N_13701,N_13476,N_13261);
or U13702 (N_13702,N_13317,N_13474);
nand U13703 (N_13703,N_13405,N_13392);
nor U13704 (N_13704,N_13497,N_13292);
or U13705 (N_13705,N_13300,N_13430);
nor U13706 (N_13706,N_13452,N_13323);
and U13707 (N_13707,N_13327,N_13381);
xor U13708 (N_13708,N_13444,N_13280);
and U13709 (N_13709,N_13345,N_13454);
and U13710 (N_13710,N_13252,N_13313);
nand U13711 (N_13711,N_13455,N_13253);
nor U13712 (N_13712,N_13284,N_13259);
and U13713 (N_13713,N_13451,N_13371);
nor U13714 (N_13714,N_13311,N_13392);
xnor U13715 (N_13715,N_13489,N_13473);
xnor U13716 (N_13716,N_13384,N_13302);
and U13717 (N_13717,N_13365,N_13334);
nor U13718 (N_13718,N_13323,N_13496);
nand U13719 (N_13719,N_13395,N_13268);
nor U13720 (N_13720,N_13484,N_13321);
nor U13721 (N_13721,N_13428,N_13408);
xnor U13722 (N_13722,N_13464,N_13344);
nor U13723 (N_13723,N_13289,N_13484);
and U13724 (N_13724,N_13342,N_13260);
or U13725 (N_13725,N_13459,N_13313);
and U13726 (N_13726,N_13496,N_13281);
and U13727 (N_13727,N_13395,N_13265);
xor U13728 (N_13728,N_13404,N_13281);
nor U13729 (N_13729,N_13252,N_13456);
or U13730 (N_13730,N_13429,N_13282);
nand U13731 (N_13731,N_13260,N_13437);
xor U13732 (N_13732,N_13283,N_13419);
nand U13733 (N_13733,N_13317,N_13343);
nor U13734 (N_13734,N_13349,N_13460);
xor U13735 (N_13735,N_13261,N_13293);
nand U13736 (N_13736,N_13259,N_13365);
nand U13737 (N_13737,N_13272,N_13275);
nand U13738 (N_13738,N_13402,N_13364);
nand U13739 (N_13739,N_13376,N_13283);
xnor U13740 (N_13740,N_13403,N_13287);
xor U13741 (N_13741,N_13400,N_13453);
xnor U13742 (N_13742,N_13413,N_13250);
or U13743 (N_13743,N_13273,N_13275);
or U13744 (N_13744,N_13275,N_13461);
and U13745 (N_13745,N_13339,N_13332);
or U13746 (N_13746,N_13258,N_13452);
nand U13747 (N_13747,N_13456,N_13258);
nor U13748 (N_13748,N_13274,N_13446);
or U13749 (N_13749,N_13337,N_13435);
nand U13750 (N_13750,N_13562,N_13693);
nand U13751 (N_13751,N_13600,N_13737);
nand U13752 (N_13752,N_13584,N_13530);
or U13753 (N_13753,N_13704,N_13747);
nor U13754 (N_13754,N_13654,N_13571);
and U13755 (N_13755,N_13527,N_13565);
and U13756 (N_13756,N_13507,N_13500);
nand U13757 (N_13757,N_13701,N_13731);
nor U13758 (N_13758,N_13505,N_13677);
and U13759 (N_13759,N_13687,N_13534);
and U13760 (N_13760,N_13626,N_13619);
or U13761 (N_13761,N_13724,N_13623);
xnor U13762 (N_13762,N_13707,N_13587);
or U13763 (N_13763,N_13667,N_13502);
and U13764 (N_13764,N_13618,N_13643);
xnor U13765 (N_13765,N_13617,N_13630);
and U13766 (N_13766,N_13504,N_13501);
xor U13767 (N_13767,N_13660,N_13717);
nor U13768 (N_13768,N_13729,N_13678);
or U13769 (N_13769,N_13748,N_13541);
or U13770 (N_13770,N_13674,N_13668);
and U13771 (N_13771,N_13593,N_13590);
xnor U13772 (N_13772,N_13629,N_13637);
and U13773 (N_13773,N_13620,N_13555);
and U13774 (N_13774,N_13563,N_13690);
nand U13775 (N_13775,N_13561,N_13653);
nand U13776 (N_13776,N_13546,N_13605);
nand U13777 (N_13777,N_13746,N_13734);
xnor U13778 (N_13778,N_13744,N_13708);
nor U13779 (N_13779,N_13514,N_13503);
or U13780 (N_13780,N_13518,N_13554);
or U13781 (N_13781,N_13664,N_13540);
or U13782 (N_13782,N_13588,N_13698);
xor U13783 (N_13783,N_13719,N_13604);
xor U13784 (N_13784,N_13589,N_13711);
nor U13785 (N_13785,N_13506,N_13718);
and U13786 (N_13786,N_13641,N_13728);
or U13787 (N_13787,N_13634,N_13566);
nand U13788 (N_13788,N_13696,N_13692);
nand U13789 (N_13789,N_13607,N_13697);
nor U13790 (N_13790,N_13648,N_13681);
and U13791 (N_13791,N_13713,N_13597);
nand U13792 (N_13792,N_13523,N_13666);
xor U13793 (N_13793,N_13513,N_13516);
xor U13794 (N_13794,N_13586,N_13661);
nand U13795 (N_13795,N_13663,N_13577);
or U13796 (N_13796,N_13627,N_13662);
xnor U13797 (N_13797,N_13550,N_13560);
nor U13798 (N_13798,N_13671,N_13631);
xnor U13799 (N_13799,N_13552,N_13596);
nand U13800 (N_13800,N_13695,N_13525);
xnor U13801 (N_13801,N_13712,N_13595);
or U13802 (N_13802,N_13510,N_13723);
or U13803 (N_13803,N_13675,N_13536);
xnor U13804 (N_13804,N_13710,N_13585);
nor U13805 (N_13805,N_13625,N_13749);
and U13806 (N_13806,N_13519,N_13745);
nor U13807 (N_13807,N_13572,N_13676);
xor U13808 (N_13808,N_13511,N_13573);
or U13809 (N_13809,N_13614,N_13699);
nand U13810 (N_13810,N_13644,N_13532);
and U13811 (N_13811,N_13659,N_13742);
nand U13812 (N_13812,N_13694,N_13715);
nand U13813 (N_13813,N_13683,N_13543);
nand U13814 (N_13814,N_13725,N_13741);
nor U13815 (N_13815,N_13551,N_13581);
or U13816 (N_13816,N_13743,N_13615);
or U13817 (N_13817,N_13578,N_13738);
or U13818 (N_13818,N_13642,N_13665);
nor U13819 (N_13819,N_13542,N_13733);
nor U13820 (N_13820,N_13640,N_13633);
nand U13821 (N_13821,N_13726,N_13716);
nand U13822 (N_13822,N_13545,N_13548);
or U13823 (N_13823,N_13685,N_13632);
nor U13824 (N_13824,N_13721,N_13569);
or U13825 (N_13825,N_13709,N_13740);
nor U13826 (N_13826,N_13606,N_13531);
xor U13827 (N_13827,N_13649,N_13591);
nand U13828 (N_13828,N_13651,N_13559);
nor U13829 (N_13829,N_13652,N_13672);
nor U13830 (N_13830,N_13739,N_13601);
nor U13831 (N_13831,N_13508,N_13655);
and U13832 (N_13832,N_13579,N_13736);
nand U13833 (N_13833,N_13730,N_13688);
xor U13834 (N_13834,N_13635,N_13558);
nor U13835 (N_13835,N_13557,N_13537);
or U13836 (N_13836,N_13533,N_13639);
and U13837 (N_13837,N_13610,N_13613);
nand U13838 (N_13838,N_13706,N_13650);
nand U13839 (N_13839,N_13575,N_13673);
or U13840 (N_13840,N_13526,N_13603);
xnor U13841 (N_13841,N_13509,N_13705);
nor U13842 (N_13842,N_13564,N_13628);
nand U13843 (N_13843,N_13646,N_13622);
and U13844 (N_13844,N_13602,N_13570);
nand U13845 (N_13845,N_13568,N_13679);
nand U13846 (N_13846,N_13702,N_13656);
nor U13847 (N_13847,N_13735,N_13529);
and U13848 (N_13848,N_13556,N_13645);
nor U13849 (N_13849,N_13515,N_13691);
or U13850 (N_13850,N_13520,N_13512);
nor U13851 (N_13851,N_13538,N_13657);
xor U13852 (N_13852,N_13553,N_13612);
and U13853 (N_13853,N_13720,N_13567);
nor U13854 (N_13854,N_13521,N_13700);
nand U13855 (N_13855,N_13582,N_13686);
nor U13856 (N_13856,N_13658,N_13616);
and U13857 (N_13857,N_13522,N_13689);
nor U13858 (N_13858,N_13576,N_13611);
xor U13859 (N_13859,N_13592,N_13647);
and U13860 (N_13860,N_13703,N_13682);
nand U13861 (N_13861,N_13580,N_13714);
nand U13862 (N_13862,N_13549,N_13583);
nor U13863 (N_13863,N_13574,N_13680);
or U13864 (N_13864,N_13594,N_13732);
nor U13865 (N_13865,N_13621,N_13624);
nor U13866 (N_13866,N_13528,N_13684);
or U13867 (N_13867,N_13669,N_13535);
xnor U13868 (N_13868,N_13609,N_13544);
nor U13869 (N_13869,N_13517,N_13727);
and U13870 (N_13870,N_13539,N_13722);
nor U13871 (N_13871,N_13547,N_13524);
nor U13872 (N_13872,N_13636,N_13608);
nand U13873 (N_13873,N_13598,N_13670);
xnor U13874 (N_13874,N_13638,N_13599);
nor U13875 (N_13875,N_13680,N_13685);
and U13876 (N_13876,N_13743,N_13521);
xnor U13877 (N_13877,N_13584,N_13528);
and U13878 (N_13878,N_13534,N_13725);
xnor U13879 (N_13879,N_13682,N_13681);
nand U13880 (N_13880,N_13531,N_13696);
nor U13881 (N_13881,N_13596,N_13664);
nand U13882 (N_13882,N_13511,N_13690);
nand U13883 (N_13883,N_13532,N_13731);
xnor U13884 (N_13884,N_13704,N_13611);
and U13885 (N_13885,N_13727,N_13639);
nand U13886 (N_13886,N_13659,N_13695);
nor U13887 (N_13887,N_13717,N_13724);
nor U13888 (N_13888,N_13537,N_13574);
nand U13889 (N_13889,N_13614,N_13735);
nor U13890 (N_13890,N_13682,N_13523);
nor U13891 (N_13891,N_13716,N_13529);
nor U13892 (N_13892,N_13582,N_13602);
xor U13893 (N_13893,N_13580,N_13699);
and U13894 (N_13894,N_13552,N_13741);
xor U13895 (N_13895,N_13601,N_13662);
nor U13896 (N_13896,N_13740,N_13654);
and U13897 (N_13897,N_13722,N_13713);
nand U13898 (N_13898,N_13655,N_13689);
and U13899 (N_13899,N_13509,N_13504);
or U13900 (N_13900,N_13708,N_13613);
and U13901 (N_13901,N_13678,N_13661);
nand U13902 (N_13902,N_13545,N_13535);
nand U13903 (N_13903,N_13683,N_13531);
or U13904 (N_13904,N_13600,N_13543);
nor U13905 (N_13905,N_13705,N_13653);
nor U13906 (N_13906,N_13558,N_13616);
and U13907 (N_13907,N_13659,N_13703);
xor U13908 (N_13908,N_13505,N_13522);
nor U13909 (N_13909,N_13687,N_13523);
nand U13910 (N_13910,N_13502,N_13702);
nand U13911 (N_13911,N_13635,N_13538);
and U13912 (N_13912,N_13653,N_13657);
nand U13913 (N_13913,N_13579,N_13689);
and U13914 (N_13914,N_13731,N_13728);
nand U13915 (N_13915,N_13557,N_13698);
or U13916 (N_13916,N_13742,N_13579);
nand U13917 (N_13917,N_13631,N_13732);
nor U13918 (N_13918,N_13688,N_13587);
nor U13919 (N_13919,N_13705,N_13693);
and U13920 (N_13920,N_13747,N_13683);
or U13921 (N_13921,N_13532,N_13502);
or U13922 (N_13922,N_13639,N_13714);
and U13923 (N_13923,N_13547,N_13718);
nand U13924 (N_13924,N_13534,N_13624);
xnor U13925 (N_13925,N_13590,N_13517);
nor U13926 (N_13926,N_13709,N_13632);
nor U13927 (N_13927,N_13664,N_13648);
and U13928 (N_13928,N_13557,N_13671);
and U13929 (N_13929,N_13728,N_13690);
nand U13930 (N_13930,N_13727,N_13634);
and U13931 (N_13931,N_13646,N_13588);
nor U13932 (N_13932,N_13678,N_13566);
xor U13933 (N_13933,N_13663,N_13690);
xnor U13934 (N_13934,N_13608,N_13507);
nand U13935 (N_13935,N_13522,N_13512);
nor U13936 (N_13936,N_13518,N_13648);
or U13937 (N_13937,N_13502,N_13738);
nor U13938 (N_13938,N_13538,N_13598);
and U13939 (N_13939,N_13572,N_13549);
and U13940 (N_13940,N_13537,N_13692);
or U13941 (N_13941,N_13634,N_13657);
or U13942 (N_13942,N_13622,N_13546);
or U13943 (N_13943,N_13524,N_13649);
nand U13944 (N_13944,N_13533,N_13630);
nor U13945 (N_13945,N_13685,N_13592);
or U13946 (N_13946,N_13573,N_13564);
nand U13947 (N_13947,N_13665,N_13714);
and U13948 (N_13948,N_13706,N_13530);
nor U13949 (N_13949,N_13729,N_13684);
or U13950 (N_13950,N_13721,N_13568);
or U13951 (N_13951,N_13748,N_13630);
or U13952 (N_13952,N_13575,N_13684);
nand U13953 (N_13953,N_13562,N_13626);
xnor U13954 (N_13954,N_13654,N_13570);
xnor U13955 (N_13955,N_13661,N_13631);
nand U13956 (N_13956,N_13701,N_13500);
nor U13957 (N_13957,N_13592,N_13738);
nand U13958 (N_13958,N_13650,N_13662);
and U13959 (N_13959,N_13693,N_13602);
nor U13960 (N_13960,N_13682,N_13723);
nand U13961 (N_13961,N_13566,N_13590);
nor U13962 (N_13962,N_13665,N_13591);
xor U13963 (N_13963,N_13726,N_13589);
nand U13964 (N_13964,N_13505,N_13631);
and U13965 (N_13965,N_13703,N_13741);
nand U13966 (N_13966,N_13731,N_13666);
and U13967 (N_13967,N_13560,N_13500);
and U13968 (N_13968,N_13534,N_13623);
and U13969 (N_13969,N_13662,N_13613);
or U13970 (N_13970,N_13585,N_13708);
nor U13971 (N_13971,N_13741,N_13734);
nor U13972 (N_13972,N_13708,N_13740);
nor U13973 (N_13973,N_13636,N_13583);
and U13974 (N_13974,N_13655,N_13677);
or U13975 (N_13975,N_13666,N_13739);
xnor U13976 (N_13976,N_13664,N_13600);
xor U13977 (N_13977,N_13543,N_13641);
nor U13978 (N_13978,N_13691,N_13533);
nand U13979 (N_13979,N_13705,N_13547);
nand U13980 (N_13980,N_13674,N_13630);
nor U13981 (N_13981,N_13687,N_13606);
nand U13982 (N_13982,N_13629,N_13672);
and U13983 (N_13983,N_13692,N_13562);
nand U13984 (N_13984,N_13648,N_13541);
or U13985 (N_13985,N_13604,N_13645);
and U13986 (N_13986,N_13736,N_13695);
xnor U13987 (N_13987,N_13693,N_13648);
xor U13988 (N_13988,N_13637,N_13562);
xor U13989 (N_13989,N_13547,N_13592);
xor U13990 (N_13990,N_13537,N_13630);
and U13991 (N_13991,N_13642,N_13711);
or U13992 (N_13992,N_13713,N_13686);
or U13993 (N_13993,N_13604,N_13599);
and U13994 (N_13994,N_13576,N_13543);
xor U13995 (N_13995,N_13710,N_13706);
or U13996 (N_13996,N_13663,N_13598);
and U13997 (N_13997,N_13652,N_13684);
and U13998 (N_13998,N_13624,N_13517);
or U13999 (N_13999,N_13594,N_13680);
nor U14000 (N_14000,N_13896,N_13844);
and U14001 (N_14001,N_13976,N_13824);
nand U14002 (N_14002,N_13873,N_13802);
or U14003 (N_14003,N_13855,N_13752);
and U14004 (N_14004,N_13806,N_13860);
or U14005 (N_14005,N_13960,N_13925);
or U14006 (N_14006,N_13811,N_13941);
nor U14007 (N_14007,N_13790,N_13977);
and U14008 (N_14008,N_13909,N_13780);
nor U14009 (N_14009,N_13820,N_13771);
or U14010 (N_14010,N_13927,N_13944);
nand U14011 (N_14011,N_13974,N_13767);
nor U14012 (N_14012,N_13763,N_13756);
and U14013 (N_14013,N_13893,N_13945);
and U14014 (N_14014,N_13829,N_13912);
nand U14015 (N_14015,N_13989,N_13905);
nor U14016 (N_14016,N_13879,N_13911);
nor U14017 (N_14017,N_13895,N_13922);
xor U14018 (N_14018,N_13789,N_13800);
nor U14019 (N_14019,N_13938,N_13981);
nand U14020 (N_14020,N_13817,N_13962);
or U14021 (N_14021,N_13902,N_13809);
and U14022 (N_14022,N_13932,N_13797);
or U14023 (N_14023,N_13973,N_13975);
and U14024 (N_14024,N_13882,N_13917);
nand U14025 (N_14025,N_13967,N_13887);
and U14026 (N_14026,N_13878,N_13803);
nand U14027 (N_14027,N_13795,N_13822);
or U14028 (N_14028,N_13951,N_13963);
nor U14029 (N_14029,N_13812,N_13834);
nand U14030 (N_14030,N_13773,N_13936);
nand U14031 (N_14031,N_13816,N_13846);
nand U14032 (N_14032,N_13928,N_13992);
or U14033 (N_14033,N_13921,N_13768);
nor U14034 (N_14034,N_13793,N_13926);
nand U14035 (N_14035,N_13871,N_13999);
and U14036 (N_14036,N_13943,N_13988);
and U14037 (N_14037,N_13875,N_13784);
xnor U14038 (N_14038,N_13866,N_13781);
or U14039 (N_14039,N_13826,N_13788);
or U14040 (N_14040,N_13987,N_13813);
and U14041 (N_14041,N_13776,N_13908);
xnor U14042 (N_14042,N_13818,N_13995);
nor U14043 (N_14043,N_13918,N_13760);
nor U14044 (N_14044,N_13799,N_13832);
nor U14045 (N_14045,N_13955,N_13897);
nor U14046 (N_14046,N_13777,N_13839);
and U14047 (N_14047,N_13954,N_13880);
nor U14048 (N_14048,N_13886,N_13968);
nand U14049 (N_14049,N_13850,N_13906);
xnor U14050 (N_14050,N_13792,N_13804);
and U14051 (N_14051,N_13863,N_13920);
nand U14052 (N_14052,N_13775,N_13762);
xnor U14053 (N_14053,N_13758,N_13979);
and U14054 (N_14054,N_13772,N_13841);
or U14055 (N_14055,N_13916,N_13845);
nor U14056 (N_14056,N_13910,N_13991);
or U14057 (N_14057,N_13894,N_13885);
nor U14058 (N_14058,N_13970,N_13934);
or U14059 (N_14059,N_13900,N_13774);
or U14060 (N_14060,N_13892,N_13755);
nor U14061 (N_14061,N_13956,N_13761);
and U14062 (N_14062,N_13924,N_13778);
or U14063 (N_14063,N_13937,N_13794);
nor U14064 (N_14064,N_13965,N_13815);
nor U14065 (N_14065,N_13969,N_13814);
xnor U14066 (N_14066,N_13913,N_13801);
nand U14067 (N_14067,N_13874,N_13980);
xnor U14068 (N_14068,N_13825,N_13754);
or U14069 (N_14069,N_13848,N_13859);
or U14070 (N_14070,N_13949,N_13864);
or U14071 (N_14071,N_13786,N_13948);
or U14072 (N_14072,N_13843,N_13808);
nor U14073 (N_14073,N_13840,N_13753);
or U14074 (N_14074,N_13872,N_13877);
nand U14075 (N_14075,N_13898,N_13983);
or U14076 (N_14076,N_13782,N_13947);
nand U14077 (N_14077,N_13883,N_13785);
nand U14078 (N_14078,N_13798,N_13901);
and U14079 (N_14079,N_13757,N_13862);
or U14080 (N_14080,N_13805,N_13854);
nand U14081 (N_14081,N_13847,N_13837);
or U14082 (N_14082,N_13942,N_13971);
nor U14083 (N_14083,N_13919,N_13997);
nor U14084 (N_14084,N_13870,N_13858);
nand U14085 (N_14085,N_13831,N_13899);
nand U14086 (N_14086,N_13851,N_13769);
xnor U14087 (N_14087,N_13994,N_13835);
nand U14088 (N_14088,N_13791,N_13868);
nor U14089 (N_14089,N_13959,N_13890);
xnor U14090 (N_14090,N_13946,N_13907);
nor U14091 (N_14091,N_13770,N_13930);
xnor U14092 (N_14092,N_13961,N_13964);
xnor U14093 (N_14093,N_13836,N_13842);
nor U14094 (N_14094,N_13931,N_13861);
and U14095 (N_14095,N_13881,N_13779);
or U14096 (N_14096,N_13750,N_13823);
nor U14097 (N_14097,N_13869,N_13903);
and U14098 (N_14098,N_13853,N_13978);
and U14099 (N_14099,N_13998,N_13810);
nand U14100 (N_14100,N_13819,N_13914);
or U14101 (N_14101,N_13993,N_13783);
or U14102 (N_14102,N_13915,N_13867);
or U14103 (N_14103,N_13857,N_13849);
nor U14104 (N_14104,N_13751,N_13996);
nor U14105 (N_14105,N_13990,N_13838);
nand U14106 (N_14106,N_13929,N_13950);
and U14107 (N_14107,N_13765,N_13827);
or U14108 (N_14108,N_13865,N_13833);
xnor U14109 (N_14109,N_13953,N_13821);
nor U14110 (N_14110,N_13796,N_13766);
nand U14111 (N_14111,N_13764,N_13985);
xor U14112 (N_14112,N_13958,N_13957);
or U14113 (N_14113,N_13856,N_13891);
xnor U14114 (N_14114,N_13982,N_13986);
xor U14115 (N_14115,N_13888,N_13876);
xnor U14116 (N_14116,N_13852,N_13830);
nand U14117 (N_14117,N_13884,N_13807);
nor U14118 (N_14118,N_13904,N_13966);
or U14119 (N_14119,N_13972,N_13935);
nand U14120 (N_14120,N_13787,N_13939);
or U14121 (N_14121,N_13889,N_13940);
nand U14122 (N_14122,N_13933,N_13984);
or U14123 (N_14123,N_13828,N_13952);
xnor U14124 (N_14124,N_13759,N_13923);
xor U14125 (N_14125,N_13795,N_13940);
nor U14126 (N_14126,N_13935,N_13901);
and U14127 (N_14127,N_13957,N_13943);
nand U14128 (N_14128,N_13971,N_13992);
and U14129 (N_14129,N_13960,N_13880);
and U14130 (N_14130,N_13979,N_13806);
xor U14131 (N_14131,N_13875,N_13946);
and U14132 (N_14132,N_13962,N_13888);
xor U14133 (N_14133,N_13845,N_13861);
nor U14134 (N_14134,N_13888,N_13848);
xnor U14135 (N_14135,N_13804,N_13828);
xnor U14136 (N_14136,N_13972,N_13861);
or U14137 (N_14137,N_13811,N_13849);
and U14138 (N_14138,N_13882,N_13814);
and U14139 (N_14139,N_13768,N_13985);
xnor U14140 (N_14140,N_13984,N_13826);
or U14141 (N_14141,N_13771,N_13975);
xnor U14142 (N_14142,N_13882,N_13823);
nand U14143 (N_14143,N_13753,N_13886);
and U14144 (N_14144,N_13931,N_13955);
or U14145 (N_14145,N_13872,N_13861);
or U14146 (N_14146,N_13901,N_13985);
or U14147 (N_14147,N_13851,N_13810);
nand U14148 (N_14148,N_13818,N_13776);
nand U14149 (N_14149,N_13819,N_13894);
xnor U14150 (N_14150,N_13807,N_13811);
xor U14151 (N_14151,N_13760,N_13884);
or U14152 (N_14152,N_13844,N_13937);
nand U14153 (N_14153,N_13830,N_13847);
nand U14154 (N_14154,N_13898,N_13891);
nand U14155 (N_14155,N_13873,N_13799);
xor U14156 (N_14156,N_13832,N_13850);
and U14157 (N_14157,N_13937,N_13866);
nor U14158 (N_14158,N_13905,N_13835);
or U14159 (N_14159,N_13958,N_13753);
and U14160 (N_14160,N_13768,N_13809);
nor U14161 (N_14161,N_13763,N_13986);
nand U14162 (N_14162,N_13986,N_13780);
xnor U14163 (N_14163,N_13794,N_13849);
xnor U14164 (N_14164,N_13905,N_13992);
xnor U14165 (N_14165,N_13988,N_13764);
nand U14166 (N_14166,N_13757,N_13849);
nand U14167 (N_14167,N_13920,N_13761);
nor U14168 (N_14168,N_13809,N_13907);
nor U14169 (N_14169,N_13758,N_13985);
nor U14170 (N_14170,N_13893,N_13950);
xnor U14171 (N_14171,N_13813,N_13949);
nand U14172 (N_14172,N_13788,N_13867);
nor U14173 (N_14173,N_13948,N_13996);
xnor U14174 (N_14174,N_13777,N_13834);
nor U14175 (N_14175,N_13955,N_13964);
and U14176 (N_14176,N_13940,N_13982);
nor U14177 (N_14177,N_13906,N_13947);
xnor U14178 (N_14178,N_13765,N_13897);
and U14179 (N_14179,N_13980,N_13971);
nand U14180 (N_14180,N_13955,N_13944);
nor U14181 (N_14181,N_13779,N_13892);
xor U14182 (N_14182,N_13931,N_13893);
xnor U14183 (N_14183,N_13998,N_13981);
or U14184 (N_14184,N_13812,N_13775);
and U14185 (N_14185,N_13852,N_13838);
or U14186 (N_14186,N_13982,N_13888);
or U14187 (N_14187,N_13801,N_13989);
and U14188 (N_14188,N_13752,N_13794);
nand U14189 (N_14189,N_13838,N_13817);
and U14190 (N_14190,N_13986,N_13879);
nor U14191 (N_14191,N_13909,N_13833);
and U14192 (N_14192,N_13891,N_13958);
xnor U14193 (N_14193,N_13773,N_13809);
nand U14194 (N_14194,N_13819,N_13992);
or U14195 (N_14195,N_13813,N_13995);
nand U14196 (N_14196,N_13755,N_13829);
and U14197 (N_14197,N_13815,N_13787);
and U14198 (N_14198,N_13991,N_13920);
and U14199 (N_14199,N_13843,N_13941);
nand U14200 (N_14200,N_13940,N_13831);
or U14201 (N_14201,N_13763,N_13794);
nand U14202 (N_14202,N_13896,N_13990);
and U14203 (N_14203,N_13843,N_13801);
and U14204 (N_14204,N_13778,N_13791);
nand U14205 (N_14205,N_13990,N_13824);
xnor U14206 (N_14206,N_13879,N_13832);
and U14207 (N_14207,N_13827,N_13770);
or U14208 (N_14208,N_13766,N_13975);
and U14209 (N_14209,N_13969,N_13900);
and U14210 (N_14210,N_13767,N_13832);
xnor U14211 (N_14211,N_13856,N_13926);
nor U14212 (N_14212,N_13972,N_13919);
or U14213 (N_14213,N_13946,N_13993);
nor U14214 (N_14214,N_13891,N_13850);
nand U14215 (N_14215,N_13847,N_13783);
xnor U14216 (N_14216,N_13780,N_13904);
or U14217 (N_14217,N_13931,N_13909);
nand U14218 (N_14218,N_13966,N_13789);
and U14219 (N_14219,N_13895,N_13871);
nor U14220 (N_14220,N_13770,N_13796);
and U14221 (N_14221,N_13932,N_13793);
and U14222 (N_14222,N_13796,N_13788);
and U14223 (N_14223,N_13956,N_13910);
or U14224 (N_14224,N_13851,N_13980);
nand U14225 (N_14225,N_13980,N_13771);
nand U14226 (N_14226,N_13997,N_13902);
or U14227 (N_14227,N_13893,N_13801);
xor U14228 (N_14228,N_13772,N_13890);
and U14229 (N_14229,N_13880,N_13987);
nor U14230 (N_14230,N_13763,N_13862);
and U14231 (N_14231,N_13845,N_13975);
nor U14232 (N_14232,N_13927,N_13872);
nor U14233 (N_14233,N_13987,N_13786);
and U14234 (N_14234,N_13750,N_13999);
nand U14235 (N_14235,N_13967,N_13778);
nor U14236 (N_14236,N_13770,N_13754);
and U14237 (N_14237,N_13830,N_13893);
nand U14238 (N_14238,N_13841,N_13930);
and U14239 (N_14239,N_13962,N_13804);
xnor U14240 (N_14240,N_13856,N_13905);
xor U14241 (N_14241,N_13837,N_13899);
nand U14242 (N_14242,N_13872,N_13804);
or U14243 (N_14243,N_13781,N_13799);
nor U14244 (N_14244,N_13935,N_13896);
and U14245 (N_14245,N_13793,N_13859);
nor U14246 (N_14246,N_13932,N_13787);
nand U14247 (N_14247,N_13938,N_13934);
nor U14248 (N_14248,N_13794,N_13952);
or U14249 (N_14249,N_13853,N_13871);
nand U14250 (N_14250,N_14180,N_14160);
or U14251 (N_14251,N_14146,N_14000);
nor U14252 (N_14252,N_14200,N_14070);
and U14253 (N_14253,N_14042,N_14228);
nor U14254 (N_14254,N_14044,N_14106);
nand U14255 (N_14255,N_14125,N_14004);
or U14256 (N_14256,N_14154,N_14054);
and U14257 (N_14257,N_14166,N_14179);
nor U14258 (N_14258,N_14178,N_14235);
xor U14259 (N_14259,N_14056,N_14082);
xor U14260 (N_14260,N_14151,N_14142);
and U14261 (N_14261,N_14080,N_14077);
and U14262 (N_14262,N_14079,N_14173);
or U14263 (N_14263,N_14061,N_14199);
and U14264 (N_14264,N_14144,N_14021);
nand U14265 (N_14265,N_14171,N_14234);
xor U14266 (N_14266,N_14205,N_14022);
and U14267 (N_14267,N_14206,N_14233);
xnor U14268 (N_14268,N_14148,N_14087);
or U14269 (N_14269,N_14204,N_14109);
nand U14270 (N_14270,N_14031,N_14203);
xnor U14271 (N_14271,N_14157,N_14005);
and U14272 (N_14272,N_14229,N_14218);
nor U14273 (N_14273,N_14115,N_14176);
nor U14274 (N_14274,N_14183,N_14138);
nor U14275 (N_14275,N_14248,N_14210);
xnor U14276 (N_14276,N_14094,N_14065);
nand U14277 (N_14277,N_14222,N_14242);
and U14278 (N_14278,N_14245,N_14165);
and U14279 (N_14279,N_14055,N_14040);
or U14280 (N_14280,N_14129,N_14091);
and U14281 (N_14281,N_14013,N_14053);
and U14282 (N_14282,N_14103,N_14038);
and U14283 (N_14283,N_14137,N_14052);
and U14284 (N_14284,N_14249,N_14023);
xnor U14285 (N_14285,N_14043,N_14036);
nand U14286 (N_14286,N_14059,N_14118);
nor U14287 (N_14287,N_14012,N_14241);
or U14288 (N_14288,N_14107,N_14064);
and U14289 (N_14289,N_14236,N_14134);
nand U14290 (N_14290,N_14223,N_14132);
and U14291 (N_14291,N_14007,N_14239);
and U14292 (N_14292,N_14133,N_14037);
nand U14293 (N_14293,N_14159,N_14126);
or U14294 (N_14294,N_14127,N_14030);
nor U14295 (N_14295,N_14175,N_14009);
xnor U14296 (N_14296,N_14045,N_14076);
and U14297 (N_14297,N_14006,N_14122);
nor U14298 (N_14298,N_14098,N_14163);
nor U14299 (N_14299,N_14237,N_14170);
nand U14300 (N_14300,N_14135,N_14075);
or U14301 (N_14301,N_14083,N_14025);
nand U14302 (N_14302,N_14208,N_14145);
or U14303 (N_14303,N_14120,N_14008);
nor U14304 (N_14304,N_14111,N_14214);
xnor U14305 (N_14305,N_14188,N_14110);
or U14306 (N_14306,N_14035,N_14168);
nand U14307 (N_14307,N_14131,N_14243);
or U14308 (N_14308,N_14071,N_14177);
and U14309 (N_14309,N_14136,N_14156);
or U14310 (N_14310,N_14017,N_14153);
nand U14311 (N_14311,N_14217,N_14169);
and U14312 (N_14312,N_14193,N_14139);
or U14313 (N_14313,N_14211,N_14224);
or U14314 (N_14314,N_14181,N_14162);
xnor U14315 (N_14315,N_14024,N_14086);
or U14316 (N_14316,N_14072,N_14119);
and U14317 (N_14317,N_14128,N_14066);
and U14318 (N_14318,N_14041,N_14124);
or U14319 (N_14319,N_14027,N_14196);
nand U14320 (N_14320,N_14194,N_14058);
xnor U14321 (N_14321,N_14112,N_14020);
or U14322 (N_14322,N_14231,N_14149);
xnor U14323 (N_14323,N_14186,N_14213);
or U14324 (N_14324,N_14247,N_14028);
nand U14325 (N_14325,N_14141,N_14039);
nand U14326 (N_14326,N_14114,N_14067);
nor U14327 (N_14327,N_14001,N_14051);
xnor U14328 (N_14328,N_14097,N_14232);
and U14329 (N_14329,N_14150,N_14197);
or U14330 (N_14330,N_14209,N_14099);
nand U14331 (N_14331,N_14090,N_14155);
or U14332 (N_14332,N_14113,N_14121);
and U14333 (N_14333,N_14172,N_14018);
and U14334 (N_14334,N_14011,N_14057);
xnor U14335 (N_14335,N_14225,N_14182);
nor U14336 (N_14336,N_14060,N_14100);
and U14337 (N_14337,N_14221,N_14085);
or U14338 (N_14338,N_14081,N_14084);
nor U14339 (N_14339,N_14198,N_14152);
nand U14340 (N_14340,N_14220,N_14201);
nor U14341 (N_14341,N_14140,N_14202);
and U14342 (N_14342,N_14029,N_14095);
or U14343 (N_14343,N_14050,N_14123);
and U14344 (N_14344,N_14074,N_14164);
xor U14345 (N_14345,N_14046,N_14010);
nand U14346 (N_14346,N_14089,N_14212);
nand U14347 (N_14347,N_14185,N_14026);
or U14348 (N_14348,N_14238,N_14063);
or U14349 (N_14349,N_14184,N_14096);
xor U14350 (N_14350,N_14230,N_14019);
nand U14351 (N_14351,N_14105,N_14032);
nand U14352 (N_14352,N_14195,N_14062);
or U14353 (N_14353,N_14190,N_14092);
and U14354 (N_14354,N_14219,N_14246);
and U14355 (N_14355,N_14014,N_14240);
nor U14356 (N_14356,N_14158,N_14130);
xor U14357 (N_14357,N_14207,N_14161);
xor U14358 (N_14358,N_14069,N_14226);
xnor U14359 (N_14359,N_14108,N_14049);
and U14360 (N_14360,N_14174,N_14102);
and U14361 (N_14361,N_14167,N_14078);
nor U14362 (N_14362,N_14048,N_14101);
and U14363 (N_14363,N_14216,N_14068);
xor U14364 (N_14364,N_14034,N_14143);
or U14365 (N_14365,N_14215,N_14016);
nor U14366 (N_14366,N_14033,N_14047);
and U14367 (N_14367,N_14192,N_14104);
xor U14368 (N_14368,N_14189,N_14191);
nand U14369 (N_14369,N_14147,N_14002);
nor U14370 (N_14370,N_14227,N_14244);
and U14371 (N_14371,N_14015,N_14116);
or U14372 (N_14372,N_14003,N_14073);
or U14373 (N_14373,N_14117,N_14187);
nand U14374 (N_14374,N_14088,N_14093);
xor U14375 (N_14375,N_14133,N_14094);
nand U14376 (N_14376,N_14165,N_14184);
nor U14377 (N_14377,N_14187,N_14007);
or U14378 (N_14378,N_14016,N_14166);
nor U14379 (N_14379,N_14102,N_14197);
and U14380 (N_14380,N_14101,N_14123);
nand U14381 (N_14381,N_14176,N_14168);
and U14382 (N_14382,N_14201,N_14211);
nor U14383 (N_14383,N_14042,N_14183);
or U14384 (N_14384,N_14071,N_14057);
nor U14385 (N_14385,N_14141,N_14197);
and U14386 (N_14386,N_14092,N_14148);
nand U14387 (N_14387,N_14213,N_14130);
nor U14388 (N_14388,N_14056,N_14055);
nor U14389 (N_14389,N_14232,N_14095);
and U14390 (N_14390,N_14006,N_14037);
xor U14391 (N_14391,N_14075,N_14061);
or U14392 (N_14392,N_14019,N_14169);
xor U14393 (N_14393,N_14224,N_14243);
nor U14394 (N_14394,N_14093,N_14004);
xor U14395 (N_14395,N_14004,N_14034);
xnor U14396 (N_14396,N_14176,N_14175);
xnor U14397 (N_14397,N_14079,N_14077);
or U14398 (N_14398,N_14203,N_14139);
or U14399 (N_14399,N_14127,N_14242);
nor U14400 (N_14400,N_14057,N_14083);
xor U14401 (N_14401,N_14014,N_14224);
xnor U14402 (N_14402,N_14207,N_14132);
xor U14403 (N_14403,N_14089,N_14084);
nor U14404 (N_14404,N_14001,N_14054);
xnor U14405 (N_14405,N_14188,N_14128);
or U14406 (N_14406,N_14166,N_14216);
and U14407 (N_14407,N_14184,N_14000);
or U14408 (N_14408,N_14235,N_14029);
and U14409 (N_14409,N_14006,N_14238);
nand U14410 (N_14410,N_14237,N_14193);
xnor U14411 (N_14411,N_14113,N_14140);
and U14412 (N_14412,N_14173,N_14130);
and U14413 (N_14413,N_14213,N_14193);
nor U14414 (N_14414,N_14004,N_14032);
or U14415 (N_14415,N_14224,N_14065);
nor U14416 (N_14416,N_14227,N_14121);
or U14417 (N_14417,N_14084,N_14204);
or U14418 (N_14418,N_14012,N_14148);
xor U14419 (N_14419,N_14047,N_14102);
and U14420 (N_14420,N_14234,N_14046);
nand U14421 (N_14421,N_14060,N_14175);
or U14422 (N_14422,N_14205,N_14061);
or U14423 (N_14423,N_14070,N_14164);
nand U14424 (N_14424,N_14200,N_14129);
nand U14425 (N_14425,N_14234,N_14039);
and U14426 (N_14426,N_14037,N_14120);
or U14427 (N_14427,N_14017,N_14150);
and U14428 (N_14428,N_14197,N_14063);
nor U14429 (N_14429,N_14131,N_14107);
xnor U14430 (N_14430,N_14131,N_14022);
and U14431 (N_14431,N_14055,N_14052);
xor U14432 (N_14432,N_14007,N_14097);
and U14433 (N_14433,N_14153,N_14159);
nand U14434 (N_14434,N_14076,N_14180);
and U14435 (N_14435,N_14120,N_14101);
or U14436 (N_14436,N_14030,N_14034);
xor U14437 (N_14437,N_14170,N_14112);
xnor U14438 (N_14438,N_14112,N_14078);
or U14439 (N_14439,N_14072,N_14040);
nor U14440 (N_14440,N_14215,N_14245);
or U14441 (N_14441,N_14001,N_14188);
nor U14442 (N_14442,N_14131,N_14144);
xor U14443 (N_14443,N_14085,N_14058);
nand U14444 (N_14444,N_14054,N_14182);
nor U14445 (N_14445,N_14016,N_14152);
nor U14446 (N_14446,N_14127,N_14090);
nand U14447 (N_14447,N_14177,N_14046);
nor U14448 (N_14448,N_14105,N_14247);
and U14449 (N_14449,N_14198,N_14221);
nor U14450 (N_14450,N_14008,N_14216);
or U14451 (N_14451,N_14179,N_14201);
or U14452 (N_14452,N_14162,N_14079);
xor U14453 (N_14453,N_14035,N_14067);
nor U14454 (N_14454,N_14116,N_14076);
nand U14455 (N_14455,N_14030,N_14141);
xor U14456 (N_14456,N_14030,N_14036);
nand U14457 (N_14457,N_14198,N_14174);
nor U14458 (N_14458,N_14065,N_14138);
nor U14459 (N_14459,N_14109,N_14143);
xnor U14460 (N_14460,N_14118,N_14107);
nand U14461 (N_14461,N_14019,N_14203);
nand U14462 (N_14462,N_14053,N_14193);
or U14463 (N_14463,N_14088,N_14013);
and U14464 (N_14464,N_14008,N_14058);
and U14465 (N_14465,N_14094,N_14046);
nand U14466 (N_14466,N_14235,N_14152);
nor U14467 (N_14467,N_14190,N_14056);
nand U14468 (N_14468,N_14034,N_14216);
nor U14469 (N_14469,N_14223,N_14238);
xnor U14470 (N_14470,N_14161,N_14123);
nand U14471 (N_14471,N_14056,N_14167);
or U14472 (N_14472,N_14069,N_14122);
nor U14473 (N_14473,N_14226,N_14126);
and U14474 (N_14474,N_14245,N_14074);
nor U14475 (N_14475,N_14101,N_14172);
nor U14476 (N_14476,N_14109,N_14181);
or U14477 (N_14477,N_14065,N_14023);
xor U14478 (N_14478,N_14148,N_14071);
nand U14479 (N_14479,N_14190,N_14047);
and U14480 (N_14480,N_14013,N_14228);
xnor U14481 (N_14481,N_14240,N_14085);
or U14482 (N_14482,N_14002,N_14222);
or U14483 (N_14483,N_14061,N_14110);
and U14484 (N_14484,N_14197,N_14165);
xor U14485 (N_14485,N_14028,N_14127);
nor U14486 (N_14486,N_14086,N_14195);
nand U14487 (N_14487,N_14111,N_14196);
nand U14488 (N_14488,N_14246,N_14087);
or U14489 (N_14489,N_14214,N_14091);
xor U14490 (N_14490,N_14035,N_14247);
xor U14491 (N_14491,N_14084,N_14119);
and U14492 (N_14492,N_14018,N_14032);
or U14493 (N_14493,N_14139,N_14076);
xor U14494 (N_14494,N_14136,N_14043);
nor U14495 (N_14495,N_14239,N_14176);
nor U14496 (N_14496,N_14150,N_14133);
or U14497 (N_14497,N_14168,N_14064);
nor U14498 (N_14498,N_14148,N_14023);
or U14499 (N_14499,N_14191,N_14053);
xor U14500 (N_14500,N_14318,N_14349);
and U14501 (N_14501,N_14292,N_14269);
nor U14502 (N_14502,N_14443,N_14267);
or U14503 (N_14503,N_14343,N_14458);
and U14504 (N_14504,N_14304,N_14351);
or U14505 (N_14505,N_14475,N_14363);
or U14506 (N_14506,N_14287,N_14310);
nand U14507 (N_14507,N_14253,N_14412);
and U14508 (N_14508,N_14383,N_14470);
nand U14509 (N_14509,N_14450,N_14407);
and U14510 (N_14510,N_14305,N_14442);
nand U14511 (N_14511,N_14497,N_14333);
or U14512 (N_14512,N_14395,N_14411);
and U14513 (N_14513,N_14452,N_14466);
xnor U14514 (N_14514,N_14430,N_14386);
nor U14515 (N_14515,N_14300,N_14439);
or U14516 (N_14516,N_14321,N_14274);
and U14517 (N_14517,N_14423,N_14424);
and U14518 (N_14518,N_14449,N_14332);
nor U14519 (N_14519,N_14499,N_14284);
nor U14520 (N_14520,N_14266,N_14422);
or U14521 (N_14521,N_14486,N_14460);
nor U14522 (N_14522,N_14484,N_14462);
and U14523 (N_14523,N_14282,N_14357);
nor U14524 (N_14524,N_14371,N_14342);
xor U14525 (N_14525,N_14431,N_14285);
xnor U14526 (N_14526,N_14329,N_14348);
nor U14527 (N_14527,N_14467,N_14252);
xnor U14528 (N_14528,N_14391,N_14438);
nor U14529 (N_14529,N_14382,N_14402);
xor U14530 (N_14530,N_14447,N_14365);
or U14531 (N_14531,N_14487,N_14378);
xor U14532 (N_14532,N_14280,N_14355);
or U14533 (N_14533,N_14405,N_14306);
and U14534 (N_14534,N_14369,N_14436);
nor U14535 (N_14535,N_14297,N_14367);
and U14536 (N_14536,N_14415,N_14250);
nor U14537 (N_14537,N_14472,N_14441);
or U14538 (N_14538,N_14334,N_14373);
xor U14539 (N_14539,N_14468,N_14320);
xor U14540 (N_14540,N_14396,N_14356);
or U14541 (N_14541,N_14265,N_14327);
nand U14542 (N_14542,N_14455,N_14276);
nor U14543 (N_14543,N_14473,N_14414);
and U14544 (N_14544,N_14485,N_14437);
and U14545 (N_14545,N_14398,N_14317);
or U14546 (N_14546,N_14393,N_14429);
xor U14547 (N_14547,N_14254,N_14289);
nor U14548 (N_14548,N_14370,N_14403);
xor U14549 (N_14549,N_14469,N_14338);
nand U14550 (N_14550,N_14433,N_14278);
or U14551 (N_14551,N_14359,N_14491);
xnor U14552 (N_14552,N_14260,N_14453);
xnor U14553 (N_14553,N_14425,N_14339);
xnor U14554 (N_14554,N_14457,N_14299);
and U14555 (N_14555,N_14296,N_14496);
xnor U14556 (N_14556,N_14319,N_14498);
and U14557 (N_14557,N_14413,N_14379);
nand U14558 (N_14558,N_14459,N_14283);
and U14559 (N_14559,N_14340,N_14481);
or U14560 (N_14560,N_14346,N_14328);
and U14561 (N_14561,N_14324,N_14388);
nor U14562 (N_14562,N_14432,N_14419);
nor U14563 (N_14563,N_14286,N_14418);
or U14564 (N_14564,N_14352,N_14477);
or U14565 (N_14565,N_14387,N_14307);
xor U14566 (N_14566,N_14313,N_14353);
xnor U14567 (N_14567,N_14344,N_14277);
or U14568 (N_14568,N_14440,N_14301);
or U14569 (N_14569,N_14456,N_14392);
or U14570 (N_14570,N_14331,N_14483);
nand U14571 (N_14571,N_14416,N_14397);
nand U14572 (N_14572,N_14314,N_14273);
and U14573 (N_14573,N_14354,N_14270);
nor U14574 (N_14574,N_14368,N_14345);
nor U14575 (N_14575,N_14364,N_14259);
and U14576 (N_14576,N_14302,N_14362);
nor U14577 (N_14577,N_14281,N_14406);
xnor U14578 (N_14578,N_14279,N_14464);
nor U14579 (N_14579,N_14463,N_14474);
nor U14580 (N_14580,N_14444,N_14336);
xnor U14581 (N_14581,N_14490,N_14295);
and U14582 (N_14582,N_14465,N_14401);
nand U14583 (N_14583,N_14476,N_14261);
xnor U14584 (N_14584,N_14291,N_14316);
nor U14585 (N_14585,N_14272,N_14445);
or U14586 (N_14586,N_14294,N_14394);
nand U14587 (N_14587,N_14375,N_14380);
nor U14588 (N_14588,N_14381,N_14374);
or U14589 (N_14589,N_14309,N_14385);
nand U14590 (N_14590,N_14493,N_14315);
nand U14591 (N_14591,N_14390,N_14410);
or U14592 (N_14592,N_14420,N_14489);
nor U14593 (N_14593,N_14461,N_14341);
nand U14594 (N_14594,N_14372,N_14262);
nand U14595 (N_14595,N_14492,N_14389);
xor U14596 (N_14596,N_14330,N_14298);
nand U14597 (N_14597,N_14399,N_14479);
nor U14598 (N_14598,N_14408,N_14358);
nand U14599 (N_14599,N_14421,N_14290);
or U14600 (N_14600,N_14360,N_14495);
or U14601 (N_14601,N_14256,N_14384);
or U14602 (N_14602,N_14488,N_14293);
and U14603 (N_14603,N_14251,N_14303);
nor U14604 (N_14604,N_14264,N_14366);
and U14605 (N_14605,N_14400,N_14478);
or U14606 (N_14606,N_14494,N_14326);
xnor U14607 (N_14607,N_14435,N_14335);
nor U14608 (N_14608,N_14312,N_14482);
nor U14609 (N_14609,N_14323,N_14451);
xor U14610 (N_14610,N_14325,N_14361);
xor U14611 (N_14611,N_14434,N_14288);
nor U14612 (N_14612,N_14322,N_14404);
xnor U14613 (N_14613,N_14257,N_14448);
nand U14614 (N_14614,N_14480,N_14337);
or U14615 (N_14615,N_14376,N_14255);
or U14616 (N_14616,N_14409,N_14311);
nand U14617 (N_14617,N_14308,N_14263);
xnor U14618 (N_14618,N_14454,N_14377);
or U14619 (N_14619,N_14347,N_14258);
nor U14620 (N_14620,N_14268,N_14426);
or U14621 (N_14621,N_14471,N_14271);
xor U14622 (N_14622,N_14428,N_14350);
xnor U14623 (N_14623,N_14275,N_14427);
nand U14624 (N_14624,N_14446,N_14417);
or U14625 (N_14625,N_14348,N_14499);
nor U14626 (N_14626,N_14301,N_14445);
nor U14627 (N_14627,N_14371,N_14496);
or U14628 (N_14628,N_14350,N_14479);
xor U14629 (N_14629,N_14380,N_14454);
and U14630 (N_14630,N_14371,N_14392);
xor U14631 (N_14631,N_14374,N_14498);
and U14632 (N_14632,N_14488,N_14315);
nand U14633 (N_14633,N_14377,N_14305);
xnor U14634 (N_14634,N_14292,N_14373);
or U14635 (N_14635,N_14420,N_14451);
and U14636 (N_14636,N_14311,N_14470);
nand U14637 (N_14637,N_14329,N_14376);
or U14638 (N_14638,N_14277,N_14408);
or U14639 (N_14639,N_14446,N_14293);
and U14640 (N_14640,N_14361,N_14405);
or U14641 (N_14641,N_14455,N_14376);
or U14642 (N_14642,N_14324,N_14316);
or U14643 (N_14643,N_14276,N_14482);
nor U14644 (N_14644,N_14285,N_14381);
nand U14645 (N_14645,N_14465,N_14359);
xnor U14646 (N_14646,N_14359,N_14407);
nor U14647 (N_14647,N_14251,N_14337);
and U14648 (N_14648,N_14381,N_14289);
or U14649 (N_14649,N_14277,N_14486);
nand U14650 (N_14650,N_14447,N_14366);
xor U14651 (N_14651,N_14316,N_14370);
xor U14652 (N_14652,N_14302,N_14329);
nor U14653 (N_14653,N_14357,N_14317);
xnor U14654 (N_14654,N_14496,N_14449);
nor U14655 (N_14655,N_14472,N_14289);
xnor U14656 (N_14656,N_14364,N_14360);
nand U14657 (N_14657,N_14437,N_14405);
xor U14658 (N_14658,N_14314,N_14258);
xor U14659 (N_14659,N_14302,N_14383);
and U14660 (N_14660,N_14268,N_14467);
or U14661 (N_14661,N_14307,N_14385);
nand U14662 (N_14662,N_14448,N_14480);
xor U14663 (N_14663,N_14415,N_14331);
nor U14664 (N_14664,N_14295,N_14419);
or U14665 (N_14665,N_14250,N_14468);
or U14666 (N_14666,N_14262,N_14369);
and U14667 (N_14667,N_14493,N_14354);
nor U14668 (N_14668,N_14472,N_14366);
nor U14669 (N_14669,N_14277,N_14474);
xor U14670 (N_14670,N_14420,N_14347);
nor U14671 (N_14671,N_14443,N_14398);
or U14672 (N_14672,N_14490,N_14396);
or U14673 (N_14673,N_14497,N_14347);
or U14674 (N_14674,N_14267,N_14286);
xor U14675 (N_14675,N_14267,N_14357);
nand U14676 (N_14676,N_14253,N_14292);
nand U14677 (N_14677,N_14324,N_14406);
nor U14678 (N_14678,N_14407,N_14334);
xor U14679 (N_14679,N_14392,N_14272);
or U14680 (N_14680,N_14338,N_14403);
nor U14681 (N_14681,N_14449,N_14295);
nor U14682 (N_14682,N_14481,N_14313);
xor U14683 (N_14683,N_14462,N_14434);
xnor U14684 (N_14684,N_14260,N_14294);
nand U14685 (N_14685,N_14470,N_14345);
and U14686 (N_14686,N_14251,N_14467);
xnor U14687 (N_14687,N_14397,N_14417);
xor U14688 (N_14688,N_14402,N_14336);
nor U14689 (N_14689,N_14349,N_14343);
nand U14690 (N_14690,N_14352,N_14414);
xnor U14691 (N_14691,N_14314,N_14297);
and U14692 (N_14692,N_14442,N_14253);
nand U14693 (N_14693,N_14282,N_14469);
xor U14694 (N_14694,N_14338,N_14320);
nor U14695 (N_14695,N_14344,N_14484);
nand U14696 (N_14696,N_14254,N_14361);
nand U14697 (N_14697,N_14494,N_14357);
nor U14698 (N_14698,N_14407,N_14321);
nand U14699 (N_14699,N_14382,N_14278);
or U14700 (N_14700,N_14416,N_14337);
and U14701 (N_14701,N_14257,N_14292);
xnor U14702 (N_14702,N_14471,N_14354);
xnor U14703 (N_14703,N_14472,N_14298);
xor U14704 (N_14704,N_14448,N_14491);
and U14705 (N_14705,N_14446,N_14257);
nand U14706 (N_14706,N_14318,N_14270);
xor U14707 (N_14707,N_14419,N_14397);
nand U14708 (N_14708,N_14443,N_14379);
xnor U14709 (N_14709,N_14393,N_14307);
nor U14710 (N_14710,N_14440,N_14441);
nor U14711 (N_14711,N_14458,N_14489);
or U14712 (N_14712,N_14308,N_14353);
xor U14713 (N_14713,N_14380,N_14470);
or U14714 (N_14714,N_14323,N_14317);
and U14715 (N_14715,N_14299,N_14377);
nand U14716 (N_14716,N_14424,N_14335);
and U14717 (N_14717,N_14441,N_14396);
nor U14718 (N_14718,N_14356,N_14323);
nand U14719 (N_14719,N_14355,N_14473);
xor U14720 (N_14720,N_14472,N_14254);
or U14721 (N_14721,N_14358,N_14348);
nor U14722 (N_14722,N_14432,N_14393);
nand U14723 (N_14723,N_14324,N_14367);
nor U14724 (N_14724,N_14451,N_14330);
nor U14725 (N_14725,N_14304,N_14382);
or U14726 (N_14726,N_14324,N_14402);
and U14727 (N_14727,N_14450,N_14303);
or U14728 (N_14728,N_14393,N_14349);
or U14729 (N_14729,N_14318,N_14354);
and U14730 (N_14730,N_14266,N_14494);
nand U14731 (N_14731,N_14384,N_14372);
xor U14732 (N_14732,N_14391,N_14490);
and U14733 (N_14733,N_14444,N_14279);
xor U14734 (N_14734,N_14270,N_14284);
xnor U14735 (N_14735,N_14343,N_14285);
nand U14736 (N_14736,N_14284,N_14420);
or U14737 (N_14737,N_14330,N_14393);
xnor U14738 (N_14738,N_14286,N_14253);
nand U14739 (N_14739,N_14496,N_14252);
or U14740 (N_14740,N_14257,N_14390);
xor U14741 (N_14741,N_14295,N_14280);
xor U14742 (N_14742,N_14290,N_14327);
nand U14743 (N_14743,N_14266,N_14416);
and U14744 (N_14744,N_14440,N_14377);
xor U14745 (N_14745,N_14436,N_14286);
nor U14746 (N_14746,N_14323,N_14310);
nor U14747 (N_14747,N_14283,N_14453);
or U14748 (N_14748,N_14333,N_14285);
nor U14749 (N_14749,N_14269,N_14489);
and U14750 (N_14750,N_14600,N_14581);
xnor U14751 (N_14751,N_14559,N_14685);
nand U14752 (N_14752,N_14553,N_14531);
and U14753 (N_14753,N_14594,N_14703);
or U14754 (N_14754,N_14572,N_14539);
or U14755 (N_14755,N_14623,N_14686);
nand U14756 (N_14756,N_14702,N_14588);
nor U14757 (N_14757,N_14620,N_14665);
nor U14758 (N_14758,N_14684,N_14676);
and U14759 (N_14759,N_14536,N_14723);
xor U14760 (N_14760,N_14564,N_14711);
or U14761 (N_14761,N_14601,N_14677);
and U14762 (N_14762,N_14640,N_14511);
xor U14763 (N_14763,N_14657,N_14687);
xnor U14764 (N_14764,N_14662,N_14726);
and U14765 (N_14765,N_14548,N_14655);
and U14766 (N_14766,N_14718,N_14603);
and U14767 (N_14767,N_14506,N_14610);
nand U14768 (N_14768,N_14527,N_14614);
nor U14769 (N_14769,N_14647,N_14627);
xnor U14770 (N_14770,N_14502,N_14645);
nor U14771 (N_14771,N_14574,N_14575);
or U14772 (N_14772,N_14613,N_14618);
nor U14773 (N_14773,N_14692,N_14570);
nand U14774 (N_14774,N_14745,N_14747);
or U14775 (N_14775,N_14681,N_14638);
and U14776 (N_14776,N_14517,N_14605);
nor U14777 (N_14777,N_14727,N_14631);
nor U14778 (N_14778,N_14519,N_14667);
nand U14779 (N_14779,N_14562,N_14652);
or U14780 (N_14780,N_14737,N_14615);
nand U14781 (N_14781,N_14543,N_14604);
nor U14782 (N_14782,N_14725,N_14617);
nand U14783 (N_14783,N_14733,N_14742);
xnor U14784 (N_14784,N_14584,N_14529);
nor U14785 (N_14785,N_14608,N_14596);
xnor U14786 (N_14786,N_14593,N_14508);
nor U14787 (N_14787,N_14509,N_14510);
xnor U14788 (N_14788,N_14670,N_14656);
nor U14789 (N_14789,N_14746,N_14609);
or U14790 (N_14790,N_14518,N_14621);
xnor U14791 (N_14791,N_14560,N_14546);
nor U14792 (N_14792,N_14644,N_14636);
nand U14793 (N_14793,N_14639,N_14635);
nor U14794 (N_14794,N_14749,N_14512);
xor U14795 (N_14795,N_14563,N_14671);
nor U14796 (N_14796,N_14629,N_14663);
and U14797 (N_14797,N_14558,N_14690);
nor U14798 (N_14798,N_14513,N_14688);
or U14799 (N_14799,N_14740,N_14541);
nor U14800 (N_14800,N_14535,N_14587);
or U14801 (N_14801,N_14622,N_14521);
nor U14802 (N_14802,N_14514,N_14646);
nand U14803 (N_14803,N_14731,N_14582);
xnor U14804 (N_14804,N_14526,N_14500);
and U14805 (N_14805,N_14547,N_14722);
and U14806 (N_14806,N_14710,N_14624);
xnor U14807 (N_14807,N_14602,N_14651);
and U14808 (N_14808,N_14701,N_14612);
or U14809 (N_14809,N_14683,N_14619);
and U14810 (N_14810,N_14532,N_14599);
or U14811 (N_14811,N_14672,N_14538);
and U14812 (N_14812,N_14598,N_14706);
nand U14813 (N_14813,N_14704,N_14632);
or U14814 (N_14814,N_14607,N_14578);
xor U14815 (N_14815,N_14567,N_14709);
and U14816 (N_14816,N_14586,N_14669);
nor U14817 (N_14817,N_14707,N_14503);
nor U14818 (N_14818,N_14679,N_14554);
and U14819 (N_14819,N_14659,N_14730);
and U14820 (N_14820,N_14520,N_14507);
and U14821 (N_14821,N_14550,N_14664);
xnor U14822 (N_14822,N_14736,N_14633);
nor U14823 (N_14823,N_14658,N_14625);
nor U14824 (N_14824,N_14649,N_14641);
nand U14825 (N_14825,N_14743,N_14589);
nor U14826 (N_14826,N_14678,N_14643);
nand U14827 (N_14827,N_14515,N_14720);
nor U14828 (N_14828,N_14525,N_14648);
xnor U14829 (N_14829,N_14561,N_14675);
nor U14830 (N_14830,N_14573,N_14650);
or U14831 (N_14831,N_14666,N_14501);
nor U14832 (N_14832,N_14583,N_14642);
xnor U14833 (N_14833,N_14698,N_14580);
or U14834 (N_14834,N_14748,N_14689);
xnor U14835 (N_14835,N_14597,N_14524);
and U14836 (N_14836,N_14533,N_14634);
or U14837 (N_14837,N_14660,N_14569);
and U14838 (N_14838,N_14566,N_14628);
or U14839 (N_14839,N_14697,N_14626);
xor U14840 (N_14840,N_14542,N_14571);
or U14841 (N_14841,N_14668,N_14616);
and U14842 (N_14842,N_14630,N_14595);
nand U14843 (N_14843,N_14549,N_14590);
nor U14844 (N_14844,N_14693,N_14721);
xor U14845 (N_14845,N_14696,N_14734);
nor U14846 (N_14846,N_14540,N_14585);
or U14847 (N_14847,N_14717,N_14592);
nor U14848 (N_14848,N_14712,N_14691);
or U14849 (N_14849,N_14744,N_14735);
or U14850 (N_14850,N_14545,N_14523);
and U14851 (N_14851,N_14714,N_14680);
or U14852 (N_14852,N_14606,N_14577);
xor U14853 (N_14853,N_14700,N_14661);
and U14854 (N_14854,N_14654,N_14534);
or U14855 (N_14855,N_14673,N_14637);
or U14856 (N_14856,N_14579,N_14708);
nor U14857 (N_14857,N_14516,N_14694);
and U14858 (N_14858,N_14528,N_14724);
and U14859 (N_14859,N_14557,N_14568);
xor U14860 (N_14860,N_14695,N_14505);
nor U14861 (N_14861,N_14719,N_14522);
nor U14862 (N_14862,N_14713,N_14544);
or U14863 (N_14863,N_14699,N_14551);
or U14864 (N_14864,N_14705,N_14611);
nor U14865 (N_14865,N_14674,N_14565);
or U14866 (N_14866,N_14715,N_14716);
and U14867 (N_14867,N_14504,N_14653);
and U14868 (N_14868,N_14738,N_14682);
nand U14869 (N_14869,N_14741,N_14552);
or U14870 (N_14870,N_14537,N_14729);
xnor U14871 (N_14871,N_14556,N_14591);
nand U14872 (N_14872,N_14739,N_14576);
nand U14873 (N_14873,N_14530,N_14732);
or U14874 (N_14874,N_14728,N_14555);
nand U14875 (N_14875,N_14600,N_14654);
nor U14876 (N_14876,N_14714,N_14595);
xnor U14877 (N_14877,N_14691,N_14558);
or U14878 (N_14878,N_14578,N_14719);
or U14879 (N_14879,N_14659,N_14519);
xor U14880 (N_14880,N_14601,N_14669);
or U14881 (N_14881,N_14504,N_14620);
nor U14882 (N_14882,N_14680,N_14532);
and U14883 (N_14883,N_14645,N_14727);
or U14884 (N_14884,N_14546,N_14531);
or U14885 (N_14885,N_14623,N_14717);
or U14886 (N_14886,N_14564,N_14669);
or U14887 (N_14887,N_14686,N_14662);
and U14888 (N_14888,N_14522,N_14546);
nor U14889 (N_14889,N_14669,N_14749);
nor U14890 (N_14890,N_14743,N_14522);
nor U14891 (N_14891,N_14728,N_14745);
xor U14892 (N_14892,N_14589,N_14742);
nand U14893 (N_14893,N_14569,N_14511);
or U14894 (N_14894,N_14702,N_14512);
nor U14895 (N_14895,N_14510,N_14644);
nor U14896 (N_14896,N_14746,N_14520);
xor U14897 (N_14897,N_14553,N_14536);
xor U14898 (N_14898,N_14735,N_14725);
nand U14899 (N_14899,N_14723,N_14720);
nor U14900 (N_14900,N_14587,N_14747);
xor U14901 (N_14901,N_14534,N_14700);
nand U14902 (N_14902,N_14515,N_14617);
or U14903 (N_14903,N_14547,N_14607);
nor U14904 (N_14904,N_14598,N_14514);
xor U14905 (N_14905,N_14689,N_14661);
xnor U14906 (N_14906,N_14563,N_14716);
and U14907 (N_14907,N_14710,N_14512);
and U14908 (N_14908,N_14648,N_14689);
xnor U14909 (N_14909,N_14693,N_14537);
nor U14910 (N_14910,N_14624,N_14739);
and U14911 (N_14911,N_14587,N_14628);
or U14912 (N_14912,N_14606,N_14617);
or U14913 (N_14913,N_14606,N_14695);
nor U14914 (N_14914,N_14648,N_14530);
or U14915 (N_14915,N_14635,N_14539);
nor U14916 (N_14916,N_14670,N_14723);
or U14917 (N_14917,N_14542,N_14553);
nand U14918 (N_14918,N_14538,N_14557);
nand U14919 (N_14919,N_14671,N_14520);
nor U14920 (N_14920,N_14746,N_14683);
or U14921 (N_14921,N_14729,N_14736);
xor U14922 (N_14922,N_14536,N_14658);
or U14923 (N_14923,N_14708,N_14711);
nand U14924 (N_14924,N_14700,N_14549);
or U14925 (N_14925,N_14592,N_14560);
and U14926 (N_14926,N_14648,N_14604);
nor U14927 (N_14927,N_14536,N_14693);
or U14928 (N_14928,N_14576,N_14635);
and U14929 (N_14929,N_14506,N_14650);
or U14930 (N_14930,N_14673,N_14526);
nor U14931 (N_14931,N_14618,N_14547);
nand U14932 (N_14932,N_14560,N_14679);
and U14933 (N_14933,N_14559,N_14582);
and U14934 (N_14934,N_14699,N_14610);
or U14935 (N_14935,N_14738,N_14597);
and U14936 (N_14936,N_14535,N_14732);
and U14937 (N_14937,N_14694,N_14638);
and U14938 (N_14938,N_14631,N_14599);
nand U14939 (N_14939,N_14710,N_14749);
and U14940 (N_14940,N_14541,N_14506);
xnor U14941 (N_14941,N_14647,N_14740);
nor U14942 (N_14942,N_14545,N_14522);
and U14943 (N_14943,N_14626,N_14610);
and U14944 (N_14944,N_14569,N_14561);
nand U14945 (N_14945,N_14623,N_14504);
nand U14946 (N_14946,N_14715,N_14536);
nor U14947 (N_14947,N_14622,N_14703);
nor U14948 (N_14948,N_14506,N_14668);
nand U14949 (N_14949,N_14585,N_14530);
or U14950 (N_14950,N_14616,N_14513);
nor U14951 (N_14951,N_14535,N_14671);
and U14952 (N_14952,N_14630,N_14522);
nand U14953 (N_14953,N_14661,N_14718);
xor U14954 (N_14954,N_14515,N_14525);
xor U14955 (N_14955,N_14502,N_14704);
and U14956 (N_14956,N_14608,N_14626);
nor U14957 (N_14957,N_14704,N_14731);
nor U14958 (N_14958,N_14546,N_14550);
nor U14959 (N_14959,N_14561,N_14593);
nand U14960 (N_14960,N_14691,N_14541);
xor U14961 (N_14961,N_14682,N_14723);
or U14962 (N_14962,N_14526,N_14682);
and U14963 (N_14963,N_14744,N_14633);
nor U14964 (N_14964,N_14504,N_14508);
or U14965 (N_14965,N_14597,N_14623);
xor U14966 (N_14966,N_14546,N_14610);
and U14967 (N_14967,N_14746,N_14527);
nor U14968 (N_14968,N_14582,N_14671);
xnor U14969 (N_14969,N_14641,N_14664);
xor U14970 (N_14970,N_14528,N_14698);
xor U14971 (N_14971,N_14505,N_14534);
and U14972 (N_14972,N_14604,N_14568);
xnor U14973 (N_14973,N_14729,N_14502);
xnor U14974 (N_14974,N_14501,N_14588);
xor U14975 (N_14975,N_14601,N_14686);
or U14976 (N_14976,N_14620,N_14746);
nand U14977 (N_14977,N_14500,N_14735);
nand U14978 (N_14978,N_14698,N_14639);
or U14979 (N_14979,N_14685,N_14671);
or U14980 (N_14980,N_14596,N_14707);
or U14981 (N_14981,N_14659,N_14588);
nand U14982 (N_14982,N_14536,N_14722);
nand U14983 (N_14983,N_14642,N_14503);
nand U14984 (N_14984,N_14686,N_14528);
nor U14985 (N_14985,N_14506,N_14611);
nor U14986 (N_14986,N_14611,N_14729);
or U14987 (N_14987,N_14734,N_14632);
or U14988 (N_14988,N_14704,N_14566);
nand U14989 (N_14989,N_14517,N_14636);
and U14990 (N_14990,N_14531,N_14623);
nor U14991 (N_14991,N_14558,N_14588);
nand U14992 (N_14992,N_14674,N_14571);
nand U14993 (N_14993,N_14561,N_14700);
xor U14994 (N_14994,N_14712,N_14620);
and U14995 (N_14995,N_14601,N_14681);
and U14996 (N_14996,N_14735,N_14527);
xor U14997 (N_14997,N_14603,N_14578);
and U14998 (N_14998,N_14509,N_14667);
or U14999 (N_14999,N_14714,N_14544);
or U15000 (N_15000,N_14876,N_14991);
nor U15001 (N_15001,N_14951,N_14999);
nand U15002 (N_15002,N_14888,N_14752);
and U15003 (N_15003,N_14887,N_14769);
nor U15004 (N_15004,N_14943,N_14911);
and U15005 (N_15005,N_14789,N_14976);
nor U15006 (N_15006,N_14962,N_14864);
nor U15007 (N_15007,N_14900,N_14776);
or U15008 (N_15008,N_14934,N_14880);
and U15009 (N_15009,N_14803,N_14751);
nand U15010 (N_15010,N_14874,N_14759);
xnor U15011 (N_15011,N_14926,N_14758);
or U15012 (N_15012,N_14784,N_14891);
xor U15013 (N_15013,N_14822,N_14760);
nand U15014 (N_15014,N_14956,N_14937);
nand U15015 (N_15015,N_14850,N_14901);
or U15016 (N_15016,N_14990,N_14871);
xnor U15017 (N_15017,N_14809,N_14863);
or U15018 (N_15018,N_14851,N_14969);
and U15019 (N_15019,N_14807,N_14763);
nor U15020 (N_15020,N_14836,N_14989);
nor U15021 (N_15021,N_14987,N_14774);
xnor U15022 (N_15022,N_14772,N_14862);
nor U15023 (N_15023,N_14840,N_14998);
xor U15024 (N_15024,N_14843,N_14810);
nand U15025 (N_15025,N_14896,N_14849);
nor U15026 (N_15026,N_14771,N_14980);
nor U15027 (N_15027,N_14915,N_14750);
and U15028 (N_15028,N_14928,N_14783);
nand U15029 (N_15029,N_14908,N_14964);
nand U15030 (N_15030,N_14965,N_14775);
and U15031 (N_15031,N_14952,N_14977);
or U15032 (N_15032,N_14885,N_14860);
or U15033 (N_15033,N_14873,N_14892);
nor U15034 (N_15034,N_14968,N_14975);
xor U15035 (N_15035,N_14893,N_14766);
xnor U15036 (N_15036,N_14800,N_14986);
and U15037 (N_15037,N_14857,N_14815);
and U15038 (N_15038,N_14811,N_14886);
nand U15039 (N_15039,N_14914,N_14827);
nor U15040 (N_15040,N_14897,N_14870);
nand U15041 (N_15041,N_14755,N_14853);
or U15042 (N_15042,N_14808,N_14921);
xnor U15043 (N_15043,N_14875,N_14916);
nand U15044 (N_15044,N_14912,N_14757);
or U15045 (N_15045,N_14942,N_14983);
and U15046 (N_15046,N_14780,N_14785);
xnor U15047 (N_15047,N_14872,N_14884);
xnor U15048 (N_15048,N_14765,N_14971);
nand U15049 (N_15049,N_14985,N_14996);
xnor U15050 (N_15050,N_14802,N_14868);
nand U15051 (N_15051,N_14754,N_14756);
nor U15052 (N_15052,N_14944,N_14818);
or U15053 (N_15053,N_14878,N_14833);
nand U15054 (N_15054,N_14922,N_14830);
xnor U15055 (N_15055,N_14966,N_14813);
or U15056 (N_15056,N_14779,N_14856);
xnor U15057 (N_15057,N_14954,N_14817);
nor U15058 (N_15058,N_14814,N_14931);
or U15059 (N_15059,N_14824,N_14826);
nor U15060 (N_15060,N_14795,N_14903);
nor U15061 (N_15061,N_14941,N_14907);
and U15062 (N_15062,N_14787,N_14819);
or U15063 (N_15063,N_14778,N_14994);
or U15064 (N_15064,N_14805,N_14923);
and U15065 (N_15065,N_14812,N_14890);
xor U15066 (N_15066,N_14919,N_14790);
xnor U15067 (N_15067,N_14777,N_14957);
nand U15068 (N_15068,N_14770,N_14904);
xnor U15069 (N_15069,N_14793,N_14792);
xnor U15070 (N_15070,N_14804,N_14972);
nand U15071 (N_15071,N_14806,N_14825);
nor U15072 (N_15072,N_14978,N_14913);
nor U15073 (N_15073,N_14859,N_14883);
xnor U15074 (N_15074,N_14847,N_14895);
xnor U15075 (N_15075,N_14981,N_14762);
and U15076 (N_15076,N_14835,N_14988);
and U15077 (N_15077,N_14917,N_14918);
or U15078 (N_15078,N_14781,N_14973);
xor U15079 (N_15079,N_14861,N_14961);
nor U15080 (N_15080,N_14949,N_14848);
or U15081 (N_15081,N_14905,N_14828);
or U15082 (N_15082,N_14950,N_14858);
or U15083 (N_15083,N_14829,N_14982);
xor U15084 (N_15084,N_14796,N_14764);
or U15085 (N_15085,N_14970,N_14823);
or U15086 (N_15086,N_14798,N_14995);
nor U15087 (N_15087,N_14816,N_14993);
or U15088 (N_15088,N_14909,N_14910);
nor U15089 (N_15089,N_14938,N_14834);
and U15090 (N_15090,N_14935,N_14906);
xor U15091 (N_15091,N_14933,N_14867);
nand U15092 (N_15092,N_14929,N_14947);
xnor U15093 (N_15093,N_14974,N_14788);
nor U15094 (N_15094,N_14997,N_14955);
and U15095 (N_15095,N_14940,N_14794);
and U15096 (N_15096,N_14846,N_14761);
and U15097 (N_15097,N_14920,N_14902);
and U15098 (N_15098,N_14753,N_14924);
nor U15099 (N_15099,N_14967,N_14979);
or U15100 (N_15100,N_14899,N_14960);
xor U15101 (N_15101,N_14821,N_14773);
nor U15102 (N_15102,N_14894,N_14854);
xnor U15103 (N_15103,N_14939,N_14838);
nand U15104 (N_15104,N_14865,N_14946);
nand U15105 (N_15105,N_14932,N_14936);
xnor U15106 (N_15106,N_14882,N_14845);
nor U15107 (N_15107,N_14786,N_14832);
xnor U15108 (N_15108,N_14799,N_14992);
nand U15109 (N_15109,N_14898,N_14984);
nor U15110 (N_15110,N_14958,N_14945);
nand U15111 (N_15111,N_14852,N_14855);
xnor U15112 (N_15112,N_14963,N_14767);
nand U15113 (N_15113,N_14881,N_14889);
or U15114 (N_15114,N_14791,N_14877);
or U15115 (N_15115,N_14768,N_14927);
and U15116 (N_15116,N_14842,N_14837);
and U15117 (N_15117,N_14866,N_14925);
or U15118 (N_15118,N_14841,N_14953);
or U15119 (N_15119,N_14782,N_14839);
and U15120 (N_15120,N_14844,N_14820);
or U15121 (N_15121,N_14797,N_14801);
xnor U15122 (N_15122,N_14879,N_14831);
or U15123 (N_15123,N_14959,N_14948);
or U15124 (N_15124,N_14930,N_14869);
or U15125 (N_15125,N_14975,N_14802);
or U15126 (N_15126,N_14827,N_14776);
xnor U15127 (N_15127,N_14780,N_14790);
nor U15128 (N_15128,N_14945,N_14796);
or U15129 (N_15129,N_14979,N_14898);
or U15130 (N_15130,N_14931,N_14947);
nand U15131 (N_15131,N_14930,N_14872);
or U15132 (N_15132,N_14975,N_14825);
and U15133 (N_15133,N_14870,N_14997);
and U15134 (N_15134,N_14995,N_14892);
nand U15135 (N_15135,N_14925,N_14909);
nand U15136 (N_15136,N_14757,N_14924);
xnor U15137 (N_15137,N_14863,N_14940);
nand U15138 (N_15138,N_14878,N_14951);
nor U15139 (N_15139,N_14880,N_14972);
nor U15140 (N_15140,N_14944,N_14972);
and U15141 (N_15141,N_14907,N_14811);
nor U15142 (N_15142,N_14952,N_14930);
or U15143 (N_15143,N_14825,N_14860);
xnor U15144 (N_15144,N_14849,N_14889);
xnor U15145 (N_15145,N_14991,N_14996);
or U15146 (N_15146,N_14750,N_14875);
or U15147 (N_15147,N_14871,N_14946);
xnor U15148 (N_15148,N_14989,N_14958);
xor U15149 (N_15149,N_14954,N_14843);
or U15150 (N_15150,N_14911,N_14965);
and U15151 (N_15151,N_14957,N_14993);
nor U15152 (N_15152,N_14817,N_14980);
xnor U15153 (N_15153,N_14921,N_14898);
and U15154 (N_15154,N_14858,N_14780);
or U15155 (N_15155,N_14846,N_14793);
xor U15156 (N_15156,N_14820,N_14971);
nand U15157 (N_15157,N_14995,N_14994);
and U15158 (N_15158,N_14756,N_14824);
xor U15159 (N_15159,N_14899,N_14999);
xor U15160 (N_15160,N_14944,N_14812);
or U15161 (N_15161,N_14840,N_14809);
nand U15162 (N_15162,N_14906,N_14828);
nand U15163 (N_15163,N_14763,N_14766);
and U15164 (N_15164,N_14835,N_14920);
nor U15165 (N_15165,N_14911,N_14923);
nand U15166 (N_15166,N_14824,N_14777);
nand U15167 (N_15167,N_14998,N_14996);
nor U15168 (N_15168,N_14854,N_14919);
xor U15169 (N_15169,N_14900,N_14860);
xor U15170 (N_15170,N_14944,N_14974);
and U15171 (N_15171,N_14906,N_14835);
and U15172 (N_15172,N_14783,N_14755);
and U15173 (N_15173,N_14841,N_14967);
and U15174 (N_15174,N_14845,N_14771);
nand U15175 (N_15175,N_14914,N_14785);
and U15176 (N_15176,N_14940,N_14758);
nor U15177 (N_15177,N_14943,N_14803);
xor U15178 (N_15178,N_14750,N_14784);
and U15179 (N_15179,N_14796,N_14918);
and U15180 (N_15180,N_14972,N_14963);
xnor U15181 (N_15181,N_14934,N_14929);
or U15182 (N_15182,N_14822,N_14888);
nor U15183 (N_15183,N_14821,N_14916);
or U15184 (N_15184,N_14767,N_14793);
or U15185 (N_15185,N_14980,N_14908);
and U15186 (N_15186,N_14883,N_14825);
nor U15187 (N_15187,N_14874,N_14796);
or U15188 (N_15188,N_14987,N_14815);
xor U15189 (N_15189,N_14773,N_14933);
xnor U15190 (N_15190,N_14971,N_14900);
or U15191 (N_15191,N_14910,N_14799);
nand U15192 (N_15192,N_14884,N_14921);
xnor U15193 (N_15193,N_14857,N_14753);
nor U15194 (N_15194,N_14988,N_14789);
nand U15195 (N_15195,N_14814,N_14810);
nand U15196 (N_15196,N_14766,N_14832);
and U15197 (N_15197,N_14884,N_14815);
nand U15198 (N_15198,N_14897,N_14968);
xnor U15199 (N_15199,N_14915,N_14879);
xnor U15200 (N_15200,N_14751,N_14768);
and U15201 (N_15201,N_14757,N_14803);
and U15202 (N_15202,N_14775,N_14884);
nand U15203 (N_15203,N_14905,N_14937);
and U15204 (N_15204,N_14981,N_14911);
xor U15205 (N_15205,N_14902,N_14911);
and U15206 (N_15206,N_14892,N_14828);
xnor U15207 (N_15207,N_14945,N_14869);
nor U15208 (N_15208,N_14876,N_14782);
or U15209 (N_15209,N_14964,N_14850);
xor U15210 (N_15210,N_14954,N_14847);
nand U15211 (N_15211,N_14988,N_14991);
nor U15212 (N_15212,N_14919,N_14782);
nand U15213 (N_15213,N_14942,N_14777);
nor U15214 (N_15214,N_14811,N_14786);
xor U15215 (N_15215,N_14898,N_14879);
or U15216 (N_15216,N_14989,N_14979);
nand U15217 (N_15217,N_14872,N_14900);
or U15218 (N_15218,N_14969,N_14830);
or U15219 (N_15219,N_14867,N_14914);
nor U15220 (N_15220,N_14884,N_14968);
nor U15221 (N_15221,N_14877,N_14842);
or U15222 (N_15222,N_14784,N_14843);
nor U15223 (N_15223,N_14751,N_14798);
nor U15224 (N_15224,N_14911,N_14884);
nor U15225 (N_15225,N_14853,N_14869);
nand U15226 (N_15226,N_14934,N_14827);
nand U15227 (N_15227,N_14938,N_14933);
and U15228 (N_15228,N_14757,N_14868);
nand U15229 (N_15229,N_14964,N_14963);
nand U15230 (N_15230,N_14864,N_14880);
and U15231 (N_15231,N_14898,N_14914);
or U15232 (N_15232,N_14895,N_14890);
xor U15233 (N_15233,N_14999,N_14856);
nor U15234 (N_15234,N_14813,N_14854);
xnor U15235 (N_15235,N_14777,N_14941);
xnor U15236 (N_15236,N_14988,N_14883);
and U15237 (N_15237,N_14902,N_14806);
and U15238 (N_15238,N_14908,N_14924);
nor U15239 (N_15239,N_14916,N_14959);
nand U15240 (N_15240,N_14767,N_14817);
nor U15241 (N_15241,N_14847,N_14796);
and U15242 (N_15242,N_14766,N_14816);
nand U15243 (N_15243,N_14845,N_14805);
and U15244 (N_15244,N_14840,N_14881);
nor U15245 (N_15245,N_14929,N_14974);
nor U15246 (N_15246,N_14873,N_14841);
xor U15247 (N_15247,N_14771,N_14880);
and U15248 (N_15248,N_14996,N_14774);
and U15249 (N_15249,N_14974,N_14825);
nor U15250 (N_15250,N_15050,N_15128);
or U15251 (N_15251,N_15076,N_15136);
or U15252 (N_15252,N_15150,N_15183);
nand U15253 (N_15253,N_15083,N_15234);
xnor U15254 (N_15254,N_15225,N_15160);
and U15255 (N_15255,N_15206,N_15187);
nor U15256 (N_15256,N_15176,N_15228);
and U15257 (N_15257,N_15079,N_15027);
or U15258 (N_15258,N_15243,N_15064);
nor U15259 (N_15259,N_15115,N_15196);
xor U15260 (N_15260,N_15000,N_15048);
nand U15261 (N_15261,N_15151,N_15034);
xnor U15262 (N_15262,N_15120,N_15114);
nand U15263 (N_15263,N_15057,N_15152);
xor U15264 (N_15264,N_15017,N_15090);
or U15265 (N_15265,N_15061,N_15153);
nor U15266 (N_15266,N_15155,N_15179);
xor U15267 (N_15267,N_15210,N_15085);
nand U15268 (N_15268,N_15108,N_15242);
xor U15269 (N_15269,N_15220,N_15065);
xnor U15270 (N_15270,N_15149,N_15002);
and U15271 (N_15271,N_15224,N_15107);
or U15272 (N_15272,N_15036,N_15014);
nor U15273 (N_15273,N_15025,N_15172);
nand U15274 (N_15274,N_15109,N_15135);
or U15275 (N_15275,N_15087,N_15181);
and U15276 (N_15276,N_15247,N_15103);
or U15277 (N_15277,N_15043,N_15200);
or U15278 (N_15278,N_15195,N_15197);
nor U15279 (N_15279,N_15012,N_15023);
and U15280 (N_15280,N_15189,N_15163);
or U15281 (N_15281,N_15072,N_15161);
nor U15282 (N_15282,N_15063,N_15098);
nor U15283 (N_15283,N_15067,N_15030);
and U15284 (N_15284,N_15159,N_15170);
nor U15285 (N_15285,N_15223,N_15029);
or U15286 (N_15286,N_15049,N_15068);
or U15287 (N_15287,N_15095,N_15248);
nand U15288 (N_15288,N_15040,N_15209);
xnor U15289 (N_15289,N_15028,N_15102);
nand U15290 (N_15290,N_15190,N_15033);
xnor U15291 (N_15291,N_15022,N_15227);
nor U15292 (N_15292,N_15171,N_15073);
nand U15293 (N_15293,N_15211,N_15217);
xnor U15294 (N_15294,N_15003,N_15111);
or U15295 (N_15295,N_15021,N_15164);
nor U15296 (N_15296,N_15180,N_15041);
and U15297 (N_15297,N_15123,N_15016);
and U15298 (N_15298,N_15047,N_15100);
or U15299 (N_15299,N_15237,N_15019);
nand U15300 (N_15300,N_15031,N_15140);
and U15301 (N_15301,N_15056,N_15122);
and U15302 (N_15302,N_15071,N_15020);
or U15303 (N_15303,N_15055,N_15167);
or U15304 (N_15304,N_15001,N_15238);
or U15305 (N_15305,N_15130,N_15219);
and U15306 (N_15306,N_15093,N_15142);
or U15307 (N_15307,N_15013,N_15112);
or U15308 (N_15308,N_15094,N_15202);
and U15309 (N_15309,N_15024,N_15044);
or U15310 (N_15310,N_15015,N_15010);
nor U15311 (N_15311,N_15166,N_15138);
or U15312 (N_15312,N_15080,N_15101);
and U15313 (N_15313,N_15091,N_15125);
nand U15314 (N_15314,N_15208,N_15204);
xor U15315 (N_15315,N_15099,N_15221);
xor U15316 (N_15316,N_15239,N_15193);
xor U15317 (N_15317,N_15032,N_15215);
and U15318 (N_15318,N_15139,N_15053);
nor U15319 (N_15319,N_15185,N_15086);
xor U15320 (N_15320,N_15232,N_15046);
nor U15321 (N_15321,N_15203,N_15124);
nor U15322 (N_15322,N_15045,N_15133);
nand U15323 (N_15323,N_15005,N_15070);
xnor U15324 (N_15324,N_15245,N_15145);
and U15325 (N_15325,N_15104,N_15110);
nor U15326 (N_15326,N_15188,N_15077);
xnor U15327 (N_15327,N_15198,N_15134);
xor U15328 (N_15328,N_15121,N_15052);
nand U15329 (N_15329,N_15218,N_15214);
nor U15330 (N_15330,N_15144,N_15141);
xor U15331 (N_15331,N_15222,N_15117);
and U15332 (N_15332,N_15075,N_15199);
nor U15333 (N_15333,N_15236,N_15231);
or U15334 (N_15334,N_15059,N_15213);
nor U15335 (N_15335,N_15186,N_15146);
nand U15336 (N_15336,N_15182,N_15039);
xnor U15337 (N_15337,N_15246,N_15212);
and U15338 (N_15338,N_15168,N_15233);
nor U15339 (N_15339,N_15105,N_15051);
or U15340 (N_15340,N_15060,N_15165);
nor U15341 (N_15341,N_15088,N_15174);
nand U15342 (N_15342,N_15240,N_15192);
nand U15343 (N_15343,N_15018,N_15092);
nor U15344 (N_15344,N_15035,N_15084);
or U15345 (N_15345,N_15129,N_15173);
or U15346 (N_15346,N_15078,N_15184);
nand U15347 (N_15347,N_15096,N_15177);
and U15348 (N_15348,N_15131,N_15201);
and U15349 (N_15349,N_15158,N_15169);
nand U15350 (N_15350,N_15241,N_15244);
and U15351 (N_15351,N_15037,N_15042);
and U15352 (N_15352,N_15226,N_15074);
nor U15353 (N_15353,N_15007,N_15006);
or U15354 (N_15354,N_15147,N_15106);
or U15355 (N_15355,N_15229,N_15066);
nand U15356 (N_15356,N_15156,N_15194);
nor U15357 (N_15357,N_15097,N_15126);
xnor U15358 (N_15358,N_15008,N_15157);
nand U15359 (N_15359,N_15132,N_15162);
and U15360 (N_15360,N_15054,N_15235);
nor U15361 (N_15361,N_15191,N_15089);
nand U15362 (N_15362,N_15249,N_15216);
nand U15363 (N_15363,N_15009,N_15143);
xnor U15364 (N_15364,N_15178,N_15118);
nand U15365 (N_15365,N_15207,N_15058);
and U15366 (N_15366,N_15062,N_15081);
xor U15367 (N_15367,N_15004,N_15119);
and U15368 (N_15368,N_15230,N_15026);
and U15369 (N_15369,N_15127,N_15011);
or U15370 (N_15370,N_15148,N_15082);
nand U15371 (N_15371,N_15137,N_15205);
nor U15372 (N_15372,N_15069,N_15038);
nor U15373 (N_15373,N_15154,N_15116);
nor U15374 (N_15374,N_15175,N_15113);
xor U15375 (N_15375,N_15220,N_15070);
or U15376 (N_15376,N_15073,N_15016);
xor U15377 (N_15377,N_15055,N_15210);
or U15378 (N_15378,N_15200,N_15215);
xnor U15379 (N_15379,N_15097,N_15110);
or U15380 (N_15380,N_15117,N_15154);
or U15381 (N_15381,N_15064,N_15170);
nand U15382 (N_15382,N_15033,N_15174);
nand U15383 (N_15383,N_15149,N_15021);
or U15384 (N_15384,N_15039,N_15101);
nor U15385 (N_15385,N_15133,N_15192);
and U15386 (N_15386,N_15238,N_15024);
nor U15387 (N_15387,N_15088,N_15099);
xnor U15388 (N_15388,N_15120,N_15045);
nand U15389 (N_15389,N_15076,N_15090);
xor U15390 (N_15390,N_15207,N_15214);
nor U15391 (N_15391,N_15034,N_15043);
nand U15392 (N_15392,N_15057,N_15185);
or U15393 (N_15393,N_15064,N_15008);
nor U15394 (N_15394,N_15057,N_15033);
nor U15395 (N_15395,N_15070,N_15195);
xor U15396 (N_15396,N_15115,N_15162);
and U15397 (N_15397,N_15247,N_15224);
xnor U15398 (N_15398,N_15086,N_15054);
or U15399 (N_15399,N_15067,N_15047);
nor U15400 (N_15400,N_15159,N_15151);
and U15401 (N_15401,N_15124,N_15100);
and U15402 (N_15402,N_15145,N_15161);
xor U15403 (N_15403,N_15062,N_15121);
xor U15404 (N_15404,N_15007,N_15146);
nand U15405 (N_15405,N_15156,N_15171);
xnor U15406 (N_15406,N_15195,N_15076);
nor U15407 (N_15407,N_15053,N_15080);
or U15408 (N_15408,N_15019,N_15109);
nand U15409 (N_15409,N_15075,N_15179);
nor U15410 (N_15410,N_15143,N_15025);
xnor U15411 (N_15411,N_15119,N_15104);
or U15412 (N_15412,N_15086,N_15146);
xnor U15413 (N_15413,N_15194,N_15114);
or U15414 (N_15414,N_15129,N_15078);
nor U15415 (N_15415,N_15142,N_15243);
and U15416 (N_15416,N_15175,N_15243);
nand U15417 (N_15417,N_15138,N_15165);
nand U15418 (N_15418,N_15215,N_15244);
nand U15419 (N_15419,N_15125,N_15011);
nor U15420 (N_15420,N_15242,N_15050);
nor U15421 (N_15421,N_15111,N_15117);
and U15422 (N_15422,N_15064,N_15067);
and U15423 (N_15423,N_15158,N_15045);
nor U15424 (N_15424,N_15112,N_15054);
or U15425 (N_15425,N_15006,N_15132);
nand U15426 (N_15426,N_15039,N_15134);
xor U15427 (N_15427,N_15046,N_15106);
nor U15428 (N_15428,N_15042,N_15168);
xnor U15429 (N_15429,N_15042,N_15172);
and U15430 (N_15430,N_15024,N_15136);
and U15431 (N_15431,N_15099,N_15153);
xor U15432 (N_15432,N_15235,N_15140);
and U15433 (N_15433,N_15091,N_15094);
nand U15434 (N_15434,N_15164,N_15200);
nand U15435 (N_15435,N_15067,N_15033);
or U15436 (N_15436,N_15214,N_15189);
and U15437 (N_15437,N_15056,N_15005);
or U15438 (N_15438,N_15136,N_15214);
nor U15439 (N_15439,N_15163,N_15012);
xor U15440 (N_15440,N_15187,N_15145);
xnor U15441 (N_15441,N_15080,N_15227);
nor U15442 (N_15442,N_15019,N_15046);
xor U15443 (N_15443,N_15111,N_15078);
nor U15444 (N_15444,N_15014,N_15069);
xor U15445 (N_15445,N_15043,N_15070);
and U15446 (N_15446,N_15093,N_15104);
and U15447 (N_15447,N_15198,N_15104);
xor U15448 (N_15448,N_15055,N_15091);
xor U15449 (N_15449,N_15103,N_15149);
xor U15450 (N_15450,N_15190,N_15203);
and U15451 (N_15451,N_15176,N_15020);
and U15452 (N_15452,N_15169,N_15165);
and U15453 (N_15453,N_15156,N_15054);
nor U15454 (N_15454,N_15232,N_15022);
or U15455 (N_15455,N_15173,N_15085);
or U15456 (N_15456,N_15001,N_15153);
and U15457 (N_15457,N_15177,N_15160);
and U15458 (N_15458,N_15141,N_15104);
or U15459 (N_15459,N_15193,N_15142);
or U15460 (N_15460,N_15088,N_15010);
or U15461 (N_15461,N_15214,N_15040);
nor U15462 (N_15462,N_15154,N_15127);
or U15463 (N_15463,N_15013,N_15246);
nand U15464 (N_15464,N_15233,N_15222);
xnor U15465 (N_15465,N_15133,N_15042);
nand U15466 (N_15466,N_15031,N_15245);
xnor U15467 (N_15467,N_15208,N_15215);
nand U15468 (N_15468,N_15240,N_15128);
or U15469 (N_15469,N_15132,N_15067);
nor U15470 (N_15470,N_15056,N_15127);
and U15471 (N_15471,N_15150,N_15092);
nand U15472 (N_15472,N_15120,N_15004);
nor U15473 (N_15473,N_15209,N_15163);
nor U15474 (N_15474,N_15106,N_15085);
and U15475 (N_15475,N_15133,N_15217);
xor U15476 (N_15476,N_15048,N_15166);
nand U15477 (N_15477,N_15022,N_15059);
or U15478 (N_15478,N_15213,N_15124);
xnor U15479 (N_15479,N_15019,N_15004);
or U15480 (N_15480,N_15042,N_15066);
nor U15481 (N_15481,N_15104,N_15037);
or U15482 (N_15482,N_15186,N_15234);
nor U15483 (N_15483,N_15064,N_15222);
and U15484 (N_15484,N_15143,N_15168);
nand U15485 (N_15485,N_15039,N_15048);
nor U15486 (N_15486,N_15186,N_15110);
xnor U15487 (N_15487,N_15223,N_15214);
nand U15488 (N_15488,N_15238,N_15143);
nor U15489 (N_15489,N_15241,N_15228);
xor U15490 (N_15490,N_15243,N_15232);
nand U15491 (N_15491,N_15028,N_15109);
nand U15492 (N_15492,N_15122,N_15040);
nor U15493 (N_15493,N_15114,N_15025);
nor U15494 (N_15494,N_15087,N_15124);
and U15495 (N_15495,N_15249,N_15096);
or U15496 (N_15496,N_15073,N_15022);
xnor U15497 (N_15497,N_15162,N_15059);
nor U15498 (N_15498,N_15047,N_15146);
or U15499 (N_15499,N_15141,N_15146);
and U15500 (N_15500,N_15323,N_15479);
nor U15501 (N_15501,N_15289,N_15465);
xor U15502 (N_15502,N_15261,N_15435);
and U15503 (N_15503,N_15287,N_15316);
nor U15504 (N_15504,N_15495,N_15278);
nor U15505 (N_15505,N_15478,N_15284);
nor U15506 (N_15506,N_15449,N_15416);
xor U15507 (N_15507,N_15496,N_15457);
xor U15508 (N_15508,N_15471,N_15336);
nor U15509 (N_15509,N_15485,N_15262);
nand U15510 (N_15510,N_15480,N_15353);
or U15511 (N_15511,N_15283,N_15327);
nor U15512 (N_15512,N_15406,N_15442);
nor U15513 (N_15513,N_15330,N_15476);
xnor U15514 (N_15514,N_15251,N_15418);
nand U15515 (N_15515,N_15466,N_15384);
and U15516 (N_15516,N_15264,N_15266);
xor U15517 (N_15517,N_15301,N_15302);
nor U15518 (N_15518,N_15324,N_15374);
xnor U15519 (N_15519,N_15426,N_15344);
and U15520 (N_15520,N_15482,N_15447);
and U15521 (N_15521,N_15497,N_15407);
and U15522 (N_15522,N_15420,N_15409);
nand U15523 (N_15523,N_15320,N_15272);
xnor U15524 (N_15524,N_15455,N_15366);
xnor U15525 (N_15525,N_15399,N_15440);
or U15526 (N_15526,N_15326,N_15292);
or U15527 (N_15527,N_15333,N_15490);
nor U15528 (N_15528,N_15367,N_15267);
nor U15529 (N_15529,N_15335,N_15310);
nand U15530 (N_15530,N_15297,N_15321);
and U15531 (N_15531,N_15257,N_15389);
nand U15532 (N_15532,N_15376,N_15274);
or U15533 (N_15533,N_15358,N_15488);
and U15534 (N_15534,N_15347,N_15296);
nor U15535 (N_15535,N_15454,N_15360);
nor U15536 (N_15536,N_15393,N_15467);
xnor U15537 (N_15537,N_15390,N_15470);
and U15538 (N_15538,N_15325,N_15487);
nand U15539 (N_15539,N_15370,N_15263);
nand U15540 (N_15540,N_15355,N_15252);
or U15541 (N_15541,N_15365,N_15295);
nand U15542 (N_15542,N_15439,N_15432);
nand U15543 (N_15543,N_15411,N_15469);
and U15544 (N_15544,N_15437,N_15332);
xnor U15545 (N_15545,N_15340,N_15375);
xor U15546 (N_15546,N_15254,N_15275);
or U15547 (N_15547,N_15304,N_15391);
xor U15548 (N_15548,N_15342,N_15423);
nor U15549 (N_15549,N_15308,N_15452);
and U15550 (N_15550,N_15349,N_15293);
and U15551 (N_15551,N_15460,N_15265);
xnor U15552 (N_15552,N_15413,N_15373);
xor U15553 (N_15553,N_15408,N_15313);
and U15554 (N_15554,N_15346,N_15392);
or U15555 (N_15555,N_15419,N_15291);
nand U15556 (N_15556,N_15491,N_15428);
and U15557 (N_15557,N_15403,N_15446);
or U15558 (N_15558,N_15282,N_15378);
xnor U15559 (N_15559,N_15362,N_15410);
nor U15560 (N_15560,N_15357,N_15350);
and U15561 (N_15561,N_15276,N_15493);
or U15562 (N_15562,N_15461,N_15288);
nor U15563 (N_15563,N_15329,N_15422);
and U15564 (N_15564,N_15381,N_15377);
xor U15565 (N_15565,N_15369,N_15337);
xnor U15566 (N_15566,N_15430,N_15394);
or U15567 (N_15567,N_15315,N_15489);
nand U15568 (N_15568,N_15398,N_15352);
and U15569 (N_15569,N_15273,N_15281);
and U15570 (N_15570,N_15492,N_15290);
xnor U15571 (N_15571,N_15277,N_15402);
nand U15572 (N_15572,N_15431,N_15280);
nand U15573 (N_15573,N_15382,N_15359);
xor U15574 (N_15574,N_15303,N_15451);
or U15575 (N_15575,N_15429,N_15400);
and U15576 (N_15576,N_15345,N_15339);
or U15577 (N_15577,N_15269,N_15404);
and U15578 (N_15578,N_15448,N_15363);
and U15579 (N_15579,N_15380,N_15425);
nor U15580 (N_15580,N_15361,N_15341);
nand U15581 (N_15581,N_15453,N_15328);
nand U15582 (N_15582,N_15364,N_15436);
or U15583 (N_15583,N_15401,N_15309);
xor U15584 (N_15584,N_15294,N_15270);
or U15585 (N_15585,N_15307,N_15322);
nand U15586 (N_15586,N_15434,N_15319);
nor U15587 (N_15587,N_15463,N_15286);
or U15588 (N_15588,N_15474,N_15458);
or U15589 (N_15589,N_15483,N_15486);
nand U15590 (N_15590,N_15395,N_15405);
nand U15591 (N_15591,N_15334,N_15268);
nand U15592 (N_15592,N_15312,N_15379);
xnor U15593 (N_15593,N_15477,N_15424);
xnor U15594 (N_15594,N_15468,N_15368);
and U15595 (N_15595,N_15300,N_15250);
and U15596 (N_15596,N_15417,N_15433);
nand U15597 (N_15597,N_15255,N_15412);
and U15598 (N_15598,N_15338,N_15414);
nor U15599 (N_15599,N_15371,N_15481);
or U15600 (N_15600,N_15271,N_15443);
xnor U15601 (N_15601,N_15298,N_15258);
or U15602 (N_15602,N_15317,N_15450);
or U15603 (N_15603,N_15259,N_15260);
nand U15604 (N_15604,N_15462,N_15385);
or U15605 (N_15605,N_15415,N_15318);
or U15606 (N_15606,N_15459,N_15331);
nor U15607 (N_15607,N_15285,N_15456);
and U15608 (N_15608,N_15475,N_15472);
and U15609 (N_15609,N_15348,N_15305);
nand U15610 (N_15610,N_15306,N_15354);
or U15611 (N_15611,N_15311,N_15299);
or U15612 (N_15612,N_15484,N_15494);
xnor U15613 (N_15613,N_15445,N_15383);
or U15614 (N_15614,N_15372,N_15438);
xnor U15615 (N_15615,N_15386,N_15498);
xnor U15616 (N_15616,N_15396,N_15499);
nor U15617 (N_15617,N_15397,N_15253);
or U15618 (N_15618,N_15343,N_15387);
nor U15619 (N_15619,N_15441,N_15279);
xor U15620 (N_15620,N_15256,N_15444);
xnor U15621 (N_15621,N_15464,N_15421);
or U15622 (N_15622,N_15356,N_15473);
nor U15623 (N_15623,N_15314,N_15351);
and U15624 (N_15624,N_15388,N_15427);
nor U15625 (N_15625,N_15361,N_15262);
or U15626 (N_15626,N_15357,N_15315);
nand U15627 (N_15627,N_15300,N_15363);
nor U15628 (N_15628,N_15352,N_15337);
and U15629 (N_15629,N_15391,N_15453);
xnor U15630 (N_15630,N_15498,N_15288);
nor U15631 (N_15631,N_15428,N_15443);
or U15632 (N_15632,N_15429,N_15263);
or U15633 (N_15633,N_15414,N_15352);
nor U15634 (N_15634,N_15473,N_15457);
and U15635 (N_15635,N_15310,N_15479);
nor U15636 (N_15636,N_15291,N_15383);
xnor U15637 (N_15637,N_15449,N_15443);
nor U15638 (N_15638,N_15376,N_15456);
nor U15639 (N_15639,N_15407,N_15427);
and U15640 (N_15640,N_15370,N_15472);
xnor U15641 (N_15641,N_15304,N_15384);
nand U15642 (N_15642,N_15374,N_15432);
or U15643 (N_15643,N_15408,N_15341);
or U15644 (N_15644,N_15451,N_15344);
nand U15645 (N_15645,N_15468,N_15355);
and U15646 (N_15646,N_15321,N_15306);
xnor U15647 (N_15647,N_15489,N_15320);
or U15648 (N_15648,N_15416,N_15451);
and U15649 (N_15649,N_15299,N_15399);
or U15650 (N_15650,N_15342,N_15309);
or U15651 (N_15651,N_15465,N_15416);
xor U15652 (N_15652,N_15447,N_15281);
and U15653 (N_15653,N_15331,N_15357);
or U15654 (N_15654,N_15484,N_15430);
nand U15655 (N_15655,N_15489,N_15384);
and U15656 (N_15656,N_15380,N_15312);
or U15657 (N_15657,N_15330,N_15425);
and U15658 (N_15658,N_15406,N_15332);
xnor U15659 (N_15659,N_15469,N_15436);
or U15660 (N_15660,N_15499,N_15455);
or U15661 (N_15661,N_15357,N_15311);
xor U15662 (N_15662,N_15455,N_15408);
or U15663 (N_15663,N_15480,N_15439);
nand U15664 (N_15664,N_15377,N_15440);
nor U15665 (N_15665,N_15289,N_15280);
and U15666 (N_15666,N_15453,N_15491);
nor U15667 (N_15667,N_15490,N_15270);
nor U15668 (N_15668,N_15450,N_15363);
nor U15669 (N_15669,N_15340,N_15470);
or U15670 (N_15670,N_15251,N_15413);
nand U15671 (N_15671,N_15419,N_15329);
nor U15672 (N_15672,N_15374,N_15386);
nand U15673 (N_15673,N_15341,N_15335);
xor U15674 (N_15674,N_15432,N_15362);
nor U15675 (N_15675,N_15388,N_15462);
nor U15676 (N_15676,N_15382,N_15363);
nor U15677 (N_15677,N_15401,N_15490);
or U15678 (N_15678,N_15251,N_15402);
nand U15679 (N_15679,N_15405,N_15472);
xor U15680 (N_15680,N_15276,N_15472);
xor U15681 (N_15681,N_15356,N_15449);
and U15682 (N_15682,N_15419,N_15349);
or U15683 (N_15683,N_15385,N_15334);
or U15684 (N_15684,N_15468,N_15478);
or U15685 (N_15685,N_15330,N_15288);
nor U15686 (N_15686,N_15288,N_15437);
nand U15687 (N_15687,N_15349,N_15433);
nand U15688 (N_15688,N_15308,N_15420);
and U15689 (N_15689,N_15407,N_15420);
xnor U15690 (N_15690,N_15369,N_15324);
and U15691 (N_15691,N_15256,N_15347);
nand U15692 (N_15692,N_15449,N_15487);
and U15693 (N_15693,N_15413,N_15390);
nor U15694 (N_15694,N_15298,N_15353);
nand U15695 (N_15695,N_15404,N_15434);
or U15696 (N_15696,N_15326,N_15361);
nor U15697 (N_15697,N_15494,N_15352);
nand U15698 (N_15698,N_15389,N_15464);
nor U15699 (N_15699,N_15287,N_15383);
nand U15700 (N_15700,N_15253,N_15347);
or U15701 (N_15701,N_15404,N_15472);
and U15702 (N_15702,N_15499,N_15490);
and U15703 (N_15703,N_15282,N_15331);
nor U15704 (N_15704,N_15349,N_15328);
nor U15705 (N_15705,N_15300,N_15428);
and U15706 (N_15706,N_15482,N_15462);
nand U15707 (N_15707,N_15397,N_15419);
and U15708 (N_15708,N_15482,N_15403);
nor U15709 (N_15709,N_15479,N_15363);
or U15710 (N_15710,N_15342,N_15486);
and U15711 (N_15711,N_15300,N_15410);
xor U15712 (N_15712,N_15294,N_15327);
nor U15713 (N_15713,N_15471,N_15289);
and U15714 (N_15714,N_15281,N_15406);
or U15715 (N_15715,N_15471,N_15273);
nand U15716 (N_15716,N_15267,N_15297);
nand U15717 (N_15717,N_15266,N_15315);
and U15718 (N_15718,N_15347,N_15260);
and U15719 (N_15719,N_15331,N_15293);
or U15720 (N_15720,N_15311,N_15355);
nand U15721 (N_15721,N_15480,N_15283);
and U15722 (N_15722,N_15266,N_15412);
nor U15723 (N_15723,N_15460,N_15276);
or U15724 (N_15724,N_15459,N_15311);
nor U15725 (N_15725,N_15293,N_15259);
nand U15726 (N_15726,N_15402,N_15291);
and U15727 (N_15727,N_15398,N_15251);
or U15728 (N_15728,N_15460,N_15493);
and U15729 (N_15729,N_15252,N_15293);
nor U15730 (N_15730,N_15269,N_15454);
nand U15731 (N_15731,N_15488,N_15476);
or U15732 (N_15732,N_15265,N_15291);
xnor U15733 (N_15733,N_15404,N_15454);
nor U15734 (N_15734,N_15255,N_15256);
nor U15735 (N_15735,N_15441,N_15395);
nand U15736 (N_15736,N_15463,N_15320);
and U15737 (N_15737,N_15368,N_15337);
or U15738 (N_15738,N_15299,N_15405);
nor U15739 (N_15739,N_15311,N_15291);
nor U15740 (N_15740,N_15387,N_15320);
nand U15741 (N_15741,N_15458,N_15408);
xor U15742 (N_15742,N_15353,N_15474);
nor U15743 (N_15743,N_15328,N_15369);
and U15744 (N_15744,N_15261,N_15254);
and U15745 (N_15745,N_15435,N_15300);
nand U15746 (N_15746,N_15388,N_15252);
xor U15747 (N_15747,N_15467,N_15276);
or U15748 (N_15748,N_15340,N_15493);
xnor U15749 (N_15749,N_15250,N_15392);
nand U15750 (N_15750,N_15592,N_15604);
or U15751 (N_15751,N_15716,N_15719);
xnor U15752 (N_15752,N_15705,N_15503);
xnor U15753 (N_15753,N_15552,N_15647);
xor U15754 (N_15754,N_15595,N_15550);
and U15755 (N_15755,N_15681,N_15529);
and U15756 (N_15756,N_15528,N_15714);
xor U15757 (N_15757,N_15574,N_15616);
and U15758 (N_15758,N_15640,N_15712);
and U15759 (N_15759,N_15600,N_15689);
nand U15760 (N_15760,N_15549,N_15664);
nand U15761 (N_15761,N_15547,N_15720);
or U15762 (N_15762,N_15546,N_15607);
nor U15763 (N_15763,N_15612,N_15690);
or U15764 (N_15764,N_15725,N_15676);
and U15765 (N_15765,N_15593,N_15562);
or U15766 (N_15766,N_15502,N_15706);
xor U15767 (N_15767,N_15649,N_15695);
and U15768 (N_15768,N_15515,N_15548);
nor U15769 (N_15769,N_15568,N_15519);
and U15770 (N_15770,N_15653,N_15687);
and U15771 (N_15771,N_15585,N_15737);
nor U15772 (N_15772,N_15735,N_15577);
nor U15773 (N_15773,N_15663,N_15511);
nor U15774 (N_15774,N_15718,N_15665);
nor U15775 (N_15775,N_15674,N_15701);
nand U15776 (N_15776,N_15742,N_15527);
xor U15777 (N_15777,N_15621,N_15504);
nand U15778 (N_15778,N_15717,N_15594);
xnor U15779 (N_15779,N_15724,N_15702);
xnor U15780 (N_15780,N_15573,N_15637);
and U15781 (N_15781,N_15516,N_15606);
or U15782 (N_15782,N_15743,N_15601);
nand U15783 (N_15783,N_15740,N_15733);
and U15784 (N_15784,N_15652,N_15668);
or U15785 (N_15785,N_15711,N_15523);
nor U15786 (N_15786,N_15708,N_15700);
xor U15787 (N_15787,N_15579,N_15698);
and U15788 (N_15788,N_15659,N_15669);
nand U15789 (N_15789,N_15541,N_15589);
nor U15790 (N_15790,N_15745,N_15605);
or U15791 (N_15791,N_15513,N_15715);
or U15792 (N_15792,N_15628,N_15746);
and U15793 (N_15793,N_15670,N_15551);
or U15794 (N_15794,N_15707,N_15591);
and U15795 (N_15795,N_15729,N_15648);
nor U15796 (N_15796,N_15538,N_15531);
nand U15797 (N_15797,N_15732,N_15630);
xnor U15798 (N_15798,N_15691,N_15713);
nor U15799 (N_15799,N_15533,N_15641);
and U15800 (N_15800,N_15747,N_15671);
nand U15801 (N_15801,N_15696,N_15726);
or U15802 (N_15802,N_15578,N_15631);
nor U15803 (N_15803,N_15704,N_15650);
xnor U15804 (N_15804,N_15673,N_15553);
and U15805 (N_15805,N_15728,N_15534);
xnor U15806 (N_15806,N_15532,N_15571);
nand U15807 (N_15807,N_15661,N_15561);
or U15808 (N_15808,N_15625,N_15727);
nor U15809 (N_15809,N_15569,N_15634);
nor U15810 (N_15810,N_15629,N_15688);
nand U15811 (N_15811,N_15748,N_15636);
and U15812 (N_15812,N_15610,N_15525);
nor U15813 (N_15813,N_15542,N_15564);
and U15814 (N_15814,N_15555,N_15570);
nand U15815 (N_15815,N_15560,N_15739);
or U15816 (N_15816,N_15638,N_15584);
or U15817 (N_15817,N_15623,N_15559);
xor U15818 (N_15818,N_15590,N_15597);
nand U15819 (N_15819,N_15656,N_15667);
or U15820 (N_15820,N_15512,N_15524);
nand U15821 (N_15821,N_15567,N_15627);
nor U15822 (N_15822,N_15526,N_15693);
or U15823 (N_15823,N_15613,N_15587);
or U15824 (N_15824,N_15723,N_15576);
xor U15825 (N_15825,N_15709,N_15566);
nand U15826 (N_15826,N_15505,N_15518);
and U15827 (N_15827,N_15643,N_15614);
nor U15828 (N_15828,N_15710,N_15507);
xor U15829 (N_15829,N_15514,N_15672);
nand U15830 (N_15830,N_15554,N_15615);
nor U15831 (N_15831,N_15572,N_15588);
or U15832 (N_15832,N_15581,N_15644);
nor U15833 (N_15833,N_15633,N_15683);
or U15834 (N_15834,N_15537,N_15635);
or U15835 (N_15835,N_15522,N_15565);
nor U15836 (N_15836,N_15685,N_15521);
and U15837 (N_15837,N_15655,N_15662);
nor U15838 (N_15838,N_15626,N_15536);
and U15839 (N_15839,N_15611,N_15563);
nand U15840 (N_15840,N_15731,N_15539);
nor U15841 (N_15841,N_15586,N_15684);
xor U15842 (N_15842,N_15558,N_15544);
and U15843 (N_15843,N_15540,N_15582);
nor U15844 (N_15844,N_15624,N_15500);
xor U15845 (N_15845,N_15741,N_15642);
nand U15846 (N_15846,N_15508,N_15680);
nand U15847 (N_15847,N_15666,N_15686);
and U15848 (N_15848,N_15510,N_15599);
xor U15849 (N_15849,N_15694,N_15620);
nor U15850 (N_15850,N_15501,N_15543);
nand U15851 (N_15851,N_15639,N_15509);
and U15852 (N_15852,N_15617,N_15520);
nor U15853 (N_15853,N_15609,N_15598);
xor U15854 (N_15854,N_15646,N_15730);
nand U15855 (N_15855,N_15506,N_15632);
nor U15856 (N_15856,N_15692,N_15618);
nor U15857 (N_15857,N_15580,N_15530);
and U15858 (N_15858,N_15651,N_15545);
nor U15859 (N_15859,N_15557,N_15622);
nor U15860 (N_15860,N_15734,N_15699);
or U15861 (N_15861,N_15749,N_15660);
and U15862 (N_15862,N_15679,N_15517);
or U15863 (N_15863,N_15703,N_15722);
nand U15864 (N_15864,N_15677,N_15608);
or U15865 (N_15865,N_15535,N_15583);
nor U15866 (N_15866,N_15602,N_15556);
nor U15867 (N_15867,N_15697,N_15619);
and U15868 (N_15868,N_15678,N_15738);
or U15869 (N_15869,N_15682,N_15657);
xor U15870 (N_15870,N_15744,N_15575);
or U15871 (N_15871,N_15603,N_15721);
or U15872 (N_15872,N_15658,N_15736);
or U15873 (N_15873,N_15596,N_15645);
nor U15874 (N_15874,N_15654,N_15675);
nor U15875 (N_15875,N_15663,N_15578);
xor U15876 (N_15876,N_15532,N_15666);
or U15877 (N_15877,N_15652,N_15542);
nor U15878 (N_15878,N_15538,N_15696);
nor U15879 (N_15879,N_15567,N_15521);
xor U15880 (N_15880,N_15596,N_15611);
nand U15881 (N_15881,N_15616,N_15696);
or U15882 (N_15882,N_15601,N_15682);
nand U15883 (N_15883,N_15676,N_15565);
nand U15884 (N_15884,N_15664,N_15518);
nor U15885 (N_15885,N_15690,N_15720);
and U15886 (N_15886,N_15617,N_15524);
nand U15887 (N_15887,N_15607,N_15629);
xnor U15888 (N_15888,N_15665,N_15506);
nor U15889 (N_15889,N_15567,N_15612);
xnor U15890 (N_15890,N_15694,N_15637);
or U15891 (N_15891,N_15609,N_15515);
xnor U15892 (N_15892,N_15716,N_15699);
or U15893 (N_15893,N_15625,N_15630);
nand U15894 (N_15894,N_15652,N_15739);
xnor U15895 (N_15895,N_15631,N_15580);
or U15896 (N_15896,N_15617,N_15541);
or U15897 (N_15897,N_15508,N_15556);
and U15898 (N_15898,N_15679,N_15611);
nand U15899 (N_15899,N_15593,N_15697);
xor U15900 (N_15900,N_15721,N_15580);
nor U15901 (N_15901,N_15589,N_15671);
nor U15902 (N_15902,N_15580,N_15704);
and U15903 (N_15903,N_15578,N_15725);
and U15904 (N_15904,N_15554,N_15666);
and U15905 (N_15905,N_15712,N_15561);
nand U15906 (N_15906,N_15737,N_15558);
and U15907 (N_15907,N_15552,N_15561);
xnor U15908 (N_15908,N_15628,N_15668);
nand U15909 (N_15909,N_15749,N_15598);
nor U15910 (N_15910,N_15705,N_15672);
and U15911 (N_15911,N_15505,N_15719);
nand U15912 (N_15912,N_15688,N_15630);
xor U15913 (N_15913,N_15602,N_15667);
nand U15914 (N_15914,N_15632,N_15630);
nand U15915 (N_15915,N_15535,N_15619);
and U15916 (N_15916,N_15729,N_15563);
and U15917 (N_15917,N_15574,N_15701);
nand U15918 (N_15918,N_15679,N_15711);
xor U15919 (N_15919,N_15624,N_15586);
xnor U15920 (N_15920,N_15557,N_15589);
xnor U15921 (N_15921,N_15546,N_15675);
and U15922 (N_15922,N_15596,N_15513);
xor U15923 (N_15923,N_15531,N_15727);
nor U15924 (N_15924,N_15500,N_15669);
or U15925 (N_15925,N_15577,N_15730);
nand U15926 (N_15926,N_15673,N_15519);
nand U15927 (N_15927,N_15586,N_15655);
or U15928 (N_15928,N_15617,N_15706);
xor U15929 (N_15929,N_15522,N_15533);
and U15930 (N_15930,N_15563,N_15646);
nand U15931 (N_15931,N_15739,N_15603);
xor U15932 (N_15932,N_15573,N_15648);
and U15933 (N_15933,N_15598,N_15593);
or U15934 (N_15934,N_15666,N_15508);
nand U15935 (N_15935,N_15742,N_15635);
xor U15936 (N_15936,N_15647,N_15727);
nand U15937 (N_15937,N_15627,N_15561);
nand U15938 (N_15938,N_15722,N_15705);
or U15939 (N_15939,N_15681,N_15637);
and U15940 (N_15940,N_15632,N_15560);
nor U15941 (N_15941,N_15656,N_15582);
nor U15942 (N_15942,N_15624,N_15642);
nor U15943 (N_15943,N_15512,N_15538);
nor U15944 (N_15944,N_15747,N_15639);
or U15945 (N_15945,N_15560,N_15510);
nor U15946 (N_15946,N_15683,N_15553);
nor U15947 (N_15947,N_15505,N_15531);
or U15948 (N_15948,N_15566,N_15648);
xnor U15949 (N_15949,N_15628,N_15612);
nand U15950 (N_15950,N_15562,N_15660);
xnor U15951 (N_15951,N_15734,N_15672);
or U15952 (N_15952,N_15508,N_15724);
nand U15953 (N_15953,N_15725,N_15723);
nor U15954 (N_15954,N_15539,N_15529);
and U15955 (N_15955,N_15596,N_15536);
nor U15956 (N_15956,N_15735,N_15686);
xor U15957 (N_15957,N_15606,N_15577);
xnor U15958 (N_15958,N_15653,N_15611);
nor U15959 (N_15959,N_15705,N_15657);
or U15960 (N_15960,N_15588,N_15546);
nand U15961 (N_15961,N_15548,N_15619);
nand U15962 (N_15962,N_15669,N_15509);
nor U15963 (N_15963,N_15539,N_15692);
xor U15964 (N_15964,N_15536,N_15717);
and U15965 (N_15965,N_15540,N_15720);
nor U15966 (N_15966,N_15591,N_15562);
or U15967 (N_15967,N_15741,N_15617);
nand U15968 (N_15968,N_15573,N_15587);
nand U15969 (N_15969,N_15682,N_15594);
nand U15970 (N_15970,N_15685,N_15583);
xnor U15971 (N_15971,N_15642,N_15589);
and U15972 (N_15972,N_15713,N_15648);
or U15973 (N_15973,N_15610,N_15651);
nand U15974 (N_15974,N_15621,N_15691);
nand U15975 (N_15975,N_15705,N_15637);
nor U15976 (N_15976,N_15592,N_15528);
xor U15977 (N_15977,N_15712,N_15544);
xnor U15978 (N_15978,N_15633,N_15738);
xnor U15979 (N_15979,N_15720,N_15525);
nand U15980 (N_15980,N_15697,N_15626);
or U15981 (N_15981,N_15636,N_15705);
nand U15982 (N_15982,N_15727,N_15522);
nor U15983 (N_15983,N_15641,N_15576);
nor U15984 (N_15984,N_15505,N_15598);
nand U15985 (N_15985,N_15744,N_15723);
or U15986 (N_15986,N_15692,N_15502);
nand U15987 (N_15987,N_15699,N_15648);
or U15988 (N_15988,N_15724,N_15588);
nor U15989 (N_15989,N_15556,N_15743);
nor U15990 (N_15990,N_15664,N_15552);
or U15991 (N_15991,N_15730,N_15503);
nand U15992 (N_15992,N_15621,N_15595);
nand U15993 (N_15993,N_15536,N_15605);
nor U15994 (N_15994,N_15630,N_15574);
nand U15995 (N_15995,N_15550,N_15671);
or U15996 (N_15996,N_15642,N_15590);
and U15997 (N_15997,N_15552,N_15729);
nor U15998 (N_15998,N_15557,N_15720);
xnor U15999 (N_15999,N_15739,N_15627);
and U16000 (N_16000,N_15991,N_15912);
and U16001 (N_16001,N_15973,N_15993);
and U16002 (N_16002,N_15946,N_15805);
nor U16003 (N_16003,N_15871,N_15932);
xor U16004 (N_16004,N_15945,N_15888);
xnor U16005 (N_16005,N_15885,N_15876);
nor U16006 (N_16006,N_15869,N_15947);
or U16007 (N_16007,N_15974,N_15793);
and U16008 (N_16008,N_15894,N_15817);
nor U16009 (N_16009,N_15948,N_15815);
and U16010 (N_16010,N_15768,N_15772);
nor U16011 (N_16011,N_15988,N_15828);
xor U16012 (N_16012,N_15832,N_15907);
xnor U16013 (N_16013,N_15780,N_15863);
or U16014 (N_16014,N_15778,N_15806);
or U16015 (N_16015,N_15783,N_15939);
or U16016 (N_16016,N_15960,N_15970);
nand U16017 (N_16017,N_15972,N_15930);
and U16018 (N_16018,N_15779,N_15767);
nor U16019 (N_16019,N_15899,N_15777);
nor U16020 (N_16020,N_15963,N_15836);
nand U16021 (N_16021,N_15957,N_15875);
nand U16022 (N_16022,N_15873,N_15854);
and U16023 (N_16023,N_15866,N_15881);
or U16024 (N_16024,N_15781,N_15756);
or U16025 (N_16025,N_15975,N_15804);
xor U16026 (N_16026,N_15757,N_15940);
nand U16027 (N_16027,N_15868,N_15814);
or U16028 (N_16028,N_15787,N_15890);
nor U16029 (N_16029,N_15799,N_15902);
nand U16030 (N_16030,N_15891,N_15898);
nor U16031 (N_16031,N_15790,N_15802);
xnor U16032 (N_16032,N_15852,N_15962);
nor U16033 (N_16033,N_15961,N_15998);
xor U16034 (N_16034,N_15809,N_15763);
and U16035 (N_16035,N_15818,N_15771);
xor U16036 (N_16036,N_15897,N_15922);
and U16037 (N_16037,N_15798,N_15859);
or U16038 (N_16038,N_15928,N_15985);
xor U16039 (N_16039,N_15864,N_15941);
nand U16040 (N_16040,N_15831,N_15917);
xor U16041 (N_16041,N_15812,N_15913);
xnor U16042 (N_16042,N_15860,N_15841);
xor U16043 (N_16043,N_15943,N_15813);
nor U16044 (N_16044,N_15807,N_15964);
nand U16045 (N_16045,N_15952,N_15782);
nand U16046 (N_16046,N_15895,N_15884);
nor U16047 (N_16047,N_15829,N_15846);
or U16048 (N_16048,N_15931,N_15791);
or U16049 (N_16049,N_15992,N_15764);
nand U16050 (N_16050,N_15944,N_15942);
xor U16051 (N_16051,N_15933,N_15879);
nor U16052 (N_16052,N_15823,N_15857);
and U16053 (N_16053,N_15851,N_15792);
xnor U16054 (N_16054,N_15853,N_15990);
and U16055 (N_16055,N_15761,N_15750);
nand U16056 (N_16056,N_15955,N_15788);
nor U16057 (N_16057,N_15977,N_15825);
nand U16058 (N_16058,N_15904,N_15819);
xor U16059 (N_16059,N_15784,N_15889);
xor U16060 (N_16060,N_15861,N_15797);
or U16061 (N_16061,N_15751,N_15980);
nand U16062 (N_16062,N_15929,N_15820);
xnor U16063 (N_16063,N_15883,N_15826);
or U16064 (N_16064,N_15915,N_15760);
or U16065 (N_16065,N_15995,N_15949);
or U16066 (N_16066,N_15858,N_15880);
or U16067 (N_16067,N_15810,N_15821);
and U16068 (N_16068,N_15919,N_15834);
nand U16069 (N_16069,N_15752,N_15900);
or U16070 (N_16070,N_15981,N_15914);
and U16071 (N_16071,N_15958,N_15837);
nand U16072 (N_16072,N_15906,N_15785);
nand U16073 (N_16073,N_15924,N_15909);
nor U16074 (N_16074,N_15968,N_15950);
nor U16075 (N_16075,N_15905,N_15822);
xor U16076 (N_16076,N_15966,N_15856);
or U16077 (N_16077,N_15753,N_15997);
and U16078 (N_16078,N_15835,N_15910);
nor U16079 (N_16079,N_15844,N_15775);
xnor U16080 (N_16080,N_15842,N_15976);
nor U16081 (N_16081,N_15867,N_15770);
nand U16082 (N_16082,N_15925,N_15971);
or U16083 (N_16083,N_15811,N_15920);
nor U16084 (N_16084,N_15978,N_15827);
nor U16085 (N_16085,N_15759,N_15923);
or U16086 (N_16086,N_15847,N_15838);
or U16087 (N_16087,N_15903,N_15773);
nor U16088 (N_16088,N_15986,N_15758);
nand U16089 (N_16089,N_15893,N_15965);
nand U16090 (N_16090,N_15855,N_15954);
xnor U16091 (N_16091,N_15896,N_15774);
xnor U16092 (N_16092,N_15795,N_15848);
nor U16093 (N_16093,N_15870,N_15808);
or U16094 (N_16094,N_15916,N_15969);
and U16095 (N_16095,N_15766,N_15927);
or U16096 (N_16096,N_15762,N_15878);
and U16097 (N_16097,N_15769,N_15934);
or U16098 (N_16098,N_15839,N_15938);
nand U16099 (N_16099,N_15953,N_15872);
or U16100 (N_16100,N_15754,N_15840);
xor U16101 (N_16101,N_15996,N_15989);
nand U16102 (N_16102,N_15824,N_15833);
xor U16103 (N_16103,N_15816,N_15882);
nor U16104 (N_16104,N_15935,N_15994);
xor U16105 (N_16105,N_15801,N_15901);
and U16106 (N_16106,N_15967,N_15999);
xnor U16107 (N_16107,N_15830,N_15979);
nand U16108 (N_16108,N_15937,N_15921);
nor U16109 (N_16109,N_15843,N_15845);
nand U16110 (N_16110,N_15796,N_15926);
nor U16111 (N_16111,N_15984,N_15983);
and U16112 (N_16112,N_15982,N_15908);
and U16113 (N_16113,N_15765,N_15959);
or U16114 (N_16114,N_15887,N_15877);
and U16115 (N_16115,N_15800,N_15786);
xnor U16116 (N_16116,N_15865,N_15755);
nand U16117 (N_16117,N_15951,N_15849);
nand U16118 (N_16118,N_15911,N_15850);
nor U16119 (N_16119,N_15918,N_15803);
or U16120 (N_16120,N_15789,N_15794);
or U16121 (N_16121,N_15874,N_15892);
xor U16122 (N_16122,N_15776,N_15886);
or U16123 (N_16123,N_15862,N_15987);
or U16124 (N_16124,N_15956,N_15936);
xnor U16125 (N_16125,N_15911,N_15786);
or U16126 (N_16126,N_15874,N_15909);
and U16127 (N_16127,N_15811,N_15862);
and U16128 (N_16128,N_15998,N_15843);
nor U16129 (N_16129,N_15917,N_15762);
xor U16130 (N_16130,N_15811,N_15885);
and U16131 (N_16131,N_15888,N_15896);
xnor U16132 (N_16132,N_15893,N_15837);
nor U16133 (N_16133,N_15950,N_15751);
and U16134 (N_16134,N_15876,N_15944);
or U16135 (N_16135,N_15824,N_15875);
or U16136 (N_16136,N_15750,N_15876);
nor U16137 (N_16137,N_15848,N_15966);
nor U16138 (N_16138,N_15947,N_15878);
nor U16139 (N_16139,N_15794,N_15803);
or U16140 (N_16140,N_15832,N_15953);
nand U16141 (N_16141,N_15930,N_15909);
nor U16142 (N_16142,N_15793,N_15795);
nor U16143 (N_16143,N_15895,N_15785);
or U16144 (N_16144,N_15780,N_15808);
xor U16145 (N_16145,N_15786,N_15804);
and U16146 (N_16146,N_15837,N_15956);
and U16147 (N_16147,N_15894,N_15821);
nor U16148 (N_16148,N_15755,N_15934);
nor U16149 (N_16149,N_15801,N_15913);
nor U16150 (N_16150,N_15811,N_15799);
or U16151 (N_16151,N_15852,N_15988);
nor U16152 (N_16152,N_15851,N_15917);
xor U16153 (N_16153,N_15763,N_15790);
nand U16154 (N_16154,N_15817,N_15841);
xor U16155 (N_16155,N_15978,N_15775);
xnor U16156 (N_16156,N_15970,N_15898);
and U16157 (N_16157,N_15936,N_15831);
xor U16158 (N_16158,N_15793,N_15850);
xor U16159 (N_16159,N_15786,N_15958);
nor U16160 (N_16160,N_15826,N_15834);
and U16161 (N_16161,N_15842,N_15820);
and U16162 (N_16162,N_15777,N_15833);
and U16163 (N_16163,N_15759,N_15798);
and U16164 (N_16164,N_15839,N_15894);
and U16165 (N_16165,N_15879,N_15951);
and U16166 (N_16166,N_15858,N_15932);
and U16167 (N_16167,N_15951,N_15913);
xor U16168 (N_16168,N_15917,N_15807);
nor U16169 (N_16169,N_15793,N_15913);
or U16170 (N_16170,N_15808,N_15896);
nor U16171 (N_16171,N_15831,N_15973);
or U16172 (N_16172,N_15902,N_15988);
nand U16173 (N_16173,N_15778,N_15834);
or U16174 (N_16174,N_15994,N_15972);
xor U16175 (N_16175,N_15822,N_15969);
and U16176 (N_16176,N_15768,N_15961);
xnor U16177 (N_16177,N_15871,N_15906);
nand U16178 (N_16178,N_15842,N_15973);
xor U16179 (N_16179,N_15850,N_15950);
nand U16180 (N_16180,N_15980,N_15892);
nor U16181 (N_16181,N_15803,N_15806);
xnor U16182 (N_16182,N_15764,N_15809);
and U16183 (N_16183,N_15812,N_15925);
xnor U16184 (N_16184,N_15854,N_15857);
nor U16185 (N_16185,N_15822,N_15882);
xnor U16186 (N_16186,N_15893,N_15854);
nor U16187 (N_16187,N_15826,N_15914);
nand U16188 (N_16188,N_15864,N_15877);
nand U16189 (N_16189,N_15761,N_15976);
and U16190 (N_16190,N_15887,N_15807);
and U16191 (N_16191,N_15881,N_15955);
xor U16192 (N_16192,N_15904,N_15783);
nor U16193 (N_16193,N_15924,N_15902);
nand U16194 (N_16194,N_15753,N_15854);
xor U16195 (N_16195,N_15996,N_15942);
nand U16196 (N_16196,N_15872,N_15818);
nand U16197 (N_16197,N_15785,N_15958);
nor U16198 (N_16198,N_15869,N_15835);
nand U16199 (N_16199,N_15867,N_15938);
xor U16200 (N_16200,N_15966,N_15905);
or U16201 (N_16201,N_15862,N_15916);
nor U16202 (N_16202,N_15991,N_15866);
and U16203 (N_16203,N_15951,N_15941);
and U16204 (N_16204,N_15852,N_15754);
and U16205 (N_16205,N_15833,N_15911);
or U16206 (N_16206,N_15946,N_15816);
nor U16207 (N_16207,N_15784,N_15903);
nor U16208 (N_16208,N_15965,N_15848);
xor U16209 (N_16209,N_15855,N_15760);
or U16210 (N_16210,N_15803,N_15943);
xnor U16211 (N_16211,N_15993,N_15980);
nor U16212 (N_16212,N_15798,N_15918);
and U16213 (N_16213,N_15894,N_15955);
nor U16214 (N_16214,N_15808,N_15917);
or U16215 (N_16215,N_15792,N_15966);
nor U16216 (N_16216,N_15852,N_15922);
or U16217 (N_16217,N_15966,N_15967);
nand U16218 (N_16218,N_15860,N_15980);
nor U16219 (N_16219,N_15870,N_15989);
or U16220 (N_16220,N_15804,N_15768);
or U16221 (N_16221,N_15993,N_15768);
nand U16222 (N_16222,N_15750,N_15994);
nand U16223 (N_16223,N_15804,N_15883);
and U16224 (N_16224,N_15993,N_15856);
xor U16225 (N_16225,N_15907,N_15947);
nand U16226 (N_16226,N_15952,N_15898);
nor U16227 (N_16227,N_15784,N_15980);
and U16228 (N_16228,N_15808,N_15914);
and U16229 (N_16229,N_15774,N_15828);
and U16230 (N_16230,N_15812,N_15873);
xnor U16231 (N_16231,N_15887,N_15865);
nor U16232 (N_16232,N_15811,N_15905);
and U16233 (N_16233,N_15965,N_15903);
and U16234 (N_16234,N_15848,N_15801);
xnor U16235 (N_16235,N_15879,N_15999);
and U16236 (N_16236,N_15936,N_15920);
and U16237 (N_16237,N_15908,N_15980);
xor U16238 (N_16238,N_15788,N_15808);
nand U16239 (N_16239,N_15883,N_15996);
xor U16240 (N_16240,N_15918,N_15977);
nand U16241 (N_16241,N_15851,N_15866);
nor U16242 (N_16242,N_15895,N_15847);
and U16243 (N_16243,N_15831,N_15929);
or U16244 (N_16244,N_15917,N_15836);
nor U16245 (N_16245,N_15807,N_15794);
nand U16246 (N_16246,N_15916,N_15818);
and U16247 (N_16247,N_15968,N_15907);
and U16248 (N_16248,N_15848,N_15877);
nand U16249 (N_16249,N_15882,N_15852);
nand U16250 (N_16250,N_16054,N_16083);
or U16251 (N_16251,N_16173,N_16104);
or U16252 (N_16252,N_16235,N_16228);
nand U16253 (N_16253,N_16074,N_16163);
xor U16254 (N_16254,N_16095,N_16194);
xnor U16255 (N_16255,N_16025,N_16124);
and U16256 (N_16256,N_16105,N_16185);
nand U16257 (N_16257,N_16200,N_16210);
nand U16258 (N_16258,N_16189,N_16192);
nor U16259 (N_16259,N_16154,N_16061);
nor U16260 (N_16260,N_16220,N_16208);
xnor U16261 (N_16261,N_16132,N_16015);
nor U16262 (N_16262,N_16140,N_16197);
nor U16263 (N_16263,N_16069,N_16227);
nor U16264 (N_16264,N_16018,N_16065);
xor U16265 (N_16265,N_16056,N_16085);
xnor U16266 (N_16266,N_16195,N_16026);
xor U16267 (N_16267,N_16012,N_16206);
xnor U16268 (N_16268,N_16032,N_16191);
and U16269 (N_16269,N_16033,N_16135);
nand U16270 (N_16270,N_16111,N_16023);
and U16271 (N_16271,N_16039,N_16179);
nor U16272 (N_16272,N_16204,N_16183);
and U16273 (N_16273,N_16157,N_16169);
nand U16274 (N_16274,N_16221,N_16171);
nand U16275 (N_16275,N_16158,N_16244);
xor U16276 (N_16276,N_16168,N_16215);
nand U16277 (N_16277,N_16145,N_16131);
nand U16278 (N_16278,N_16050,N_16003);
and U16279 (N_16279,N_16116,N_16029);
and U16280 (N_16280,N_16062,N_16136);
xnor U16281 (N_16281,N_16068,N_16151);
nand U16282 (N_16282,N_16028,N_16106);
nor U16283 (N_16283,N_16038,N_16059);
xnor U16284 (N_16284,N_16188,N_16232);
and U16285 (N_16285,N_16128,N_16034);
and U16286 (N_16286,N_16207,N_16109);
nor U16287 (N_16287,N_16222,N_16230);
and U16288 (N_16288,N_16091,N_16149);
and U16289 (N_16289,N_16092,N_16156);
nor U16290 (N_16290,N_16182,N_16066);
nand U16291 (N_16291,N_16180,N_16042);
xnor U16292 (N_16292,N_16159,N_16184);
xnor U16293 (N_16293,N_16239,N_16078);
xnor U16294 (N_16294,N_16088,N_16129);
or U16295 (N_16295,N_16112,N_16102);
nand U16296 (N_16296,N_16031,N_16130);
xor U16297 (N_16297,N_16080,N_16119);
and U16298 (N_16298,N_16087,N_16127);
xnor U16299 (N_16299,N_16234,N_16202);
nand U16300 (N_16300,N_16160,N_16090);
and U16301 (N_16301,N_16107,N_16123);
and U16302 (N_16302,N_16043,N_16082);
or U16303 (N_16303,N_16233,N_16084);
xnor U16304 (N_16304,N_16108,N_16120);
or U16305 (N_16305,N_16040,N_16203);
or U16306 (N_16306,N_16075,N_16133);
and U16307 (N_16307,N_16216,N_16242);
and U16308 (N_16308,N_16167,N_16096);
and U16309 (N_16309,N_16086,N_16057);
xor U16310 (N_16310,N_16113,N_16079);
and U16311 (N_16311,N_16243,N_16010);
and U16312 (N_16312,N_16170,N_16049);
nand U16313 (N_16313,N_16046,N_16247);
xnor U16314 (N_16314,N_16001,N_16166);
or U16315 (N_16315,N_16245,N_16209);
nand U16316 (N_16316,N_16030,N_16110);
or U16317 (N_16317,N_16076,N_16052);
nand U16318 (N_16318,N_16053,N_16051);
and U16319 (N_16319,N_16213,N_16024);
or U16320 (N_16320,N_16081,N_16060);
xor U16321 (N_16321,N_16117,N_16186);
or U16322 (N_16322,N_16205,N_16201);
and U16323 (N_16323,N_16240,N_16000);
nor U16324 (N_16324,N_16008,N_16193);
xor U16325 (N_16325,N_16199,N_16198);
or U16326 (N_16326,N_16225,N_16218);
xor U16327 (N_16327,N_16045,N_16021);
xnor U16328 (N_16328,N_16067,N_16236);
nand U16329 (N_16329,N_16217,N_16002);
nor U16330 (N_16330,N_16044,N_16125);
or U16331 (N_16331,N_16098,N_16126);
or U16332 (N_16332,N_16141,N_16137);
and U16333 (N_16333,N_16237,N_16099);
and U16334 (N_16334,N_16150,N_16100);
nor U16335 (N_16335,N_16037,N_16161);
or U16336 (N_16336,N_16249,N_16147);
nand U16337 (N_16337,N_16071,N_16115);
or U16338 (N_16338,N_16196,N_16174);
xor U16339 (N_16339,N_16172,N_16229);
and U16340 (N_16340,N_16016,N_16006);
or U16341 (N_16341,N_16155,N_16089);
nand U16342 (N_16342,N_16020,N_16055);
or U16343 (N_16343,N_16072,N_16231);
xnor U16344 (N_16344,N_16211,N_16004);
nand U16345 (N_16345,N_16223,N_16142);
or U16346 (N_16346,N_16238,N_16073);
or U16347 (N_16347,N_16162,N_16118);
nand U16348 (N_16348,N_16047,N_16121);
nor U16349 (N_16349,N_16063,N_16022);
nor U16350 (N_16350,N_16094,N_16219);
nor U16351 (N_16351,N_16048,N_16093);
and U16352 (N_16352,N_16019,N_16097);
nor U16353 (N_16353,N_16187,N_16009);
xnor U16354 (N_16354,N_16214,N_16103);
and U16355 (N_16355,N_16041,N_16241);
and U16356 (N_16356,N_16134,N_16146);
nor U16357 (N_16357,N_16143,N_16139);
or U16358 (N_16358,N_16144,N_16005);
nor U16359 (N_16359,N_16152,N_16148);
xnor U16360 (N_16360,N_16176,N_16122);
and U16361 (N_16361,N_16246,N_16070);
nand U16362 (N_16362,N_16153,N_16011);
and U16363 (N_16363,N_16077,N_16064);
or U16364 (N_16364,N_16017,N_16013);
nor U16365 (N_16365,N_16178,N_16164);
nand U16366 (N_16366,N_16175,N_16248);
nand U16367 (N_16367,N_16138,N_16058);
or U16368 (N_16368,N_16114,N_16036);
nand U16369 (N_16369,N_16190,N_16027);
xnor U16370 (N_16370,N_16224,N_16014);
nand U16371 (N_16371,N_16007,N_16212);
and U16372 (N_16372,N_16035,N_16101);
and U16373 (N_16373,N_16181,N_16177);
xor U16374 (N_16374,N_16226,N_16165);
nand U16375 (N_16375,N_16145,N_16048);
or U16376 (N_16376,N_16136,N_16029);
and U16377 (N_16377,N_16236,N_16191);
xor U16378 (N_16378,N_16195,N_16222);
xor U16379 (N_16379,N_16192,N_16060);
nor U16380 (N_16380,N_16040,N_16174);
xnor U16381 (N_16381,N_16201,N_16003);
xnor U16382 (N_16382,N_16014,N_16148);
nand U16383 (N_16383,N_16027,N_16117);
or U16384 (N_16384,N_16135,N_16058);
nor U16385 (N_16385,N_16022,N_16242);
and U16386 (N_16386,N_16008,N_16107);
xnor U16387 (N_16387,N_16209,N_16032);
and U16388 (N_16388,N_16219,N_16081);
nor U16389 (N_16389,N_16150,N_16229);
xor U16390 (N_16390,N_16089,N_16243);
nor U16391 (N_16391,N_16234,N_16167);
nor U16392 (N_16392,N_16139,N_16036);
nand U16393 (N_16393,N_16198,N_16109);
and U16394 (N_16394,N_16188,N_16019);
or U16395 (N_16395,N_16232,N_16109);
or U16396 (N_16396,N_16013,N_16079);
and U16397 (N_16397,N_16084,N_16241);
or U16398 (N_16398,N_16137,N_16123);
and U16399 (N_16399,N_16008,N_16017);
nand U16400 (N_16400,N_16235,N_16129);
nor U16401 (N_16401,N_16100,N_16022);
nand U16402 (N_16402,N_16249,N_16012);
nand U16403 (N_16403,N_16174,N_16055);
nor U16404 (N_16404,N_16139,N_16131);
xor U16405 (N_16405,N_16145,N_16202);
or U16406 (N_16406,N_16154,N_16226);
nand U16407 (N_16407,N_16041,N_16159);
nor U16408 (N_16408,N_16015,N_16095);
nand U16409 (N_16409,N_16135,N_16193);
xor U16410 (N_16410,N_16164,N_16127);
and U16411 (N_16411,N_16162,N_16101);
or U16412 (N_16412,N_16241,N_16158);
or U16413 (N_16413,N_16108,N_16077);
nor U16414 (N_16414,N_16067,N_16220);
xor U16415 (N_16415,N_16150,N_16120);
or U16416 (N_16416,N_16080,N_16212);
or U16417 (N_16417,N_16036,N_16051);
or U16418 (N_16418,N_16048,N_16157);
and U16419 (N_16419,N_16065,N_16119);
or U16420 (N_16420,N_16057,N_16230);
and U16421 (N_16421,N_16226,N_16186);
nor U16422 (N_16422,N_16092,N_16114);
nor U16423 (N_16423,N_16235,N_16053);
or U16424 (N_16424,N_16081,N_16228);
xor U16425 (N_16425,N_16131,N_16128);
and U16426 (N_16426,N_16126,N_16237);
or U16427 (N_16427,N_16233,N_16196);
xor U16428 (N_16428,N_16026,N_16037);
and U16429 (N_16429,N_16172,N_16095);
or U16430 (N_16430,N_16011,N_16027);
and U16431 (N_16431,N_16116,N_16122);
and U16432 (N_16432,N_16064,N_16199);
nor U16433 (N_16433,N_16165,N_16114);
or U16434 (N_16434,N_16182,N_16114);
nor U16435 (N_16435,N_16003,N_16131);
nor U16436 (N_16436,N_16044,N_16000);
xor U16437 (N_16437,N_16165,N_16221);
and U16438 (N_16438,N_16061,N_16232);
and U16439 (N_16439,N_16192,N_16153);
or U16440 (N_16440,N_16115,N_16092);
xnor U16441 (N_16441,N_16202,N_16043);
nor U16442 (N_16442,N_16249,N_16120);
nor U16443 (N_16443,N_16222,N_16070);
or U16444 (N_16444,N_16117,N_16041);
or U16445 (N_16445,N_16120,N_16105);
and U16446 (N_16446,N_16094,N_16153);
and U16447 (N_16447,N_16032,N_16229);
xnor U16448 (N_16448,N_16105,N_16219);
and U16449 (N_16449,N_16178,N_16053);
nand U16450 (N_16450,N_16141,N_16220);
nor U16451 (N_16451,N_16083,N_16003);
or U16452 (N_16452,N_16194,N_16073);
or U16453 (N_16453,N_16164,N_16100);
or U16454 (N_16454,N_16053,N_16000);
nor U16455 (N_16455,N_16127,N_16050);
or U16456 (N_16456,N_16158,N_16061);
xor U16457 (N_16457,N_16048,N_16212);
nor U16458 (N_16458,N_16216,N_16107);
nor U16459 (N_16459,N_16065,N_16078);
xnor U16460 (N_16460,N_16149,N_16087);
nand U16461 (N_16461,N_16242,N_16217);
and U16462 (N_16462,N_16183,N_16167);
or U16463 (N_16463,N_16037,N_16223);
xor U16464 (N_16464,N_16187,N_16221);
xor U16465 (N_16465,N_16045,N_16046);
or U16466 (N_16466,N_16246,N_16185);
and U16467 (N_16467,N_16156,N_16076);
nor U16468 (N_16468,N_16127,N_16124);
xnor U16469 (N_16469,N_16201,N_16125);
and U16470 (N_16470,N_16184,N_16025);
nor U16471 (N_16471,N_16219,N_16210);
nor U16472 (N_16472,N_16248,N_16068);
and U16473 (N_16473,N_16160,N_16003);
nand U16474 (N_16474,N_16119,N_16016);
and U16475 (N_16475,N_16203,N_16189);
or U16476 (N_16476,N_16001,N_16144);
xor U16477 (N_16477,N_16157,N_16032);
nand U16478 (N_16478,N_16157,N_16156);
and U16479 (N_16479,N_16189,N_16029);
and U16480 (N_16480,N_16013,N_16011);
and U16481 (N_16481,N_16008,N_16043);
and U16482 (N_16482,N_16153,N_16146);
nor U16483 (N_16483,N_16054,N_16174);
xnor U16484 (N_16484,N_16006,N_16221);
xor U16485 (N_16485,N_16174,N_16100);
or U16486 (N_16486,N_16150,N_16073);
and U16487 (N_16487,N_16031,N_16171);
xnor U16488 (N_16488,N_16053,N_16183);
nand U16489 (N_16489,N_16221,N_16155);
nor U16490 (N_16490,N_16233,N_16027);
or U16491 (N_16491,N_16090,N_16135);
nand U16492 (N_16492,N_16192,N_16131);
and U16493 (N_16493,N_16212,N_16248);
or U16494 (N_16494,N_16101,N_16161);
nor U16495 (N_16495,N_16150,N_16055);
or U16496 (N_16496,N_16035,N_16056);
or U16497 (N_16497,N_16136,N_16227);
or U16498 (N_16498,N_16024,N_16096);
xor U16499 (N_16499,N_16005,N_16203);
nand U16500 (N_16500,N_16429,N_16493);
nand U16501 (N_16501,N_16387,N_16448);
and U16502 (N_16502,N_16406,N_16295);
and U16503 (N_16503,N_16446,N_16273);
or U16504 (N_16504,N_16361,N_16411);
xnor U16505 (N_16505,N_16302,N_16359);
and U16506 (N_16506,N_16324,N_16407);
nor U16507 (N_16507,N_16274,N_16421);
or U16508 (N_16508,N_16316,N_16272);
or U16509 (N_16509,N_16357,N_16384);
nor U16510 (N_16510,N_16415,N_16325);
or U16511 (N_16511,N_16263,N_16354);
and U16512 (N_16512,N_16313,N_16306);
and U16513 (N_16513,N_16380,N_16327);
nand U16514 (N_16514,N_16457,N_16307);
nand U16515 (N_16515,N_16365,N_16386);
xnor U16516 (N_16516,N_16443,N_16401);
nor U16517 (N_16517,N_16485,N_16499);
xnor U16518 (N_16518,N_16342,N_16343);
or U16519 (N_16519,N_16285,N_16293);
and U16520 (N_16520,N_16439,N_16334);
or U16521 (N_16521,N_16312,N_16492);
xor U16522 (N_16522,N_16400,N_16351);
nand U16523 (N_16523,N_16290,N_16482);
or U16524 (N_16524,N_16367,N_16321);
and U16525 (N_16525,N_16438,N_16283);
nand U16526 (N_16526,N_16434,N_16275);
nand U16527 (N_16527,N_16371,N_16314);
and U16528 (N_16528,N_16425,N_16322);
and U16529 (N_16529,N_16483,N_16481);
and U16530 (N_16530,N_16479,N_16254);
nor U16531 (N_16531,N_16397,N_16336);
nand U16532 (N_16532,N_16301,N_16494);
nand U16533 (N_16533,N_16497,N_16463);
nor U16534 (N_16534,N_16284,N_16427);
xor U16535 (N_16535,N_16491,N_16424);
nor U16536 (N_16536,N_16432,N_16416);
nand U16537 (N_16537,N_16253,N_16330);
or U16538 (N_16538,N_16375,N_16468);
nand U16539 (N_16539,N_16474,N_16445);
xor U16540 (N_16540,N_16399,N_16475);
or U16541 (N_16541,N_16454,N_16394);
nand U16542 (N_16542,N_16477,N_16345);
or U16543 (N_16543,N_16320,N_16369);
nand U16544 (N_16544,N_16298,N_16389);
and U16545 (N_16545,N_16435,N_16402);
xor U16546 (N_16546,N_16323,N_16413);
nor U16547 (N_16547,N_16417,N_16318);
and U16548 (N_16548,N_16469,N_16376);
nor U16549 (N_16549,N_16256,N_16431);
xnor U16550 (N_16550,N_16259,N_16348);
nor U16551 (N_16551,N_16419,N_16317);
or U16552 (N_16552,N_16490,N_16266);
and U16553 (N_16553,N_16442,N_16255);
nor U16554 (N_16554,N_16264,N_16453);
nand U16555 (N_16555,N_16370,N_16449);
or U16556 (N_16556,N_16260,N_16422);
and U16557 (N_16557,N_16391,N_16309);
nand U16558 (N_16558,N_16360,N_16430);
or U16559 (N_16559,N_16478,N_16456);
nor U16560 (N_16560,N_16498,N_16332);
nor U16561 (N_16561,N_16296,N_16339);
and U16562 (N_16562,N_16465,N_16441);
nand U16563 (N_16563,N_16395,N_16372);
nand U16564 (N_16564,N_16258,N_16269);
xnor U16565 (N_16565,N_16329,N_16414);
or U16566 (N_16566,N_16251,N_16282);
xnor U16567 (N_16567,N_16458,N_16262);
or U16568 (N_16568,N_16250,N_16393);
nor U16569 (N_16569,N_16385,N_16356);
or U16570 (N_16570,N_16310,N_16381);
and U16571 (N_16571,N_16358,N_16473);
xor U16572 (N_16572,N_16488,N_16418);
and U16573 (N_16573,N_16455,N_16464);
xor U16574 (N_16574,N_16412,N_16279);
nor U16575 (N_16575,N_16467,N_16319);
xnor U16576 (N_16576,N_16362,N_16462);
or U16577 (N_16577,N_16363,N_16396);
nor U16578 (N_16578,N_16436,N_16460);
or U16579 (N_16579,N_16305,N_16486);
nand U16580 (N_16580,N_16252,N_16461);
nor U16581 (N_16581,N_16423,N_16480);
and U16582 (N_16582,N_16466,N_16338);
or U16583 (N_16583,N_16374,N_16489);
or U16584 (N_16584,N_16335,N_16409);
nor U16585 (N_16585,N_16308,N_16286);
nand U16586 (N_16586,N_16487,N_16315);
nor U16587 (N_16587,N_16333,N_16257);
nand U16588 (N_16588,N_16300,N_16398);
or U16589 (N_16589,N_16472,N_16404);
or U16590 (N_16590,N_16261,N_16366);
and U16591 (N_16591,N_16297,N_16270);
and U16592 (N_16592,N_16368,N_16470);
nor U16593 (N_16593,N_16484,N_16288);
nor U16594 (N_16594,N_16344,N_16340);
and U16595 (N_16595,N_16265,N_16352);
nor U16596 (N_16596,N_16382,N_16495);
or U16597 (N_16597,N_16311,N_16268);
nand U16598 (N_16598,N_16331,N_16353);
xnor U16599 (N_16599,N_16388,N_16291);
nand U16600 (N_16600,N_16303,N_16428);
nand U16601 (N_16601,N_16355,N_16346);
nor U16602 (N_16602,N_16377,N_16405);
or U16603 (N_16603,N_16292,N_16277);
or U16604 (N_16604,N_16390,N_16337);
nand U16605 (N_16605,N_16450,N_16281);
or U16606 (N_16606,N_16276,N_16341);
and U16607 (N_16607,N_16392,N_16471);
xnor U16608 (N_16608,N_16403,N_16459);
or U16609 (N_16609,N_16289,N_16299);
and U16610 (N_16610,N_16433,N_16383);
nand U16611 (N_16611,N_16294,N_16326);
nor U16612 (N_16612,N_16287,N_16378);
and U16613 (N_16613,N_16476,N_16349);
and U16614 (N_16614,N_16280,N_16447);
nor U16615 (N_16615,N_16420,N_16452);
xor U16616 (N_16616,N_16364,N_16426);
or U16617 (N_16617,N_16451,N_16408);
and U16618 (N_16618,N_16271,N_16437);
nor U16619 (N_16619,N_16444,N_16278);
xor U16620 (N_16620,N_16350,N_16410);
and U16621 (N_16621,N_16328,N_16379);
nor U16622 (N_16622,N_16304,N_16267);
or U16623 (N_16623,N_16496,N_16373);
nor U16624 (N_16624,N_16347,N_16440);
nor U16625 (N_16625,N_16318,N_16307);
xor U16626 (N_16626,N_16300,N_16306);
nand U16627 (N_16627,N_16494,N_16348);
and U16628 (N_16628,N_16432,N_16268);
and U16629 (N_16629,N_16456,N_16380);
and U16630 (N_16630,N_16471,N_16389);
nor U16631 (N_16631,N_16336,N_16300);
nor U16632 (N_16632,N_16278,N_16291);
xor U16633 (N_16633,N_16378,N_16268);
nand U16634 (N_16634,N_16255,N_16258);
and U16635 (N_16635,N_16271,N_16384);
and U16636 (N_16636,N_16443,N_16447);
nand U16637 (N_16637,N_16490,N_16485);
nand U16638 (N_16638,N_16297,N_16328);
xor U16639 (N_16639,N_16267,N_16456);
and U16640 (N_16640,N_16391,N_16371);
xor U16641 (N_16641,N_16256,N_16438);
and U16642 (N_16642,N_16441,N_16314);
and U16643 (N_16643,N_16262,N_16321);
xor U16644 (N_16644,N_16440,N_16289);
nand U16645 (N_16645,N_16322,N_16437);
xor U16646 (N_16646,N_16390,N_16310);
nand U16647 (N_16647,N_16417,N_16351);
and U16648 (N_16648,N_16320,N_16304);
and U16649 (N_16649,N_16389,N_16392);
and U16650 (N_16650,N_16353,N_16295);
xnor U16651 (N_16651,N_16357,N_16316);
nor U16652 (N_16652,N_16463,N_16416);
or U16653 (N_16653,N_16296,N_16491);
or U16654 (N_16654,N_16477,N_16336);
xnor U16655 (N_16655,N_16301,N_16347);
xnor U16656 (N_16656,N_16397,N_16317);
or U16657 (N_16657,N_16468,N_16252);
nand U16658 (N_16658,N_16265,N_16261);
nand U16659 (N_16659,N_16387,N_16383);
nor U16660 (N_16660,N_16387,N_16266);
xnor U16661 (N_16661,N_16264,N_16365);
xor U16662 (N_16662,N_16393,N_16383);
or U16663 (N_16663,N_16287,N_16499);
xor U16664 (N_16664,N_16476,N_16400);
and U16665 (N_16665,N_16452,N_16480);
nand U16666 (N_16666,N_16334,N_16368);
and U16667 (N_16667,N_16440,N_16498);
or U16668 (N_16668,N_16283,N_16412);
xor U16669 (N_16669,N_16460,N_16499);
xor U16670 (N_16670,N_16257,N_16336);
nor U16671 (N_16671,N_16371,N_16479);
and U16672 (N_16672,N_16291,N_16467);
xnor U16673 (N_16673,N_16424,N_16496);
xor U16674 (N_16674,N_16464,N_16319);
and U16675 (N_16675,N_16455,N_16271);
nor U16676 (N_16676,N_16250,N_16470);
and U16677 (N_16677,N_16455,N_16398);
or U16678 (N_16678,N_16494,N_16255);
or U16679 (N_16679,N_16449,N_16445);
xor U16680 (N_16680,N_16401,N_16307);
or U16681 (N_16681,N_16413,N_16382);
or U16682 (N_16682,N_16486,N_16366);
nand U16683 (N_16683,N_16415,N_16483);
nor U16684 (N_16684,N_16446,N_16296);
nor U16685 (N_16685,N_16255,N_16322);
nand U16686 (N_16686,N_16286,N_16366);
or U16687 (N_16687,N_16255,N_16486);
nand U16688 (N_16688,N_16414,N_16302);
or U16689 (N_16689,N_16313,N_16255);
xor U16690 (N_16690,N_16479,N_16352);
nand U16691 (N_16691,N_16377,N_16412);
and U16692 (N_16692,N_16266,N_16261);
xnor U16693 (N_16693,N_16348,N_16474);
or U16694 (N_16694,N_16319,N_16305);
or U16695 (N_16695,N_16333,N_16403);
or U16696 (N_16696,N_16385,N_16285);
nor U16697 (N_16697,N_16465,N_16445);
and U16698 (N_16698,N_16326,N_16403);
nand U16699 (N_16699,N_16337,N_16419);
nor U16700 (N_16700,N_16338,N_16461);
or U16701 (N_16701,N_16491,N_16490);
nor U16702 (N_16702,N_16315,N_16326);
and U16703 (N_16703,N_16373,N_16259);
and U16704 (N_16704,N_16346,N_16261);
nand U16705 (N_16705,N_16295,N_16327);
nand U16706 (N_16706,N_16447,N_16309);
xor U16707 (N_16707,N_16339,N_16270);
or U16708 (N_16708,N_16295,N_16405);
nor U16709 (N_16709,N_16266,N_16384);
and U16710 (N_16710,N_16267,N_16262);
or U16711 (N_16711,N_16339,N_16461);
or U16712 (N_16712,N_16432,N_16483);
nand U16713 (N_16713,N_16473,N_16418);
nor U16714 (N_16714,N_16414,N_16458);
nand U16715 (N_16715,N_16459,N_16381);
or U16716 (N_16716,N_16272,N_16315);
or U16717 (N_16717,N_16421,N_16395);
and U16718 (N_16718,N_16333,N_16411);
xnor U16719 (N_16719,N_16264,N_16417);
or U16720 (N_16720,N_16276,N_16259);
and U16721 (N_16721,N_16449,N_16422);
and U16722 (N_16722,N_16328,N_16295);
nor U16723 (N_16723,N_16289,N_16252);
nor U16724 (N_16724,N_16412,N_16429);
and U16725 (N_16725,N_16293,N_16358);
xnor U16726 (N_16726,N_16379,N_16357);
and U16727 (N_16727,N_16285,N_16297);
nor U16728 (N_16728,N_16388,N_16486);
nor U16729 (N_16729,N_16377,N_16421);
and U16730 (N_16730,N_16460,N_16328);
xor U16731 (N_16731,N_16336,N_16496);
nand U16732 (N_16732,N_16473,N_16291);
or U16733 (N_16733,N_16431,N_16409);
and U16734 (N_16734,N_16283,N_16331);
nor U16735 (N_16735,N_16453,N_16306);
nand U16736 (N_16736,N_16297,N_16423);
and U16737 (N_16737,N_16461,N_16317);
nor U16738 (N_16738,N_16287,N_16324);
and U16739 (N_16739,N_16301,N_16478);
nand U16740 (N_16740,N_16340,N_16311);
nor U16741 (N_16741,N_16319,N_16332);
nand U16742 (N_16742,N_16463,N_16298);
xor U16743 (N_16743,N_16438,N_16304);
or U16744 (N_16744,N_16387,N_16490);
nand U16745 (N_16745,N_16457,N_16256);
xor U16746 (N_16746,N_16270,N_16464);
nand U16747 (N_16747,N_16338,N_16253);
and U16748 (N_16748,N_16340,N_16269);
xnor U16749 (N_16749,N_16384,N_16432);
xor U16750 (N_16750,N_16700,N_16747);
nor U16751 (N_16751,N_16578,N_16689);
xnor U16752 (N_16752,N_16584,N_16685);
and U16753 (N_16753,N_16543,N_16749);
nor U16754 (N_16754,N_16613,N_16646);
xor U16755 (N_16755,N_16673,N_16528);
nand U16756 (N_16756,N_16538,N_16540);
or U16757 (N_16757,N_16710,N_16644);
or U16758 (N_16758,N_16722,N_16683);
xor U16759 (N_16759,N_16593,N_16654);
xnor U16760 (N_16760,N_16585,N_16723);
nand U16761 (N_16761,N_16653,N_16628);
or U16762 (N_16762,N_16731,N_16676);
and U16763 (N_16763,N_16535,N_16674);
and U16764 (N_16764,N_16506,N_16642);
and U16765 (N_16765,N_16717,N_16640);
xnor U16766 (N_16766,N_16504,N_16730);
or U16767 (N_16767,N_16698,N_16550);
or U16768 (N_16768,N_16576,N_16627);
or U16769 (N_16769,N_16630,N_16726);
xnor U16770 (N_16770,N_16574,N_16580);
and U16771 (N_16771,N_16546,N_16520);
xnor U16772 (N_16772,N_16526,N_16609);
nor U16773 (N_16773,N_16664,N_16519);
nor U16774 (N_16774,N_16541,N_16510);
and U16775 (N_16775,N_16706,N_16547);
or U16776 (N_16776,N_16732,N_16744);
nor U16777 (N_16777,N_16632,N_16745);
or U16778 (N_16778,N_16662,N_16645);
nor U16779 (N_16779,N_16599,N_16678);
or U16780 (N_16780,N_16572,N_16603);
and U16781 (N_16781,N_16587,N_16512);
nand U16782 (N_16782,N_16513,N_16622);
nand U16783 (N_16783,N_16514,N_16637);
xor U16784 (N_16784,N_16690,N_16701);
and U16785 (N_16785,N_16534,N_16610);
xnor U16786 (N_16786,N_16625,N_16537);
nand U16787 (N_16787,N_16518,N_16557);
nor U16788 (N_16788,N_16607,N_16500);
xnor U16789 (N_16789,N_16523,N_16525);
and U16790 (N_16790,N_16524,N_16527);
and U16791 (N_16791,N_16687,N_16624);
nor U16792 (N_16792,N_16581,N_16503);
and U16793 (N_16793,N_16591,N_16606);
nand U16794 (N_16794,N_16565,N_16635);
nor U16795 (N_16795,N_16571,N_16661);
nor U16796 (N_16796,N_16704,N_16545);
or U16797 (N_16797,N_16663,N_16739);
xnor U16798 (N_16798,N_16595,N_16737);
nand U16799 (N_16799,N_16551,N_16522);
nor U16800 (N_16800,N_16566,N_16619);
and U16801 (N_16801,N_16552,N_16604);
xnor U16802 (N_16802,N_16539,N_16583);
and U16803 (N_16803,N_16532,N_16564);
or U16804 (N_16804,N_16602,N_16684);
nor U16805 (N_16805,N_16562,N_16659);
xor U16806 (N_16806,N_16612,N_16691);
nor U16807 (N_16807,N_16725,N_16636);
and U16808 (N_16808,N_16736,N_16743);
nor U16809 (N_16809,N_16719,N_16507);
nor U16810 (N_16810,N_16594,N_16544);
nor U16811 (N_16811,N_16548,N_16573);
nand U16812 (N_16812,N_16748,N_16615);
and U16813 (N_16813,N_16579,N_16600);
nand U16814 (N_16814,N_16575,N_16742);
nor U16815 (N_16815,N_16665,N_16643);
xor U16816 (N_16816,N_16715,N_16569);
nor U16817 (N_16817,N_16657,N_16598);
nor U16818 (N_16818,N_16582,N_16656);
and U16819 (N_16819,N_16631,N_16530);
nor U16820 (N_16820,N_16555,N_16711);
nor U16821 (N_16821,N_16658,N_16505);
nand U16822 (N_16822,N_16716,N_16618);
or U16823 (N_16823,N_16517,N_16589);
nor U16824 (N_16824,N_16511,N_16556);
xnor U16825 (N_16825,N_16601,N_16713);
and U16826 (N_16826,N_16570,N_16721);
nor U16827 (N_16827,N_16516,N_16536);
xor U16828 (N_16828,N_16633,N_16634);
and U16829 (N_16829,N_16533,N_16734);
nor U16830 (N_16830,N_16738,N_16681);
and U16831 (N_16831,N_16670,N_16655);
nand U16832 (N_16832,N_16679,N_16720);
and U16833 (N_16833,N_16741,N_16592);
nor U16834 (N_16834,N_16703,N_16702);
nor U16835 (N_16835,N_16672,N_16515);
and U16836 (N_16836,N_16647,N_16509);
nand U16837 (N_16837,N_16596,N_16669);
nor U16838 (N_16838,N_16699,N_16568);
nor U16839 (N_16839,N_16696,N_16677);
xnor U16840 (N_16840,N_16553,N_16746);
xor U16841 (N_16841,N_16559,N_16688);
xnor U16842 (N_16842,N_16626,N_16707);
and U16843 (N_16843,N_16652,N_16629);
nor U16844 (N_16844,N_16692,N_16542);
xnor U16845 (N_16845,N_16708,N_16529);
or U16846 (N_16846,N_16686,N_16709);
nand U16847 (N_16847,N_16668,N_16616);
xor U16848 (N_16848,N_16660,N_16560);
nor U16849 (N_16849,N_16567,N_16693);
xnor U16850 (N_16850,N_16608,N_16531);
xor U16851 (N_16851,N_16617,N_16697);
and U16852 (N_16852,N_16705,N_16590);
nor U16853 (N_16853,N_16623,N_16638);
nand U16854 (N_16854,N_16501,N_16727);
nor U16855 (N_16855,N_16521,N_16641);
nor U16856 (N_16856,N_16714,N_16680);
or U16857 (N_16857,N_16671,N_16586);
nand U16858 (N_16858,N_16729,N_16728);
nand U16859 (N_16859,N_16740,N_16724);
nand U16860 (N_16860,N_16577,N_16666);
and U16861 (N_16861,N_16667,N_16651);
or U16862 (N_16862,N_16588,N_16718);
and U16863 (N_16863,N_16611,N_16614);
and U16864 (N_16864,N_16694,N_16549);
or U16865 (N_16865,N_16563,N_16620);
and U16866 (N_16866,N_16621,N_16733);
xor U16867 (N_16867,N_16502,N_16558);
or U16868 (N_16868,N_16650,N_16508);
or U16869 (N_16869,N_16605,N_16712);
nand U16870 (N_16870,N_16597,N_16682);
nand U16871 (N_16871,N_16675,N_16561);
nor U16872 (N_16872,N_16649,N_16735);
and U16873 (N_16873,N_16554,N_16648);
or U16874 (N_16874,N_16639,N_16695);
and U16875 (N_16875,N_16595,N_16677);
nand U16876 (N_16876,N_16514,N_16708);
nor U16877 (N_16877,N_16544,N_16700);
and U16878 (N_16878,N_16739,N_16707);
nand U16879 (N_16879,N_16635,N_16689);
or U16880 (N_16880,N_16715,N_16580);
xor U16881 (N_16881,N_16679,N_16501);
xor U16882 (N_16882,N_16636,N_16685);
xnor U16883 (N_16883,N_16558,N_16556);
and U16884 (N_16884,N_16738,N_16711);
or U16885 (N_16885,N_16684,N_16507);
and U16886 (N_16886,N_16705,N_16688);
xor U16887 (N_16887,N_16596,N_16645);
nor U16888 (N_16888,N_16611,N_16661);
or U16889 (N_16889,N_16515,N_16543);
or U16890 (N_16890,N_16629,N_16737);
and U16891 (N_16891,N_16622,N_16616);
or U16892 (N_16892,N_16509,N_16639);
or U16893 (N_16893,N_16636,N_16622);
nand U16894 (N_16894,N_16519,N_16606);
nor U16895 (N_16895,N_16606,N_16739);
nor U16896 (N_16896,N_16712,N_16695);
or U16897 (N_16897,N_16664,N_16742);
xnor U16898 (N_16898,N_16681,N_16500);
or U16899 (N_16899,N_16728,N_16519);
xnor U16900 (N_16900,N_16519,N_16504);
nor U16901 (N_16901,N_16500,N_16590);
nand U16902 (N_16902,N_16718,N_16698);
and U16903 (N_16903,N_16615,N_16584);
or U16904 (N_16904,N_16702,N_16658);
and U16905 (N_16905,N_16608,N_16655);
xor U16906 (N_16906,N_16713,N_16560);
xor U16907 (N_16907,N_16578,N_16632);
or U16908 (N_16908,N_16587,N_16688);
xor U16909 (N_16909,N_16599,N_16598);
and U16910 (N_16910,N_16602,N_16634);
and U16911 (N_16911,N_16639,N_16678);
and U16912 (N_16912,N_16532,N_16572);
nand U16913 (N_16913,N_16573,N_16630);
or U16914 (N_16914,N_16577,N_16639);
nand U16915 (N_16915,N_16501,N_16618);
xor U16916 (N_16916,N_16694,N_16681);
nor U16917 (N_16917,N_16687,N_16701);
xnor U16918 (N_16918,N_16717,N_16699);
and U16919 (N_16919,N_16669,N_16698);
or U16920 (N_16920,N_16547,N_16534);
or U16921 (N_16921,N_16561,N_16540);
nand U16922 (N_16922,N_16700,N_16650);
or U16923 (N_16923,N_16522,N_16503);
xnor U16924 (N_16924,N_16572,N_16525);
nor U16925 (N_16925,N_16693,N_16557);
or U16926 (N_16926,N_16734,N_16650);
xnor U16927 (N_16927,N_16612,N_16565);
and U16928 (N_16928,N_16509,N_16580);
nand U16929 (N_16929,N_16507,N_16583);
or U16930 (N_16930,N_16528,N_16649);
or U16931 (N_16931,N_16741,N_16616);
and U16932 (N_16932,N_16530,N_16655);
or U16933 (N_16933,N_16591,N_16647);
or U16934 (N_16934,N_16617,N_16508);
nand U16935 (N_16935,N_16622,N_16515);
xnor U16936 (N_16936,N_16693,N_16649);
or U16937 (N_16937,N_16611,N_16578);
nand U16938 (N_16938,N_16593,N_16627);
or U16939 (N_16939,N_16505,N_16694);
or U16940 (N_16940,N_16614,N_16680);
or U16941 (N_16941,N_16562,N_16711);
nor U16942 (N_16942,N_16722,N_16570);
nor U16943 (N_16943,N_16551,N_16719);
xnor U16944 (N_16944,N_16729,N_16559);
or U16945 (N_16945,N_16544,N_16540);
or U16946 (N_16946,N_16748,N_16519);
and U16947 (N_16947,N_16665,N_16725);
or U16948 (N_16948,N_16527,N_16672);
xnor U16949 (N_16949,N_16568,N_16559);
and U16950 (N_16950,N_16693,N_16601);
nor U16951 (N_16951,N_16717,N_16518);
or U16952 (N_16952,N_16657,N_16500);
nor U16953 (N_16953,N_16513,N_16637);
and U16954 (N_16954,N_16588,N_16580);
or U16955 (N_16955,N_16532,N_16736);
xor U16956 (N_16956,N_16525,N_16594);
nor U16957 (N_16957,N_16535,N_16603);
xor U16958 (N_16958,N_16694,N_16716);
or U16959 (N_16959,N_16587,N_16639);
nor U16960 (N_16960,N_16561,N_16629);
xnor U16961 (N_16961,N_16644,N_16604);
xnor U16962 (N_16962,N_16688,N_16655);
nand U16963 (N_16963,N_16611,N_16606);
xnor U16964 (N_16964,N_16504,N_16656);
and U16965 (N_16965,N_16721,N_16565);
nand U16966 (N_16966,N_16671,N_16654);
or U16967 (N_16967,N_16738,N_16532);
xor U16968 (N_16968,N_16719,N_16643);
or U16969 (N_16969,N_16657,N_16665);
xnor U16970 (N_16970,N_16661,N_16647);
and U16971 (N_16971,N_16508,N_16561);
nor U16972 (N_16972,N_16711,N_16698);
or U16973 (N_16973,N_16656,N_16692);
nor U16974 (N_16974,N_16541,N_16559);
or U16975 (N_16975,N_16580,N_16591);
nor U16976 (N_16976,N_16629,N_16745);
and U16977 (N_16977,N_16682,N_16541);
xor U16978 (N_16978,N_16530,N_16667);
nor U16979 (N_16979,N_16578,N_16699);
xor U16980 (N_16980,N_16670,N_16500);
and U16981 (N_16981,N_16587,N_16669);
nor U16982 (N_16982,N_16731,N_16581);
or U16983 (N_16983,N_16546,N_16702);
nand U16984 (N_16984,N_16634,N_16512);
xnor U16985 (N_16985,N_16570,N_16566);
xor U16986 (N_16986,N_16533,N_16597);
and U16987 (N_16987,N_16537,N_16504);
xnor U16988 (N_16988,N_16728,N_16577);
nand U16989 (N_16989,N_16739,N_16630);
nor U16990 (N_16990,N_16566,N_16581);
nand U16991 (N_16991,N_16674,N_16657);
and U16992 (N_16992,N_16583,N_16551);
nor U16993 (N_16993,N_16534,N_16688);
xor U16994 (N_16994,N_16623,N_16729);
xor U16995 (N_16995,N_16735,N_16596);
and U16996 (N_16996,N_16636,N_16532);
nor U16997 (N_16997,N_16654,N_16641);
nand U16998 (N_16998,N_16513,N_16598);
nor U16999 (N_16999,N_16532,N_16519);
nand U17000 (N_17000,N_16832,N_16828);
and U17001 (N_17001,N_16790,N_16997);
xor U17002 (N_17002,N_16895,N_16958);
nor U17003 (N_17003,N_16835,N_16773);
or U17004 (N_17004,N_16827,N_16865);
nand U17005 (N_17005,N_16785,N_16826);
or U17006 (N_17006,N_16989,N_16899);
and U17007 (N_17007,N_16880,N_16769);
nor U17008 (N_17008,N_16890,N_16882);
and U17009 (N_17009,N_16933,N_16888);
nor U17010 (N_17010,N_16876,N_16981);
nor U17011 (N_17011,N_16818,N_16753);
nor U17012 (N_17012,N_16988,N_16868);
nor U17013 (N_17013,N_16794,N_16853);
and U17014 (N_17014,N_16873,N_16952);
or U17015 (N_17015,N_16795,N_16805);
or U17016 (N_17016,N_16966,N_16938);
xnor U17017 (N_17017,N_16979,N_16846);
nand U17018 (N_17018,N_16945,N_16812);
or U17019 (N_17019,N_16934,N_16816);
nor U17020 (N_17020,N_16810,N_16807);
xnor U17021 (N_17021,N_16841,N_16776);
and U17022 (N_17022,N_16964,N_16842);
nor U17023 (N_17023,N_16834,N_16990);
xnor U17024 (N_17024,N_16922,N_16781);
nor U17025 (N_17025,N_16970,N_16800);
xnor U17026 (N_17026,N_16968,N_16869);
and U17027 (N_17027,N_16931,N_16960);
or U17028 (N_17028,N_16896,N_16954);
nor U17029 (N_17029,N_16949,N_16774);
and U17030 (N_17030,N_16892,N_16768);
and U17031 (N_17031,N_16755,N_16914);
or U17032 (N_17032,N_16983,N_16856);
and U17033 (N_17033,N_16920,N_16811);
and U17034 (N_17034,N_16925,N_16986);
nand U17035 (N_17035,N_16940,N_16959);
xor U17036 (N_17036,N_16994,N_16961);
and U17037 (N_17037,N_16845,N_16760);
and U17038 (N_17038,N_16916,N_16849);
xnor U17039 (N_17039,N_16917,N_16763);
or U17040 (N_17040,N_16972,N_16829);
nand U17041 (N_17041,N_16782,N_16991);
nor U17042 (N_17042,N_16787,N_16900);
nand U17043 (N_17043,N_16867,N_16973);
or U17044 (N_17044,N_16801,N_16766);
nand U17045 (N_17045,N_16941,N_16779);
xnor U17046 (N_17046,N_16935,N_16798);
and U17047 (N_17047,N_16944,N_16783);
nor U17048 (N_17048,N_16859,N_16775);
or U17049 (N_17049,N_16885,N_16955);
or U17050 (N_17050,N_16919,N_16975);
nand U17051 (N_17051,N_16759,N_16854);
xnor U17052 (N_17052,N_16821,N_16861);
nand U17053 (N_17053,N_16967,N_16943);
nor U17054 (N_17054,N_16850,N_16843);
and U17055 (N_17055,N_16847,N_16809);
and U17056 (N_17056,N_16980,N_16995);
nand U17057 (N_17057,N_16878,N_16784);
xnor U17058 (N_17058,N_16956,N_16864);
or U17059 (N_17059,N_16751,N_16984);
xnor U17060 (N_17060,N_16871,N_16824);
and U17061 (N_17061,N_16965,N_16802);
and U17062 (N_17062,N_16905,N_16918);
nand U17063 (N_17063,N_16806,N_16953);
or U17064 (N_17064,N_16761,N_16901);
xnor U17065 (N_17065,N_16870,N_16887);
nor U17066 (N_17066,N_16808,N_16894);
and U17067 (N_17067,N_16881,N_16862);
or U17068 (N_17068,N_16912,N_16891);
xnor U17069 (N_17069,N_16921,N_16998);
nand U17070 (N_17070,N_16874,N_16903);
nor U17071 (N_17071,N_16839,N_16976);
or U17072 (N_17072,N_16883,N_16996);
and U17073 (N_17073,N_16822,N_16758);
nor U17074 (N_17074,N_16957,N_16772);
and U17075 (N_17075,N_16978,N_16778);
xnor U17076 (N_17076,N_16908,N_16992);
xor U17077 (N_17077,N_16804,N_16770);
or U17078 (N_17078,N_16937,N_16797);
and U17079 (N_17079,N_16926,N_16942);
nor U17080 (N_17080,N_16929,N_16857);
and U17081 (N_17081,N_16757,N_16993);
and U17082 (N_17082,N_16789,N_16982);
nor U17083 (N_17083,N_16844,N_16928);
xnor U17084 (N_17084,N_16788,N_16915);
nand U17085 (N_17085,N_16792,N_16819);
or U17086 (N_17086,N_16863,N_16820);
nand U17087 (N_17087,N_16963,N_16813);
and U17088 (N_17088,N_16750,N_16754);
and U17089 (N_17089,N_16879,N_16799);
or U17090 (N_17090,N_16791,N_16907);
nor U17091 (N_17091,N_16947,N_16817);
nand U17092 (N_17092,N_16971,N_16946);
nor U17093 (N_17093,N_16950,N_16803);
nand U17094 (N_17094,N_16756,N_16927);
or U17095 (N_17095,N_16889,N_16886);
xnor U17096 (N_17096,N_16974,N_16777);
or U17097 (N_17097,N_16999,N_16877);
and U17098 (N_17098,N_16830,N_16767);
nor U17099 (N_17099,N_16765,N_16969);
and U17100 (N_17100,N_16904,N_16884);
nor U17101 (N_17101,N_16897,N_16898);
nand U17102 (N_17102,N_16815,N_16902);
nor U17103 (N_17103,N_16825,N_16823);
and U17104 (N_17104,N_16923,N_16780);
and U17105 (N_17105,N_16848,N_16793);
or U17106 (N_17106,N_16911,N_16858);
and U17107 (N_17107,N_16936,N_16932);
nor U17108 (N_17108,N_16930,N_16831);
xnor U17109 (N_17109,N_16962,N_16939);
xor U17110 (N_17110,N_16771,N_16764);
and U17111 (N_17111,N_16837,N_16836);
xor U17112 (N_17112,N_16893,N_16906);
xor U17113 (N_17113,N_16987,N_16948);
or U17114 (N_17114,N_16866,N_16833);
nor U17115 (N_17115,N_16838,N_16977);
and U17116 (N_17116,N_16796,N_16851);
nand U17117 (N_17117,N_16924,N_16951);
nor U17118 (N_17118,N_16762,N_16840);
or U17119 (N_17119,N_16855,N_16909);
xnor U17120 (N_17120,N_16913,N_16910);
nor U17121 (N_17121,N_16875,N_16985);
and U17122 (N_17122,N_16872,N_16752);
xor U17123 (N_17123,N_16814,N_16786);
nand U17124 (N_17124,N_16860,N_16852);
xnor U17125 (N_17125,N_16883,N_16782);
and U17126 (N_17126,N_16928,N_16977);
nor U17127 (N_17127,N_16900,N_16923);
xor U17128 (N_17128,N_16959,N_16750);
and U17129 (N_17129,N_16950,N_16984);
nand U17130 (N_17130,N_16992,N_16979);
and U17131 (N_17131,N_16854,N_16831);
or U17132 (N_17132,N_16972,N_16760);
nand U17133 (N_17133,N_16887,N_16908);
or U17134 (N_17134,N_16996,N_16800);
or U17135 (N_17135,N_16791,N_16995);
xor U17136 (N_17136,N_16961,N_16931);
xor U17137 (N_17137,N_16858,N_16914);
nor U17138 (N_17138,N_16996,N_16918);
nor U17139 (N_17139,N_16971,N_16783);
and U17140 (N_17140,N_16980,N_16881);
or U17141 (N_17141,N_16788,N_16784);
or U17142 (N_17142,N_16761,N_16843);
nand U17143 (N_17143,N_16759,N_16792);
or U17144 (N_17144,N_16855,N_16908);
nand U17145 (N_17145,N_16768,N_16983);
or U17146 (N_17146,N_16925,N_16820);
xor U17147 (N_17147,N_16920,N_16753);
nor U17148 (N_17148,N_16961,N_16964);
and U17149 (N_17149,N_16949,N_16813);
or U17150 (N_17150,N_16947,N_16989);
or U17151 (N_17151,N_16977,N_16948);
xor U17152 (N_17152,N_16892,N_16985);
or U17153 (N_17153,N_16930,N_16975);
nand U17154 (N_17154,N_16843,N_16926);
nand U17155 (N_17155,N_16794,N_16968);
xnor U17156 (N_17156,N_16994,N_16819);
nand U17157 (N_17157,N_16846,N_16805);
or U17158 (N_17158,N_16928,N_16920);
and U17159 (N_17159,N_16864,N_16981);
or U17160 (N_17160,N_16989,N_16893);
or U17161 (N_17161,N_16821,N_16937);
or U17162 (N_17162,N_16760,N_16910);
nand U17163 (N_17163,N_16839,N_16856);
nor U17164 (N_17164,N_16943,N_16879);
nor U17165 (N_17165,N_16975,N_16757);
nor U17166 (N_17166,N_16781,N_16949);
nand U17167 (N_17167,N_16829,N_16999);
and U17168 (N_17168,N_16783,N_16787);
and U17169 (N_17169,N_16826,N_16967);
nand U17170 (N_17170,N_16868,N_16898);
or U17171 (N_17171,N_16755,N_16800);
nor U17172 (N_17172,N_16758,N_16812);
nand U17173 (N_17173,N_16935,N_16814);
nor U17174 (N_17174,N_16950,N_16773);
or U17175 (N_17175,N_16915,N_16845);
nor U17176 (N_17176,N_16870,N_16944);
xor U17177 (N_17177,N_16994,N_16891);
or U17178 (N_17178,N_16830,N_16772);
and U17179 (N_17179,N_16771,N_16854);
xor U17180 (N_17180,N_16960,N_16777);
and U17181 (N_17181,N_16770,N_16821);
nor U17182 (N_17182,N_16910,N_16872);
xor U17183 (N_17183,N_16873,N_16808);
or U17184 (N_17184,N_16851,N_16808);
or U17185 (N_17185,N_16772,N_16865);
or U17186 (N_17186,N_16790,N_16974);
nor U17187 (N_17187,N_16983,N_16955);
nor U17188 (N_17188,N_16973,N_16926);
and U17189 (N_17189,N_16976,N_16885);
xnor U17190 (N_17190,N_16965,N_16757);
and U17191 (N_17191,N_16760,N_16927);
and U17192 (N_17192,N_16977,N_16786);
and U17193 (N_17193,N_16879,N_16828);
and U17194 (N_17194,N_16927,N_16976);
nand U17195 (N_17195,N_16832,N_16919);
and U17196 (N_17196,N_16793,N_16866);
nand U17197 (N_17197,N_16972,N_16865);
nand U17198 (N_17198,N_16825,N_16992);
nor U17199 (N_17199,N_16976,N_16856);
xnor U17200 (N_17200,N_16923,N_16915);
nor U17201 (N_17201,N_16991,N_16913);
or U17202 (N_17202,N_16946,N_16768);
or U17203 (N_17203,N_16950,N_16763);
nand U17204 (N_17204,N_16864,N_16960);
nor U17205 (N_17205,N_16821,N_16767);
and U17206 (N_17206,N_16948,N_16879);
nand U17207 (N_17207,N_16963,N_16822);
nor U17208 (N_17208,N_16875,N_16906);
nand U17209 (N_17209,N_16971,N_16850);
nand U17210 (N_17210,N_16828,N_16972);
and U17211 (N_17211,N_16844,N_16904);
or U17212 (N_17212,N_16917,N_16916);
nor U17213 (N_17213,N_16789,N_16973);
nor U17214 (N_17214,N_16893,N_16837);
nand U17215 (N_17215,N_16814,N_16788);
nand U17216 (N_17216,N_16765,N_16986);
or U17217 (N_17217,N_16987,N_16883);
nor U17218 (N_17218,N_16859,N_16943);
nor U17219 (N_17219,N_16853,N_16846);
and U17220 (N_17220,N_16927,N_16968);
xnor U17221 (N_17221,N_16928,N_16934);
or U17222 (N_17222,N_16765,N_16949);
and U17223 (N_17223,N_16804,N_16924);
and U17224 (N_17224,N_16778,N_16841);
xnor U17225 (N_17225,N_16964,N_16760);
xnor U17226 (N_17226,N_16953,N_16957);
and U17227 (N_17227,N_16906,N_16946);
nor U17228 (N_17228,N_16937,N_16855);
or U17229 (N_17229,N_16818,N_16825);
xnor U17230 (N_17230,N_16902,N_16794);
nor U17231 (N_17231,N_16751,N_16880);
or U17232 (N_17232,N_16956,N_16959);
nand U17233 (N_17233,N_16750,N_16954);
nand U17234 (N_17234,N_16858,N_16842);
or U17235 (N_17235,N_16818,N_16913);
or U17236 (N_17236,N_16787,N_16997);
and U17237 (N_17237,N_16805,N_16928);
and U17238 (N_17238,N_16973,N_16846);
xnor U17239 (N_17239,N_16948,N_16953);
nand U17240 (N_17240,N_16815,N_16833);
nand U17241 (N_17241,N_16979,N_16761);
and U17242 (N_17242,N_16840,N_16826);
xnor U17243 (N_17243,N_16971,N_16858);
nor U17244 (N_17244,N_16789,N_16957);
or U17245 (N_17245,N_16923,N_16869);
nor U17246 (N_17246,N_16758,N_16911);
nor U17247 (N_17247,N_16846,N_16912);
and U17248 (N_17248,N_16985,N_16954);
nand U17249 (N_17249,N_16758,N_16999);
xor U17250 (N_17250,N_17171,N_17190);
or U17251 (N_17251,N_17203,N_17202);
or U17252 (N_17252,N_17162,N_17241);
nor U17253 (N_17253,N_17160,N_17245);
nand U17254 (N_17254,N_17169,N_17006);
nand U17255 (N_17255,N_17211,N_17034);
and U17256 (N_17256,N_17213,N_17007);
xor U17257 (N_17257,N_17189,N_17037);
nor U17258 (N_17258,N_17236,N_17217);
nand U17259 (N_17259,N_17188,N_17041);
and U17260 (N_17260,N_17095,N_17094);
or U17261 (N_17261,N_17248,N_17170);
or U17262 (N_17262,N_17100,N_17051);
xor U17263 (N_17263,N_17042,N_17050);
nand U17264 (N_17264,N_17043,N_17145);
nor U17265 (N_17265,N_17087,N_17226);
or U17266 (N_17266,N_17018,N_17085);
and U17267 (N_17267,N_17235,N_17101);
and U17268 (N_17268,N_17026,N_17147);
and U17269 (N_17269,N_17175,N_17194);
nand U17270 (N_17270,N_17127,N_17104);
nand U17271 (N_17271,N_17179,N_17080);
nand U17272 (N_17272,N_17205,N_17193);
nor U17273 (N_17273,N_17128,N_17238);
nand U17274 (N_17274,N_17022,N_17064);
or U17275 (N_17275,N_17218,N_17216);
xnor U17276 (N_17276,N_17137,N_17232);
and U17277 (N_17277,N_17060,N_17125);
nor U17278 (N_17278,N_17174,N_17068);
and U17279 (N_17279,N_17053,N_17163);
or U17280 (N_17280,N_17224,N_17052);
and U17281 (N_17281,N_17214,N_17161);
nand U17282 (N_17282,N_17001,N_17013);
or U17283 (N_17283,N_17230,N_17075);
nor U17284 (N_17284,N_17021,N_17110);
and U17285 (N_17285,N_17047,N_17166);
and U17286 (N_17286,N_17143,N_17221);
nor U17287 (N_17287,N_17005,N_17196);
xor U17288 (N_17288,N_17112,N_17209);
or U17289 (N_17289,N_17126,N_17197);
and U17290 (N_17290,N_17191,N_17144);
and U17291 (N_17291,N_17164,N_17182);
and U17292 (N_17292,N_17054,N_17017);
nand U17293 (N_17293,N_17072,N_17219);
nor U17294 (N_17294,N_17183,N_17186);
nand U17295 (N_17295,N_17132,N_17176);
nand U17296 (N_17296,N_17228,N_17082);
nand U17297 (N_17297,N_17098,N_17071);
nor U17298 (N_17298,N_17012,N_17016);
nor U17299 (N_17299,N_17033,N_17124);
and U17300 (N_17300,N_17195,N_17215);
xor U17301 (N_17301,N_17056,N_17222);
nor U17302 (N_17302,N_17247,N_17220);
xnor U17303 (N_17303,N_17208,N_17008);
and U17304 (N_17304,N_17011,N_17078);
xor U17305 (N_17305,N_17083,N_17185);
and U17306 (N_17306,N_17158,N_17246);
nand U17307 (N_17307,N_17045,N_17129);
xor U17308 (N_17308,N_17058,N_17069);
and U17309 (N_17309,N_17155,N_17131);
nand U17310 (N_17310,N_17115,N_17146);
or U17311 (N_17311,N_17009,N_17020);
or U17312 (N_17312,N_17172,N_17181);
nor U17313 (N_17313,N_17210,N_17074);
nor U17314 (N_17314,N_17107,N_17136);
nand U17315 (N_17315,N_17059,N_17118);
nand U17316 (N_17316,N_17027,N_17184);
xor U17317 (N_17317,N_17010,N_17204);
xor U17318 (N_17318,N_17229,N_17103);
or U17319 (N_17319,N_17000,N_17138);
or U17320 (N_17320,N_17063,N_17057);
and U17321 (N_17321,N_17201,N_17105);
nor U17322 (N_17322,N_17106,N_17091);
nand U17323 (N_17323,N_17242,N_17200);
or U17324 (N_17324,N_17090,N_17154);
nand U17325 (N_17325,N_17240,N_17140);
nor U17326 (N_17326,N_17055,N_17117);
xor U17327 (N_17327,N_17157,N_17062);
or U17328 (N_17328,N_17130,N_17123);
and U17329 (N_17329,N_17156,N_17014);
or U17330 (N_17330,N_17116,N_17084);
xor U17331 (N_17331,N_17111,N_17077);
xnor U17332 (N_17332,N_17233,N_17113);
nor U17333 (N_17333,N_17225,N_17038);
nand U17334 (N_17334,N_17023,N_17119);
or U17335 (N_17335,N_17092,N_17249);
or U17336 (N_17336,N_17120,N_17093);
or U17337 (N_17337,N_17173,N_17108);
nor U17338 (N_17338,N_17079,N_17243);
xnor U17339 (N_17339,N_17048,N_17046);
xor U17340 (N_17340,N_17061,N_17036);
and U17341 (N_17341,N_17040,N_17028);
nand U17342 (N_17342,N_17044,N_17151);
and U17343 (N_17343,N_17168,N_17002);
xor U17344 (N_17344,N_17035,N_17134);
xnor U17345 (N_17345,N_17153,N_17109);
nand U17346 (N_17346,N_17239,N_17025);
nor U17347 (N_17347,N_17207,N_17029);
or U17348 (N_17348,N_17159,N_17133);
nor U17349 (N_17349,N_17081,N_17142);
xnor U17350 (N_17350,N_17032,N_17167);
nand U17351 (N_17351,N_17148,N_17076);
nor U17352 (N_17352,N_17073,N_17070);
nor U17353 (N_17353,N_17019,N_17024);
xnor U17354 (N_17354,N_17198,N_17097);
xor U17355 (N_17355,N_17122,N_17030);
or U17356 (N_17356,N_17199,N_17152);
xnor U17357 (N_17357,N_17244,N_17089);
nand U17358 (N_17358,N_17031,N_17227);
xnor U17359 (N_17359,N_17150,N_17065);
or U17360 (N_17360,N_17141,N_17223);
nand U17361 (N_17361,N_17212,N_17165);
or U17362 (N_17362,N_17237,N_17187);
nand U17363 (N_17363,N_17067,N_17139);
and U17364 (N_17364,N_17234,N_17102);
nand U17365 (N_17365,N_17192,N_17206);
xnor U17366 (N_17366,N_17177,N_17114);
or U17367 (N_17367,N_17088,N_17231);
and U17368 (N_17368,N_17178,N_17099);
nand U17369 (N_17369,N_17003,N_17049);
nand U17370 (N_17370,N_17039,N_17066);
nand U17371 (N_17371,N_17135,N_17015);
nand U17372 (N_17372,N_17121,N_17096);
xnor U17373 (N_17373,N_17149,N_17086);
or U17374 (N_17374,N_17180,N_17004);
nand U17375 (N_17375,N_17088,N_17096);
or U17376 (N_17376,N_17210,N_17006);
or U17377 (N_17377,N_17098,N_17000);
or U17378 (N_17378,N_17118,N_17035);
nor U17379 (N_17379,N_17150,N_17082);
or U17380 (N_17380,N_17034,N_17188);
nor U17381 (N_17381,N_17113,N_17144);
nor U17382 (N_17382,N_17073,N_17247);
nand U17383 (N_17383,N_17092,N_17056);
or U17384 (N_17384,N_17108,N_17098);
nand U17385 (N_17385,N_17021,N_17209);
xnor U17386 (N_17386,N_17167,N_17152);
and U17387 (N_17387,N_17143,N_17215);
nor U17388 (N_17388,N_17007,N_17164);
or U17389 (N_17389,N_17082,N_17135);
xnor U17390 (N_17390,N_17026,N_17217);
or U17391 (N_17391,N_17001,N_17188);
or U17392 (N_17392,N_17043,N_17098);
nor U17393 (N_17393,N_17235,N_17088);
or U17394 (N_17394,N_17218,N_17009);
or U17395 (N_17395,N_17024,N_17158);
nand U17396 (N_17396,N_17078,N_17213);
and U17397 (N_17397,N_17066,N_17124);
xnor U17398 (N_17398,N_17121,N_17230);
nand U17399 (N_17399,N_17082,N_17249);
nand U17400 (N_17400,N_17213,N_17032);
xor U17401 (N_17401,N_17152,N_17046);
and U17402 (N_17402,N_17212,N_17043);
xor U17403 (N_17403,N_17219,N_17165);
nor U17404 (N_17404,N_17072,N_17249);
and U17405 (N_17405,N_17058,N_17205);
xor U17406 (N_17406,N_17218,N_17214);
xor U17407 (N_17407,N_17193,N_17153);
nor U17408 (N_17408,N_17204,N_17232);
and U17409 (N_17409,N_17167,N_17103);
nor U17410 (N_17410,N_17246,N_17077);
or U17411 (N_17411,N_17146,N_17087);
nor U17412 (N_17412,N_17094,N_17103);
xnor U17413 (N_17413,N_17041,N_17224);
xor U17414 (N_17414,N_17100,N_17078);
or U17415 (N_17415,N_17094,N_17062);
or U17416 (N_17416,N_17206,N_17012);
nor U17417 (N_17417,N_17019,N_17020);
and U17418 (N_17418,N_17242,N_17219);
and U17419 (N_17419,N_17027,N_17054);
nor U17420 (N_17420,N_17246,N_17206);
nor U17421 (N_17421,N_17071,N_17041);
nor U17422 (N_17422,N_17013,N_17036);
nand U17423 (N_17423,N_17109,N_17031);
nand U17424 (N_17424,N_17043,N_17172);
or U17425 (N_17425,N_17020,N_17134);
xnor U17426 (N_17426,N_17080,N_17222);
nor U17427 (N_17427,N_17202,N_17024);
or U17428 (N_17428,N_17219,N_17019);
xnor U17429 (N_17429,N_17107,N_17013);
nand U17430 (N_17430,N_17031,N_17058);
and U17431 (N_17431,N_17088,N_17114);
or U17432 (N_17432,N_17178,N_17146);
nor U17433 (N_17433,N_17216,N_17046);
and U17434 (N_17434,N_17160,N_17156);
or U17435 (N_17435,N_17197,N_17165);
nand U17436 (N_17436,N_17021,N_17211);
xnor U17437 (N_17437,N_17197,N_17007);
xnor U17438 (N_17438,N_17171,N_17002);
or U17439 (N_17439,N_17022,N_17194);
nand U17440 (N_17440,N_17087,N_17015);
or U17441 (N_17441,N_17189,N_17123);
or U17442 (N_17442,N_17198,N_17021);
or U17443 (N_17443,N_17036,N_17022);
nand U17444 (N_17444,N_17118,N_17040);
nor U17445 (N_17445,N_17196,N_17042);
or U17446 (N_17446,N_17105,N_17005);
and U17447 (N_17447,N_17044,N_17129);
nand U17448 (N_17448,N_17019,N_17176);
nor U17449 (N_17449,N_17225,N_17216);
or U17450 (N_17450,N_17216,N_17021);
xnor U17451 (N_17451,N_17181,N_17230);
nand U17452 (N_17452,N_17126,N_17147);
xor U17453 (N_17453,N_17179,N_17037);
xnor U17454 (N_17454,N_17221,N_17061);
xnor U17455 (N_17455,N_17222,N_17059);
nor U17456 (N_17456,N_17101,N_17023);
or U17457 (N_17457,N_17113,N_17055);
nor U17458 (N_17458,N_17239,N_17121);
xnor U17459 (N_17459,N_17091,N_17126);
nand U17460 (N_17460,N_17191,N_17079);
nor U17461 (N_17461,N_17062,N_17153);
and U17462 (N_17462,N_17171,N_17018);
nor U17463 (N_17463,N_17197,N_17074);
nor U17464 (N_17464,N_17183,N_17065);
and U17465 (N_17465,N_17053,N_17216);
and U17466 (N_17466,N_17098,N_17238);
nor U17467 (N_17467,N_17083,N_17222);
xor U17468 (N_17468,N_17008,N_17085);
or U17469 (N_17469,N_17070,N_17124);
nand U17470 (N_17470,N_17189,N_17091);
nand U17471 (N_17471,N_17210,N_17094);
nor U17472 (N_17472,N_17117,N_17236);
nor U17473 (N_17473,N_17248,N_17115);
or U17474 (N_17474,N_17100,N_17046);
or U17475 (N_17475,N_17177,N_17174);
nand U17476 (N_17476,N_17163,N_17000);
nor U17477 (N_17477,N_17091,N_17132);
xor U17478 (N_17478,N_17055,N_17232);
xnor U17479 (N_17479,N_17049,N_17130);
or U17480 (N_17480,N_17161,N_17038);
or U17481 (N_17481,N_17001,N_17116);
xor U17482 (N_17482,N_17028,N_17073);
and U17483 (N_17483,N_17168,N_17219);
and U17484 (N_17484,N_17213,N_17022);
nand U17485 (N_17485,N_17043,N_17190);
and U17486 (N_17486,N_17165,N_17143);
nor U17487 (N_17487,N_17048,N_17137);
or U17488 (N_17488,N_17162,N_17187);
nand U17489 (N_17489,N_17057,N_17126);
xor U17490 (N_17490,N_17032,N_17106);
or U17491 (N_17491,N_17140,N_17018);
nor U17492 (N_17492,N_17014,N_17141);
or U17493 (N_17493,N_17231,N_17035);
or U17494 (N_17494,N_17205,N_17137);
xor U17495 (N_17495,N_17026,N_17081);
and U17496 (N_17496,N_17111,N_17084);
or U17497 (N_17497,N_17034,N_17125);
or U17498 (N_17498,N_17045,N_17052);
or U17499 (N_17499,N_17006,N_17080);
xor U17500 (N_17500,N_17338,N_17299);
nor U17501 (N_17501,N_17297,N_17319);
or U17502 (N_17502,N_17381,N_17369);
nor U17503 (N_17503,N_17336,N_17474);
nor U17504 (N_17504,N_17291,N_17422);
and U17505 (N_17505,N_17451,N_17473);
nor U17506 (N_17506,N_17435,N_17288);
nor U17507 (N_17507,N_17421,N_17441);
or U17508 (N_17508,N_17337,N_17427);
xor U17509 (N_17509,N_17402,N_17325);
nand U17510 (N_17510,N_17386,N_17418);
or U17511 (N_17511,N_17498,N_17412);
and U17512 (N_17512,N_17356,N_17497);
or U17513 (N_17513,N_17290,N_17493);
nor U17514 (N_17514,N_17256,N_17433);
nand U17515 (N_17515,N_17476,N_17255);
xnor U17516 (N_17516,N_17387,N_17280);
and U17517 (N_17517,N_17283,N_17431);
and U17518 (N_17518,N_17357,N_17376);
and U17519 (N_17519,N_17355,N_17490);
xnor U17520 (N_17520,N_17467,N_17317);
nor U17521 (N_17521,N_17274,N_17465);
or U17522 (N_17522,N_17460,N_17442);
and U17523 (N_17523,N_17349,N_17411);
xor U17524 (N_17524,N_17443,N_17273);
or U17525 (N_17525,N_17437,N_17482);
or U17526 (N_17526,N_17454,N_17373);
or U17527 (N_17527,N_17420,N_17471);
nor U17528 (N_17528,N_17271,N_17446);
xnor U17529 (N_17529,N_17258,N_17466);
nor U17530 (N_17530,N_17259,N_17453);
or U17531 (N_17531,N_17368,N_17250);
and U17532 (N_17532,N_17254,N_17415);
and U17533 (N_17533,N_17408,N_17303);
or U17534 (N_17534,N_17417,N_17392);
and U17535 (N_17535,N_17276,N_17331);
nor U17536 (N_17536,N_17360,N_17456);
nor U17537 (N_17537,N_17486,N_17322);
nand U17538 (N_17538,N_17472,N_17440);
and U17539 (N_17539,N_17345,N_17404);
and U17540 (N_17540,N_17300,N_17333);
nor U17541 (N_17541,N_17313,N_17372);
or U17542 (N_17542,N_17301,N_17398);
and U17543 (N_17543,N_17439,N_17270);
and U17544 (N_17544,N_17455,N_17468);
and U17545 (N_17545,N_17265,N_17430);
and U17546 (N_17546,N_17298,N_17310);
or U17547 (N_17547,N_17496,N_17307);
xnor U17548 (N_17548,N_17449,N_17461);
xnor U17549 (N_17549,N_17479,N_17304);
nor U17550 (N_17550,N_17399,N_17475);
or U17551 (N_17551,N_17395,N_17286);
or U17552 (N_17552,N_17306,N_17414);
and U17553 (N_17553,N_17374,N_17406);
nand U17554 (N_17554,N_17393,N_17292);
xnor U17555 (N_17555,N_17407,N_17269);
or U17556 (N_17556,N_17302,N_17428);
nand U17557 (N_17557,N_17383,N_17278);
nor U17558 (N_17558,N_17483,N_17409);
xor U17559 (N_17559,N_17293,N_17457);
nand U17560 (N_17560,N_17448,N_17309);
nand U17561 (N_17561,N_17429,N_17257);
nor U17562 (N_17562,N_17295,N_17321);
nor U17563 (N_17563,N_17346,N_17312);
nand U17564 (N_17564,N_17328,N_17339);
xor U17565 (N_17565,N_17492,N_17423);
and U17566 (N_17566,N_17327,N_17389);
and U17567 (N_17567,N_17330,N_17268);
nor U17568 (N_17568,N_17315,N_17401);
nor U17569 (N_17569,N_17463,N_17484);
nor U17570 (N_17570,N_17350,N_17478);
xor U17571 (N_17571,N_17397,N_17488);
and U17572 (N_17572,N_17489,N_17445);
xnor U17573 (N_17573,N_17450,N_17294);
and U17574 (N_17574,N_17491,N_17400);
or U17575 (N_17575,N_17361,N_17377);
nand U17576 (N_17576,N_17348,N_17385);
nor U17577 (N_17577,N_17436,N_17284);
xor U17578 (N_17578,N_17470,N_17364);
and U17579 (N_17579,N_17260,N_17316);
or U17580 (N_17580,N_17266,N_17391);
xnor U17581 (N_17581,N_17394,N_17359);
nor U17582 (N_17582,N_17324,N_17379);
xnor U17583 (N_17583,N_17252,N_17424);
xnor U17584 (N_17584,N_17494,N_17347);
nand U17585 (N_17585,N_17326,N_17480);
and U17586 (N_17586,N_17426,N_17267);
and U17587 (N_17587,N_17481,N_17447);
or U17588 (N_17588,N_17287,N_17277);
nand U17589 (N_17589,N_17363,N_17279);
or U17590 (N_17590,N_17344,N_17444);
and U17591 (N_17591,N_17434,N_17485);
nand U17592 (N_17592,N_17469,N_17341);
or U17593 (N_17593,N_17495,N_17419);
nand U17594 (N_17594,N_17318,N_17308);
and U17595 (N_17595,N_17464,N_17378);
and U17596 (N_17596,N_17261,N_17388);
or U17597 (N_17597,N_17438,N_17281);
or U17598 (N_17598,N_17410,N_17452);
and U17599 (N_17599,N_17329,N_17396);
and U17600 (N_17600,N_17499,N_17371);
or U17601 (N_17601,N_17262,N_17384);
and U17602 (N_17602,N_17366,N_17289);
nand U17603 (N_17603,N_17403,N_17311);
nor U17604 (N_17604,N_17251,N_17390);
nor U17605 (N_17605,N_17365,N_17405);
nand U17606 (N_17606,N_17352,N_17370);
nand U17607 (N_17607,N_17354,N_17351);
or U17608 (N_17608,N_17432,N_17358);
and U17609 (N_17609,N_17416,N_17314);
or U17610 (N_17610,N_17272,N_17342);
or U17611 (N_17611,N_17425,N_17282);
or U17612 (N_17612,N_17263,N_17459);
xor U17613 (N_17613,N_17477,N_17380);
xor U17614 (N_17614,N_17296,N_17320);
nand U17615 (N_17615,N_17264,N_17343);
and U17616 (N_17616,N_17275,N_17305);
nand U17617 (N_17617,N_17462,N_17323);
xor U17618 (N_17618,N_17340,N_17382);
xor U17619 (N_17619,N_17367,N_17353);
and U17620 (N_17620,N_17285,N_17334);
xnor U17621 (N_17621,N_17253,N_17487);
nor U17622 (N_17622,N_17458,N_17375);
xor U17623 (N_17623,N_17332,N_17413);
or U17624 (N_17624,N_17362,N_17335);
nand U17625 (N_17625,N_17338,N_17487);
nor U17626 (N_17626,N_17433,N_17253);
and U17627 (N_17627,N_17276,N_17359);
or U17628 (N_17628,N_17447,N_17367);
or U17629 (N_17629,N_17366,N_17491);
nor U17630 (N_17630,N_17466,N_17380);
nand U17631 (N_17631,N_17471,N_17433);
nand U17632 (N_17632,N_17293,N_17452);
and U17633 (N_17633,N_17318,N_17430);
nor U17634 (N_17634,N_17275,N_17294);
nand U17635 (N_17635,N_17476,N_17392);
and U17636 (N_17636,N_17427,N_17289);
or U17637 (N_17637,N_17498,N_17291);
or U17638 (N_17638,N_17474,N_17297);
nand U17639 (N_17639,N_17263,N_17311);
xnor U17640 (N_17640,N_17282,N_17461);
nand U17641 (N_17641,N_17309,N_17390);
and U17642 (N_17642,N_17278,N_17252);
nor U17643 (N_17643,N_17455,N_17312);
xor U17644 (N_17644,N_17340,N_17339);
and U17645 (N_17645,N_17468,N_17297);
nor U17646 (N_17646,N_17412,N_17318);
nand U17647 (N_17647,N_17398,N_17378);
and U17648 (N_17648,N_17383,N_17352);
nor U17649 (N_17649,N_17292,N_17308);
nor U17650 (N_17650,N_17398,N_17423);
or U17651 (N_17651,N_17387,N_17407);
xnor U17652 (N_17652,N_17410,N_17311);
nor U17653 (N_17653,N_17395,N_17291);
nand U17654 (N_17654,N_17280,N_17307);
or U17655 (N_17655,N_17333,N_17378);
nand U17656 (N_17656,N_17348,N_17381);
nand U17657 (N_17657,N_17384,N_17402);
and U17658 (N_17658,N_17424,N_17422);
xor U17659 (N_17659,N_17483,N_17449);
nand U17660 (N_17660,N_17250,N_17280);
nor U17661 (N_17661,N_17431,N_17338);
xnor U17662 (N_17662,N_17295,N_17336);
or U17663 (N_17663,N_17379,N_17442);
nor U17664 (N_17664,N_17325,N_17354);
and U17665 (N_17665,N_17472,N_17460);
and U17666 (N_17666,N_17455,N_17473);
xor U17667 (N_17667,N_17425,N_17428);
nand U17668 (N_17668,N_17379,N_17268);
and U17669 (N_17669,N_17285,N_17354);
xor U17670 (N_17670,N_17470,N_17405);
nand U17671 (N_17671,N_17362,N_17255);
and U17672 (N_17672,N_17356,N_17363);
nand U17673 (N_17673,N_17335,N_17468);
nor U17674 (N_17674,N_17297,N_17407);
xnor U17675 (N_17675,N_17491,N_17474);
nor U17676 (N_17676,N_17408,N_17358);
or U17677 (N_17677,N_17254,N_17459);
xor U17678 (N_17678,N_17278,N_17326);
nand U17679 (N_17679,N_17323,N_17482);
or U17680 (N_17680,N_17475,N_17285);
nor U17681 (N_17681,N_17252,N_17256);
or U17682 (N_17682,N_17324,N_17345);
and U17683 (N_17683,N_17468,N_17318);
nand U17684 (N_17684,N_17414,N_17421);
and U17685 (N_17685,N_17440,N_17483);
or U17686 (N_17686,N_17348,N_17481);
nand U17687 (N_17687,N_17402,N_17454);
and U17688 (N_17688,N_17399,N_17491);
nor U17689 (N_17689,N_17314,N_17474);
nand U17690 (N_17690,N_17383,N_17260);
xor U17691 (N_17691,N_17309,N_17345);
or U17692 (N_17692,N_17289,N_17363);
and U17693 (N_17693,N_17334,N_17318);
or U17694 (N_17694,N_17317,N_17338);
or U17695 (N_17695,N_17298,N_17386);
or U17696 (N_17696,N_17369,N_17430);
xor U17697 (N_17697,N_17358,N_17286);
or U17698 (N_17698,N_17484,N_17353);
nand U17699 (N_17699,N_17444,N_17433);
xor U17700 (N_17700,N_17393,N_17389);
xor U17701 (N_17701,N_17369,N_17469);
xnor U17702 (N_17702,N_17333,N_17370);
nor U17703 (N_17703,N_17393,N_17361);
or U17704 (N_17704,N_17443,N_17374);
or U17705 (N_17705,N_17371,N_17254);
nor U17706 (N_17706,N_17334,N_17353);
and U17707 (N_17707,N_17271,N_17492);
and U17708 (N_17708,N_17252,N_17375);
xnor U17709 (N_17709,N_17260,N_17360);
nand U17710 (N_17710,N_17356,N_17402);
or U17711 (N_17711,N_17349,N_17378);
nand U17712 (N_17712,N_17283,N_17406);
nor U17713 (N_17713,N_17365,N_17281);
nor U17714 (N_17714,N_17259,N_17293);
and U17715 (N_17715,N_17393,N_17420);
and U17716 (N_17716,N_17293,N_17288);
xnor U17717 (N_17717,N_17368,N_17284);
or U17718 (N_17718,N_17402,N_17483);
nor U17719 (N_17719,N_17438,N_17374);
nor U17720 (N_17720,N_17428,N_17301);
nor U17721 (N_17721,N_17259,N_17487);
nand U17722 (N_17722,N_17379,N_17304);
or U17723 (N_17723,N_17345,N_17335);
or U17724 (N_17724,N_17423,N_17475);
or U17725 (N_17725,N_17273,N_17292);
nor U17726 (N_17726,N_17454,N_17445);
xnor U17727 (N_17727,N_17436,N_17456);
or U17728 (N_17728,N_17373,N_17309);
xnor U17729 (N_17729,N_17494,N_17394);
xnor U17730 (N_17730,N_17445,N_17494);
and U17731 (N_17731,N_17267,N_17283);
nor U17732 (N_17732,N_17434,N_17489);
or U17733 (N_17733,N_17360,N_17371);
and U17734 (N_17734,N_17448,N_17477);
xnor U17735 (N_17735,N_17253,N_17310);
and U17736 (N_17736,N_17416,N_17477);
nor U17737 (N_17737,N_17418,N_17320);
and U17738 (N_17738,N_17400,N_17406);
nor U17739 (N_17739,N_17348,N_17354);
xnor U17740 (N_17740,N_17280,N_17492);
or U17741 (N_17741,N_17472,N_17403);
nor U17742 (N_17742,N_17368,N_17455);
nor U17743 (N_17743,N_17295,N_17446);
nor U17744 (N_17744,N_17301,N_17364);
xor U17745 (N_17745,N_17361,N_17364);
nor U17746 (N_17746,N_17432,N_17286);
nand U17747 (N_17747,N_17316,N_17431);
and U17748 (N_17748,N_17417,N_17483);
and U17749 (N_17749,N_17406,N_17309);
and U17750 (N_17750,N_17611,N_17582);
and U17751 (N_17751,N_17558,N_17547);
nor U17752 (N_17752,N_17703,N_17520);
and U17753 (N_17753,N_17551,N_17503);
nand U17754 (N_17754,N_17726,N_17614);
nor U17755 (N_17755,N_17683,N_17584);
and U17756 (N_17756,N_17612,N_17524);
nand U17757 (N_17757,N_17549,N_17710);
and U17758 (N_17758,N_17579,N_17572);
or U17759 (N_17759,N_17660,N_17727);
or U17760 (N_17760,N_17533,N_17525);
and U17761 (N_17761,N_17637,N_17633);
or U17762 (N_17762,N_17597,N_17639);
xor U17763 (N_17763,N_17748,N_17634);
nand U17764 (N_17764,N_17737,N_17513);
nand U17765 (N_17765,N_17638,N_17643);
nand U17766 (N_17766,N_17546,N_17521);
and U17767 (N_17767,N_17655,N_17528);
or U17768 (N_17768,N_17535,N_17729);
nor U17769 (N_17769,N_17606,N_17539);
nand U17770 (N_17770,N_17702,N_17570);
xor U17771 (N_17771,N_17509,N_17661);
xnor U17772 (N_17772,N_17591,N_17502);
xnor U17773 (N_17773,N_17736,N_17515);
or U17774 (N_17774,N_17517,N_17730);
and U17775 (N_17775,N_17556,N_17742);
or U17776 (N_17776,N_17530,N_17615);
nor U17777 (N_17777,N_17552,N_17585);
nand U17778 (N_17778,N_17563,N_17649);
and U17779 (N_17779,N_17644,N_17571);
xor U17780 (N_17780,N_17733,N_17632);
or U17781 (N_17781,N_17577,N_17745);
xnor U17782 (N_17782,N_17642,N_17707);
or U17783 (N_17783,N_17668,N_17540);
or U17784 (N_17784,N_17523,N_17709);
nor U17785 (N_17785,N_17747,N_17657);
or U17786 (N_17786,N_17601,N_17522);
and U17787 (N_17787,N_17575,N_17687);
xor U17788 (N_17788,N_17731,N_17548);
or U17789 (N_17789,N_17629,N_17567);
xor U17790 (N_17790,N_17700,N_17659);
nand U17791 (N_17791,N_17718,N_17685);
or U17792 (N_17792,N_17721,N_17722);
xnor U17793 (N_17793,N_17593,N_17550);
or U17794 (N_17794,N_17555,N_17566);
nor U17795 (N_17795,N_17699,N_17746);
nor U17796 (N_17796,N_17623,N_17543);
nor U17797 (N_17797,N_17646,N_17663);
xnor U17798 (N_17798,N_17607,N_17568);
and U17799 (N_17799,N_17719,N_17538);
xnor U17800 (N_17800,N_17620,N_17672);
nor U17801 (N_17801,N_17507,N_17514);
xnor U17802 (N_17802,N_17595,N_17588);
nand U17803 (N_17803,N_17602,N_17676);
and U17804 (N_17804,N_17704,N_17576);
xnor U17805 (N_17805,N_17527,N_17616);
xnor U17806 (N_17806,N_17599,N_17664);
xor U17807 (N_17807,N_17689,N_17715);
and U17808 (N_17808,N_17670,N_17600);
nand U17809 (N_17809,N_17708,N_17675);
and U17810 (N_17810,N_17627,N_17603);
and U17811 (N_17811,N_17716,N_17744);
or U17812 (N_17812,N_17724,N_17504);
xnor U17813 (N_17813,N_17698,N_17741);
and U17814 (N_17814,N_17622,N_17723);
or U17815 (N_17815,N_17604,N_17658);
xor U17816 (N_17816,N_17749,N_17656);
nand U17817 (N_17817,N_17586,N_17506);
or U17818 (N_17818,N_17662,N_17587);
xnor U17819 (N_17819,N_17667,N_17743);
nor U17820 (N_17820,N_17684,N_17621);
nand U17821 (N_17821,N_17714,N_17650);
xor U17822 (N_17822,N_17681,N_17692);
xnor U17823 (N_17823,N_17605,N_17531);
and U17824 (N_17824,N_17677,N_17544);
xor U17825 (N_17825,N_17693,N_17564);
and U17826 (N_17826,N_17665,N_17711);
nand U17827 (N_17827,N_17580,N_17583);
nor U17828 (N_17828,N_17536,N_17694);
and U17829 (N_17829,N_17569,N_17574);
nor U17830 (N_17830,N_17688,N_17560);
nand U17831 (N_17831,N_17640,N_17508);
nor U17832 (N_17832,N_17512,N_17728);
xnor U17833 (N_17833,N_17613,N_17740);
and U17834 (N_17834,N_17636,N_17669);
nor U17835 (N_17835,N_17609,N_17701);
nand U17836 (N_17836,N_17618,N_17537);
xor U17837 (N_17837,N_17651,N_17635);
or U17838 (N_17838,N_17690,N_17581);
or U17839 (N_17839,N_17697,N_17559);
nand U17840 (N_17840,N_17619,N_17732);
and U17841 (N_17841,N_17691,N_17695);
and U17842 (N_17842,N_17501,N_17526);
and U17843 (N_17843,N_17565,N_17671);
and U17844 (N_17844,N_17519,N_17735);
and U17845 (N_17845,N_17545,N_17696);
or U17846 (N_17846,N_17712,N_17626);
nand U17847 (N_17847,N_17630,N_17518);
and U17848 (N_17848,N_17674,N_17541);
and U17849 (N_17849,N_17717,N_17720);
or U17850 (N_17850,N_17608,N_17678);
or U17851 (N_17851,N_17641,N_17589);
and U17852 (N_17852,N_17542,N_17554);
nand U17853 (N_17853,N_17534,N_17653);
or U17854 (N_17854,N_17673,N_17598);
and U17855 (N_17855,N_17738,N_17573);
xnor U17856 (N_17856,N_17592,N_17590);
nor U17857 (N_17857,N_17624,N_17578);
or U17858 (N_17858,N_17561,N_17617);
nor U17859 (N_17859,N_17510,N_17739);
or U17860 (N_17860,N_17645,N_17596);
or U17861 (N_17861,N_17725,N_17680);
nor U17862 (N_17862,N_17682,N_17631);
nor U17863 (N_17863,N_17706,N_17679);
nor U17864 (N_17864,N_17713,N_17505);
nand U17865 (N_17865,N_17654,N_17628);
or U17866 (N_17866,N_17500,N_17532);
and U17867 (N_17867,N_17562,N_17610);
nor U17868 (N_17868,N_17686,N_17648);
and U17869 (N_17869,N_17511,N_17553);
or U17870 (N_17870,N_17647,N_17734);
or U17871 (N_17871,N_17594,N_17516);
nand U17872 (N_17872,N_17652,N_17705);
or U17873 (N_17873,N_17666,N_17557);
or U17874 (N_17874,N_17529,N_17625);
xor U17875 (N_17875,N_17649,N_17588);
nand U17876 (N_17876,N_17503,N_17706);
xor U17877 (N_17877,N_17558,N_17500);
nand U17878 (N_17878,N_17724,N_17507);
or U17879 (N_17879,N_17542,N_17519);
and U17880 (N_17880,N_17622,N_17696);
nand U17881 (N_17881,N_17748,N_17741);
or U17882 (N_17882,N_17574,N_17502);
nor U17883 (N_17883,N_17715,N_17545);
xor U17884 (N_17884,N_17651,N_17539);
xor U17885 (N_17885,N_17572,N_17610);
nor U17886 (N_17886,N_17695,N_17697);
xor U17887 (N_17887,N_17519,N_17646);
xnor U17888 (N_17888,N_17649,N_17604);
nand U17889 (N_17889,N_17738,N_17641);
nand U17890 (N_17890,N_17544,N_17732);
and U17891 (N_17891,N_17548,N_17619);
and U17892 (N_17892,N_17654,N_17537);
nand U17893 (N_17893,N_17570,N_17546);
or U17894 (N_17894,N_17657,N_17553);
nand U17895 (N_17895,N_17650,N_17721);
and U17896 (N_17896,N_17697,N_17661);
nand U17897 (N_17897,N_17604,N_17532);
xnor U17898 (N_17898,N_17745,N_17540);
nand U17899 (N_17899,N_17672,N_17619);
nand U17900 (N_17900,N_17748,N_17717);
xnor U17901 (N_17901,N_17728,N_17576);
nor U17902 (N_17902,N_17679,N_17589);
and U17903 (N_17903,N_17593,N_17600);
xor U17904 (N_17904,N_17638,N_17535);
nand U17905 (N_17905,N_17635,N_17572);
xor U17906 (N_17906,N_17672,N_17623);
or U17907 (N_17907,N_17578,N_17744);
or U17908 (N_17908,N_17568,N_17524);
or U17909 (N_17909,N_17676,N_17612);
or U17910 (N_17910,N_17527,N_17717);
xnor U17911 (N_17911,N_17704,N_17671);
nand U17912 (N_17912,N_17519,N_17636);
or U17913 (N_17913,N_17600,N_17594);
or U17914 (N_17914,N_17633,N_17742);
and U17915 (N_17915,N_17684,N_17638);
and U17916 (N_17916,N_17747,N_17679);
or U17917 (N_17917,N_17678,N_17622);
or U17918 (N_17918,N_17610,N_17635);
xnor U17919 (N_17919,N_17652,N_17562);
or U17920 (N_17920,N_17647,N_17745);
nand U17921 (N_17921,N_17559,N_17746);
and U17922 (N_17922,N_17511,N_17599);
xnor U17923 (N_17923,N_17636,N_17557);
and U17924 (N_17924,N_17677,N_17723);
and U17925 (N_17925,N_17512,N_17635);
nor U17926 (N_17926,N_17660,N_17638);
and U17927 (N_17927,N_17535,N_17585);
nor U17928 (N_17928,N_17553,N_17701);
or U17929 (N_17929,N_17519,N_17716);
xor U17930 (N_17930,N_17721,N_17701);
and U17931 (N_17931,N_17660,N_17586);
or U17932 (N_17932,N_17690,N_17714);
and U17933 (N_17933,N_17592,N_17689);
nor U17934 (N_17934,N_17651,N_17652);
or U17935 (N_17935,N_17566,N_17553);
nand U17936 (N_17936,N_17519,N_17596);
nand U17937 (N_17937,N_17559,N_17641);
nand U17938 (N_17938,N_17622,N_17652);
or U17939 (N_17939,N_17737,N_17609);
nand U17940 (N_17940,N_17589,N_17681);
nand U17941 (N_17941,N_17520,N_17632);
and U17942 (N_17942,N_17596,N_17742);
xnor U17943 (N_17943,N_17647,N_17625);
nand U17944 (N_17944,N_17744,N_17634);
or U17945 (N_17945,N_17608,N_17729);
or U17946 (N_17946,N_17507,N_17650);
and U17947 (N_17947,N_17571,N_17725);
and U17948 (N_17948,N_17688,N_17554);
xor U17949 (N_17949,N_17644,N_17547);
nor U17950 (N_17950,N_17663,N_17588);
nor U17951 (N_17951,N_17573,N_17555);
xor U17952 (N_17952,N_17590,N_17584);
and U17953 (N_17953,N_17687,N_17697);
and U17954 (N_17954,N_17594,N_17734);
nor U17955 (N_17955,N_17601,N_17590);
nand U17956 (N_17956,N_17717,N_17590);
and U17957 (N_17957,N_17625,N_17561);
nand U17958 (N_17958,N_17595,N_17543);
nand U17959 (N_17959,N_17653,N_17527);
nor U17960 (N_17960,N_17680,N_17513);
and U17961 (N_17961,N_17611,N_17741);
nor U17962 (N_17962,N_17715,N_17680);
or U17963 (N_17963,N_17523,N_17568);
xnor U17964 (N_17964,N_17688,N_17632);
or U17965 (N_17965,N_17594,N_17672);
and U17966 (N_17966,N_17575,N_17603);
nor U17967 (N_17967,N_17552,N_17711);
and U17968 (N_17968,N_17736,N_17541);
nor U17969 (N_17969,N_17653,N_17747);
or U17970 (N_17970,N_17687,N_17618);
nand U17971 (N_17971,N_17517,N_17570);
and U17972 (N_17972,N_17612,N_17517);
xor U17973 (N_17973,N_17626,N_17749);
or U17974 (N_17974,N_17671,N_17723);
xnor U17975 (N_17975,N_17600,N_17609);
or U17976 (N_17976,N_17663,N_17630);
nand U17977 (N_17977,N_17538,N_17561);
and U17978 (N_17978,N_17508,N_17696);
or U17979 (N_17979,N_17564,N_17552);
and U17980 (N_17980,N_17685,N_17501);
nor U17981 (N_17981,N_17577,N_17550);
and U17982 (N_17982,N_17573,N_17673);
nand U17983 (N_17983,N_17703,N_17641);
nand U17984 (N_17984,N_17639,N_17675);
or U17985 (N_17985,N_17710,N_17565);
xor U17986 (N_17986,N_17568,N_17722);
and U17987 (N_17987,N_17651,N_17700);
xor U17988 (N_17988,N_17575,N_17565);
or U17989 (N_17989,N_17524,N_17648);
nand U17990 (N_17990,N_17744,N_17508);
xor U17991 (N_17991,N_17516,N_17714);
xnor U17992 (N_17992,N_17673,N_17634);
and U17993 (N_17993,N_17660,N_17503);
xnor U17994 (N_17994,N_17594,N_17741);
nand U17995 (N_17995,N_17528,N_17584);
and U17996 (N_17996,N_17667,N_17610);
nor U17997 (N_17997,N_17740,N_17737);
nor U17998 (N_17998,N_17743,N_17531);
or U17999 (N_17999,N_17634,N_17521);
and U18000 (N_18000,N_17893,N_17939);
xnor U18001 (N_18001,N_17794,N_17921);
xnor U18002 (N_18002,N_17813,N_17889);
and U18003 (N_18003,N_17752,N_17999);
nor U18004 (N_18004,N_17928,N_17830);
and U18005 (N_18005,N_17766,N_17777);
and U18006 (N_18006,N_17877,N_17887);
and U18007 (N_18007,N_17832,N_17858);
nor U18008 (N_18008,N_17817,N_17849);
or U18009 (N_18009,N_17979,N_17776);
and U18010 (N_18010,N_17751,N_17845);
or U18011 (N_18011,N_17764,N_17905);
or U18012 (N_18012,N_17774,N_17988);
and U18013 (N_18013,N_17837,N_17855);
xor U18014 (N_18014,N_17750,N_17985);
or U18015 (N_18015,N_17891,N_17758);
xor U18016 (N_18016,N_17782,N_17789);
and U18017 (N_18017,N_17872,N_17866);
xnor U18018 (N_18018,N_17952,N_17983);
or U18019 (N_18019,N_17756,N_17820);
or U18020 (N_18020,N_17904,N_17807);
and U18021 (N_18021,N_17827,N_17951);
nand U18022 (N_18022,N_17969,N_17907);
xnor U18023 (N_18023,N_17883,N_17784);
and U18024 (N_18024,N_17990,N_17882);
xnor U18025 (N_18025,N_17765,N_17942);
xnor U18026 (N_18026,N_17790,N_17851);
and U18027 (N_18027,N_17971,N_17930);
nor U18028 (N_18028,N_17839,N_17792);
nor U18029 (N_18029,N_17918,N_17812);
nor U18030 (N_18030,N_17779,N_17909);
xor U18031 (N_18031,N_17811,N_17825);
and U18032 (N_18032,N_17838,N_17800);
xor U18033 (N_18033,N_17967,N_17911);
or U18034 (N_18034,N_17934,N_17836);
and U18035 (N_18035,N_17834,N_17910);
and U18036 (N_18036,N_17932,N_17901);
nor U18037 (N_18037,N_17981,N_17862);
xor U18038 (N_18038,N_17968,N_17857);
or U18039 (N_18039,N_17998,N_17846);
xnor U18040 (N_18040,N_17821,N_17896);
or U18041 (N_18041,N_17785,N_17874);
nor U18042 (N_18042,N_17991,N_17864);
xnor U18043 (N_18043,N_17875,N_17980);
or U18044 (N_18044,N_17850,N_17987);
nand U18045 (N_18045,N_17860,N_17953);
nand U18046 (N_18046,N_17814,N_17954);
xor U18047 (N_18047,N_17994,N_17895);
and U18048 (N_18048,N_17788,N_17960);
nand U18049 (N_18049,N_17878,N_17898);
or U18050 (N_18050,N_17966,N_17879);
xnor U18051 (N_18051,N_17854,N_17955);
or U18052 (N_18052,N_17767,N_17768);
and U18053 (N_18053,N_17859,N_17974);
or U18054 (N_18054,N_17970,N_17945);
xnor U18055 (N_18055,N_17853,N_17925);
or U18056 (N_18056,N_17977,N_17780);
xnor U18057 (N_18057,N_17835,N_17936);
and U18058 (N_18058,N_17848,N_17871);
and U18059 (N_18059,N_17831,N_17926);
xor U18060 (N_18060,N_17840,N_17947);
xor U18061 (N_18061,N_17941,N_17783);
or U18062 (N_18062,N_17885,N_17829);
and U18063 (N_18063,N_17982,N_17989);
xor U18064 (N_18064,N_17797,N_17841);
nor U18065 (N_18065,N_17861,N_17852);
or U18066 (N_18066,N_17822,N_17931);
nand U18067 (N_18067,N_17903,N_17880);
nor U18068 (N_18068,N_17972,N_17769);
and U18069 (N_18069,N_17916,N_17856);
and U18070 (N_18070,N_17787,N_17844);
and U18071 (N_18071,N_17973,N_17781);
nor U18072 (N_18072,N_17757,N_17847);
nand U18073 (N_18073,N_17922,N_17763);
and U18074 (N_18074,N_17935,N_17770);
or U18075 (N_18075,N_17753,N_17876);
or U18076 (N_18076,N_17957,N_17808);
and U18077 (N_18077,N_17992,N_17984);
nand U18078 (N_18078,N_17863,N_17892);
and U18079 (N_18079,N_17773,N_17819);
and U18080 (N_18080,N_17826,N_17908);
nand U18081 (N_18081,N_17943,N_17997);
nor U18082 (N_18082,N_17755,N_17786);
nor U18083 (N_18083,N_17920,N_17940);
or U18084 (N_18084,N_17965,N_17886);
nor U18085 (N_18085,N_17890,N_17865);
xnor U18086 (N_18086,N_17917,N_17805);
xnor U18087 (N_18087,N_17978,N_17796);
nand U18088 (N_18088,N_17995,N_17843);
xnor U18089 (N_18089,N_17937,N_17906);
nor U18090 (N_18090,N_17801,N_17806);
nand U18091 (N_18091,N_17964,N_17810);
or U18092 (N_18092,N_17944,N_17950);
nor U18093 (N_18093,N_17772,N_17828);
xnor U18094 (N_18094,N_17924,N_17815);
or U18095 (N_18095,N_17833,N_17760);
nand U18096 (N_18096,N_17884,N_17946);
nand U18097 (N_18097,N_17959,N_17762);
or U18098 (N_18098,N_17949,N_17956);
xor U18099 (N_18099,N_17888,N_17993);
and U18100 (N_18100,N_17894,N_17919);
nand U18101 (N_18101,N_17902,N_17799);
and U18102 (N_18102,N_17938,N_17816);
and U18103 (N_18103,N_17986,N_17996);
or U18104 (N_18104,N_17912,N_17899);
nand U18105 (N_18105,N_17754,N_17870);
nand U18106 (N_18106,N_17881,N_17927);
or U18107 (N_18107,N_17791,N_17868);
or U18108 (N_18108,N_17823,N_17867);
nor U18109 (N_18109,N_17775,N_17869);
and U18110 (N_18110,N_17793,N_17961);
nand U18111 (N_18111,N_17933,N_17900);
nor U18112 (N_18112,N_17958,N_17923);
and U18113 (N_18113,N_17771,N_17976);
nor U18114 (N_18114,N_17804,N_17929);
nor U18115 (N_18115,N_17913,N_17798);
and U18116 (N_18116,N_17778,N_17842);
xnor U18117 (N_18117,N_17873,N_17759);
nor U18118 (N_18118,N_17795,N_17761);
nand U18119 (N_18119,N_17948,N_17963);
nor U18120 (N_18120,N_17962,N_17802);
nor U18121 (N_18121,N_17975,N_17803);
nand U18122 (N_18122,N_17915,N_17914);
nor U18123 (N_18123,N_17824,N_17809);
nand U18124 (N_18124,N_17897,N_17818);
nand U18125 (N_18125,N_17816,N_17915);
nor U18126 (N_18126,N_17899,N_17930);
nor U18127 (N_18127,N_17808,N_17861);
xnor U18128 (N_18128,N_17821,N_17967);
and U18129 (N_18129,N_17928,N_17941);
nand U18130 (N_18130,N_17963,N_17902);
nand U18131 (N_18131,N_17802,N_17966);
or U18132 (N_18132,N_17896,N_17863);
xor U18133 (N_18133,N_17840,N_17917);
xnor U18134 (N_18134,N_17795,N_17862);
nor U18135 (N_18135,N_17902,N_17995);
xor U18136 (N_18136,N_17998,N_17884);
and U18137 (N_18137,N_17911,N_17879);
xor U18138 (N_18138,N_17852,N_17958);
or U18139 (N_18139,N_17957,N_17879);
nor U18140 (N_18140,N_17815,N_17978);
and U18141 (N_18141,N_17918,N_17755);
or U18142 (N_18142,N_17824,N_17960);
xor U18143 (N_18143,N_17952,N_17823);
or U18144 (N_18144,N_17924,N_17796);
and U18145 (N_18145,N_17973,N_17875);
xnor U18146 (N_18146,N_17755,N_17754);
nor U18147 (N_18147,N_17974,N_17828);
nor U18148 (N_18148,N_17954,N_17820);
and U18149 (N_18149,N_17940,N_17838);
nor U18150 (N_18150,N_17994,N_17843);
nand U18151 (N_18151,N_17930,N_17986);
nand U18152 (N_18152,N_17788,N_17768);
or U18153 (N_18153,N_17962,N_17898);
xnor U18154 (N_18154,N_17850,N_17926);
xnor U18155 (N_18155,N_17827,N_17835);
nand U18156 (N_18156,N_17933,N_17952);
nand U18157 (N_18157,N_17920,N_17803);
nand U18158 (N_18158,N_17988,N_17799);
nor U18159 (N_18159,N_17913,N_17891);
xor U18160 (N_18160,N_17848,N_17886);
and U18161 (N_18161,N_17982,N_17875);
xnor U18162 (N_18162,N_17869,N_17778);
nand U18163 (N_18163,N_17879,N_17788);
or U18164 (N_18164,N_17781,N_17868);
and U18165 (N_18165,N_17829,N_17843);
and U18166 (N_18166,N_17961,N_17939);
and U18167 (N_18167,N_17821,N_17992);
xor U18168 (N_18168,N_17859,N_17908);
nor U18169 (N_18169,N_17796,N_17789);
and U18170 (N_18170,N_17858,N_17932);
xor U18171 (N_18171,N_17856,N_17759);
nand U18172 (N_18172,N_17830,N_17867);
and U18173 (N_18173,N_17994,N_17877);
nor U18174 (N_18174,N_17883,N_17911);
or U18175 (N_18175,N_17908,N_17906);
nor U18176 (N_18176,N_17784,N_17858);
or U18177 (N_18177,N_17928,N_17773);
nand U18178 (N_18178,N_17914,N_17801);
xnor U18179 (N_18179,N_17998,N_17978);
nand U18180 (N_18180,N_17759,N_17774);
nor U18181 (N_18181,N_17999,N_17849);
or U18182 (N_18182,N_17833,N_17828);
xnor U18183 (N_18183,N_17987,N_17886);
xnor U18184 (N_18184,N_17904,N_17968);
xor U18185 (N_18185,N_17752,N_17957);
nand U18186 (N_18186,N_17824,N_17766);
nor U18187 (N_18187,N_17831,N_17836);
and U18188 (N_18188,N_17917,N_17909);
nand U18189 (N_18189,N_17886,N_17876);
nand U18190 (N_18190,N_17791,N_17917);
nor U18191 (N_18191,N_17830,N_17943);
and U18192 (N_18192,N_17758,N_17766);
nor U18193 (N_18193,N_17913,N_17980);
and U18194 (N_18194,N_17904,N_17844);
xnor U18195 (N_18195,N_17874,N_17980);
xor U18196 (N_18196,N_17898,N_17795);
or U18197 (N_18197,N_17793,N_17791);
nor U18198 (N_18198,N_17901,N_17974);
xor U18199 (N_18199,N_17826,N_17970);
and U18200 (N_18200,N_17794,N_17912);
xnor U18201 (N_18201,N_17782,N_17962);
and U18202 (N_18202,N_17847,N_17884);
nor U18203 (N_18203,N_17860,N_17954);
xnor U18204 (N_18204,N_17955,N_17998);
xor U18205 (N_18205,N_17804,N_17889);
nand U18206 (N_18206,N_17939,N_17925);
nand U18207 (N_18207,N_17910,N_17821);
nor U18208 (N_18208,N_17781,N_17931);
and U18209 (N_18209,N_17928,N_17754);
and U18210 (N_18210,N_17953,N_17980);
nand U18211 (N_18211,N_17810,N_17817);
and U18212 (N_18212,N_17968,N_17789);
nand U18213 (N_18213,N_17869,N_17982);
nor U18214 (N_18214,N_17857,N_17986);
nor U18215 (N_18215,N_17888,N_17951);
nor U18216 (N_18216,N_17963,N_17872);
xnor U18217 (N_18217,N_17964,N_17989);
nor U18218 (N_18218,N_17948,N_17959);
xor U18219 (N_18219,N_17848,N_17790);
nand U18220 (N_18220,N_17942,N_17799);
or U18221 (N_18221,N_17876,N_17918);
xor U18222 (N_18222,N_17765,N_17962);
or U18223 (N_18223,N_17935,N_17936);
xor U18224 (N_18224,N_17894,N_17985);
xnor U18225 (N_18225,N_17949,N_17878);
xnor U18226 (N_18226,N_17809,N_17836);
and U18227 (N_18227,N_17781,N_17915);
or U18228 (N_18228,N_17805,N_17892);
nand U18229 (N_18229,N_17968,N_17753);
nand U18230 (N_18230,N_17961,N_17872);
or U18231 (N_18231,N_17969,N_17955);
or U18232 (N_18232,N_17754,N_17977);
nor U18233 (N_18233,N_17795,N_17906);
xnor U18234 (N_18234,N_17847,N_17762);
or U18235 (N_18235,N_17963,N_17938);
and U18236 (N_18236,N_17821,N_17829);
and U18237 (N_18237,N_17817,N_17876);
xnor U18238 (N_18238,N_17913,N_17835);
xor U18239 (N_18239,N_17814,N_17762);
and U18240 (N_18240,N_17810,N_17970);
xor U18241 (N_18241,N_17769,N_17999);
and U18242 (N_18242,N_17794,N_17943);
nand U18243 (N_18243,N_17816,N_17881);
or U18244 (N_18244,N_17867,N_17841);
xnor U18245 (N_18245,N_17893,N_17755);
nand U18246 (N_18246,N_17975,N_17945);
and U18247 (N_18247,N_17993,N_17835);
nand U18248 (N_18248,N_17997,N_17877);
xor U18249 (N_18249,N_17913,N_17832);
or U18250 (N_18250,N_18043,N_18228);
nor U18251 (N_18251,N_18088,N_18177);
nor U18252 (N_18252,N_18089,N_18192);
and U18253 (N_18253,N_18005,N_18006);
or U18254 (N_18254,N_18144,N_18174);
nor U18255 (N_18255,N_18167,N_18029);
xnor U18256 (N_18256,N_18063,N_18048);
nor U18257 (N_18257,N_18133,N_18092);
nand U18258 (N_18258,N_18171,N_18212);
nor U18259 (N_18259,N_18095,N_18070);
and U18260 (N_18260,N_18002,N_18195);
or U18261 (N_18261,N_18200,N_18180);
xor U18262 (N_18262,N_18113,N_18033);
and U18263 (N_18263,N_18050,N_18231);
and U18264 (N_18264,N_18016,N_18163);
or U18265 (N_18265,N_18205,N_18120);
xnor U18266 (N_18266,N_18001,N_18085);
xnor U18267 (N_18267,N_18238,N_18248);
or U18268 (N_18268,N_18111,N_18143);
and U18269 (N_18269,N_18162,N_18196);
nor U18270 (N_18270,N_18184,N_18225);
nor U18271 (N_18271,N_18181,N_18012);
and U18272 (N_18272,N_18026,N_18216);
or U18273 (N_18273,N_18169,N_18185);
nand U18274 (N_18274,N_18054,N_18104);
xor U18275 (N_18275,N_18037,N_18229);
xnor U18276 (N_18276,N_18160,N_18064);
and U18277 (N_18277,N_18081,N_18051);
nor U18278 (N_18278,N_18135,N_18204);
or U18279 (N_18279,N_18145,N_18115);
and U18280 (N_18280,N_18208,N_18147);
or U18281 (N_18281,N_18096,N_18217);
nor U18282 (N_18282,N_18125,N_18084);
and U18283 (N_18283,N_18189,N_18197);
and U18284 (N_18284,N_18067,N_18232);
or U18285 (N_18285,N_18211,N_18102);
and U18286 (N_18286,N_18236,N_18045);
and U18287 (N_18287,N_18154,N_18061);
and U18288 (N_18288,N_18039,N_18047);
and U18289 (N_18289,N_18224,N_18024);
nand U18290 (N_18290,N_18086,N_18017);
nor U18291 (N_18291,N_18237,N_18114);
nor U18292 (N_18292,N_18166,N_18244);
nor U18293 (N_18293,N_18093,N_18025);
or U18294 (N_18294,N_18027,N_18003);
nand U18295 (N_18295,N_18191,N_18100);
nand U18296 (N_18296,N_18159,N_18056);
nand U18297 (N_18297,N_18032,N_18087);
or U18298 (N_18298,N_18082,N_18157);
or U18299 (N_18299,N_18140,N_18128);
nand U18300 (N_18300,N_18146,N_18233);
nor U18301 (N_18301,N_18198,N_18069);
xnor U18302 (N_18302,N_18053,N_18090);
nor U18303 (N_18303,N_18249,N_18235);
or U18304 (N_18304,N_18239,N_18020);
nand U18305 (N_18305,N_18116,N_18179);
nor U18306 (N_18306,N_18246,N_18134);
or U18307 (N_18307,N_18187,N_18164);
xor U18308 (N_18308,N_18172,N_18141);
or U18309 (N_18309,N_18117,N_18074);
and U18310 (N_18310,N_18161,N_18188);
nand U18311 (N_18311,N_18156,N_18023);
nand U18312 (N_18312,N_18108,N_18209);
nor U18313 (N_18313,N_18126,N_18097);
nand U18314 (N_18314,N_18136,N_18046);
xor U18315 (N_18315,N_18013,N_18122);
nand U18316 (N_18316,N_18098,N_18007);
nor U18317 (N_18317,N_18077,N_18094);
and U18318 (N_18318,N_18139,N_18057);
nor U18319 (N_18319,N_18014,N_18130);
or U18320 (N_18320,N_18215,N_18036);
or U18321 (N_18321,N_18132,N_18121);
and U18322 (N_18322,N_18153,N_18137);
nor U18323 (N_18323,N_18011,N_18071);
nor U18324 (N_18324,N_18219,N_18178);
nand U18325 (N_18325,N_18038,N_18091);
xnor U18326 (N_18326,N_18044,N_18222);
nor U18327 (N_18327,N_18151,N_18107);
xnor U18328 (N_18328,N_18127,N_18176);
and U18329 (N_18329,N_18138,N_18103);
xor U18330 (N_18330,N_18221,N_18123);
nand U18331 (N_18331,N_18105,N_18042);
nand U18332 (N_18332,N_18101,N_18247);
nand U18333 (N_18333,N_18009,N_18000);
nor U18334 (N_18334,N_18186,N_18058);
and U18335 (N_18335,N_18099,N_18119);
nor U18336 (N_18336,N_18110,N_18004);
and U18337 (N_18337,N_18008,N_18041);
xor U18338 (N_18338,N_18234,N_18214);
and U18339 (N_18339,N_18220,N_18124);
or U18340 (N_18340,N_18242,N_18201);
xnor U18341 (N_18341,N_18106,N_18158);
xnor U18342 (N_18342,N_18059,N_18052);
or U18343 (N_18343,N_18018,N_18118);
xor U18344 (N_18344,N_18079,N_18165);
nor U18345 (N_18345,N_18072,N_18223);
nand U18346 (N_18346,N_18068,N_18076);
or U18347 (N_18347,N_18173,N_18022);
nand U18348 (N_18348,N_18170,N_18240);
and U18349 (N_18349,N_18019,N_18112);
and U18350 (N_18350,N_18131,N_18021);
nor U18351 (N_18351,N_18035,N_18183);
nand U18352 (N_18352,N_18075,N_18028);
and U18353 (N_18353,N_18065,N_18227);
and U18354 (N_18354,N_18073,N_18010);
nand U18355 (N_18355,N_18243,N_18210);
nand U18356 (N_18356,N_18129,N_18207);
or U18357 (N_18357,N_18109,N_18245);
or U18358 (N_18358,N_18241,N_18193);
or U18359 (N_18359,N_18203,N_18152);
nor U18360 (N_18360,N_18066,N_18040);
or U18361 (N_18361,N_18080,N_18206);
or U18362 (N_18362,N_18060,N_18150);
or U18363 (N_18363,N_18168,N_18034);
nor U18364 (N_18364,N_18175,N_18202);
and U18365 (N_18365,N_18218,N_18078);
and U18366 (N_18366,N_18015,N_18148);
and U18367 (N_18367,N_18062,N_18049);
xor U18368 (N_18368,N_18190,N_18194);
and U18369 (N_18369,N_18030,N_18149);
or U18370 (N_18370,N_18142,N_18226);
and U18371 (N_18371,N_18055,N_18182);
xor U18372 (N_18372,N_18155,N_18213);
nand U18373 (N_18373,N_18199,N_18031);
nor U18374 (N_18374,N_18230,N_18083);
and U18375 (N_18375,N_18173,N_18202);
and U18376 (N_18376,N_18003,N_18102);
xor U18377 (N_18377,N_18039,N_18049);
nand U18378 (N_18378,N_18144,N_18176);
or U18379 (N_18379,N_18089,N_18199);
and U18380 (N_18380,N_18208,N_18037);
xor U18381 (N_18381,N_18231,N_18200);
nor U18382 (N_18382,N_18186,N_18090);
nor U18383 (N_18383,N_18066,N_18221);
xor U18384 (N_18384,N_18182,N_18218);
nor U18385 (N_18385,N_18200,N_18085);
nor U18386 (N_18386,N_18155,N_18135);
xor U18387 (N_18387,N_18229,N_18216);
nand U18388 (N_18388,N_18163,N_18112);
xnor U18389 (N_18389,N_18226,N_18046);
nor U18390 (N_18390,N_18058,N_18110);
nand U18391 (N_18391,N_18008,N_18223);
nand U18392 (N_18392,N_18242,N_18088);
or U18393 (N_18393,N_18203,N_18048);
nor U18394 (N_18394,N_18056,N_18120);
nand U18395 (N_18395,N_18225,N_18204);
or U18396 (N_18396,N_18025,N_18189);
and U18397 (N_18397,N_18117,N_18243);
or U18398 (N_18398,N_18181,N_18090);
xor U18399 (N_18399,N_18015,N_18157);
xor U18400 (N_18400,N_18141,N_18223);
nor U18401 (N_18401,N_18039,N_18036);
nand U18402 (N_18402,N_18197,N_18069);
xor U18403 (N_18403,N_18198,N_18205);
and U18404 (N_18404,N_18125,N_18135);
nand U18405 (N_18405,N_18174,N_18145);
or U18406 (N_18406,N_18139,N_18175);
nor U18407 (N_18407,N_18053,N_18028);
and U18408 (N_18408,N_18029,N_18086);
xor U18409 (N_18409,N_18095,N_18071);
or U18410 (N_18410,N_18120,N_18103);
xnor U18411 (N_18411,N_18029,N_18105);
or U18412 (N_18412,N_18029,N_18133);
nor U18413 (N_18413,N_18027,N_18124);
or U18414 (N_18414,N_18100,N_18043);
and U18415 (N_18415,N_18098,N_18092);
xor U18416 (N_18416,N_18121,N_18149);
or U18417 (N_18417,N_18058,N_18000);
and U18418 (N_18418,N_18214,N_18116);
xor U18419 (N_18419,N_18029,N_18090);
nand U18420 (N_18420,N_18169,N_18179);
nor U18421 (N_18421,N_18113,N_18025);
xnor U18422 (N_18422,N_18175,N_18227);
nand U18423 (N_18423,N_18163,N_18126);
nor U18424 (N_18424,N_18138,N_18142);
and U18425 (N_18425,N_18090,N_18202);
and U18426 (N_18426,N_18232,N_18140);
xor U18427 (N_18427,N_18225,N_18062);
nor U18428 (N_18428,N_18214,N_18015);
xor U18429 (N_18429,N_18125,N_18137);
and U18430 (N_18430,N_18183,N_18124);
or U18431 (N_18431,N_18076,N_18041);
and U18432 (N_18432,N_18003,N_18038);
nor U18433 (N_18433,N_18005,N_18229);
and U18434 (N_18434,N_18061,N_18131);
xnor U18435 (N_18435,N_18043,N_18056);
nand U18436 (N_18436,N_18020,N_18128);
nand U18437 (N_18437,N_18057,N_18149);
and U18438 (N_18438,N_18166,N_18101);
and U18439 (N_18439,N_18041,N_18038);
nor U18440 (N_18440,N_18176,N_18142);
and U18441 (N_18441,N_18055,N_18227);
nand U18442 (N_18442,N_18178,N_18046);
or U18443 (N_18443,N_18013,N_18016);
xnor U18444 (N_18444,N_18233,N_18105);
nand U18445 (N_18445,N_18212,N_18044);
nand U18446 (N_18446,N_18132,N_18056);
nor U18447 (N_18447,N_18145,N_18248);
and U18448 (N_18448,N_18228,N_18077);
nor U18449 (N_18449,N_18172,N_18023);
xor U18450 (N_18450,N_18078,N_18176);
xor U18451 (N_18451,N_18139,N_18122);
xor U18452 (N_18452,N_18057,N_18077);
or U18453 (N_18453,N_18175,N_18200);
nand U18454 (N_18454,N_18072,N_18245);
nor U18455 (N_18455,N_18173,N_18034);
or U18456 (N_18456,N_18239,N_18043);
or U18457 (N_18457,N_18182,N_18044);
and U18458 (N_18458,N_18019,N_18014);
and U18459 (N_18459,N_18052,N_18168);
nand U18460 (N_18460,N_18046,N_18223);
and U18461 (N_18461,N_18187,N_18000);
and U18462 (N_18462,N_18040,N_18184);
nand U18463 (N_18463,N_18052,N_18211);
nor U18464 (N_18464,N_18096,N_18060);
nor U18465 (N_18465,N_18002,N_18109);
xor U18466 (N_18466,N_18007,N_18244);
xor U18467 (N_18467,N_18242,N_18034);
or U18468 (N_18468,N_18147,N_18015);
nor U18469 (N_18469,N_18066,N_18236);
xnor U18470 (N_18470,N_18227,N_18177);
or U18471 (N_18471,N_18200,N_18058);
nand U18472 (N_18472,N_18229,N_18048);
xnor U18473 (N_18473,N_18117,N_18087);
and U18474 (N_18474,N_18248,N_18010);
nor U18475 (N_18475,N_18241,N_18019);
or U18476 (N_18476,N_18209,N_18058);
nor U18477 (N_18477,N_18085,N_18233);
and U18478 (N_18478,N_18234,N_18005);
xnor U18479 (N_18479,N_18190,N_18034);
or U18480 (N_18480,N_18188,N_18043);
nor U18481 (N_18481,N_18183,N_18205);
xor U18482 (N_18482,N_18246,N_18171);
or U18483 (N_18483,N_18120,N_18088);
xor U18484 (N_18484,N_18152,N_18089);
nand U18485 (N_18485,N_18212,N_18180);
xnor U18486 (N_18486,N_18246,N_18208);
or U18487 (N_18487,N_18183,N_18143);
or U18488 (N_18488,N_18051,N_18102);
and U18489 (N_18489,N_18182,N_18001);
nand U18490 (N_18490,N_18101,N_18230);
nor U18491 (N_18491,N_18029,N_18062);
xnor U18492 (N_18492,N_18220,N_18040);
or U18493 (N_18493,N_18185,N_18091);
and U18494 (N_18494,N_18223,N_18099);
xor U18495 (N_18495,N_18031,N_18135);
nor U18496 (N_18496,N_18001,N_18185);
nor U18497 (N_18497,N_18245,N_18002);
and U18498 (N_18498,N_18013,N_18203);
nand U18499 (N_18499,N_18071,N_18171);
or U18500 (N_18500,N_18294,N_18492);
or U18501 (N_18501,N_18389,N_18252);
and U18502 (N_18502,N_18458,N_18431);
or U18503 (N_18503,N_18330,N_18289);
xor U18504 (N_18504,N_18425,N_18280);
xnor U18505 (N_18505,N_18450,N_18446);
or U18506 (N_18506,N_18263,N_18408);
nand U18507 (N_18507,N_18435,N_18442);
or U18508 (N_18508,N_18430,N_18296);
or U18509 (N_18509,N_18368,N_18268);
nor U18510 (N_18510,N_18281,N_18436);
or U18511 (N_18511,N_18316,N_18467);
and U18512 (N_18512,N_18272,N_18270);
nand U18513 (N_18513,N_18299,N_18343);
and U18514 (N_18514,N_18312,N_18424);
or U18515 (N_18515,N_18279,N_18264);
nor U18516 (N_18516,N_18367,N_18336);
and U18517 (N_18517,N_18423,N_18354);
or U18518 (N_18518,N_18426,N_18421);
and U18519 (N_18519,N_18455,N_18388);
or U18520 (N_18520,N_18490,N_18329);
or U18521 (N_18521,N_18398,N_18314);
or U18522 (N_18522,N_18303,N_18325);
nor U18523 (N_18523,N_18440,N_18350);
nor U18524 (N_18524,N_18444,N_18499);
xnor U18525 (N_18525,N_18413,N_18478);
nor U18526 (N_18526,N_18382,N_18456);
nand U18527 (N_18527,N_18394,N_18432);
nor U18528 (N_18528,N_18461,N_18441);
or U18529 (N_18529,N_18472,N_18332);
nand U18530 (N_18530,N_18286,N_18291);
nor U18531 (N_18531,N_18342,N_18417);
nor U18532 (N_18532,N_18352,N_18341);
or U18533 (N_18533,N_18459,N_18292);
xor U18534 (N_18534,N_18403,N_18428);
nand U18535 (N_18535,N_18414,N_18273);
xor U18536 (N_18536,N_18322,N_18290);
or U18537 (N_18537,N_18372,N_18400);
or U18538 (N_18538,N_18357,N_18380);
and U18539 (N_18539,N_18462,N_18359);
and U18540 (N_18540,N_18257,N_18392);
xnor U18541 (N_18541,N_18419,N_18447);
nor U18542 (N_18542,N_18420,N_18277);
xor U18543 (N_18543,N_18401,N_18407);
and U18544 (N_18544,N_18338,N_18384);
or U18545 (N_18545,N_18259,N_18267);
nand U18546 (N_18546,N_18463,N_18269);
and U18547 (N_18547,N_18410,N_18363);
nor U18548 (N_18548,N_18437,N_18346);
or U18549 (N_18549,N_18295,N_18283);
nand U18550 (N_18550,N_18261,N_18371);
nor U18551 (N_18551,N_18433,N_18323);
nand U18552 (N_18552,N_18351,N_18487);
nor U18553 (N_18553,N_18497,N_18297);
nor U18554 (N_18554,N_18443,N_18493);
xnor U18555 (N_18555,N_18376,N_18300);
and U18556 (N_18556,N_18474,N_18434);
nand U18557 (N_18557,N_18482,N_18310);
nor U18558 (N_18558,N_18355,N_18457);
or U18559 (N_18559,N_18370,N_18360);
nand U18560 (N_18560,N_18362,N_18464);
nand U18561 (N_18561,N_18475,N_18375);
or U18562 (N_18562,N_18439,N_18427);
nor U18563 (N_18563,N_18485,N_18311);
xor U18564 (N_18564,N_18483,N_18466);
nand U18565 (N_18565,N_18397,N_18258);
or U18566 (N_18566,N_18344,N_18302);
or U18567 (N_18567,N_18307,N_18345);
xnor U18568 (N_18568,N_18275,N_18491);
and U18569 (N_18569,N_18313,N_18395);
nor U18570 (N_18570,N_18284,N_18469);
and U18571 (N_18571,N_18470,N_18326);
nand U18572 (N_18572,N_18301,N_18481);
nor U18573 (N_18573,N_18324,N_18495);
nand U18574 (N_18574,N_18361,N_18452);
xnor U18575 (N_18575,N_18287,N_18364);
or U18576 (N_18576,N_18451,N_18253);
xnor U18577 (N_18577,N_18429,N_18448);
nor U18578 (N_18578,N_18406,N_18356);
or U18579 (N_18579,N_18282,N_18468);
nand U18580 (N_18580,N_18396,N_18318);
and U18581 (N_18581,N_18304,N_18305);
and U18582 (N_18582,N_18339,N_18373);
and U18583 (N_18583,N_18489,N_18480);
nand U18584 (N_18584,N_18473,N_18479);
nand U18585 (N_18585,N_18349,N_18317);
xor U18586 (N_18586,N_18404,N_18254);
nor U18587 (N_18587,N_18265,N_18320);
nor U18588 (N_18588,N_18471,N_18327);
and U18589 (N_18589,N_18315,N_18422);
and U18590 (N_18590,N_18379,N_18353);
nand U18591 (N_18591,N_18337,N_18366);
or U18592 (N_18592,N_18331,N_18328);
nor U18593 (N_18593,N_18308,N_18465);
or U18594 (N_18594,N_18486,N_18271);
or U18595 (N_18595,N_18365,N_18293);
xnor U18596 (N_18596,N_18276,N_18309);
or U18597 (N_18597,N_18498,N_18477);
and U18598 (N_18598,N_18333,N_18399);
and U18599 (N_18599,N_18418,N_18262);
nor U18600 (N_18600,N_18386,N_18496);
or U18601 (N_18601,N_18393,N_18484);
nand U18602 (N_18602,N_18385,N_18369);
nor U18603 (N_18603,N_18391,N_18383);
xor U18604 (N_18604,N_18460,N_18378);
xor U18605 (N_18605,N_18340,N_18319);
and U18606 (N_18606,N_18347,N_18381);
xnor U18607 (N_18607,N_18390,N_18488);
xor U18608 (N_18608,N_18377,N_18476);
nand U18609 (N_18609,N_18494,N_18453);
xor U18610 (N_18610,N_18405,N_18415);
nand U18611 (N_18611,N_18278,N_18285);
nand U18612 (N_18612,N_18266,N_18260);
nor U18613 (N_18613,N_18411,N_18412);
xnor U18614 (N_18614,N_18306,N_18416);
nand U18615 (N_18615,N_18454,N_18409);
and U18616 (N_18616,N_18358,N_18256);
nand U18617 (N_18617,N_18250,N_18449);
nand U18618 (N_18618,N_18288,N_18402);
xor U18619 (N_18619,N_18251,N_18348);
and U18620 (N_18620,N_18298,N_18374);
nand U18621 (N_18621,N_18255,N_18445);
and U18622 (N_18622,N_18321,N_18335);
and U18623 (N_18623,N_18274,N_18387);
nor U18624 (N_18624,N_18334,N_18438);
or U18625 (N_18625,N_18291,N_18264);
nor U18626 (N_18626,N_18383,N_18319);
or U18627 (N_18627,N_18475,N_18418);
and U18628 (N_18628,N_18288,N_18357);
and U18629 (N_18629,N_18479,N_18360);
and U18630 (N_18630,N_18410,N_18470);
nand U18631 (N_18631,N_18372,N_18475);
nor U18632 (N_18632,N_18395,N_18440);
or U18633 (N_18633,N_18383,N_18429);
nand U18634 (N_18634,N_18357,N_18493);
and U18635 (N_18635,N_18287,N_18311);
and U18636 (N_18636,N_18445,N_18338);
xor U18637 (N_18637,N_18322,N_18448);
nor U18638 (N_18638,N_18397,N_18349);
or U18639 (N_18639,N_18497,N_18265);
and U18640 (N_18640,N_18454,N_18336);
nand U18641 (N_18641,N_18369,N_18362);
nor U18642 (N_18642,N_18377,N_18458);
nor U18643 (N_18643,N_18303,N_18269);
or U18644 (N_18644,N_18483,N_18408);
nand U18645 (N_18645,N_18325,N_18306);
and U18646 (N_18646,N_18378,N_18346);
nor U18647 (N_18647,N_18317,N_18321);
or U18648 (N_18648,N_18332,N_18296);
nor U18649 (N_18649,N_18423,N_18364);
or U18650 (N_18650,N_18486,N_18498);
xor U18651 (N_18651,N_18491,N_18494);
and U18652 (N_18652,N_18444,N_18302);
nor U18653 (N_18653,N_18374,N_18379);
and U18654 (N_18654,N_18349,N_18376);
or U18655 (N_18655,N_18442,N_18269);
xnor U18656 (N_18656,N_18408,N_18460);
nor U18657 (N_18657,N_18294,N_18448);
or U18658 (N_18658,N_18459,N_18300);
nor U18659 (N_18659,N_18447,N_18292);
nand U18660 (N_18660,N_18451,N_18332);
or U18661 (N_18661,N_18474,N_18461);
nor U18662 (N_18662,N_18275,N_18421);
and U18663 (N_18663,N_18365,N_18392);
xnor U18664 (N_18664,N_18493,N_18256);
nand U18665 (N_18665,N_18278,N_18270);
nand U18666 (N_18666,N_18329,N_18388);
or U18667 (N_18667,N_18296,N_18279);
nor U18668 (N_18668,N_18324,N_18488);
or U18669 (N_18669,N_18301,N_18459);
nand U18670 (N_18670,N_18315,N_18375);
nand U18671 (N_18671,N_18447,N_18397);
and U18672 (N_18672,N_18344,N_18460);
nand U18673 (N_18673,N_18437,N_18291);
nand U18674 (N_18674,N_18357,N_18417);
xnor U18675 (N_18675,N_18451,N_18302);
or U18676 (N_18676,N_18420,N_18472);
or U18677 (N_18677,N_18332,N_18477);
and U18678 (N_18678,N_18287,N_18345);
xor U18679 (N_18679,N_18340,N_18484);
and U18680 (N_18680,N_18347,N_18276);
or U18681 (N_18681,N_18397,N_18316);
xor U18682 (N_18682,N_18468,N_18450);
xnor U18683 (N_18683,N_18355,N_18311);
xor U18684 (N_18684,N_18362,N_18298);
xor U18685 (N_18685,N_18363,N_18409);
and U18686 (N_18686,N_18275,N_18384);
nand U18687 (N_18687,N_18439,N_18276);
xor U18688 (N_18688,N_18397,N_18357);
or U18689 (N_18689,N_18443,N_18475);
or U18690 (N_18690,N_18445,N_18306);
and U18691 (N_18691,N_18285,N_18455);
or U18692 (N_18692,N_18333,N_18351);
nor U18693 (N_18693,N_18284,N_18410);
xor U18694 (N_18694,N_18267,N_18292);
nor U18695 (N_18695,N_18292,N_18451);
xnor U18696 (N_18696,N_18306,N_18422);
nand U18697 (N_18697,N_18446,N_18324);
and U18698 (N_18698,N_18487,N_18329);
nand U18699 (N_18699,N_18256,N_18398);
nand U18700 (N_18700,N_18390,N_18325);
and U18701 (N_18701,N_18374,N_18482);
xnor U18702 (N_18702,N_18260,N_18497);
nand U18703 (N_18703,N_18455,N_18373);
or U18704 (N_18704,N_18265,N_18391);
nand U18705 (N_18705,N_18410,N_18273);
nand U18706 (N_18706,N_18444,N_18463);
xnor U18707 (N_18707,N_18480,N_18499);
nor U18708 (N_18708,N_18497,N_18362);
nand U18709 (N_18709,N_18301,N_18441);
nand U18710 (N_18710,N_18445,N_18293);
or U18711 (N_18711,N_18465,N_18368);
or U18712 (N_18712,N_18323,N_18476);
xor U18713 (N_18713,N_18413,N_18324);
xnor U18714 (N_18714,N_18426,N_18332);
and U18715 (N_18715,N_18363,N_18355);
nand U18716 (N_18716,N_18408,N_18464);
nand U18717 (N_18717,N_18399,N_18362);
and U18718 (N_18718,N_18412,N_18312);
or U18719 (N_18719,N_18330,N_18280);
nand U18720 (N_18720,N_18423,N_18478);
and U18721 (N_18721,N_18421,N_18250);
or U18722 (N_18722,N_18318,N_18387);
nand U18723 (N_18723,N_18360,N_18329);
and U18724 (N_18724,N_18346,N_18328);
or U18725 (N_18725,N_18266,N_18484);
xnor U18726 (N_18726,N_18479,N_18405);
xor U18727 (N_18727,N_18373,N_18467);
xor U18728 (N_18728,N_18335,N_18423);
nor U18729 (N_18729,N_18272,N_18467);
nor U18730 (N_18730,N_18301,N_18365);
and U18731 (N_18731,N_18340,N_18292);
nand U18732 (N_18732,N_18309,N_18334);
nor U18733 (N_18733,N_18428,N_18350);
and U18734 (N_18734,N_18444,N_18254);
xnor U18735 (N_18735,N_18384,N_18343);
xor U18736 (N_18736,N_18382,N_18316);
nor U18737 (N_18737,N_18494,N_18307);
and U18738 (N_18738,N_18308,N_18284);
nor U18739 (N_18739,N_18483,N_18306);
nor U18740 (N_18740,N_18279,N_18441);
or U18741 (N_18741,N_18339,N_18381);
or U18742 (N_18742,N_18257,N_18318);
nor U18743 (N_18743,N_18353,N_18358);
nor U18744 (N_18744,N_18404,N_18382);
and U18745 (N_18745,N_18278,N_18447);
and U18746 (N_18746,N_18270,N_18448);
or U18747 (N_18747,N_18369,N_18403);
nand U18748 (N_18748,N_18424,N_18417);
nand U18749 (N_18749,N_18434,N_18385);
nand U18750 (N_18750,N_18700,N_18731);
nand U18751 (N_18751,N_18712,N_18665);
nand U18752 (N_18752,N_18702,N_18629);
nand U18753 (N_18753,N_18695,N_18652);
or U18754 (N_18754,N_18696,N_18694);
nor U18755 (N_18755,N_18707,N_18518);
xor U18756 (N_18756,N_18595,N_18587);
nor U18757 (N_18757,N_18542,N_18739);
or U18758 (N_18758,N_18504,N_18687);
xor U18759 (N_18759,N_18507,N_18586);
xnor U18760 (N_18760,N_18566,N_18506);
nor U18761 (N_18761,N_18666,N_18724);
xor U18762 (N_18762,N_18670,N_18641);
or U18763 (N_18763,N_18512,N_18502);
or U18764 (N_18764,N_18647,N_18588);
nand U18765 (N_18765,N_18740,N_18612);
or U18766 (N_18766,N_18668,N_18598);
and U18767 (N_18767,N_18547,N_18727);
nor U18768 (N_18768,N_18624,N_18720);
nand U18769 (N_18769,N_18683,N_18725);
or U18770 (N_18770,N_18619,N_18555);
xnor U18771 (N_18771,N_18645,N_18519);
or U18772 (N_18772,N_18600,N_18563);
xnor U18773 (N_18773,N_18510,N_18523);
nand U18774 (N_18774,N_18620,N_18582);
and U18775 (N_18775,N_18734,N_18508);
or U18776 (N_18776,N_18562,N_18597);
and U18777 (N_18777,N_18591,N_18560);
and U18778 (N_18778,N_18548,N_18608);
xnor U18779 (N_18779,N_18743,N_18556);
or U18780 (N_18780,N_18644,N_18660);
xnor U18781 (N_18781,N_18579,N_18524);
and U18782 (N_18782,N_18703,N_18733);
nand U18783 (N_18783,N_18708,N_18677);
nor U18784 (N_18784,N_18564,N_18594);
and U18785 (N_18785,N_18747,N_18517);
xnor U18786 (N_18786,N_18537,N_18672);
nand U18787 (N_18787,N_18623,N_18601);
xor U18788 (N_18788,N_18546,N_18651);
nand U18789 (N_18789,N_18583,N_18580);
and U18790 (N_18790,N_18554,N_18749);
xor U18791 (N_18791,N_18643,N_18704);
nand U18792 (N_18792,N_18678,N_18661);
nor U18793 (N_18793,N_18689,N_18551);
xor U18794 (N_18794,N_18646,N_18557);
and U18795 (N_18795,N_18549,N_18540);
nor U18796 (N_18796,N_18627,N_18631);
xor U18797 (N_18797,N_18584,N_18536);
and U18798 (N_18798,N_18658,N_18729);
nor U18799 (N_18799,N_18710,N_18685);
nand U18800 (N_18800,N_18552,N_18717);
or U18801 (N_18801,N_18680,N_18625);
or U18802 (N_18802,N_18573,N_18669);
or U18803 (N_18803,N_18663,N_18539);
nand U18804 (N_18804,N_18513,N_18633);
nand U18805 (N_18805,N_18576,N_18714);
nor U18806 (N_18806,N_18701,N_18721);
nor U18807 (N_18807,N_18742,N_18691);
xor U18808 (N_18808,N_18569,N_18514);
xnor U18809 (N_18809,N_18533,N_18745);
nor U18810 (N_18810,N_18532,N_18527);
and U18811 (N_18811,N_18520,N_18607);
and U18812 (N_18812,N_18500,N_18503);
xor U18813 (N_18813,N_18692,N_18738);
nand U18814 (N_18814,N_18662,N_18626);
nor U18815 (N_18815,N_18723,N_18737);
nor U18816 (N_18816,N_18654,N_18715);
or U18817 (N_18817,N_18559,N_18541);
or U18818 (N_18818,N_18719,N_18611);
xor U18819 (N_18819,N_18693,N_18642);
or U18820 (N_18820,N_18574,N_18679);
or U18821 (N_18821,N_18614,N_18675);
and U18822 (N_18822,N_18676,N_18593);
and U18823 (N_18823,N_18565,N_18671);
nor U18824 (N_18824,N_18570,N_18516);
xnor U18825 (N_18825,N_18705,N_18572);
and U18826 (N_18826,N_18634,N_18613);
nand U18827 (N_18827,N_18610,N_18553);
and U18828 (N_18828,N_18728,N_18726);
or U18829 (N_18829,N_18630,N_18699);
and U18830 (N_18830,N_18718,N_18592);
nand U18831 (N_18831,N_18684,N_18505);
or U18832 (N_18832,N_18578,N_18618);
xnor U18833 (N_18833,N_18509,N_18511);
nor U18834 (N_18834,N_18674,N_18664);
nor U18835 (N_18835,N_18711,N_18690);
and U18836 (N_18836,N_18697,N_18653);
xor U18837 (N_18837,N_18709,N_18655);
or U18838 (N_18838,N_18659,N_18713);
or U18839 (N_18839,N_18628,N_18602);
xor U18840 (N_18840,N_18575,N_18730);
or U18841 (N_18841,N_18648,N_18637);
or U18842 (N_18842,N_18609,N_18535);
or U18843 (N_18843,N_18525,N_18617);
xor U18844 (N_18844,N_18673,N_18567);
xor U18845 (N_18845,N_18688,N_18615);
xnor U18846 (N_18846,N_18568,N_18522);
xnor U18847 (N_18847,N_18736,N_18589);
nand U18848 (N_18848,N_18649,N_18526);
and U18849 (N_18849,N_18521,N_18744);
nor U18850 (N_18850,N_18545,N_18550);
nor U18851 (N_18851,N_18732,N_18590);
or U18852 (N_18852,N_18616,N_18530);
nand U18853 (N_18853,N_18501,N_18640);
nand U18854 (N_18854,N_18621,N_18558);
nand U18855 (N_18855,N_18635,N_18622);
or U18856 (N_18856,N_18604,N_18686);
nand U18857 (N_18857,N_18638,N_18657);
nor U18858 (N_18858,N_18741,N_18561);
xor U18859 (N_18859,N_18603,N_18528);
and U18860 (N_18860,N_18538,N_18599);
nand U18861 (N_18861,N_18639,N_18534);
or U18862 (N_18862,N_18636,N_18735);
or U18863 (N_18863,N_18605,N_18722);
nor U18864 (N_18864,N_18606,N_18581);
nor U18865 (N_18865,N_18682,N_18746);
and U18866 (N_18866,N_18632,N_18543);
xnor U18867 (N_18867,N_18596,N_18706);
nand U18868 (N_18868,N_18585,N_18650);
and U18869 (N_18869,N_18544,N_18656);
or U18870 (N_18870,N_18577,N_18667);
or U18871 (N_18871,N_18571,N_18698);
xor U18872 (N_18872,N_18515,N_18748);
xor U18873 (N_18873,N_18531,N_18716);
xnor U18874 (N_18874,N_18529,N_18681);
or U18875 (N_18875,N_18739,N_18679);
nand U18876 (N_18876,N_18720,N_18517);
nor U18877 (N_18877,N_18520,N_18564);
and U18878 (N_18878,N_18644,N_18503);
nor U18879 (N_18879,N_18668,N_18623);
xnor U18880 (N_18880,N_18525,N_18627);
nor U18881 (N_18881,N_18578,N_18598);
and U18882 (N_18882,N_18664,N_18513);
xnor U18883 (N_18883,N_18576,N_18667);
or U18884 (N_18884,N_18586,N_18624);
or U18885 (N_18885,N_18534,N_18740);
xnor U18886 (N_18886,N_18749,N_18659);
nor U18887 (N_18887,N_18704,N_18520);
xor U18888 (N_18888,N_18660,N_18610);
or U18889 (N_18889,N_18719,N_18615);
nand U18890 (N_18890,N_18569,N_18593);
xnor U18891 (N_18891,N_18607,N_18667);
nand U18892 (N_18892,N_18733,N_18644);
and U18893 (N_18893,N_18599,N_18525);
or U18894 (N_18894,N_18691,N_18656);
and U18895 (N_18895,N_18680,N_18510);
xnor U18896 (N_18896,N_18733,N_18746);
nor U18897 (N_18897,N_18532,N_18695);
or U18898 (N_18898,N_18535,N_18511);
nand U18899 (N_18899,N_18645,N_18672);
or U18900 (N_18900,N_18714,N_18520);
nor U18901 (N_18901,N_18686,N_18589);
and U18902 (N_18902,N_18609,N_18579);
nand U18903 (N_18903,N_18581,N_18667);
nand U18904 (N_18904,N_18629,N_18605);
and U18905 (N_18905,N_18748,N_18543);
and U18906 (N_18906,N_18537,N_18504);
and U18907 (N_18907,N_18594,N_18694);
or U18908 (N_18908,N_18679,N_18636);
nor U18909 (N_18909,N_18732,N_18531);
and U18910 (N_18910,N_18589,N_18720);
xor U18911 (N_18911,N_18696,N_18546);
nand U18912 (N_18912,N_18510,N_18679);
and U18913 (N_18913,N_18673,N_18711);
nor U18914 (N_18914,N_18502,N_18570);
nor U18915 (N_18915,N_18611,N_18515);
and U18916 (N_18916,N_18565,N_18531);
and U18917 (N_18917,N_18536,N_18674);
xnor U18918 (N_18918,N_18527,N_18647);
or U18919 (N_18919,N_18500,N_18685);
and U18920 (N_18920,N_18706,N_18568);
nand U18921 (N_18921,N_18711,N_18506);
and U18922 (N_18922,N_18550,N_18592);
xor U18923 (N_18923,N_18574,N_18558);
or U18924 (N_18924,N_18535,N_18557);
nor U18925 (N_18925,N_18702,N_18581);
xnor U18926 (N_18926,N_18696,N_18640);
and U18927 (N_18927,N_18655,N_18664);
or U18928 (N_18928,N_18692,N_18520);
xor U18929 (N_18929,N_18545,N_18748);
nand U18930 (N_18930,N_18640,N_18657);
and U18931 (N_18931,N_18715,N_18688);
nand U18932 (N_18932,N_18613,N_18560);
nor U18933 (N_18933,N_18668,N_18523);
xnor U18934 (N_18934,N_18671,N_18623);
xor U18935 (N_18935,N_18690,N_18731);
nand U18936 (N_18936,N_18693,N_18533);
nand U18937 (N_18937,N_18666,N_18678);
nor U18938 (N_18938,N_18554,N_18525);
or U18939 (N_18939,N_18501,N_18684);
nor U18940 (N_18940,N_18704,N_18616);
nand U18941 (N_18941,N_18682,N_18558);
nor U18942 (N_18942,N_18632,N_18680);
and U18943 (N_18943,N_18560,N_18678);
or U18944 (N_18944,N_18519,N_18685);
nand U18945 (N_18945,N_18723,N_18711);
and U18946 (N_18946,N_18740,N_18524);
xor U18947 (N_18947,N_18590,N_18555);
or U18948 (N_18948,N_18635,N_18722);
xor U18949 (N_18949,N_18574,N_18672);
and U18950 (N_18950,N_18742,N_18672);
or U18951 (N_18951,N_18547,N_18633);
xnor U18952 (N_18952,N_18658,N_18725);
nor U18953 (N_18953,N_18556,N_18718);
and U18954 (N_18954,N_18563,N_18710);
and U18955 (N_18955,N_18673,N_18509);
or U18956 (N_18956,N_18640,N_18553);
and U18957 (N_18957,N_18550,N_18732);
and U18958 (N_18958,N_18602,N_18714);
nand U18959 (N_18959,N_18535,N_18626);
xor U18960 (N_18960,N_18537,N_18577);
nand U18961 (N_18961,N_18515,N_18626);
nand U18962 (N_18962,N_18690,N_18737);
nand U18963 (N_18963,N_18539,N_18649);
or U18964 (N_18964,N_18555,N_18596);
and U18965 (N_18965,N_18551,N_18742);
or U18966 (N_18966,N_18696,N_18628);
nand U18967 (N_18967,N_18636,N_18580);
xor U18968 (N_18968,N_18603,N_18734);
nor U18969 (N_18969,N_18727,N_18555);
or U18970 (N_18970,N_18611,N_18555);
or U18971 (N_18971,N_18702,N_18566);
and U18972 (N_18972,N_18510,N_18644);
nor U18973 (N_18973,N_18628,N_18605);
xnor U18974 (N_18974,N_18737,N_18558);
nor U18975 (N_18975,N_18582,N_18534);
nor U18976 (N_18976,N_18716,N_18679);
or U18977 (N_18977,N_18701,N_18639);
xnor U18978 (N_18978,N_18538,N_18734);
nor U18979 (N_18979,N_18603,N_18649);
and U18980 (N_18980,N_18749,N_18719);
or U18981 (N_18981,N_18730,N_18629);
xnor U18982 (N_18982,N_18520,N_18659);
nor U18983 (N_18983,N_18667,N_18741);
nand U18984 (N_18984,N_18590,N_18502);
or U18985 (N_18985,N_18555,N_18545);
nor U18986 (N_18986,N_18532,N_18538);
or U18987 (N_18987,N_18509,N_18703);
and U18988 (N_18988,N_18698,N_18616);
and U18989 (N_18989,N_18523,N_18695);
nand U18990 (N_18990,N_18637,N_18631);
nand U18991 (N_18991,N_18502,N_18546);
nand U18992 (N_18992,N_18744,N_18702);
or U18993 (N_18993,N_18650,N_18648);
xnor U18994 (N_18994,N_18624,N_18651);
xor U18995 (N_18995,N_18629,N_18652);
or U18996 (N_18996,N_18744,N_18567);
nor U18997 (N_18997,N_18502,N_18566);
and U18998 (N_18998,N_18647,N_18742);
nor U18999 (N_18999,N_18610,N_18699);
nand U19000 (N_19000,N_18881,N_18892);
and U19001 (N_19001,N_18987,N_18767);
and U19002 (N_19002,N_18945,N_18832);
or U19003 (N_19003,N_18970,N_18776);
nor U19004 (N_19004,N_18915,N_18791);
xor U19005 (N_19005,N_18806,N_18789);
xor U19006 (N_19006,N_18836,N_18998);
nand U19007 (N_19007,N_18982,N_18751);
nand U19008 (N_19008,N_18844,N_18980);
nor U19009 (N_19009,N_18777,N_18922);
nand U19010 (N_19010,N_18882,N_18939);
or U19011 (N_19011,N_18925,N_18961);
nor U19012 (N_19012,N_18808,N_18784);
or U19013 (N_19013,N_18849,N_18774);
or U19014 (N_19014,N_18753,N_18921);
or U19015 (N_19015,N_18920,N_18802);
or U19016 (N_19016,N_18821,N_18977);
nand U19017 (N_19017,N_18887,N_18861);
nand U19018 (N_19018,N_18933,N_18799);
and U19019 (N_19019,N_18962,N_18807);
or U19020 (N_19020,N_18830,N_18828);
nor U19021 (N_19021,N_18946,N_18877);
and U19022 (N_19022,N_18983,N_18816);
and U19023 (N_19023,N_18827,N_18984);
nand U19024 (N_19024,N_18842,N_18848);
nand U19025 (N_19025,N_18936,N_18876);
nor U19026 (N_19026,N_18964,N_18800);
nand U19027 (N_19027,N_18905,N_18896);
or U19028 (N_19028,N_18752,N_18953);
nand U19029 (N_19029,N_18888,N_18912);
nor U19030 (N_19030,N_18768,N_18759);
nand U19031 (N_19031,N_18902,N_18914);
nand U19032 (N_19032,N_18763,N_18911);
nor U19033 (N_19033,N_18760,N_18762);
xnor U19034 (N_19034,N_18958,N_18804);
or U19035 (N_19035,N_18875,N_18974);
nor U19036 (N_19036,N_18972,N_18909);
or U19037 (N_19037,N_18997,N_18989);
nand U19038 (N_19038,N_18996,N_18765);
nor U19039 (N_19039,N_18831,N_18908);
nand U19040 (N_19040,N_18840,N_18867);
xor U19041 (N_19041,N_18822,N_18856);
or U19042 (N_19042,N_18775,N_18754);
nor U19043 (N_19043,N_18895,N_18868);
and U19044 (N_19044,N_18750,N_18801);
and U19045 (N_19045,N_18793,N_18779);
nor U19046 (N_19046,N_18937,N_18930);
or U19047 (N_19047,N_18986,N_18812);
nor U19048 (N_19048,N_18969,N_18992);
nor U19049 (N_19049,N_18883,N_18786);
and U19050 (N_19050,N_18813,N_18924);
nor U19051 (N_19051,N_18947,N_18963);
or U19052 (N_19052,N_18880,N_18764);
xnor U19053 (N_19053,N_18820,N_18917);
or U19054 (N_19054,N_18761,N_18913);
and U19055 (N_19055,N_18781,N_18951);
nor U19056 (N_19056,N_18771,N_18841);
and U19057 (N_19057,N_18959,N_18859);
nand U19058 (N_19058,N_18973,N_18919);
nand U19059 (N_19059,N_18783,N_18843);
or U19060 (N_19060,N_18787,N_18966);
or U19061 (N_19061,N_18854,N_18770);
or U19062 (N_19062,N_18901,N_18869);
xor U19063 (N_19063,N_18978,N_18906);
nand U19064 (N_19064,N_18810,N_18870);
and U19065 (N_19065,N_18903,N_18805);
nand U19066 (N_19066,N_18798,N_18904);
or U19067 (N_19067,N_18889,N_18772);
and U19068 (N_19068,N_18845,N_18999);
or U19069 (N_19069,N_18858,N_18857);
nand U19070 (N_19070,N_18835,N_18834);
and U19071 (N_19071,N_18872,N_18886);
or U19072 (N_19072,N_18795,N_18991);
and U19073 (N_19073,N_18851,N_18866);
and U19074 (N_19074,N_18935,N_18934);
nor U19075 (N_19075,N_18954,N_18850);
nand U19076 (N_19076,N_18757,N_18780);
and U19077 (N_19077,N_18817,N_18910);
and U19078 (N_19078,N_18981,N_18988);
nor U19079 (N_19079,N_18918,N_18773);
nand U19080 (N_19080,N_18847,N_18826);
or U19081 (N_19081,N_18769,N_18891);
xnor U19082 (N_19082,N_18790,N_18976);
nor U19083 (N_19083,N_18879,N_18894);
or U19084 (N_19084,N_18927,N_18949);
nand U19085 (N_19085,N_18893,N_18907);
nand U19086 (N_19086,N_18846,N_18792);
nand U19087 (N_19087,N_18853,N_18803);
and U19088 (N_19088,N_18852,N_18766);
or U19089 (N_19089,N_18755,N_18855);
nand U19090 (N_19090,N_18956,N_18985);
and U19091 (N_19091,N_18758,N_18990);
or U19092 (N_19092,N_18897,N_18878);
or U19093 (N_19093,N_18952,N_18885);
nor U19094 (N_19094,N_18943,N_18873);
nor U19095 (N_19095,N_18971,N_18899);
nand U19096 (N_19096,N_18965,N_18818);
nor U19097 (N_19097,N_18837,N_18829);
xnor U19098 (N_19098,N_18950,N_18957);
nand U19099 (N_19099,N_18900,N_18928);
nor U19100 (N_19100,N_18926,N_18898);
nand U19101 (N_19101,N_18788,N_18944);
nor U19102 (N_19102,N_18890,N_18811);
nor U19103 (N_19103,N_18860,N_18923);
and U19104 (N_19104,N_18838,N_18871);
and U19105 (N_19105,N_18929,N_18815);
or U19106 (N_19106,N_18825,N_18993);
or U19107 (N_19107,N_18824,N_18864);
xor U19108 (N_19108,N_18931,N_18782);
nor U19109 (N_19109,N_18809,N_18916);
and U19110 (N_19110,N_18975,N_18932);
and U19111 (N_19111,N_18955,N_18833);
and U19112 (N_19112,N_18863,N_18823);
or U19113 (N_19113,N_18968,N_18814);
nand U19114 (N_19114,N_18778,N_18960);
nor U19115 (N_19115,N_18865,N_18884);
nand U19116 (N_19116,N_18948,N_18862);
or U19117 (N_19117,N_18967,N_18796);
xnor U19118 (N_19118,N_18756,N_18819);
or U19119 (N_19119,N_18785,N_18839);
nor U19120 (N_19120,N_18874,N_18794);
or U19121 (N_19121,N_18940,N_18995);
nand U19122 (N_19122,N_18994,N_18941);
xor U19123 (N_19123,N_18942,N_18797);
nor U19124 (N_19124,N_18979,N_18938);
xnor U19125 (N_19125,N_18846,N_18912);
xnor U19126 (N_19126,N_18840,N_18958);
or U19127 (N_19127,N_18968,N_18813);
nor U19128 (N_19128,N_18950,N_18993);
nor U19129 (N_19129,N_18855,N_18978);
xnor U19130 (N_19130,N_18807,N_18894);
xor U19131 (N_19131,N_18798,N_18976);
nor U19132 (N_19132,N_18893,N_18971);
nor U19133 (N_19133,N_18883,N_18973);
or U19134 (N_19134,N_18908,N_18878);
xnor U19135 (N_19135,N_18773,N_18789);
nand U19136 (N_19136,N_18759,N_18773);
nor U19137 (N_19137,N_18860,N_18925);
nand U19138 (N_19138,N_18984,N_18798);
or U19139 (N_19139,N_18900,N_18884);
xor U19140 (N_19140,N_18806,N_18881);
or U19141 (N_19141,N_18932,N_18877);
and U19142 (N_19142,N_18940,N_18957);
nor U19143 (N_19143,N_18955,N_18818);
and U19144 (N_19144,N_18986,N_18939);
xor U19145 (N_19145,N_18764,N_18872);
nor U19146 (N_19146,N_18843,N_18930);
xnor U19147 (N_19147,N_18954,N_18859);
or U19148 (N_19148,N_18902,N_18979);
nand U19149 (N_19149,N_18897,N_18894);
nand U19150 (N_19150,N_18919,N_18917);
xnor U19151 (N_19151,N_18762,N_18757);
nand U19152 (N_19152,N_18779,N_18993);
and U19153 (N_19153,N_18856,N_18945);
or U19154 (N_19154,N_18969,N_18803);
and U19155 (N_19155,N_18829,N_18756);
nor U19156 (N_19156,N_18917,N_18929);
and U19157 (N_19157,N_18892,N_18782);
nand U19158 (N_19158,N_18828,N_18847);
xnor U19159 (N_19159,N_18885,N_18761);
nor U19160 (N_19160,N_18790,N_18905);
nand U19161 (N_19161,N_18996,N_18907);
or U19162 (N_19162,N_18867,N_18860);
nor U19163 (N_19163,N_18977,N_18797);
or U19164 (N_19164,N_18953,N_18781);
nand U19165 (N_19165,N_18800,N_18812);
or U19166 (N_19166,N_18955,N_18896);
nor U19167 (N_19167,N_18916,N_18837);
and U19168 (N_19168,N_18969,N_18864);
xor U19169 (N_19169,N_18984,N_18755);
nand U19170 (N_19170,N_18853,N_18955);
nand U19171 (N_19171,N_18805,N_18772);
and U19172 (N_19172,N_18900,N_18848);
or U19173 (N_19173,N_18899,N_18756);
xnor U19174 (N_19174,N_18954,N_18884);
and U19175 (N_19175,N_18997,N_18855);
and U19176 (N_19176,N_18903,N_18852);
nand U19177 (N_19177,N_18931,N_18865);
and U19178 (N_19178,N_18820,N_18810);
or U19179 (N_19179,N_18807,N_18757);
xor U19180 (N_19180,N_18948,N_18958);
nand U19181 (N_19181,N_18867,N_18871);
and U19182 (N_19182,N_18832,N_18969);
and U19183 (N_19183,N_18924,N_18910);
nor U19184 (N_19184,N_18986,N_18753);
or U19185 (N_19185,N_18886,N_18859);
nor U19186 (N_19186,N_18985,N_18860);
xor U19187 (N_19187,N_18969,N_18822);
or U19188 (N_19188,N_18802,N_18889);
or U19189 (N_19189,N_18911,N_18844);
nor U19190 (N_19190,N_18958,N_18824);
xnor U19191 (N_19191,N_18775,N_18799);
and U19192 (N_19192,N_18984,N_18931);
nand U19193 (N_19193,N_18903,N_18899);
or U19194 (N_19194,N_18841,N_18968);
nand U19195 (N_19195,N_18954,N_18991);
or U19196 (N_19196,N_18760,N_18781);
nand U19197 (N_19197,N_18937,N_18774);
and U19198 (N_19198,N_18818,N_18854);
and U19199 (N_19199,N_18901,N_18788);
or U19200 (N_19200,N_18866,N_18872);
and U19201 (N_19201,N_18950,N_18953);
nor U19202 (N_19202,N_18876,N_18861);
nor U19203 (N_19203,N_18807,N_18765);
nand U19204 (N_19204,N_18904,N_18960);
nor U19205 (N_19205,N_18971,N_18964);
xnor U19206 (N_19206,N_18878,N_18792);
nor U19207 (N_19207,N_18914,N_18946);
or U19208 (N_19208,N_18835,N_18884);
xor U19209 (N_19209,N_18848,N_18840);
nor U19210 (N_19210,N_18878,N_18791);
nand U19211 (N_19211,N_18841,N_18898);
xnor U19212 (N_19212,N_18911,N_18776);
nor U19213 (N_19213,N_18949,N_18982);
or U19214 (N_19214,N_18750,N_18924);
xnor U19215 (N_19215,N_18937,N_18888);
nor U19216 (N_19216,N_18765,N_18929);
or U19217 (N_19217,N_18917,N_18838);
and U19218 (N_19218,N_18848,N_18898);
and U19219 (N_19219,N_18889,N_18912);
nand U19220 (N_19220,N_18778,N_18994);
nor U19221 (N_19221,N_18794,N_18840);
or U19222 (N_19222,N_18937,N_18932);
nand U19223 (N_19223,N_18957,N_18805);
nand U19224 (N_19224,N_18783,N_18761);
or U19225 (N_19225,N_18769,N_18953);
or U19226 (N_19226,N_18755,N_18834);
or U19227 (N_19227,N_18968,N_18822);
nor U19228 (N_19228,N_18955,N_18899);
nand U19229 (N_19229,N_18782,N_18834);
nand U19230 (N_19230,N_18781,N_18873);
xnor U19231 (N_19231,N_18783,N_18940);
nor U19232 (N_19232,N_18911,N_18851);
nor U19233 (N_19233,N_18869,N_18975);
and U19234 (N_19234,N_18832,N_18778);
xnor U19235 (N_19235,N_18860,N_18911);
or U19236 (N_19236,N_18840,N_18758);
nor U19237 (N_19237,N_18814,N_18755);
nor U19238 (N_19238,N_18904,N_18926);
and U19239 (N_19239,N_18835,N_18839);
and U19240 (N_19240,N_18872,N_18774);
or U19241 (N_19241,N_18967,N_18868);
nand U19242 (N_19242,N_18981,N_18908);
xnor U19243 (N_19243,N_18907,N_18837);
nor U19244 (N_19244,N_18798,N_18988);
nor U19245 (N_19245,N_18934,N_18781);
nand U19246 (N_19246,N_18822,N_18752);
xor U19247 (N_19247,N_18883,N_18932);
and U19248 (N_19248,N_18793,N_18762);
xnor U19249 (N_19249,N_18993,N_18812);
and U19250 (N_19250,N_19117,N_19087);
xnor U19251 (N_19251,N_19057,N_19081);
and U19252 (N_19252,N_19116,N_19180);
nor U19253 (N_19253,N_19068,N_19203);
or U19254 (N_19254,N_19131,N_19166);
or U19255 (N_19255,N_19167,N_19055);
xor U19256 (N_19256,N_19237,N_19066);
or U19257 (N_19257,N_19128,N_19205);
nand U19258 (N_19258,N_19224,N_19101);
nand U19259 (N_19259,N_19236,N_19230);
nor U19260 (N_19260,N_19215,N_19130);
or U19261 (N_19261,N_19077,N_19126);
or U19262 (N_19262,N_19218,N_19233);
or U19263 (N_19263,N_19226,N_19085);
nor U19264 (N_19264,N_19151,N_19178);
and U19265 (N_19265,N_19073,N_19204);
nand U19266 (N_19266,N_19028,N_19051);
and U19267 (N_19267,N_19111,N_19125);
xor U19268 (N_19268,N_19133,N_19071);
and U19269 (N_19269,N_19026,N_19056);
nand U19270 (N_19270,N_19023,N_19162);
nand U19271 (N_19271,N_19053,N_19084);
or U19272 (N_19272,N_19090,N_19222);
nor U19273 (N_19273,N_19198,N_19091);
or U19274 (N_19274,N_19083,N_19160);
xnor U19275 (N_19275,N_19105,N_19127);
xnor U19276 (N_19276,N_19246,N_19059);
and U19277 (N_19277,N_19248,N_19199);
nor U19278 (N_19278,N_19074,N_19046);
xor U19279 (N_19279,N_19016,N_19145);
nand U19280 (N_19280,N_19197,N_19219);
or U19281 (N_19281,N_19123,N_19153);
and U19282 (N_19282,N_19165,N_19100);
and U19283 (N_19283,N_19006,N_19141);
xor U19284 (N_19284,N_19072,N_19092);
xnor U19285 (N_19285,N_19062,N_19168);
and U19286 (N_19286,N_19142,N_19060);
and U19287 (N_19287,N_19047,N_19192);
nor U19288 (N_19288,N_19030,N_19078);
or U19289 (N_19289,N_19098,N_19177);
and U19290 (N_19290,N_19052,N_19185);
and U19291 (N_19291,N_19103,N_19225);
nor U19292 (N_19292,N_19147,N_19058);
nand U19293 (N_19293,N_19120,N_19208);
nor U19294 (N_19294,N_19044,N_19106);
and U19295 (N_19295,N_19234,N_19093);
or U19296 (N_19296,N_19201,N_19174);
nand U19297 (N_19297,N_19029,N_19207);
and U19298 (N_19298,N_19002,N_19136);
or U19299 (N_19299,N_19036,N_19137);
nor U19300 (N_19300,N_19012,N_19021);
xor U19301 (N_19301,N_19183,N_19070);
or U19302 (N_19302,N_19027,N_19195);
or U19303 (N_19303,N_19176,N_19249);
and U19304 (N_19304,N_19164,N_19159);
nor U19305 (N_19305,N_19170,N_19034);
nor U19306 (N_19306,N_19194,N_19099);
nor U19307 (N_19307,N_19188,N_19042);
nor U19308 (N_19308,N_19200,N_19080);
nor U19309 (N_19309,N_19015,N_19220);
and U19310 (N_19310,N_19112,N_19228);
xor U19311 (N_19311,N_19017,N_19157);
xnor U19312 (N_19312,N_19007,N_19108);
nand U19313 (N_19313,N_19181,N_19206);
or U19314 (N_19314,N_19132,N_19152);
or U19315 (N_19315,N_19020,N_19032);
and U19316 (N_19316,N_19033,N_19114);
or U19317 (N_19317,N_19229,N_19003);
nor U19318 (N_19318,N_19129,N_19172);
or U19319 (N_19319,N_19216,N_19061);
nor U19320 (N_19320,N_19113,N_19109);
nand U19321 (N_19321,N_19156,N_19211);
and U19322 (N_19322,N_19054,N_19049);
and U19323 (N_19323,N_19094,N_19191);
nand U19324 (N_19324,N_19031,N_19223);
or U19325 (N_19325,N_19134,N_19050);
or U19326 (N_19326,N_19144,N_19155);
or U19327 (N_19327,N_19014,N_19227);
nand U19328 (N_19328,N_19244,N_19004);
and U19329 (N_19329,N_19102,N_19019);
xor U19330 (N_19330,N_19063,N_19231);
nand U19331 (N_19331,N_19115,N_19107);
nor U19332 (N_19332,N_19139,N_19124);
nand U19333 (N_19333,N_19213,N_19212);
nand U19334 (N_19334,N_19193,N_19140);
or U19335 (N_19335,N_19008,N_19182);
nand U19336 (N_19336,N_19005,N_19149);
or U19337 (N_19337,N_19158,N_19175);
and U19338 (N_19338,N_19122,N_19187);
or U19339 (N_19339,N_19035,N_19095);
or U19340 (N_19340,N_19240,N_19039);
nand U19341 (N_19341,N_19179,N_19064);
and U19342 (N_19342,N_19082,N_19041);
nand U19343 (N_19343,N_19243,N_19138);
or U19344 (N_19344,N_19119,N_19186);
xnor U19345 (N_19345,N_19086,N_19096);
nand U19346 (N_19346,N_19067,N_19245);
xor U19347 (N_19347,N_19239,N_19121);
or U19348 (N_19348,N_19089,N_19171);
or U19349 (N_19349,N_19018,N_19075);
or U19350 (N_19350,N_19214,N_19011);
nand U19351 (N_19351,N_19169,N_19010);
or U19352 (N_19352,N_19242,N_19146);
and U19353 (N_19353,N_19163,N_19210);
nor U19354 (N_19354,N_19076,N_19104);
and U19355 (N_19355,N_19097,N_19196);
nor U19356 (N_19356,N_19154,N_19217);
or U19357 (N_19357,N_19048,N_19079);
xor U19358 (N_19358,N_19024,N_19161);
nand U19359 (N_19359,N_19173,N_19135);
xor U19360 (N_19360,N_19110,N_19000);
xnor U19361 (N_19361,N_19088,N_19241);
and U19362 (N_19362,N_19025,N_19209);
nor U19363 (N_19363,N_19221,N_19148);
or U19364 (N_19364,N_19069,N_19013);
and U19365 (N_19365,N_19001,N_19143);
or U19366 (N_19366,N_19065,N_19202);
or U19367 (N_19367,N_19118,N_19043);
and U19368 (N_19368,N_19038,N_19235);
xor U19369 (N_19369,N_19040,N_19009);
and U19370 (N_19370,N_19190,N_19037);
and U19371 (N_19371,N_19247,N_19232);
and U19372 (N_19372,N_19238,N_19022);
nor U19373 (N_19373,N_19045,N_19150);
nor U19374 (N_19374,N_19189,N_19184);
nor U19375 (N_19375,N_19220,N_19054);
nand U19376 (N_19376,N_19045,N_19235);
nand U19377 (N_19377,N_19211,N_19086);
nand U19378 (N_19378,N_19066,N_19247);
or U19379 (N_19379,N_19115,N_19077);
xor U19380 (N_19380,N_19244,N_19097);
nor U19381 (N_19381,N_19156,N_19229);
or U19382 (N_19382,N_19039,N_19089);
nand U19383 (N_19383,N_19096,N_19156);
xor U19384 (N_19384,N_19197,N_19224);
and U19385 (N_19385,N_19180,N_19066);
or U19386 (N_19386,N_19141,N_19117);
nor U19387 (N_19387,N_19024,N_19184);
nand U19388 (N_19388,N_19227,N_19243);
or U19389 (N_19389,N_19044,N_19063);
nor U19390 (N_19390,N_19065,N_19218);
xor U19391 (N_19391,N_19109,N_19155);
xnor U19392 (N_19392,N_19108,N_19200);
and U19393 (N_19393,N_19230,N_19241);
or U19394 (N_19394,N_19183,N_19205);
nor U19395 (N_19395,N_19081,N_19185);
and U19396 (N_19396,N_19029,N_19083);
nand U19397 (N_19397,N_19162,N_19174);
or U19398 (N_19398,N_19026,N_19117);
nand U19399 (N_19399,N_19024,N_19145);
and U19400 (N_19400,N_19023,N_19198);
and U19401 (N_19401,N_19052,N_19206);
nor U19402 (N_19402,N_19214,N_19009);
and U19403 (N_19403,N_19044,N_19242);
and U19404 (N_19404,N_19130,N_19056);
nor U19405 (N_19405,N_19001,N_19004);
and U19406 (N_19406,N_19214,N_19126);
or U19407 (N_19407,N_19013,N_19034);
nand U19408 (N_19408,N_19051,N_19009);
nand U19409 (N_19409,N_19002,N_19184);
xnor U19410 (N_19410,N_19206,N_19243);
xor U19411 (N_19411,N_19077,N_19189);
xnor U19412 (N_19412,N_19088,N_19177);
nand U19413 (N_19413,N_19021,N_19142);
xnor U19414 (N_19414,N_19127,N_19012);
nand U19415 (N_19415,N_19207,N_19034);
xor U19416 (N_19416,N_19125,N_19208);
nor U19417 (N_19417,N_19166,N_19045);
nand U19418 (N_19418,N_19057,N_19077);
nand U19419 (N_19419,N_19229,N_19116);
nor U19420 (N_19420,N_19015,N_19196);
nand U19421 (N_19421,N_19088,N_19024);
or U19422 (N_19422,N_19177,N_19167);
and U19423 (N_19423,N_19113,N_19083);
nor U19424 (N_19424,N_19245,N_19212);
nand U19425 (N_19425,N_19026,N_19241);
and U19426 (N_19426,N_19240,N_19011);
or U19427 (N_19427,N_19060,N_19105);
xnor U19428 (N_19428,N_19048,N_19050);
or U19429 (N_19429,N_19195,N_19215);
nor U19430 (N_19430,N_19058,N_19137);
nor U19431 (N_19431,N_19101,N_19225);
or U19432 (N_19432,N_19082,N_19241);
nor U19433 (N_19433,N_19162,N_19062);
xnor U19434 (N_19434,N_19045,N_19159);
nand U19435 (N_19435,N_19096,N_19069);
and U19436 (N_19436,N_19055,N_19077);
and U19437 (N_19437,N_19006,N_19136);
nand U19438 (N_19438,N_19083,N_19145);
and U19439 (N_19439,N_19007,N_19110);
or U19440 (N_19440,N_19004,N_19157);
nand U19441 (N_19441,N_19196,N_19213);
or U19442 (N_19442,N_19176,N_19175);
nand U19443 (N_19443,N_19126,N_19051);
nand U19444 (N_19444,N_19178,N_19071);
xnor U19445 (N_19445,N_19178,N_19072);
or U19446 (N_19446,N_19033,N_19058);
and U19447 (N_19447,N_19238,N_19171);
nor U19448 (N_19448,N_19178,N_19191);
and U19449 (N_19449,N_19015,N_19158);
xnor U19450 (N_19450,N_19035,N_19013);
xor U19451 (N_19451,N_19025,N_19085);
xnor U19452 (N_19452,N_19211,N_19206);
nor U19453 (N_19453,N_19011,N_19212);
nor U19454 (N_19454,N_19080,N_19120);
and U19455 (N_19455,N_19151,N_19110);
or U19456 (N_19456,N_19220,N_19026);
or U19457 (N_19457,N_19173,N_19191);
xor U19458 (N_19458,N_19185,N_19206);
and U19459 (N_19459,N_19120,N_19222);
nand U19460 (N_19460,N_19092,N_19002);
or U19461 (N_19461,N_19158,N_19033);
or U19462 (N_19462,N_19113,N_19191);
nor U19463 (N_19463,N_19194,N_19171);
or U19464 (N_19464,N_19174,N_19176);
xor U19465 (N_19465,N_19227,N_19138);
xor U19466 (N_19466,N_19189,N_19245);
xnor U19467 (N_19467,N_19182,N_19063);
nand U19468 (N_19468,N_19172,N_19064);
or U19469 (N_19469,N_19195,N_19050);
or U19470 (N_19470,N_19132,N_19155);
or U19471 (N_19471,N_19008,N_19053);
xor U19472 (N_19472,N_19225,N_19131);
xnor U19473 (N_19473,N_19071,N_19008);
and U19474 (N_19474,N_19139,N_19184);
or U19475 (N_19475,N_19175,N_19177);
nand U19476 (N_19476,N_19004,N_19014);
and U19477 (N_19477,N_19040,N_19007);
and U19478 (N_19478,N_19035,N_19231);
or U19479 (N_19479,N_19072,N_19025);
and U19480 (N_19480,N_19226,N_19063);
and U19481 (N_19481,N_19164,N_19219);
nand U19482 (N_19482,N_19232,N_19121);
or U19483 (N_19483,N_19184,N_19128);
and U19484 (N_19484,N_19189,N_19230);
xor U19485 (N_19485,N_19216,N_19108);
and U19486 (N_19486,N_19104,N_19163);
xor U19487 (N_19487,N_19161,N_19148);
and U19488 (N_19488,N_19110,N_19107);
or U19489 (N_19489,N_19059,N_19242);
or U19490 (N_19490,N_19247,N_19069);
xnor U19491 (N_19491,N_19208,N_19108);
and U19492 (N_19492,N_19202,N_19053);
xnor U19493 (N_19493,N_19061,N_19023);
and U19494 (N_19494,N_19052,N_19169);
xnor U19495 (N_19495,N_19054,N_19010);
nor U19496 (N_19496,N_19086,N_19057);
and U19497 (N_19497,N_19000,N_19220);
xnor U19498 (N_19498,N_19108,N_19093);
nand U19499 (N_19499,N_19185,N_19116);
or U19500 (N_19500,N_19331,N_19265);
xnor U19501 (N_19501,N_19372,N_19389);
nor U19502 (N_19502,N_19479,N_19374);
and U19503 (N_19503,N_19392,N_19493);
nand U19504 (N_19504,N_19343,N_19406);
xor U19505 (N_19505,N_19390,N_19395);
and U19506 (N_19506,N_19269,N_19301);
or U19507 (N_19507,N_19413,N_19358);
and U19508 (N_19508,N_19405,N_19329);
xor U19509 (N_19509,N_19397,N_19283);
or U19510 (N_19510,N_19286,N_19289);
nor U19511 (N_19511,N_19474,N_19279);
nand U19512 (N_19512,N_19380,N_19250);
nand U19513 (N_19513,N_19381,N_19398);
xor U19514 (N_19514,N_19436,N_19464);
nor U19515 (N_19515,N_19432,N_19400);
nand U19516 (N_19516,N_19257,N_19290);
or U19517 (N_19517,N_19480,N_19498);
xor U19518 (N_19518,N_19363,N_19385);
nand U19519 (N_19519,N_19354,N_19259);
xor U19520 (N_19520,N_19294,N_19359);
xor U19521 (N_19521,N_19316,N_19458);
nand U19522 (N_19522,N_19306,N_19333);
nor U19523 (N_19523,N_19293,N_19414);
or U19524 (N_19524,N_19328,N_19373);
nor U19525 (N_19525,N_19460,N_19394);
xor U19526 (N_19526,N_19303,N_19305);
nand U19527 (N_19527,N_19443,N_19351);
or U19528 (N_19528,N_19320,N_19318);
nor U19529 (N_19529,N_19272,N_19496);
or U19530 (N_19530,N_19456,N_19492);
or U19531 (N_19531,N_19285,N_19455);
nor U19532 (N_19532,N_19391,N_19384);
xor U19533 (N_19533,N_19417,N_19271);
nor U19534 (N_19534,N_19468,N_19326);
or U19535 (N_19535,N_19368,N_19416);
or U19536 (N_19536,N_19438,N_19304);
and U19537 (N_19537,N_19298,N_19415);
or U19538 (N_19538,N_19495,N_19253);
nor U19539 (N_19539,N_19422,N_19487);
or U19540 (N_19540,N_19309,N_19434);
nor U19541 (N_19541,N_19375,N_19457);
and U19542 (N_19542,N_19267,N_19335);
nand U19543 (N_19543,N_19378,N_19428);
nor U19544 (N_19544,N_19486,N_19332);
and U19545 (N_19545,N_19476,N_19449);
or U19546 (N_19546,N_19348,N_19256);
and U19547 (N_19547,N_19383,N_19497);
nand U19548 (N_19548,N_19308,N_19323);
xnor U19549 (N_19549,N_19403,N_19297);
nor U19550 (N_19550,N_19361,N_19282);
nand U19551 (N_19551,N_19313,N_19437);
nor U19552 (N_19552,N_19302,N_19345);
xnor U19553 (N_19553,N_19388,N_19469);
xor U19554 (N_19554,N_19360,N_19273);
xor U19555 (N_19555,N_19441,N_19473);
and U19556 (N_19556,N_19451,N_19288);
nor U19557 (N_19557,N_19393,N_19412);
or U19558 (N_19558,N_19430,N_19296);
nor U19559 (N_19559,N_19338,N_19418);
and U19560 (N_19560,N_19263,N_19357);
or U19561 (N_19561,N_19252,N_19467);
nor U19562 (N_19562,N_19340,N_19324);
and U19563 (N_19563,N_19491,N_19404);
nand U19564 (N_19564,N_19268,N_19330);
nand U19565 (N_19565,N_19299,N_19355);
nor U19566 (N_19566,N_19494,N_19466);
and U19567 (N_19567,N_19260,N_19447);
or U19568 (N_19568,N_19435,N_19445);
or U19569 (N_19569,N_19261,N_19454);
and U19570 (N_19570,N_19488,N_19425);
nor U19571 (N_19571,N_19295,N_19342);
nand U19572 (N_19572,N_19459,N_19353);
nor U19573 (N_19573,N_19386,N_19266);
xnor U19574 (N_19574,N_19376,N_19419);
xor U19575 (N_19575,N_19367,N_19281);
and U19576 (N_19576,N_19490,N_19287);
and U19577 (N_19577,N_19423,N_19364);
nor U19578 (N_19578,N_19396,N_19321);
nor U19579 (N_19579,N_19300,N_19485);
nand U19580 (N_19580,N_19349,N_19408);
xnor U19581 (N_19581,N_19429,N_19278);
nand U19582 (N_19582,N_19379,N_19475);
nand U19583 (N_19583,N_19387,N_19433);
xor U19584 (N_19584,N_19382,N_19312);
nand U19585 (N_19585,N_19276,N_19410);
nor U19586 (N_19586,N_19284,N_19452);
or U19587 (N_19587,N_19270,N_19366);
nand U19588 (N_19588,N_19325,N_19499);
or U19589 (N_19589,N_19489,N_19439);
and U19590 (N_19590,N_19370,N_19471);
and U19591 (N_19591,N_19450,N_19377);
nand U19592 (N_19592,N_19448,N_19356);
xnor U19593 (N_19593,N_19258,N_19350);
nand U19594 (N_19594,N_19319,N_19346);
xnor U19595 (N_19595,N_19472,N_19334);
nor U19596 (N_19596,N_19264,N_19255);
nor U19597 (N_19597,N_19402,N_19327);
nor U19598 (N_19598,N_19341,N_19462);
and U19599 (N_19599,N_19274,N_19291);
nor U19600 (N_19600,N_19482,N_19369);
xnor U19601 (N_19601,N_19315,N_19275);
nor U19602 (N_19602,N_19277,N_19292);
nor U19603 (N_19603,N_19431,N_19322);
nand U19604 (N_19604,N_19401,N_19280);
nor U19605 (N_19605,N_19477,N_19424);
nor U19606 (N_19606,N_19254,N_19465);
nor U19607 (N_19607,N_19446,N_19420);
nor U19608 (N_19608,N_19310,N_19371);
nand U19609 (N_19609,N_19314,N_19409);
or U19610 (N_19610,N_19365,N_19453);
and U19611 (N_19611,N_19442,N_19311);
xor U19612 (N_19612,N_19427,N_19251);
nor U19613 (N_19613,N_19399,N_19407);
nand U19614 (N_19614,N_19470,N_19484);
xnor U19615 (N_19615,N_19352,N_19362);
and U19616 (N_19616,N_19421,N_19426);
xor U19617 (N_19617,N_19262,N_19307);
or U19618 (N_19618,N_19440,N_19461);
and U19619 (N_19619,N_19347,N_19483);
xnor U19620 (N_19620,N_19317,N_19444);
and U19621 (N_19621,N_19336,N_19344);
xor U19622 (N_19622,N_19337,N_19478);
nand U19623 (N_19623,N_19463,N_19481);
nand U19624 (N_19624,N_19411,N_19339);
nor U19625 (N_19625,N_19424,N_19457);
xnor U19626 (N_19626,N_19407,N_19383);
nand U19627 (N_19627,N_19270,N_19476);
and U19628 (N_19628,N_19369,N_19465);
or U19629 (N_19629,N_19350,N_19256);
or U19630 (N_19630,N_19476,N_19428);
and U19631 (N_19631,N_19392,N_19421);
and U19632 (N_19632,N_19366,N_19396);
nand U19633 (N_19633,N_19438,N_19373);
or U19634 (N_19634,N_19466,N_19386);
nand U19635 (N_19635,N_19396,N_19399);
and U19636 (N_19636,N_19276,N_19365);
nand U19637 (N_19637,N_19483,N_19472);
or U19638 (N_19638,N_19462,N_19395);
xor U19639 (N_19639,N_19301,N_19440);
and U19640 (N_19640,N_19374,N_19493);
and U19641 (N_19641,N_19437,N_19412);
nor U19642 (N_19642,N_19303,N_19317);
xor U19643 (N_19643,N_19300,N_19421);
xor U19644 (N_19644,N_19455,N_19418);
xor U19645 (N_19645,N_19334,N_19378);
nor U19646 (N_19646,N_19323,N_19427);
nand U19647 (N_19647,N_19449,N_19493);
or U19648 (N_19648,N_19289,N_19414);
nor U19649 (N_19649,N_19445,N_19393);
nand U19650 (N_19650,N_19453,N_19313);
xor U19651 (N_19651,N_19359,N_19252);
and U19652 (N_19652,N_19455,N_19315);
nor U19653 (N_19653,N_19468,N_19448);
or U19654 (N_19654,N_19360,N_19435);
nor U19655 (N_19655,N_19414,N_19438);
and U19656 (N_19656,N_19256,N_19421);
nor U19657 (N_19657,N_19495,N_19327);
nor U19658 (N_19658,N_19357,N_19366);
nor U19659 (N_19659,N_19279,N_19378);
nand U19660 (N_19660,N_19361,N_19433);
nand U19661 (N_19661,N_19340,N_19257);
or U19662 (N_19662,N_19458,N_19467);
xnor U19663 (N_19663,N_19421,N_19266);
and U19664 (N_19664,N_19354,N_19463);
nand U19665 (N_19665,N_19443,N_19470);
nand U19666 (N_19666,N_19312,N_19401);
nor U19667 (N_19667,N_19474,N_19440);
or U19668 (N_19668,N_19251,N_19433);
xnor U19669 (N_19669,N_19435,N_19312);
xor U19670 (N_19670,N_19324,N_19384);
xor U19671 (N_19671,N_19452,N_19487);
nand U19672 (N_19672,N_19261,N_19483);
nor U19673 (N_19673,N_19422,N_19333);
xor U19674 (N_19674,N_19277,N_19353);
nor U19675 (N_19675,N_19488,N_19498);
xnor U19676 (N_19676,N_19322,N_19410);
nand U19677 (N_19677,N_19424,N_19470);
nor U19678 (N_19678,N_19316,N_19272);
and U19679 (N_19679,N_19319,N_19422);
and U19680 (N_19680,N_19324,N_19378);
or U19681 (N_19681,N_19470,N_19353);
or U19682 (N_19682,N_19354,N_19435);
nand U19683 (N_19683,N_19336,N_19369);
or U19684 (N_19684,N_19404,N_19444);
nor U19685 (N_19685,N_19334,N_19296);
and U19686 (N_19686,N_19495,N_19411);
xnor U19687 (N_19687,N_19303,N_19360);
xnor U19688 (N_19688,N_19354,N_19369);
and U19689 (N_19689,N_19256,N_19363);
nor U19690 (N_19690,N_19434,N_19449);
xor U19691 (N_19691,N_19401,N_19266);
nor U19692 (N_19692,N_19285,N_19443);
or U19693 (N_19693,N_19381,N_19325);
nand U19694 (N_19694,N_19293,N_19410);
and U19695 (N_19695,N_19455,N_19354);
or U19696 (N_19696,N_19437,N_19429);
or U19697 (N_19697,N_19365,N_19430);
and U19698 (N_19698,N_19472,N_19373);
or U19699 (N_19699,N_19491,N_19378);
and U19700 (N_19700,N_19449,N_19395);
xnor U19701 (N_19701,N_19462,N_19455);
and U19702 (N_19702,N_19262,N_19270);
xnor U19703 (N_19703,N_19311,N_19287);
nand U19704 (N_19704,N_19332,N_19437);
and U19705 (N_19705,N_19255,N_19312);
nor U19706 (N_19706,N_19354,N_19371);
nor U19707 (N_19707,N_19301,N_19451);
nor U19708 (N_19708,N_19485,N_19282);
and U19709 (N_19709,N_19381,N_19272);
xor U19710 (N_19710,N_19265,N_19461);
nor U19711 (N_19711,N_19296,N_19367);
nor U19712 (N_19712,N_19326,N_19369);
nor U19713 (N_19713,N_19447,N_19332);
nand U19714 (N_19714,N_19483,N_19376);
nand U19715 (N_19715,N_19397,N_19383);
xnor U19716 (N_19716,N_19437,N_19275);
or U19717 (N_19717,N_19251,N_19466);
nand U19718 (N_19718,N_19453,N_19498);
and U19719 (N_19719,N_19417,N_19416);
nand U19720 (N_19720,N_19407,N_19254);
or U19721 (N_19721,N_19254,N_19252);
and U19722 (N_19722,N_19341,N_19480);
and U19723 (N_19723,N_19313,N_19256);
nand U19724 (N_19724,N_19466,N_19275);
xnor U19725 (N_19725,N_19362,N_19479);
nand U19726 (N_19726,N_19459,N_19373);
nand U19727 (N_19727,N_19304,N_19463);
or U19728 (N_19728,N_19319,N_19270);
xor U19729 (N_19729,N_19416,N_19258);
nand U19730 (N_19730,N_19310,N_19262);
nor U19731 (N_19731,N_19469,N_19439);
xor U19732 (N_19732,N_19397,N_19300);
nand U19733 (N_19733,N_19365,N_19275);
nor U19734 (N_19734,N_19386,N_19492);
nand U19735 (N_19735,N_19456,N_19375);
xor U19736 (N_19736,N_19429,N_19454);
xor U19737 (N_19737,N_19399,N_19282);
and U19738 (N_19738,N_19448,N_19329);
or U19739 (N_19739,N_19273,N_19492);
or U19740 (N_19740,N_19417,N_19405);
nor U19741 (N_19741,N_19481,N_19265);
or U19742 (N_19742,N_19470,N_19250);
nor U19743 (N_19743,N_19387,N_19265);
and U19744 (N_19744,N_19274,N_19265);
and U19745 (N_19745,N_19262,N_19281);
xor U19746 (N_19746,N_19400,N_19409);
nor U19747 (N_19747,N_19374,N_19343);
nand U19748 (N_19748,N_19311,N_19398);
nor U19749 (N_19749,N_19269,N_19282);
and U19750 (N_19750,N_19501,N_19518);
or U19751 (N_19751,N_19589,N_19622);
or U19752 (N_19752,N_19540,N_19742);
xor U19753 (N_19753,N_19709,N_19646);
or U19754 (N_19754,N_19548,N_19541);
or U19755 (N_19755,N_19650,N_19537);
xor U19756 (N_19756,N_19712,N_19556);
xnor U19757 (N_19757,N_19619,N_19656);
nor U19758 (N_19758,N_19711,N_19603);
and U19759 (N_19759,N_19515,N_19608);
and U19760 (N_19760,N_19555,N_19660);
xnor U19761 (N_19761,N_19610,N_19734);
nor U19762 (N_19762,N_19591,N_19704);
and U19763 (N_19763,N_19698,N_19701);
or U19764 (N_19764,N_19651,N_19631);
nand U19765 (N_19765,N_19636,N_19719);
xnor U19766 (N_19766,N_19749,N_19569);
nand U19767 (N_19767,N_19510,N_19658);
nor U19768 (N_19768,N_19578,N_19668);
nand U19769 (N_19769,N_19640,N_19615);
and U19770 (N_19770,N_19652,N_19692);
and U19771 (N_19771,N_19593,N_19679);
nor U19772 (N_19772,N_19581,N_19544);
nand U19773 (N_19773,N_19624,N_19545);
and U19774 (N_19774,N_19592,N_19504);
nand U19775 (N_19775,N_19635,N_19509);
xnor U19776 (N_19776,N_19604,N_19746);
xnor U19777 (N_19777,N_19655,N_19572);
nand U19778 (N_19778,N_19745,N_19525);
or U19779 (N_19779,N_19554,N_19715);
xor U19780 (N_19780,N_19519,N_19539);
xor U19781 (N_19781,N_19620,N_19690);
and U19782 (N_19782,N_19649,N_19594);
nor U19783 (N_19783,N_19676,N_19667);
or U19784 (N_19784,N_19687,N_19724);
and U19785 (N_19785,N_19577,N_19664);
xnor U19786 (N_19786,N_19527,N_19741);
nand U19787 (N_19787,N_19549,N_19670);
xnor U19788 (N_19788,N_19506,N_19534);
xnor U19789 (N_19789,N_19740,N_19576);
nand U19790 (N_19790,N_19588,N_19623);
and U19791 (N_19791,N_19643,N_19607);
nand U19792 (N_19792,N_19672,N_19561);
and U19793 (N_19793,N_19703,N_19505);
or U19794 (N_19794,N_19552,N_19503);
and U19795 (N_19795,N_19508,N_19606);
xor U19796 (N_19796,N_19562,N_19553);
and U19797 (N_19797,N_19700,N_19706);
and U19798 (N_19798,N_19677,N_19617);
nand U19799 (N_19799,N_19579,N_19626);
nand U19800 (N_19800,N_19521,N_19637);
and U19801 (N_19801,N_19502,N_19653);
or U19802 (N_19802,N_19601,N_19714);
xor U19803 (N_19803,N_19736,N_19543);
nor U19804 (N_19804,N_19682,N_19696);
nor U19805 (N_19805,N_19586,N_19523);
nor U19806 (N_19806,N_19748,N_19547);
or U19807 (N_19807,N_19718,N_19570);
xnor U19808 (N_19808,N_19633,N_19705);
or U19809 (N_19809,N_19590,N_19729);
xor U19810 (N_19810,N_19744,N_19516);
or U19811 (N_19811,N_19699,N_19550);
and U19812 (N_19812,N_19730,N_19693);
and U19813 (N_19813,N_19738,N_19512);
nand U19814 (N_19814,N_19708,N_19595);
or U19815 (N_19815,N_19725,N_19680);
or U19816 (N_19816,N_19684,N_19683);
or U19817 (N_19817,N_19691,N_19551);
nor U19818 (N_19818,N_19634,N_19565);
or U19819 (N_19819,N_19574,N_19732);
or U19820 (N_19820,N_19612,N_19728);
and U19821 (N_19821,N_19743,N_19710);
and U19822 (N_19822,N_19522,N_19566);
and U19823 (N_19823,N_19618,N_19722);
nand U19824 (N_19824,N_19674,N_19507);
nand U19825 (N_19825,N_19582,N_19542);
nand U19826 (N_19826,N_19611,N_19597);
nand U19827 (N_19827,N_19675,N_19697);
nand U19828 (N_19828,N_19694,N_19678);
nor U19829 (N_19829,N_19535,N_19560);
and U19830 (N_19830,N_19721,N_19669);
xor U19831 (N_19831,N_19557,N_19530);
nor U19832 (N_19832,N_19531,N_19702);
or U19833 (N_19833,N_19575,N_19647);
and U19834 (N_19834,N_19644,N_19642);
nand U19835 (N_19835,N_19733,N_19673);
xor U19836 (N_19836,N_19529,N_19671);
nand U19837 (N_19837,N_19666,N_19723);
nand U19838 (N_19838,N_19632,N_19686);
nand U19839 (N_19839,N_19726,N_19716);
and U19840 (N_19840,N_19641,N_19571);
and U19841 (N_19841,N_19681,N_19609);
or U19842 (N_19842,N_19524,N_19665);
nand U19843 (N_19843,N_19526,N_19583);
nor U19844 (N_19844,N_19513,N_19727);
xor U19845 (N_19845,N_19645,N_19599);
nor U19846 (N_19846,N_19500,N_19639);
xor U19847 (N_19847,N_19585,N_19707);
xor U19848 (N_19848,N_19532,N_19628);
and U19849 (N_19849,N_19567,N_19685);
and U19850 (N_19850,N_19514,N_19528);
nand U19851 (N_19851,N_19735,N_19538);
and U19852 (N_19852,N_19747,N_19638);
nand U19853 (N_19853,N_19616,N_19661);
and U19854 (N_19854,N_19559,N_19659);
and U19855 (N_19855,N_19605,N_19596);
nor U19856 (N_19856,N_19717,N_19573);
or U19857 (N_19857,N_19689,N_19657);
nor U19858 (N_19858,N_19731,N_19739);
nor U19859 (N_19859,N_19713,N_19630);
or U19860 (N_19860,N_19520,N_19598);
and U19861 (N_19861,N_19648,N_19533);
xnor U19862 (N_19862,N_19558,N_19627);
and U19863 (N_19863,N_19621,N_19517);
xor U19864 (N_19864,N_19587,N_19564);
xor U19865 (N_19865,N_19720,N_19580);
xnor U19866 (N_19866,N_19602,N_19546);
xor U19867 (N_19867,N_19600,N_19654);
nand U19868 (N_19868,N_19629,N_19614);
and U19869 (N_19869,N_19613,N_19695);
and U19870 (N_19870,N_19536,N_19511);
or U19871 (N_19871,N_19568,N_19688);
nor U19872 (N_19872,N_19663,N_19625);
nand U19873 (N_19873,N_19584,N_19737);
nor U19874 (N_19874,N_19563,N_19662);
and U19875 (N_19875,N_19733,N_19541);
nand U19876 (N_19876,N_19718,N_19636);
xnor U19877 (N_19877,N_19705,N_19630);
or U19878 (N_19878,N_19558,N_19730);
or U19879 (N_19879,N_19507,N_19659);
nand U19880 (N_19880,N_19665,N_19719);
nand U19881 (N_19881,N_19559,N_19542);
xor U19882 (N_19882,N_19648,N_19732);
and U19883 (N_19883,N_19538,N_19617);
or U19884 (N_19884,N_19628,N_19618);
or U19885 (N_19885,N_19711,N_19700);
and U19886 (N_19886,N_19642,N_19597);
nand U19887 (N_19887,N_19551,N_19616);
nand U19888 (N_19888,N_19531,N_19513);
nand U19889 (N_19889,N_19730,N_19620);
and U19890 (N_19890,N_19640,N_19531);
and U19891 (N_19891,N_19726,N_19585);
and U19892 (N_19892,N_19652,N_19598);
nand U19893 (N_19893,N_19567,N_19636);
nor U19894 (N_19894,N_19600,N_19706);
nand U19895 (N_19895,N_19557,N_19703);
or U19896 (N_19896,N_19614,N_19684);
nor U19897 (N_19897,N_19684,N_19743);
xor U19898 (N_19898,N_19535,N_19534);
and U19899 (N_19899,N_19627,N_19525);
or U19900 (N_19900,N_19557,N_19579);
nor U19901 (N_19901,N_19558,N_19743);
and U19902 (N_19902,N_19580,N_19638);
and U19903 (N_19903,N_19741,N_19711);
or U19904 (N_19904,N_19522,N_19701);
xnor U19905 (N_19905,N_19735,N_19695);
xor U19906 (N_19906,N_19582,N_19566);
or U19907 (N_19907,N_19708,N_19656);
nand U19908 (N_19908,N_19606,N_19730);
or U19909 (N_19909,N_19584,N_19576);
nor U19910 (N_19910,N_19587,N_19557);
and U19911 (N_19911,N_19725,N_19599);
nand U19912 (N_19912,N_19701,N_19520);
nor U19913 (N_19913,N_19622,N_19581);
nand U19914 (N_19914,N_19585,N_19694);
xor U19915 (N_19915,N_19584,N_19517);
nand U19916 (N_19916,N_19685,N_19523);
or U19917 (N_19917,N_19521,N_19575);
and U19918 (N_19918,N_19744,N_19739);
nand U19919 (N_19919,N_19572,N_19660);
nand U19920 (N_19920,N_19738,N_19582);
xor U19921 (N_19921,N_19559,N_19746);
and U19922 (N_19922,N_19586,N_19731);
nand U19923 (N_19923,N_19527,N_19589);
nor U19924 (N_19924,N_19535,N_19675);
or U19925 (N_19925,N_19731,N_19676);
nor U19926 (N_19926,N_19721,N_19501);
and U19927 (N_19927,N_19614,N_19679);
or U19928 (N_19928,N_19724,N_19726);
nor U19929 (N_19929,N_19747,N_19714);
nand U19930 (N_19930,N_19694,N_19516);
nor U19931 (N_19931,N_19710,N_19714);
or U19932 (N_19932,N_19646,N_19543);
and U19933 (N_19933,N_19606,N_19505);
nand U19934 (N_19934,N_19617,N_19606);
nor U19935 (N_19935,N_19534,N_19740);
and U19936 (N_19936,N_19651,N_19563);
nand U19937 (N_19937,N_19504,N_19717);
xnor U19938 (N_19938,N_19595,N_19533);
nor U19939 (N_19939,N_19608,N_19534);
and U19940 (N_19940,N_19626,N_19659);
nor U19941 (N_19941,N_19552,N_19539);
nor U19942 (N_19942,N_19651,N_19686);
xnor U19943 (N_19943,N_19705,N_19723);
or U19944 (N_19944,N_19598,N_19544);
xnor U19945 (N_19945,N_19594,N_19581);
nor U19946 (N_19946,N_19594,N_19517);
nand U19947 (N_19947,N_19701,N_19662);
nand U19948 (N_19948,N_19735,N_19577);
nor U19949 (N_19949,N_19647,N_19551);
nand U19950 (N_19950,N_19680,N_19561);
xnor U19951 (N_19951,N_19512,N_19586);
nor U19952 (N_19952,N_19601,N_19528);
xor U19953 (N_19953,N_19624,N_19706);
nand U19954 (N_19954,N_19689,N_19651);
xor U19955 (N_19955,N_19730,N_19536);
nor U19956 (N_19956,N_19641,N_19522);
and U19957 (N_19957,N_19582,N_19626);
and U19958 (N_19958,N_19506,N_19698);
nand U19959 (N_19959,N_19654,N_19592);
or U19960 (N_19960,N_19691,N_19534);
xnor U19961 (N_19961,N_19640,N_19638);
xnor U19962 (N_19962,N_19729,N_19511);
and U19963 (N_19963,N_19612,N_19562);
xor U19964 (N_19964,N_19713,N_19528);
nor U19965 (N_19965,N_19631,N_19527);
nand U19966 (N_19966,N_19646,N_19707);
or U19967 (N_19967,N_19688,N_19544);
nor U19968 (N_19968,N_19583,N_19615);
and U19969 (N_19969,N_19522,N_19642);
xnor U19970 (N_19970,N_19561,N_19515);
xor U19971 (N_19971,N_19731,N_19507);
or U19972 (N_19972,N_19668,N_19710);
nor U19973 (N_19973,N_19635,N_19562);
nand U19974 (N_19974,N_19605,N_19684);
xnor U19975 (N_19975,N_19736,N_19650);
nor U19976 (N_19976,N_19513,N_19652);
and U19977 (N_19977,N_19717,N_19629);
nand U19978 (N_19978,N_19569,N_19597);
and U19979 (N_19979,N_19667,N_19708);
or U19980 (N_19980,N_19584,N_19738);
nand U19981 (N_19981,N_19522,N_19685);
and U19982 (N_19982,N_19529,N_19675);
xor U19983 (N_19983,N_19695,N_19728);
or U19984 (N_19984,N_19650,N_19665);
or U19985 (N_19985,N_19709,N_19694);
or U19986 (N_19986,N_19536,N_19653);
xnor U19987 (N_19987,N_19572,N_19672);
and U19988 (N_19988,N_19697,N_19624);
xor U19989 (N_19989,N_19660,N_19580);
xor U19990 (N_19990,N_19722,N_19732);
or U19991 (N_19991,N_19642,N_19613);
or U19992 (N_19992,N_19614,N_19661);
or U19993 (N_19993,N_19584,N_19554);
or U19994 (N_19994,N_19579,N_19584);
or U19995 (N_19995,N_19501,N_19505);
nand U19996 (N_19996,N_19591,N_19623);
or U19997 (N_19997,N_19611,N_19745);
or U19998 (N_19998,N_19605,N_19547);
xor U19999 (N_19999,N_19695,N_19733);
and UO_0 (O_0,N_19863,N_19922);
xnor UO_1 (O_1,N_19952,N_19993);
or UO_2 (O_2,N_19895,N_19949);
and UO_3 (O_3,N_19814,N_19780);
nor UO_4 (O_4,N_19934,N_19970);
and UO_5 (O_5,N_19824,N_19899);
or UO_6 (O_6,N_19832,N_19976);
xor UO_7 (O_7,N_19782,N_19785);
nand UO_8 (O_8,N_19916,N_19891);
xor UO_9 (O_9,N_19930,N_19790);
or UO_10 (O_10,N_19857,N_19803);
xnor UO_11 (O_11,N_19996,N_19950);
or UO_12 (O_12,N_19966,N_19858);
and UO_13 (O_13,N_19939,N_19795);
xor UO_14 (O_14,N_19909,N_19870);
xor UO_15 (O_15,N_19779,N_19771);
nor UO_16 (O_16,N_19854,N_19998);
or UO_17 (O_17,N_19750,N_19764);
nand UO_18 (O_18,N_19888,N_19936);
or UO_19 (O_19,N_19894,N_19864);
and UO_20 (O_20,N_19942,N_19969);
nor UO_21 (O_21,N_19752,N_19827);
nand UO_22 (O_22,N_19921,N_19849);
or UO_23 (O_23,N_19751,N_19826);
or UO_24 (O_24,N_19935,N_19829);
and UO_25 (O_25,N_19890,N_19997);
nand UO_26 (O_26,N_19992,N_19798);
nor UO_27 (O_27,N_19962,N_19974);
or UO_28 (O_28,N_19940,N_19768);
nor UO_29 (O_29,N_19817,N_19906);
nor UO_30 (O_30,N_19926,N_19758);
nand UO_31 (O_31,N_19905,N_19839);
nand UO_32 (O_32,N_19884,N_19968);
nor UO_33 (O_33,N_19965,N_19765);
or UO_34 (O_34,N_19871,N_19853);
xnor UO_35 (O_35,N_19873,N_19862);
nand UO_36 (O_36,N_19920,N_19860);
nor UO_37 (O_37,N_19914,N_19800);
or UO_38 (O_38,N_19988,N_19772);
nand UO_39 (O_39,N_19763,N_19809);
or UO_40 (O_40,N_19842,N_19855);
nand UO_41 (O_41,N_19769,N_19818);
or UO_42 (O_42,N_19999,N_19807);
and UO_43 (O_43,N_19836,N_19980);
nor UO_44 (O_44,N_19844,N_19877);
and UO_45 (O_45,N_19897,N_19778);
or UO_46 (O_46,N_19959,N_19866);
xor UO_47 (O_47,N_19947,N_19972);
and UO_48 (O_48,N_19956,N_19835);
and UO_49 (O_49,N_19971,N_19963);
and UO_50 (O_50,N_19754,N_19874);
nor UO_51 (O_51,N_19841,N_19887);
xor UO_52 (O_52,N_19961,N_19903);
nor UO_53 (O_53,N_19912,N_19924);
or UO_54 (O_54,N_19840,N_19957);
xnor UO_55 (O_55,N_19911,N_19883);
nand UO_56 (O_56,N_19933,N_19872);
xnor UO_57 (O_57,N_19805,N_19923);
xor UO_58 (O_58,N_19901,N_19865);
or UO_59 (O_59,N_19981,N_19793);
nand UO_60 (O_60,N_19919,N_19876);
and UO_61 (O_61,N_19896,N_19989);
nor UO_62 (O_62,N_19964,N_19910);
nand UO_63 (O_63,N_19978,N_19845);
and UO_64 (O_64,N_19830,N_19918);
or UO_65 (O_65,N_19927,N_19893);
nor UO_66 (O_66,N_19789,N_19759);
xnor UO_67 (O_67,N_19928,N_19767);
nand UO_68 (O_68,N_19838,N_19848);
nor UO_69 (O_69,N_19755,N_19958);
xor UO_70 (O_70,N_19784,N_19786);
xnor UO_71 (O_71,N_19820,N_19831);
nand UO_72 (O_72,N_19879,N_19788);
xor UO_73 (O_73,N_19846,N_19889);
or UO_74 (O_74,N_19796,N_19753);
or UO_75 (O_75,N_19945,N_19794);
nor UO_76 (O_76,N_19868,N_19955);
xnor UO_77 (O_77,N_19946,N_19900);
or UO_78 (O_78,N_19878,N_19954);
nor UO_79 (O_79,N_19787,N_19932);
or UO_80 (O_80,N_19825,N_19977);
or UO_81 (O_81,N_19931,N_19856);
and UO_82 (O_82,N_19984,N_19967);
and UO_83 (O_83,N_19843,N_19881);
and UO_84 (O_84,N_19847,N_19851);
xor UO_85 (O_85,N_19761,N_19822);
nor UO_86 (O_86,N_19948,N_19762);
nand UO_87 (O_87,N_19833,N_19867);
or UO_88 (O_88,N_19917,N_19875);
xor UO_89 (O_89,N_19951,N_19783);
nor UO_90 (O_90,N_19938,N_19801);
nor UO_91 (O_91,N_19806,N_19834);
nor UO_92 (O_92,N_19915,N_19799);
xor UO_93 (O_93,N_19960,N_19797);
nor UO_94 (O_94,N_19902,N_19819);
and UO_95 (O_95,N_19975,N_19944);
and UO_96 (O_96,N_19908,N_19837);
and UO_97 (O_97,N_19812,N_19886);
xor UO_98 (O_98,N_19777,N_19773);
or UO_99 (O_99,N_19987,N_19776);
xor UO_100 (O_100,N_19990,N_19760);
xor UO_101 (O_101,N_19986,N_19811);
nor UO_102 (O_102,N_19953,N_19985);
and UO_103 (O_103,N_19816,N_19994);
and UO_104 (O_104,N_19859,N_19804);
nand UO_105 (O_105,N_19898,N_19775);
xnor UO_106 (O_106,N_19757,N_19766);
and UO_107 (O_107,N_19802,N_19943);
or UO_108 (O_108,N_19979,N_19869);
xor UO_109 (O_109,N_19885,N_19774);
xor UO_110 (O_110,N_19791,N_19823);
nand UO_111 (O_111,N_19882,N_19828);
nand UO_112 (O_112,N_19852,N_19983);
xor UO_113 (O_113,N_19913,N_19973);
or UO_114 (O_114,N_19781,N_19821);
nor UO_115 (O_115,N_19810,N_19941);
nor UO_116 (O_116,N_19892,N_19904);
nor UO_117 (O_117,N_19907,N_19982);
xnor UO_118 (O_118,N_19929,N_19815);
xor UO_119 (O_119,N_19880,N_19850);
and UO_120 (O_120,N_19808,N_19792);
nand UO_121 (O_121,N_19756,N_19925);
and UO_122 (O_122,N_19861,N_19813);
nand UO_123 (O_123,N_19770,N_19995);
nand UO_124 (O_124,N_19937,N_19991);
nand UO_125 (O_125,N_19869,N_19925);
nand UO_126 (O_126,N_19912,N_19982);
nand UO_127 (O_127,N_19831,N_19793);
and UO_128 (O_128,N_19886,N_19787);
nor UO_129 (O_129,N_19837,N_19842);
and UO_130 (O_130,N_19886,N_19878);
and UO_131 (O_131,N_19832,N_19889);
and UO_132 (O_132,N_19976,N_19765);
and UO_133 (O_133,N_19951,N_19876);
xor UO_134 (O_134,N_19792,N_19826);
and UO_135 (O_135,N_19929,N_19763);
nand UO_136 (O_136,N_19940,N_19946);
nor UO_137 (O_137,N_19790,N_19846);
nand UO_138 (O_138,N_19752,N_19868);
or UO_139 (O_139,N_19878,N_19757);
nor UO_140 (O_140,N_19792,N_19905);
or UO_141 (O_141,N_19909,N_19905);
xor UO_142 (O_142,N_19778,N_19771);
and UO_143 (O_143,N_19885,N_19762);
nor UO_144 (O_144,N_19960,N_19783);
xor UO_145 (O_145,N_19791,N_19948);
nand UO_146 (O_146,N_19824,N_19970);
and UO_147 (O_147,N_19881,N_19750);
nor UO_148 (O_148,N_19753,N_19925);
xor UO_149 (O_149,N_19838,N_19878);
nand UO_150 (O_150,N_19927,N_19821);
nor UO_151 (O_151,N_19932,N_19900);
or UO_152 (O_152,N_19844,N_19873);
and UO_153 (O_153,N_19949,N_19798);
or UO_154 (O_154,N_19817,N_19851);
or UO_155 (O_155,N_19973,N_19942);
or UO_156 (O_156,N_19999,N_19792);
or UO_157 (O_157,N_19873,N_19819);
nor UO_158 (O_158,N_19932,N_19948);
xor UO_159 (O_159,N_19997,N_19842);
xnor UO_160 (O_160,N_19947,N_19959);
and UO_161 (O_161,N_19797,N_19795);
and UO_162 (O_162,N_19960,N_19953);
nand UO_163 (O_163,N_19860,N_19804);
or UO_164 (O_164,N_19872,N_19849);
xnor UO_165 (O_165,N_19824,N_19794);
or UO_166 (O_166,N_19825,N_19917);
xor UO_167 (O_167,N_19963,N_19890);
nand UO_168 (O_168,N_19980,N_19958);
nor UO_169 (O_169,N_19986,N_19871);
and UO_170 (O_170,N_19809,N_19900);
or UO_171 (O_171,N_19892,N_19811);
or UO_172 (O_172,N_19859,N_19968);
or UO_173 (O_173,N_19773,N_19956);
or UO_174 (O_174,N_19830,N_19756);
nor UO_175 (O_175,N_19893,N_19928);
and UO_176 (O_176,N_19940,N_19776);
xnor UO_177 (O_177,N_19842,N_19796);
or UO_178 (O_178,N_19765,N_19905);
xor UO_179 (O_179,N_19763,N_19874);
or UO_180 (O_180,N_19846,N_19810);
xor UO_181 (O_181,N_19853,N_19948);
or UO_182 (O_182,N_19844,N_19789);
nor UO_183 (O_183,N_19858,N_19897);
nand UO_184 (O_184,N_19809,N_19949);
and UO_185 (O_185,N_19790,N_19939);
xnor UO_186 (O_186,N_19923,N_19931);
and UO_187 (O_187,N_19765,N_19885);
nand UO_188 (O_188,N_19995,N_19813);
or UO_189 (O_189,N_19891,N_19986);
or UO_190 (O_190,N_19826,N_19941);
xnor UO_191 (O_191,N_19892,N_19866);
and UO_192 (O_192,N_19853,N_19852);
nor UO_193 (O_193,N_19924,N_19966);
and UO_194 (O_194,N_19841,N_19943);
nor UO_195 (O_195,N_19750,N_19836);
nor UO_196 (O_196,N_19969,N_19999);
xnor UO_197 (O_197,N_19877,N_19866);
xor UO_198 (O_198,N_19848,N_19997);
xor UO_199 (O_199,N_19859,N_19928);
nand UO_200 (O_200,N_19859,N_19773);
nor UO_201 (O_201,N_19922,N_19948);
xnor UO_202 (O_202,N_19832,N_19916);
nand UO_203 (O_203,N_19760,N_19880);
nand UO_204 (O_204,N_19951,N_19974);
xor UO_205 (O_205,N_19953,N_19980);
xor UO_206 (O_206,N_19994,N_19996);
nor UO_207 (O_207,N_19930,N_19919);
nand UO_208 (O_208,N_19775,N_19890);
xor UO_209 (O_209,N_19907,N_19969);
or UO_210 (O_210,N_19957,N_19968);
and UO_211 (O_211,N_19852,N_19806);
and UO_212 (O_212,N_19830,N_19825);
nand UO_213 (O_213,N_19859,N_19827);
nor UO_214 (O_214,N_19958,N_19794);
xor UO_215 (O_215,N_19805,N_19866);
xor UO_216 (O_216,N_19973,N_19831);
xnor UO_217 (O_217,N_19798,N_19807);
xnor UO_218 (O_218,N_19799,N_19964);
nand UO_219 (O_219,N_19929,N_19946);
or UO_220 (O_220,N_19951,N_19764);
or UO_221 (O_221,N_19891,N_19923);
nand UO_222 (O_222,N_19890,N_19952);
or UO_223 (O_223,N_19956,N_19982);
nor UO_224 (O_224,N_19842,N_19808);
nor UO_225 (O_225,N_19967,N_19881);
and UO_226 (O_226,N_19945,N_19763);
and UO_227 (O_227,N_19916,N_19827);
and UO_228 (O_228,N_19852,N_19940);
or UO_229 (O_229,N_19916,N_19873);
or UO_230 (O_230,N_19935,N_19999);
nor UO_231 (O_231,N_19832,N_19750);
or UO_232 (O_232,N_19921,N_19993);
and UO_233 (O_233,N_19980,N_19830);
nor UO_234 (O_234,N_19884,N_19754);
nor UO_235 (O_235,N_19911,N_19774);
nor UO_236 (O_236,N_19849,N_19909);
nand UO_237 (O_237,N_19971,N_19875);
xor UO_238 (O_238,N_19793,N_19887);
xor UO_239 (O_239,N_19780,N_19942);
xnor UO_240 (O_240,N_19783,N_19869);
or UO_241 (O_241,N_19999,N_19885);
xnor UO_242 (O_242,N_19991,N_19765);
nor UO_243 (O_243,N_19990,N_19829);
and UO_244 (O_244,N_19825,N_19760);
nor UO_245 (O_245,N_19993,N_19787);
nand UO_246 (O_246,N_19987,N_19948);
nand UO_247 (O_247,N_19888,N_19901);
and UO_248 (O_248,N_19930,N_19854);
and UO_249 (O_249,N_19991,N_19892);
nand UO_250 (O_250,N_19896,N_19914);
nor UO_251 (O_251,N_19868,N_19913);
xor UO_252 (O_252,N_19815,N_19978);
or UO_253 (O_253,N_19753,N_19841);
nor UO_254 (O_254,N_19936,N_19927);
or UO_255 (O_255,N_19772,N_19766);
and UO_256 (O_256,N_19821,N_19793);
or UO_257 (O_257,N_19873,N_19880);
and UO_258 (O_258,N_19843,N_19829);
or UO_259 (O_259,N_19783,N_19752);
nand UO_260 (O_260,N_19783,N_19967);
and UO_261 (O_261,N_19975,N_19797);
or UO_262 (O_262,N_19952,N_19831);
nand UO_263 (O_263,N_19888,N_19751);
xnor UO_264 (O_264,N_19902,N_19870);
nor UO_265 (O_265,N_19916,N_19791);
or UO_266 (O_266,N_19761,N_19790);
xor UO_267 (O_267,N_19939,N_19869);
and UO_268 (O_268,N_19779,N_19906);
or UO_269 (O_269,N_19985,N_19914);
nand UO_270 (O_270,N_19969,N_19862);
and UO_271 (O_271,N_19924,N_19859);
and UO_272 (O_272,N_19814,N_19839);
xnor UO_273 (O_273,N_19998,N_19896);
and UO_274 (O_274,N_19879,N_19941);
and UO_275 (O_275,N_19808,N_19893);
nand UO_276 (O_276,N_19774,N_19929);
or UO_277 (O_277,N_19755,N_19872);
or UO_278 (O_278,N_19794,N_19970);
or UO_279 (O_279,N_19813,N_19868);
xor UO_280 (O_280,N_19996,N_19886);
and UO_281 (O_281,N_19988,N_19804);
nor UO_282 (O_282,N_19940,N_19785);
nand UO_283 (O_283,N_19770,N_19977);
nand UO_284 (O_284,N_19856,N_19900);
nor UO_285 (O_285,N_19915,N_19876);
and UO_286 (O_286,N_19982,N_19896);
nor UO_287 (O_287,N_19890,N_19832);
xor UO_288 (O_288,N_19982,N_19766);
xnor UO_289 (O_289,N_19815,N_19812);
or UO_290 (O_290,N_19950,N_19860);
nor UO_291 (O_291,N_19957,N_19950);
and UO_292 (O_292,N_19901,N_19936);
and UO_293 (O_293,N_19832,N_19887);
nor UO_294 (O_294,N_19920,N_19825);
nand UO_295 (O_295,N_19908,N_19899);
xor UO_296 (O_296,N_19984,N_19927);
xor UO_297 (O_297,N_19814,N_19983);
or UO_298 (O_298,N_19818,N_19952);
and UO_299 (O_299,N_19982,N_19925);
nor UO_300 (O_300,N_19879,N_19866);
nor UO_301 (O_301,N_19874,N_19927);
and UO_302 (O_302,N_19820,N_19938);
and UO_303 (O_303,N_19959,N_19863);
nand UO_304 (O_304,N_19758,N_19904);
nor UO_305 (O_305,N_19866,N_19999);
nor UO_306 (O_306,N_19942,N_19968);
nand UO_307 (O_307,N_19836,N_19819);
and UO_308 (O_308,N_19998,N_19815);
nor UO_309 (O_309,N_19756,N_19872);
nand UO_310 (O_310,N_19823,N_19754);
or UO_311 (O_311,N_19973,N_19773);
or UO_312 (O_312,N_19961,N_19841);
nand UO_313 (O_313,N_19921,N_19775);
xor UO_314 (O_314,N_19998,N_19986);
xnor UO_315 (O_315,N_19888,N_19761);
xnor UO_316 (O_316,N_19839,N_19763);
xnor UO_317 (O_317,N_19938,N_19844);
or UO_318 (O_318,N_19760,N_19805);
xnor UO_319 (O_319,N_19966,N_19825);
and UO_320 (O_320,N_19790,N_19984);
and UO_321 (O_321,N_19963,N_19966);
xor UO_322 (O_322,N_19932,N_19970);
nand UO_323 (O_323,N_19971,N_19988);
nand UO_324 (O_324,N_19994,N_19849);
and UO_325 (O_325,N_19855,N_19921);
xnor UO_326 (O_326,N_19828,N_19860);
nand UO_327 (O_327,N_19952,N_19926);
nor UO_328 (O_328,N_19988,N_19981);
xnor UO_329 (O_329,N_19914,N_19787);
and UO_330 (O_330,N_19933,N_19805);
and UO_331 (O_331,N_19821,N_19918);
nand UO_332 (O_332,N_19869,N_19787);
nor UO_333 (O_333,N_19847,N_19888);
nand UO_334 (O_334,N_19927,N_19938);
nor UO_335 (O_335,N_19803,N_19847);
and UO_336 (O_336,N_19757,N_19812);
nand UO_337 (O_337,N_19936,N_19757);
or UO_338 (O_338,N_19758,N_19865);
nand UO_339 (O_339,N_19827,N_19824);
nor UO_340 (O_340,N_19987,N_19890);
nor UO_341 (O_341,N_19890,N_19848);
nand UO_342 (O_342,N_19754,N_19762);
nor UO_343 (O_343,N_19916,N_19913);
nand UO_344 (O_344,N_19989,N_19970);
or UO_345 (O_345,N_19933,N_19802);
or UO_346 (O_346,N_19966,N_19770);
or UO_347 (O_347,N_19942,N_19832);
xnor UO_348 (O_348,N_19972,N_19767);
nor UO_349 (O_349,N_19953,N_19863);
and UO_350 (O_350,N_19759,N_19939);
nor UO_351 (O_351,N_19762,N_19916);
nor UO_352 (O_352,N_19969,N_19848);
and UO_353 (O_353,N_19929,N_19997);
xnor UO_354 (O_354,N_19818,N_19763);
nand UO_355 (O_355,N_19926,N_19960);
xnor UO_356 (O_356,N_19894,N_19907);
and UO_357 (O_357,N_19950,N_19841);
and UO_358 (O_358,N_19866,N_19881);
nor UO_359 (O_359,N_19853,N_19985);
xnor UO_360 (O_360,N_19761,N_19880);
nor UO_361 (O_361,N_19794,N_19759);
or UO_362 (O_362,N_19938,N_19848);
and UO_363 (O_363,N_19870,N_19799);
and UO_364 (O_364,N_19989,N_19763);
xnor UO_365 (O_365,N_19920,N_19813);
nand UO_366 (O_366,N_19936,N_19846);
or UO_367 (O_367,N_19939,N_19887);
nand UO_368 (O_368,N_19986,N_19878);
and UO_369 (O_369,N_19780,N_19977);
xor UO_370 (O_370,N_19883,N_19798);
or UO_371 (O_371,N_19867,N_19995);
nand UO_372 (O_372,N_19897,N_19971);
or UO_373 (O_373,N_19930,N_19992);
and UO_374 (O_374,N_19830,N_19974);
xor UO_375 (O_375,N_19937,N_19881);
and UO_376 (O_376,N_19772,N_19797);
nor UO_377 (O_377,N_19773,N_19784);
nand UO_378 (O_378,N_19752,N_19806);
xor UO_379 (O_379,N_19994,N_19756);
nor UO_380 (O_380,N_19753,N_19991);
nor UO_381 (O_381,N_19951,N_19918);
or UO_382 (O_382,N_19872,N_19942);
xnor UO_383 (O_383,N_19810,N_19798);
nor UO_384 (O_384,N_19903,N_19913);
and UO_385 (O_385,N_19843,N_19758);
and UO_386 (O_386,N_19907,N_19763);
and UO_387 (O_387,N_19854,N_19912);
nand UO_388 (O_388,N_19823,N_19997);
nand UO_389 (O_389,N_19782,N_19760);
nand UO_390 (O_390,N_19818,N_19906);
nor UO_391 (O_391,N_19757,N_19858);
and UO_392 (O_392,N_19837,N_19992);
nor UO_393 (O_393,N_19927,N_19830);
nor UO_394 (O_394,N_19907,N_19873);
nor UO_395 (O_395,N_19779,N_19785);
or UO_396 (O_396,N_19752,N_19892);
nor UO_397 (O_397,N_19807,N_19978);
or UO_398 (O_398,N_19881,N_19907);
or UO_399 (O_399,N_19771,N_19755);
nand UO_400 (O_400,N_19903,N_19957);
nor UO_401 (O_401,N_19931,N_19948);
xnor UO_402 (O_402,N_19852,N_19857);
or UO_403 (O_403,N_19822,N_19866);
and UO_404 (O_404,N_19963,N_19922);
or UO_405 (O_405,N_19894,N_19763);
or UO_406 (O_406,N_19884,N_19912);
xor UO_407 (O_407,N_19903,N_19942);
and UO_408 (O_408,N_19781,N_19857);
xnor UO_409 (O_409,N_19894,N_19934);
xnor UO_410 (O_410,N_19753,N_19912);
nor UO_411 (O_411,N_19902,N_19800);
or UO_412 (O_412,N_19862,N_19899);
or UO_413 (O_413,N_19813,N_19864);
nand UO_414 (O_414,N_19945,N_19929);
and UO_415 (O_415,N_19794,N_19881);
nor UO_416 (O_416,N_19840,N_19789);
nor UO_417 (O_417,N_19969,N_19788);
and UO_418 (O_418,N_19838,N_19982);
xnor UO_419 (O_419,N_19981,N_19898);
or UO_420 (O_420,N_19769,N_19791);
xnor UO_421 (O_421,N_19839,N_19913);
and UO_422 (O_422,N_19923,N_19826);
xor UO_423 (O_423,N_19859,N_19915);
xnor UO_424 (O_424,N_19775,N_19860);
nor UO_425 (O_425,N_19911,N_19915);
nor UO_426 (O_426,N_19841,N_19872);
xnor UO_427 (O_427,N_19856,N_19788);
and UO_428 (O_428,N_19986,N_19953);
nand UO_429 (O_429,N_19844,N_19890);
nor UO_430 (O_430,N_19753,N_19795);
or UO_431 (O_431,N_19801,N_19812);
nor UO_432 (O_432,N_19835,N_19994);
xnor UO_433 (O_433,N_19786,N_19889);
or UO_434 (O_434,N_19833,N_19909);
xor UO_435 (O_435,N_19869,N_19894);
nor UO_436 (O_436,N_19963,N_19997);
or UO_437 (O_437,N_19986,N_19932);
nand UO_438 (O_438,N_19931,N_19911);
nor UO_439 (O_439,N_19936,N_19796);
or UO_440 (O_440,N_19798,N_19799);
xor UO_441 (O_441,N_19999,N_19759);
nor UO_442 (O_442,N_19863,N_19753);
nand UO_443 (O_443,N_19770,N_19951);
and UO_444 (O_444,N_19918,N_19892);
or UO_445 (O_445,N_19988,N_19761);
xnor UO_446 (O_446,N_19753,N_19977);
xnor UO_447 (O_447,N_19848,N_19798);
xor UO_448 (O_448,N_19922,N_19779);
nor UO_449 (O_449,N_19962,N_19856);
nand UO_450 (O_450,N_19786,N_19864);
or UO_451 (O_451,N_19874,N_19813);
xnor UO_452 (O_452,N_19943,N_19906);
xnor UO_453 (O_453,N_19796,N_19901);
and UO_454 (O_454,N_19869,N_19981);
nand UO_455 (O_455,N_19853,N_19942);
xnor UO_456 (O_456,N_19929,N_19750);
nor UO_457 (O_457,N_19924,N_19823);
or UO_458 (O_458,N_19892,N_19938);
nor UO_459 (O_459,N_19917,N_19914);
or UO_460 (O_460,N_19789,N_19956);
nor UO_461 (O_461,N_19816,N_19820);
or UO_462 (O_462,N_19882,N_19840);
or UO_463 (O_463,N_19874,N_19911);
and UO_464 (O_464,N_19785,N_19877);
nand UO_465 (O_465,N_19791,N_19892);
xor UO_466 (O_466,N_19835,N_19753);
nor UO_467 (O_467,N_19879,N_19787);
nand UO_468 (O_468,N_19751,N_19882);
or UO_469 (O_469,N_19892,N_19849);
xnor UO_470 (O_470,N_19876,N_19870);
nor UO_471 (O_471,N_19755,N_19837);
nand UO_472 (O_472,N_19774,N_19790);
nand UO_473 (O_473,N_19940,N_19994);
xor UO_474 (O_474,N_19957,N_19974);
nor UO_475 (O_475,N_19971,N_19968);
xnor UO_476 (O_476,N_19940,N_19901);
nor UO_477 (O_477,N_19937,N_19791);
or UO_478 (O_478,N_19802,N_19789);
nor UO_479 (O_479,N_19770,N_19885);
nor UO_480 (O_480,N_19914,N_19821);
and UO_481 (O_481,N_19836,N_19900);
nor UO_482 (O_482,N_19930,N_19832);
nand UO_483 (O_483,N_19783,N_19804);
nor UO_484 (O_484,N_19983,N_19840);
xor UO_485 (O_485,N_19776,N_19822);
and UO_486 (O_486,N_19925,N_19955);
nor UO_487 (O_487,N_19910,N_19928);
xnor UO_488 (O_488,N_19795,N_19901);
nor UO_489 (O_489,N_19833,N_19879);
nand UO_490 (O_490,N_19855,N_19753);
and UO_491 (O_491,N_19932,N_19756);
xnor UO_492 (O_492,N_19914,N_19930);
nand UO_493 (O_493,N_19961,N_19784);
or UO_494 (O_494,N_19828,N_19990);
or UO_495 (O_495,N_19861,N_19905);
nor UO_496 (O_496,N_19798,N_19867);
xnor UO_497 (O_497,N_19892,N_19810);
xnor UO_498 (O_498,N_19937,N_19977);
nand UO_499 (O_499,N_19855,N_19954);
nand UO_500 (O_500,N_19923,N_19927);
and UO_501 (O_501,N_19970,N_19905);
or UO_502 (O_502,N_19834,N_19771);
or UO_503 (O_503,N_19858,N_19836);
nor UO_504 (O_504,N_19967,N_19914);
nor UO_505 (O_505,N_19909,N_19934);
and UO_506 (O_506,N_19762,N_19765);
nand UO_507 (O_507,N_19986,N_19855);
nand UO_508 (O_508,N_19904,N_19788);
xor UO_509 (O_509,N_19763,N_19959);
xnor UO_510 (O_510,N_19767,N_19958);
or UO_511 (O_511,N_19765,N_19795);
nand UO_512 (O_512,N_19923,N_19872);
and UO_513 (O_513,N_19879,N_19996);
nor UO_514 (O_514,N_19870,N_19910);
xor UO_515 (O_515,N_19789,N_19824);
nand UO_516 (O_516,N_19844,N_19906);
nor UO_517 (O_517,N_19945,N_19999);
nor UO_518 (O_518,N_19766,N_19966);
xnor UO_519 (O_519,N_19932,N_19808);
and UO_520 (O_520,N_19839,N_19977);
nand UO_521 (O_521,N_19846,N_19841);
and UO_522 (O_522,N_19903,N_19765);
nor UO_523 (O_523,N_19945,N_19785);
nand UO_524 (O_524,N_19889,N_19927);
and UO_525 (O_525,N_19992,N_19764);
or UO_526 (O_526,N_19791,N_19993);
nand UO_527 (O_527,N_19818,N_19985);
or UO_528 (O_528,N_19934,N_19993);
xnor UO_529 (O_529,N_19867,N_19963);
xnor UO_530 (O_530,N_19972,N_19930);
nand UO_531 (O_531,N_19948,N_19770);
or UO_532 (O_532,N_19910,N_19983);
xnor UO_533 (O_533,N_19771,N_19898);
nand UO_534 (O_534,N_19826,N_19889);
or UO_535 (O_535,N_19751,N_19886);
or UO_536 (O_536,N_19893,N_19776);
or UO_537 (O_537,N_19797,N_19789);
or UO_538 (O_538,N_19753,N_19939);
nand UO_539 (O_539,N_19852,N_19839);
or UO_540 (O_540,N_19786,N_19782);
and UO_541 (O_541,N_19775,N_19881);
or UO_542 (O_542,N_19938,N_19978);
or UO_543 (O_543,N_19806,N_19935);
or UO_544 (O_544,N_19875,N_19953);
or UO_545 (O_545,N_19843,N_19867);
and UO_546 (O_546,N_19844,N_19911);
or UO_547 (O_547,N_19955,N_19992);
nor UO_548 (O_548,N_19918,N_19787);
or UO_549 (O_549,N_19913,N_19814);
or UO_550 (O_550,N_19865,N_19935);
and UO_551 (O_551,N_19874,N_19823);
nor UO_552 (O_552,N_19896,N_19789);
nand UO_553 (O_553,N_19889,N_19821);
or UO_554 (O_554,N_19771,N_19989);
nor UO_555 (O_555,N_19769,N_19782);
nand UO_556 (O_556,N_19896,N_19968);
nand UO_557 (O_557,N_19762,N_19876);
xnor UO_558 (O_558,N_19983,N_19783);
and UO_559 (O_559,N_19877,N_19970);
nor UO_560 (O_560,N_19885,N_19914);
or UO_561 (O_561,N_19967,N_19908);
nor UO_562 (O_562,N_19967,N_19972);
nand UO_563 (O_563,N_19832,N_19943);
nor UO_564 (O_564,N_19883,N_19764);
xor UO_565 (O_565,N_19752,N_19813);
xor UO_566 (O_566,N_19965,N_19840);
nand UO_567 (O_567,N_19884,N_19818);
nand UO_568 (O_568,N_19902,N_19937);
xor UO_569 (O_569,N_19756,N_19968);
and UO_570 (O_570,N_19857,N_19992);
nor UO_571 (O_571,N_19753,N_19957);
nor UO_572 (O_572,N_19921,N_19909);
or UO_573 (O_573,N_19984,N_19909);
or UO_574 (O_574,N_19978,N_19821);
xor UO_575 (O_575,N_19908,N_19935);
and UO_576 (O_576,N_19753,N_19856);
or UO_577 (O_577,N_19960,N_19786);
nand UO_578 (O_578,N_19858,N_19845);
xnor UO_579 (O_579,N_19810,N_19907);
or UO_580 (O_580,N_19871,N_19987);
nor UO_581 (O_581,N_19764,N_19959);
and UO_582 (O_582,N_19991,N_19986);
and UO_583 (O_583,N_19858,N_19872);
xnor UO_584 (O_584,N_19902,N_19909);
nor UO_585 (O_585,N_19957,N_19898);
nand UO_586 (O_586,N_19804,N_19793);
or UO_587 (O_587,N_19836,N_19983);
xnor UO_588 (O_588,N_19833,N_19997);
or UO_589 (O_589,N_19940,N_19904);
nand UO_590 (O_590,N_19841,N_19779);
and UO_591 (O_591,N_19990,N_19924);
xnor UO_592 (O_592,N_19840,N_19915);
nand UO_593 (O_593,N_19834,N_19972);
or UO_594 (O_594,N_19789,N_19990);
or UO_595 (O_595,N_19809,N_19830);
and UO_596 (O_596,N_19900,N_19957);
xor UO_597 (O_597,N_19926,N_19868);
and UO_598 (O_598,N_19777,N_19835);
xor UO_599 (O_599,N_19833,N_19842);
or UO_600 (O_600,N_19844,N_19836);
and UO_601 (O_601,N_19929,N_19853);
and UO_602 (O_602,N_19826,N_19916);
xnor UO_603 (O_603,N_19888,N_19994);
and UO_604 (O_604,N_19837,N_19836);
xor UO_605 (O_605,N_19956,N_19964);
or UO_606 (O_606,N_19797,N_19968);
nand UO_607 (O_607,N_19827,N_19974);
or UO_608 (O_608,N_19988,N_19996);
and UO_609 (O_609,N_19903,N_19895);
nor UO_610 (O_610,N_19970,N_19863);
and UO_611 (O_611,N_19841,N_19952);
or UO_612 (O_612,N_19848,N_19828);
nand UO_613 (O_613,N_19813,N_19834);
nand UO_614 (O_614,N_19865,N_19965);
nor UO_615 (O_615,N_19844,N_19960);
or UO_616 (O_616,N_19923,N_19981);
or UO_617 (O_617,N_19929,N_19937);
nor UO_618 (O_618,N_19922,N_19883);
nor UO_619 (O_619,N_19929,N_19920);
xor UO_620 (O_620,N_19868,N_19947);
nand UO_621 (O_621,N_19863,N_19815);
nor UO_622 (O_622,N_19976,N_19755);
and UO_623 (O_623,N_19827,N_19981);
nor UO_624 (O_624,N_19781,N_19878);
xnor UO_625 (O_625,N_19767,N_19760);
or UO_626 (O_626,N_19911,N_19799);
xor UO_627 (O_627,N_19817,N_19833);
xnor UO_628 (O_628,N_19778,N_19882);
and UO_629 (O_629,N_19829,N_19991);
and UO_630 (O_630,N_19913,N_19964);
and UO_631 (O_631,N_19805,N_19806);
and UO_632 (O_632,N_19867,N_19830);
and UO_633 (O_633,N_19954,N_19774);
nand UO_634 (O_634,N_19895,N_19995);
or UO_635 (O_635,N_19798,N_19879);
or UO_636 (O_636,N_19803,N_19794);
xnor UO_637 (O_637,N_19913,N_19886);
xnor UO_638 (O_638,N_19921,N_19815);
nand UO_639 (O_639,N_19907,N_19841);
and UO_640 (O_640,N_19781,N_19912);
and UO_641 (O_641,N_19826,N_19998);
nand UO_642 (O_642,N_19769,N_19776);
nor UO_643 (O_643,N_19984,N_19824);
nand UO_644 (O_644,N_19759,N_19812);
xnor UO_645 (O_645,N_19982,N_19970);
xor UO_646 (O_646,N_19776,N_19910);
xnor UO_647 (O_647,N_19865,N_19806);
nor UO_648 (O_648,N_19751,N_19832);
and UO_649 (O_649,N_19892,N_19927);
xnor UO_650 (O_650,N_19906,N_19977);
nor UO_651 (O_651,N_19816,N_19962);
or UO_652 (O_652,N_19904,N_19858);
nor UO_653 (O_653,N_19830,N_19936);
or UO_654 (O_654,N_19883,N_19898);
nand UO_655 (O_655,N_19846,N_19766);
and UO_656 (O_656,N_19780,N_19946);
nand UO_657 (O_657,N_19995,N_19850);
nor UO_658 (O_658,N_19890,N_19862);
xnor UO_659 (O_659,N_19904,N_19962);
nor UO_660 (O_660,N_19867,N_19988);
or UO_661 (O_661,N_19814,N_19980);
nor UO_662 (O_662,N_19851,N_19986);
and UO_663 (O_663,N_19913,N_19873);
nor UO_664 (O_664,N_19894,N_19942);
xor UO_665 (O_665,N_19832,N_19934);
and UO_666 (O_666,N_19897,N_19786);
or UO_667 (O_667,N_19957,N_19975);
or UO_668 (O_668,N_19903,N_19947);
xnor UO_669 (O_669,N_19808,N_19777);
and UO_670 (O_670,N_19886,N_19947);
and UO_671 (O_671,N_19926,N_19946);
or UO_672 (O_672,N_19848,N_19978);
nor UO_673 (O_673,N_19812,N_19887);
or UO_674 (O_674,N_19837,N_19890);
nand UO_675 (O_675,N_19861,N_19777);
and UO_676 (O_676,N_19885,N_19841);
xnor UO_677 (O_677,N_19905,N_19959);
and UO_678 (O_678,N_19950,N_19894);
nor UO_679 (O_679,N_19966,N_19939);
nand UO_680 (O_680,N_19941,N_19995);
nor UO_681 (O_681,N_19817,N_19863);
nor UO_682 (O_682,N_19780,N_19888);
nor UO_683 (O_683,N_19778,N_19793);
xor UO_684 (O_684,N_19816,N_19853);
xnor UO_685 (O_685,N_19750,N_19854);
and UO_686 (O_686,N_19888,N_19783);
xnor UO_687 (O_687,N_19894,N_19866);
and UO_688 (O_688,N_19858,N_19963);
and UO_689 (O_689,N_19779,N_19999);
nand UO_690 (O_690,N_19808,N_19856);
nor UO_691 (O_691,N_19762,N_19818);
xnor UO_692 (O_692,N_19814,N_19760);
xor UO_693 (O_693,N_19833,N_19791);
or UO_694 (O_694,N_19778,N_19928);
and UO_695 (O_695,N_19866,N_19976);
or UO_696 (O_696,N_19861,N_19994);
xnor UO_697 (O_697,N_19777,N_19949);
xor UO_698 (O_698,N_19987,N_19980);
nor UO_699 (O_699,N_19997,N_19813);
xor UO_700 (O_700,N_19854,N_19862);
nor UO_701 (O_701,N_19817,N_19964);
nor UO_702 (O_702,N_19845,N_19983);
nand UO_703 (O_703,N_19867,N_19855);
and UO_704 (O_704,N_19808,N_19890);
nand UO_705 (O_705,N_19953,N_19942);
nand UO_706 (O_706,N_19903,N_19770);
nand UO_707 (O_707,N_19834,N_19790);
and UO_708 (O_708,N_19989,N_19868);
nand UO_709 (O_709,N_19926,N_19783);
xor UO_710 (O_710,N_19964,N_19983);
xnor UO_711 (O_711,N_19936,N_19871);
nor UO_712 (O_712,N_19949,N_19784);
nand UO_713 (O_713,N_19836,N_19767);
nand UO_714 (O_714,N_19987,N_19913);
xor UO_715 (O_715,N_19903,N_19762);
or UO_716 (O_716,N_19801,N_19750);
nand UO_717 (O_717,N_19871,N_19755);
nand UO_718 (O_718,N_19762,N_19944);
xor UO_719 (O_719,N_19895,N_19825);
nor UO_720 (O_720,N_19864,N_19923);
nor UO_721 (O_721,N_19997,N_19958);
nor UO_722 (O_722,N_19915,N_19982);
nor UO_723 (O_723,N_19994,N_19821);
nand UO_724 (O_724,N_19991,N_19901);
nor UO_725 (O_725,N_19890,N_19941);
and UO_726 (O_726,N_19992,N_19883);
and UO_727 (O_727,N_19865,N_19964);
nand UO_728 (O_728,N_19815,N_19782);
or UO_729 (O_729,N_19969,N_19863);
nand UO_730 (O_730,N_19982,N_19853);
and UO_731 (O_731,N_19799,N_19822);
or UO_732 (O_732,N_19835,N_19820);
or UO_733 (O_733,N_19809,N_19829);
nor UO_734 (O_734,N_19819,N_19828);
xnor UO_735 (O_735,N_19885,N_19916);
and UO_736 (O_736,N_19846,N_19825);
nor UO_737 (O_737,N_19931,N_19940);
nand UO_738 (O_738,N_19896,N_19769);
and UO_739 (O_739,N_19915,N_19753);
nand UO_740 (O_740,N_19937,N_19882);
or UO_741 (O_741,N_19954,N_19980);
nor UO_742 (O_742,N_19819,N_19912);
nand UO_743 (O_743,N_19765,N_19794);
nand UO_744 (O_744,N_19941,N_19778);
or UO_745 (O_745,N_19753,N_19774);
or UO_746 (O_746,N_19874,N_19820);
nor UO_747 (O_747,N_19903,N_19829);
or UO_748 (O_748,N_19896,N_19826);
nor UO_749 (O_749,N_19880,N_19796);
and UO_750 (O_750,N_19919,N_19899);
nand UO_751 (O_751,N_19988,N_19750);
nor UO_752 (O_752,N_19859,N_19872);
xnor UO_753 (O_753,N_19784,N_19911);
nand UO_754 (O_754,N_19874,N_19834);
nor UO_755 (O_755,N_19940,N_19801);
xnor UO_756 (O_756,N_19822,N_19838);
and UO_757 (O_757,N_19824,N_19840);
or UO_758 (O_758,N_19851,N_19970);
or UO_759 (O_759,N_19913,N_19929);
nand UO_760 (O_760,N_19902,N_19886);
and UO_761 (O_761,N_19767,N_19896);
nand UO_762 (O_762,N_19844,N_19754);
xnor UO_763 (O_763,N_19962,N_19827);
xor UO_764 (O_764,N_19916,N_19983);
or UO_765 (O_765,N_19955,N_19989);
nor UO_766 (O_766,N_19859,N_19908);
xor UO_767 (O_767,N_19863,N_19864);
xnor UO_768 (O_768,N_19905,N_19859);
xor UO_769 (O_769,N_19924,N_19978);
nand UO_770 (O_770,N_19845,N_19948);
or UO_771 (O_771,N_19874,N_19913);
nor UO_772 (O_772,N_19762,N_19945);
xnor UO_773 (O_773,N_19970,N_19975);
nand UO_774 (O_774,N_19835,N_19750);
nor UO_775 (O_775,N_19836,N_19855);
or UO_776 (O_776,N_19793,N_19765);
and UO_777 (O_777,N_19787,N_19899);
or UO_778 (O_778,N_19942,N_19949);
xor UO_779 (O_779,N_19813,N_19880);
xnor UO_780 (O_780,N_19885,N_19913);
and UO_781 (O_781,N_19956,N_19885);
nor UO_782 (O_782,N_19915,N_19807);
nor UO_783 (O_783,N_19950,N_19885);
and UO_784 (O_784,N_19853,N_19771);
or UO_785 (O_785,N_19991,N_19853);
nand UO_786 (O_786,N_19872,N_19988);
nand UO_787 (O_787,N_19975,N_19983);
and UO_788 (O_788,N_19979,N_19981);
xor UO_789 (O_789,N_19937,N_19862);
nor UO_790 (O_790,N_19891,N_19778);
xnor UO_791 (O_791,N_19900,N_19760);
and UO_792 (O_792,N_19999,N_19830);
and UO_793 (O_793,N_19800,N_19889);
and UO_794 (O_794,N_19933,N_19970);
xnor UO_795 (O_795,N_19858,N_19823);
xor UO_796 (O_796,N_19959,N_19867);
nand UO_797 (O_797,N_19980,N_19867);
and UO_798 (O_798,N_19932,N_19845);
nor UO_799 (O_799,N_19974,N_19753);
and UO_800 (O_800,N_19914,N_19817);
and UO_801 (O_801,N_19958,N_19758);
xnor UO_802 (O_802,N_19898,N_19901);
or UO_803 (O_803,N_19820,N_19854);
or UO_804 (O_804,N_19926,N_19777);
xnor UO_805 (O_805,N_19923,N_19883);
nand UO_806 (O_806,N_19992,N_19956);
nand UO_807 (O_807,N_19982,N_19987);
or UO_808 (O_808,N_19865,N_19986);
nor UO_809 (O_809,N_19791,N_19965);
nand UO_810 (O_810,N_19863,N_19814);
nand UO_811 (O_811,N_19768,N_19944);
nand UO_812 (O_812,N_19960,N_19780);
and UO_813 (O_813,N_19843,N_19927);
or UO_814 (O_814,N_19886,N_19950);
or UO_815 (O_815,N_19856,N_19821);
and UO_816 (O_816,N_19833,N_19975);
or UO_817 (O_817,N_19836,N_19797);
nor UO_818 (O_818,N_19753,N_19983);
nand UO_819 (O_819,N_19951,N_19856);
and UO_820 (O_820,N_19824,N_19961);
nor UO_821 (O_821,N_19777,N_19889);
and UO_822 (O_822,N_19998,N_19969);
nand UO_823 (O_823,N_19812,N_19983);
and UO_824 (O_824,N_19958,N_19889);
and UO_825 (O_825,N_19835,N_19858);
nand UO_826 (O_826,N_19764,N_19762);
or UO_827 (O_827,N_19951,N_19987);
and UO_828 (O_828,N_19921,N_19982);
and UO_829 (O_829,N_19830,N_19919);
xor UO_830 (O_830,N_19993,N_19755);
nand UO_831 (O_831,N_19780,N_19794);
nor UO_832 (O_832,N_19892,N_19859);
or UO_833 (O_833,N_19967,N_19916);
xor UO_834 (O_834,N_19791,N_19904);
or UO_835 (O_835,N_19768,N_19979);
or UO_836 (O_836,N_19822,N_19971);
or UO_837 (O_837,N_19808,N_19913);
xor UO_838 (O_838,N_19955,N_19808);
xor UO_839 (O_839,N_19796,N_19809);
xnor UO_840 (O_840,N_19974,N_19990);
and UO_841 (O_841,N_19841,N_19832);
and UO_842 (O_842,N_19822,N_19951);
nor UO_843 (O_843,N_19831,N_19808);
xnor UO_844 (O_844,N_19993,N_19780);
and UO_845 (O_845,N_19837,N_19838);
or UO_846 (O_846,N_19788,N_19909);
nor UO_847 (O_847,N_19883,N_19944);
nor UO_848 (O_848,N_19932,N_19903);
xor UO_849 (O_849,N_19818,N_19951);
xor UO_850 (O_850,N_19903,N_19959);
nor UO_851 (O_851,N_19790,N_19839);
nand UO_852 (O_852,N_19767,N_19909);
or UO_853 (O_853,N_19955,N_19778);
xnor UO_854 (O_854,N_19805,N_19774);
xor UO_855 (O_855,N_19902,N_19790);
nand UO_856 (O_856,N_19937,N_19863);
nor UO_857 (O_857,N_19896,N_19962);
xor UO_858 (O_858,N_19767,N_19916);
or UO_859 (O_859,N_19867,N_19840);
nor UO_860 (O_860,N_19922,N_19925);
nand UO_861 (O_861,N_19828,N_19792);
xor UO_862 (O_862,N_19802,N_19947);
or UO_863 (O_863,N_19840,N_19946);
and UO_864 (O_864,N_19866,N_19759);
and UO_865 (O_865,N_19868,N_19780);
or UO_866 (O_866,N_19982,N_19929);
and UO_867 (O_867,N_19827,N_19894);
nand UO_868 (O_868,N_19958,N_19874);
nand UO_869 (O_869,N_19945,N_19947);
nand UO_870 (O_870,N_19762,N_19902);
xor UO_871 (O_871,N_19849,N_19821);
and UO_872 (O_872,N_19855,N_19823);
nand UO_873 (O_873,N_19852,N_19979);
nand UO_874 (O_874,N_19906,N_19848);
nand UO_875 (O_875,N_19910,N_19841);
or UO_876 (O_876,N_19887,N_19925);
xor UO_877 (O_877,N_19845,N_19809);
or UO_878 (O_878,N_19776,N_19926);
or UO_879 (O_879,N_19897,N_19796);
xnor UO_880 (O_880,N_19800,N_19831);
and UO_881 (O_881,N_19877,N_19856);
or UO_882 (O_882,N_19802,N_19865);
xnor UO_883 (O_883,N_19773,N_19888);
or UO_884 (O_884,N_19849,N_19891);
and UO_885 (O_885,N_19938,N_19774);
and UO_886 (O_886,N_19850,N_19945);
nor UO_887 (O_887,N_19854,N_19758);
and UO_888 (O_888,N_19944,N_19923);
or UO_889 (O_889,N_19873,N_19970);
nor UO_890 (O_890,N_19869,N_19903);
nand UO_891 (O_891,N_19843,N_19924);
or UO_892 (O_892,N_19872,N_19922);
and UO_893 (O_893,N_19899,N_19970);
nand UO_894 (O_894,N_19940,N_19937);
nor UO_895 (O_895,N_19986,N_19854);
or UO_896 (O_896,N_19956,N_19751);
xor UO_897 (O_897,N_19760,N_19994);
and UO_898 (O_898,N_19905,N_19918);
and UO_899 (O_899,N_19841,N_19992);
xnor UO_900 (O_900,N_19884,N_19984);
xnor UO_901 (O_901,N_19860,N_19789);
nand UO_902 (O_902,N_19845,N_19810);
and UO_903 (O_903,N_19966,N_19968);
xor UO_904 (O_904,N_19815,N_19853);
and UO_905 (O_905,N_19818,N_19832);
nand UO_906 (O_906,N_19792,N_19767);
nor UO_907 (O_907,N_19827,N_19784);
nor UO_908 (O_908,N_19933,N_19793);
nand UO_909 (O_909,N_19875,N_19802);
xnor UO_910 (O_910,N_19960,N_19917);
or UO_911 (O_911,N_19954,N_19771);
or UO_912 (O_912,N_19819,N_19954);
nor UO_913 (O_913,N_19975,N_19839);
xnor UO_914 (O_914,N_19890,N_19901);
nor UO_915 (O_915,N_19888,N_19804);
or UO_916 (O_916,N_19762,N_19772);
nand UO_917 (O_917,N_19793,N_19972);
or UO_918 (O_918,N_19910,N_19916);
or UO_919 (O_919,N_19798,N_19991);
and UO_920 (O_920,N_19875,N_19906);
or UO_921 (O_921,N_19794,N_19902);
nand UO_922 (O_922,N_19752,N_19933);
xnor UO_923 (O_923,N_19937,N_19778);
or UO_924 (O_924,N_19863,N_19801);
nand UO_925 (O_925,N_19840,N_19802);
xnor UO_926 (O_926,N_19897,N_19902);
xor UO_927 (O_927,N_19812,N_19977);
nor UO_928 (O_928,N_19878,N_19792);
xnor UO_929 (O_929,N_19753,N_19809);
nor UO_930 (O_930,N_19918,N_19956);
or UO_931 (O_931,N_19788,N_19997);
nand UO_932 (O_932,N_19937,N_19755);
and UO_933 (O_933,N_19912,N_19851);
or UO_934 (O_934,N_19915,N_19975);
or UO_935 (O_935,N_19808,N_19989);
and UO_936 (O_936,N_19870,N_19847);
or UO_937 (O_937,N_19975,N_19836);
xor UO_938 (O_938,N_19758,N_19750);
nand UO_939 (O_939,N_19828,N_19946);
xor UO_940 (O_940,N_19946,N_19762);
and UO_941 (O_941,N_19982,N_19941);
nand UO_942 (O_942,N_19770,N_19935);
nor UO_943 (O_943,N_19771,N_19951);
nor UO_944 (O_944,N_19760,N_19797);
xnor UO_945 (O_945,N_19858,N_19775);
nand UO_946 (O_946,N_19838,N_19928);
or UO_947 (O_947,N_19873,N_19910);
and UO_948 (O_948,N_19898,N_19864);
or UO_949 (O_949,N_19893,N_19805);
xnor UO_950 (O_950,N_19907,N_19868);
nand UO_951 (O_951,N_19920,N_19959);
and UO_952 (O_952,N_19785,N_19925);
nor UO_953 (O_953,N_19754,N_19880);
xor UO_954 (O_954,N_19975,N_19929);
and UO_955 (O_955,N_19801,N_19787);
and UO_956 (O_956,N_19756,N_19926);
nor UO_957 (O_957,N_19985,N_19865);
xor UO_958 (O_958,N_19829,N_19973);
xnor UO_959 (O_959,N_19885,N_19761);
or UO_960 (O_960,N_19869,N_19988);
nand UO_961 (O_961,N_19827,N_19946);
xor UO_962 (O_962,N_19812,N_19926);
nand UO_963 (O_963,N_19996,N_19833);
nand UO_964 (O_964,N_19809,N_19952);
and UO_965 (O_965,N_19773,N_19829);
nand UO_966 (O_966,N_19776,N_19800);
xnor UO_967 (O_967,N_19760,N_19969);
nor UO_968 (O_968,N_19866,N_19816);
nor UO_969 (O_969,N_19911,N_19967);
and UO_970 (O_970,N_19788,N_19816);
nand UO_971 (O_971,N_19909,N_19939);
xor UO_972 (O_972,N_19872,N_19831);
xnor UO_973 (O_973,N_19762,N_19782);
nand UO_974 (O_974,N_19823,N_19991);
nor UO_975 (O_975,N_19925,N_19811);
and UO_976 (O_976,N_19864,N_19990);
xor UO_977 (O_977,N_19832,N_19944);
nand UO_978 (O_978,N_19892,N_19983);
nand UO_979 (O_979,N_19863,N_19966);
xor UO_980 (O_980,N_19758,N_19914);
nor UO_981 (O_981,N_19976,N_19987);
and UO_982 (O_982,N_19857,N_19967);
nand UO_983 (O_983,N_19920,N_19994);
nor UO_984 (O_984,N_19815,N_19856);
nor UO_985 (O_985,N_19932,N_19782);
xor UO_986 (O_986,N_19761,N_19927);
xnor UO_987 (O_987,N_19901,N_19887);
xor UO_988 (O_988,N_19942,N_19994);
xor UO_989 (O_989,N_19915,N_19939);
nand UO_990 (O_990,N_19990,N_19912);
xor UO_991 (O_991,N_19885,N_19998);
xor UO_992 (O_992,N_19757,N_19969);
and UO_993 (O_993,N_19911,N_19830);
xnor UO_994 (O_994,N_19929,N_19905);
nand UO_995 (O_995,N_19759,N_19777);
xor UO_996 (O_996,N_19951,N_19966);
nand UO_997 (O_997,N_19873,N_19859);
or UO_998 (O_998,N_19778,N_19770);
or UO_999 (O_999,N_19814,N_19971);
nand UO_1000 (O_1000,N_19828,N_19935);
and UO_1001 (O_1001,N_19801,N_19830);
xor UO_1002 (O_1002,N_19908,N_19925);
or UO_1003 (O_1003,N_19816,N_19967);
and UO_1004 (O_1004,N_19764,N_19948);
nand UO_1005 (O_1005,N_19844,N_19942);
nand UO_1006 (O_1006,N_19916,N_19785);
nand UO_1007 (O_1007,N_19788,N_19925);
xor UO_1008 (O_1008,N_19889,N_19964);
nor UO_1009 (O_1009,N_19885,N_19907);
or UO_1010 (O_1010,N_19854,N_19819);
xor UO_1011 (O_1011,N_19856,N_19811);
xor UO_1012 (O_1012,N_19932,N_19821);
nand UO_1013 (O_1013,N_19814,N_19910);
xor UO_1014 (O_1014,N_19757,N_19937);
or UO_1015 (O_1015,N_19847,N_19937);
xnor UO_1016 (O_1016,N_19844,N_19759);
nor UO_1017 (O_1017,N_19751,N_19952);
nor UO_1018 (O_1018,N_19898,N_19842);
or UO_1019 (O_1019,N_19835,N_19889);
and UO_1020 (O_1020,N_19936,N_19756);
xnor UO_1021 (O_1021,N_19970,N_19767);
xnor UO_1022 (O_1022,N_19809,N_19962);
or UO_1023 (O_1023,N_19989,N_19954);
or UO_1024 (O_1024,N_19840,N_19798);
nor UO_1025 (O_1025,N_19969,N_19991);
and UO_1026 (O_1026,N_19990,N_19790);
xor UO_1027 (O_1027,N_19916,N_19815);
xnor UO_1028 (O_1028,N_19821,N_19891);
nand UO_1029 (O_1029,N_19927,N_19754);
xor UO_1030 (O_1030,N_19759,N_19984);
xnor UO_1031 (O_1031,N_19794,N_19997);
nor UO_1032 (O_1032,N_19951,N_19971);
or UO_1033 (O_1033,N_19936,N_19999);
or UO_1034 (O_1034,N_19881,N_19800);
nand UO_1035 (O_1035,N_19772,N_19777);
xnor UO_1036 (O_1036,N_19873,N_19946);
nand UO_1037 (O_1037,N_19773,N_19952);
nor UO_1038 (O_1038,N_19871,N_19751);
nand UO_1039 (O_1039,N_19839,N_19968);
nand UO_1040 (O_1040,N_19879,N_19861);
nor UO_1041 (O_1041,N_19957,N_19824);
xnor UO_1042 (O_1042,N_19839,N_19932);
nand UO_1043 (O_1043,N_19963,N_19893);
and UO_1044 (O_1044,N_19781,N_19841);
nor UO_1045 (O_1045,N_19911,N_19847);
and UO_1046 (O_1046,N_19824,N_19766);
and UO_1047 (O_1047,N_19811,N_19924);
or UO_1048 (O_1048,N_19764,N_19929);
or UO_1049 (O_1049,N_19884,N_19772);
nand UO_1050 (O_1050,N_19941,N_19836);
or UO_1051 (O_1051,N_19854,N_19851);
nor UO_1052 (O_1052,N_19786,N_19888);
xnor UO_1053 (O_1053,N_19776,N_19752);
xnor UO_1054 (O_1054,N_19982,N_19953);
nor UO_1055 (O_1055,N_19786,N_19826);
nor UO_1056 (O_1056,N_19804,N_19848);
nand UO_1057 (O_1057,N_19835,N_19904);
xnor UO_1058 (O_1058,N_19875,N_19819);
nand UO_1059 (O_1059,N_19854,N_19818);
nor UO_1060 (O_1060,N_19906,N_19770);
xnor UO_1061 (O_1061,N_19916,N_19760);
nor UO_1062 (O_1062,N_19950,N_19784);
nand UO_1063 (O_1063,N_19764,N_19913);
and UO_1064 (O_1064,N_19922,N_19893);
nand UO_1065 (O_1065,N_19857,N_19854);
nand UO_1066 (O_1066,N_19874,N_19894);
xnor UO_1067 (O_1067,N_19776,N_19922);
xor UO_1068 (O_1068,N_19826,N_19897);
or UO_1069 (O_1069,N_19888,N_19840);
nand UO_1070 (O_1070,N_19942,N_19989);
or UO_1071 (O_1071,N_19872,N_19935);
and UO_1072 (O_1072,N_19965,N_19892);
or UO_1073 (O_1073,N_19849,N_19893);
nor UO_1074 (O_1074,N_19970,N_19768);
or UO_1075 (O_1075,N_19752,N_19951);
and UO_1076 (O_1076,N_19787,N_19890);
xor UO_1077 (O_1077,N_19961,N_19982);
nor UO_1078 (O_1078,N_19992,N_19854);
and UO_1079 (O_1079,N_19789,N_19807);
nand UO_1080 (O_1080,N_19867,N_19910);
and UO_1081 (O_1081,N_19844,N_19876);
or UO_1082 (O_1082,N_19838,N_19933);
nor UO_1083 (O_1083,N_19965,N_19799);
nand UO_1084 (O_1084,N_19783,N_19920);
and UO_1085 (O_1085,N_19910,N_19771);
nor UO_1086 (O_1086,N_19835,N_19842);
xor UO_1087 (O_1087,N_19986,N_19861);
nor UO_1088 (O_1088,N_19837,N_19798);
or UO_1089 (O_1089,N_19969,N_19768);
or UO_1090 (O_1090,N_19977,N_19859);
nand UO_1091 (O_1091,N_19811,N_19999);
nor UO_1092 (O_1092,N_19771,N_19851);
and UO_1093 (O_1093,N_19757,N_19943);
and UO_1094 (O_1094,N_19926,N_19781);
nand UO_1095 (O_1095,N_19890,N_19816);
and UO_1096 (O_1096,N_19883,N_19761);
xor UO_1097 (O_1097,N_19758,N_19794);
nand UO_1098 (O_1098,N_19857,N_19820);
nor UO_1099 (O_1099,N_19989,N_19937);
and UO_1100 (O_1100,N_19923,N_19979);
nor UO_1101 (O_1101,N_19764,N_19862);
xor UO_1102 (O_1102,N_19814,N_19998);
nand UO_1103 (O_1103,N_19989,N_19816);
nor UO_1104 (O_1104,N_19887,N_19865);
and UO_1105 (O_1105,N_19879,N_19750);
xor UO_1106 (O_1106,N_19937,N_19946);
nor UO_1107 (O_1107,N_19777,N_19998);
nor UO_1108 (O_1108,N_19929,N_19987);
nand UO_1109 (O_1109,N_19841,N_19851);
xor UO_1110 (O_1110,N_19924,N_19996);
and UO_1111 (O_1111,N_19762,N_19936);
and UO_1112 (O_1112,N_19787,N_19903);
and UO_1113 (O_1113,N_19956,N_19909);
nor UO_1114 (O_1114,N_19810,N_19897);
or UO_1115 (O_1115,N_19991,N_19879);
nor UO_1116 (O_1116,N_19895,N_19916);
nand UO_1117 (O_1117,N_19849,N_19865);
nand UO_1118 (O_1118,N_19833,N_19852);
nor UO_1119 (O_1119,N_19954,N_19806);
nor UO_1120 (O_1120,N_19834,N_19947);
nand UO_1121 (O_1121,N_19792,N_19834);
nor UO_1122 (O_1122,N_19997,N_19934);
nor UO_1123 (O_1123,N_19820,N_19908);
nor UO_1124 (O_1124,N_19766,N_19965);
xnor UO_1125 (O_1125,N_19968,N_19934);
and UO_1126 (O_1126,N_19969,N_19756);
or UO_1127 (O_1127,N_19754,N_19975);
or UO_1128 (O_1128,N_19883,N_19777);
and UO_1129 (O_1129,N_19923,N_19849);
nand UO_1130 (O_1130,N_19935,N_19996);
nand UO_1131 (O_1131,N_19990,N_19885);
or UO_1132 (O_1132,N_19821,N_19899);
xor UO_1133 (O_1133,N_19928,N_19892);
xnor UO_1134 (O_1134,N_19865,N_19952);
xnor UO_1135 (O_1135,N_19929,N_19991);
xnor UO_1136 (O_1136,N_19981,N_19973);
and UO_1137 (O_1137,N_19889,N_19870);
xor UO_1138 (O_1138,N_19956,N_19899);
or UO_1139 (O_1139,N_19799,N_19853);
or UO_1140 (O_1140,N_19947,N_19793);
or UO_1141 (O_1141,N_19890,N_19792);
nand UO_1142 (O_1142,N_19757,N_19909);
and UO_1143 (O_1143,N_19773,N_19827);
xor UO_1144 (O_1144,N_19809,N_19948);
nand UO_1145 (O_1145,N_19991,N_19850);
or UO_1146 (O_1146,N_19987,N_19989);
or UO_1147 (O_1147,N_19796,N_19969);
xor UO_1148 (O_1148,N_19844,N_19778);
nor UO_1149 (O_1149,N_19902,N_19844);
nor UO_1150 (O_1150,N_19798,N_19841);
or UO_1151 (O_1151,N_19893,N_19866);
and UO_1152 (O_1152,N_19870,N_19826);
or UO_1153 (O_1153,N_19870,N_19757);
and UO_1154 (O_1154,N_19990,N_19819);
or UO_1155 (O_1155,N_19896,N_19832);
and UO_1156 (O_1156,N_19804,N_19905);
nor UO_1157 (O_1157,N_19996,N_19812);
nand UO_1158 (O_1158,N_19807,N_19908);
nor UO_1159 (O_1159,N_19929,N_19957);
nor UO_1160 (O_1160,N_19976,N_19781);
and UO_1161 (O_1161,N_19984,N_19866);
and UO_1162 (O_1162,N_19971,N_19799);
nand UO_1163 (O_1163,N_19877,N_19879);
or UO_1164 (O_1164,N_19847,N_19766);
xor UO_1165 (O_1165,N_19851,N_19897);
nor UO_1166 (O_1166,N_19894,N_19756);
xor UO_1167 (O_1167,N_19883,N_19950);
nor UO_1168 (O_1168,N_19944,N_19998);
xnor UO_1169 (O_1169,N_19968,N_19786);
and UO_1170 (O_1170,N_19769,N_19965);
nand UO_1171 (O_1171,N_19759,N_19768);
xnor UO_1172 (O_1172,N_19849,N_19903);
or UO_1173 (O_1173,N_19837,N_19788);
or UO_1174 (O_1174,N_19764,N_19763);
xor UO_1175 (O_1175,N_19802,N_19835);
nand UO_1176 (O_1176,N_19994,N_19900);
and UO_1177 (O_1177,N_19918,N_19773);
nand UO_1178 (O_1178,N_19880,N_19814);
or UO_1179 (O_1179,N_19869,N_19767);
and UO_1180 (O_1180,N_19842,N_19952);
and UO_1181 (O_1181,N_19982,N_19835);
xor UO_1182 (O_1182,N_19770,N_19813);
and UO_1183 (O_1183,N_19945,N_19765);
xor UO_1184 (O_1184,N_19759,N_19915);
nand UO_1185 (O_1185,N_19907,N_19857);
nor UO_1186 (O_1186,N_19768,N_19786);
or UO_1187 (O_1187,N_19950,N_19995);
or UO_1188 (O_1188,N_19786,N_19753);
xor UO_1189 (O_1189,N_19767,N_19800);
or UO_1190 (O_1190,N_19918,N_19961);
xnor UO_1191 (O_1191,N_19956,N_19894);
xnor UO_1192 (O_1192,N_19907,N_19786);
and UO_1193 (O_1193,N_19968,N_19904);
nor UO_1194 (O_1194,N_19766,N_19931);
xnor UO_1195 (O_1195,N_19841,N_19942);
or UO_1196 (O_1196,N_19830,N_19957);
or UO_1197 (O_1197,N_19886,N_19906);
xnor UO_1198 (O_1198,N_19933,N_19887);
nand UO_1199 (O_1199,N_19816,N_19963);
or UO_1200 (O_1200,N_19877,N_19964);
or UO_1201 (O_1201,N_19781,N_19995);
and UO_1202 (O_1202,N_19893,N_19973);
nand UO_1203 (O_1203,N_19863,N_19796);
xor UO_1204 (O_1204,N_19784,N_19882);
or UO_1205 (O_1205,N_19799,N_19796);
xnor UO_1206 (O_1206,N_19951,N_19781);
or UO_1207 (O_1207,N_19815,N_19970);
nand UO_1208 (O_1208,N_19973,N_19807);
xnor UO_1209 (O_1209,N_19914,N_19776);
and UO_1210 (O_1210,N_19888,N_19928);
or UO_1211 (O_1211,N_19799,N_19919);
nand UO_1212 (O_1212,N_19871,N_19791);
nand UO_1213 (O_1213,N_19899,N_19988);
nand UO_1214 (O_1214,N_19892,N_19901);
and UO_1215 (O_1215,N_19846,N_19984);
xnor UO_1216 (O_1216,N_19757,N_19935);
nand UO_1217 (O_1217,N_19971,N_19789);
xor UO_1218 (O_1218,N_19847,N_19751);
xor UO_1219 (O_1219,N_19964,N_19814);
xor UO_1220 (O_1220,N_19968,N_19891);
xor UO_1221 (O_1221,N_19786,N_19853);
and UO_1222 (O_1222,N_19796,N_19776);
and UO_1223 (O_1223,N_19919,N_19775);
nor UO_1224 (O_1224,N_19810,N_19778);
xnor UO_1225 (O_1225,N_19902,N_19922);
and UO_1226 (O_1226,N_19848,N_19783);
or UO_1227 (O_1227,N_19760,N_19763);
nor UO_1228 (O_1228,N_19795,N_19756);
nor UO_1229 (O_1229,N_19866,N_19981);
or UO_1230 (O_1230,N_19806,N_19899);
or UO_1231 (O_1231,N_19986,N_19985);
nor UO_1232 (O_1232,N_19768,N_19862);
nor UO_1233 (O_1233,N_19841,N_19815);
nor UO_1234 (O_1234,N_19934,N_19773);
nand UO_1235 (O_1235,N_19974,N_19857);
and UO_1236 (O_1236,N_19998,N_19929);
nor UO_1237 (O_1237,N_19887,N_19805);
or UO_1238 (O_1238,N_19952,N_19825);
nor UO_1239 (O_1239,N_19909,N_19938);
nor UO_1240 (O_1240,N_19981,N_19797);
nor UO_1241 (O_1241,N_19983,N_19978);
nand UO_1242 (O_1242,N_19858,N_19788);
xnor UO_1243 (O_1243,N_19816,N_19899);
nand UO_1244 (O_1244,N_19954,N_19918);
and UO_1245 (O_1245,N_19771,N_19766);
xor UO_1246 (O_1246,N_19904,N_19995);
nand UO_1247 (O_1247,N_19956,N_19853);
xnor UO_1248 (O_1248,N_19998,N_19852);
nand UO_1249 (O_1249,N_19990,N_19918);
nand UO_1250 (O_1250,N_19767,N_19758);
or UO_1251 (O_1251,N_19936,N_19809);
xnor UO_1252 (O_1252,N_19915,N_19875);
nor UO_1253 (O_1253,N_19853,N_19819);
and UO_1254 (O_1254,N_19985,N_19836);
nand UO_1255 (O_1255,N_19961,N_19907);
nor UO_1256 (O_1256,N_19986,N_19794);
and UO_1257 (O_1257,N_19986,N_19899);
xor UO_1258 (O_1258,N_19972,N_19837);
nand UO_1259 (O_1259,N_19922,N_19924);
nand UO_1260 (O_1260,N_19783,N_19895);
nand UO_1261 (O_1261,N_19901,N_19806);
nand UO_1262 (O_1262,N_19923,N_19956);
nand UO_1263 (O_1263,N_19764,N_19949);
nand UO_1264 (O_1264,N_19924,N_19845);
and UO_1265 (O_1265,N_19909,N_19859);
xnor UO_1266 (O_1266,N_19820,N_19972);
or UO_1267 (O_1267,N_19913,N_19931);
or UO_1268 (O_1268,N_19832,N_19804);
nor UO_1269 (O_1269,N_19936,N_19937);
and UO_1270 (O_1270,N_19812,N_19986);
nor UO_1271 (O_1271,N_19750,N_19894);
nor UO_1272 (O_1272,N_19949,N_19906);
and UO_1273 (O_1273,N_19821,N_19896);
and UO_1274 (O_1274,N_19841,N_19837);
nor UO_1275 (O_1275,N_19805,N_19913);
nor UO_1276 (O_1276,N_19904,N_19862);
nor UO_1277 (O_1277,N_19788,N_19927);
and UO_1278 (O_1278,N_19813,N_19779);
nand UO_1279 (O_1279,N_19901,N_19899);
and UO_1280 (O_1280,N_19967,N_19921);
nand UO_1281 (O_1281,N_19912,N_19860);
nor UO_1282 (O_1282,N_19787,N_19853);
or UO_1283 (O_1283,N_19795,N_19807);
nor UO_1284 (O_1284,N_19995,N_19912);
and UO_1285 (O_1285,N_19770,N_19888);
and UO_1286 (O_1286,N_19894,N_19928);
nor UO_1287 (O_1287,N_19990,N_19846);
and UO_1288 (O_1288,N_19871,N_19840);
and UO_1289 (O_1289,N_19877,N_19795);
and UO_1290 (O_1290,N_19765,N_19807);
nor UO_1291 (O_1291,N_19973,N_19881);
nor UO_1292 (O_1292,N_19924,N_19760);
xor UO_1293 (O_1293,N_19815,N_19935);
nor UO_1294 (O_1294,N_19829,N_19851);
xnor UO_1295 (O_1295,N_19782,N_19993);
or UO_1296 (O_1296,N_19913,N_19986);
nor UO_1297 (O_1297,N_19956,N_19753);
xnor UO_1298 (O_1298,N_19778,N_19782);
xor UO_1299 (O_1299,N_19798,N_19864);
xnor UO_1300 (O_1300,N_19802,N_19986);
xnor UO_1301 (O_1301,N_19848,N_19780);
nor UO_1302 (O_1302,N_19867,N_19786);
xnor UO_1303 (O_1303,N_19925,N_19863);
nand UO_1304 (O_1304,N_19956,N_19768);
or UO_1305 (O_1305,N_19996,N_19923);
nand UO_1306 (O_1306,N_19804,N_19872);
xnor UO_1307 (O_1307,N_19959,N_19931);
nand UO_1308 (O_1308,N_19804,N_19819);
nor UO_1309 (O_1309,N_19961,N_19783);
xor UO_1310 (O_1310,N_19880,N_19802);
xor UO_1311 (O_1311,N_19778,N_19913);
and UO_1312 (O_1312,N_19985,N_19912);
and UO_1313 (O_1313,N_19880,N_19903);
and UO_1314 (O_1314,N_19968,N_19958);
or UO_1315 (O_1315,N_19876,N_19826);
or UO_1316 (O_1316,N_19815,N_19764);
xor UO_1317 (O_1317,N_19924,N_19758);
or UO_1318 (O_1318,N_19834,N_19943);
nor UO_1319 (O_1319,N_19824,N_19885);
and UO_1320 (O_1320,N_19822,N_19973);
nor UO_1321 (O_1321,N_19930,N_19920);
and UO_1322 (O_1322,N_19957,N_19896);
and UO_1323 (O_1323,N_19768,N_19794);
nor UO_1324 (O_1324,N_19945,N_19857);
nand UO_1325 (O_1325,N_19825,N_19983);
or UO_1326 (O_1326,N_19988,N_19925);
xnor UO_1327 (O_1327,N_19969,N_19847);
nor UO_1328 (O_1328,N_19884,N_19861);
or UO_1329 (O_1329,N_19779,N_19968);
nand UO_1330 (O_1330,N_19816,N_19802);
and UO_1331 (O_1331,N_19763,N_19845);
and UO_1332 (O_1332,N_19762,N_19783);
nand UO_1333 (O_1333,N_19751,N_19967);
xor UO_1334 (O_1334,N_19951,N_19806);
or UO_1335 (O_1335,N_19812,N_19944);
nor UO_1336 (O_1336,N_19768,N_19796);
nand UO_1337 (O_1337,N_19778,N_19859);
xor UO_1338 (O_1338,N_19847,N_19970);
and UO_1339 (O_1339,N_19908,N_19919);
nand UO_1340 (O_1340,N_19947,N_19919);
xor UO_1341 (O_1341,N_19970,N_19875);
or UO_1342 (O_1342,N_19777,N_19755);
nand UO_1343 (O_1343,N_19837,N_19792);
and UO_1344 (O_1344,N_19904,N_19983);
nand UO_1345 (O_1345,N_19946,N_19959);
or UO_1346 (O_1346,N_19816,N_19974);
nand UO_1347 (O_1347,N_19839,N_19918);
nand UO_1348 (O_1348,N_19959,N_19807);
nor UO_1349 (O_1349,N_19839,N_19771);
xor UO_1350 (O_1350,N_19884,N_19987);
and UO_1351 (O_1351,N_19965,N_19981);
nand UO_1352 (O_1352,N_19983,N_19807);
nor UO_1353 (O_1353,N_19828,N_19803);
or UO_1354 (O_1354,N_19853,N_19847);
and UO_1355 (O_1355,N_19981,N_19971);
and UO_1356 (O_1356,N_19971,N_19836);
xor UO_1357 (O_1357,N_19799,N_19993);
nor UO_1358 (O_1358,N_19843,N_19942);
or UO_1359 (O_1359,N_19845,N_19791);
nor UO_1360 (O_1360,N_19753,N_19825);
xnor UO_1361 (O_1361,N_19905,N_19838);
nor UO_1362 (O_1362,N_19793,N_19882);
xnor UO_1363 (O_1363,N_19804,N_19833);
xnor UO_1364 (O_1364,N_19850,N_19828);
and UO_1365 (O_1365,N_19849,N_19856);
and UO_1366 (O_1366,N_19993,N_19831);
xor UO_1367 (O_1367,N_19868,N_19759);
nand UO_1368 (O_1368,N_19944,N_19899);
xor UO_1369 (O_1369,N_19918,N_19762);
or UO_1370 (O_1370,N_19894,N_19972);
xnor UO_1371 (O_1371,N_19858,N_19849);
or UO_1372 (O_1372,N_19812,N_19932);
nor UO_1373 (O_1373,N_19774,N_19780);
nor UO_1374 (O_1374,N_19926,N_19914);
or UO_1375 (O_1375,N_19997,N_19942);
nor UO_1376 (O_1376,N_19939,N_19862);
nand UO_1377 (O_1377,N_19839,N_19978);
xor UO_1378 (O_1378,N_19784,N_19941);
nand UO_1379 (O_1379,N_19762,N_19868);
xor UO_1380 (O_1380,N_19853,N_19796);
xnor UO_1381 (O_1381,N_19978,N_19873);
or UO_1382 (O_1382,N_19882,N_19907);
and UO_1383 (O_1383,N_19831,N_19963);
xnor UO_1384 (O_1384,N_19984,N_19764);
nor UO_1385 (O_1385,N_19778,N_19877);
nor UO_1386 (O_1386,N_19861,N_19781);
nor UO_1387 (O_1387,N_19978,N_19886);
xor UO_1388 (O_1388,N_19776,N_19753);
nor UO_1389 (O_1389,N_19801,N_19996);
nor UO_1390 (O_1390,N_19977,N_19773);
and UO_1391 (O_1391,N_19759,N_19913);
xnor UO_1392 (O_1392,N_19984,N_19879);
xor UO_1393 (O_1393,N_19920,N_19972);
or UO_1394 (O_1394,N_19993,N_19947);
nor UO_1395 (O_1395,N_19957,N_19832);
nor UO_1396 (O_1396,N_19988,N_19801);
or UO_1397 (O_1397,N_19918,N_19819);
or UO_1398 (O_1398,N_19797,N_19988);
xnor UO_1399 (O_1399,N_19861,N_19964);
or UO_1400 (O_1400,N_19862,N_19848);
nand UO_1401 (O_1401,N_19930,N_19885);
nand UO_1402 (O_1402,N_19986,N_19790);
xnor UO_1403 (O_1403,N_19847,N_19824);
nor UO_1404 (O_1404,N_19773,N_19793);
or UO_1405 (O_1405,N_19932,N_19991);
nor UO_1406 (O_1406,N_19990,N_19936);
nor UO_1407 (O_1407,N_19942,N_19813);
nor UO_1408 (O_1408,N_19959,N_19927);
or UO_1409 (O_1409,N_19784,N_19843);
nor UO_1410 (O_1410,N_19955,N_19830);
nor UO_1411 (O_1411,N_19928,N_19904);
nor UO_1412 (O_1412,N_19891,N_19978);
xnor UO_1413 (O_1413,N_19890,N_19962);
and UO_1414 (O_1414,N_19908,N_19889);
xnor UO_1415 (O_1415,N_19825,N_19877);
nor UO_1416 (O_1416,N_19938,N_19839);
or UO_1417 (O_1417,N_19852,N_19873);
xnor UO_1418 (O_1418,N_19808,N_19790);
nand UO_1419 (O_1419,N_19914,N_19867);
xnor UO_1420 (O_1420,N_19890,N_19935);
nor UO_1421 (O_1421,N_19917,N_19824);
nor UO_1422 (O_1422,N_19896,N_19774);
and UO_1423 (O_1423,N_19871,N_19883);
and UO_1424 (O_1424,N_19999,N_19810);
xor UO_1425 (O_1425,N_19944,N_19947);
nor UO_1426 (O_1426,N_19956,N_19807);
nand UO_1427 (O_1427,N_19990,N_19899);
xor UO_1428 (O_1428,N_19854,N_19938);
xor UO_1429 (O_1429,N_19968,N_19771);
and UO_1430 (O_1430,N_19903,N_19756);
nor UO_1431 (O_1431,N_19969,N_19779);
xnor UO_1432 (O_1432,N_19814,N_19859);
or UO_1433 (O_1433,N_19908,N_19853);
xor UO_1434 (O_1434,N_19953,N_19949);
xor UO_1435 (O_1435,N_19843,N_19797);
or UO_1436 (O_1436,N_19780,N_19896);
nand UO_1437 (O_1437,N_19790,N_19817);
and UO_1438 (O_1438,N_19990,N_19836);
or UO_1439 (O_1439,N_19946,N_19819);
or UO_1440 (O_1440,N_19896,N_19800);
and UO_1441 (O_1441,N_19975,N_19778);
nand UO_1442 (O_1442,N_19949,N_19885);
nand UO_1443 (O_1443,N_19839,N_19853);
and UO_1444 (O_1444,N_19865,N_19773);
nor UO_1445 (O_1445,N_19861,N_19828);
nand UO_1446 (O_1446,N_19918,N_19989);
nand UO_1447 (O_1447,N_19980,N_19899);
nand UO_1448 (O_1448,N_19980,N_19919);
and UO_1449 (O_1449,N_19877,N_19998);
xor UO_1450 (O_1450,N_19995,N_19901);
nand UO_1451 (O_1451,N_19855,N_19875);
nor UO_1452 (O_1452,N_19876,N_19964);
or UO_1453 (O_1453,N_19919,N_19772);
nor UO_1454 (O_1454,N_19854,N_19915);
nand UO_1455 (O_1455,N_19974,N_19965);
and UO_1456 (O_1456,N_19796,N_19812);
nand UO_1457 (O_1457,N_19933,N_19850);
or UO_1458 (O_1458,N_19769,N_19841);
nand UO_1459 (O_1459,N_19966,N_19945);
xnor UO_1460 (O_1460,N_19755,N_19859);
or UO_1461 (O_1461,N_19838,N_19882);
xor UO_1462 (O_1462,N_19838,N_19829);
or UO_1463 (O_1463,N_19923,N_19860);
nor UO_1464 (O_1464,N_19978,N_19896);
nand UO_1465 (O_1465,N_19898,N_19885);
or UO_1466 (O_1466,N_19985,N_19889);
and UO_1467 (O_1467,N_19900,N_19778);
or UO_1468 (O_1468,N_19836,N_19905);
and UO_1469 (O_1469,N_19773,N_19919);
nand UO_1470 (O_1470,N_19904,N_19994);
xnor UO_1471 (O_1471,N_19868,N_19876);
xnor UO_1472 (O_1472,N_19755,N_19787);
and UO_1473 (O_1473,N_19936,N_19924);
and UO_1474 (O_1474,N_19930,N_19788);
nand UO_1475 (O_1475,N_19887,N_19976);
xnor UO_1476 (O_1476,N_19865,N_19934);
nand UO_1477 (O_1477,N_19894,N_19780);
nor UO_1478 (O_1478,N_19785,N_19913);
and UO_1479 (O_1479,N_19852,N_19941);
or UO_1480 (O_1480,N_19966,N_19818);
or UO_1481 (O_1481,N_19905,N_19875);
and UO_1482 (O_1482,N_19808,N_19903);
xor UO_1483 (O_1483,N_19909,N_19928);
or UO_1484 (O_1484,N_19844,N_19858);
nand UO_1485 (O_1485,N_19852,N_19997);
xnor UO_1486 (O_1486,N_19818,N_19971);
or UO_1487 (O_1487,N_19868,N_19999);
xor UO_1488 (O_1488,N_19972,N_19772);
xnor UO_1489 (O_1489,N_19842,N_19968);
and UO_1490 (O_1490,N_19846,N_19829);
or UO_1491 (O_1491,N_19927,N_19778);
nor UO_1492 (O_1492,N_19887,N_19780);
xor UO_1493 (O_1493,N_19897,N_19785);
and UO_1494 (O_1494,N_19852,N_19954);
nor UO_1495 (O_1495,N_19923,N_19763);
nor UO_1496 (O_1496,N_19993,N_19853);
xnor UO_1497 (O_1497,N_19778,N_19902);
and UO_1498 (O_1498,N_19909,N_19781);
or UO_1499 (O_1499,N_19900,N_19828);
and UO_1500 (O_1500,N_19891,N_19814);
xor UO_1501 (O_1501,N_19819,N_19979);
xor UO_1502 (O_1502,N_19826,N_19821);
nand UO_1503 (O_1503,N_19928,N_19930);
or UO_1504 (O_1504,N_19945,N_19949);
nand UO_1505 (O_1505,N_19807,N_19812);
nor UO_1506 (O_1506,N_19968,N_19997);
or UO_1507 (O_1507,N_19769,N_19921);
or UO_1508 (O_1508,N_19984,N_19779);
nor UO_1509 (O_1509,N_19805,N_19811);
nor UO_1510 (O_1510,N_19997,N_19959);
nand UO_1511 (O_1511,N_19757,N_19898);
or UO_1512 (O_1512,N_19837,N_19775);
and UO_1513 (O_1513,N_19929,N_19765);
or UO_1514 (O_1514,N_19852,N_19969);
and UO_1515 (O_1515,N_19917,N_19864);
or UO_1516 (O_1516,N_19810,N_19783);
nand UO_1517 (O_1517,N_19889,N_19946);
and UO_1518 (O_1518,N_19851,N_19886);
nand UO_1519 (O_1519,N_19933,N_19903);
or UO_1520 (O_1520,N_19885,N_19871);
and UO_1521 (O_1521,N_19769,N_19792);
and UO_1522 (O_1522,N_19986,N_19758);
or UO_1523 (O_1523,N_19888,N_19889);
or UO_1524 (O_1524,N_19810,N_19998);
and UO_1525 (O_1525,N_19991,N_19862);
and UO_1526 (O_1526,N_19759,N_19829);
nand UO_1527 (O_1527,N_19757,N_19849);
nor UO_1528 (O_1528,N_19944,N_19999);
xor UO_1529 (O_1529,N_19815,N_19843);
nand UO_1530 (O_1530,N_19771,N_19919);
xor UO_1531 (O_1531,N_19891,N_19939);
and UO_1532 (O_1532,N_19887,N_19978);
nor UO_1533 (O_1533,N_19857,N_19836);
nor UO_1534 (O_1534,N_19992,N_19777);
xor UO_1535 (O_1535,N_19991,N_19794);
nor UO_1536 (O_1536,N_19979,N_19868);
xnor UO_1537 (O_1537,N_19818,N_19771);
or UO_1538 (O_1538,N_19961,N_19886);
or UO_1539 (O_1539,N_19939,N_19941);
xor UO_1540 (O_1540,N_19907,N_19947);
nor UO_1541 (O_1541,N_19977,N_19824);
nor UO_1542 (O_1542,N_19954,N_19753);
and UO_1543 (O_1543,N_19758,N_19832);
or UO_1544 (O_1544,N_19917,N_19859);
nand UO_1545 (O_1545,N_19838,N_19920);
nor UO_1546 (O_1546,N_19784,N_19915);
xor UO_1547 (O_1547,N_19774,N_19875);
and UO_1548 (O_1548,N_19912,N_19869);
or UO_1549 (O_1549,N_19996,N_19901);
or UO_1550 (O_1550,N_19960,N_19977);
and UO_1551 (O_1551,N_19821,N_19917);
nand UO_1552 (O_1552,N_19915,N_19767);
xor UO_1553 (O_1553,N_19901,N_19878);
nor UO_1554 (O_1554,N_19809,N_19969);
xor UO_1555 (O_1555,N_19939,N_19827);
xor UO_1556 (O_1556,N_19893,N_19878);
nand UO_1557 (O_1557,N_19932,N_19809);
xnor UO_1558 (O_1558,N_19951,N_19750);
xor UO_1559 (O_1559,N_19844,N_19845);
or UO_1560 (O_1560,N_19976,N_19806);
xor UO_1561 (O_1561,N_19812,N_19965);
nand UO_1562 (O_1562,N_19797,N_19873);
nand UO_1563 (O_1563,N_19800,N_19883);
xnor UO_1564 (O_1564,N_19817,N_19825);
or UO_1565 (O_1565,N_19927,N_19965);
nor UO_1566 (O_1566,N_19832,N_19895);
and UO_1567 (O_1567,N_19917,N_19913);
or UO_1568 (O_1568,N_19884,N_19878);
xor UO_1569 (O_1569,N_19912,N_19944);
and UO_1570 (O_1570,N_19780,N_19793);
or UO_1571 (O_1571,N_19763,N_19856);
or UO_1572 (O_1572,N_19777,N_19986);
xor UO_1573 (O_1573,N_19783,N_19794);
and UO_1574 (O_1574,N_19772,N_19980);
nor UO_1575 (O_1575,N_19893,N_19943);
xor UO_1576 (O_1576,N_19827,N_19761);
or UO_1577 (O_1577,N_19774,N_19861);
or UO_1578 (O_1578,N_19887,N_19935);
and UO_1579 (O_1579,N_19989,N_19867);
and UO_1580 (O_1580,N_19828,N_19798);
xor UO_1581 (O_1581,N_19865,N_19949);
nor UO_1582 (O_1582,N_19871,N_19889);
or UO_1583 (O_1583,N_19848,N_19860);
nand UO_1584 (O_1584,N_19857,N_19762);
and UO_1585 (O_1585,N_19928,N_19884);
and UO_1586 (O_1586,N_19756,N_19818);
and UO_1587 (O_1587,N_19857,N_19951);
or UO_1588 (O_1588,N_19946,N_19998);
and UO_1589 (O_1589,N_19823,N_19854);
xnor UO_1590 (O_1590,N_19980,N_19912);
and UO_1591 (O_1591,N_19915,N_19974);
or UO_1592 (O_1592,N_19917,N_19964);
xnor UO_1593 (O_1593,N_19777,N_19854);
nand UO_1594 (O_1594,N_19877,N_19937);
nor UO_1595 (O_1595,N_19882,N_19974);
nor UO_1596 (O_1596,N_19910,N_19900);
nor UO_1597 (O_1597,N_19831,N_19890);
nor UO_1598 (O_1598,N_19818,N_19783);
and UO_1599 (O_1599,N_19991,N_19777);
and UO_1600 (O_1600,N_19831,N_19770);
and UO_1601 (O_1601,N_19908,N_19864);
nand UO_1602 (O_1602,N_19754,N_19935);
xnor UO_1603 (O_1603,N_19789,N_19817);
or UO_1604 (O_1604,N_19970,N_19859);
and UO_1605 (O_1605,N_19947,N_19880);
or UO_1606 (O_1606,N_19878,N_19787);
nor UO_1607 (O_1607,N_19779,N_19939);
nor UO_1608 (O_1608,N_19908,N_19961);
nand UO_1609 (O_1609,N_19921,N_19836);
or UO_1610 (O_1610,N_19772,N_19824);
nand UO_1611 (O_1611,N_19980,N_19998);
xnor UO_1612 (O_1612,N_19829,N_19879);
and UO_1613 (O_1613,N_19897,N_19843);
nor UO_1614 (O_1614,N_19767,N_19889);
nor UO_1615 (O_1615,N_19916,N_19894);
xor UO_1616 (O_1616,N_19941,N_19850);
or UO_1617 (O_1617,N_19834,N_19886);
xnor UO_1618 (O_1618,N_19816,N_19930);
or UO_1619 (O_1619,N_19894,N_19758);
nor UO_1620 (O_1620,N_19980,N_19932);
nand UO_1621 (O_1621,N_19794,N_19914);
nand UO_1622 (O_1622,N_19932,N_19774);
nor UO_1623 (O_1623,N_19912,N_19874);
and UO_1624 (O_1624,N_19956,N_19805);
xnor UO_1625 (O_1625,N_19779,N_19774);
and UO_1626 (O_1626,N_19918,N_19924);
or UO_1627 (O_1627,N_19843,N_19780);
nand UO_1628 (O_1628,N_19915,N_19885);
xor UO_1629 (O_1629,N_19974,N_19840);
and UO_1630 (O_1630,N_19811,N_19904);
or UO_1631 (O_1631,N_19862,N_19913);
nand UO_1632 (O_1632,N_19900,N_19941);
xnor UO_1633 (O_1633,N_19984,N_19943);
nand UO_1634 (O_1634,N_19999,N_19949);
and UO_1635 (O_1635,N_19758,N_19932);
nand UO_1636 (O_1636,N_19965,N_19854);
and UO_1637 (O_1637,N_19958,N_19992);
nor UO_1638 (O_1638,N_19881,N_19784);
xor UO_1639 (O_1639,N_19923,N_19988);
xor UO_1640 (O_1640,N_19774,N_19833);
nor UO_1641 (O_1641,N_19965,N_19860);
xor UO_1642 (O_1642,N_19831,N_19966);
and UO_1643 (O_1643,N_19839,N_19987);
or UO_1644 (O_1644,N_19888,N_19873);
nand UO_1645 (O_1645,N_19766,N_19881);
xor UO_1646 (O_1646,N_19968,N_19973);
nor UO_1647 (O_1647,N_19812,N_19904);
and UO_1648 (O_1648,N_19982,N_19822);
xor UO_1649 (O_1649,N_19941,N_19758);
and UO_1650 (O_1650,N_19759,N_19852);
and UO_1651 (O_1651,N_19823,N_19817);
xor UO_1652 (O_1652,N_19750,N_19959);
nor UO_1653 (O_1653,N_19938,N_19952);
xor UO_1654 (O_1654,N_19981,N_19886);
xor UO_1655 (O_1655,N_19846,N_19812);
and UO_1656 (O_1656,N_19790,N_19853);
or UO_1657 (O_1657,N_19934,N_19961);
nand UO_1658 (O_1658,N_19891,N_19792);
or UO_1659 (O_1659,N_19758,N_19905);
and UO_1660 (O_1660,N_19880,N_19763);
nand UO_1661 (O_1661,N_19804,N_19840);
or UO_1662 (O_1662,N_19891,N_19955);
xnor UO_1663 (O_1663,N_19920,N_19821);
xnor UO_1664 (O_1664,N_19811,N_19831);
xnor UO_1665 (O_1665,N_19918,N_19967);
nand UO_1666 (O_1666,N_19879,N_19918);
nor UO_1667 (O_1667,N_19954,N_19856);
xnor UO_1668 (O_1668,N_19898,N_19824);
nand UO_1669 (O_1669,N_19994,N_19772);
and UO_1670 (O_1670,N_19805,N_19908);
nand UO_1671 (O_1671,N_19875,N_19798);
nand UO_1672 (O_1672,N_19810,N_19915);
and UO_1673 (O_1673,N_19824,N_19927);
xnor UO_1674 (O_1674,N_19838,N_19771);
or UO_1675 (O_1675,N_19883,N_19830);
or UO_1676 (O_1676,N_19973,N_19817);
or UO_1677 (O_1677,N_19917,N_19792);
and UO_1678 (O_1678,N_19976,N_19823);
nor UO_1679 (O_1679,N_19889,N_19828);
xnor UO_1680 (O_1680,N_19907,N_19977);
and UO_1681 (O_1681,N_19836,N_19846);
or UO_1682 (O_1682,N_19763,N_19786);
or UO_1683 (O_1683,N_19953,N_19782);
nor UO_1684 (O_1684,N_19818,N_19980);
nor UO_1685 (O_1685,N_19930,N_19934);
or UO_1686 (O_1686,N_19813,N_19849);
nor UO_1687 (O_1687,N_19914,N_19900);
nor UO_1688 (O_1688,N_19988,N_19832);
nor UO_1689 (O_1689,N_19972,N_19788);
and UO_1690 (O_1690,N_19915,N_19947);
nor UO_1691 (O_1691,N_19956,N_19791);
xor UO_1692 (O_1692,N_19782,N_19832);
or UO_1693 (O_1693,N_19965,N_19988);
nand UO_1694 (O_1694,N_19903,N_19931);
and UO_1695 (O_1695,N_19871,N_19886);
xnor UO_1696 (O_1696,N_19928,N_19960);
nor UO_1697 (O_1697,N_19908,N_19916);
and UO_1698 (O_1698,N_19914,N_19927);
nand UO_1699 (O_1699,N_19771,N_19878);
and UO_1700 (O_1700,N_19758,N_19940);
or UO_1701 (O_1701,N_19761,N_19798);
and UO_1702 (O_1702,N_19863,N_19853);
nor UO_1703 (O_1703,N_19964,N_19840);
or UO_1704 (O_1704,N_19945,N_19905);
xor UO_1705 (O_1705,N_19957,N_19779);
xnor UO_1706 (O_1706,N_19900,N_19861);
nor UO_1707 (O_1707,N_19860,N_19984);
or UO_1708 (O_1708,N_19972,N_19975);
or UO_1709 (O_1709,N_19851,N_19989);
nand UO_1710 (O_1710,N_19852,N_19858);
and UO_1711 (O_1711,N_19960,N_19879);
nor UO_1712 (O_1712,N_19835,N_19843);
or UO_1713 (O_1713,N_19923,N_19887);
xor UO_1714 (O_1714,N_19860,N_19902);
or UO_1715 (O_1715,N_19753,N_19837);
and UO_1716 (O_1716,N_19790,N_19991);
nor UO_1717 (O_1717,N_19999,N_19815);
and UO_1718 (O_1718,N_19908,N_19832);
nand UO_1719 (O_1719,N_19884,N_19759);
xnor UO_1720 (O_1720,N_19822,N_19817);
xor UO_1721 (O_1721,N_19937,N_19849);
nor UO_1722 (O_1722,N_19831,N_19844);
xor UO_1723 (O_1723,N_19855,N_19979);
nor UO_1724 (O_1724,N_19979,N_19930);
and UO_1725 (O_1725,N_19937,N_19876);
and UO_1726 (O_1726,N_19763,N_19968);
nor UO_1727 (O_1727,N_19971,N_19811);
xor UO_1728 (O_1728,N_19813,N_19856);
xnor UO_1729 (O_1729,N_19930,N_19981);
nor UO_1730 (O_1730,N_19829,N_19794);
xor UO_1731 (O_1731,N_19775,N_19751);
and UO_1732 (O_1732,N_19802,N_19884);
or UO_1733 (O_1733,N_19934,N_19991);
nand UO_1734 (O_1734,N_19889,N_19757);
or UO_1735 (O_1735,N_19963,N_19987);
xor UO_1736 (O_1736,N_19988,N_19866);
and UO_1737 (O_1737,N_19796,N_19994);
nor UO_1738 (O_1738,N_19914,N_19948);
xnor UO_1739 (O_1739,N_19832,N_19947);
or UO_1740 (O_1740,N_19784,N_19847);
xnor UO_1741 (O_1741,N_19789,N_19973);
nor UO_1742 (O_1742,N_19809,N_19793);
nand UO_1743 (O_1743,N_19855,N_19774);
nor UO_1744 (O_1744,N_19932,N_19979);
nand UO_1745 (O_1745,N_19753,N_19919);
xnor UO_1746 (O_1746,N_19777,N_19782);
and UO_1747 (O_1747,N_19946,N_19922);
nor UO_1748 (O_1748,N_19864,N_19804);
nand UO_1749 (O_1749,N_19900,N_19934);
or UO_1750 (O_1750,N_19775,N_19801);
nor UO_1751 (O_1751,N_19906,N_19792);
nor UO_1752 (O_1752,N_19822,N_19908);
nor UO_1753 (O_1753,N_19913,N_19930);
nand UO_1754 (O_1754,N_19860,N_19969);
and UO_1755 (O_1755,N_19848,N_19904);
nand UO_1756 (O_1756,N_19834,N_19811);
xnor UO_1757 (O_1757,N_19764,N_19819);
nand UO_1758 (O_1758,N_19974,N_19881);
or UO_1759 (O_1759,N_19759,N_19872);
or UO_1760 (O_1760,N_19753,N_19942);
nand UO_1761 (O_1761,N_19808,N_19945);
and UO_1762 (O_1762,N_19802,N_19890);
xnor UO_1763 (O_1763,N_19906,N_19772);
or UO_1764 (O_1764,N_19976,N_19853);
nor UO_1765 (O_1765,N_19751,N_19868);
nor UO_1766 (O_1766,N_19970,N_19766);
nand UO_1767 (O_1767,N_19859,N_19982);
xor UO_1768 (O_1768,N_19793,N_19829);
xor UO_1769 (O_1769,N_19926,N_19925);
nand UO_1770 (O_1770,N_19840,N_19954);
xor UO_1771 (O_1771,N_19925,N_19940);
and UO_1772 (O_1772,N_19871,N_19841);
or UO_1773 (O_1773,N_19830,N_19933);
nor UO_1774 (O_1774,N_19999,N_19780);
or UO_1775 (O_1775,N_19937,N_19911);
xnor UO_1776 (O_1776,N_19772,N_19790);
nand UO_1777 (O_1777,N_19938,N_19834);
and UO_1778 (O_1778,N_19821,N_19841);
xnor UO_1779 (O_1779,N_19827,N_19943);
and UO_1780 (O_1780,N_19841,N_19785);
nor UO_1781 (O_1781,N_19772,N_19911);
xor UO_1782 (O_1782,N_19924,N_19863);
nor UO_1783 (O_1783,N_19983,N_19793);
nand UO_1784 (O_1784,N_19894,N_19841);
or UO_1785 (O_1785,N_19970,N_19927);
and UO_1786 (O_1786,N_19936,N_19827);
xnor UO_1787 (O_1787,N_19799,N_19991);
xnor UO_1788 (O_1788,N_19921,N_19878);
nand UO_1789 (O_1789,N_19783,N_19816);
xor UO_1790 (O_1790,N_19895,N_19914);
or UO_1791 (O_1791,N_19956,N_19862);
xor UO_1792 (O_1792,N_19786,N_19865);
and UO_1793 (O_1793,N_19976,N_19776);
nand UO_1794 (O_1794,N_19904,N_19929);
or UO_1795 (O_1795,N_19761,N_19754);
nor UO_1796 (O_1796,N_19880,N_19931);
and UO_1797 (O_1797,N_19789,N_19917);
xnor UO_1798 (O_1798,N_19925,N_19875);
nand UO_1799 (O_1799,N_19994,N_19843);
and UO_1800 (O_1800,N_19965,N_19905);
nand UO_1801 (O_1801,N_19799,N_19912);
xor UO_1802 (O_1802,N_19822,N_19770);
nand UO_1803 (O_1803,N_19992,N_19953);
nor UO_1804 (O_1804,N_19820,N_19965);
and UO_1805 (O_1805,N_19801,N_19804);
or UO_1806 (O_1806,N_19844,N_19940);
or UO_1807 (O_1807,N_19814,N_19843);
xnor UO_1808 (O_1808,N_19920,N_19767);
nand UO_1809 (O_1809,N_19876,N_19940);
nand UO_1810 (O_1810,N_19927,N_19861);
xnor UO_1811 (O_1811,N_19865,N_19819);
or UO_1812 (O_1812,N_19799,N_19961);
nor UO_1813 (O_1813,N_19933,N_19898);
and UO_1814 (O_1814,N_19948,N_19833);
and UO_1815 (O_1815,N_19934,N_19980);
nor UO_1816 (O_1816,N_19955,N_19963);
or UO_1817 (O_1817,N_19834,N_19983);
xor UO_1818 (O_1818,N_19990,N_19926);
nand UO_1819 (O_1819,N_19785,N_19912);
and UO_1820 (O_1820,N_19946,N_19851);
nand UO_1821 (O_1821,N_19753,N_19857);
nor UO_1822 (O_1822,N_19774,N_19946);
or UO_1823 (O_1823,N_19914,N_19751);
and UO_1824 (O_1824,N_19870,N_19992);
xor UO_1825 (O_1825,N_19795,N_19767);
nor UO_1826 (O_1826,N_19994,N_19990);
and UO_1827 (O_1827,N_19815,N_19872);
nor UO_1828 (O_1828,N_19818,N_19772);
or UO_1829 (O_1829,N_19779,N_19866);
and UO_1830 (O_1830,N_19950,N_19982);
and UO_1831 (O_1831,N_19859,N_19844);
nand UO_1832 (O_1832,N_19889,N_19852);
xor UO_1833 (O_1833,N_19853,N_19923);
nor UO_1834 (O_1834,N_19921,N_19969);
nor UO_1835 (O_1835,N_19789,N_19826);
nand UO_1836 (O_1836,N_19876,N_19756);
nor UO_1837 (O_1837,N_19855,N_19899);
or UO_1838 (O_1838,N_19922,N_19844);
nand UO_1839 (O_1839,N_19759,N_19801);
and UO_1840 (O_1840,N_19938,N_19823);
nor UO_1841 (O_1841,N_19905,N_19883);
or UO_1842 (O_1842,N_19788,N_19990);
or UO_1843 (O_1843,N_19902,N_19768);
xor UO_1844 (O_1844,N_19951,N_19817);
or UO_1845 (O_1845,N_19832,N_19898);
nand UO_1846 (O_1846,N_19831,N_19836);
or UO_1847 (O_1847,N_19981,N_19872);
or UO_1848 (O_1848,N_19900,N_19838);
nand UO_1849 (O_1849,N_19999,N_19925);
xnor UO_1850 (O_1850,N_19962,N_19981);
nand UO_1851 (O_1851,N_19917,N_19807);
nand UO_1852 (O_1852,N_19808,N_19898);
xor UO_1853 (O_1853,N_19948,N_19888);
xnor UO_1854 (O_1854,N_19803,N_19947);
or UO_1855 (O_1855,N_19881,N_19940);
and UO_1856 (O_1856,N_19878,N_19943);
nand UO_1857 (O_1857,N_19808,N_19787);
or UO_1858 (O_1858,N_19918,N_19791);
nand UO_1859 (O_1859,N_19898,N_19752);
or UO_1860 (O_1860,N_19842,N_19878);
xnor UO_1861 (O_1861,N_19979,N_19762);
nor UO_1862 (O_1862,N_19866,N_19750);
xor UO_1863 (O_1863,N_19884,N_19809);
xnor UO_1864 (O_1864,N_19930,N_19775);
or UO_1865 (O_1865,N_19778,N_19934);
nand UO_1866 (O_1866,N_19887,N_19894);
and UO_1867 (O_1867,N_19773,N_19983);
nand UO_1868 (O_1868,N_19794,N_19827);
and UO_1869 (O_1869,N_19940,N_19954);
and UO_1870 (O_1870,N_19943,N_19903);
xnor UO_1871 (O_1871,N_19866,N_19878);
nand UO_1872 (O_1872,N_19940,N_19861);
or UO_1873 (O_1873,N_19806,N_19916);
nor UO_1874 (O_1874,N_19937,N_19807);
nand UO_1875 (O_1875,N_19752,N_19852);
nand UO_1876 (O_1876,N_19965,N_19803);
and UO_1877 (O_1877,N_19943,N_19918);
nand UO_1878 (O_1878,N_19990,N_19886);
or UO_1879 (O_1879,N_19935,N_19765);
and UO_1880 (O_1880,N_19944,N_19902);
nand UO_1881 (O_1881,N_19969,N_19881);
and UO_1882 (O_1882,N_19999,N_19801);
nand UO_1883 (O_1883,N_19952,N_19900);
xor UO_1884 (O_1884,N_19989,N_19839);
xnor UO_1885 (O_1885,N_19884,N_19892);
and UO_1886 (O_1886,N_19813,N_19836);
nand UO_1887 (O_1887,N_19920,N_19887);
nor UO_1888 (O_1888,N_19943,N_19824);
nor UO_1889 (O_1889,N_19860,N_19857);
xnor UO_1890 (O_1890,N_19760,N_19909);
nor UO_1891 (O_1891,N_19777,N_19850);
and UO_1892 (O_1892,N_19763,N_19802);
nor UO_1893 (O_1893,N_19774,N_19953);
or UO_1894 (O_1894,N_19899,N_19885);
nand UO_1895 (O_1895,N_19852,N_19893);
nand UO_1896 (O_1896,N_19898,N_19802);
and UO_1897 (O_1897,N_19959,N_19772);
xnor UO_1898 (O_1898,N_19992,N_19965);
xor UO_1899 (O_1899,N_19820,N_19798);
or UO_1900 (O_1900,N_19976,N_19861);
nand UO_1901 (O_1901,N_19985,N_19763);
and UO_1902 (O_1902,N_19887,N_19787);
xor UO_1903 (O_1903,N_19862,N_19855);
xor UO_1904 (O_1904,N_19827,N_19851);
or UO_1905 (O_1905,N_19841,N_19963);
nor UO_1906 (O_1906,N_19876,N_19759);
xnor UO_1907 (O_1907,N_19796,N_19973);
nor UO_1908 (O_1908,N_19793,N_19996);
nand UO_1909 (O_1909,N_19917,N_19991);
nand UO_1910 (O_1910,N_19885,N_19892);
xnor UO_1911 (O_1911,N_19795,N_19835);
nor UO_1912 (O_1912,N_19767,N_19936);
and UO_1913 (O_1913,N_19783,N_19887);
or UO_1914 (O_1914,N_19936,N_19964);
nand UO_1915 (O_1915,N_19976,N_19810);
or UO_1916 (O_1916,N_19815,N_19997);
or UO_1917 (O_1917,N_19896,N_19796);
nor UO_1918 (O_1918,N_19997,N_19981);
xnor UO_1919 (O_1919,N_19874,N_19923);
nand UO_1920 (O_1920,N_19992,N_19784);
xnor UO_1921 (O_1921,N_19908,N_19973);
nor UO_1922 (O_1922,N_19787,N_19776);
nor UO_1923 (O_1923,N_19876,N_19840);
and UO_1924 (O_1924,N_19813,N_19939);
xor UO_1925 (O_1925,N_19888,N_19988);
and UO_1926 (O_1926,N_19750,N_19897);
and UO_1927 (O_1927,N_19921,N_19997);
xor UO_1928 (O_1928,N_19799,N_19754);
nand UO_1929 (O_1929,N_19959,N_19860);
nor UO_1930 (O_1930,N_19981,N_19921);
nor UO_1931 (O_1931,N_19877,N_19950);
or UO_1932 (O_1932,N_19953,N_19760);
xnor UO_1933 (O_1933,N_19836,N_19824);
nor UO_1934 (O_1934,N_19850,N_19878);
nor UO_1935 (O_1935,N_19898,N_19841);
or UO_1936 (O_1936,N_19882,N_19855);
or UO_1937 (O_1937,N_19834,N_19995);
nor UO_1938 (O_1938,N_19810,N_19905);
and UO_1939 (O_1939,N_19931,N_19808);
nor UO_1940 (O_1940,N_19982,N_19998);
and UO_1941 (O_1941,N_19789,N_19837);
or UO_1942 (O_1942,N_19992,N_19858);
nand UO_1943 (O_1943,N_19785,N_19907);
xor UO_1944 (O_1944,N_19886,N_19985);
xor UO_1945 (O_1945,N_19948,N_19960);
and UO_1946 (O_1946,N_19806,N_19779);
nor UO_1947 (O_1947,N_19839,N_19868);
or UO_1948 (O_1948,N_19833,N_19931);
nand UO_1949 (O_1949,N_19975,N_19842);
and UO_1950 (O_1950,N_19845,N_19949);
and UO_1951 (O_1951,N_19928,N_19984);
and UO_1952 (O_1952,N_19951,N_19998);
nand UO_1953 (O_1953,N_19856,N_19831);
nor UO_1954 (O_1954,N_19998,N_19979);
nand UO_1955 (O_1955,N_19878,N_19810);
and UO_1956 (O_1956,N_19980,N_19835);
nand UO_1957 (O_1957,N_19986,N_19822);
xor UO_1958 (O_1958,N_19984,N_19897);
and UO_1959 (O_1959,N_19819,N_19792);
and UO_1960 (O_1960,N_19832,N_19836);
nand UO_1961 (O_1961,N_19903,N_19902);
and UO_1962 (O_1962,N_19996,N_19904);
nand UO_1963 (O_1963,N_19956,N_19843);
nand UO_1964 (O_1964,N_19889,N_19851);
and UO_1965 (O_1965,N_19815,N_19801);
xnor UO_1966 (O_1966,N_19894,N_19905);
nand UO_1967 (O_1967,N_19865,N_19762);
and UO_1968 (O_1968,N_19921,N_19853);
nor UO_1969 (O_1969,N_19923,N_19788);
or UO_1970 (O_1970,N_19907,N_19771);
and UO_1971 (O_1971,N_19881,N_19763);
xnor UO_1972 (O_1972,N_19941,N_19958);
xor UO_1973 (O_1973,N_19917,N_19780);
nand UO_1974 (O_1974,N_19888,N_19967);
or UO_1975 (O_1975,N_19792,N_19754);
and UO_1976 (O_1976,N_19792,N_19774);
xor UO_1977 (O_1977,N_19861,N_19962);
and UO_1978 (O_1978,N_19992,N_19917);
xnor UO_1979 (O_1979,N_19895,N_19761);
or UO_1980 (O_1980,N_19799,N_19750);
nor UO_1981 (O_1981,N_19888,N_19763);
nor UO_1982 (O_1982,N_19995,N_19784);
xnor UO_1983 (O_1983,N_19812,N_19914);
nor UO_1984 (O_1984,N_19752,N_19932);
and UO_1985 (O_1985,N_19866,N_19865);
or UO_1986 (O_1986,N_19751,N_19792);
or UO_1987 (O_1987,N_19918,N_19827);
and UO_1988 (O_1988,N_19908,N_19900);
nor UO_1989 (O_1989,N_19750,N_19882);
nand UO_1990 (O_1990,N_19916,N_19857);
nor UO_1991 (O_1991,N_19823,N_19917);
and UO_1992 (O_1992,N_19946,N_19967);
or UO_1993 (O_1993,N_19763,N_19940);
xnor UO_1994 (O_1994,N_19919,N_19778);
nand UO_1995 (O_1995,N_19939,N_19879);
or UO_1996 (O_1996,N_19756,N_19902);
or UO_1997 (O_1997,N_19895,N_19913);
and UO_1998 (O_1998,N_19936,N_19976);
and UO_1999 (O_1999,N_19987,N_19878);
or UO_2000 (O_2000,N_19777,N_19894);
nor UO_2001 (O_2001,N_19795,N_19774);
nor UO_2002 (O_2002,N_19860,N_19878);
nor UO_2003 (O_2003,N_19972,N_19878);
xor UO_2004 (O_2004,N_19943,N_19923);
xor UO_2005 (O_2005,N_19902,N_19793);
xor UO_2006 (O_2006,N_19830,N_19954);
and UO_2007 (O_2007,N_19778,N_19758);
and UO_2008 (O_2008,N_19792,N_19768);
or UO_2009 (O_2009,N_19808,N_19788);
xnor UO_2010 (O_2010,N_19971,N_19762);
and UO_2011 (O_2011,N_19790,N_19934);
nand UO_2012 (O_2012,N_19948,N_19983);
and UO_2013 (O_2013,N_19820,N_19780);
and UO_2014 (O_2014,N_19769,N_19890);
nand UO_2015 (O_2015,N_19751,N_19958);
or UO_2016 (O_2016,N_19974,N_19849);
xnor UO_2017 (O_2017,N_19846,N_19930);
or UO_2018 (O_2018,N_19762,N_19755);
xor UO_2019 (O_2019,N_19845,N_19764);
xnor UO_2020 (O_2020,N_19916,N_19912);
xor UO_2021 (O_2021,N_19847,N_19921);
or UO_2022 (O_2022,N_19977,N_19998);
or UO_2023 (O_2023,N_19788,N_19867);
nand UO_2024 (O_2024,N_19766,N_19857);
and UO_2025 (O_2025,N_19768,N_19885);
nand UO_2026 (O_2026,N_19769,N_19828);
and UO_2027 (O_2027,N_19968,N_19862);
and UO_2028 (O_2028,N_19983,N_19779);
nor UO_2029 (O_2029,N_19919,N_19935);
xor UO_2030 (O_2030,N_19887,N_19860);
nand UO_2031 (O_2031,N_19950,N_19771);
nor UO_2032 (O_2032,N_19821,N_19767);
nand UO_2033 (O_2033,N_19930,N_19954);
and UO_2034 (O_2034,N_19890,N_19917);
nand UO_2035 (O_2035,N_19862,N_19787);
xor UO_2036 (O_2036,N_19812,N_19952);
or UO_2037 (O_2037,N_19996,N_19820);
or UO_2038 (O_2038,N_19821,N_19895);
nor UO_2039 (O_2039,N_19907,N_19975);
nand UO_2040 (O_2040,N_19966,N_19809);
nand UO_2041 (O_2041,N_19839,N_19761);
and UO_2042 (O_2042,N_19795,N_19876);
and UO_2043 (O_2043,N_19997,N_19766);
nor UO_2044 (O_2044,N_19950,N_19977);
and UO_2045 (O_2045,N_19950,N_19887);
and UO_2046 (O_2046,N_19788,N_19975);
and UO_2047 (O_2047,N_19993,N_19941);
nor UO_2048 (O_2048,N_19885,N_19821);
or UO_2049 (O_2049,N_19761,N_19831);
xor UO_2050 (O_2050,N_19873,N_19827);
and UO_2051 (O_2051,N_19820,N_19870);
nor UO_2052 (O_2052,N_19820,N_19951);
nor UO_2053 (O_2053,N_19759,N_19994);
nor UO_2054 (O_2054,N_19977,N_19866);
and UO_2055 (O_2055,N_19836,N_19803);
or UO_2056 (O_2056,N_19875,N_19886);
xnor UO_2057 (O_2057,N_19814,N_19996);
xnor UO_2058 (O_2058,N_19964,N_19931);
nor UO_2059 (O_2059,N_19943,N_19960);
or UO_2060 (O_2060,N_19932,N_19865);
nor UO_2061 (O_2061,N_19887,N_19902);
and UO_2062 (O_2062,N_19909,N_19808);
xnor UO_2063 (O_2063,N_19896,N_19937);
and UO_2064 (O_2064,N_19923,N_19779);
and UO_2065 (O_2065,N_19754,N_19841);
xor UO_2066 (O_2066,N_19869,N_19919);
and UO_2067 (O_2067,N_19869,N_19794);
xor UO_2068 (O_2068,N_19790,N_19766);
or UO_2069 (O_2069,N_19934,N_19842);
xor UO_2070 (O_2070,N_19833,N_19824);
and UO_2071 (O_2071,N_19763,N_19795);
xor UO_2072 (O_2072,N_19883,N_19907);
nand UO_2073 (O_2073,N_19901,N_19762);
or UO_2074 (O_2074,N_19763,N_19783);
xnor UO_2075 (O_2075,N_19973,N_19914);
nor UO_2076 (O_2076,N_19950,N_19916);
xor UO_2077 (O_2077,N_19778,N_19946);
nand UO_2078 (O_2078,N_19954,N_19815);
and UO_2079 (O_2079,N_19968,N_19801);
nand UO_2080 (O_2080,N_19950,N_19781);
nor UO_2081 (O_2081,N_19844,N_19767);
xor UO_2082 (O_2082,N_19883,N_19977);
and UO_2083 (O_2083,N_19792,N_19812);
or UO_2084 (O_2084,N_19870,N_19760);
and UO_2085 (O_2085,N_19852,N_19835);
or UO_2086 (O_2086,N_19811,N_19861);
or UO_2087 (O_2087,N_19823,N_19893);
nand UO_2088 (O_2088,N_19925,N_19854);
or UO_2089 (O_2089,N_19751,N_19840);
or UO_2090 (O_2090,N_19758,N_19922);
or UO_2091 (O_2091,N_19802,N_19966);
xnor UO_2092 (O_2092,N_19876,N_19885);
nand UO_2093 (O_2093,N_19890,N_19819);
or UO_2094 (O_2094,N_19994,N_19913);
nor UO_2095 (O_2095,N_19976,N_19759);
xor UO_2096 (O_2096,N_19826,N_19933);
nand UO_2097 (O_2097,N_19982,N_19791);
xnor UO_2098 (O_2098,N_19969,N_19802);
nand UO_2099 (O_2099,N_19890,N_19821);
nand UO_2100 (O_2100,N_19759,N_19779);
and UO_2101 (O_2101,N_19905,N_19805);
xor UO_2102 (O_2102,N_19762,N_19824);
nor UO_2103 (O_2103,N_19944,N_19925);
or UO_2104 (O_2104,N_19776,N_19978);
xnor UO_2105 (O_2105,N_19849,N_19751);
nor UO_2106 (O_2106,N_19786,N_19892);
and UO_2107 (O_2107,N_19820,N_19915);
nor UO_2108 (O_2108,N_19828,N_19755);
nor UO_2109 (O_2109,N_19997,N_19827);
nor UO_2110 (O_2110,N_19779,N_19827);
nand UO_2111 (O_2111,N_19791,N_19888);
or UO_2112 (O_2112,N_19914,N_19899);
xor UO_2113 (O_2113,N_19851,N_19898);
xor UO_2114 (O_2114,N_19871,N_19969);
xor UO_2115 (O_2115,N_19912,N_19891);
xnor UO_2116 (O_2116,N_19926,N_19850);
and UO_2117 (O_2117,N_19880,N_19807);
and UO_2118 (O_2118,N_19953,N_19850);
xnor UO_2119 (O_2119,N_19813,N_19888);
or UO_2120 (O_2120,N_19774,N_19828);
nand UO_2121 (O_2121,N_19923,N_19958);
xor UO_2122 (O_2122,N_19759,N_19991);
and UO_2123 (O_2123,N_19875,N_19839);
xor UO_2124 (O_2124,N_19798,N_19997);
nand UO_2125 (O_2125,N_19847,N_19830);
xor UO_2126 (O_2126,N_19778,N_19781);
xnor UO_2127 (O_2127,N_19947,N_19998);
or UO_2128 (O_2128,N_19824,N_19801);
xor UO_2129 (O_2129,N_19914,N_19779);
and UO_2130 (O_2130,N_19808,N_19889);
xor UO_2131 (O_2131,N_19833,N_19907);
nor UO_2132 (O_2132,N_19877,N_19898);
xor UO_2133 (O_2133,N_19896,N_19999);
xnor UO_2134 (O_2134,N_19882,N_19953);
and UO_2135 (O_2135,N_19877,N_19926);
xor UO_2136 (O_2136,N_19875,N_19955);
xor UO_2137 (O_2137,N_19786,N_19759);
and UO_2138 (O_2138,N_19967,N_19836);
xnor UO_2139 (O_2139,N_19967,N_19840);
nand UO_2140 (O_2140,N_19989,N_19764);
nand UO_2141 (O_2141,N_19932,N_19850);
nor UO_2142 (O_2142,N_19773,N_19972);
nand UO_2143 (O_2143,N_19777,N_19848);
or UO_2144 (O_2144,N_19868,N_19934);
xnor UO_2145 (O_2145,N_19937,N_19979);
or UO_2146 (O_2146,N_19805,N_19984);
nor UO_2147 (O_2147,N_19853,N_19851);
nor UO_2148 (O_2148,N_19821,N_19869);
or UO_2149 (O_2149,N_19848,N_19954);
and UO_2150 (O_2150,N_19773,N_19752);
nor UO_2151 (O_2151,N_19770,N_19868);
nor UO_2152 (O_2152,N_19869,N_19867);
and UO_2153 (O_2153,N_19907,N_19890);
xor UO_2154 (O_2154,N_19826,N_19881);
nand UO_2155 (O_2155,N_19773,N_19948);
and UO_2156 (O_2156,N_19786,N_19958);
nor UO_2157 (O_2157,N_19936,N_19795);
and UO_2158 (O_2158,N_19985,N_19974);
nand UO_2159 (O_2159,N_19835,N_19915);
or UO_2160 (O_2160,N_19899,N_19783);
and UO_2161 (O_2161,N_19972,N_19858);
or UO_2162 (O_2162,N_19906,N_19845);
xnor UO_2163 (O_2163,N_19828,N_19794);
nand UO_2164 (O_2164,N_19793,N_19989);
nand UO_2165 (O_2165,N_19913,N_19887);
nand UO_2166 (O_2166,N_19859,N_19766);
nor UO_2167 (O_2167,N_19803,N_19793);
xor UO_2168 (O_2168,N_19915,N_19800);
nand UO_2169 (O_2169,N_19976,N_19802);
nand UO_2170 (O_2170,N_19782,N_19849);
nor UO_2171 (O_2171,N_19851,N_19935);
xnor UO_2172 (O_2172,N_19960,N_19915);
nor UO_2173 (O_2173,N_19871,N_19930);
and UO_2174 (O_2174,N_19752,N_19935);
or UO_2175 (O_2175,N_19812,N_19900);
and UO_2176 (O_2176,N_19916,N_19787);
nand UO_2177 (O_2177,N_19752,N_19921);
or UO_2178 (O_2178,N_19975,N_19961);
nor UO_2179 (O_2179,N_19834,N_19997);
nand UO_2180 (O_2180,N_19957,N_19886);
nand UO_2181 (O_2181,N_19859,N_19943);
or UO_2182 (O_2182,N_19792,N_19755);
xor UO_2183 (O_2183,N_19820,N_19878);
and UO_2184 (O_2184,N_19861,N_19831);
xnor UO_2185 (O_2185,N_19775,N_19819);
and UO_2186 (O_2186,N_19894,N_19918);
and UO_2187 (O_2187,N_19971,N_19926);
xnor UO_2188 (O_2188,N_19915,N_19778);
nand UO_2189 (O_2189,N_19881,N_19959);
nand UO_2190 (O_2190,N_19941,N_19978);
nand UO_2191 (O_2191,N_19812,N_19861);
and UO_2192 (O_2192,N_19869,N_19927);
nor UO_2193 (O_2193,N_19787,N_19970);
and UO_2194 (O_2194,N_19938,N_19906);
nor UO_2195 (O_2195,N_19906,N_19828);
or UO_2196 (O_2196,N_19809,N_19995);
and UO_2197 (O_2197,N_19850,N_19906);
nand UO_2198 (O_2198,N_19875,N_19883);
nor UO_2199 (O_2199,N_19800,N_19804);
and UO_2200 (O_2200,N_19819,N_19896);
nor UO_2201 (O_2201,N_19979,N_19851);
and UO_2202 (O_2202,N_19978,N_19788);
nor UO_2203 (O_2203,N_19817,N_19842);
xor UO_2204 (O_2204,N_19847,N_19999);
nor UO_2205 (O_2205,N_19817,N_19872);
nand UO_2206 (O_2206,N_19794,N_19932);
or UO_2207 (O_2207,N_19834,N_19904);
nor UO_2208 (O_2208,N_19767,N_19856);
and UO_2209 (O_2209,N_19898,N_19819);
xor UO_2210 (O_2210,N_19785,N_19895);
nor UO_2211 (O_2211,N_19761,N_19786);
or UO_2212 (O_2212,N_19802,N_19971);
xor UO_2213 (O_2213,N_19938,N_19775);
or UO_2214 (O_2214,N_19791,N_19908);
nand UO_2215 (O_2215,N_19929,N_19844);
nor UO_2216 (O_2216,N_19829,N_19781);
or UO_2217 (O_2217,N_19903,N_19835);
or UO_2218 (O_2218,N_19831,N_19829);
xnor UO_2219 (O_2219,N_19875,N_19914);
xor UO_2220 (O_2220,N_19845,N_19862);
xnor UO_2221 (O_2221,N_19965,N_19940);
or UO_2222 (O_2222,N_19986,N_19974);
nor UO_2223 (O_2223,N_19753,N_19788);
xor UO_2224 (O_2224,N_19908,N_19793);
xnor UO_2225 (O_2225,N_19768,N_19798);
or UO_2226 (O_2226,N_19783,N_19956);
nand UO_2227 (O_2227,N_19883,N_19889);
xnor UO_2228 (O_2228,N_19908,N_19871);
xor UO_2229 (O_2229,N_19924,N_19879);
nor UO_2230 (O_2230,N_19944,N_19811);
or UO_2231 (O_2231,N_19955,N_19995);
nor UO_2232 (O_2232,N_19830,N_19897);
and UO_2233 (O_2233,N_19798,N_19958);
nor UO_2234 (O_2234,N_19819,N_19953);
xor UO_2235 (O_2235,N_19856,N_19914);
nand UO_2236 (O_2236,N_19948,N_19890);
and UO_2237 (O_2237,N_19823,N_19837);
nand UO_2238 (O_2238,N_19934,N_19929);
and UO_2239 (O_2239,N_19966,N_19957);
xor UO_2240 (O_2240,N_19968,N_19974);
xor UO_2241 (O_2241,N_19882,N_19879);
nor UO_2242 (O_2242,N_19928,N_19936);
nand UO_2243 (O_2243,N_19765,N_19964);
xnor UO_2244 (O_2244,N_19851,N_19821);
nor UO_2245 (O_2245,N_19809,N_19897);
nand UO_2246 (O_2246,N_19811,N_19827);
nor UO_2247 (O_2247,N_19918,N_19950);
nor UO_2248 (O_2248,N_19978,N_19775);
or UO_2249 (O_2249,N_19958,N_19865);
xor UO_2250 (O_2250,N_19888,N_19987);
xnor UO_2251 (O_2251,N_19985,N_19764);
or UO_2252 (O_2252,N_19772,N_19918);
nand UO_2253 (O_2253,N_19882,N_19930);
xor UO_2254 (O_2254,N_19914,N_19936);
xnor UO_2255 (O_2255,N_19933,N_19881);
and UO_2256 (O_2256,N_19965,N_19945);
nor UO_2257 (O_2257,N_19916,N_19825);
and UO_2258 (O_2258,N_19762,N_19853);
nor UO_2259 (O_2259,N_19808,N_19758);
nor UO_2260 (O_2260,N_19915,N_19803);
and UO_2261 (O_2261,N_19944,N_19870);
nand UO_2262 (O_2262,N_19753,N_19930);
and UO_2263 (O_2263,N_19921,N_19863);
nand UO_2264 (O_2264,N_19805,N_19881);
nand UO_2265 (O_2265,N_19836,N_19901);
nand UO_2266 (O_2266,N_19873,N_19994);
nor UO_2267 (O_2267,N_19964,N_19777);
nor UO_2268 (O_2268,N_19990,N_19998);
nor UO_2269 (O_2269,N_19900,N_19833);
nand UO_2270 (O_2270,N_19932,N_19931);
or UO_2271 (O_2271,N_19873,N_19806);
and UO_2272 (O_2272,N_19910,N_19808);
nor UO_2273 (O_2273,N_19788,N_19795);
and UO_2274 (O_2274,N_19893,N_19807);
and UO_2275 (O_2275,N_19771,N_19866);
nor UO_2276 (O_2276,N_19811,N_19973);
nand UO_2277 (O_2277,N_19983,N_19887);
or UO_2278 (O_2278,N_19991,N_19768);
and UO_2279 (O_2279,N_19994,N_19997);
nand UO_2280 (O_2280,N_19776,N_19885);
or UO_2281 (O_2281,N_19814,N_19877);
xnor UO_2282 (O_2282,N_19809,N_19756);
nor UO_2283 (O_2283,N_19772,N_19792);
xor UO_2284 (O_2284,N_19903,N_19911);
or UO_2285 (O_2285,N_19899,N_19941);
nor UO_2286 (O_2286,N_19962,N_19851);
nor UO_2287 (O_2287,N_19928,N_19945);
or UO_2288 (O_2288,N_19785,N_19875);
or UO_2289 (O_2289,N_19951,N_19785);
and UO_2290 (O_2290,N_19804,N_19865);
nand UO_2291 (O_2291,N_19978,N_19954);
and UO_2292 (O_2292,N_19908,N_19786);
nor UO_2293 (O_2293,N_19833,N_19899);
nand UO_2294 (O_2294,N_19754,N_19759);
xor UO_2295 (O_2295,N_19990,N_19999);
nor UO_2296 (O_2296,N_19984,N_19935);
nand UO_2297 (O_2297,N_19946,N_19936);
and UO_2298 (O_2298,N_19884,N_19891);
and UO_2299 (O_2299,N_19947,N_19913);
or UO_2300 (O_2300,N_19877,N_19904);
nand UO_2301 (O_2301,N_19828,N_19953);
nand UO_2302 (O_2302,N_19836,N_19777);
nor UO_2303 (O_2303,N_19779,N_19773);
and UO_2304 (O_2304,N_19876,N_19892);
or UO_2305 (O_2305,N_19977,N_19841);
or UO_2306 (O_2306,N_19894,N_19783);
or UO_2307 (O_2307,N_19851,N_19871);
nor UO_2308 (O_2308,N_19913,N_19837);
xor UO_2309 (O_2309,N_19812,N_19935);
or UO_2310 (O_2310,N_19922,N_19882);
nand UO_2311 (O_2311,N_19867,N_19906);
and UO_2312 (O_2312,N_19868,N_19889);
nor UO_2313 (O_2313,N_19943,N_19839);
and UO_2314 (O_2314,N_19764,N_19900);
xor UO_2315 (O_2315,N_19869,N_19873);
nand UO_2316 (O_2316,N_19834,N_19898);
and UO_2317 (O_2317,N_19868,N_19805);
nor UO_2318 (O_2318,N_19907,N_19979);
or UO_2319 (O_2319,N_19834,N_19864);
or UO_2320 (O_2320,N_19815,N_19959);
nand UO_2321 (O_2321,N_19824,N_19750);
xor UO_2322 (O_2322,N_19812,N_19928);
or UO_2323 (O_2323,N_19881,N_19917);
nor UO_2324 (O_2324,N_19860,N_19796);
nor UO_2325 (O_2325,N_19828,N_19924);
xor UO_2326 (O_2326,N_19963,N_19942);
and UO_2327 (O_2327,N_19807,N_19761);
nand UO_2328 (O_2328,N_19816,N_19822);
nor UO_2329 (O_2329,N_19932,N_19797);
nand UO_2330 (O_2330,N_19830,N_19792);
nand UO_2331 (O_2331,N_19759,N_19809);
xnor UO_2332 (O_2332,N_19772,N_19795);
nor UO_2333 (O_2333,N_19930,N_19758);
nor UO_2334 (O_2334,N_19945,N_19866);
xnor UO_2335 (O_2335,N_19967,N_19866);
nor UO_2336 (O_2336,N_19983,N_19939);
nor UO_2337 (O_2337,N_19890,N_19878);
or UO_2338 (O_2338,N_19775,N_19834);
and UO_2339 (O_2339,N_19924,N_19841);
nand UO_2340 (O_2340,N_19960,N_19857);
xnor UO_2341 (O_2341,N_19995,N_19887);
or UO_2342 (O_2342,N_19780,N_19815);
xnor UO_2343 (O_2343,N_19791,N_19927);
and UO_2344 (O_2344,N_19820,N_19810);
or UO_2345 (O_2345,N_19954,N_19974);
nand UO_2346 (O_2346,N_19822,N_19811);
nor UO_2347 (O_2347,N_19804,N_19974);
nor UO_2348 (O_2348,N_19822,N_19984);
or UO_2349 (O_2349,N_19923,N_19888);
or UO_2350 (O_2350,N_19827,N_19790);
or UO_2351 (O_2351,N_19941,N_19940);
nand UO_2352 (O_2352,N_19893,N_19762);
xor UO_2353 (O_2353,N_19980,N_19949);
and UO_2354 (O_2354,N_19770,N_19782);
and UO_2355 (O_2355,N_19843,N_19967);
nand UO_2356 (O_2356,N_19783,N_19984);
or UO_2357 (O_2357,N_19984,N_19978);
nor UO_2358 (O_2358,N_19937,N_19808);
xnor UO_2359 (O_2359,N_19781,N_19902);
and UO_2360 (O_2360,N_19967,N_19912);
nand UO_2361 (O_2361,N_19895,N_19770);
nor UO_2362 (O_2362,N_19989,N_19961);
nor UO_2363 (O_2363,N_19815,N_19851);
xor UO_2364 (O_2364,N_19810,N_19888);
and UO_2365 (O_2365,N_19988,N_19792);
and UO_2366 (O_2366,N_19797,N_19799);
xor UO_2367 (O_2367,N_19861,N_19789);
or UO_2368 (O_2368,N_19953,N_19856);
nand UO_2369 (O_2369,N_19968,N_19894);
or UO_2370 (O_2370,N_19777,N_19997);
xor UO_2371 (O_2371,N_19770,N_19883);
nor UO_2372 (O_2372,N_19960,N_19889);
and UO_2373 (O_2373,N_19763,N_19869);
or UO_2374 (O_2374,N_19770,N_19869);
nand UO_2375 (O_2375,N_19786,N_19801);
and UO_2376 (O_2376,N_19806,N_19808);
nand UO_2377 (O_2377,N_19955,N_19867);
xor UO_2378 (O_2378,N_19927,N_19850);
xor UO_2379 (O_2379,N_19799,N_19933);
xor UO_2380 (O_2380,N_19777,N_19957);
and UO_2381 (O_2381,N_19880,N_19872);
xnor UO_2382 (O_2382,N_19833,N_19985);
or UO_2383 (O_2383,N_19971,N_19856);
or UO_2384 (O_2384,N_19855,N_19765);
xor UO_2385 (O_2385,N_19952,N_19761);
xor UO_2386 (O_2386,N_19978,N_19956);
nor UO_2387 (O_2387,N_19991,N_19936);
nor UO_2388 (O_2388,N_19858,N_19958);
xor UO_2389 (O_2389,N_19814,N_19949);
nor UO_2390 (O_2390,N_19918,N_19771);
or UO_2391 (O_2391,N_19822,N_19884);
and UO_2392 (O_2392,N_19802,N_19804);
nand UO_2393 (O_2393,N_19864,N_19759);
nor UO_2394 (O_2394,N_19976,N_19800);
nor UO_2395 (O_2395,N_19760,N_19906);
or UO_2396 (O_2396,N_19874,N_19910);
and UO_2397 (O_2397,N_19995,N_19844);
and UO_2398 (O_2398,N_19849,N_19979);
nand UO_2399 (O_2399,N_19826,N_19842);
xnor UO_2400 (O_2400,N_19808,N_19814);
xor UO_2401 (O_2401,N_19788,N_19823);
or UO_2402 (O_2402,N_19861,N_19955);
or UO_2403 (O_2403,N_19956,N_19987);
xnor UO_2404 (O_2404,N_19971,N_19796);
and UO_2405 (O_2405,N_19886,N_19867);
or UO_2406 (O_2406,N_19979,N_19885);
nor UO_2407 (O_2407,N_19886,N_19905);
nor UO_2408 (O_2408,N_19848,N_19786);
nand UO_2409 (O_2409,N_19866,N_19758);
or UO_2410 (O_2410,N_19775,N_19866);
or UO_2411 (O_2411,N_19849,N_19904);
xnor UO_2412 (O_2412,N_19859,N_19933);
or UO_2413 (O_2413,N_19767,N_19806);
and UO_2414 (O_2414,N_19962,N_19793);
xor UO_2415 (O_2415,N_19757,N_19963);
nand UO_2416 (O_2416,N_19869,N_19815);
or UO_2417 (O_2417,N_19752,N_19782);
nor UO_2418 (O_2418,N_19911,N_19840);
xor UO_2419 (O_2419,N_19812,N_19920);
xor UO_2420 (O_2420,N_19752,N_19976);
and UO_2421 (O_2421,N_19926,N_19824);
nand UO_2422 (O_2422,N_19848,N_19929);
nand UO_2423 (O_2423,N_19971,N_19907);
or UO_2424 (O_2424,N_19960,N_19992);
and UO_2425 (O_2425,N_19905,N_19785);
nor UO_2426 (O_2426,N_19989,N_19933);
and UO_2427 (O_2427,N_19806,N_19960);
xnor UO_2428 (O_2428,N_19949,N_19891);
xnor UO_2429 (O_2429,N_19891,N_19920);
nor UO_2430 (O_2430,N_19856,N_19908);
nor UO_2431 (O_2431,N_19780,N_19861);
nand UO_2432 (O_2432,N_19935,N_19855);
nor UO_2433 (O_2433,N_19881,N_19859);
xor UO_2434 (O_2434,N_19893,N_19813);
and UO_2435 (O_2435,N_19891,N_19798);
or UO_2436 (O_2436,N_19943,N_19848);
or UO_2437 (O_2437,N_19980,N_19791);
or UO_2438 (O_2438,N_19941,N_19873);
nor UO_2439 (O_2439,N_19869,N_19862);
nand UO_2440 (O_2440,N_19922,N_19978);
nand UO_2441 (O_2441,N_19770,N_19893);
and UO_2442 (O_2442,N_19946,N_19979);
or UO_2443 (O_2443,N_19969,N_19872);
nor UO_2444 (O_2444,N_19953,N_19940);
and UO_2445 (O_2445,N_19943,N_19904);
nand UO_2446 (O_2446,N_19922,N_19837);
xor UO_2447 (O_2447,N_19845,N_19775);
or UO_2448 (O_2448,N_19870,N_19970);
or UO_2449 (O_2449,N_19818,N_19867);
and UO_2450 (O_2450,N_19908,N_19796);
and UO_2451 (O_2451,N_19980,N_19951);
nand UO_2452 (O_2452,N_19883,N_19807);
nor UO_2453 (O_2453,N_19970,N_19823);
nand UO_2454 (O_2454,N_19908,N_19890);
nor UO_2455 (O_2455,N_19850,N_19956);
xor UO_2456 (O_2456,N_19815,N_19949);
nor UO_2457 (O_2457,N_19869,N_19985);
nand UO_2458 (O_2458,N_19811,N_19813);
nand UO_2459 (O_2459,N_19942,N_19944);
xnor UO_2460 (O_2460,N_19750,N_19751);
nor UO_2461 (O_2461,N_19966,N_19958);
or UO_2462 (O_2462,N_19766,N_19993);
nor UO_2463 (O_2463,N_19931,N_19772);
nand UO_2464 (O_2464,N_19882,N_19900);
nor UO_2465 (O_2465,N_19846,N_19778);
nand UO_2466 (O_2466,N_19757,N_19939);
or UO_2467 (O_2467,N_19821,N_19993);
and UO_2468 (O_2468,N_19869,N_19959);
nor UO_2469 (O_2469,N_19878,N_19848);
xor UO_2470 (O_2470,N_19911,N_19971);
or UO_2471 (O_2471,N_19916,N_19816);
nand UO_2472 (O_2472,N_19993,N_19836);
and UO_2473 (O_2473,N_19969,N_19903);
nand UO_2474 (O_2474,N_19865,N_19913);
and UO_2475 (O_2475,N_19965,N_19980);
nor UO_2476 (O_2476,N_19837,N_19806);
or UO_2477 (O_2477,N_19834,N_19935);
xnor UO_2478 (O_2478,N_19970,N_19906);
nand UO_2479 (O_2479,N_19925,N_19815);
or UO_2480 (O_2480,N_19855,N_19976);
nor UO_2481 (O_2481,N_19794,N_19883);
nand UO_2482 (O_2482,N_19798,N_19760);
xnor UO_2483 (O_2483,N_19858,N_19777);
and UO_2484 (O_2484,N_19953,N_19870);
and UO_2485 (O_2485,N_19781,N_19986);
or UO_2486 (O_2486,N_19836,N_19864);
and UO_2487 (O_2487,N_19877,N_19968);
nor UO_2488 (O_2488,N_19887,N_19778);
nand UO_2489 (O_2489,N_19884,N_19864);
or UO_2490 (O_2490,N_19967,N_19935);
or UO_2491 (O_2491,N_19769,N_19989);
xor UO_2492 (O_2492,N_19965,N_19843);
and UO_2493 (O_2493,N_19972,N_19883);
xor UO_2494 (O_2494,N_19779,N_19842);
and UO_2495 (O_2495,N_19865,N_19943);
nand UO_2496 (O_2496,N_19980,N_19909);
nand UO_2497 (O_2497,N_19928,N_19805);
nor UO_2498 (O_2498,N_19901,N_19754);
nand UO_2499 (O_2499,N_19999,N_19791);
endmodule