module basic_750_5000_1000_10_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_164,In_170);
nor U1 (N_1,In_322,In_662);
and U2 (N_2,In_236,In_114);
or U3 (N_3,In_713,In_36);
and U4 (N_4,In_188,In_231);
and U5 (N_5,In_400,In_470);
nor U6 (N_6,In_746,In_417);
xor U7 (N_7,In_7,In_660);
nand U8 (N_8,In_159,In_690);
and U9 (N_9,In_351,In_222);
nor U10 (N_10,In_520,In_545);
nand U11 (N_11,In_743,In_323);
or U12 (N_12,In_386,In_262);
or U13 (N_13,In_488,In_367);
nor U14 (N_14,In_326,In_511);
xnor U15 (N_15,In_65,In_600);
and U16 (N_16,In_183,In_287);
nand U17 (N_17,In_736,In_16);
and U18 (N_18,In_666,In_144);
and U19 (N_19,In_514,In_361);
nor U20 (N_20,In_580,In_204);
nand U21 (N_21,In_434,In_366);
or U22 (N_22,In_609,In_695);
and U23 (N_23,In_329,In_350);
nand U24 (N_24,In_415,In_633);
nor U25 (N_25,In_435,In_349);
nand U26 (N_26,In_293,In_86);
nor U27 (N_27,In_186,In_64);
and U28 (N_28,In_503,In_557);
nand U29 (N_29,In_75,In_76);
or U30 (N_30,In_558,In_411);
nor U31 (N_31,In_334,In_310);
nand U32 (N_32,In_523,In_740);
nor U33 (N_33,In_725,In_416);
nor U34 (N_34,In_10,In_431);
and U35 (N_35,In_501,In_370);
nor U36 (N_36,In_150,In_702);
and U37 (N_37,In_160,In_3);
or U38 (N_38,In_474,In_289);
nor U39 (N_39,In_549,In_252);
nor U40 (N_40,In_172,In_165);
nand U41 (N_41,In_308,In_699);
nor U42 (N_42,In_572,In_612);
and U43 (N_43,In_254,In_583);
and U44 (N_44,In_13,In_111);
or U45 (N_45,In_54,In_304);
xnor U46 (N_46,In_371,In_149);
nand U47 (N_47,In_700,In_177);
nor U48 (N_48,In_680,In_180);
or U49 (N_49,In_709,In_229);
and U50 (N_50,In_378,In_197);
nor U51 (N_51,In_429,In_279);
or U52 (N_52,In_585,In_43);
nor U53 (N_53,In_487,In_185);
and U54 (N_54,In_729,In_642);
nand U55 (N_55,In_701,In_171);
or U56 (N_56,In_352,In_283);
nor U57 (N_57,In_527,In_586);
nand U58 (N_58,In_344,In_452);
xnor U59 (N_59,In_407,In_201);
or U60 (N_60,In_207,In_607);
nand U61 (N_61,In_749,In_577);
and U62 (N_62,In_74,In_317);
nand U63 (N_63,In_747,In_90);
nand U64 (N_64,In_221,In_656);
and U65 (N_65,In_681,In_273);
and U66 (N_66,In_151,In_405);
nor U67 (N_67,In_524,In_140);
xor U68 (N_68,In_668,In_47);
and U69 (N_69,In_509,In_34);
and U70 (N_70,In_248,In_399);
and U71 (N_71,In_345,In_696);
and U72 (N_72,In_637,In_512);
and U73 (N_73,In_497,In_398);
nor U74 (N_74,In_240,In_384);
xnor U75 (N_75,In_596,In_375);
xor U76 (N_76,In_423,In_259);
or U77 (N_77,In_122,In_234);
or U78 (N_78,In_670,In_300);
or U79 (N_79,In_357,In_581);
and U80 (N_80,In_176,In_672);
or U81 (N_81,In_95,In_335);
or U82 (N_82,In_539,In_602);
nor U83 (N_83,In_529,In_8);
or U84 (N_84,In_296,In_493);
or U85 (N_85,In_80,In_288);
nor U86 (N_86,In_473,In_395);
and U87 (N_87,In_69,In_358);
nor U88 (N_88,In_320,In_167);
and U89 (N_89,In_142,In_694);
and U90 (N_90,In_362,In_475);
or U91 (N_91,In_465,In_742);
nand U92 (N_92,In_428,In_265);
nand U93 (N_93,In_129,In_98);
and U94 (N_94,In_741,In_313);
and U95 (N_95,In_44,In_675);
nor U96 (N_96,In_267,In_181);
nor U97 (N_97,In_522,In_246);
xnor U98 (N_98,In_679,In_71);
and U99 (N_99,In_591,In_360);
or U100 (N_100,In_404,In_528);
nand U101 (N_101,In_286,In_682);
and U102 (N_102,In_157,In_104);
and U103 (N_103,In_318,In_714);
or U104 (N_104,In_193,In_394);
nor U105 (N_105,In_618,In_573);
nand U106 (N_106,In_225,In_309);
and U107 (N_107,In_518,In_110);
nand U108 (N_108,In_206,In_734);
nand U109 (N_109,In_677,In_35);
or U110 (N_110,In_505,In_608);
and U111 (N_111,In_464,In_224);
or U112 (N_112,In_564,In_719);
xnor U113 (N_113,In_218,In_632);
and U114 (N_114,In_133,In_385);
nand U115 (N_115,In_712,In_55);
nand U116 (N_116,In_516,In_26);
nand U117 (N_117,In_626,In_29);
nand U118 (N_118,In_61,In_409);
nor U119 (N_119,In_315,In_565);
nor U120 (N_120,In_587,In_364);
xnor U121 (N_121,In_346,In_108);
or U122 (N_122,In_593,In_578);
or U123 (N_123,In_223,In_548);
or U124 (N_124,In_575,In_368);
and U125 (N_125,In_715,In_169);
or U126 (N_126,In_175,In_732);
nor U127 (N_127,In_247,In_698);
or U128 (N_128,In_15,In_588);
nor U129 (N_129,In_629,In_388);
nor U130 (N_130,In_673,In_93);
nand U131 (N_131,In_392,In_621);
xnor U132 (N_132,In_570,In_494);
xor U133 (N_133,In_726,In_406);
nor U134 (N_134,In_195,In_282);
or U135 (N_135,In_517,In_359);
nor U136 (N_136,In_619,In_363);
nor U137 (N_137,In_635,In_622);
and U138 (N_138,In_121,In_214);
nand U139 (N_139,In_525,In_651);
and U140 (N_140,In_555,In_678);
and U141 (N_141,In_30,In_657);
and U142 (N_142,In_544,In_650);
xnor U143 (N_143,In_492,In_597);
and U144 (N_144,In_307,In_716);
or U145 (N_145,In_532,In_63);
nand U146 (N_146,In_628,In_124);
and U147 (N_147,In_275,In_274);
nand U148 (N_148,In_336,In_128);
xnor U149 (N_149,In_264,In_245);
nand U150 (N_150,In_21,In_208);
nand U151 (N_151,In_613,In_82);
and U152 (N_152,In_354,In_448);
nor U153 (N_153,In_125,In_707);
nor U154 (N_154,In_89,In_546);
nor U155 (N_155,In_298,In_102);
or U156 (N_156,In_625,In_724);
or U157 (N_157,In_325,In_687);
nand U158 (N_158,In_58,In_620);
nor U159 (N_159,In_11,In_212);
and U160 (N_160,In_569,In_495);
xnor U161 (N_161,In_705,In_135);
nor U162 (N_162,In_105,In_439);
and U163 (N_163,In_182,In_605);
nand U164 (N_164,In_466,In_402);
and U165 (N_165,In_271,In_198);
and U166 (N_166,In_137,In_28);
or U167 (N_167,In_4,In_241);
nor U168 (N_168,In_373,In_737);
and U169 (N_169,In_50,In_674);
nor U170 (N_170,In_303,In_266);
and U171 (N_171,In_278,In_515);
and U172 (N_172,In_189,In_56);
xnor U173 (N_173,In_256,In_243);
and U174 (N_174,In_220,In_314);
nand U175 (N_175,In_215,In_382);
or U176 (N_176,In_255,In_594);
or U177 (N_177,In_441,In_531);
xnor U178 (N_178,In_79,In_192);
or U179 (N_179,In_377,In_1);
nand U180 (N_180,In_295,In_134);
nand U181 (N_181,In_476,In_645);
xnor U182 (N_182,In_285,In_51);
xnor U183 (N_183,In_263,In_92);
nor U184 (N_184,In_77,In_141);
and U185 (N_185,In_209,In_504);
nand U186 (N_186,In_59,In_299);
nor U187 (N_187,In_67,In_735);
or U188 (N_188,In_120,In_312);
nand U189 (N_189,In_233,In_490);
nor U190 (N_190,In_393,In_353);
nand U191 (N_191,In_601,In_32);
and U192 (N_192,In_199,In_553);
nand U193 (N_193,In_540,In_667);
nor U194 (N_194,In_669,In_574);
or U195 (N_195,In_106,In_109);
nor U196 (N_196,In_457,In_389);
nand U197 (N_197,In_194,In_576);
nand U198 (N_198,In_592,In_408);
xnor U199 (N_199,In_62,In_538);
nand U200 (N_200,In_455,In_306);
nand U201 (N_201,In_571,In_467);
or U202 (N_202,In_97,In_365);
xor U203 (N_203,In_284,In_444);
or U204 (N_204,In_603,In_691);
nor U205 (N_205,In_671,In_33);
nand U206 (N_206,In_658,In_268);
xor U207 (N_207,In_584,In_319);
nor U208 (N_208,In_328,In_533);
nand U209 (N_209,In_294,In_130);
or U210 (N_210,In_210,In_132);
and U211 (N_211,In_692,In_611);
nand U212 (N_212,In_462,In_23);
or U213 (N_213,In_148,In_450);
and U214 (N_214,In_610,In_723);
nand U215 (N_215,In_433,In_347);
or U216 (N_216,In_57,In_145);
or U217 (N_217,In_340,In_20);
nor U218 (N_218,In_653,In_419);
nor U219 (N_219,In_414,In_127);
and U220 (N_220,In_341,In_463);
and U221 (N_221,In_327,In_253);
and U222 (N_222,In_468,In_269);
nand U223 (N_223,In_412,In_648);
and U224 (N_224,In_708,In_281);
and U225 (N_225,In_230,In_117);
and U226 (N_226,In_506,In_242);
or U227 (N_227,In_153,In_472);
nand U228 (N_228,In_280,In_561);
or U229 (N_229,In_301,In_324);
and U230 (N_230,In_291,In_566);
nor U231 (N_231,In_277,In_445);
nand U232 (N_232,In_717,In_582);
nor U233 (N_233,In_261,In_238);
or U234 (N_234,In_630,In_482);
and U235 (N_235,In_397,In_202);
nor U236 (N_236,In_720,In_526);
or U237 (N_237,In_748,In_342);
nor U238 (N_238,In_676,In_9);
and U239 (N_239,In_537,In_541);
and U240 (N_240,In_211,In_659);
nand U241 (N_241,In_731,In_100);
nand U242 (N_242,In_119,In_706);
nor U243 (N_243,In_152,In_446);
xor U244 (N_244,In_72,In_604);
nand U245 (N_245,In_103,In_166);
nand U246 (N_246,In_547,In_646);
xnor U247 (N_247,In_639,In_118);
or U248 (N_248,In_237,In_0);
or U249 (N_249,In_391,In_543);
nor U250 (N_250,In_499,In_239);
and U251 (N_251,In_232,In_449);
or U252 (N_252,In_556,In_5);
nor U253 (N_253,In_19,In_401);
nor U254 (N_254,In_711,In_249);
or U255 (N_255,In_739,In_437);
nor U256 (N_256,In_410,In_420);
or U257 (N_257,In_250,In_728);
and U258 (N_258,In_738,In_745);
xor U259 (N_259,In_112,In_443);
or U260 (N_260,In_688,In_251);
nor U261 (N_261,In_131,In_78);
nor U262 (N_262,In_217,In_49);
nor U263 (N_263,In_614,In_46);
nand U264 (N_264,In_421,In_73);
and U265 (N_265,In_477,In_91);
nand U266 (N_266,In_478,In_685);
nor U267 (N_267,In_403,In_203);
or U268 (N_268,In_235,In_722);
and U269 (N_269,In_52,In_427);
nand U270 (N_270,In_458,In_115);
nor U271 (N_271,In_53,In_432);
nor U272 (N_272,In_302,In_6);
nand U273 (N_273,In_321,In_116);
nand U274 (N_274,In_96,In_638);
xnor U275 (N_275,In_480,In_94);
and U276 (N_276,In_507,In_213);
nand U277 (N_277,In_519,In_343);
and U278 (N_278,In_390,In_661);
or U279 (N_279,In_107,In_684);
or U280 (N_280,In_491,In_40);
and U281 (N_281,In_483,In_156);
and U282 (N_282,In_190,In_81);
or U283 (N_283,In_330,In_196);
nor U284 (N_284,In_471,In_42);
nand U285 (N_285,In_551,In_697);
nor U286 (N_286,In_615,In_184);
xor U287 (N_287,In_589,In_647);
nand U288 (N_288,In_710,In_356);
xor U289 (N_289,In_568,In_617);
or U290 (N_290,In_606,In_101);
nand U291 (N_291,In_70,In_14);
or U292 (N_292,In_616,In_559);
or U293 (N_293,In_644,In_704);
and U294 (N_294,In_590,In_454);
or U295 (N_295,In_258,In_479);
nand U296 (N_296,In_634,In_60);
nor U297 (N_297,In_461,In_599);
nand U298 (N_298,In_228,In_598);
nor U299 (N_299,In_372,In_496);
nand U300 (N_300,In_567,In_502);
and U301 (N_301,In_655,In_290);
or U302 (N_302,In_536,In_147);
or U303 (N_303,In_689,In_530);
nand U304 (N_304,In_721,In_88);
nor U305 (N_305,In_643,In_380);
or U306 (N_306,In_66,In_422);
nand U307 (N_307,In_418,In_693);
nor U308 (N_308,In_562,In_355);
nor U309 (N_309,In_376,In_649);
or U310 (N_310,In_139,In_162);
xor U311 (N_311,In_163,In_31);
and U312 (N_312,In_276,In_272);
or U313 (N_313,In_718,In_636);
and U314 (N_314,In_513,In_550);
xnor U315 (N_315,In_730,In_168);
and U316 (N_316,In_436,In_369);
or U317 (N_317,In_424,In_498);
nor U318 (N_318,In_126,In_640);
and U319 (N_319,In_12,In_703);
nand U320 (N_320,In_683,In_316);
xor U321 (N_321,In_257,In_641);
nor U322 (N_322,In_534,In_396);
nor U323 (N_323,In_453,In_311);
nor U324 (N_324,In_332,In_469);
xnor U325 (N_325,In_664,In_348);
nand U326 (N_326,In_22,In_87);
and U327 (N_327,In_339,In_48);
and U328 (N_328,In_654,In_27);
and U329 (N_329,In_146,In_459);
nand U330 (N_330,In_624,In_579);
nand U331 (N_331,In_216,In_508);
or U332 (N_332,In_425,In_297);
nand U333 (N_333,In_205,In_143);
and U334 (N_334,In_270,In_554);
or U335 (N_335,In_484,In_563);
and U336 (N_336,In_542,In_292);
nor U337 (N_337,In_623,In_627);
and U338 (N_338,In_173,In_84);
nor U339 (N_339,In_331,In_430);
nor U340 (N_340,In_38,In_174);
nand U341 (N_341,In_727,In_387);
or U342 (N_342,In_460,In_227);
nand U343 (N_343,In_83,In_521);
or U344 (N_344,In_226,In_161);
or U345 (N_345,In_631,In_456);
nor U346 (N_346,In_45,In_37);
nand U347 (N_347,In_485,In_39);
and U348 (N_348,In_244,In_744);
nor U349 (N_349,In_136,In_305);
or U350 (N_350,In_686,In_191);
and U351 (N_351,In_200,In_219);
and U352 (N_352,In_25,In_442);
or U353 (N_353,In_333,In_510);
and U354 (N_354,In_426,In_113);
nand U355 (N_355,In_383,In_338);
and U356 (N_356,In_486,In_438);
nor U357 (N_357,In_2,In_138);
xnor U358 (N_358,In_451,In_123);
or U359 (N_359,In_379,In_381);
and U360 (N_360,In_68,In_663);
and U361 (N_361,In_18,In_158);
and U362 (N_362,In_481,In_440);
nor U363 (N_363,In_552,In_535);
nand U364 (N_364,In_595,In_85);
or U365 (N_365,In_413,In_155);
nand U366 (N_366,In_489,In_17);
nor U367 (N_367,In_260,In_337);
xnor U368 (N_368,In_41,In_733);
nand U369 (N_369,In_560,In_665);
or U370 (N_370,In_24,In_154);
nor U371 (N_371,In_187,In_374);
and U372 (N_372,In_179,In_178);
xor U373 (N_373,In_99,In_652);
or U374 (N_374,In_447,In_500);
or U375 (N_375,In_606,In_79);
nand U376 (N_376,In_437,In_232);
and U377 (N_377,In_113,In_602);
or U378 (N_378,In_13,In_364);
nor U379 (N_379,In_107,In_476);
and U380 (N_380,In_320,In_172);
nor U381 (N_381,In_465,In_615);
nor U382 (N_382,In_488,In_375);
xnor U383 (N_383,In_268,In_167);
nor U384 (N_384,In_329,In_717);
xnor U385 (N_385,In_678,In_199);
and U386 (N_386,In_236,In_350);
or U387 (N_387,In_302,In_736);
or U388 (N_388,In_634,In_256);
nand U389 (N_389,In_537,In_343);
xnor U390 (N_390,In_96,In_643);
xnor U391 (N_391,In_239,In_638);
nor U392 (N_392,In_602,In_704);
and U393 (N_393,In_82,In_133);
nand U394 (N_394,In_709,In_202);
nand U395 (N_395,In_444,In_114);
and U396 (N_396,In_272,In_81);
or U397 (N_397,In_678,In_644);
xnor U398 (N_398,In_66,In_681);
and U399 (N_399,In_17,In_333);
and U400 (N_400,In_664,In_478);
nor U401 (N_401,In_328,In_420);
and U402 (N_402,In_348,In_92);
xor U403 (N_403,In_682,In_35);
xor U404 (N_404,In_682,In_458);
nor U405 (N_405,In_145,In_436);
and U406 (N_406,In_563,In_43);
nor U407 (N_407,In_100,In_617);
nand U408 (N_408,In_586,In_644);
nand U409 (N_409,In_362,In_628);
nor U410 (N_410,In_730,In_505);
nor U411 (N_411,In_719,In_605);
or U412 (N_412,In_336,In_171);
nor U413 (N_413,In_303,In_401);
nand U414 (N_414,In_473,In_162);
nor U415 (N_415,In_108,In_714);
nand U416 (N_416,In_458,In_92);
and U417 (N_417,In_254,In_536);
xnor U418 (N_418,In_543,In_714);
or U419 (N_419,In_71,In_39);
nand U420 (N_420,In_40,In_460);
nand U421 (N_421,In_274,In_633);
and U422 (N_422,In_739,In_358);
nand U423 (N_423,In_536,In_368);
nand U424 (N_424,In_124,In_460);
and U425 (N_425,In_251,In_415);
nand U426 (N_426,In_84,In_393);
or U427 (N_427,In_52,In_203);
xor U428 (N_428,In_678,In_677);
or U429 (N_429,In_44,In_557);
nor U430 (N_430,In_358,In_743);
xor U431 (N_431,In_473,In_630);
and U432 (N_432,In_217,In_80);
or U433 (N_433,In_251,In_648);
or U434 (N_434,In_441,In_289);
and U435 (N_435,In_189,In_525);
nand U436 (N_436,In_176,In_554);
nor U437 (N_437,In_368,In_237);
nor U438 (N_438,In_243,In_427);
or U439 (N_439,In_721,In_364);
and U440 (N_440,In_372,In_216);
nor U441 (N_441,In_343,In_77);
nand U442 (N_442,In_57,In_180);
or U443 (N_443,In_587,In_35);
nor U444 (N_444,In_705,In_35);
and U445 (N_445,In_372,In_529);
nor U446 (N_446,In_220,In_293);
nor U447 (N_447,In_63,In_315);
or U448 (N_448,In_729,In_411);
nand U449 (N_449,In_491,In_101);
or U450 (N_450,In_319,In_546);
nor U451 (N_451,In_517,In_117);
nor U452 (N_452,In_480,In_214);
nor U453 (N_453,In_643,In_74);
nor U454 (N_454,In_606,In_494);
xnor U455 (N_455,In_575,In_614);
xor U456 (N_456,In_624,In_659);
or U457 (N_457,In_57,In_0);
and U458 (N_458,In_618,In_530);
and U459 (N_459,In_266,In_389);
nor U460 (N_460,In_567,In_280);
nor U461 (N_461,In_510,In_195);
nand U462 (N_462,In_531,In_423);
nand U463 (N_463,In_204,In_632);
nand U464 (N_464,In_353,In_667);
and U465 (N_465,In_664,In_688);
nand U466 (N_466,In_369,In_59);
and U467 (N_467,In_723,In_330);
or U468 (N_468,In_156,In_492);
or U469 (N_469,In_545,In_285);
or U470 (N_470,In_286,In_279);
or U471 (N_471,In_436,In_270);
nand U472 (N_472,In_420,In_40);
and U473 (N_473,In_483,In_79);
and U474 (N_474,In_315,In_278);
and U475 (N_475,In_4,In_568);
nor U476 (N_476,In_418,In_103);
nor U477 (N_477,In_51,In_625);
and U478 (N_478,In_390,In_405);
nand U479 (N_479,In_269,In_604);
and U480 (N_480,In_348,In_4);
or U481 (N_481,In_680,In_540);
xnor U482 (N_482,In_3,In_358);
or U483 (N_483,In_366,In_340);
nor U484 (N_484,In_345,In_88);
nor U485 (N_485,In_718,In_694);
nand U486 (N_486,In_283,In_281);
nor U487 (N_487,In_11,In_720);
and U488 (N_488,In_584,In_221);
and U489 (N_489,In_86,In_204);
and U490 (N_490,In_575,In_400);
nand U491 (N_491,In_303,In_742);
or U492 (N_492,In_164,In_14);
or U493 (N_493,In_685,In_407);
and U494 (N_494,In_694,In_684);
nor U495 (N_495,In_176,In_570);
and U496 (N_496,In_679,In_709);
nand U497 (N_497,In_95,In_477);
or U498 (N_498,In_142,In_35);
nor U499 (N_499,In_181,In_623);
and U500 (N_500,N_423,N_55);
or U501 (N_501,N_18,N_344);
and U502 (N_502,N_8,N_380);
xnor U503 (N_503,N_425,N_435);
nand U504 (N_504,N_292,N_485);
or U505 (N_505,N_258,N_346);
nand U506 (N_506,N_280,N_16);
nor U507 (N_507,N_491,N_327);
nand U508 (N_508,N_216,N_359);
and U509 (N_509,N_125,N_471);
and U510 (N_510,N_391,N_294);
xnor U511 (N_511,N_308,N_137);
nor U512 (N_512,N_28,N_301);
nand U513 (N_513,N_191,N_393);
or U514 (N_514,N_37,N_401);
and U515 (N_515,N_404,N_204);
xor U516 (N_516,N_326,N_94);
xnor U517 (N_517,N_453,N_56);
nand U518 (N_518,N_402,N_383);
nand U519 (N_519,N_26,N_236);
xor U520 (N_520,N_349,N_493);
nand U521 (N_521,N_31,N_469);
and U522 (N_522,N_376,N_63);
nand U523 (N_523,N_46,N_73);
nand U524 (N_524,N_40,N_281);
nand U525 (N_525,N_190,N_377);
xor U526 (N_526,N_405,N_218);
or U527 (N_527,N_316,N_84);
xor U528 (N_528,N_355,N_450);
nand U529 (N_529,N_411,N_487);
or U530 (N_530,N_59,N_368);
or U531 (N_531,N_282,N_345);
xnor U532 (N_532,N_240,N_388);
nor U533 (N_533,N_34,N_177);
nand U534 (N_534,N_472,N_168);
nor U535 (N_535,N_263,N_203);
nor U536 (N_536,N_489,N_441);
nor U537 (N_537,N_74,N_224);
nand U538 (N_538,N_429,N_181);
xor U539 (N_539,N_211,N_473);
or U540 (N_540,N_217,N_398);
xnor U541 (N_541,N_445,N_322);
and U542 (N_542,N_71,N_418);
xor U543 (N_543,N_185,N_342);
nand U544 (N_544,N_307,N_65);
and U545 (N_545,N_114,N_156);
xnor U546 (N_546,N_428,N_335);
and U547 (N_547,N_357,N_225);
or U548 (N_548,N_486,N_439);
and U549 (N_549,N_314,N_188);
nand U550 (N_550,N_146,N_27);
and U551 (N_551,N_331,N_262);
or U552 (N_552,N_430,N_350);
and U553 (N_553,N_436,N_298);
nand U554 (N_554,N_247,N_70);
and U555 (N_555,N_139,N_4);
and U556 (N_556,N_271,N_272);
nor U557 (N_557,N_78,N_482);
or U558 (N_558,N_348,N_295);
or U559 (N_559,N_132,N_309);
nor U560 (N_560,N_245,N_52);
and U561 (N_561,N_235,N_264);
nor U562 (N_562,N_417,N_1);
and U563 (N_563,N_149,N_494);
or U564 (N_564,N_303,N_497);
xor U565 (N_565,N_250,N_67);
xnor U566 (N_566,N_124,N_186);
and U567 (N_567,N_289,N_174);
nand U568 (N_568,N_25,N_150);
nand U569 (N_569,N_131,N_286);
nor U570 (N_570,N_479,N_363);
and U571 (N_571,N_440,N_385);
and U572 (N_572,N_318,N_9);
nand U573 (N_573,N_33,N_134);
nand U574 (N_574,N_437,N_302);
nor U575 (N_575,N_47,N_374);
and U576 (N_576,N_154,N_324);
nor U577 (N_577,N_347,N_477);
or U578 (N_578,N_396,N_300);
nor U579 (N_579,N_136,N_45);
and U580 (N_580,N_296,N_449);
and U581 (N_581,N_317,N_241);
xnor U582 (N_582,N_305,N_413);
and U583 (N_583,N_448,N_118);
and U584 (N_584,N_228,N_170);
and U585 (N_585,N_351,N_36);
nor U586 (N_586,N_115,N_457);
nand U587 (N_587,N_279,N_192);
nor U588 (N_588,N_127,N_284);
nand U589 (N_589,N_256,N_283);
and U590 (N_590,N_287,N_189);
and U591 (N_591,N_242,N_173);
nor U592 (N_592,N_277,N_29);
nor U593 (N_593,N_179,N_382);
nor U594 (N_594,N_323,N_220);
or U595 (N_595,N_111,N_468);
xnor U596 (N_596,N_432,N_315);
nand U597 (N_597,N_231,N_395);
and U598 (N_598,N_381,N_13);
or U599 (N_599,N_2,N_7);
nor U600 (N_600,N_147,N_336);
or U601 (N_601,N_144,N_109);
or U602 (N_602,N_354,N_130);
and U603 (N_603,N_332,N_321);
and U604 (N_604,N_403,N_379);
nor U605 (N_605,N_495,N_265);
or U606 (N_606,N_199,N_213);
xor U607 (N_607,N_145,N_400);
xnor U608 (N_608,N_105,N_461);
nand U609 (N_609,N_244,N_416);
and U610 (N_610,N_194,N_122);
and U611 (N_611,N_397,N_82);
or U612 (N_612,N_483,N_157);
and U613 (N_613,N_51,N_169);
nand U614 (N_614,N_103,N_64);
nor U615 (N_615,N_361,N_434);
nor U616 (N_616,N_358,N_340);
nand U617 (N_617,N_455,N_15);
nand U618 (N_618,N_375,N_338);
and U619 (N_619,N_66,N_30);
or U620 (N_620,N_221,N_88);
and U621 (N_621,N_227,N_79);
nor U622 (N_622,N_492,N_95);
xnor U623 (N_623,N_270,N_38);
nand U624 (N_624,N_3,N_238);
or U625 (N_625,N_275,N_72);
xnor U626 (N_626,N_460,N_198);
and U627 (N_627,N_389,N_116);
or U628 (N_628,N_446,N_32);
and U629 (N_629,N_129,N_50);
or U630 (N_630,N_373,N_113);
nor U631 (N_631,N_320,N_499);
nor U632 (N_632,N_454,N_6);
nand U633 (N_633,N_133,N_187);
nor U634 (N_634,N_343,N_80);
nand U635 (N_635,N_176,N_442);
nand U636 (N_636,N_152,N_269);
nand U637 (N_637,N_77,N_310);
or U638 (N_638,N_219,N_490);
nand U639 (N_639,N_274,N_232);
xor U640 (N_640,N_162,N_339);
and U641 (N_641,N_107,N_180);
nand U642 (N_642,N_370,N_41);
or U643 (N_643,N_178,N_172);
nand U644 (N_644,N_255,N_311);
or U645 (N_645,N_252,N_478);
xnor U646 (N_646,N_0,N_160);
nand U647 (N_647,N_313,N_239);
nor U648 (N_648,N_365,N_366);
and U649 (N_649,N_42,N_447);
nand U650 (N_650,N_43,N_22);
nor U651 (N_651,N_337,N_424);
xnor U652 (N_652,N_452,N_49);
xnor U653 (N_653,N_155,N_249);
and U654 (N_654,N_202,N_387);
nand U655 (N_655,N_85,N_293);
and U656 (N_656,N_167,N_119);
or U657 (N_657,N_319,N_267);
xnor U658 (N_658,N_62,N_128);
nor U659 (N_659,N_98,N_438);
xnor U660 (N_660,N_456,N_421);
or U661 (N_661,N_422,N_215);
and U662 (N_662,N_356,N_17);
or U663 (N_663,N_341,N_234);
nand U664 (N_664,N_390,N_212);
nand U665 (N_665,N_81,N_183);
or U666 (N_666,N_104,N_54);
or U667 (N_667,N_407,N_158);
nand U668 (N_668,N_386,N_151);
nor U669 (N_669,N_19,N_58);
or U670 (N_670,N_75,N_384);
nor U671 (N_671,N_117,N_196);
or U672 (N_672,N_44,N_106);
nor U673 (N_673,N_325,N_10);
or U674 (N_674,N_53,N_299);
nor U675 (N_675,N_312,N_378);
or U676 (N_676,N_12,N_142);
or U677 (N_677,N_304,N_463);
nor U678 (N_678,N_171,N_352);
xor U679 (N_679,N_99,N_92);
nand U680 (N_680,N_222,N_254);
nand U681 (N_681,N_251,N_223);
nand U682 (N_682,N_433,N_409);
and U683 (N_683,N_306,N_166);
and U684 (N_684,N_243,N_89);
and U685 (N_685,N_48,N_464);
or U686 (N_686,N_290,N_291);
nor U687 (N_687,N_498,N_60);
nand U688 (N_688,N_467,N_431);
nor U689 (N_689,N_21,N_259);
nand U690 (N_690,N_392,N_209);
and U691 (N_691,N_35,N_394);
xor U692 (N_692,N_253,N_5);
or U693 (N_693,N_362,N_276);
nor U694 (N_694,N_237,N_419);
nor U695 (N_695,N_484,N_288);
xnor U696 (N_696,N_474,N_148);
nand U697 (N_697,N_201,N_123);
or U698 (N_698,N_61,N_260);
nor U699 (N_699,N_11,N_112);
nor U700 (N_700,N_462,N_120);
nor U701 (N_701,N_90,N_143);
and U702 (N_702,N_161,N_475);
nand U703 (N_703,N_412,N_257);
or U704 (N_704,N_76,N_86);
nor U705 (N_705,N_233,N_268);
or U706 (N_706,N_23,N_426);
nand U707 (N_707,N_207,N_83);
nand U708 (N_708,N_476,N_246);
nor U709 (N_709,N_87,N_206);
nand U710 (N_710,N_229,N_138);
or U711 (N_711,N_427,N_184);
xnor U712 (N_712,N_488,N_163);
or U713 (N_713,N_214,N_333);
and U714 (N_714,N_415,N_153);
and U715 (N_715,N_208,N_459);
nor U716 (N_716,N_101,N_197);
and U717 (N_717,N_367,N_226);
nor U718 (N_718,N_372,N_328);
nand U719 (N_719,N_285,N_443);
or U720 (N_720,N_91,N_39);
nor U721 (N_721,N_68,N_480);
xnor U722 (N_722,N_110,N_266);
nor U723 (N_723,N_414,N_193);
xor U724 (N_724,N_248,N_444);
or U725 (N_725,N_273,N_108);
or U726 (N_726,N_466,N_399);
nand U727 (N_727,N_165,N_278);
nand U728 (N_728,N_126,N_195);
or U729 (N_729,N_353,N_102);
or U730 (N_730,N_205,N_408);
and U731 (N_731,N_330,N_135);
and U732 (N_732,N_369,N_141);
nor U733 (N_733,N_334,N_420);
nand U734 (N_734,N_121,N_261);
nand U735 (N_735,N_200,N_140);
or U736 (N_736,N_451,N_97);
nor U737 (N_737,N_360,N_297);
nand U738 (N_738,N_496,N_406);
nand U739 (N_739,N_24,N_329);
nor U740 (N_740,N_57,N_96);
and U741 (N_741,N_159,N_182);
xnor U742 (N_742,N_410,N_69);
and U743 (N_743,N_210,N_175);
and U744 (N_744,N_470,N_481);
nand U745 (N_745,N_458,N_465);
or U746 (N_746,N_371,N_364);
or U747 (N_747,N_20,N_230);
or U748 (N_748,N_93,N_164);
and U749 (N_749,N_14,N_100);
or U750 (N_750,N_484,N_63);
nor U751 (N_751,N_291,N_408);
and U752 (N_752,N_407,N_316);
nand U753 (N_753,N_233,N_413);
nand U754 (N_754,N_45,N_177);
and U755 (N_755,N_205,N_442);
or U756 (N_756,N_118,N_170);
nand U757 (N_757,N_145,N_299);
or U758 (N_758,N_124,N_85);
or U759 (N_759,N_129,N_393);
nor U760 (N_760,N_464,N_209);
nand U761 (N_761,N_200,N_292);
xor U762 (N_762,N_461,N_413);
and U763 (N_763,N_324,N_484);
or U764 (N_764,N_85,N_133);
and U765 (N_765,N_319,N_36);
or U766 (N_766,N_161,N_92);
and U767 (N_767,N_148,N_297);
nand U768 (N_768,N_380,N_44);
and U769 (N_769,N_75,N_388);
nand U770 (N_770,N_275,N_492);
nor U771 (N_771,N_173,N_164);
nand U772 (N_772,N_332,N_245);
nor U773 (N_773,N_365,N_319);
nand U774 (N_774,N_138,N_317);
or U775 (N_775,N_414,N_485);
nor U776 (N_776,N_424,N_131);
and U777 (N_777,N_369,N_248);
nor U778 (N_778,N_148,N_28);
nand U779 (N_779,N_78,N_55);
and U780 (N_780,N_240,N_184);
and U781 (N_781,N_48,N_222);
nand U782 (N_782,N_447,N_406);
nor U783 (N_783,N_370,N_454);
or U784 (N_784,N_16,N_69);
and U785 (N_785,N_299,N_232);
nand U786 (N_786,N_183,N_42);
and U787 (N_787,N_83,N_466);
nor U788 (N_788,N_87,N_319);
xnor U789 (N_789,N_175,N_96);
or U790 (N_790,N_164,N_355);
nor U791 (N_791,N_305,N_442);
nand U792 (N_792,N_42,N_109);
and U793 (N_793,N_168,N_45);
xnor U794 (N_794,N_425,N_298);
and U795 (N_795,N_155,N_213);
or U796 (N_796,N_496,N_368);
nor U797 (N_797,N_40,N_139);
nand U798 (N_798,N_335,N_363);
nand U799 (N_799,N_284,N_347);
nor U800 (N_800,N_106,N_486);
nor U801 (N_801,N_327,N_435);
nor U802 (N_802,N_499,N_305);
nand U803 (N_803,N_61,N_83);
or U804 (N_804,N_233,N_84);
nand U805 (N_805,N_434,N_36);
nand U806 (N_806,N_304,N_275);
nor U807 (N_807,N_19,N_470);
xor U808 (N_808,N_407,N_499);
nor U809 (N_809,N_168,N_288);
nor U810 (N_810,N_151,N_81);
or U811 (N_811,N_181,N_470);
and U812 (N_812,N_127,N_171);
and U813 (N_813,N_377,N_463);
xor U814 (N_814,N_328,N_388);
nand U815 (N_815,N_47,N_144);
xor U816 (N_816,N_217,N_215);
and U817 (N_817,N_468,N_400);
or U818 (N_818,N_72,N_245);
nor U819 (N_819,N_178,N_468);
xnor U820 (N_820,N_483,N_55);
nand U821 (N_821,N_22,N_38);
nor U822 (N_822,N_56,N_33);
and U823 (N_823,N_463,N_383);
xnor U824 (N_824,N_56,N_70);
nor U825 (N_825,N_37,N_133);
or U826 (N_826,N_308,N_31);
nor U827 (N_827,N_67,N_77);
nor U828 (N_828,N_265,N_161);
nand U829 (N_829,N_421,N_193);
nor U830 (N_830,N_321,N_77);
and U831 (N_831,N_427,N_108);
or U832 (N_832,N_172,N_198);
or U833 (N_833,N_457,N_396);
nor U834 (N_834,N_403,N_457);
and U835 (N_835,N_78,N_437);
nor U836 (N_836,N_206,N_61);
nor U837 (N_837,N_106,N_192);
nand U838 (N_838,N_259,N_453);
nand U839 (N_839,N_454,N_426);
or U840 (N_840,N_395,N_264);
xor U841 (N_841,N_41,N_75);
xnor U842 (N_842,N_426,N_340);
nor U843 (N_843,N_163,N_50);
nor U844 (N_844,N_477,N_251);
nand U845 (N_845,N_138,N_432);
nor U846 (N_846,N_175,N_335);
or U847 (N_847,N_55,N_76);
xnor U848 (N_848,N_266,N_250);
or U849 (N_849,N_185,N_340);
nor U850 (N_850,N_461,N_144);
or U851 (N_851,N_129,N_69);
and U852 (N_852,N_333,N_373);
and U853 (N_853,N_218,N_313);
or U854 (N_854,N_325,N_394);
and U855 (N_855,N_155,N_368);
nor U856 (N_856,N_171,N_368);
or U857 (N_857,N_351,N_468);
and U858 (N_858,N_152,N_331);
nand U859 (N_859,N_181,N_312);
or U860 (N_860,N_79,N_300);
and U861 (N_861,N_239,N_226);
nor U862 (N_862,N_140,N_137);
or U863 (N_863,N_225,N_335);
or U864 (N_864,N_3,N_255);
nand U865 (N_865,N_414,N_49);
nand U866 (N_866,N_147,N_20);
nand U867 (N_867,N_72,N_336);
xnor U868 (N_868,N_315,N_373);
or U869 (N_869,N_171,N_273);
nor U870 (N_870,N_483,N_222);
nand U871 (N_871,N_266,N_189);
and U872 (N_872,N_432,N_306);
or U873 (N_873,N_4,N_460);
and U874 (N_874,N_433,N_302);
or U875 (N_875,N_292,N_14);
xnor U876 (N_876,N_168,N_1);
nand U877 (N_877,N_217,N_4);
xnor U878 (N_878,N_323,N_474);
and U879 (N_879,N_402,N_145);
or U880 (N_880,N_265,N_388);
or U881 (N_881,N_497,N_124);
nand U882 (N_882,N_355,N_209);
or U883 (N_883,N_498,N_25);
or U884 (N_884,N_380,N_93);
nand U885 (N_885,N_6,N_246);
nand U886 (N_886,N_360,N_38);
or U887 (N_887,N_245,N_266);
nand U888 (N_888,N_198,N_332);
nor U889 (N_889,N_70,N_168);
nor U890 (N_890,N_2,N_106);
and U891 (N_891,N_282,N_38);
nand U892 (N_892,N_289,N_339);
nor U893 (N_893,N_367,N_75);
or U894 (N_894,N_166,N_325);
nor U895 (N_895,N_381,N_185);
nand U896 (N_896,N_122,N_457);
nor U897 (N_897,N_496,N_300);
nand U898 (N_898,N_174,N_414);
or U899 (N_899,N_50,N_42);
xor U900 (N_900,N_429,N_269);
nand U901 (N_901,N_103,N_171);
nor U902 (N_902,N_271,N_146);
nand U903 (N_903,N_314,N_328);
nor U904 (N_904,N_463,N_494);
and U905 (N_905,N_381,N_453);
and U906 (N_906,N_124,N_245);
nand U907 (N_907,N_164,N_407);
xnor U908 (N_908,N_294,N_83);
nor U909 (N_909,N_245,N_434);
and U910 (N_910,N_107,N_30);
nand U911 (N_911,N_340,N_222);
nor U912 (N_912,N_499,N_461);
xor U913 (N_913,N_56,N_25);
and U914 (N_914,N_319,N_195);
and U915 (N_915,N_498,N_258);
xor U916 (N_916,N_53,N_250);
nand U917 (N_917,N_213,N_63);
nand U918 (N_918,N_404,N_2);
or U919 (N_919,N_84,N_374);
nand U920 (N_920,N_46,N_215);
nor U921 (N_921,N_416,N_279);
or U922 (N_922,N_469,N_411);
or U923 (N_923,N_267,N_247);
or U924 (N_924,N_259,N_34);
xnor U925 (N_925,N_488,N_63);
or U926 (N_926,N_472,N_336);
nand U927 (N_927,N_74,N_79);
nor U928 (N_928,N_231,N_287);
or U929 (N_929,N_314,N_127);
nor U930 (N_930,N_151,N_315);
xor U931 (N_931,N_442,N_297);
nand U932 (N_932,N_337,N_390);
nor U933 (N_933,N_492,N_325);
nor U934 (N_934,N_416,N_326);
and U935 (N_935,N_230,N_163);
nand U936 (N_936,N_29,N_344);
and U937 (N_937,N_171,N_210);
nand U938 (N_938,N_21,N_468);
nor U939 (N_939,N_144,N_176);
or U940 (N_940,N_300,N_428);
nor U941 (N_941,N_338,N_464);
nor U942 (N_942,N_294,N_157);
xor U943 (N_943,N_122,N_186);
and U944 (N_944,N_140,N_85);
xor U945 (N_945,N_448,N_119);
and U946 (N_946,N_489,N_238);
xor U947 (N_947,N_142,N_277);
nand U948 (N_948,N_421,N_199);
nor U949 (N_949,N_285,N_164);
nand U950 (N_950,N_242,N_467);
nor U951 (N_951,N_347,N_183);
nor U952 (N_952,N_115,N_279);
or U953 (N_953,N_430,N_464);
nand U954 (N_954,N_271,N_483);
nor U955 (N_955,N_361,N_100);
nand U956 (N_956,N_227,N_420);
nand U957 (N_957,N_477,N_205);
and U958 (N_958,N_425,N_323);
nand U959 (N_959,N_359,N_260);
or U960 (N_960,N_184,N_387);
nor U961 (N_961,N_373,N_94);
nand U962 (N_962,N_224,N_424);
nand U963 (N_963,N_476,N_60);
or U964 (N_964,N_280,N_361);
or U965 (N_965,N_233,N_290);
nor U966 (N_966,N_224,N_219);
nand U967 (N_967,N_386,N_301);
nand U968 (N_968,N_422,N_94);
or U969 (N_969,N_296,N_476);
xor U970 (N_970,N_478,N_480);
or U971 (N_971,N_246,N_350);
and U972 (N_972,N_378,N_494);
nor U973 (N_973,N_100,N_8);
nor U974 (N_974,N_195,N_68);
nor U975 (N_975,N_4,N_43);
nor U976 (N_976,N_338,N_52);
or U977 (N_977,N_232,N_204);
or U978 (N_978,N_323,N_308);
and U979 (N_979,N_383,N_175);
xnor U980 (N_980,N_308,N_213);
or U981 (N_981,N_385,N_109);
nor U982 (N_982,N_481,N_350);
or U983 (N_983,N_363,N_226);
xnor U984 (N_984,N_332,N_362);
and U985 (N_985,N_95,N_355);
nand U986 (N_986,N_483,N_434);
nor U987 (N_987,N_200,N_382);
xnor U988 (N_988,N_160,N_415);
nand U989 (N_989,N_282,N_247);
nand U990 (N_990,N_439,N_79);
or U991 (N_991,N_128,N_325);
nor U992 (N_992,N_449,N_468);
and U993 (N_993,N_349,N_377);
or U994 (N_994,N_160,N_20);
nand U995 (N_995,N_281,N_35);
and U996 (N_996,N_469,N_57);
and U997 (N_997,N_413,N_373);
or U998 (N_998,N_222,N_62);
nand U999 (N_999,N_2,N_147);
nor U1000 (N_1000,N_965,N_919);
nand U1001 (N_1001,N_916,N_608);
nor U1002 (N_1002,N_977,N_819);
and U1003 (N_1003,N_893,N_783);
nor U1004 (N_1004,N_818,N_800);
nor U1005 (N_1005,N_744,N_983);
xnor U1006 (N_1006,N_659,N_935);
nor U1007 (N_1007,N_778,N_793);
nand U1008 (N_1008,N_904,N_578);
xor U1009 (N_1009,N_998,N_545);
and U1010 (N_1010,N_816,N_680);
nor U1011 (N_1011,N_588,N_634);
xor U1012 (N_1012,N_502,N_698);
nor U1013 (N_1013,N_687,N_939);
nand U1014 (N_1014,N_693,N_604);
nand U1015 (N_1015,N_932,N_947);
xnor U1016 (N_1016,N_573,N_596);
xnor U1017 (N_1017,N_673,N_937);
and U1018 (N_1018,N_838,N_665);
and U1019 (N_1019,N_973,N_789);
xor U1020 (N_1020,N_576,N_841);
nand U1021 (N_1021,N_592,N_533);
and U1022 (N_1022,N_513,N_548);
nand U1023 (N_1023,N_745,N_913);
xnor U1024 (N_1024,N_633,N_637);
and U1025 (N_1025,N_942,N_833);
xnor U1026 (N_1026,N_832,N_717);
nor U1027 (N_1027,N_929,N_541);
nand U1028 (N_1028,N_820,N_674);
and U1029 (N_1029,N_572,N_992);
nand U1030 (N_1030,N_714,N_503);
and U1031 (N_1031,N_658,N_955);
xnor U1032 (N_1032,N_875,N_722);
and U1033 (N_1033,N_975,N_842);
or U1034 (N_1034,N_761,N_809);
nand U1035 (N_1035,N_969,N_663);
nand U1036 (N_1036,N_974,N_537);
xnor U1037 (N_1037,N_524,N_516);
nor U1038 (N_1038,N_856,N_890);
nor U1039 (N_1039,N_515,N_870);
nand U1040 (N_1040,N_643,N_544);
and U1041 (N_1041,N_551,N_797);
or U1042 (N_1042,N_688,N_689);
nand U1043 (N_1043,N_764,N_917);
and U1044 (N_1044,N_521,N_854);
nand U1045 (N_1045,N_962,N_641);
nand U1046 (N_1046,N_991,N_821);
nor U1047 (N_1047,N_682,N_827);
and U1048 (N_1048,N_812,N_859);
nand U1049 (N_1049,N_964,N_584);
and U1050 (N_1050,N_702,N_766);
and U1051 (N_1051,N_653,N_520);
nand U1052 (N_1052,N_956,N_599);
or U1053 (N_1053,N_712,N_569);
nand U1054 (N_1054,N_678,N_774);
nor U1055 (N_1055,N_945,N_750);
or U1056 (N_1056,N_899,N_640);
nand U1057 (N_1057,N_928,N_598);
nor U1058 (N_1058,N_925,N_754);
or U1059 (N_1059,N_726,N_924);
and U1060 (N_1060,N_857,N_853);
or U1061 (N_1061,N_861,N_669);
and U1062 (N_1062,N_755,N_705);
or U1063 (N_1063,N_996,N_926);
nor U1064 (N_1064,N_664,N_948);
nor U1065 (N_1065,N_655,N_751);
or U1066 (N_1066,N_614,N_791);
nand U1067 (N_1067,N_798,N_512);
nand U1068 (N_1068,N_867,N_619);
nand U1069 (N_1069,N_910,N_999);
or U1070 (N_1070,N_523,N_970);
nor U1071 (N_1071,N_632,N_574);
xor U1072 (N_1072,N_748,N_518);
nor U1073 (N_1073,N_933,N_708);
nor U1074 (N_1074,N_994,N_906);
nor U1075 (N_1075,N_963,N_782);
nand U1076 (N_1076,N_718,N_550);
or U1077 (N_1077,N_629,N_630);
and U1078 (N_1078,N_880,N_651);
nand U1079 (N_1079,N_891,N_567);
nor U1080 (N_1080,N_773,N_577);
or U1081 (N_1081,N_734,N_605);
nor U1082 (N_1082,N_677,N_845);
nand U1083 (N_1083,N_603,N_834);
nor U1084 (N_1084,N_786,N_531);
or U1085 (N_1085,N_601,N_609);
nor U1086 (N_1086,N_727,N_644);
nor U1087 (N_1087,N_894,N_912);
and U1088 (N_1088,N_730,N_522);
and U1089 (N_1089,N_990,N_892);
or U1090 (N_1090,N_679,N_954);
or U1091 (N_1091,N_539,N_606);
nor U1092 (N_1092,N_989,N_529);
xnor U1093 (N_1093,N_792,N_984);
nor U1094 (N_1094,N_799,N_938);
or U1095 (N_1095,N_525,N_556);
nor U1096 (N_1096,N_626,N_780);
and U1097 (N_1097,N_728,N_535);
and U1098 (N_1098,N_873,N_957);
and U1099 (N_1099,N_628,N_565);
nand U1100 (N_1100,N_887,N_918);
nand U1101 (N_1101,N_920,N_570);
nor U1102 (N_1102,N_966,N_874);
or U1103 (N_1103,N_901,N_807);
nor U1104 (N_1104,N_746,N_769);
or U1105 (N_1105,N_639,N_528);
and U1106 (N_1106,N_747,N_757);
and U1107 (N_1107,N_784,N_546);
nand U1108 (N_1108,N_506,N_622);
nand U1109 (N_1109,N_949,N_505);
xor U1110 (N_1110,N_787,N_772);
or U1111 (N_1111,N_790,N_828);
and U1112 (N_1112,N_504,N_931);
xnor U1113 (N_1113,N_770,N_645);
xnor U1114 (N_1114,N_553,N_972);
nor U1115 (N_1115,N_624,N_552);
nor U1116 (N_1116,N_858,N_872);
nand U1117 (N_1117,N_701,N_566);
and U1118 (N_1118,N_796,N_612);
nand U1119 (N_1119,N_547,N_840);
or U1120 (N_1120,N_923,N_709);
nor U1121 (N_1121,N_871,N_716);
xor U1122 (N_1122,N_738,N_971);
and U1123 (N_1123,N_638,N_952);
or U1124 (N_1124,N_559,N_767);
nand U1125 (N_1125,N_811,N_666);
and U1126 (N_1126,N_720,N_826);
or U1127 (N_1127,N_921,N_978);
nand U1128 (N_1128,N_562,N_731);
and U1129 (N_1129,N_776,N_788);
nand U1130 (N_1130,N_876,N_940);
and U1131 (N_1131,N_986,N_697);
xor U1132 (N_1132,N_930,N_543);
and U1133 (N_1133,N_713,N_737);
or U1134 (N_1134,N_768,N_909);
xor U1135 (N_1135,N_941,N_946);
nand U1136 (N_1136,N_879,N_944);
nand U1137 (N_1137,N_882,N_808);
or U1138 (N_1138,N_775,N_943);
nor U1139 (N_1139,N_736,N_813);
nand U1140 (N_1140,N_690,N_881);
and U1141 (N_1141,N_648,N_863);
or U1142 (N_1142,N_895,N_685);
nand U1143 (N_1143,N_560,N_777);
and U1144 (N_1144,N_922,N_691);
nand U1145 (N_1145,N_968,N_883);
nor U1146 (N_1146,N_810,N_517);
and U1147 (N_1147,N_710,N_707);
xor U1148 (N_1148,N_900,N_934);
and U1149 (N_1149,N_620,N_993);
nor U1150 (N_1150,N_927,N_670);
or U1151 (N_1151,N_740,N_607);
nand U1152 (N_1152,N_958,N_613);
nand U1153 (N_1153,N_616,N_844);
nor U1154 (N_1154,N_846,N_959);
nor U1155 (N_1155,N_950,N_597);
and U1156 (N_1156,N_721,N_802);
xor U1157 (N_1157,N_835,N_866);
and U1158 (N_1158,N_815,N_695);
nor U1159 (N_1159,N_555,N_985);
nor U1160 (N_1160,N_650,N_580);
nand U1161 (N_1161,N_635,N_885);
or U1162 (N_1162,N_563,N_785);
and U1163 (N_1163,N_649,N_660);
nor U1164 (N_1164,N_829,N_571);
and U1165 (N_1165,N_536,N_724);
nor U1166 (N_1166,N_739,N_500);
or U1167 (N_1167,N_590,N_549);
xnor U1168 (N_1168,N_997,N_527);
nor U1169 (N_1169,N_915,N_749);
nor U1170 (N_1170,N_814,N_756);
or U1171 (N_1171,N_869,N_804);
or U1172 (N_1172,N_723,N_836);
and U1173 (N_1173,N_557,N_847);
nand U1174 (N_1174,N_631,N_532);
or U1175 (N_1175,N_591,N_843);
nor U1176 (N_1176,N_661,N_684);
or U1177 (N_1177,N_611,N_903);
nor U1178 (N_1178,N_558,N_621);
xnor U1179 (N_1179,N_850,N_568);
or U1180 (N_1180,N_686,N_675);
and U1181 (N_1181,N_610,N_822);
nand U1182 (N_1182,N_507,N_907);
and U1183 (N_1183,N_823,N_575);
and U1184 (N_1184,N_715,N_762);
xnor U1185 (N_1185,N_781,N_884);
nor U1186 (N_1186,N_540,N_526);
nor U1187 (N_1187,N_699,N_760);
nor U1188 (N_1188,N_729,N_554);
nor U1189 (N_1189,N_636,N_831);
or U1190 (N_1190,N_752,N_511);
or U1191 (N_1191,N_771,N_877);
nor U1192 (N_1192,N_742,N_676);
or U1193 (N_1193,N_642,N_741);
xnor U1194 (N_1194,N_806,N_896);
or U1195 (N_1195,N_595,N_681);
or U1196 (N_1196,N_719,N_706);
xnor U1197 (N_1197,N_646,N_898);
and U1198 (N_1198,N_615,N_561);
and U1199 (N_1199,N_743,N_980);
or U1200 (N_1200,N_839,N_855);
or U1201 (N_1201,N_667,N_837);
nand U1202 (N_1202,N_662,N_967);
nor U1203 (N_1203,N_542,N_509);
and U1204 (N_1204,N_888,N_514);
nor U1205 (N_1205,N_886,N_510);
nand U1206 (N_1206,N_586,N_794);
or U1207 (N_1207,N_803,N_725);
or U1208 (N_1208,N_585,N_961);
nor U1209 (N_1209,N_936,N_825);
nand U1210 (N_1210,N_652,N_902);
nor U1211 (N_1211,N_765,N_617);
or U1212 (N_1212,N_897,N_795);
nor U1213 (N_1213,N_703,N_735);
and U1214 (N_1214,N_733,N_779);
and U1215 (N_1215,N_647,N_700);
nand U1216 (N_1216,N_995,N_911);
or U1217 (N_1217,N_711,N_732);
nand U1218 (N_1218,N_696,N_704);
nor U1219 (N_1219,N_564,N_582);
nor U1220 (N_1220,N_805,N_979);
and U1221 (N_1221,N_865,N_981);
and U1222 (N_1222,N_530,N_683);
and U1223 (N_1223,N_976,N_951);
xor U1224 (N_1224,N_623,N_692);
and U1225 (N_1225,N_587,N_908);
nand U1226 (N_1226,N_593,N_538);
or U1227 (N_1227,N_657,N_753);
xor U1228 (N_1228,N_914,N_519);
or U1229 (N_1229,N_579,N_982);
nor U1230 (N_1230,N_589,N_656);
and U1231 (N_1231,N_824,N_878);
and U1232 (N_1232,N_988,N_583);
and U1233 (N_1233,N_868,N_758);
nor U1234 (N_1234,N_671,N_594);
nor U1235 (N_1235,N_501,N_694);
xor U1236 (N_1236,N_860,N_801);
and U1237 (N_1237,N_848,N_600);
and U1238 (N_1238,N_960,N_618);
nand U1239 (N_1239,N_864,N_602);
nand U1240 (N_1240,N_889,N_852);
nand U1241 (N_1241,N_849,N_830);
xor U1242 (N_1242,N_668,N_654);
or U1243 (N_1243,N_672,N_862);
nand U1244 (N_1244,N_987,N_627);
nand U1245 (N_1245,N_817,N_851);
or U1246 (N_1246,N_508,N_625);
nor U1247 (N_1247,N_763,N_581);
and U1248 (N_1248,N_534,N_759);
xnor U1249 (N_1249,N_953,N_905);
nor U1250 (N_1250,N_881,N_910);
nor U1251 (N_1251,N_897,N_891);
nand U1252 (N_1252,N_513,N_657);
or U1253 (N_1253,N_509,N_752);
or U1254 (N_1254,N_847,N_927);
or U1255 (N_1255,N_828,N_824);
nor U1256 (N_1256,N_553,N_889);
nor U1257 (N_1257,N_544,N_823);
nand U1258 (N_1258,N_815,N_796);
and U1259 (N_1259,N_775,N_778);
nor U1260 (N_1260,N_680,N_760);
or U1261 (N_1261,N_650,N_835);
or U1262 (N_1262,N_704,N_644);
or U1263 (N_1263,N_875,N_640);
xor U1264 (N_1264,N_500,N_950);
and U1265 (N_1265,N_745,N_915);
nand U1266 (N_1266,N_860,N_541);
or U1267 (N_1267,N_764,N_747);
nand U1268 (N_1268,N_562,N_585);
and U1269 (N_1269,N_656,N_791);
or U1270 (N_1270,N_998,N_976);
nand U1271 (N_1271,N_911,N_853);
nand U1272 (N_1272,N_807,N_525);
and U1273 (N_1273,N_949,N_628);
xnor U1274 (N_1274,N_881,N_957);
nor U1275 (N_1275,N_615,N_866);
or U1276 (N_1276,N_953,N_537);
and U1277 (N_1277,N_677,N_929);
or U1278 (N_1278,N_808,N_512);
nor U1279 (N_1279,N_751,N_969);
nand U1280 (N_1280,N_737,N_780);
and U1281 (N_1281,N_995,N_527);
and U1282 (N_1282,N_647,N_530);
and U1283 (N_1283,N_913,N_721);
and U1284 (N_1284,N_987,N_557);
and U1285 (N_1285,N_605,N_543);
nor U1286 (N_1286,N_743,N_608);
nor U1287 (N_1287,N_537,N_874);
nand U1288 (N_1288,N_989,N_659);
nand U1289 (N_1289,N_523,N_746);
and U1290 (N_1290,N_526,N_963);
nand U1291 (N_1291,N_817,N_681);
nor U1292 (N_1292,N_739,N_766);
or U1293 (N_1293,N_879,N_950);
nor U1294 (N_1294,N_740,N_505);
or U1295 (N_1295,N_634,N_671);
nor U1296 (N_1296,N_888,N_524);
or U1297 (N_1297,N_896,N_636);
or U1298 (N_1298,N_737,N_925);
nand U1299 (N_1299,N_554,N_547);
nor U1300 (N_1300,N_755,N_766);
nand U1301 (N_1301,N_684,N_565);
or U1302 (N_1302,N_514,N_901);
or U1303 (N_1303,N_873,N_562);
nand U1304 (N_1304,N_610,N_756);
xor U1305 (N_1305,N_915,N_833);
or U1306 (N_1306,N_590,N_504);
or U1307 (N_1307,N_593,N_649);
and U1308 (N_1308,N_812,N_986);
and U1309 (N_1309,N_689,N_554);
nor U1310 (N_1310,N_880,N_698);
and U1311 (N_1311,N_567,N_763);
nand U1312 (N_1312,N_656,N_926);
and U1313 (N_1313,N_693,N_912);
nand U1314 (N_1314,N_933,N_794);
and U1315 (N_1315,N_787,N_668);
and U1316 (N_1316,N_730,N_830);
or U1317 (N_1317,N_789,N_991);
or U1318 (N_1318,N_928,N_873);
or U1319 (N_1319,N_898,N_701);
and U1320 (N_1320,N_840,N_910);
or U1321 (N_1321,N_620,N_709);
or U1322 (N_1322,N_985,N_783);
or U1323 (N_1323,N_555,N_796);
and U1324 (N_1324,N_523,N_959);
or U1325 (N_1325,N_960,N_708);
nor U1326 (N_1326,N_856,N_769);
or U1327 (N_1327,N_772,N_581);
nor U1328 (N_1328,N_806,N_604);
nand U1329 (N_1329,N_885,N_642);
xnor U1330 (N_1330,N_944,N_740);
nor U1331 (N_1331,N_564,N_569);
xnor U1332 (N_1332,N_522,N_578);
and U1333 (N_1333,N_773,N_951);
nor U1334 (N_1334,N_785,N_950);
nand U1335 (N_1335,N_860,N_668);
and U1336 (N_1336,N_510,N_688);
or U1337 (N_1337,N_597,N_898);
or U1338 (N_1338,N_516,N_753);
nand U1339 (N_1339,N_669,N_902);
nand U1340 (N_1340,N_963,N_854);
nand U1341 (N_1341,N_647,N_692);
nor U1342 (N_1342,N_521,N_532);
or U1343 (N_1343,N_775,N_874);
or U1344 (N_1344,N_926,N_771);
or U1345 (N_1345,N_518,N_558);
nand U1346 (N_1346,N_904,N_594);
and U1347 (N_1347,N_817,N_934);
nor U1348 (N_1348,N_873,N_603);
and U1349 (N_1349,N_899,N_884);
nand U1350 (N_1350,N_601,N_943);
or U1351 (N_1351,N_897,N_703);
or U1352 (N_1352,N_581,N_608);
or U1353 (N_1353,N_774,N_760);
nand U1354 (N_1354,N_919,N_500);
and U1355 (N_1355,N_751,N_766);
and U1356 (N_1356,N_636,N_710);
or U1357 (N_1357,N_892,N_878);
and U1358 (N_1358,N_634,N_710);
or U1359 (N_1359,N_894,N_755);
xnor U1360 (N_1360,N_686,N_727);
nor U1361 (N_1361,N_526,N_623);
nor U1362 (N_1362,N_690,N_750);
nand U1363 (N_1363,N_901,N_654);
nand U1364 (N_1364,N_679,N_817);
or U1365 (N_1365,N_813,N_925);
nand U1366 (N_1366,N_951,N_954);
xor U1367 (N_1367,N_892,N_970);
and U1368 (N_1368,N_707,N_925);
and U1369 (N_1369,N_812,N_969);
or U1370 (N_1370,N_661,N_630);
nor U1371 (N_1371,N_685,N_578);
and U1372 (N_1372,N_904,N_563);
and U1373 (N_1373,N_795,N_626);
nand U1374 (N_1374,N_644,N_539);
and U1375 (N_1375,N_629,N_872);
xor U1376 (N_1376,N_904,N_509);
nand U1377 (N_1377,N_824,N_869);
nand U1378 (N_1378,N_721,N_874);
and U1379 (N_1379,N_960,N_709);
or U1380 (N_1380,N_938,N_782);
and U1381 (N_1381,N_797,N_970);
nor U1382 (N_1382,N_515,N_672);
and U1383 (N_1383,N_682,N_761);
or U1384 (N_1384,N_865,N_842);
and U1385 (N_1385,N_963,N_960);
nor U1386 (N_1386,N_879,N_501);
nor U1387 (N_1387,N_725,N_932);
or U1388 (N_1388,N_953,N_612);
or U1389 (N_1389,N_710,N_541);
xor U1390 (N_1390,N_504,N_776);
nand U1391 (N_1391,N_729,N_569);
and U1392 (N_1392,N_755,N_889);
and U1393 (N_1393,N_851,N_738);
nor U1394 (N_1394,N_518,N_762);
or U1395 (N_1395,N_663,N_968);
nand U1396 (N_1396,N_687,N_870);
and U1397 (N_1397,N_534,N_953);
and U1398 (N_1398,N_766,N_677);
or U1399 (N_1399,N_534,N_666);
nor U1400 (N_1400,N_802,N_616);
nor U1401 (N_1401,N_720,N_864);
nand U1402 (N_1402,N_793,N_859);
nor U1403 (N_1403,N_649,N_881);
or U1404 (N_1404,N_505,N_697);
or U1405 (N_1405,N_622,N_658);
nand U1406 (N_1406,N_689,N_927);
nor U1407 (N_1407,N_611,N_671);
and U1408 (N_1408,N_560,N_602);
and U1409 (N_1409,N_862,N_911);
nor U1410 (N_1410,N_503,N_829);
nand U1411 (N_1411,N_912,N_537);
xor U1412 (N_1412,N_937,N_993);
nand U1413 (N_1413,N_526,N_882);
and U1414 (N_1414,N_526,N_917);
nor U1415 (N_1415,N_849,N_543);
and U1416 (N_1416,N_607,N_599);
nand U1417 (N_1417,N_546,N_561);
and U1418 (N_1418,N_633,N_832);
or U1419 (N_1419,N_786,N_998);
and U1420 (N_1420,N_930,N_937);
and U1421 (N_1421,N_801,N_737);
xor U1422 (N_1422,N_784,N_831);
and U1423 (N_1423,N_758,N_696);
or U1424 (N_1424,N_533,N_593);
or U1425 (N_1425,N_758,N_534);
xnor U1426 (N_1426,N_975,N_771);
nor U1427 (N_1427,N_558,N_884);
xor U1428 (N_1428,N_930,N_654);
nand U1429 (N_1429,N_983,N_745);
xor U1430 (N_1430,N_544,N_517);
xnor U1431 (N_1431,N_834,N_959);
nand U1432 (N_1432,N_733,N_792);
nor U1433 (N_1433,N_732,N_817);
nand U1434 (N_1434,N_998,N_662);
or U1435 (N_1435,N_849,N_876);
nand U1436 (N_1436,N_778,N_959);
or U1437 (N_1437,N_657,N_976);
nand U1438 (N_1438,N_757,N_687);
xnor U1439 (N_1439,N_552,N_529);
nor U1440 (N_1440,N_527,N_729);
nor U1441 (N_1441,N_775,N_833);
nand U1442 (N_1442,N_996,N_703);
nor U1443 (N_1443,N_653,N_634);
nand U1444 (N_1444,N_532,N_595);
xnor U1445 (N_1445,N_952,N_724);
nor U1446 (N_1446,N_837,N_840);
and U1447 (N_1447,N_826,N_740);
nor U1448 (N_1448,N_715,N_819);
or U1449 (N_1449,N_626,N_850);
or U1450 (N_1450,N_867,N_869);
and U1451 (N_1451,N_635,N_794);
nand U1452 (N_1452,N_685,N_940);
and U1453 (N_1453,N_692,N_703);
nor U1454 (N_1454,N_908,N_606);
and U1455 (N_1455,N_912,N_532);
and U1456 (N_1456,N_695,N_657);
or U1457 (N_1457,N_562,N_996);
nand U1458 (N_1458,N_805,N_576);
nand U1459 (N_1459,N_789,N_513);
nor U1460 (N_1460,N_718,N_636);
nand U1461 (N_1461,N_673,N_597);
nand U1462 (N_1462,N_718,N_683);
or U1463 (N_1463,N_538,N_838);
nand U1464 (N_1464,N_762,N_948);
xnor U1465 (N_1465,N_503,N_746);
and U1466 (N_1466,N_539,N_651);
nor U1467 (N_1467,N_993,N_939);
nor U1468 (N_1468,N_908,N_815);
nor U1469 (N_1469,N_548,N_559);
and U1470 (N_1470,N_804,N_860);
or U1471 (N_1471,N_603,N_579);
nand U1472 (N_1472,N_935,N_588);
and U1473 (N_1473,N_886,N_928);
nand U1474 (N_1474,N_843,N_889);
xnor U1475 (N_1475,N_939,N_858);
nor U1476 (N_1476,N_855,N_993);
and U1477 (N_1477,N_588,N_662);
or U1478 (N_1478,N_754,N_508);
or U1479 (N_1479,N_590,N_955);
or U1480 (N_1480,N_777,N_625);
nand U1481 (N_1481,N_711,N_627);
xnor U1482 (N_1482,N_927,N_890);
and U1483 (N_1483,N_706,N_811);
nor U1484 (N_1484,N_664,N_927);
nor U1485 (N_1485,N_790,N_848);
or U1486 (N_1486,N_927,N_586);
nand U1487 (N_1487,N_568,N_748);
xor U1488 (N_1488,N_645,N_534);
xnor U1489 (N_1489,N_910,N_795);
or U1490 (N_1490,N_512,N_943);
nand U1491 (N_1491,N_503,N_631);
xor U1492 (N_1492,N_635,N_773);
nor U1493 (N_1493,N_729,N_595);
nand U1494 (N_1494,N_882,N_727);
and U1495 (N_1495,N_534,N_902);
and U1496 (N_1496,N_668,N_948);
and U1497 (N_1497,N_849,N_678);
nor U1498 (N_1498,N_856,N_536);
nand U1499 (N_1499,N_564,N_778);
nor U1500 (N_1500,N_1025,N_1496);
nor U1501 (N_1501,N_1429,N_1142);
nand U1502 (N_1502,N_1180,N_1056);
nor U1503 (N_1503,N_1086,N_1304);
nand U1504 (N_1504,N_1062,N_1239);
or U1505 (N_1505,N_1139,N_1439);
xor U1506 (N_1506,N_1355,N_1223);
nand U1507 (N_1507,N_1430,N_1396);
nor U1508 (N_1508,N_1410,N_1263);
and U1509 (N_1509,N_1104,N_1254);
or U1510 (N_1510,N_1407,N_1319);
or U1511 (N_1511,N_1315,N_1466);
or U1512 (N_1512,N_1372,N_1053);
or U1513 (N_1513,N_1117,N_1061);
or U1514 (N_1514,N_1494,N_1081);
nor U1515 (N_1515,N_1371,N_1099);
and U1516 (N_1516,N_1215,N_1312);
nand U1517 (N_1517,N_1066,N_1487);
nand U1518 (N_1518,N_1005,N_1275);
or U1519 (N_1519,N_1115,N_1365);
and U1520 (N_1520,N_1435,N_1051);
nor U1521 (N_1521,N_1128,N_1064);
and U1522 (N_1522,N_1185,N_1240);
or U1523 (N_1523,N_1266,N_1002);
and U1524 (N_1524,N_1159,N_1210);
nor U1525 (N_1525,N_1233,N_1307);
and U1526 (N_1526,N_1369,N_1190);
or U1527 (N_1527,N_1088,N_1375);
or U1528 (N_1528,N_1188,N_1449);
nor U1529 (N_1529,N_1224,N_1301);
or U1530 (N_1530,N_1406,N_1399);
and U1531 (N_1531,N_1322,N_1381);
nand U1532 (N_1532,N_1325,N_1391);
and U1533 (N_1533,N_1423,N_1149);
nand U1534 (N_1534,N_1334,N_1231);
nor U1535 (N_1535,N_1182,N_1045);
nand U1536 (N_1536,N_1294,N_1124);
nor U1537 (N_1537,N_1076,N_1237);
or U1538 (N_1538,N_1111,N_1329);
nor U1539 (N_1539,N_1168,N_1013);
or U1540 (N_1540,N_1242,N_1136);
or U1541 (N_1541,N_1065,N_1326);
nand U1542 (N_1542,N_1485,N_1132);
and U1543 (N_1543,N_1107,N_1152);
nor U1544 (N_1544,N_1349,N_1024);
or U1545 (N_1545,N_1269,N_1367);
nand U1546 (N_1546,N_1361,N_1453);
and U1547 (N_1547,N_1141,N_1267);
nor U1548 (N_1548,N_1386,N_1226);
nor U1549 (N_1549,N_1402,N_1222);
nor U1550 (N_1550,N_1278,N_1044);
nand U1551 (N_1551,N_1444,N_1205);
and U1552 (N_1552,N_1379,N_1320);
nand U1553 (N_1553,N_1426,N_1020);
or U1554 (N_1554,N_1360,N_1486);
nor U1555 (N_1555,N_1057,N_1036);
and U1556 (N_1556,N_1248,N_1131);
nand U1557 (N_1557,N_1404,N_1467);
and U1558 (N_1558,N_1472,N_1134);
nor U1559 (N_1559,N_1140,N_1105);
nor U1560 (N_1560,N_1192,N_1475);
nand U1561 (N_1561,N_1255,N_1236);
and U1562 (N_1562,N_1495,N_1470);
or U1563 (N_1563,N_1434,N_1323);
nor U1564 (N_1564,N_1091,N_1345);
nor U1565 (N_1565,N_1098,N_1284);
xor U1566 (N_1566,N_1079,N_1194);
or U1567 (N_1567,N_1452,N_1110);
or U1568 (N_1568,N_1012,N_1216);
or U1569 (N_1569,N_1148,N_1212);
or U1570 (N_1570,N_1422,N_1469);
nand U1571 (N_1571,N_1401,N_1471);
and U1572 (N_1572,N_1283,N_1127);
nor U1573 (N_1573,N_1211,N_1377);
and U1574 (N_1574,N_1067,N_1077);
or U1575 (N_1575,N_1010,N_1374);
nand U1576 (N_1576,N_1271,N_1094);
or U1577 (N_1577,N_1041,N_1172);
and U1578 (N_1578,N_1021,N_1418);
nand U1579 (N_1579,N_1455,N_1290);
nor U1580 (N_1580,N_1464,N_1123);
or U1581 (N_1581,N_1314,N_1093);
or U1582 (N_1582,N_1074,N_1060);
nor U1583 (N_1583,N_1357,N_1114);
nor U1584 (N_1584,N_1150,N_1202);
or U1585 (N_1585,N_1156,N_1438);
nand U1586 (N_1586,N_1293,N_1287);
and U1587 (N_1587,N_1052,N_1414);
and U1588 (N_1588,N_1341,N_1247);
nor U1589 (N_1589,N_1316,N_1209);
nand U1590 (N_1590,N_1344,N_1338);
nor U1591 (N_1591,N_1340,N_1151);
or U1592 (N_1592,N_1299,N_1004);
nand U1593 (N_1593,N_1261,N_1229);
nand U1594 (N_1594,N_1243,N_1448);
nand U1595 (N_1595,N_1443,N_1143);
nor U1596 (N_1596,N_1351,N_1199);
nor U1597 (N_1597,N_1085,N_1161);
nand U1598 (N_1598,N_1029,N_1462);
nand U1599 (N_1599,N_1238,N_1116);
or U1600 (N_1600,N_1480,N_1303);
xor U1601 (N_1601,N_1245,N_1405);
xor U1602 (N_1602,N_1482,N_1441);
xor U1603 (N_1603,N_1001,N_1167);
xor U1604 (N_1604,N_1108,N_1273);
nand U1605 (N_1605,N_1397,N_1125);
nand U1606 (N_1606,N_1217,N_1321);
nand U1607 (N_1607,N_1258,N_1280);
and U1608 (N_1608,N_1183,N_1252);
nor U1609 (N_1609,N_1144,N_1276);
nor U1610 (N_1610,N_1154,N_1129);
and U1611 (N_1611,N_1031,N_1121);
nor U1612 (N_1612,N_1461,N_1366);
xnor U1613 (N_1613,N_1311,N_1090);
and U1614 (N_1614,N_1174,N_1409);
nand U1615 (N_1615,N_1084,N_1383);
nor U1616 (N_1616,N_1011,N_1291);
nand U1617 (N_1617,N_1055,N_1384);
or U1618 (N_1618,N_1126,N_1219);
or U1619 (N_1619,N_1412,N_1416);
and U1620 (N_1620,N_1333,N_1389);
nand U1621 (N_1621,N_1499,N_1153);
nand U1622 (N_1622,N_1437,N_1063);
xnor U1623 (N_1623,N_1264,N_1417);
nor U1624 (N_1624,N_1003,N_1112);
nand U1625 (N_1625,N_1309,N_1100);
or U1626 (N_1626,N_1419,N_1176);
nand U1627 (N_1627,N_1335,N_1048);
nor U1628 (N_1628,N_1122,N_1350);
nor U1629 (N_1629,N_1428,N_1481);
nand U1630 (N_1630,N_1042,N_1353);
and U1631 (N_1631,N_1440,N_1498);
nand U1632 (N_1632,N_1257,N_1208);
or U1633 (N_1633,N_1017,N_1162);
xor U1634 (N_1634,N_1220,N_1015);
nor U1635 (N_1635,N_1187,N_1196);
nand U1636 (N_1636,N_1206,N_1008);
nand U1637 (N_1637,N_1476,N_1424);
nor U1638 (N_1638,N_1398,N_1033);
xnor U1639 (N_1639,N_1177,N_1119);
xnor U1640 (N_1640,N_1071,N_1352);
and U1641 (N_1641,N_1038,N_1392);
or U1642 (N_1642,N_1030,N_1478);
or U1643 (N_1643,N_1225,N_1007);
nand U1644 (N_1644,N_1382,N_1368);
nor U1645 (N_1645,N_1483,N_1492);
and U1646 (N_1646,N_1014,N_1059);
and U1647 (N_1647,N_1343,N_1347);
or U1648 (N_1648,N_1373,N_1427);
nor U1649 (N_1649,N_1262,N_1195);
xnor U1650 (N_1650,N_1274,N_1477);
and U1651 (N_1651,N_1137,N_1318);
nor U1652 (N_1652,N_1327,N_1479);
nand U1653 (N_1653,N_1028,N_1490);
or U1654 (N_1654,N_1456,N_1250);
nand U1655 (N_1655,N_1302,N_1336);
xor U1656 (N_1656,N_1032,N_1000);
or U1657 (N_1657,N_1027,N_1169);
and U1658 (N_1658,N_1468,N_1200);
and U1659 (N_1659,N_1408,N_1308);
nor U1660 (N_1660,N_1420,N_1281);
and U1661 (N_1661,N_1022,N_1346);
or U1662 (N_1662,N_1259,N_1400);
nand U1663 (N_1663,N_1037,N_1279);
nor U1664 (N_1664,N_1376,N_1109);
nand U1665 (N_1665,N_1364,N_1157);
nand U1666 (N_1666,N_1049,N_1313);
nor U1667 (N_1667,N_1181,N_1458);
nand U1668 (N_1668,N_1046,N_1463);
nor U1669 (N_1669,N_1354,N_1043);
or U1670 (N_1670,N_1337,N_1241);
nand U1671 (N_1671,N_1227,N_1097);
nand U1672 (N_1672,N_1083,N_1268);
nor U1673 (N_1673,N_1106,N_1145);
or U1674 (N_1674,N_1411,N_1256);
nand U1675 (N_1675,N_1070,N_1454);
nand U1676 (N_1676,N_1228,N_1034);
and U1677 (N_1677,N_1207,N_1166);
nor U1678 (N_1678,N_1249,N_1186);
nand U1679 (N_1679,N_1101,N_1324);
xnor U1680 (N_1680,N_1089,N_1246);
nand U1681 (N_1681,N_1073,N_1425);
and U1682 (N_1682,N_1019,N_1380);
nor U1683 (N_1683,N_1288,N_1035);
nor U1684 (N_1684,N_1331,N_1253);
xor U1685 (N_1685,N_1431,N_1270);
and U1686 (N_1686,N_1120,N_1218);
xnor U1687 (N_1687,N_1446,N_1072);
xor U1688 (N_1688,N_1138,N_1232);
nor U1689 (N_1689,N_1460,N_1197);
nand U1690 (N_1690,N_1491,N_1272);
and U1691 (N_1691,N_1433,N_1473);
or U1692 (N_1692,N_1450,N_1047);
nand U1693 (N_1693,N_1054,N_1413);
nor U1694 (N_1694,N_1265,N_1078);
xor U1695 (N_1695,N_1358,N_1451);
xor U1696 (N_1696,N_1395,N_1163);
nor U1697 (N_1697,N_1135,N_1075);
and U1698 (N_1698,N_1295,N_1393);
nand U1699 (N_1699,N_1296,N_1175);
and U1700 (N_1700,N_1362,N_1378);
xor U1701 (N_1701,N_1289,N_1103);
xor U1702 (N_1702,N_1363,N_1442);
or U1703 (N_1703,N_1356,N_1221);
and U1704 (N_1704,N_1080,N_1415);
or U1705 (N_1705,N_1390,N_1488);
and U1706 (N_1706,N_1370,N_1191);
nand U1707 (N_1707,N_1465,N_1178);
and U1708 (N_1708,N_1130,N_1213);
nand U1709 (N_1709,N_1204,N_1493);
or U1710 (N_1710,N_1040,N_1147);
xor U1711 (N_1711,N_1459,N_1421);
nand U1712 (N_1712,N_1388,N_1069);
nand U1713 (N_1713,N_1171,N_1203);
nand U1714 (N_1714,N_1244,N_1118);
nand U1715 (N_1715,N_1230,N_1006);
nor U1716 (N_1716,N_1277,N_1058);
nand U1717 (N_1717,N_1018,N_1387);
and U1718 (N_1718,N_1050,N_1317);
or U1719 (N_1719,N_1260,N_1026);
or U1720 (N_1720,N_1039,N_1474);
and U1721 (N_1721,N_1348,N_1328);
or U1722 (N_1722,N_1087,N_1068);
nor U1723 (N_1723,N_1234,N_1385);
nand U1724 (N_1724,N_1447,N_1342);
or U1725 (N_1725,N_1160,N_1432);
nor U1726 (N_1726,N_1023,N_1193);
nor U1727 (N_1727,N_1306,N_1394);
nor U1728 (N_1728,N_1297,N_1146);
nand U1729 (N_1729,N_1305,N_1164);
nand U1730 (N_1730,N_1403,N_1359);
and U1731 (N_1731,N_1095,N_1158);
nor U1732 (N_1732,N_1184,N_1170);
nor U1733 (N_1733,N_1092,N_1285);
and U1734 (N_1734,N_1489,N_1133);
and U1735 (N_1735,N_1165,N_1082);
and U1736 (N_1736,N_1339,N_1310);
nor U1737 (N_1737,N_1300,N_1332);
or U1738 (N_1738,N_1251,N_1214);
and U1739 (N_1739,N_1445,N_1484);
nor U1740 (N_1740,N_1282,N_1457);
nor U1741 (N_1741,N_1102,N_1330);
nand U1742 (N_1742,N_1113,N_1298);
and U1743 (N_1743,N_1292,N_1009);
xnor U1744 (N_1744,N_1235,N_1096);
or U1745 (N_1745,N_1198,N_1173);
nand U1746 (N_1746,N_1497,N_1179);
nand U1747 (N_1747,N_1436,N_1201);
or U1748 (N_1748,N_1189,N_1016);
or U1749 (N_1749,N_1286,N_1155);
or U1750 (N_1750,N_1341,N_1197);
xnor U1751 (N_1751,N_1413,N_1201);
and U1752 (N_1752,N_1469,N_1361);
and U1753 (N_1753,N_1406,N_1322);
nor U1754 (N_1754,N_1035,N_1022);
nor U1755 (N_1755,N_1187,N_1346);
nor U1756 (N_1756,N_1259,N_1255);
or U1757 (N_1757,N_1229,N_1315);
or U1758 (N_1758,N_1190,N_1335);
nor U1759 (N_1759,N_1421,N_1192);
and U1760 (N_1760,N_1327,N_1326);
xor U1761 (N_1761,N_1324,N_1200);
nand U1762 (N_1762,N_1379,N_1483);
nand U1763 (N_1763,N_1339,N_1118);
nand U1764 (N_1764,N_1064,N_1158);
or U1765 (N_1765,N_1021,N_1326);
xnor U1766 (N_1766,N_1333,N_1011);
nand U1767 (N_1767,N_1425,N_1481);
and U1768 (N_1768,N_1069,N_1472);
nand U1769 (N_1769,N_1249,N_1255);
xor U1770 (N_1770,N_1444,N_1309);
xor U1771 (N_1771,N_1483,N_1311);
nand U1772 (N_1772,N_1464,N_1129);
nand U1773 (N_1773,N_1399,N_1402);
nand U1774 (N_1774,N_1125,N_1439);
xnor U1775 (N_1775,N_1079,N_1461);
or U1776 (N_1776,N_1035,N_1314);
nand U1777 (N_1777,N_1469,N_1382);
nor U1778 (N_1778,N_1060,N_1336);
and U1779 (N_1779,N_1414,N_1369);
xor U1780 (N_1780,N_1282,N_1377);
and U1781 (N_1781,N_1436,N_1174);
nor U1782 (N_1782,N_1012,N_1402);
xnor U1783 (N_1783,N_1021,N_1340);
xnor U1784 (N_1784,N_1373,N_1112);
and U1785 (N_1785,N_1096,N_1164);
nor U1786 (N_1786,N_1498,N_1027);
xnor U1787 (N_1787,N_1391,N_1292);
or U1788 (N_1788,N_1063,N_1480);
and U1789 (N_1789,N_1368,N_1304);
or U1790 (N_1790,N_1161,N_1431);
xnor U1791 (N_1791,N_1288,N_1022);
nor U1792 (N_1792,N_1156,N_1106);
nor U1793 (N_1793,N_1252,N_1132);
or U1794 (N_1794,N_1357,N_1152);
xnor U1795 (N_1795,N_1130,N_1320);
and U1796 (N_1796,N_1220,N_1266);
or U1797 (N_1797,N_1326,N_1336);
nor U1798 (N_1798,N_1199,N_1119);
and U1799 (N_1799,N_1440,N_1356);
nand U1800 (N_1800,N_1221,N_1009);
and U1801 (N_1801,N_1296,N_1022);
nand U1802 (N_1802,N_1223,N_1406);
and U1803 (N_1803,N_1300,N_1015);
and U1804 (N_1804,N_1243,N_1224);
and U1805 (N_1805,N_1494,N_1211);
and U1806 (N_1806,N_1237,N_1085);
nor U1807 (N_1807,N_1273,N_1142);
nor U1808 (N_1808,N_1086,N_1208);
and U1809 (N_1809,N_1386,N_1065);
and U1810 (N_1810,N_1388,N_1424);
nor U1811 (N_1811,N_1190,N_1248);
and U1812 (N_1812,N_1109,N_1478);
nand U1813 (N_1813,N_1354,N_1321);
or U1814 (N_1814,N_1308,N_1198);
nor U1815 (N_1815,N_1050,N_1485);
nand U1816 (N_1816,N_1428,N_1291);
xor U1817 (N_1817,N_1370,N_1017);
or U1818 (N_1818,N_1230,N_1350);
or U1819 (N_1819,N_1273,N_1150);
nand U1820 (N_1820,N_1016,N_1065);
nand U1821 (N_1821,N_1207,N_1205);
or U1822 (N_1822,N_1277,N_1038);
xnor U1823 (N_1823,N_1321,N_1249);
nand U1824 (N_1824,N_1209,N_1381);
nand U1825 (N_1825,N_1063,N_1234);
xnor U1826 (N_1826,N_1447,N_1077);
nor U1827 (N_1827,N_1165,N_1127);
and U1828 (N_1828,N_1241,N_1055);
xor U1829 (N_1829,N_1352,N_1457);
or U1830 (N_1830,N_1331,N_1439);
nand U1831 (N_1831,N_1172,N_1337);
or U1832 (N_1832,N_1379,N_1347);
nand U1833 (N_1833,N_1209,N_1283);
xor U1834 (N_1834,N_1259,N_1022);
nor U1835 (N_1835,N_1212,N_1241);
and U1836 (N_1836,N_1416,N_1472);
nor U1837 (N_1837,N_1314,N_1254);
or U1838 (N_1838,N_1388,N_1201);
nand U1839 (N_1839,N_1067,N_1135);
or U1840 (N_1840,N_1015,N_1468);
nand U1841 (N_1841,N_1309,N_1409);
or U1842 (N_1842,N_1432,N_1228);
xnor U1843 (N_1843,N_1346,N_1303);
and U1844 (N_1844,N_1469,N_1320);
or U1845 (N_1845,N_1408,N_1022);
nor U1846 (N_1846,N_1084,N_1356);
and U1847 (N_1847,N_1343,N_1238);
nand U1848 (N_1848,N_1482,N_1460);
nor U1849 (N_1849,N_1285,N_1145);
and U1850 (N_1850,N_1382,N_1365);
and U1851 (N_1851,N_1362,N_1102);
nor U1852 (N_1852,N_1046,N_1068);
and U1853 (N_1853,N_1491,N_1043);
or U1854 (N_1854,N_1233,N_1312);
and U1855 (N_1855,N_1093,N_1486);
and U1856 (N_1856,N_1436,N_1106);
or U1857 (N_1857,N_1231,N_1404);
and U1858 (N_1858,N_1385,N_1486);
nor U1859 (N_1859,N_1324,N_1407);
nor U1860 (N_1860,N_1372,N_1409);
nor U1861 (N_1861,N_1130,N_1056);
nor U1862 (N_1862,N_1374,N_1362);
nand U1863 (N_1863,N_1253,N_1326);
nand U1864 (N_1864,N_1072,N_1470);
and U1865 (N_1865,N_1443,N_1244);
nor U1866 (N_1866,N_1448,N_1454);
and U1867 (N_1867,N_1034,N_1061);
and U1868 (N_1868,N_1332,N_1412);
nor U1869 (N_1869,N_1332,N_1136);
nor U1870 (N_1870,N_1009,N_1263);
nor U1871 (N_1871,N_1201,N_1205);
nand U1872 (N_1872,N_1353,N_1261);
nand U1873 (N_1873,N_1164,N_1117);
xnor U1874 (N_1874,N_1445,N_1037);
or U1875 (N_1875,N_1221,N_1029);
or U1876 (N_1876,N_1455,N_1452);
nor U1877 (N_1877,N_1412,N_1285);
nor U1878 (N_1878,N_1181,N_1269);
xor U1879 (N_1879,N_1220,N_1144);
and U1880 (N_1880,N_1319,N_1363);
nor U1881 (N_1881,N_1314,N_1391);
nand U1882 (N_1882,N_1437,N_1114);
xnor U1883 (N_1883,N_1210,N_1109);
or U1884 (N_1884,N_1008,N_1364);
xor U1885 (N_1885,N_1187,N_1389);
and U1886 (N_1886,N_1465,N_1401);
or U1887 (N_1887,N_1255,N_1028);
and U1888 (N_1888,N_1304,N_1436);
or U1889 (N_1889,N_1251,N_1388);
or U1890 (N_1890,N_1291,N_1452);
and U1891 (N_1891,N_1491,N_1475);
and U1892 (N_1892,N_1125,N_1189);
xnor U1893 (N_1893,N_1171,N_1445);
nor U1894 (N_1894,N_1132,N_1358);
nor U1895 (N_1895,N_1387,N_1213);
xnor U1896 (N_1896,N_1394,N_1397);
nor U1897 (N_1897,N_1345,N_1131);
and U1898 (N_1898,N_1033,N_1418);
and U1899 (N_1899,N_1353,N_1026);
and U1900 (N_1900,N_1338,N_1093);
nor U1901 (N_1901,N_1469,N_1104);
or U1902 (N_1902,N_1321,N_1011);
nor U1903 (N_1903,N_1455,N_1223);
and U1904 (N_1904,N_1341,N_1161);
or U1905 (N_1905,N_1373,N_1267);
nand U1906 (N_1906,N_1152,N_1047);
nand U1907 (N_1907,N_1022,N_1129);
nand U1908 (N_1908,N_1394,N_1020);
or U1909 (N_1909,N_1100,N_1396);
and U1910 (N_1910,N_1040,N_1220);
and U1911 (N_1911,N_1294,N_1426);
or U1912 (N_1912,N_1163,N_1315);
and U1913 (N_1913,N_1195,N_1162);
nand U1914 (N_1914,N_1374,N_1268);
xor U1915 (N_1915,N_1351,N_1188);
or U1916 (N_1916,N_1171,N_1200);
or U1917 (N_1917,N_1341,N_1181);
and U1918 (N_1918,N_1165,N_1168);
nand U1919 (N_1919,N_1153,N_1079);
and U1920 (N_1920,N_1233,N_1067);
or U1921 (N_1921,N_1037,N_1306);
nand U1922 (N_1922,N_1330,N_1164);
nor U1923 (N_1923,N_1260,N_1364);
nand U1924 (N_1924,N_1310,N_1185);
xor U1925 (N_1925,N_1193,N_1107);
or U1926 (N_1926,N_1270,N_1293);
nand U1927 (N_1927,N_1425,N_1027);
nor U1928 (N_1928,N_1003,N_1005);
nand U1929 (N_1929,N_1420,N_1308);
nand U1930 (N_1930,N_1286,N_1013);
or U1931 (N_1931,N_1145,N_1413);
nand U1932 (N_1932,N_1361,N_1006);
nor U1933 (N_1933,N_1054,N_1363);
and U1934 (N_1934,N_1491,N_1331);
nand U1935 (N_1935,N_1234,N_1478);
and U1936 (N_1936,N_1177,N_1156);
nand U1937 (N_1937,N_1241,N_1462);
nor U1938 (N_1938,N_1129,N_1286);
and U1939 (N_1939,N_1369,N_1217);
nor U1940 (N_1940,N_1276,N_1244);
or U1941 (N_1941,N_1038,N_1194);
nand U1942 (N_1942,N_1331,N_1355);
nor U1943 (N_1943,N_1474,N_1162);
or U1944 (N_1944,N_1082,N_1358);
and U1945 (N_1945,N_1176,N_1106);
xor U1946 (N_1946,N_1120,N_1396);
or U1947 (N_1947,N_1097,N_1093);
nor U1948 (N_1948,N_1379,N_1241);
xor U1949 (N_1949,N_1435,N_1371);
or U1950 (N_1950,N_1301,N_1066);
or U1951 (N_1951,N_1051,N_1497);
nand U1952 (N_1952,N_1319,N_1429);
nor U1953 (N_1953,N_1328,N_1487);
and U1954 (N_1954,N_1074,N_1028);
nor U1955 (N_1955,N_1338,N_1397);
nor U1956 (N_1956,N_1344,N_1388);
and U1957 (N_1957,N_1111,N_1069);
nor U1958 (N_1958,N_1400,N_1392);
and U1959 (N_1959,N_1222,N_1073);
and U1960 (N_1960,N_1269,N_1111);
and U1961 (N_1961,N_1387,N_1276);
or U1962 (N_1962,N_1272,N_1216);
nand U1963 (N_1963,N_1441,N_1357);
nand U1964 (N_1964,N_1472,N_1383);
and U1965 (N_1965,N_1497,N_1439);
xor U1966 (N_1966,N_1002,N_1228);
nor U1967 (N_1967,N_1341,N_1217);
and U1968 (N_1968,N_1071,N_1004);
nand U1969 (N_1969,N_1090,N_1496);
nor U1970 (N_1970,N_1381,N_1030);
nor U1971 (N_1971,N_1162,N_1081);
nor U1972 (N_1972,N_1450,N_1362);
xor U1973 (N_1973,N_1231,N_1138);
nor U1974 (N_1974,N_1474,N_1404);
nor U1975 (N_1975,N_1133,N_1449);
nand U1976 (N_1976,N_1016,N_1220);
nor U1977 (N_1977,N_1261,N_1060);
nand U1978 (N_1978,N_1261,N_1038);
or U1979 (N_1979,N_1076,N_1459);
or U1980 (N_1980,N_1294,N_1211);
or U1981 (N_1981,N_1199,N_1095);
xor U1982 (N_1982,N_1219,N_1001);
or U1983 (N_1983,N_1105,N_1489);
nand U1984 (N_1984,N_1344,N_1277);
or U1985 (N_1985,N_1152,N_1069);
xnor U1986 (N_1986,N_1061,N_1144);
nor U1987 (N_1987,N_1443,N_1416);
or U1988 (N_1988,N_1055,N_1372);
or U1989 (N_1989,N_1157,N_1188);
or U1990 (N_1990,N_1181,N_1214);
nand U1991 (N_1991,N_1350,N_1402);
nand U1992 (N_1992,N_1164,N_1354);
and U1993 (N_1993,N_1182,N_1092);
and U1994 (N_1994,N_1283,N_1152);
nand U1995 (N_1995,N_1469,N_1006);
nor U1996 (N_1996,N_1096,N_1142);
and U1997 (N_1997,N_1467,N_1311);
and U1998 (N_1998,N_1438,N_1272);
nor U1999 (N_1999,N_1293,N_1129);
nor U2000 (N_2000,N_1637,N_1528);
and U2001 (N_2001,N_1527,N_1849);
and U2002 (N_2002,N_1788,N_1787);
nor U2003 (N_2003,N_1615,N_1928);
or U2004 (N_2004,N_1634,N_1845);
nand U2005 (N_2005,N_1728,N_1673);
or U2006 (N_2006,N_1661,N_1540);
nor U2007 (N_2007,N_1850,N_1853);
and U2008 (N_2008,N_1708,N_1639);
nor U2009 (N_2009,N_1726,N_1650);
xor U2010 (N_2010,N_1569,N_1821);
nor U2011 (N_2011,N_1858,N_1838);
or U2012 (N_2012,N_1716,N_1738);
or U2013 (N_2013,N_1502,N_1987);
and U2014 (N_2014,N_1605,N_1971);
or U2015 (N_2015,N_1877,N_1684);
or U2016 (N_2016,N_1686,N_1769);
nor U2017 (N_2017,N_1626,N_1953);
nor U2018 (N_2018,N_1718,N_1669);
nand U2019 (N_2019,N_1553,N_1740);
nor U2020 (N_2020,N_1798,N_1510);
nand U2021 (N_2021,N_1520,N_1882);
nand U2022 (N_2022,N_1517,N_1620);
xor U2023 (N_2023,N_1888,N_1980);
nand U2024 (N_2024,N_1733,N_1938);
or U2025 (N_2025,N_1700,N_1796);
nor U2026 (N_2026,N_1759,N_1644);
or U2027 (N_2027,N_1952,N_1786);
and U2028 (N_2028,N_1709,N_1560);
and U2029 (N_2029,N_1568,N_1590);
xor U2030 (N_2030,N_1775,N_1734);
or U2031 (N_2031,N_1864,N_1833);
xor U2032 (N_2032,N_1997,N_1694);
xnor U2033 (N_2033,N_1596,N_1710);
nand U2034 (N_2034,N_1704,N_1585);
nand U2035 (N_2035,N_1978,N_1957);
nand U2036 (N_2036,N_1837,N_1830);
or U2037 (N_2037,N_1998,N_1848);
nor U2038 (N_2038,N_1809,N_1766);
and U2039 (N_2039,N_1599,N_1544);
and U2040 (N_2040,N_1917,N_1536);
or U2041 (N_2041,N_1555,N_1617);
or U2042 (N_2042,N_1688,N_1697);
or U2043 (N_2043,N_1816,N_1801);
nor U2044 (N_2044,N_1587,N_1960);
nand U2045 (N_2045,N_1547,N_1676);
xnor U2046 (N_2046,N_1966,N_1757);
xnor U2047 (N_2047,N_1623,N_1862);
nor U2048 (N_2048,N_1643,N_1925);
or U2049 (N_2049,N_1532,N_1949);
xor U2050 (N_2050,N_1780,N_1525);
xor U2051 (N_2051,N_1577,N_1937);
nor U2052 (N_2052,N_1999,N_1667);
and U2053 (N_2053,N_1974,N_1994);
or U2054 (N_2054,N_1655,N_1905);
nand U2055 (N_2055,N_1526,N_1995);
nand U2056 (N_2056,N_1926,N_1660);
nor U2057 (N_2057,N_1530,N_1887);
xnor U2058 (N_2058,N_1979,N_1598);
nand U2059 (N_2059,N_1556,N_1880);
xor U2060 (N_2060,N_1785,N_1879);
nand U2061 (N_2061,N_1873,N_1962);
and U2062 (N_2062,N_1619,N_1976);
and U2063 (N_2063,N_1600,N_1903);
nor U2064 (N_2064,N_1606,N_1981);
nand U2065 (N_2065,N_1610,N_1908);
nor U2066 (N_2066,N_1703,N_1752);
nand U2067 (N_2067,N_1621,N_1648);
xnor U2068 (N_2068,N_1731,N_1834);
and U2069 (N_2069,N_1561,N_1947);
or U2070 (N_2070,N_1509,N_1699);
nor U2071 (N_2071,N_1940,N_1870);
nand U2072 (N_2072,N_1674,N_1549);
and U2073 (N_2073,N_1725,N_1616);
or U2074 (N_2074,N_1827,N_1678);
and U2075 (N_2075,N_1758,N_1899);
nor U2076 (N_2076,N_1892,N_1832);
nor U2077 (N_2077,N_1854,N_1972);
and U2078 (N_2078,N_1677,N_1931);
nor U2079 (N_2079,N_1872,N_1954);
nand U2080 (N_2080,N_1773,N_1652);
nor U2081 (N_2081,N_1671,N_1601);
and U2082 (N_2082,N_1589,N_1765);
xor U2083 (N_2083,N_1632,N_1715);
and U2084 (N_2084,N_1507,N_1625);
or U2085 (N_2085,N_1665,N_1800);
and U2086 (N_2086,N_1713,N_1578);
and U2087 (N_2087,N_1618,N_1916);
and U2088 (N_2088,N_1878,N_1609);
nor U2089 (N_2089,N_1820,N_1583);
or U2090 (N_2090,N_1542,N_1656);
nand U2091 (N_2091,N_1815,N_1896);
nand U2092 (N_2092,N_1804,N_1777);
or U2093 (N_2093,N_1638,N_1914);
nand U2094 (N_2094,N_1680,N_1748);
or U2095 (N_2095,N_1982,N_1658);
and U2096 (N_2096,N_1582,N_1662);
nand U2097 (N_2097,N_1512,N_1524);
nand U2098 (N_2098,N_1706,N_1941);
and U2099 (N_2099,N_1727,N_1562);
nor U2100 (N_2100,N_1546,N_1965);
nand U2101 (N_2101,N_1581,N_1946);
nor U2102 (N_2102,N_1554,N_1614);
nand U2103 (N_2103,N_1818,N_1519);
and U2104 (N_2104,N_1742,N_1921);
xor U2105 (N_2105,N_1822,N_1831);
or U2106 (N_2106,N_1584,N_1755);
and U2107 (N_2107,N_1735,N_1576);
nor U2108 (N_2108,N_1891,N_1959);
nand U2109 (N_2109,N_1645,N_1557);
nand U2110 (N_2110,N_1642,N_1653);
or U2111 (N_2111,N_1983,N_1746);
xor U2112 (N_2112,N_1712,N_1550);
nand U2113 (N_2113,N_1861,N_1779);
or U2114 (N_2114,N_1573,N_1575);
nor U2115 (N_2115,N_1539,N_1607);
xor U2116 (N_2116,N_1685,N_1679);
and U2117 (N_2117,N_1841,N_1996);
and U2118 (N_2118,N_1548,N_1624);
xor U2119 (N_2119,N_1693,N_1737);
nor U2120 (N_2120,N_1764,N_1687);
xnor U2121 (N_2121,N_1681,N_1958);
or U2122 (N_2122,N_1629,N_1789);
or U2123 (N_2123,N_1967,N_1511);
nand U2124 (N_2124,N_1778,N_1529);
or U2125 (N_2125,N_1729,N_1839);
or U2126 (N_2126,N_1672,N_1935);
or U2127 (N_2127,N_1574,N_1724);
and U2128 (N_2128,N_1559,N_1961);
nand U2129 (N_2129,N_1631,N_1720);
nand U2130 (N_2130,N_1835,N_1739);
or U2131 (N_2131,N_1943,N_1696);
nor U2132 (N_2132,N_1707,N_1771);
nand U2133 (N_2133,N_1889,N_1593);
or U2134 (N_2134,N_1927,N_1945);
nand U2135 (N_2135,N_1791,N_1723);
or U2136 (N_2136,N_1751,N_1866);
or U2137 (N_2137,N_1500,N_1814);
or U2138 (N_2138,N_1990,N_1741);
xnor U2139 (N_2139,N_1803,N_1933);
nand U2140 (N_2140,N_1790,N_1749);
nor U2141 (N_2141,N_1992,N_1613);
nor U2142 (N_2142,N_1915,N_1855);
xor U2143 (N_2143,N_1852,N_1819);
nor U2144 (N_2144,N_1692,N_1951);
and U2145 (N_2145,N_1984,N_1522);
or U2146 (N_2146,N_1719,N_1505);
and U2147 (N_2147,N_1823,N_1942);
and U2148 (N_2148,N_1794,N_1701);
nor U2149 (N_2149,N_1571,N_1840);
and U2150 (N_2150,N_1635,N_1767);
nand U2151 (N_2151,N_1770,N_1811);
or U2152 (N_2152,N_1760,N_1847);
nor U2153 (N_2153,N_1973,N_1813);
or U2154 (N_2154,N_1747,N_1647);
nand U2155 (N_2155,N_1881,N_1675);
nand U2156 (N_2156,N_1913,N_1923);
and U2157 (N_2157,N_1977,N_1970);
nor U2158 (N_2158,N_1641,N_1910);
or U2159 (N_2159,N_1912,N_1893);
and U2160 (N_2160,N_1664,N_1566);
and U2161 (N_2161,N_1843,N_1986);
nand U2162 (N_2162,N_1579,N_1659);
nand U2163 (N_2163,N_1863,N_1636);
and U2164 (N_2164,N_1886,N_1909);
or U2165 (N_2165,N_1963,N_1969);
nor U2166 (N_2166,N_1508,N_1936);
and U2167 (N_2167,N_1776,N_1504);
nand U2168 (N_2168,N_1898,N_1924);
or U2169 (N_2169,N_1572,N_1772);
nand U2170 (N_2170,N_1894,N_1543);
nand U2171 (N_2171,N_1763,N_1901);
or U2172 (N_2172,N_1993,N_1867);
and U2173 (N_2173,N_1663,N_1657);
and U2174 (N_2174,N_1792,N_1603);
nand U2175 (N_2175,N_1782,N_1717);
and U2176 (N_2176,N_1869,N_1797);
nor U2177 (N_2177,N_1828,N_1918);
and U2178 (N_2178,N_1859,N_1812);
xor U2179 (N_2179,N_1907,N_1846);
or U2180 (N_2180,N_1874,N_1513);
nor U2181 (N_2181,N_1552,N_1989);
nand U2182 (N_2182,N_1531,N_1670);
or U2183 (N_2183,N_1691,N_1762);
nor U2184 (N_2184,N_1868,N_1876);
nand U2185 (N_2185,N_1955,N_1934);
nor U2186 (N_2186,N_1690,N_1906);
xnor U2187 (N_2187,N_1612,N_1991);
or U2188 (N_2188,N_1783,N_1950);
and U2189 (N_2189,N_1714,N_1591);
nor U2190 (N_2190,N_1654,N_1922);
and U2191 (N_2191,N_1930,N_1551);
nand U2192 (N_2192,N_1988,N_1948);
nand U2193 (N_2193,N_1829,N_1808);
and U2194 (N_2194,N_1883,N_1856);
or U2195 (N_2195,N_1754,N_1836);
and U2196 (N_2196,N_1592,N_1506);
nand U2197 (N_2197,N_1570,N_1501);
nor U2198 (N_2198,N_1865,N_1793);
or U2199 (N_2199,N_1695,N_1774);
nand U2200 (N_2200,N_1900,N_1781);
or U2201 (N_2201,N_1721,N_1622);
nand U2202 (N_2202,N_1683,N_1649);
nor U2203 (N_2203,N_1968,N_1911);
nand U2204 (N_2204,N_1689,N_1627);
xor U2205 (N_2205,N_1595,N_1975);
or U2206 (N_2206,N_1736,N_1784);
nand U2207 (N_2207,N_1956,N_1515);
or U2208 (N_2208,N_1857,N_1563);
and U2209 (N_2209,N_1860,N_1630);
nor U2210 (N_2210,N_1932,N_1824);
or U2211 (N_2211,N_1698,N_1514);
nor U2212 (N_2212,N_1964,N_1929);
or U2213 (N_2213,N_1985,N_1732);
and U2214 (N_2214,N_1795,N_1640);
nor U2215 (N_2215,N_1939,N_1588);
nor U2216 (N_2216,N_1885,N_1711);
nand U2217 (N_2217,N_1521,N_1537);
or U2218 (N_2218,N_1545,N_1651);
and U2219 (N_2219,N_1602,N_1702);
or U2220 (N_2220,N_1851,N_1810);
nand U2221 (N_2221,N_1753,N_1750);
xor U2222 (N_2222,N_1541,N_1807);
xor U2223 (N_2223,N_1705,N_1565);
nor U2224 (N_2224,N_1730,N_1523);
xor U2225 (N_2225,N_1902,N_1564);
nor U2226 (N_2226,N_1668,N_1567);
nand U2227 (N_2227,N_1920,N_1682);
nand U2228 (N_2228,N_1826,N_1518);
nand U2229 (N_2229,N_1745,N_1756);
xnor U2230 (N_2230,N_1744,N_1761);
nand U2231 (N_2231,N_1628,N_1944);
nor U2232 (N_2232,N_1897,N_1594);
and U2233 (N_2233,N_1597,N_1806);
nor U2234 (N_2234,N_1608,N_1633);
nand U2235 (N_2235,N_1534,N_1799);
or U2236 (N_2236,N_1802,N_1604);
nand U2237 (N_2237,N_1895,N_1611);
or U2238 (N_2238,N_1646,N_1884);
and U2239 (N_2239,N_1825,N_1503);
and U2240 (N_2240,N_1580,N_1871);
and U2241 (N_2241,N_1890,N_1904);
nor U2242 (N_2242,N_1805,N_1558);
xor U2243 (N_2243,N_1722,N_1817);
nor U2244 (N_2244,N_1516,N_1844);
nor U2245 (N_2245,N_1743,N_1666);
and U2246 (N_2246,N_1533,N_1535);
nor U2247 (N_2247,N_1538,N_1842);
or U2248 (N_2248,N_1768,N_1875);
nand U2249 (N_2249,N_1586,N_1919);
nor U2250 (N_2250,N_1816,N_1709);
nand U2251 (N_2251,N_1517,N_1913);
nand U2252 (N_2252,N_1814,N_1970);
nand U2253 (N_2253,N_1634,N_1778);
or U2254 (N_2254,N_1537,N_1788);
and U2255 (N_2255,N_1807,N_1513);
and U2256 (N_2256,N_1908,N_1975);
or U2257 (N_2257,N_1753,N_1839);
nand U2258 (N_2258,N_1950,N_1627);
nand U2259 (N_2259,N_1874,N_1612);
and U2260 (N_2260,N_1802,N_1622);
and U2261 (N_2261,N_1545,N_1993);
nand U2262 (N_2262,N_1971,N_1940);
nand U2263 (N_2263,N_1591,N_1772);
and U2264 (N_2264,N_1847,N_1950);
nand U2265 (N_2265,N_1621,N_1828);
or U2266 (N_2266,N_1930,N_1644);
and U2267 (N_2267,N_1780,N_1524);
or U2268 (N_2268,N_1868,N_1506);
or U2269 (N_2269,N_1932,N_1872);
nor U2270 (N_2270,N_1850,N_1606);
nand U2271 (N_2271,N_1809,N_1713);
xnor U2272 (N_2272,N_1679,N_1660);
or U2273 (N_2273,N_1808,N_1525);
and U2274 (N_2274,N_1857,N_1940);
or U2275 (N_2275,N_1904,N_1534);
nand U2276 (N_2276,N_1858,N_1857);
and U2277 (N_2277,N_1851,N_1842);
or U2278 (N_2278,N_1795,N_1980);
nand U2279 (N_2279,N_1800,N_1924);
and U2280 (N_2280,N_1686,N_1866);
and U2281 (N_2281,N_1562,N_1883);
nor U2282 (N_2282,N_1709,N_1820);
nand U2283 (N_2283,N_1692,N_1533);
nor U2284 (N_2284,N_1763,N_1573);
xor U2285 (N_2285,N_1805,N_1914);
and U2286 (N_2286,N_1579,N_1722);
or U2287 (N_2287,N_1563,N_1574);
nor U2288 (N_2288,N_1661,N_1552);
nor U2289 (N_2289,N_1817,N_1872);
and U2290 (N_2290,N_1741,N_1879);
and U2291 (N_2291,N_1804,N_1763);
or U2292 (N_2292,N_1697,N_1875);
nor U2293 (N_2293,N_1840,N_1993);
and U2294 (N_2294,N_1502,N_1875);
nor U2295 (N_2295,N_1659,N_1980);
xor U2296 (N_2296,N_1765,N_1637);
or U2297 (N_2297,N_1920,N_1680);
or U2298 (N_2298,N_1575,N_1840);
nor U2299 (N_2299,N_1645,N_1542);
or U2300 (N_2300,N_1551,N_1851);
or U2301 (N_2301,N_1505,N_1818);
nand U2302 (N_2302,N_1804,N_1863);
or U2303 (N_2303,N_1541,N_1937);
or U2304 (N_2304,N_1794,N_1852);
nand U2305 (N_2305,N_1612,N_1901);
xor U2306 (N_2306,N_1528,N_1919);
or U2307 (N_2307,N_1536,N_1533);
nand U2308 (N_2308,N_1573,N_1854);
xor U2309 (N_2309,N_1643,N_1988);
xor U2310 (N_2310,N_1973,N_1673);
or U2311 (N_2311,N_1822,N_1931);
nor U2312 (N_2312,N_1882,N_1700);
nand U2313 (N_2313,N_1797,N_1763);
and U2314 (N_2314,N_1975,N_1555);
and U2315 (N_2315,N_1553,N_1833);
nand U2316 (N_2316,N_1850,N_1906);
nor U2317 (N_2317,N_1661,N_1648);
nor U2318 (N_2318,N_1954,N_1506);
or U2319 (N_2319,N_1522,N_1861);
and U2320 (N_2320,N_1544,N_1688);
and U2321 (N_2321,N_1950,N_1933);
nand U2322 (N_2322,N_1849,N_1772);
nand U2323 (N_2323,N_1805,N_1877);
or U2324 (N_2324,N_1760,N_1934);
nand U2325 (N_2325,N_1881,N_1624);
nor U2326 (N_2326,N_1818,N_1908);
nor U2327 (N_2327,N_1650,N_1756);
and U2328 (N_2328,N_1792,N_1523);
and U2329 (N_2329,N_1731,N_1648);
and U2330 (N_2330,N_1937,N_1827);
or U2331 (N_2331,N_1889,N_1536);
nand U2332 (N_2332,N_1862,N_1975);
and U2333 (N_2333,N_1955,N_1627);
or U2334 (N_2334,N_1981,N_1926);
and U2335 (N_2335,N_1642,N_1701);
or U2336 (N_2336,N_1995,N_1949);
nor U2337 (N_2337,N_1718,N_1842);
xnor U2338 (N_2338,N_1893,N_1834);
or U2339 (N_2339,N_1565,N_1907);
and U2340 (N_2340,N_1960,N_1825);
nor U2341 (N_2341,N_1961,N_1865);
nor U2342 (N_2342,N_1775,N_1526);
and U2343 (N_2343,N_1655,N_1836);
nand U2344 (N_2344,N_1866,N_1659);
nand U2345 (N_2345,N_1613,N_1660);
and U2346 (N_2346,N_1522,N_1571);
nand U2347 (N_2347,N_1889,N_1820);
or U2348 (N_2348,N_1663,N_1857);
nand U2349 (N_2349,N_1765,N_1548);
nor U2350 (N_2350,N_1822,N_1525);
or U2351 (N_2351,N_1918,N_1976);
nand U2352 (N_2352,N_1743,N_1599);
or U2353 (N_2353,N_1605,N_1746);
and U2354 (N_2354,N_1774,N_1623);
nor U2355 (N_2355,N_1891,N_1708);
or U2356 (N_2356,N_1798,N_1955);
and U2357 (N_2357,N_1841,N_1917);
and U2358 (N_2358,N_1946,N_1585);
nand U2359 (N_2359,N_1500,N_1778);
or U2360 (N_2360,N_1500,N_1713);
nand U2361 (N_2361,N_1994,N_1629);
and U2362 (N_2362,N_1726,N_1755);
and U2363 (N_2363,N_1626,N_1586);
or U2364 (N_2364,N_1862,N_1954);
or U2365 (N_2365,N_1928,N_1949);
and U2366 (N_2366,N_1657,N_1900);
and U2367 (N_2367,N_1952,N_1724);
and U2368 (N_2368,N_1716,N_1517);
or U2369 (N_2369,N_1567,N_1731);
nor U2370 (N_2370,N_1658,N_1749);
nor U2371 (N_2371,N_1650,N_1899);
nor U2372 (N_2372,N_1756,N_1771);
and U2373 (N_2373,N_1717,N_1698);
nor U2374 (N_2374,N_1856,N_1655);
nand U2375 (N_2375,N_1833,N_1534);
nor U2376 (N_2376,N_1655,N_1852);
or U2377 (N_2377,N_1989,N_1589);
and U2378 (N_2378,N_1703,N_1979);
nor U2379 (N_2379,N_1996,N_1606);
and U2380 (N_2380,N_1701,N_1980);
nand U2381 (N_2381,N_1626,N_1503);
or U2382 (N_2382,N_1549,N_1841);
nor U2383 (N_2383,N_1649,N_1598);
or U2384 (N_2384,N_1631,N_1760);
or U2385 (N_2385,N_1765,N_1726);
or U2386 (N_2386,N_1869,N_1603);
nand U2387 (N_2387,N_1891,N_1965);
nand U2388 (N_2388,N_1879,N_1601);
or U2389 (N_2389,N_1959,N_1752);
and U2390 (N_2390,N_1605,N_1941);
and U2391 (N_2391,N_1770,N_1888);
xor U2392 (N_2392,N_1951,N_1933);
and U2393 (N_2393,N_1806,N_1968);
or U2394 (N_2394,N_1526,N_1653);
and U2395 (N_2395,N_1706,N_1641);
nor U2396 (N_2396,N_1567,N_1992);
and U2397 (N_2397,N_1944,N_1951);
or U2398 (N_2398,N_1561,N_1981);
xor U2399 (N_2399,N_1846,N_1863);
xor U2400 (N_2400,N_1580,N_1579);
and U2401 (N_2401,N_1927,N_1626);
xor U2402 (N_2402,N_1519,N_1729);
and U2403 (N_2403,N_1966,N_1669);
nor U2404 (N_2404,N_1598,N_1657);
and U2405 (N_2405,N_1585,N_1817);
and U2406 (N_2406,N_1675,N_1521);
and U2407 (N_2407,N_1748,N_1731);
xor U2408 (N_2408,N_1824,N_1718);
or U2409 (N_2409,N_1869,N_1881);
nand U2410 (N_2410,N_1650,N_1942);
and U2411 (N_2411,N_1641,N_1767);
nand U2412 (N_2412,N_1957,N_1578);
nor U2413 (N_2413,N_1619,N_1555);
and U2414 (N_2414,N_1862,N_1721);
nor U2415 (N_2415,N_1789,N_1898);
or U2416 (N_2416,N_1688,N_1897);
xnor U2417 (N_2417,N_1593,N_1573);
nand U2418 (N_2418,N_1596,N_1548);
and U2419 (N_2419,N_1886,N_1658);
or U2420 (N_2420,N_1964,N_1838);
nand U2421 (N_2421,N_1962,N_1718);
nor U2422 (N_2422,N_1951,N_1770);
nand U2423 (N_2423,N_1997,N_1862);
nand U2424 (N_2424,N_1563,N_1887);
or U2425 (N_2425,N_1556,N_1953);
nand U2426 (N_2426,N_1808,N_1545);
xor U2427 (N_2427,N_1527,N_1991);
nor U2428 (N_2428,N_1649,N_1946);
nor U2429 (N_2429,N_1779,N_1830);
nand U2430 (N_2430,N_1846,N_1690);
nor U2431 (N_2431,N_1930,N_1592);
nand U2432 (N_2432,N_1523,N_1545);
nand U2433 (N_2433,N_1722,N_1636);
and U2434 (N_2434,N_1974,N_1907);
nand U2435 (N_2435,N_1547,N_1548);
or U2436 (N_2436,N_1683,N_1553);
or U2437 (N_2437,N_1609,N_1962);
or U2438 (N_2438,N_1505,N_1766);
or U2439 (N_2439,N_1706,N_1714);
and U2440 (N_2440,N_1721,N_1579);
nor U2441 (N_2441,N_1615,N_1555);
xnor U2442 (N_2442,N_1928,N_1867);
and U2443 (N_2443,N_1565,N_1921);
or U2444 (N_2444,N_1838,N_1859);
xnor U2445 (N_2445,N_1809,N_1602);
or U2446 (N_2446,N_1557,N_1989);
nand U2447 (N_2447,N_1679,N_1925);
xnor U2448 (N_2448,N_1762,N_1649);
xor U2449 (N_2449,N_1803,N_1846);
and U2450 (N_2450,N_1912,N_1665);
or U2451 (N_2451,N_1772,N_1990);
or U2452 (N_2452,N_1865,N_1638);
xor U2453 (N_2453,N_1851,N_1618);
and U2454 (N_2454,N_1586,N_1861);
or U2455 (N_2455,N_1914,N_1867);
nand U2456 (N_2456,N_1508,N_1838);
or U2457 (N_2457,N_1958,N_1989);
nand U2458 (N_2458,N_1852,N_1754);
nand U2459 (N_2459,N_1677,N_1599);
nor U2460 (N_2460,N_1552,N_1950);
nor U2461 (N_2461,N_1776,N_1625);
nand U2462 (N_2462,N_1848,N_1698);
and U2463 (N_2463,N_1591,N_1785);
nand U2464 (N_2464,N_1679,N_1610);
and U2465 (N_2465,N_1786,N_1981);
nand U2466 (N_2466,N_1629,N_1988);
nor U2467 (N_2467,N_1959,N_1925);
xnor U2468 (N_2468,N_1563,N_1924);
or U2469 (N_2469,N_1772,N_1686);
nor U2470 (N_2470,N_1780,N_1830);
or U2471 (N_2471,N_1990,N_1791);
and U2472 (N_2472,N_1656,N_1720);
nor U2473 (N_2473,N_1662,N_1593);
and U2474 (N_2474,N_1605,N_1821);
nor U2475 (N_2475,N_1836,N_1612);
nor U2476 (N_2476,N_1921,N_1958);
and U2477 (N_2477,N_1835,N_1964);
or U2478 (N_2478,N_1705,N_1806);
nor U2479 (N_2479,N_1925,N_1932);
and U2480 (N_2480,N_1700,N_1988);
nor U2481 (N_2481,N_1838,N_1517);
nor U2482 (N_2482,N_1685,N_1673);
and U2483 (N_2483,N_1520,N_1605);
nand U2484 (N_2484,N_1973,N_1902);
nand U2485 (N_2485,N_1698,N_1941);
nor U2486 (N_2486,N_1848,N_1828);
or U2487 (N_2487,N_1988,N_1753);
xor U2488 (N_2488,N_1996,N_1912);
or U2489 (N_2489,N_1989,N_1777);
nand U2490 (N_2490,N_1773,N_1860);
nor U2491 (N_2491,N_1504,N_1517);
and U2492 (N_2492,N_1930,N_1758);
and U2493 (N_2493,N_1509,N_1821);
and U2494 (N_2494,N_1566,N_1574);
and U2495 (N_2495,N_1806,N_1920);
nor U2496 (N_2496,N_1749,N_1607);
and U2497 (N_2497,N_1944,N_1580);
nor U2498 (N_2498,N_1965,N_1643);
nor U2499 (N_2499,N_1586,N_1970);
xnor U2500 (N_2500,N_2412,N_2023);
and U2501 (N_2501,N_2131,N_2244);
nor U2502 (N_2502,N_2209,N_2175);
or U2503 (N_2503,N_2036,N_2124);
or U2504 (N_2504,N_2317,N_2246);
and U2505 (N_2505,N_2233,N_2190);
nand U2506 (N_2506,N_2204,N_2088);
nand U2507 (N_2507,N_2105,N_2118);
xor U2508 (N_2508,N_2495,N_2197);
or U2509 (N_2509,N_2193,N_2458);
and U2510 (N_2510,N_2098,N_2147);
and U2511 (N_2511,N_2289,N_2433);
xor U2512 (N_2512,N_2082,N_2135);
and U2513 (N_2513,N_2189,N_2092);
or U2514 (N_2514,N_2400,N_2372);
or U2515 (N_2515,N_2043,N_2336);
xor U2516 (N_2516,N_2203,N_2451);
nand U2517 (N_2517,N_2148,N_2079);
nor U2518 (N_2518,N_2051,N_2308);
nand U2519 (N_2519,N_2397,N_2068);
or U2520 (N_2520,N_2060,N_2460);
or U2521 (N_2521,N_2096,N_2008);
nor U2522 (N_2522,N_2173,N_2213);
or U2523 (N_2523,N_2295,N_2125);
nand U2524 (N_2524,N_2026,N_2466);
and U2525 (N_2525,N_2150,N_2112);
nor U2526 (N_2526,N_2083,N_2180);
or U2527 (N_2527,N_2496,N_2330);
nor U2528 (N_2528,N_2354,N_2347);
nor U2529 (N_2529,N_2455,N_2360);
nand U2530 (N_2530,N_2469,N_2061);
or U2531 (N_2531,N_2220,N_2107);
nand U2532 (N_2532,N_2409,N_2086);
nor U2533 (N_2533,N_2375,N_2390);
nor U2534 (N_2534,N_2278,N_2377);
and U2535 (N_2535,N_2471,N_2258);
nand U2536 (N_2536,N_2093,N_2311);
nand U2537 (N_2537,N_2494,N_2369);
and U2538 (N_2538,N_2095,N_2444);
xnor U2539 (N_2539,N_2352,N_2445);
and U2540 (N_2540,N_2235,N_2226);
and U2541 (N_2541,N_2262,N_2172);
nor U2542 (N_2542,N_2000,N_2481);
and U2543 (N_2543,N_2426,N_2006);
nor U2544 (N_2544,N_2356,N_2156);
and U2545 (N_2545,N_2248,N_2241);
nor U2546 (N_2546,N_2019,N_2247);
nor U2547 (N_2547,N_2363,N_2114);
and U2548 (N_2548,N_2253,N_2089);
and U2549 (N_2549,N_2138,N_2414);
or U2550 (N_2550,N_2298,N_2242);
nor U2551 (N_2551,N_2382,N_2130);
nor U2552 (N_2552,N_2070,N_2398);
and U2553 (N_2553,N_2110,N_2475);
nand U2554 (N_2554,N_2388,N_2222);
nand U2555 (N_2555,N_2228,N_2099);
or U2556 (N_2556,N_2044,N_2321);
nand U2557 (N_2557,N_2153,N_2046);
nor U2558 (N_2558,N_2076,N_2304);
nor U2559 (N_2559,N_2436,N_2231);
nand U2560 (N_2560,N_2306,N_2021);
xor U2561 (N_2561,N_2257,N_2421);
nor U2562 (N_2562,N_2208,N_2211);
or U2563 (N_2563,N_2296,N_2029);
nor U2564 (N_2564,N_2492,N_2161);
or U2565 (N_2565,N_2254,N_2285);
nor U2566 (N_2566,N_2126,N_2264);
and U2567 (N_2567,N_2376,N_2343);
or U2568 (N_2568,N_2256,N_2259);
nand U2569 (N_2569,N_2432,N_2178);
nor U2570 (N_2570,N_2380,N_2165);
nand U2571 (N_2571,N_2340,N_2232);
nor U2572 (N_2572,N_2212,N_2443);
nor U2573 (N_2573,N_2215,N_2005);
and U2574 (N_2574,N_2338,N_2195);
nor U2575 (N_2575,N_2462,N_2129);
or U2576 (N_2576,N_2151,N_2411);
or U2577 (N_2577,N_2279,N_2144);
and U2578 (N_2578,N_2163,N_2077);
or U2579 (N_2579,N_2310,N_2162);
or U2580 (N_2580,N_2386,N_2169);
nand U2581 (N_2581,N_2065,N_2030);
nand U2582 (N_2582,N_2331,N_2011);
xnor U2583 (N_2583,N_2478,N_2196);
and U2584 (N_2584,N_2049,N_2337);
or U2585 (N_2585,N_2265,N_2309);
nand U2586 (N_2586,N_2263,N_2188);
nand U2587 (N_2587,N_2355,N_2056);
and U2588 (N_2588,N_2468,N_2224);
nor U2589 (N_2589,N_2484,N_2479);
or U2590 (N_2590,N_2216,N_2450);
nor U2591 (N_2591,N_2305,N_2314);
and U2592 (N_2592,N_2243,N_2123);
nand U2593 (N_2593,N_2327,N_2486);
or U2594 (N_2594,N_2452,N_2234);
nand U2595 (N_2595,N_2250,N_2358);
or U2596 (N_2596,N_2419,N_2498);
and U2597 (N_2597,N_2395,N_2187);
nor U2598 (N_2598,N_2391,N_2072);
xor U2599 (N_2599,N_2361,N_2393);
and U2600 (N_2600,N_2218,N_2035);
and U2601 (N_2601,N_2430,N_2127);
and U2602 (N_2602,N_2027,N_2456);
and U2603 (N_2603,N_2446,N_2183);
and U2604 (N_2604,N_2090,N_2273);
and U2605 (N_2605,N_2344,N_2037);
or U2606 (N_2606,N_2063,N_2066);
xor U2607 (N_2607,N_2128,N_2313);
xnor U2608 (N_2608,N_2202,N_2418);
nand U2609 (N_2609,N_2081,N_2302);
nor U2610 (N_2610,N_2345,N_2389);
and U2611 (N_2611,N_2320,N_2185);
and U2612 (N_2612,N_2240,N_2073);
nor U2613 (N_2613,N_2055,N_2293);
nand U2614 (N_2614,N_2283,N_2157);
or U2615 (N_2615,N_2402,N_2370);
or U2616 (N_2616,N_2275,N_2111);
and U2617 (N_2617,N_2013,N_2424);
and U2618 (N_2618,N_2119,N_2245);
nand U2619 (N_2619,N_2483,N_2058);
and U2620 (N_2620,N_2316,N_2490);
and U2621 (N_2621,N_2297,N_2270);
nor U2622 (N_2622,N_2230,N_2237);
nor U2623 (N_2623,N_2152,N_2015);
and U2624 (N_2624,N_2179,N_2171);
and U2625 (N_2625,N_2201,N_2274);
or U2626 (N_2626,N_2467,N_2214);
and U2627 (N_2627,N_2371,N_2261);
and U2628 (N_2628,N_2407,N_2476);
and U2629 (N_2629,N_2007,N_2210);
xnor U2630 (N_2630,N_2009,N_2342);
or U2631 (N_2631,N_2477,N_2417);
nand U2632 (N_2632,N_2001,N_2227);
and U2633 (N_2633,N_2004,N_2223);
and U2634 (N_2634,N_2074,N_2025);
nor U2635 (N_2635,N_2164,N_2472);
and U2636 (N_2636,N_2034,N_2192);
or U2637 (N_2637,N_2387,N_2016);
or U2638 (N_2638,N_2286,N_2047);
or U2639 (N_2639,N_2453,N_2420);
or U2640 (N_2640,N_2367,N_2206);
or U2641 (N_2641,N_2457,N_2174);
and U2642 (N_2642,N_2441,N_2062);
nor U2643 (N_2643,N_2260,N_2399);
nand U2644 (N_2644,N_2413,N_2143);
nand U2645 (N_2645,N_2291,N_2362);
and U2646 (N_2646,N_2454,N_2028);
nand U2647 (N_2647,N_2113,N_2385);
and U2648 (N_2648,N_2415,N_2022);
or U2649 (N_2649,N_2101,N_2473);
or U2650 (N_2650,N_2280,N_2396);
nand U2651 (N_2651,N_2149,N_2315);
or U2652 (N_2652,N_2348,N_2042);
xnor U2653 (N_2653,N_2333,N_2239);
xor U2654 (N_2654,N_2064,N_2040);
nand U2655 (N_2655,N_2229,N_2039);
or U2656 (N_2656,N_2122,N_2488);
nand U2657 (N_2657,N_2091,N_2405);
or U2658 (N_2658,N_2017,N_2299);
or U2659 (N_2659,N_2429,N_2176);
xor U2660 (N_2660,N_2168,N_2236);
and U2661 (N_2661,N_2085,N_2438);
and U2662 (N_2662,N_2084,N_2384);
nand U2663 (N_2663,N_2133,N_2106);
or U2664 (N_2664,N_2394,N_2136);
and U2665 (N_2665,N_2108,N_2422);
or U2666 (N_2666,N_2109,N_2050);
nand U2667 (N_2667,N_2404,N_2281);
nor U2668 (N_2668,N_2431,N_2470);
and U2669 (N_2669,N_2373,N_2434);
or U2670 (N_2670,N_2020,N_2166);
nor U2671 (N_2671,N_2078,N_2251);
or U2672 (N_2672,N_2031,N_2087);
nand U2673 (N_2673,N_2097,N_2057);
and U2674 (N_2674,N_2284,N_2485);
or U2675 (N_2675,N_2491,N_2059);
nand U2676 (N_2676,N_2219,N_2053);
or U2677 (N_2677,N_2205,N_2014);
and U2678 (N_2678,N_2115,N_2155);
xor U2679 (N_2679,N_2427,N_2252);
nand U2680 (N_2680,N_2401,N_2300);
and U2681 (N_2681,N_2416,N_2364);
nand U2682 (N_2682,N_2403,N_2069);
nand U2683 (N_2683,N_2440,N_2328);
or U2684 (N_2684,N_2071,N_2410);
and U2685 (N_2685,N_2350,N_2121);
or U2686 (N_2686,N_2080,N_2288);
nor U2687 (N_2687,N_2378,N_2447);
nor U2688 (N_2688,N_2357,N_2104);
or U2689 (N_2689,N_2041,N_2489);
and U2690 (N_2690,N_2266,N_2480);
xnor U2691 (N_2691,N_2272,N_2351);
nand U2692 (N_2692,N_2381,N_2319);
and U2693 (N_2693,N_2010,N_2353);
and U2694 (N_2694,N_2465,N_2499);
xnor U2695 (N_2695,N_2103,N_2249);
nor U2696 (N_2696,N_2474,N_2045);
or U2697 (N_2697,N_2437,N_2329);
nand U2698 (N_2698,N_2366,N_2383);
and U2699 (N_2699,N_2221,N_2032);
nand U2700 (N_2700,N_2406,N_2318);
or U2701 (N_2701,N_2054,N_2449);
or U2702 (N_2702,N_2335,N_2100);
nor U2703 (N_2703,N_2238,N_2067);
nand U2704 (N_2704,N_2170,N_2307);
or U2705 (N_2705,N_2198,N_2448);
nand U2706 (N_2706,N_2024,N_2312);
and U2707 (N_2707,N_2167,N_2132);
and U2708 (N_2708,N_2269,N_2374);
and U2709 (N_2709,N_2339,N_2139);
xnor U2710 (N_2710,N_2018,N_2487);
and U2711 (N_2711,N_2075,N_2459);
and U2712 (N_2712,N_2463,N_2217);
or U2713 (N_2713,N_2292,N_2276);
nor U2714 (N_2714,N_2428,N_2365);
nand U2715 (N_2715,N_2181,N_2048);
nand U2716 (N_2716,N_2116,N_2287);
or U2717 (N_2717,N_2301,N_2146);
nand U2718 (N_2718,N_2332,N_2303);
xor U2719 (N_2719,N_2033,N_2094);
and U2720 (N_2720,N_2324,N_2482);
nor U2721 (N_2721,N_2154,N_2493);
or U2722 (N_2722,N_2359,N_2191);
nor U2723 (N_2723,N_2294,N_2497);
or U2724 (N_2724,N_2158,N_2326);
nand U2725 (N_2725,N_2177,N_2439);
nor U2726 (N_2726,N_2282,N_2277);
and U2727 (N_2727,N_2267,N_2145);
xor U2728 (N_2728,N_2159,N_2102);
nand U2729 (N_2729,N_2425,N_2160);
or U2730 (N_2730,N_2200,N_2120);
xnor U2731 (N_2731,N_2117,N_2134);
or U2732 (N_2732,N_2002,N_2290);
nand U2733 (N_2733,N_2408,N_2349);
and U2734 (N_2734,N_2271,N_2140);
or U2735 (N_2735,N_2012,N_2186);
and U2736 (N_2736,N_2141,N_2184);
and U2737 (N_2737,N_2038,N_2182);
or U2738 (N_2738,N_2334,N_2052);
or U2739 (N_2739,N_2142,N_2207);
xor U2740 (N_2740,N_2268,N_2323);
nor U2741 (N_2741,N_2368,N_2325);
nand U2742 (N_2742,N_2423,N_2194);
xor U2743 (N_2743,N_2322,N_2225);
and U2744 (N_2744,N_2461,N_2341);
or U2745 (N_2745,N_2392,N_2464);
and U2746 (N_2746,N_2003,N_2379);
nor U2747 (N_2747,N_2435,N_2442);
xnor U2748 (N_2748,N_2346,N_2137);
and U2749 (N_2749,N_2199,N_2255);
nand U2750 (N_2750,N_2086,N_2252);
nand U2751 (N_2751,N_2395,N_2226);
and U2752 (N_2752,N_2430,N_2212);
nor U2753 (N_2753,N_2163,N_2233);
nand U2754 (N_2754,N_2077,N_2158);
nand U2755 (N_2755,N_2195,N_2255);
or U2756 (N_2756,N_2251,N_2041);
and U2757 (N_2757,N_2269,N_2051);
xnor U2758 (N_2758,N_2244,N_2332);
and U2759 (N_2759,N_2053,N_2457);
nand U2760 (N_2760,N_2416,N_2117);
and U2761 (N_2761,N_2459,N_2428);
nor U2762 (N_2762,N_2469,N_2362);
and U2763 (N_2763,N_2435,N_2036);
nor U2764 (N_2764,N_2002,N_2013);
and U2765 (N_2765,N_2026,N_2420);
nand U2766 (N_2766,N_2127,N_2329);
nand U2767 (N_2767,N_2431,N_2021);
nor U2768 (N_2768,N_2027,N_2177);
nor U2769 (N_2769,N_2231,N_2287);
nand U2770 (N_2770,N_2308,N_2069);
nand U2771 (N_2771,N_2305,N_2076);
nor U2772 (N_2772,N_2230,N_2161);
and U2773 (N_2773,N_2261,N_2407);
or U2774 (N_2774,N_2465,N_2124);
nand U2775 (N_2775,N_2018,N_2127);
nor U2776 (N_2776,N_2044,N_2438);
nor U2777 (N_2777,N_2181,N_2350);
or U2778 (N_2778,N_2265,N_2278);
and U2779 (N_2779,N_2086,N_2238);
xor U2780 (N_2780,N_2455,N_2330);
or U2781 (N_2781,N_2432,N_2320);
and U2782 (N_2782,N_2014,N_2156);
and U2783 (N_2783,N_2082,N_2487);
nor U2784 (N_2784,N_2074,N_2140);
xor U2785 (N_2785,N_2104,N_2150);
xnor U2786 (N_2786,N_2177,N_2230);
nand U2787 (N_2787,N_2279,N_2282);
or U2788 (N_2788,N_2220,N_2198);
or U2789 (N_2789,N_2204,N_2491);
nand U2790 (N_2790,N_2201,N_2352);
and U2791 (N_2791,N_2120,N_2382);
nand U2792 (N_2792,N_2392,N_2289);
xnor U2793 (N_2793,N_2443,N_2371);
nand U2794 (N_2794,N_2002,N_2061);
and U2795 (N_2795,N_2010,N_2484);
and U2796 (N_2796,N_2406,N_2272);
xnor U2797 (N_2797,N_2035,N_2428);
nor U2798 (N_2798,N_2294,N_2439);
and U2799 (N_2799,N_2380,N_2079);
nor U2800 (N_2800,N_2177,N_2443);
or U2801 (N_2801,N_2316,N_2326);
or U2802 (N_2802,N_2317,N_2082);
and U2803 (N_2803,N_2007,N_2085);
nand U2804 (N_2804,N_2330,N_2061);
nand U2805 (N_2805,N_2184,N_2481);
and U2806 (N_2806,N_2427,N_2177);
xor U2807 (N_2807,N_2146,N_2311);
or U2808 (N_2808,N_2130,N_2235);
or U2809 (N_2809,N_2151,N_2337);
or U2810 (N_2810,N_2106,N_2425);
nor U2811 (N_2811,N_2287,N_2054);
or U2812 (N_2812,N_2106,N_2464);
and U2813 (N_2813,N_2388,N_2282);
or U2814 (N_2814,N_2053,N_2149);
nand U2815 (N_2815,N_2237,N_2077);
nand U2816 (N_2816,N_2082,N_2352);
and U2817 (N_2817,N_2285,N_2170);
and U2818 (N_2818,N_2335,N_2475);
nand U2819 (N_2819,N_2011,N_2438);
nor U2820 (N_2820,N_2417,N_2497);
and U2821 (N_2821,N_2203,N_2297);
xnor U2822 (N_2822,N_2417,N_2182);
nand U2823 (N_2823,N_2081,N_2462);
xor U2824 (N_2824,N_2296,N_2344);
nand U2825 (N_2825,N_2412,N_2105);
and U2826 (N_2826,N_2322,N_2259);
or U2827 (N_2827,N_2422,N_2411);
nor U2828 (N_2828,N_2046,N_2065);
or U2829 (N_2829,N_2401,N_2243);
and U2830 (N_2830,N_2293,N_2062);
nor U2831 (N_2831,N_2005,N_2308);
nor U2832 (N_2832,N_2453,N_2305);
nor U2833 (N_2833,N_2076,N_2460);
xnor U2834 (N_2834,N_2301,N_2205);
xor U2835 (N_2835,N_2160,N_2025);
or U2836 (N_2836,N_2420,N_2032);
nor U2837 (N_2837,N_2163,N_2385);
nor U2838 (N_2838,N_2433,N_2276);
nand U2839 (N_2839,N_2305,N_2172);
nand U2840 (N_2840,N_2292,N_2484);
nor U2841 (N_2841,N_2426,N_2110);
or U2842 (N_2842,N_2132,N_2434);
nand U2843 (N_2843,N_2219,N_2254);
nand U2844 (N_2844,N_2094,N_2254);
and U2845 (N_2845,N_2483,N_2329);
xnor U2846 (N_2846,N_2000,N_2054);
nand U2847 (N_2847,N_2012,N_2040);
or U2848 (N_2848,N_2314,N_2147);
nor U2849 (N_2849,N_2060,N_2009);
xor U2850 (N_2850,N_2022,N_2469);
or U2851 (N_2851,N_2086,N_2305);
xor U2852 (N_2852,N_2264,N_2292);
and U2853 (N_2853,N_2236,N_2287);
nand U2854 (N_2854,N_2233,N_2236);
or U2855 (N_2855,N_2494,N_2391);
nand U2856 (N_2856,N_2026,N_2393);
or U2857 (N_2857,N_2446,N_2167);
nor U2858 (N_2858,N_2439,N_2422);
xnor U2859 (N_2859,N_2023,N_2089);
nand U2860 (N_2860,N_2177,N_2287);
nor U2861 (N_2861,N_2436,N_2299);
or U2862 (N_2862,N_2333,N_2283);
nor U2863 (N_2863,N_2279,N_2286);
or U2864 (N_2864,N_2316,N_2480);
nand U2865 (N_2865,N_2373,N_2061);
or U2866 (N_2866,N_2068,N_2272);
nor U2867 (N_2867,N_2111,N_2212);
nor U2868 (N_2868,N_2009,N_2067);
nand U2869 (N_2869,N_2270,N_2397);
nand U2870 (N_2870,N_2452,N_2356);
and U2871 (N_2871,N_2055,N_2494);
and U2872 (N_2872,N_2305,N_2171);
or U2873 (N_2873,N_2064,N_2174);
nand U2874 (N_2874,N_2396,N_2442);
nor U2875 (N_2875,N_2194,N_2356);
nor U2876 (N_2876,N_2398,N_2199);
nand U2877 (N_2877,N_2064,N_2336);
xnor U2878 (N_2878,N_2339,N_2103);
or U2879 (N_2879,N_2362,N_2432);
and U2880 (N_2880,N_2380,N_2309);
or U2881 (N_2881,N_2191,N_2160);
nand U2882 (N_2882,N_2126,N_2054);
xor U2883 (N_2883,N_2296,N_2096);
and U2884 (N_2884,N_2277,N_2083);
and U2885 (N_2885,N_2301,N_2468);
xnor U2886 (N_2886,N_2174,N_2483);
or U2887 (N_2887,N_2093,N_2095);
nand U2888 (N_2888,N_2067,N_2292);
nor U2889 (N_2889,N_2433,N_2305);
and U2890 (N_2890,N_2301,N_2418);
xnor U2891 (N_2891,N_2413,N_2075);
or U2892 (N_2892,N_2352,N_2105);
or U2893 (N_2893,N_2435,N_2232);
nand U2894 (N_2894,N_2497,N_2372);
or U2895 (N_2895,N_2079,N_2067);
nor U2896 (N_2896,N_2315,N_2283);
nand U2897 (N_2897,N_2125,N_2450);
and U2898 (N_2898,N_2306,N_2067);
or U2899 (N_2899,N_2066,N_2292);
nand U2900 (N_2900,N_2414,N_2217);
nand U2901 (N_2901,N_2404,N_2495);
nor U2902 (N_2902,N_2419,N_2302);
xor U2903 (N_2903,N_2225,N_2105);
nand U2904 (N_2904,N_2357,N_2176);
nor U2905 (N_2905,N_2447,N_2188);
nand U2906 (N_2906,N_2197,N_2166);
and U2907 (N_2907,N_2228,N_2258);
nor U2908 (N_2908,N_2035,N_2437);
or U2909 (N_2909,N_2417,N_2008);
nor U2910 (N_2910,N_2133,N_2187);
or U2911 (N_2911,N_2282,N_2362);
nand U2912 (N_2912,N_2076,N_2186);
or U2913 (N_2913,N_2402,N_2361);
nor U2914 (N_2914,N_2108,N_2106);
xor U2915 (N_2915,N_2477,N_2302);
nand U2916 (N_2916,N_2218,N_2461);
and U2917 (N_2917,N_2455,N_2248);
nor U2918 (N_2918,N_2042,N_2437);
and U2919 (N_2919,N_2285,N_2184);
or U2920 (N_2920,N_2003,N_2119);
and U2921 (N_2921,N_2278,N_2052);
or U2922 (N_2922,N_2283,N_2323);
xnor U2923 (N_2923,N_2326,N_2264);
nand U2924 (N_2924,N_2372,N_2192);
or U2925 (N_2925,N_2472,N_2182);
nand U2926 (N_2926,N_2432,N_2077);
or U2927 (N_2927,N_2253,N_2161);
and U2928 (N_2928,N_2145,N_2483);
or U2929 (N_2929,N_2264,N_2062);
and U2930 (N_2930,N_2446,N_2371);
nand U2931 (N_2931,N_2388,N_2000);
xnor U2932 (N_2932,N_2111,N_2318);
and U2933 (N_2933,N_2467,N_2031);
and U2934 (N_2934,N_2112,N_2347);
nor U2935 (N_2935,N_2050,N_2048);
nand U2936 (N_2936,N_2151,N_2080);
and U2937 (N_2937,N_2415,N_2031);
nand U2938 (N_2938,N_2410,N_2024);
or U2939 (N_2939,N_2482,N_2340);
nor U2940 (N_2940,N_2358,N_2300);
nor U2941 (N_2941,N_2342,N_2387);
nor U2942 (N_2942,N_2431,N_2276);
nand U2943 (N_2943,N_2010,N_2381);
nand U2944 (N_2944,N_2323,N_2176);
or U2945 (N_2945,N_2480,N_2479);
nand U2946 (N_2946,N_2087,N_2047);
xor U2947 (N_2947,N_2139,N_2143);
nand U2948 (N_2948,N_2271,N_2179);
nand U2949 (N_2949,N_2093,N_2294);
nor U2950 (N_2950,N_2415,N_2000);
or U2951 (N_2951,N_2322,N_2114);
and U2952 (N_2952,N_2066,N_2465);
nand U2953 (N_2953,N_2250,N_2244);
nand U2954 (N_2954,N_2028,N_2259);
nand U2955 (N_2955,N_2336,N_2180);
nor U2956 (N_2956,N_2066,N_2381);
xor U2957 (N_2957,N_2427,N_2066);
nor U2958 (N_2958,N_2124,N_2092);
nand U2959 (N_2959,N_2157,N_2191);
and U2960 (N_2960,N_2082,N_2490);
xor U2961 (N_2961,N_2086,N_2399);
nor U2962 (N_2962,N_2403,N_2184);
nor U2963 (N_2963,N_2235,N_2234);
or U2964 (N_2964,N_2422,N_2458);
and U2965 (N_2965,N_2024,N_2079);
or U2966 (N_2966,N_2032,N_2113);
xnor U2967 (N_2967,N_2383,N_2203);
or U2968 (N_2968,N_2127,N_2405);
nor U2969 (N_2969,N_2132,N_2210);
or U2970 (N_2970,N_2278,N_2007);
xor U2971 (N_2971,N_2328,N_2478);
or U2972 (N_2972,N_2220,N_2466);
xnor U2973 (N_2973,N_2206,N_2422);
nor U2974 (N_2974,N_2164,N_2241);
nand U2975 (N_2975,N_2372,N_2213);
or U2976 (N_2976,N_2068,N_2053);
and U2977 (N_2977,N_2180,N_2009);
or U2978 (N_2978,N_2495,N_2274);
nor U2979 (N_2979,N_2396,N_2307);
nand U2980 (N_2980,N_2173,N_2379);
and U2981 (N_2981,N_2380,N_2417);
nor U2982 (N_2982,N_2488,N_2372);
and U2983 (N_2983,N_2386,N_2142);
xnor U2984 (N_2984,N_2023,N_2447);
or U2985 (N_2985,N_2254,N_2267);
or U2986 (N_2986,N_2319,N_2265);
nor U2987 (N_2987,N_2235,N_2455);
and U2988 (N_2988,N_2244,N_2027);
and U2989 (N_2989,N_2352,N_2011);
nand U2990 (N_2990,N_2060,N_2144);
nor U2991 (N_2991,N_2307,N_2113);
and U2992 (N_2992,N_2084,N_2321);
nand U2993 (N_2993,N_2149,N_2335);
or U2994 (N_2994,N_2191,N_2463);
xor U2995 (N_2995,N_2224,N_2128);
nor U2996 (N_2996,N_2304,N_2062);
and U2997 (N_2997,N_2179,N_2309);
or U2998 (N_2998,N_2337,N_2183);
or U2999 (N_2999,N_2319,N_2151);
nand U3000 (N_3000,N_2509,N_2609);
or U3001 (N_3001,N_2815,N_2947);
xnor U3002 (N_3002,N_2805,N_2533);
or U3003 (N_3003,N_2573,N_2576);
xor U3004 (N_3004,N_2714,N_2799);
nor U3005 (N_3005,N_2830,N_2593);
xnor U3006 (N_3006,N_2787,N_2933);
or U3007 (N_3007,N_2530,N_2878);
or U3008 (N_3008,N_2606,N_2750);
xnor U3009 (N_3009,N_2546,N_2776);
nand U3010 (N_3010,N_2884,N_2702);
and U3011 (N_3011,N_2508,N_2529);
nor U3012 (N_3012,N_2595,N_2746);
nand U3013 (N_3013,N_2832,N_2782);
and U3014 (N_3014,N_2558,N_2737);
or U3015 (N_3015,N_2734,N_2517);
nor U3016 (N_3016,N_2999,N_2589);
nor U3017 (N_3017,N_2564,N_2591);
nand U3018 (N_3018,N_2671,N_2722);
or U3019 (N_3019,N_2888,N_2630);
and U3020 (N_3020,N_2553,N_2755);
xnor U3021 (N_3021,N_2911,N_2792);
nand U3022 (N_3022,N_2917,N_2940);
xor U3023 (N_3023,N_2550,N_2623);
and U3024 (N_3024,N_2730,N_2869);
nor U3025 (N_3025,N_2883,N_2524);
nor U3026 (N_3026,N_2932,N_2634);
nand U3027 (N_3027,N_2675,N_2541);
and U3028 (N_3028,N_2763,N_2982);
nand U3029 (N_3029,N_2708,N_2682);
nand U3030 (N_3030,N_2626,N_2753);
or U3031 (N_3031,N_2861,N_2959);
xor U3032 (N_3032,N_2752,N_2654);
xor U3033 (N_3033,N_2621,N_2724);
xnor U3034 (N_3034,N_2871,N_2960);
nor U3035 (N_3035,N_2681,N_2662);
nor U3036 (N_3036,N_2742,N_2653);
and U3037 (N_3037,N_2731,N_2904);
nand U3038 (N_3038,N_2759,N_2797);
or U3039 (N_3039,N_2539,N_2928);
nand U3040 (N_3040,N_2818,N_2918);
nand U3041 (N_3041,N_2645,N_2608);
and U3042 (N_3042,N_2984,N_2758);
and U3043 (N_3043,N_2780,N_2810);
nor U3044 (N_3044,N_2605,N_2976);
nor U3045 (N_3045,N_2680,N_2774);
and U3046 (N_3046,N_2728,N_2821);
and U3047 (N_3047,N_2851,N_2747);
nor U3048 (N_3048,N_2824,N_2924);
and U3049 (N_3049,N_2813,N_2899);
and U3050 (N_3050,N_2562,N_2538);
and U3051 (N_3051,N_2971,N_2685);
nor U3052 (N_3052,N_2537,N_2577);
or U3053 (N_3053,N_2751,N_2580);
nand U3054 (N_3054,N_2555,N_2726);
nor U3055 (N_3055,N_2571,N_2563);
xor U3056 (N_3056,N_2578,N_2594);
xnor U3057 (N_3057,N_2567,N_2514);
and U3058 (N_3058,N_2570,N_2798);
nor U3059 (N_3059,N_2891,N_2738);
nor U3060 (N_3060,N_2896,N_2543);
or U3061 (N_3061,N_2867,N_2895);
or U3062 (N_3062,N_2913,N_2996);
nand U3063 (N_3063,N_2856,N_2719);
or U3064 (N_3064,N_2831,N_2523);
or U3065 (N_3065,N_2819,N_2705);
and U3066 (N_3066,N_2762,N_2767);
xnor U3067 (N_3067,N_2893,N_2687);
nand U3068 (N_3068,N_2993,N_2968);
xnor U3069 (N_3069,N_2784,N_2688);
nor U3070 (N_3070,N_2859,N_2502);
and U3071 (N_3071,N_2709,N_2790);
and U3072 (N_3072,N_2603,N_2644);
xor U3073 (N_3073,N_2711,N_2771);
nand U3074 (N_3074,N_2665,N_2789);
or U3075 (N_3075,N_2733,N_2816);
and U3076 (N_3076,N_2693,N_2811);
xnor U3077 (N_3077,N_2710,N_2812);
xnor U3078 (N_3078,N_2766,N_2833);
nand U3079 (N_3079,N_2900,N_2663);
nor U3080 (N_3080,N_2761,N_2616);
or U3081 (N_3081,N_2857,N_2977);
and U3082 (N_3082,N_2631,N_2843);
nor U3083 (N_3083,N_2721,N_2949);
and U3084 (N_3084,N_2920,N_2997);
nor U3085 (N_3085,N_2720,N_2732);
nand U3086 (N_3086,N_2638,N_2951);
nor U3087 (N_3087,N_2527,N_2979);
and U3088 (N_3088,N_2690,N_2848);
or U3089 (N_3089,N_2660,N_2769);
and U3090 (N_3090,N_2736,N_2903);
nand U3091 (N_3091,N_2651,N_2703);
or U3092 (N_3092,N_2611,N_2520);
and U3093 (N_3093,N_2600,N_2559);
xor U3094 (N_3094,N_2915,N_2985);
and U3095 (N_3095,N_2568,N_2822);
nand U3096 (N_3096,N_2599,N_2664);
nor U3097 (N_3097,N_2872,N_2828);
xor U3098 (N_3098,N_2873,N_2936);
or U3099 (N_3099,N_2639,N_2975);
nor U3100 (N_3100,N_2672,N_2522);
nor U3101 (N_3101,N_2542,N_2670);
or U3102 (N_3102,N_2518,N_2863);
xor U3103 (N_3103,N_2881,N_2916);
nor U3104 (N_3104,N_2588,N_2998);
xnor U3105 (N_3105,N_2614,N_2788);
or U3106 (N_3106,N_2974,N_2640);
or U3107 (N_3107,N_2648,N_2908);
and U3108 (N_3108,N_2513,N_2622);
or U3109 (N_3109,N_2768,N_2849);
nor U3110 (N_3110,N_2879,N_2992);
nand U3111 (N_3111,N_2507,N_2842);
xnor U3112 (N_3112,N_2596,N_2938);
nand U3113 (N_3113,N_2673,N_2519);
nor U3114 (N_3114,N_2739,N_2749);
and U3115 (N_3115,N_2583,N_2607);
and U3116 (N_3116,N_2549,N_2910);
nand U3117 (N_3117,N_2635,N_2686);
and U3118 (N_3118,N_2579,N_2852);
nand U3119 (N_3119,N_2696,N_2661);
xor U3120 (N_3120,N_2692,N_2882);
or U3121 (N_3121,N_2793,N_2941);
or U3122 (N_3122,N_2946,N_2741);
xor U3123 (N_3123,N_2735,N_2919);
or U3124 (N_3124,N_2590,N_2862);
nand U3125 (N_3125,N_2802,N_2560);
and U3126 (N_3126,N_2887,N_2500);
or U3127 (N_3127,N_2937,N_2796);
or U3128 (N_3128,N_2547,N_2925);
or U3129 (N_3129,N_2566,N_2698);
nor U3130 (N_3130,N_2987,N_2855);
nand U3131 (N_3131,N_2952,N_2966);
and U3132 (N_3132,N_2674,N_2958);
nand U3133 (N_3133,N_2876,N_2647);
nor U3134 (N_3134,N_2834,N_2754);
nor U3135 (N_3135,N_2597,N_2505);
or U3136 (N_3136,N_2934,N_2850);
nand U3137 (N_3137,N_2989,N_2886);
and U3138 (N_3138,N_2545,N_2953);
nor U3139 (N_3139,N_2718,N_2874);
or U3140 (N_3140,N_2858,N_2864);
and U3141 (N_3141,N_2572,N_2620);
xor U3142 (N_3142,N_2526,N_2967);
xnor U3143 (N_3143,N_2624,N_2561);
and U3144 (N_3144,N_2649,N_2748);
or U3145 (N_3145,N_2652,N_2847);
or U3146 (N_3146,N_2534,N_2585);
nor U3147 (N_3147,N_2957,N_2961);
or U3148 (N_3148,N_2945,N_2898);
or U3149 (N_3149,N_2825,N_2897);
xor U3150 (N_3150,N_2785,N_2803);
xnor U3151 (N_3151,N_2677,N_2691);
or U3152 (N_3152,N_2689,N_2587);
and U3153 (N_3153,N_2723,N_2781);
nor U3154 (N_3154,N_2978,N_2844);
nor U3155 (N_3155,N_2808,N_2980);
nand U3156 (N_3156,N_2865,N_2536);
nor U3157 (N_3157,N_2618,N_2637);
or U3158 (N_3158,N_2613,N_2772);
and U3159 (N_3159,N_2981,N_2632);
nand U3160 (N_3160,N_2551,N_2922);
or U3161 (N_3161,N_2679,N_2729);
xnor U3162 (N_3162,N_2791,N_2592);
nor U3163 (N_3163,N_2773,N_2510);
nand U3164 (N_3164,N_2656,N_2697);
xor U3165 (N_3165,N_2806,N_2795);
or U3166 (N_3166,N_2535,N_2659);
xnor U3167 (N_3167,N_2939,N_2716);
or U3168 (N_3168,N_2826,N_2854);
or U3169 (N_3169,N_2612,N_2926);
or U3170 (N_3170,N_2646,N_2501);
nor U3171 (N_3171,N_2744,N_2516);
nand U3172 (N_3172,N_2548,N_2515);
nor U3173 (N_3173,N_2923,N_2950);
nor U3174 (N_3174,N_2701,N_2610);
or U3175 (N_3175,N_2912,N_2694);
nor U3176 (N_3176,N_2617,N_2704);
nor U3177 (N_3177,N_2964,N_2540);
nand U3178 (N_3178,N_2633,N_2707);
nor U3179 (N_3179,N_2532,N_2713);
nor U3180 (N_3180,N_2853,N_2629);
and U3181 (N_3181,N_2521,N_2511);
nand U3182 (N_3182,N_2699,N_2875);
nand U3183 (N_3183,N_2846,N_2779);
and U3184 (N_3184,N_2804,N_2667);
nand U3185 (N_3185,N_2777,N_2956);
or U3186 (N_3186,N_2727,N_2948);
or U3187 (N_3187,N_2942,N_2764);
xnor U3188 (N_3188,N_2683,N_2581);
and U3189 (N_3189,N_2955,N_2914);
nand U3190 (N_3190,N_2909,N_2760);
or U3191 (N_3191,N_2794,N_2885);
nor U3192 (N_3192,N_2829,N_2642);
xnor U3193 (N_3193,N_2528,N_2552);
and U3194 (N_3194,N_2625,N_2531);
and U3195 (N_3195,N_2817,N_2866);
or U3196 (N_3196,N_2569,N_2619);
or U3197 (N_3197,N_2725,N_2770);
xor U3198 (N_3198,N_2657,N_2706);
and U3199 (N_3199,N_2839,N_2930);
or U3200 (N_3200,N_2889,N_2901);
or U3201 (N_3201,N_2666,N_2743);
or U3202 (N_3202,N_2860,N_2944);
or U3203 (N_3203,N_2700,N_2991);
or U3204 (N_3204,N_2927,N_2756);
and U3205 (N_3205,N_2807,N_2963);
or U3206 (N_3206,N_2643,N_2604);
and U3207 (N_3207,N_2943,N_2668);
nand U3208 (N_3208,N_2557,N_2814);
or U3209 (N_3209,N_2827,N_2972);
xnor U3210 (N_3210,N_2877,N_2929);
xor U3211 (N_3211,N_2506,N_2835);
nand U3212 (N_3212,N_2954,N_2973);
and U3213 (N_3213,N_2868,N_2601);
or U3214 (N_3214,N_2556,N_2554);
and U3215 (N_3215,N_2503,N_2575);
nor U3216 (N_3216,N_2740,N_2931);
nand U3217 (N_3217,N_2783,N_2598);
nor U3218 (N_3218,N_2820,N_2717);
and U3219 (N_3219,N_2650,N_2544);
nor U3220 (N_3220,N_2676,N_2584);
or U3221 (N_3221,N_2836,N_2907);
xor U3222 (N_3222,N_2986,N_2837);
and U3223 (N_3223,N_2655,N_2983);
nand U3224 (N_3224,N_2669,N_2905);
nand U3225 (N_3225,N_2512,N_2628);
nand U3226 (N_3226,N_2602,N_2880);
and U3227 (N_3227,N_2800,N_2765);
nand U3228 (N_3228,N_2823,N_2935);
nor U3229 (N_3229,N_2775,N_2894);
or U3230 (N_3230,N_2890,N_2565);
and U3231 (N_3231,N_2962,N_2641);
or U3232 (N_3232,N_2525,N_2838);
and U3233 (N_3233,N_2586,N_2684);
or U3234 (N_3234,N_2615,N_2845);
nor U3235 (N_3235,N_2636,N_2921);
nor U3236 (N_3236,N_2574,N_2582);
nor U3237 (N_3237,N_2840,N_2627);
nand U3238 (N_3238,N_2990,N_2892);
nor U3239 (N_3239,N_2994,N_2786);
and U3240 (N_3240,N_2801,N_2841);
and U3241 (N_3241,N_2970,N_2712);
nor U3242 (N_3242,N_2715,N_2965);
and U3243 (N_3243,N_2745,N_2969);
nor U3244 (N_3244,N_2988,N_2902);
and U3245 (N_3245,N_2504,N_2757);
and U3246 (N_3246,N_2809,N_2778);
or U3247 (N_3247,N_2870,N_2995);
or U3248 (N_3248,N_2678,N_2695);
xor U3249 (N_3249,N_2906,N_2658);
or U3250 (N_3250,N_2871,N_2596);
and U3251 (N_3251,N_2524,N_2780);
xnor U3252 (N_3252,N_2659,N_2770);
nor U3253 (N_3253,N_2964,N_2959);
nor U3254 (N_3254,N_2993,N_2521);
or U3255 (N_3255,N_2644,N_2676);
or U3256 (N_3256,N_2519,N_2540);
and U3257 (N_3257,N_2806,N_2523);
nand U3258 (N_3258,N_2921,N_2538);
nand U3259 (N_3259,N_2769,N_2535);
nand U3260 (N_3260,N_2880,N_2724);
nor U3261 (N_3261,N_2713,N_2738);
and U3262 (N_3262,N_2922,N_2736);
nor U3263 (N_3263,N_2886,N_2981);
or U3264 (N_3264,N_2720,N_2731);
nand U3265 (N_3265,N_2999,N_2638);
nand U3266 (N_3266,N_2567,N_2693);
and U3267 (N_3267,N_2922,N_2564);
nor U3268 (N_3268,N_2791,N_2810);
and U3269 (N_3269,N_2618,N_2997);
nand U3270 (N_3270,N_2603,N_2824);
or U3271 (N_3271,N_2947,N_2629);
and U3272 (N_3272,N_2729,N_2947);
or U3273 (N_3273,N_2666,N_2718);
or U3274 (N_3274,N_2610,N_2537);
nand U3275 (N_3275,N_2741,N_2710);
or U3276 (N_3276,N_2517,N_2738);
nor U3277 (N_3277,N_2934,N_2542);
or U3278 (N_3278,N_2701,N_2578);
nand U3279 (N_3279,N_2912,N_2719);
nand U3280 (N_3280,N_2707,N_2732);
and U3281 (N_3281,N_2833,N_2587);
xnor U3282 (N_3282,N_2867,N_2871);
or U3283 (N_3283,N_2577,N_2757);
and U3284 (N_3284,N_2558,N_2661);
nand U3285 (N_3285,N_2994,N_2711);
nand U3286 (N_3286,N_2625,N_2647);
or U3287 (N_3287,N_2595,N_2683);
or U3288 (N_3288,N_2686,N_2674);
nor U3289 (N_3289,N_2776,N_2812);
nor U3290 (N_3290,N_2714,N_2666);
nand U3291 (N_3291,N_2636,N_2830);
nand U3292 (N_3292,N_2752,N_2639);
and U3293 (N_3293,N_2782,N_2664);
nand U3294 (N_3294,N_2626,N_2575);
and U3295 (N_3295,N_2678,N_2757);
nand U3296 (N_3296,N_2564,N_2819);
and U3297 (N_3297,N_2500,N_2853);
nor U3298 (N_3298,N_2867,N_2646);
or U3299 (N_3299,N_2985,N_2884);
nor U3300 (N_3300,N_2638,N_2570);
nor U3301 (N_3301,N_2541,N_2602);
and U3302 (N_3302,N_2956,N_2703);
or U3303 (N_3303,N_2621,N_2957);
xnor U3304 (N_3304,N_2778,N_2595);
xnor U3305 (N_3305,N_2919,N_2806);
or U3306 (N_3306,N_2527,N_2538);
xnor U3307 (N_3307,N_2955,N_2661);
nor U3308 (N_3308,N_2669,N_2874);
nand U3309 (N_3309,N_2709,N_2880);
nor U3310 (N_3310,N_2898,N_2849);
or U3311 (N_3311,N_2643,N_2645);
xor U3312 (N_3312,N_2643,N_2894);
and U3313 (N_3313,N_2975,N_2680);
nand U3314 (N_3314,N_2681,N_2643);
nand U3315 (N_3315,N_2967,N_2548);
and U3316 (N_3316,N_2785,N_2844);
and U3317 (N_3317,N_2749,N_2623);
and U3318 (N_3318,N_2568,N_2833);
nand U3319 (N_3319,N_2935,N_2929);
nor U3320 (N_3320,N_2949,N_2607);
and U3321 (N_3321,N_2856,N_2919);
nand U3322 (N_3322,N_2862,N_2800);
or U3323 (N_3323,N_2818,N_2990);
and U3324 (N_3324,N_2591,N_2931);
nand U3325 (N_3325,N_2510,N_2863);
nor U3326 (N_3326,N_2615,N_2735);
nand U3327 (N_3327,N_2649,N_2977);
nand U3328 (N_3328,N_2850,N_2829);
nand U3329 (N_3329,N_2508,N_2777);
or U3330 (N_3330,N_2732,N_2690);
or U3331 (N_3331,N_2826,N_2815);
nor U3332 (N_3332,N_2666,N_2747);
nor U3333 (N_3333,N_2553,N_2862);
or U3334 (N_3334,N_2989,N_2623);
and U3335 (N_3335,N_2764,N_2974);
and U3336 (N_3336,N_2885,N_2591);
xor U3337 (N_3337,N_2640,N_2560);
or U3338 (N_3338,N_2649,N_2880);
nand U3339 (N_3339,N_2555,N_2703);
nand U3340 (N_3340,N_2677,N_2762);
and U3341 (N_3341,N_2703,N_2671);
and U3342 (N_3342,N_2581,N_2781);
nor U3343 (N_3343,N_2520,N_2516);
nor U3344 (N_3344,N_2989,N_2927);
nand U3345 (N_3345,N_2563,N_2576);
nand U3346 (N_3346,N_2608,N_2605);
or U3347 (N_3347,N_2934,N_2870);
and U3348 (N_3348,N_2702,N_2911);
xnor U3349 (N_3349,N_2540,N_2929);
xor U3350 (N_3350,N_2693,N_2699);
nand U3351 (N_3351,N_2775,N_2670);
nor U3352 (N_3352,N_2607,N_2689);
or U3353 (N_3353,N_2573,N_2804);
nand U3354 (N_3354,N_2989,N_2890);
and U3355 (N_3355,N_2858,N_2667);
nor U3356 (N_3356,N_2880,N_2502);
and U3357 (N_3357,N_2617,N_2511);
xor U3358 (N_3358,N_2906,N_2776);
nand U3359 (N_3359,N_2843,N_2687);
or U3360 (N_3360,N_2856,N_2969);
and U3361 (N_3361,N_2726,N_2529);
and U3362 (N_3362,N_2863,N_2785);
or U3363 (N_3363,N_2776,N_2755);
xnor U3364 (N_3364,N_2614,N_2684);
nand U3365 (N_3365,N_2606,N_2541);
nor U3366 (N_3366,N_2806,N_2812);
nor U3367 (N_3367,N_2834,N_2569);
and U3368 (N_3368,N_2737,N_2733);
and U3369 (N_3369,N_2828,N_2853);
nor U3370 (N_3370,N_2747,N_2587);
nand U3371 (N_3371,N_2892,N_2907);
nand U3372 (N_3372,N_2719,N_2529);
or U3373 (N_3373,N_2823,N_2769);
nand U3374 (N_3374,N_2731,N_2817);
nand U3375 (N_3375,N_2901,N_2580);
and U3376 (N_3376,N_2663,N_2672);
or U3377 (N_3377,N_2931,N_2948);
and U3378 (N_3378,N_2900,N_2541);
or U3379 (N_3379,N_2646,N_2550);
and U3380 (N_3380,N_2972,N_2533);
nand U3381 (N_3381,N_2886,N_2687);
or U3382 (N_3382,N_2518,N_2657);
nand U3383 (N_3383,N_2902,N_2989);
nor U3384 (N_3384,N_2745,N_2821);
nor U3385 (N_3385,N_2945,N_2757);
xnor U3386 (N_3386,N_2882,N_2878);
nand U3387 (N_3387,N_2707,N_2690);
nor U3388 (N_3388,N_2698,N_2512);
nand U3389 (N_3389,N_2929,N_2988);
or U3390 (N_3390,N_2902,N_2558);
xnor U3391 (N_3391,N_2875,N_2513);
and U3392 (N_3392,N_2859,N_2824);
and U3393 (N_3393,N_2878,N_2962);
and U3394 (N_3394,N_2870,N_2697);
nand U3395 (N_3395,N_2629,N_2773);
or U3396 (N_3396,N_2986,N_2852);
nor U3397 (N_3397,N_2665,N_2637);
or U3398 (N_3398,N_2948,N_2776);
nand U3399 (N_3399,N_2749,N_2555);
and U3400 (N_3400,N_2771,N_2551);
nor U3401 (N_3401,N_2726,N_2505);
and U3402 (N_3402,N_2680,N_2789);
or U3403 (N_3403,N_2889,N_2764);
and U3404 (N_3404,N_2737,N_2517);
nor U3405 (N_3405,N_2739,N_2667);
or U3406 (N_3406,N_2830,N_2581);
xor U3407 (N_3407,N_2657,N_2504);
or U3408 (N_3408,N_2949,N_2565);
nand U3409 (N_3409,N_2505,N_2731);
nand U3410 (N_3410,N_2780,N_2579);
and U3411 (N_3411,N_2774,N_2912);
xor U3412 (N_3412,N_2620,N_2967);
nand U3413 (N_3413,N_2774,N_2734);
xor U3414 (N_3414,N_2894,N_2779);
nor U3415 (N_3415,N_2951,N_2598);
or U3416 (N_3416,N_2568,N_2694);
and U3417 (N_3417,N_2534,N_2550);
nand U3418 (N_3418,N_2507,N_2850);
nor U3419 (N_3419,N_2919,N_2594);
and U3420 (N_3420,N_2832,N_2939);
nand U3421 (N_3421,N_2701,N_2722);
or U3422 (N_3422,N_2577,N_2689);
and U3423 (N_3423,N_2808,N_2682);
and U3424 (N_3424,N_2961,N_2954);
or U3425 (N_3425,N_2552,N_2963);
or U3426 (N_3426,N_2589,N_2907);
nand U3427 (N_3427,N_2643,N_2620);
or U3428 (N_3428,N_2939,N_2907);
nand U3429 (N_3429,N_2738,N_2686);
nor U3430 (N_3430,N_2929,N_2541);
or U3431 (N_3431,N_2790,N_2528);
and U3432 (N_3432,N_2571,N_2510);
and U3433 (N_3433,N_2565,N_2576);
and U3434 (N_3434,N_2910,N_2554);
or U3435 (N_3435,N_2579,N_2688);
and U3436 (N_3436,N_2756,N_2812);
and U3437 (N_3437,N_2921,N_2704);
and U3438 (N_3438,N_2665,N_2851);
nand U3439 (N_3439,N_2761,N_2884);
nor U3440 (N_3440,N_2833,N_2856);
nand U3441 (N_3441,N_2935,N_2647);
or U3442 (N_3442,N_2808,N_2578);
or U3443 (N_3443,N_2946,N_2699);
nor U3444 (N_3444,N_2589,N_2657);
or U3445 (N_3445,N_2819,N_2615);
nor U3446 (N_3446,N_2747,N_2631);
and U3447 (N_3447,N_2713,N_2550);
nor U3448 (N_3448,N_2609,N_2947);
xnor U3449 (N_3449,N_2604,N_2572);
nand U3450 (N_3450,N_2770,N_2645);
or U3451 (N_3451,N_2939,N_2913);
nor U3452 (N_3452,N_2992,N_2980);
and U3453 (N_3453,N_2701,N_2695);
or U3454 (N_3454,N_2842,N_2873);
nor U3455 (N_3455,N_2522,N_2819);
and U3456 (N_3456,N_2601,N_2910);
or U3457 (N_3457,N_2669,N_2764);
nand U3458 (N_3458,N_2761,N_2680);
nor U3459 (N_3459,N_2755,N_2506);
nor U3460 (N_3460,N_2962,N_2889);
xnor U3461 (N_3461,N_2912,N_2862);
or U3462 (N_3462,N_2608,N_2954);
nand U3463 (N_3463,N_2955,N_2779);
nand U3464 (N_3464,N_2800,N_2576);
xor U3465 (N_3465,N_2881,N_2863);
xnor U3466 (N_3466,N_2781,N_2580);
xnor U3467 (N_3467,N_2822,N_2793);
nand U3468 (N_3468,N_2714,N_2621);
xnor U3469 (N_3469,N_2693,N_2566);
or U3470 (N_3470,N_2987,N_2506);
and U3471 (N_3471,N_2789,N_2572);
nor U3472 (N_3472,N_2896,N_2591);
xnor U3473 (N_3473,N_2675,N_2782);
and U3474 (N_3474,N_2520,N_2808);
or U3475 (N_3475,N_2671,N_2934);
nor U3476 (N_3476,N_2538,N_2827);
or U3477 (N_3477,N_2756,N_2750);
or U3478 (N_3478,N_2604,N_2748);
and U3479 (N_3479,N_2920,N_2766);
nand U3480 (N_3480,N_2973,N_2774);
and U3481 (N_3481,N_2509,N_2521);
nor U3482 (N_3482,N_2783,N_2914);
nor U3483 (N_3483,N_2536,N_2806);
nand U3484 (N_3484,N_2515,N_2564);
xnor U3485 (N_3485,N_2597,N_2899);
or U3486 (N_3486,N_2751,N_2833);
nand U3487 (N_3487,N_2694,N_2945);
or U3488 (N_3488,N_2732,N_2593);
nor U3489 (N_3489,N_2858,N_2756);
and U3490 (N_3490,N_2983,N_2984);
nor U3491 (N_3491,N_2791,N_2940);
or U3492 (N_3492,N_2784,N_2577);
or U3493 (N_3493,N_2622,N_2535);
nand U3494 (N_3494,N_2511,N_2746);
and U3495 (N_3495,N_2661,N_2580);
nor U3496 (N_3496,N_2649,N_2891);
nand U3497 (N_3497,N_2560,N_2521);
nor U3498 (N_3498,N_2886,N_2776);
nand U3499 (N_3499,N_2592,N_2767);
nand U3500 (N_3500,N_3263,N_3049);
nor U3501 (N_3501,N_3383,N_3408);
and U3502 (N_3502,N_3352,N_3468);
nand U3503 (N_3503,N_3216,N_3256);
nand U3504 (N_3504,N_3079,N_3211);
or U3505 (N_3505,N_3258,N_3285);
or U3506 (N_3506,N_3025,N_3172);
nand U3507 (N_3507,N_3117,N_3231);
or U3508 (N_3508,N_3370,N_3469);
nand U3509 (N_3509,N_3336,N_3186);
xor U3510 (N_3510,N_3323,N_3347);
or U3511 (N_3511,N_3277,N_3241);
or U3512 (N_3512,N_3297,N_3324);
or U3513 (N_3513,N_3445,N_3078);
nor U3514 (N_3514,N_3380,N_3162);
nand U3515 (N_3515,N_3213,N_3459);
nand U3516 (N_3516,N_3108,N_3421);
xor U3517 (N_3517,N_3464,N_3091);
or U3518 (N_3518,N_3032,N_3082);
or U3519 (N_3519,N_3354,N_3153);
xor U3520 (N_3520,N_3362,N_3453);
and U3521 (N_3521,N_3062,N_3406);
nand U3522 (N_3522,N_3447,N_3060);
nor U3523 (N_3523,N_3373,N_3010);
or U3524 (N_3524,N_3470,N_3425);
xnor U3525 (N_3525,N_3335,N_3145);
and U3526 (N_3526,N_3109,N_3189);
and U3527 (N_3527,N_3287,N_3157);
nor U3528 (N_3528,N_3332,N_3034);
and U3529 (N_3529,N_3257,N_3291);
nor U3530 (N_3530,N_3143,N_3279);
xnor U3531 (N_3531,N_3003,N_3321);
nand U3532 (N_3532,N_3286,N_3350);
or U3533 (N_3533,N_3466,N_3016);
nand U3534 (N_3534,N_3358,N_3181);
xnor U3535 (N_3535,N_3133,N_3377);
nand U3536 (N_3536,N_3372,N_3412);
xnor U3537 (N_3537,N_3471,N_3301);
or U3538 (N_3538,N_3110,N_3274);
or U3539 (N_3539,N_3012,N_3273);
or U3540 (N_3540,N_3473,N_3138);
or U3541 (N_3541,N_3268,N_3151);
nor U3542 (N_3542,N_3127,N_3044);
or U3543 (N_3543,N_3365,N_3340);
or U3544 (N_3544,N_3461,N_3167);
nand U3545 (N_3545,N_3289,N_3465);
nor U3546 (N_3546,N_3409,N_3064);
or U3547 (N_3547,N_3472,N_3485);
and U3548 (N_3548,N_3440,N_3233);
and U3549 (N_3549,N_3033,N_3306);
and U3550 (N_3550,N_3066,N_3477);
xnor U3551 (N_3551,N_3024,N_3148);
or U3552 (N_3552,N_3169,N_3232);
and U3553 (N_3553,N_3028,N_3396);
xor U3554 (N_3554,N_3042,N_3330);
nand U3555 (N_3555,N_3229,N_3441);
nand U3556 (N_3556,N_3410,N_3234);
and U3557 (N_3557,N_3249,N_3391);
and U3558 (N_3558,N_3367,N_3096);
nor U3559 (N_3559,N_3065,N_3077);
xnor U3560 (N_3560,N_3224,N_3009);
nor U3561 (N_3561,N_3221,N_3059);
or U3562 (N_3562,N_3013,N_3051);
nand U3563 (N_3563,N_3317,N_3192);
xnor U3564 (N_3564,N_3411,N_3008);
nor U3565 (N_3565,N_3443,N_3124);
and U3566 (N_3566,N_3021,N_3228);
nor U3567 (N_3567,N_3293,N_3270);
and U3568 (N_3568,N_3299,N_3206);
nor U3569 (N_3569,N_3191,N_3264);
nor U3570 (N_3570,N_3444,N_3111);
or U3571 (N_3571,N_3119,N_3305);
or U3572 (N_3572,N_3056,N_3045);
nor U3573 (N_3573,N_3495,N_3093);
xor U3574 (N_3574,N_3463,N_3161);
nor U3575 (N_3575,N_3276,N_3239);
or U3576 (N_3576,N_3415,N_3386);
or U3577 (N_3577,N_3460,N_3392);
xnor U3578 (N_3578,N_3399,N_3202);
nor U3579 (N_3579,N_3481,N_3403);
xnor U3580 (N_3580,N_3329,N_3075);
nor U3581 (N_3581,N_3413,N_3081);
xnor U3582 (N_3582,N_3176,N_3292);
nor U3583 (N_3583,N_3490,N_3338);
and U3584 (N_3584,N_3382,N_3307);
nor U3585 (N_3585,N_3251,N_3222);
or U3586 (N_3586,N_3300,N_3183);
or U3587 (N_3587,N_3499,N_3070);
nor U3588 (N_3588,N_3250,N_3462);
nor U3589 (N_3589,N_3026,N_3337);
or U3590 (N_3590,N_3437,N_3067);
nand U3591 (N_3591,N_3101,N_3043);
nand U3592 (N_3592,N_3493,N_3047);
and U3593 (N_3593,N_3318,N_3178);
nand U3594 (N_3594,N_3379,N_3141);
nor U3595 (N_3595,N_3435,N_3058);
or U3596 (N_3596,N_3416,N_3422);
nor U3597 (N_3597,N_3095,N_3227);
or U3598 (N_3598,N_3104,N_3209);
nor U3599 (N_3599,N_3004,N_3061);
nand U3600 (N_3600,N_3128,N_3255);
nand U3601 (N_3601,N_3381,N_3036);
nor U3602 (N_3602,N_3107,N_3375);
or U3603 (N_3603,N_3328,N_3195);
nor U3604 (N_3604,N_3269,N_3098);
or U3605 (N_3605,N_3099,N_3456);
nand U3606 (N_3606,N_3030,N_3219);
nor U3607 (N_3607,N_3105,N_3357);
nand U3608 (N_3608,N_3041,N_3387);
or U3609 (N_3609,N_3414,N_3121);
or U3610 (N_3610,N_3163,N_3245);
nor U3611 (N_3611,N_3368,N_3427);
and U3612 (N_3612,N_3244,N_3046);
or U3613 (N_3613,N_3311,N_3031);
or U3614 (N_3614,N_3247,N_3288);
nor U3615 (N_3615,N_3319,N_3184);
and U3616 (N_3616,N_3140,N_3334);
or U3617 (N_3617,N_3243,N_3130);
nand U3618 (N_3618,N_3165,N_3068);
nand U3619 (N_3619,N_3448,N_3089);
and U3620 (N_3620,N_3230,N_3074);
and U3621 (N_3621,N_3198,N_3146);
and U3622 (N_3622,N_3080,N_3439);
and U3623 (N_3623,N_3260,N_3149);
and U3624 (N_3624,N_3492,N_3309);
xor U3625 (N_3625,N_3226,N_3083);
nor U3626 (N_3626,N_3267,N_3103);
and U3627 (N_3627,N_3187,N_3147);
and U3628 (N_3628,N_3280,N_3112);
xor U3629 (N_3629,N_3316,N_3405);
nor U3630 (N_3630,N_3175,N_3160);
or U3631 (N_3631,N_3458,N_3038);
or U3632 (N_3632,N_3039,N_3424);
and U3633 (N_3633,N_3040,N_3100);
and U3634 (N_3634,N_3011,N_3142);
nand U3635 (N_3635,N_3423,N_3394);
nand U3636 (N_3636,N_3308,N_3407);
nand U3637 (N_3637,N_3005,N_3353);
and U3638 (N_3638,N_3237,N_3339);
nand U3639 (N_3639,N_3451,N_3125);
or U3640 (N_3640,N_3006,N_3310);
nand U3641 (N_3641,N_3428,N_3019);
xnor U3642 (N_3642,N_3196,N_3491);
or U3643 (N_3643,N_3356,N_3343);
nor U3644 (N_3644,N_3197,N_3348);
and U3645 (N_3645,N_3017,N_3238);
and U3646 (N_3646,N_3090,N_3304);
or U3647 (N_3647,N_3434,N_3055);
or U3648 (N_3648,N_3432,N_3205);
and U3649 (N_3649,N_3320,N_3092);
and U3650 (N_3650,N_3193,N_3361);
nor U3651 (N_3651,N_3253,N_3223);
nor U3652 (N_3652,N_3488,N_3217);
xor U3653 (N_3653,N_3312,N_3378);
nand U3654 (N_3654,N_3275,N_3053);
nor U3655 (N_3655,N_3129,N_3072);
nand U3656 (N_3656,N_3489,N_3155);
xor U3657 (N_3657,N_3054,N_3388);
nand U3658 (N_3658,N_3063,N_3097);
nand U3659 (N_3659,N_3159,N_3235);
nand U3660 (N_3660,N_3371,N_3050);
or U3661 (N_3661,N_3333,N_3262);
xnor U3662 (N_3662,N_3271,N_3120);
nor U3663 (N_3663,N_3171,N_3182);
nand U3664 (N_3664,N_3210,N_3020);
or U3665 (N_3665,N_3389,N_3442);
and U3666 (N_3666,N_3266,N_3457);
nor U3667 (N_3667,N_3190,N_3325);
nor U3668 (N_3668,N_3294,N_3179);
xor U3669 (N_3669,N_3152,N_3418);
and U3670 (N_3670,N_3154,N_3113);
and U3671 (N_3671,N_3430,N_3071);
nor U3672 (N_3672,N_3474,N_3131);
nand U3673 (N_3673,N_3076,N_3144);
nor U3674 (N_3674,N_3173,N_3484);
nand U3675 (N_3675,N_3327,N_3002);
and U3676 (N_3676,N_3214,N_3450);
and U3677 (N_3677,N_3174,N_3369);
nor U3678 (N_3678,N_3037,N_3207);
or U3679 (N_3679,N_3236,N_3482);
and U3680 (N_3680,N_3115,N_3073);
or U3681 (N_3681,N_3118,N_3326);
and U3682 (N_3682,N_3385,N_3242);
xnor U3683 (N_3683,N_3166,N_3139);
xnor U3684 (N_3684,N_3164,N_3436);
and U3685 (N_3685,N_3475,N_3454);
or U3686 (N_3686,N_3265,N_3027);
nand U3687 (N_3687,N_3342,N_3200);
nand U3688 (N_3688,N_3194,N_3252);
nand U3689 (N_3689,N_3479,N_3069);
nand U3690 (N_3690,N_3384,N_3498);
or U3691 (N_3691,N_3156,N_3106);
and U3692 (N_3692,N_3331,N_3126);
nand U3693 (N_3693,N_3259,N_3199);
and U3694 (N_3694,N_3086,N_3341);
and U3695 (N_3695,N_3283,N_3029);
xnor U3696 (N_3696,N_3303,N_3204);
or U3697 (N_3697,N_3346,N_3246);
and U3698 (N_3698,N_3429,N_3376);
nand U3699 (N_3699,N_3048,N_3446);
nor U3700 (N_3700,N_3170,N_3497);
nor U3701 (N_3701,N_3349,N_3000);
xor U3702 (N_3702,N_3296,N_3208);
nand U3703 (N_3703,N_3483,N_3278);
xor U3704 (N_3704,N_3018,N_3168);
and U3705 (N_3705,N_3359,N_3220);
nand U3706 (N_3706,N_3136,N_3360);
and U3707 (N_3707,N_3281,N_3203);
nand U3708 (N_3708,N_3322,N_3015);
or U3709 (N_3709,N_3158,N_3177);
or U3710 (N_3710,N_3272,N_3185);
nand U3711 (N_3711,N_3001,N_3390);
and U3712 (N_3712,N_3052,N_3035);
nor U3713 (N_3713,N_3134,N_3395);
and U3714 (N_3714,N_3426,N_3135);
nand U3715 (N_3715,N_3431,N_3023);
nand U3716 (N_3716,N_3188,N_3402);
nand U3717 (N_3717,N_3240,N_3397);
nor U3718 (N_3718,N_3433,N_3314);
and U3719 (N_3719,N_3302,N_3088);
xor U3720 (N_3720,N_3398,N_3022);
nand U3721 (N_3721,N_3212,N_3487);
nand U3722 (N_3722,N_3345,N_3467);
nand U3723 (N_3723,N_3123,N_3084);
and U3724 (N_3724,N_3225,N_3419);
nand U3725 (N_3725,N_3282,N_3085);
nor U3726 (N_3726,N_3417,N_3452);
and U3727 (N_3727,N_3298,N_3449);
nor U3728 (N_3728,N_3137,N_3315);
or U3729 (N_3729,N_3132,N_3496);
nand U3730 (N_3730,N_3364,N_3393);
xor U3731 (N_3731,N_3401,N_3438);
or U3732 (N_3732,N_3215,N_3400);
xor U3733 (N_3733,N_3180,N_3102);
or U3734 (N_3734,N_3248,N_3122);
or U3735 (N_3735,N_3116,N_3014);
nor U3736 (N_3736,N_3150,N_3094);
and U3737 (N_3737,N_3366,N_3057);
xor U3738 (N_3738,N_3404,N_3114);
nand U3739 (N_3739,N_3494,N_3313);
nand U3740 (N_3740,N_3344,N_3254);
nor U3741 (N_3741,N_3363,N_3351);
nand U3742 (N_3742,N_3374,N_3201);
nand U3743 (N_3743,N_3420,N_3295);
nor U3744 (N_3744,N_3486,N_3087);
nor U3745 (N_3745,N_3476,N_3480);
and U3746 (N_3746,N_3455,N_3218);
and U3747 (N_3747,N_3284,N_3261);
and U3748 (N_3748,N_3007,N_3355);
nand U3749 (N_3749,N_3290,N_3478);
nor U3750 (N_3750,N_3339,N_3086);
xor U3751 (N_3751,N_3110,N_3099);
nand U3752 (N_3752,N_3258,N_3064);
xnor U3753 (N_3753,N_3288,N_3299);
or U3754 (N_3754,N_3426,N_3493);
and U3755 (N_3755,N_3107,N_3404);
xor U3756 (N_3756,N_3497,N_3483);
and U3757 (N_3757,N_3213,N_3473);
xor U3758 (N_3758,N_3354,N_3364);
nor U3759 (N_3759,N_3133,N_3047);
or U3760 (N_3760,N_3195,N_3415);
xor U3761 (N_3761,N_3268,N_3022);
nand U3762 (N_3762,N_3458,N_3104);
nor U3763 (N_3763,N_3489,N_3095);
nand U3764 (N_3764,N_3470,N_3284);
and U3765 (N_3765,N_3485,N_3448);
nor U3766 (N_3766,N_3313,N_3260);
xor U3767 (N_3767,N_3434,N_3122);
xnor U3768 (N_3768,N_3068,N_3494);
nor U3769 (N_3769,N_3172,N_3141);
and U3770 (N_3770,N_3182,N_3169);
nor U3771 (N_3771,N_3111,N_3283);
nor U3772 (N_3772,N_3320,N_3109);
nand U3773 (N_3773,N_3117,N_3056);
xnor U3774 (N_3774,N_3197,N_3193);
nor U3775 (N_3775,N_3020,N_3025);
nand U3776 (N_3776,N_3495,N_3390);
nor U3777 (N_3777,N_3222,N_3439);
and U3778 (N_3778,N_3480,N_3233);
nor U3779 (N_3779,N_3250,N_3007);
or U3780 (N_3780,N_3048,N_3164);
nand U3781 (N_3781,N_3453,N_3319);
and U3782 (N_3782,N_3450,N_3286);
or U3783 (N_3783,N_3260,N_3494);
and U3784 (N_3784,N_3400,N_3136);
nand U3785 (N_3785,N_3034,N_3347);
nand U3786 (N_3786,N_3078,N_3123);
or U3787 (N_3787,N_3480,N_3206);
nor U3788 (N_3788,N_3174,N_3054);
nor U3789 (N_3789,N_3058,N_3137);
and U3790 (N_3790,N_3103,N_3371);
nand U3791 (N_3791,N_3295,N_3256);
or U3792 (N_3792,N_3498,N_3422);
nand U3793 (N_3793,N_3076,N_3249);
or U3794 (N_3794,N_3102,N_3232);
and U3795 (N_3795,N_3153,N_3008);
xor U3796 (N_3796,N_3470,N_3041);
nand U3797 (N_3797,N_3385,N_3150);
and U3798 (N_3798,N_3152,N_3434);
nand U3799 (N_3799,N_3078,N_3263);
or U3800 (N_3800,N_3351,N_3109);
and U3801 (N_3801,N_3210,N_3300);
nand U3802 (N_3802,N_3106,N_3117);
or U3803 (N_3803,N_3398,N_3154);
xnor U3804 (N_3804,N_3052,N_3144);
and U3805 (N_3805,N_3272,N_3436);
nor U3806 (N_3806,N_3487,N_3243);
nor U3807 (N_3807,N_3406,N_3034);
xor U3808 (N_3808,N_3365,N_3359);
xor U3809 (N_3809,N_3403,N_3061);
nand U3810 (N_3810,N_3333,N_3447);
nand U3811 (N_3811,N_3076,N_3200);
xnor U3812 (N_3812,N_3471,N_3134);
or U3813 (N_3813,N_3277,N_3002);
xor U3814 (N_3814,N_3272,N_3190);
xnor U3815 (N_3815,N_3459,N_3482);
nand U3816 (N_3816,N_3325,N_3473);
nor U3817 (N_3817,N_3443,N_3007);
and U3818 (N_3818,N_3045,N_3488);
xnor U3819 (N_3819,N_3331,N_3452);
nand U3820 (N_3820,N_3419,N_3145);
nor U3821 (N_3821,N_3131,N_3418);
nand U3822 (N_3822,N_3168,N_3488);
nand U3823 (N_3823,N_3496,N_3176);
or U3824 (N_3824,N_3300,N_3366);
or U3825 (N_3825,N_3396,N_3184);
nand U3826 (N_3826,N_3385,N_3180);
nor U3827 (N_3827,N_3393,N_3434);
nor U3828 (N_3828,N_3440,N_3305);
or U3829 (N_3829,N_3159,N_3014);
and U3830 (N_3830,N_3014,N_3418);
or U3831 (N_3831,N_3001,N_3244);
nand U3832 (N_3832,N_3196,N_3173);
and U3833 (N_3833,N_3187,N_3366);
nand U3834 (N_3834,N_3178,N_3208);
xnor U3835 (N_3835,N_3210,N_3457);
nand U3836 (N_3836,N_3428,N_3093);
xor U3837 (N_3837,N_3271,N_3071);
and U3838 (N_3838,N_3129,N_3226);
or U3839 (N_3839,N_3316,N_3268);
and U3840 (N_3840,N_3488,N_3055);
and U3841 (N_3841,N_3116,N_3312);
or U3842 (N_3842,N_3486,N_3479);
nand U3843 (N_3843,N_3271,N_3446);
and U3844 (N_3844,N_3003,N_3481);
or U3845 (N_3845,N_3333,N_3437);
or U3846 (N_3846,N_3369,N_3412);
nor U3847 (N_3847,N_3242,N_3317);
and U3848 (N_3848,N_3089,N_3487);
and U3849 (N_3849,N_3009,N_3356);
and U3850 (N_3850,N_3476,N_3035);
or U3851 (N_3851,N_3176,N_3219);
nand U3852 (N_3852,N_3086,N_3106);
nor U3853 (N_3853,N_3293,N_3235);
nor U3854 (N_3854,N_3423,N_3059);
nor U3855 (N_3855,N_3492,N_3119);
xor U3856 (N_3856,N_3340,N_3081);
nand U3857 (N_3857,N_3340,N_3229);
nand U3858 (N_3858,N_3492,N_3481);
and U3859 (N_3859,N_3274,N_3327);
and U3860 (N_3860,N_3138,N_3285);
and U3861 (N_3861,N_3246,N_3394);
nor U3862 (N_3862,N_3186,N_3195);
nand U3863 (N_3863,N_3467,N_3476);
or U3864 (N_3864,N_3083,N_3201);
and U3865 (N_3865,N_3434,N_3454);
or U3866 (N_3866,N_3038,N_3343);
and U3867 (N_3867,N_3064,N_3084);
or U3868 (N_3868,N_3227,N_3124);
or U3869 (N_3869,N_3466,N_3399);
nor U3870 (N_3870,N_3318,N_3428);
nor U3871 (N_3871,N_3372,N_3122);
or U3872 (N_3872,N_3187,N_3468);
or U3873 (N_3873,N_3424,N_3239);
nand U3874 (N_3874,N_3488,N_3334);
or U3875 (N_3875,N_3123,N_3488);
nor U3876 (N_3876,N_3471,N_3366);
nor U3877 (N_3877,N_3011,N_3282);
xor U3878 (N_3878,N_3364,N_3055);
and U3879 (N_3879,N_3434,N_3284);
nor U3880 (N_3880,N_3460,N_3405);
nand U3881 (N_3881,N_3289,N_3215);
or U3882 (N_3882,N_3110,N_3148);
nor U3883 (N_3883,N_3169,N_3427);
or U3884 (N_3884,N_3013,N_3400);
and U3885 (N_3885,N_3492,N_3144);
or U3886 (N_3886,N_3457,N_3075);
and U3887 (N_3887,N_3162,N_3272);
and U3888 (N_3888,N_3391,N_3238);
nand U3889 (N_3889,N_3475,N_3391);
or U3890 (N_3890,N_3004,N_3226);
nor U3891 (N_3891,N_3283,N_3085);
xnor U3892 (N_3892,N_3444,N_3498);
xnor U3893 (N_3893,N_3265,N_3128);
and U3894 (N_3894,N_3191,N_3334);
or U3895 (N_3895,N_3050,N_3002);
nand U3896 (N_3896,N_3167,N_3296);
nand U3897 (N_3897,N_3358,N_3144);
nor U3898 (N_3898,N_3222,N_3116);
and U3899 (N_3899,N_3021,N_3285);
nand U3900 (N_3900,N_3112,N_3428);
nor U3901 (N_3901,N_3264,N_3132);
or U3902 (N_3902,N_3492,N_3134);
and U3903 (N_3903,N_3427,N_3025);
nand U3904 (N_3904,N_3122,N_3343);
or U3905 (N_3905,N_3246,N_3050);
and U3906 (N_3906,N_3054,N_3119);
and U3907 (N_3907,N_3220,N_3270);
or U3908 (N_3908,N_3340,N_3079);
nand U3909 (N_3909,N_3183,N_3012);
nor U3910 (N_3910,N_3321,N_3033);
or U3911 (N_3911,N_3102,N_3366);
and U3912 (N_3912,N_3498,N_3379);
nor U3913 (N_3913,N_3254,N_3459);
nor U3914 (N_3914,N_3429,N_3280);
or U3915 (N_3915,N_3233,N_3365);
nand U3916 (N_3916,N_3138,N_3466);
nor U3917 (N_3917,N_3170,N_3081);
nand U3918 (N_3918,N_3493,N_3277);
nand U3919 (N_3919,N_3003,N_3049);
nor U3920 (N_3920,N_3214,N_3384);
nand U3921 (N_3921,N_3343,N_3059);
or U3922 (N_3922,N_3419,N_3182);
nor U3923 (N_3923,N_3274,N_3445);
nand U3924 (N_3924,N_3308,N_3394);
nor U3925 (N_3925,N_3034,N_3076);
nand U3926 (N_3926,N_3186,N_3434);
or U3927 (N_3927,N_3143,N_3334);
nand U3928 (N_3928,N_3471,N_3433);
and U3929 (N_3929,N_3236,N_3248);
nor U3930 (N_3930,N_3026,N_3148);
or U3931 (N_3931,N_3160,N_3010);
and U3932 (N_3932,N_3038,N_3477);
xor U3933 (N_3933,N_3215,N_3207);
or U3934 (N_3934,N_3450,N_3014);
nor U3935 (N_3935,N_3191,N_3422);
nor U3936 (N_3936,N_3182,N_3272);
nand U3937 (N_3937,N_3219,N_3121);
and U3938 (N_3938,N_3161,N_3334);
or U3939 (N_3939,N_3290,N_3140);
nor U3940 (N_3940,N_3387,N_3281);
xnor U3941 (N_3941,N_3478,N_3226);
and U3942 (N_3942,N_3184,N_3121);
nand U3943 (N_3943,N_3332,N_3423);
nor U3944 (N_3944,N_3275,N_3081);
nand U3945 (N_3945,N_3244,N_3335);
nand U3946 (N_3946,N_3275,N_3400);
or U3947 (N_3947,N_3479,N_3168);
and U3948 (N_3948,N_3247,N_3150);
and U3949 (N_3949,N_3417,N_3224);
or U3950 (N_3950,N_3135,N_3277);
or U3951 (N_3951,N_3369,N_3051);
nand U3952 (N_3952,N_3398,N_3492);
and U3953 (N_3953,N_3045,N_3286);
or U3954 (N_3954,N_3213,N_3257);
xor U3955 (N_3955,N_3048,N_3440);
nor U3956 (N_3956,N_3008,N_3129);
or U3957 (N_3957,N_3103,N_3250);
or U3958 (N_3958,N_3307,N_3254);
xor U3959 (N_3959,N_3017,N_3133);
nand U3960 (N_3960,N_3459,N_3139);
nand U3961 (N_3961,N_3013,N_3425);
nor U3962 (N_3962,N_3469,N_3094);
or U3963 (N_3963,N_3495,N_3160);
or U3964 (N_3964,N_3414,N_3471);
or U3965 (N_3965,N_3497,N_3340);
nor U3966 (N_3966,N_3052,N_3449);
nand U3967 (N_3967,N_3152,N_3300);
xor U3968 (N_3968,N_3260,N_3069);
or U3969 (N_3969,N_3309,N_3073);
or U3970 (N_3970,N_3007,N_3482);
or U3971 (N_3971,N_3097,N_3407);
and U3972 (N_3972,N_3220,N_3461);
nor U3973 (N_3973,N_3115,N_3011);
nand U3974 (N_3974,N_3461,N_3208);
xnor U3975 (N_3975,N_3029,N_3115);
and U3976 (N_3976,N_3420,N_3284);
xnor U3977 (N_3977,N_3313,N_3438);
nand U3978 (N_3978,N_3090,N_3297);
or U3979 (N_3979,N_3052,N_3475);
xnor U3980 (N_3980,N_3208,N_3126);
nor U3981 (N_3981,N_3392,N_3182);
or U3982 (N_3982,N_3149,N_3306);
xor U3983 (N_3983,N_3128,N_3359);
nor U3984 (N_3984,N_3270,N_3450);
nor U3985 (N_3985,N_3196,N_3008);
nor U3986 (N_3986,N_3065,N_3097);
or U3987 (N_3987,N_3499,N_3469);
nor U3988 (N_3988,N_3307,N_3000);
nor U3989 (N_3989,N_3484,N_3250);
nand U3990 (N_3990,N_3255,N_3239);
nand U3991 (N_3991,N_3336,N_3349);
xnor U3992 (N_3992,N_3021,N_3259);
nor U3993 (N_3993,N_3079,N_3422);
nand U3994 (N_3994,N_3122,N_3358);
xor U3995 (N_3995,N_3319,N_3294);
nand U3996 (N_3996,N_3256,N_3073);
or U3997 (N_3997,N_3488,N_3304);
nor U3998 (N_3998,N_3038,N_3445);
and U3999 (N_3999,N_3387,N_3411);
nand U4000 (N_4000,N_3791,N_3807);
nor U4001 (N_4001,N_3922,N_3947);
nor U4002 (N_4002,N_3795,N_3908);
and U4003 (N_4003,N_3659,N_3620);
nand U4004 (N_4004,N_3631,N_3966);
and U4005 (N_4005,N_3579,N_3646);
nand U4006 (N_4006,N_3600,N_3906);
or U4007 (N_4007,N_3762,N_3825);
xnor U4008 (N_4008,N_3777,N_3633);
or U4009 (N_4009,N_3813,N_3712);
and U4010 (N_4010,N_3532,N_3604);
or U4011 (N_4011,N_3970,N_3953);
or U4012 (N_4012,N_3786,N_3982);
nor U4013 (N_4013,N_3874,N_3591);
and U4014 (N_4014,N_3886,N_3958);
and U4015 (N_4015,N_3590,N_3548);
and U4016 (N_4016,N_3747,N_3972);
or U4017 (N_4017,N_3519,N_3632);
nand U4018 (N_4018,N_3715,N_3944);
and U4019 (N_4019,N_3510,N_3509);
or U4020 (N_4020,N_3834,N_3885);
nor U4021 (N_4021,N_3962,N_3597);
xnor U4022 (N_4022,N_3576,N_3569);
nor U4023 (N_4023,N_3746,N_3948);
nand U4024 (N_4024,N_3860,N_3657);
nor U4025 (N_4025,N_3960,N_3702);
nor U4026 (N_4026,N_3552,N_3687);
and U4027 (N_4027,N_3606,N_3835);
nand U4028 (N_4028,N_3816,N_3545);
and U4029 (N_4029,N_3826,N_3580);
nand U4030 (N_4030,N_3800,N_3678);
nand U4031 (N_4031,N_3768,N_3693);
or U4032 (N_4032,N_3821,N_3751);
nand U4033 (N_4033,N_3806,N_3793);
xnor U4034 (N_4034,N_3598,N_3555);
or U4035 (N_4035,N_3901,N_3750);
nand U4036 (N_4036,N_3538,N_3518);
nand U4037 (N_4037,N_3973,N_3849);
nand U4038 (N_4038,N_3898,N_3823);
and U4039 (N_4039,N_3796,N_3686);
nor U4040 (N_4040,N_3998,N_3797);
and U4041 (N_4041,N_3773,N_3771);
or U4042 (N_4042,N_3879,N_3649);
nor U4043 (N_4043,N_3848,N_3924);
and U4044 (N_4044,N_3938,N_3524);
and U4045 (N_4045,N_3596,N_3805);
and U4046 (N_4046,N_3918,N_3820);
or U4047 (N_4047,N_3933,N_3581);
or U4048 (N_4048,N_3977,N_3881);
nand U4049 (N_4049,N_3640,N_3586);
or U4050 (N_4050,N_3585,N_3584);
nor U4051 (N_4051,N_3997,N_3913);
nor U4052 (N_4052,N_3971,N_3957);
xnor U4053 (N_4053,N_3529,N_3949);
nand U4054 (N_4054,N_3843,N_3900);
nor U4055 (N_4055,N_3814,N_3878);
nand U4056 (N_4056,N_3551,N_3740);
and U4057 (N_4057,N_3688,N_3719);
or U4058 (N_4058,N_3671,N_3999);
or U4059 (N_4059,N_3903,N_3703);
and U4060 (N_4060,N_3954,N_3699);
and U4061 (N_4061,N_3522,N_3929);
nand U4062 (N_4062,N_3931,N_3838);
nand U4063 (N_4063,N_3701,N_3996);
xnor U4064 (N_4064,N_3945,N_3742);
and U4065 (N_4065,N_3883,N_3562);
or U4066 (N_4066,N_3675,N_3912);
and U4067 (N_4067,N_3840,N_3790);
or U4068 (N_4068,N_3910,N_3622);
and U4069 (N_4069,N_3905,N_3560);
and U4070 (N_4070,N_3717,N_3914);
nand U4071 (N_4071,N_3547,N_3575);
nor U4072 (N_4072,N_3978,N_3639);
and U4073 (N_4073,N_3753,N_3828);
nand U4074 (N_4074,N_3617,N_3810);
and U4075 (N_4075,N_3526,N_3549);
nand U4076 (N_4076,N_3844,N_3644);
nand U4077 (N_4077,N_3691,N_3680);
nand U4078 (N_4078,N_3963,N_3694);
nor U4079 (N_4079,N_3899,N_3511);
nand U4080 (N_4080,N_3544,N_3809);
nand U4081 (N_4081,N_3818,N_3634);
and U4082 (N_4082,N_3515,N_3781);
nand U4083 (N_4083,N_3616,N_3779);
and U4084 (N_4084,N_3625,N_3561);
and U4085 (N_4085,N_3830,N_3984);
nor U4086 (N_4086,N_3605,N_3744);
nor U4087 (N_4087,N_3643,N_3799);
and U4088 (N_4088,N_3660,N_3683);
nand U4089 (N_4089,N_3917,N_3767);
xnor U4090 (N_4090,N_3697,N_3578);
nor U4091 (N_4091,N_3871,N_3864);
nor U4092 (N_4092,N_3872,N_3558);
nor U4093 (N_4093,N_3556,N_3761);
or U4094 (N_4094,N_3819,N_3685);
nor U4095 (N_4095,N_3775,N_3690);
nor U4096 (N_4096,N_3695,N_3884);
and U4097 (N_4097,N_3500,N_3845);
nor U4098 (N_4098,N_3629,N_3939);
nand U4099 (N_4099,N_3772,N_3647);
and U4100 (N_4100,N_3974,N_3850);
and U4101 (N_4101,N_3778,N_3855);
or U4102 (N_4102,N_3756,N_3943);
and U4103 (N_4103,N_3749,N_3537);
nor U4104 (N_4104,N_3921,N_3983);
and U4105 (N_4105,N_3927,N_3714);
and U4106 (N_4106,N_3904,N_3967);
or U4107 (N_4107,N_3593,N_3546);
xor U4108 (N_4108,N_3655,N_3706);
or U4109 (N_4109,N_3987,N_3776);
nor U4110 (N_4110,N_3928,N_3567);
and U4111 (N_4111,N_3663,N_3780);
nor U4112 (N_4112,N_3824,N_3641);
or U4113 (N_4113,N_3648,N_3976);
nor U4114 (N_4114,N_3990,N_3618);
nand U4115 (N_4115,N_3504,N_3950);
or U4116 (N_4116,N_3802,N_3923);
and U4117 (N_4117,N_3669,N_3677);
nand U4118 (N_4118,N_3572,N_3915);
or U4119 (N_4119,N_3527,N_3888);
xor U4120 (N_4120,N_3539,N_3863);
nand U4121 (N_4121,N_3925,N_3969);
or U4122 (N_4122,N_3865,N_3523);
nor U4123 (N_4123,N_3952,N_3782);
nor U4124 (N_4124,N_3568,N_3979);
nor U4125 (N_4125,N_3731,N_3808);
and U4126 (N_4126,N_3839,N_3512);
and U4127 (N_4127,N_3672,N_3829);
nor U4128 (N_4128,N_3501,N_3517);
nand U4129 (N_4129,N_3533,N_3670);
nor U4130 (N_4130,N_3946,N_3866);
or U4131 (N_4131,N_3896,N_3728);
or U4132 (N_4132,N_3566,N_3877);
and U4133 (N_4133,N_3557,N_3891);
or U4134 (N_4134,N_3815,N_3563);
nor U4135 (N_4135,N_3602,N_3801);
nor U4136 (N_4136,N_3530,N_3592);
nor U4137 (N_4137,N_3986,N_3708);
and U4138 (N_4138,N_3736,N_3705);
nor U4139 (N_4139,N_3502,N_3769);
xor U4140 (N_4140,N_3964,N_3737);
or U4141 (N_4141,N_3540,N_3867);
and U4142 (N_4142,N_3862,N_3599);
and U4143 (N_4143,N_3991,N_3892);
xnor U4144 (N_4144,N_3889,N_3609);
and U4145 (N_4145,N_3926,N_3763);
or U4146 (N_4146,N_3794,N_3774);
nand U4147 (N_4147,N_3822,N_3505);
nor U4148 (N_4148,N_3851,N_3857);
and U4149 (N_4149,N_3937,N_3506);
nand U4150 (N_4150,N_3650,N_3528);
or U4151 (N_4151,N_3662,N_3738);
or U4152 (N_4152,N_3890,N_3789);
nand U4153 (N_4153,N_3985,N_3536);
and U4154 (N_4154,N_3610,N_3729);
nor U4155 (N_4155,N_3748,N_3674);
and U4156 (N_4156,N_3992,N_3621);
nor U4157 (N_4157,N_3619,N_3804);
and U4158 (N_4158,N_3847,N_3932);
nand U4159 (N_4159,N_3732,N_3909);
nor U4160 (N_4160,N_3995,N_3817);
nand U4161 (N_4161,N_3870,N_3920);
or U4162 (N_4162,N_3652,N_3711);
or U4163 (N_4163,N_3770,N_3836);
nand U4164 (N_4164,N_3955,N_3897);
and U4165 (N_4165,N_3503,N_3664);
nor U4166 (N_4166,N_3521,N_3696);
and U4167 (N_4167,N_3853,N_3868);
and U4168 (N_4168,N_3713,N_3667);
nor U4169 (N_4169,N_3676,N_3707);
nand U4170 (N_4170,N_3934,N_3757);
nor U4171 (N_4171,N_3535,N_3607);
and U4172 (N_4172,N_3859,N_3792);
nand U4173 (N_4173,N_3842,N_3832);
nand U4174 (N_4174,N_3612,N_3959);
nor U4175 (N_4175,N_3559,N_3887);
or U4176 (N_4176,N_3666,N_3827);
xor U4177 (N_4177,N_3726,N_3743);
nor U4178 (N_4178,N_3722,N_3550);
or U4179 (N_4179,N_3710,N_3873);
nand U4180 (N_4180,N_3811,N_3930);
xor U4181 (N_4181,N_3601,N_3727);
nand U4182 (N_4182,N_3583,N_3759);
nand U4183 (N_4183,N_3852,N_3733);
nor U4184 (N_4184,N_3785,N_3681);
xor U4185 (N_4185,N_3783,N_3615);
and U4186 (N_4186,N_3841,N_3542);
and U4187 (N_4187,N_3554,N_3725);
xnor U4188 (N_4188,N_3833,N_3624);
nand U4189 (N_4189,N_3875,N_3916);
nand U4190 (N_4190,N_3935,N_3961);
and U4191 (N_4191,N_3638,N_3981);
or U4192 (N_4192,N_3894,N_3658);
and U4193 (N_4193,N_3942,N_3861);
nor U4194 (N_4194,N_3764,N_3895);
and U4195 (N_4195,N_3661,N_3788);
and U4196 (N_4196,N_3752,N_3721);
nand U4197 (N_4197,N_3936,N_3831);
nor U4198 (N_4198,N_3692,N_3543);
or U4199 (N_4199,N_3513,N_3516);
xnor U4200 (N_4200,N_3541,N_3635);
nor U4201 (N_4201,N_3668,N_3653);
nor U4202 (N_4202,N_3758,N_3654);
or U4203 (N_4203,N_3595,N_3812);
nor U4204 (N_4204,N_3739,N_3755);
nand U4205 (N_4205,N_3594,N_3956);
and U4206 (N_4206,N_3988,N_3698);
nand U4207 (N_4207,N_3893,N_3628);
and U4208 (N_4208,N_3951,N_3627);
nand U4209 (N_4209,N_3614,N_3574);
nand U4210 (N_4210,N_3637,N_3760);
nand U4211 (N_4211,N_3684,N_3798);
xnor U4212 (N_4212,N_3704,N_3507);
nor U4213 (N_4213,N_3534,N_3784);
xor U4214 (N_4214,N_3837,N_3919);
nor U4215 (N_4215,N_3745,N_3673);
or U4216 (N_4216,N_3630,N_3709);
or U4217 (N_4217,N_3608,N_3882);
nand U4218 (N_4218,N_3968,N_3626);
nor U4219 (N_4219,N_3803,N_3907);
nor U4220 (N_4220,N_3980,N_3553);
nor U4221 (N_4221,N_3754,N_3645);
nand U4222 (N_4222,N_3573,N_3724);
nand U4223 (N_4223,N_3514,N_3989);
xnor U4224 (N_4224,N_3577,N_3623);
nor U4225 (N_4225,N_3734,N_3582);
xnor U4226 (N_4226,N_3651,N_3603);
or U4227 (N_4227,N_3718,N_3656);
or U4228 (N_4228,N_3911,N_3720);
nand U4229 (N_4229,N_3587,N_3858);
nand U4230 (N_4230,N_3508,N_3570);
and U4231 (N_4231,N_3846,N_3588);
nor U4232 (N_4232,N_3741,N_3902);
or U4233 (N_4233,N_3876,N_3679);
nor U4234 (N_4234,N_3765,N_3941);
and U4235 (N_4235,N_3880,N_3940);
nor U4236 (N_4236,N_3689,N_3723);
nor U4237 (N_4237,N_3571,N_3965);
or U4238 (N_4238,N_3564,N_3665);
xor U4239 (N_4239,N_3531,N_3611);
nand U4240 (N_4240,N_3869,N_3716);
and U4241 (N_4241,N_3766,N_3735);
nand U4242 (N_4242,N_3854,N_3525);
nor U4243 (N_4243,N_3642,N_3993);
or U4244 (N_4244,N_3636,N_3613);
nor U4245 (N_4245,N_3700,N_3730);
nand U4246 (N_4246,N_3975,N_3994);
nand U4247 (N_4247,N_3520,N_3565);
nor U4248 (N_4248,N_3787,N_3589);
or U4249 (N_4249,N_3682,N_3856);
or U4250 (N_4250,N_3627,N_3892);
nor U4251 (N_4251,N_3876,N_3643);
or U4252 (N_4252,N_3991,N_3905);
nand U4253 (N_4253,N_3682,N_3701);
or U4254 (N_4254,N_3518,N_3818);
and U4255 (N_4255,N_3724,N_3515);
xor U4256 (N_4256,N_3638,N_3622);
nand U4257 (N_4257,N_3855,N_3766);
and U4258 (N_4258,N_3574,N_3780);
nand U4259 (N_4259,N_3723,N_3757);
xnor U4260 (N_4260,N_3896,N_3890);
and U4261 (N_4261,N_3786,N_3750);
nor U4262 (N_4262,N_3806,N_3617);
and U4263 (N_4263,N_3872,N_3504);
nor U4264 (N_4264,N_3942,N_3576);
nor U4265 (N_4265,N_3994,N_3703);
nor U4266 (N_4266,N_3591,N_3670);
nand U4267 (N_4267,N_3961,N_3665);
or U4268 (N_4268,N_3538,N_3895);
or U4269 (N_4269,N_3678,N_3743);
or U4270 (N_4270,N_3510,N_3711);
xor U4271 (N_4271,N_3833,N_3844);
nor U4272 (N_4272,N_3571,N_3925);
nand U4273 (N_4273,N_3746,N_3808);
or U4274 (N_4274,N_3686,N_3884);
and U4275 (N_4275,N_3651,N_3983);
nor U4276 (N_4276,N_3612,N_3939);
nand U4277 (N_4277,N_3598,N_3880);
and U4278 (N_4278,N_3656,N_3784);
or U4279 (N_4279,N_3800,N_3506);
nor U4280 (N_4280,N_3794,N_3887);
nand U4281 (N_4281,N_3811,N_3588);
or U4282 (N_4282,N_3895,N_3661);
nor U4283 (N_4283,N_3937,N_3901);
nand U4284 (N_4284,N_3515,N_3647);
nor U4285 (N_4285,N_3698,N_3986);
and U4286 (N_4286,N_3550,N_3829);
and U4287 (N_4287,N_3922,N_3891);
or U4288 (N_4288,N_3701,N_3951);
or U4289 (N_4289,N_3866,N_3740);
nand U4290 (N_4290,N_3931,N_3614);
and U4291 (N_4291,N_3579,N_3738);
nand U4292 (N_4292,N_3643,N_3576);
and U4293 (N_4293,N_3815,N_3611);
nand U4294 (N_4294,N_3504,N_3730);
or U4295 (N_4295,N_3779,N_3531);
nand U4296 (N_4296,N_3722,N_3825);
nor U4297 (N_4297,N_3940,N_3881);
nor U4298 (N_4298,N_3909,N_3629);
or U4299 (N_4299,N_3690,N_3864);
nand U4300 (N_4300,N_3991,N_3664);
nand U4301 (N_4301,N_3639,N_3973);
and U4302 (N_4302,N_3880,N_3586);
or U4303 (N_4303,N_3959,N_3942);
or U4304 (N_4304,N_3904,N_3885);
and U4305 (N_4305,N_3900,N_3789);
or U4306 (N_4306,N_3823,N_3899);
or U4307 (N_4307,N_3796,N_3842);
or U4308 (N_4308,N_3959,N_3590);
nor U4309 (N_4309,N_3942,N_3845);
and U4310 (N_4310,N_3518,N_3579);
nand U4311 (N_4311,N_3850,N_3549);
or U4312 (N_4312,N_3872,N_3879);
nand U4313 (N_4313,N_3821,N_3927);
or U4314 (N_4314,N_3543,N_3596);
and U4315 (N_4315,N_3875,N_3781);
nor U4316 (N_4316,N_3548,N_3871);
nand U4317 (N_4317,N_3578,N_3757);
and U4318 (N_4318,N_3993,N_3894);
nand U4319 (N_4319,N_3927,N_3684);
or U4320 (N_4320,N_3779,N_3795);
nor U4321 (N_4321,N_3654,N_3608);
or U4322 (N_4322,N_3611,N_3955);
or U4323 (N_4323,N_3766,N_3597);
and U4324 (N_4324,N_3503,N_3640);
and U4325 (N_4325,N_3982,N_3679);
and U4326 (N_4326,N_3592,N_3622);
or U4327 (N_4327,N_3659,N_3799);
nand U4328 (N_4328,N_3987,N_3656);
or U4329 (N_4329,N_3576,N_3608);
nor U4330 (N_4330,N_3825,N_3513);
or U4331 (N_4331,N_3730,N_3627);
xor U4332 (N_4332,N_3564,N_3538);
nor U4333 (N_4333,N_3903,N_3881);
nand U4334 (N_4334,N_3636,N_3801);
nand U4335 (N_4335,N_3748,N_3571);
nand U4336 (N_4336,N_3541,N_3766);
nand U4337 (N_4337,N_3908,N_3821);
nand U4338 (N_4338,N_3799,N_3613);
nor U4339 (N_4339,N_3794,N_3583);
or U4340 (N_4340,N_3721,N_3975);
or U4341 (N_4341,N_3870,N_3633);
nand U4342 (N_4342,N_3584,N_3647);
and U4343 (N_4343,N_3589,N_3687);
and U4344 (N_4344,N_3602,N_3819);
nand U4345 (N_4345,N_3815,N_3763);
nand U4346 (N_4346,N_3592,N_3809);
nor U4347 (N_4347,N_3645,N_3950);
nand U4348 (N_4348,N_3658,N_3910);
nand U4349 (N_4349,N_3520,N_3668);
nor U4350 (N_4350,N_3905,N_3939);
xnor U4351 (N_4351,N_3505,N_3557);
and U4352 (N_4352,N_3978,N_3804);
nor U4353 (N_4353,N_3917,N_3795);
nor U4354 (N_4354,N_3773,N_3920);
nor U4355 (N_4355,N_3851,N_3825);
nand U4356 (N_4356,N_3526,N_3788);
or U4357 (N_4357,N_3893,N_3539);
nand U4358 (N_4358,N_3850,N_3940);
or U4359 (N_4359,N_3734,N_3752);
nor U4360 (N_4360,N_3508,N_3819);
nor U4361 (N_4361,N_3502,N_3645);
and U4362 (N_4362,N_3526,N_3957);
nor U4363 (N_4363,N_3887,N_3688);
nand U4364 (N_4364,N_3797,N_3518);
nor U4365 (N_4365,N_3743,N_3659);
and U4366 (N_4366,N_3592,N_3600);
or U4367 (N_4367,N_3984,N_3696);
nand U4368 (N_4368,N_3735,N_3582);
nand U4369 (N_4369,N_3675,N_3752);
nand U4370 (N_4370,N_3954,N_3860);
nor U4371 (N_4371,N_3759,N_3689);
nand U4372 (N_4372,N_3604,N_3872);
and U4373 (N_4373,N_3841,N_3885);
nand U4374 (N_4374,N_3508,N_3655);
nand U4375 (N_4375,N_3766,N_3752);
xnor U4376 (N_4376,N_3586,N_3552);
or U4377 (N_4377,N_3718,N_3677);
or U4378 (N_4378,N_3586,N_3821);
nor U4379 (N_4379,N_3807,N_3965);
and U4380 (N_4380,N_3865,N_3818);
nor U4381 (N_4381,N_3582,N_3829);
nor U4382 (N_4382,N_3677,N_3829);
and U4383 (N_4383,N_3968,N_3738);
or U4384 (N_4384,N_3950,N_3753);
or U4385 (N_4385,N_3619,N_3945);
or U4386 (N_4386,N_3883,N_3920);
xor U4387 (N_4387,N_3657,N_3516);
xnor U4388 (N_4388,N_3672,N_3980);
nor U4389 (N_4389,N_3886,N_3864);
xor U4390 (N_4390,N_3711,N_3869);
xor U4391 (N_4391,N_3823,N_3914);
nor U4392 (N_4392,N_3997,N_3548);
nor U4393 (N_4393,N_3921,N_3542);
and U4394 (N_4394,N_3620,N_3952);
nand U4395 (N_4395,N_3617,N_3784);
nand U4396 (N_4396,N_3856,N_3880);
or U4397 (N_4397,N_3757,N_3995);
or U4398 (N_4398,N_3996,N_3729);
or U4399 (N_4399,N_3738,N_3971);
and U4400 (N_4400,N_3832,N_3548);
and U4401 (N_4401,N_3692,N_3965);
or U4402 (N_4402,N_3803,N_3933);
xnor U4403 (N_4403,N_3678,N_3734);
nor U4404 (N_4404,N_3977,N_3891);
or U4405 (N_4405,N_3875,N_3829);
nand U4406 (N_4406,N_3626,N_3843);
or U4407 (N_4407,N_3753,N_3769);
and U4408 (N_4408,N_3697,N_3638);
nor U4409 (N_4409,N_3959,N_3722);
or U4410 (N_4410,N_3808,N_3701);
xnor U4411 (N_4411,N_3981,N_3660);
or U4412 (N_4412,N_3926,N_3990);
xnor U4413 (N_4413,N_3558,N_3896);
nand U4414 (N_4414,N_3605,N_3904);
or U4415 (N_4415,N_3592,N_3905);
or U4416 (N_4416,N_3725,N_3718);
and U4417 (N_4417,N_3761,N_3521);
or U4418 (N_4418,N_3574,N_3911);
nor U4419 (N_4419,N_3509,N_3958);
xnor U4420 (N_4420,N_3508,N_3741);
and U4421 (N_4421,N_3635,N_3582);
xor U4422 (N_4422,N_3936,N_3528);
xor U4423 (N_4423,N_3577,N_3839);
or U4424 (N_4424,N_3874,N_3714);
nor U4425 (N_4425,N_3784,N_3863);
nand U4426 (N_4426,N_3733,N_3655);
and U4427 (N_4427,N_3672,N_3868);
xor U4428 (N_4428,N_3693,N_3672);
nand U4429 (N_4429,N_3507,N_3761);
or U4430 (N_4430,N_3958,N_3956);
nor U4431 (N_4431,N_3577,N_3988);
and U4432 (N_4432,N_3828,N_3884);
nor U4433 (N_4433,N_3565,N_3633);
nor U4434 (N_4434,N_3839,N_3992);
nand U4435 (N_4435,N_3823,N_3863);
nand U4436 (N_4436,N_3800,N_3566);
nand U4437 (N_4437,N_3772,N_3984);
or U4438 (N_4438,N_3534,N_3761);
xor U4439 (N_4439,N_3691,N_3956);
nand U4440 (N_4440,N_3797,N_3760);
nor U4441 (N_4441,N_3709,N_3507);
or U4442 (N_4442,N_3861,N_3648);
or U4443 (N_4443,N_3776,N_3917);
or U4444 (N_4444,N_3690,N_3517);
xor U4445 (N_4445,N_3839,N_3574);
or U4446 (N_4446,N_3551,N_3802);
nor U4447 (N_4447,N_3928,N_3882);
nor U4448 (N_4448,N_3577,N_3854);
nand U4449 (N_4449,N_3846,N_3756);
or U4450 (N_4450,N_3792,N_3690);
and U4451 (N_4451,N_3519,N_3595);
or U4452 (N_4452,N_3625,N_3965);
and U4453 (N_4453,N_3776,N_3826);
nor U4454 (N_4454,N_3969,N_3730);
nor U4455 (N_4455,N_3628,N_3885);
nand U4456 (N_4456,N_3832,N_3802);
or U4457 (N_4457,N_3621,N_3664);
nor U4458 (N_4458,N_3919,N_3989);
or U4459 (N_4459,N_3651,N_3746);
or U4460 (N_4460,N_3629,N_3795);
nand U4461 (N_4461,N_3948,N_3716);
nor U4462 (N_4462,N_3778,N_3720);
nand U4463 (N_4463,N_3506,N_3952);
and U4464 (N_4464,N_3618,N_3766);
and U4465 (N_4465,N_3629,N_3709);
nand U4466 (N_4466,N_3642,N_3726);
xnor U4467 (N_4467,N_3812,N_3937);
or U4468 (N_4468,N_3863,N_3942);
nand U4469 (N_4469,N_3755,N_3626);
and U4470 (N_4470,N_3880,N_3695);
nor U4471 (N_4471,N_3931,N_3732);
nand U4472 (N_4472,N_3666,N_3505);
xnor U4473 (N_4473,N_3998,N_3983);
xor U4474 (N_4474,N_3835,N_3685);
or U4475 (N_4475,N_3504,N_3602);
nand U4476 (N_4476,N_3688,N_3721);
xnor U4477 (N_4477,N_3521,N_3944);
nor U4478 (N_4478,N_3555,N_3966);
and U4479 (N_4479,N_3750,N_3906);
or U4480 (N_4480,N_3896,N_3980);
nor U4481 (N_4481,N_3976,N_3707);
nand U4482 (N_4482,N_3886,N_3717);
nand U4483 (N_4483,N_3669,N_3534);
and U4484 (N_4484,N_3962,N_3692);
xnor U4485 (N_4485,N_3838,N_3974);
or U4486 (N_4486,N_3615,N_3871);
nor U4487 (N_4487,N_3633,N_3907);
nand U4488 (N_4488,N_3733,N_3950);
nand U4489 (N_4489,N_3520,N_3515);
and U4490 (N_4490,N_3576,N_3777);
nor U4491 (N_4491,N_3636,N_3664);
or U4492 (N_4492,N_3851,N_3598);
nand U4493 (N_4493,N_3562,N_3623);
and U4494 (N_4494,N_3809,N_3598);
or U4495 (N_4495,N_3690,N_3664);
or U4496 (N_4496,N_3907,N_3909);
nor U4497 (N_4497,N_3694,N_3511);
xnor U4498 (N_4498,N_3898,N_3877);
xor U4499 (N_4499,N_3862,N_3856);
or U4500 (N_4500,N_4462,N_4461);
and U4501 (N_4501,N_4355,N_4379);
and U4502 (N_4502,N_4369,N_4258);
and U4503 (N_4503,N_4497,N_4053);
and U4504 (N_4504,N_4122,N_4101);
nand U4505 (N_4505,N_4309,N_4029);
xor U4506 (N_4506,N_4374,N_4399);
xnor U4507 (N_4507,N_4092,N_4103);
nor U4508 (N_4508,N_4175,N_4297);
nor U4509 (N_4509,N_4460,N_4128);
xor U4510 (N_4510,N_4123,N_4260);
and U4511 (N_4511,N_4179,N_4271);
xnor U4512 (N_4512,N_4344,N_4014);
nand U4513 (N_4513,N_4071,N_4219);
and U4514 (N_4514,N_4323,N_4320);
nor U4515 (N_4515,N_4276,N_4499);
and U4516 (N_4516,N_4305,N_4495);
and U4517 (N_4517,N_4069,N_4111);
xor U4518 (N_4518,N_4381,N_4050);
nand U4519 (N_4519,N_4058,N_4424);
nor U4520 (N_4520,N_4042,N_4070);
or U4521 (N_4521,N_4486,N_4159);
and U4522 (N_4522,N_4080,N_4131);
nor U4523 (N_4523,N_4075,N_4021);
or U4524 (N_4524,N_4234,N_4097);
xnor U4525 (N_4525,N_4190,N_4372);
xnor U4526 (N_4526,N_4206,N_4353);
xor U4527 (N_4527,N_4149,N_4456);
xnor U4528 (N_4528,N_4248,N_4140);
and U4529 (N_4529,N_4425,N_4384);
or U4530 (N_4530,N_4173,N_4336);
nor U4531 (N_4531,N_4283,N_4094);
or U4532 (N_4532,N_4154,N_4318);
nand U4533 (N_4533,N_4005,N_4221);
and U4534 (N_4534,N_4265,N_4035);
nand U4535 (N_4535,N_4196,N_4286);
xnor U4536 (N_4536,N_4376,N_4082);
nand U4537 (N_4537,N_4300,N_4361);
nand U4538 (N_4538,N_4441,N_4316);
and U4539 (N_4539,N_4394,N_4099);
or U4540 (N_4540,N_4423,N_4213);
and U4541 (N_4541,N_4409,N_4064);
or U4542 (N_4542,N_4313,N_4060);
and U4543 (N_4543,N_4270,N_4378);
xor U4544 (N_4544,N_4367,N_4209);
nor U4545 (N_4545,N_4051,N_4141);
nor U4546 (N_4546,N_4404,N_4467);
nand U4547 (N_4547,N_4208,N_4390);
or U4548 (N_4548,N_4307,N_4341);
nor U4549 (N_4549,N_4285,N_4397);
xnor U4550 (N_4550,N_4350,N_4298);
and U4551 (N_4551,N_4304,N_4192);
and U4552 (N_4552,N_4322,N_4373);
or U4553 (N_4553,N_4088,N_4231);
nor U4554 (N_4554,N_4411,N_4228);
nand U4555 (N_4555,N_4440,N_4072);
nor U4556 (N_4556,N_4057,N_4020);
nor U4557 (N_4557,N_4280,N_4161);
and U4558 (N_4558,N_4279,N_4427);
and U4559 (N_4559,N_4125,N_4386);
or U4560 (N_4560,N_4043,N_4056);
xor U4561 (N_4561,N_4335,N_4249);
or U4562 (N_4562,N_4430,N_4211);
nor U4563 (N_4563,N_4413,N_4330);
or U4564 (N_4564,N_4188,N_4337);
nor U4565 (N_4565,N_4429,N_4315);
nor U4566 (N_4566,N_4485,N_4358);
nor U4567 (N_4567,N_4025,N_4242);
and U4568 (N_4568,N_4135,N_4327);
xor U4569 (N_4569,N_4437,N_4257);
and U4570 (N_4570,N_4478,N_4116);
nand U4571 (N_4571,N_4143,N_4389);
xnor U4572 (N_4572,N_4172,N_4155);
nand U4573 (N_4573,N_4421,N_4366);
nor U4574 (N_4574,N_4450,N_4296);
or U4575 (N_4575,N_4026,N_4107);
nor U4576 (N_4576,N_4011,N_4459);
nand U4577 (N_4577,N_4292,N_4112);
and U4578 (N_4578,N_4207,N_4455);
nand U4579 (N_4579,N_4165,N_4266);
or U4580 (N_4580,N_4137,N_4342);
and U4581 (N_4581,N_4278,N_4045);
or U4582 (N_4582,N_4015,N_4134);
nand U4583 (N_4583,N_4079,N_4084);
and U4584 (N_4584,N_4040,N_4245);
xnor U4585 (N_4585,N_4465,N_4287);
and U4586 (N_4586,N_4244,N_4473);
and U4587 (N_4587,N_4120,N_4133);
or U4588 (N_4588,N_4181,N_4147);
nor U4589 (N_4589,N_4167,N_4275);
or U4590 (N_4590,N_4272,N_4210);
xor U4591 (N_4591,N_4252,N_4212);
or U4592 (N_4592,N_4146,N_4185);
or U4593 (N_4593,N_4180,N_4448);
xor U4594 (N_4594,N_4127,N_4178);
xnor U4595 (N_4595,N_4477,N_4375);
nor U4596 (N_4596,N_4498,N_4452);
xnor U4597 (N_4597,N_4062,N_4222);
or U4598 (N_4598,N_4301,N_4083);
nor U4599 (N_4599,N_4204,N_4326);
and U4600 (N_4600,N_4162,N_4281);
and U4601 (N_4601,N_4193,N_4293);
nor U4602 (N_4602,N_4377,N_4312);
or U4603 (N_4603,N_4205,N_4360);
or U4604 (N_4604,N_4481,N_4371);
and U4605 (N_4605,N_4416,N_4420);
or U4606 (N_4606,N_4008,N_4494);
or U4607 (N_4607,N_4232,N_4218);
nand U4608 (N_4608,N_4446,N_4152);
and U4609 (N_4609,N_4028,N_4226);
nor U4610 (N_4610,N_4233,N_4038);
and U4611 (N_4611,N_4264,N_4129);
nor U4612 (N_4612,N_4415,N_4414);
and U4613 (N_4613,N_4352,N_4151);
nand U4614 (N_4614,N_4086,N_4024);
nand U4615 (N_4615,N_4434,N_4000);
and U4616 (N_4616,N_4239,N_4447);
or U4617 (N_4617,N_4184,N_4200);
nand U4618 (N_4618,N_4321,N_4009);
and U4619 (N_4619,N_4126,N_4417);
nor U4620 (N_4620,N_4166,N_4194);
nor U4621 (N_4621,N_4302,N_4090);
and U4622 (N_4622,N_4346,N_4010);
or U4623 (N_4623,N_4001,N_4357);
nand U4624 (N_4624,N_4142,N_4263);
nor U4625 (N_4625,N_4401,N_4383);
or U4626 (N_4626,N_4457,N_4325);
and U4627 (N_4627,N_4453,N_4255);
nor U4628 (N_4628,N_4359,N_4023);
and U4629 (N_4629,N_4338,N_4018);
or U4630 (N_4630,N_4109,N_4114);
and U4631 (N_4631,N_4334,N_4468);
nor U4632 (N_4632,N_4329,N_4443);
or U4633 (N_4633,N_4382,N_4199);
nand U4634 (N_4634,N_4254,N_4105);
and U4635 (N_4635,N_4007,N_4391);
and U4636 (N_4636,N_4380,N_4076);
nand U4637 (N_4637,N_4354,N_4484);
nor U4638 (N_4638,N_4095,N_4170);
xor U4639 (N_4639,N_4136,N_4362);
or U4640 (N_4640,N_4093,N_4428);
nand U4641 (N_4641,N_4236,N_4482);
nand U4642 (N_4642,N_4130,N_4291);
nand U4643 (N_4643,N_4396,N_4229);
nor U4644 (N_4644,N_4235,N_4224);
nor U4645 (N_4645,N_4163,N_4253);
nand U4646 (N_4646,N_4066,N_4438);
or U4647 (N_4647,N_4158,N_4187);
nand U4648 (N_4648,N_4108,N_4124);
nor U4649 (N_4649,N_4483,N_4288);
or U4650 (N_4650,N_4189,N_4085);
and U4651 (N_4651,N_4032,N_4348);
or U4652 (N_4652,N_4393,N_4174);
or U4653 (N_4653,N_4282,N_4006);
or U4654 (N_4654,N_4148,N_4031);
nor U4655 (N_4655,N_4299,N_4306);
or U4656 (N_4656,N_4458,N_4488);
nand U4657 (N_4657,N_4487,N_4351);
and U4658 (N_4658,N_4104,N_4087);
or U4659 (N_4659,N_4017,N_4197);
nor U4660 (N_4660,N_4089,N_4356);
xnor U4661 (N_4661,N_4433,N_4345);
and U4662 (N_4662,N_4033,N_4418);
nor U4663 (N_4663,N_4160,N_4328);
or U4664 (N_4664,N_4308,N_4220);
xor U4665 (N_4665,N_4493,N_4157);
nor U4666 (N_4666,N_4259,N_4183);
nand U4667 (N_4667,N_4268,N_4339);
or U4668 (N_4668,N_4022,N_4474);
and U4669 (N_4669,N_4445,N_4340);
nand U4670 (N_4670,N_4150,N_4365);
and U4671 (N_4671,N_4078,N_4169);
or U4672 (N_4672,N_4289,N_4153);
nand U4673 (N_4673,N_4191,N_4041);
or U4674 (N_4674,N_4454,N_4449);
and U4675 (N_4675,N_4496,N_4403);
nand U4676 (N_4676,N_4004,N_4240);
xor U4677 (N_4677,N_4492,N_4223);
nand U4678 (N_4678,N_4471,N_4049);
or U4679 (N_4679,N_4177,N_4246);
nor U4680 (N_4680,N_4227,N_4171);
and U4681 (N_4681,N_4466,N_4347);
xor U4682 (N_4682,N_4214,N_4139);
nor U4683 (N_4683,N_4364,N_4310);
nor U4684 (N_4684,N_4113,N_4405);
or U4685 (N_4685,N_4479,N_4256);
nand U4686 (N_4686,N_4463,N_4324);
nor U4687 (N_4687,N_4491,N_4052);
or U4688 (N_4688,N_4034,N_4182);
or U4689 (N_4689,N_4048,N_4274);
nand U4690 (N_4690,N_4406,N_4277);
nand U4691 (N_4691,N_4115,N_4439);
and U4692 (N_4692,N_4030,N_4349);
xor U4693 (N_4693,N_4431,N_4398);
nand U4694 (N_4694,N_4370,N_4436);
nor U4695 (N_4695,N_4238,N_4016);
nor U4696 (N_4696,N_4273,N_4201);
nand U4697 (N_4697,N_4117,N_4261);
or U4698 (N_4698,N_4119,N_4480);
nand U4699 (N_4699,N_4195,N_4395);
nor U4700 (N_4700,N_4444,N_4419);
nand U4701 (N_4701,N_4055,N_4046);
nand U4702 (N_4702,N_4217,N_4290);
and U4703 (N_4703,N_4475,N_4063);
nor U4704 (N_4704,N_4145,N_4392);
nand U4705 (N_4705,N_4077,N_4451);
and U4706 (N_4706,N_4102,N_4317);
and U4707 (N_4707,N_4118,N_4247);
or U4708 (N_4708,N_4412,N_4402);
or U4709 (N_4709,N_4216,N_4138);
nand U4710 (N_4710,N_4472,N_4039);
and U4711 (N_4711,N_4303,N_4490);
nor U4712 (N_4712,N_4203,N_4269);
nor U4713 (N_4713,N_4435,N_4100);
or U4714 (N_4714,N_4110,N_4091);
nand U4715 (N_4715,N_4002,N_4476);
or U4716 (N_4716,N_4343,N_4262);
or U4717 (N_4717,N_4284,N_4098);
nand U4718 (N_4718,N_4164,N_4037);
nand U4719 (N_4719,N_4408,N_4132);
nor U4720 (N_4720,N_4106,N_4096);
or U4721 (N_4721,N_4363,N_4202);
and U4722 (N_4722,N_4225,N_4065);
nand U4723 (N_4723,N_4019,N_4168);
and U4724 (N_4724,N_4144,N_4311);
or U4725 (N_4725,N_4027,N_4410);
nor U4726 (N_4726,N_4426,N_4368);
or U4727 (N_4727,N_4059,N_4003);
nor U4728 (N_4728,N_4044,N_4176);
or U4729 (N_4729,N_4388,N_4156);
nor U4730 (N_4730,N_4295,N_4422);
or U4731 (N_4731,N_4469,N_4121);
or U4732 (N_4732,N_4067,N_4333);
nor U4733 (N_4733,N_4314,N_4387);
and U4734 (N_4734,N_4215,N_4250);
nor U4735 (N_4735,N_4385,N_4251);
nand U4736 (N_4736,N_4186,N_4332);
nor U4737 (N_4737,N_4237,N_4036);
nand U4738 (N_4738,N_4241,N_4068);
and U4739 (N_4739,N_4267,N_4073);
nor U4740 (N_4740,N_4230,N_4081);
or U4741 (N_4741,N_4331,N_4061);
and U4742 (N_4742,N_4407,N_4400);
or U4743 (N_4743,N_4432,N_4054);
nor U4744 (N_4744,N_4319,N_4243);
xor U4745 (N_4745,N_4442,N_4489);
nand U4746 (N_4746,N_4012,N_4047);
or U4747 (N_4747,N_4464,N_4074);
or U4748 (N_4748,N_4294,N_4198);
nor U4749 (N_4749,N_4470,N_4013);
nor U4750 (N_4750,N_4220,N_4474);
nand U4751 (N_4751,N_4002,N_4352);
and U4752 (N_4752,N_4408,N_4489);
or U4753 (N_4753,N_4336,N_4389);
nand U4754 (N_4754,N_4383,N_4145);
nor U4755 (N_4755,N_4289,N_4269);
nor U4756 (N_4756,N_4200,N_4085);
or U4757 (N_4757,N_4491,N_4317);
and U4758 (N_4758,N_4407,N_4013);
nor U4759 (N_4759,N_4323,N_4073);
nor U4760 (N_4760,N_4138,N_4286);
xnor U4761 (N_4761,N_4008,N_4240);
xor U4762 (N_4762,N_4164,N_4443);
or U4763 (N_4763,N_4172,N_4118);
or U4764 (N_4764,N_4318,N_4291);
or U4765 (N_4765,N_4365,N_4050);
nand U4766 (N_4766,N_4293,N_4106);
or U4767 (N_4767,N_4130,N_4365);
nand U4768 (N_4768,N_4075,N_4495);
nor U4769 (N_4769,N_4261,N_4343);
nor U4770 (N_4770,N_4445,N_4087);
or U4771 (N_4771,N_4427,N_4186);
and U4772 (N_4772,N_4042,N_4429);
or U4773 (N_4773,N_4275,N_4294);
and U4774 (N_4774,N_4456,N_4002);
or U4775 (N_4775,N_4160,N_4488);
xor U4776 (N_4776,N_4298,N_4269);
nor U4777 (N_4777,N_4103,N_4459);
nand U4778 (N_4778,N_4095,N_4275);
or U4779 (N_4779,N_4495,N_4419);
and U4780 (N_4780,N_4352,N_4147);
nand U4781 (N_4781,N_4385,N_4188);
nor U4782 (N_4782,N_4192,N_4346);
nor U4783 (N_4783,N_4348,N_4081);
or U4784 (N_4784,N_4221,N_4282);
nor U4785 (N_4785,N_4393,N_4346);
nand U4786 (N_4786,N_4033,N_4417);
nor U4787 (N_4787,N_4354,N_4282);
xor U4788 (N_4788,N_4165,N_4398);
xnor U4789 (N_4789,N_4321,N_4418);
and U4790 (N_4790,N_4159,N_4327);
or U4791 (N_4791,N_4423,N_4498);
nand U4792 (N_4792,N_4391,N_4231);
nand U4793 (N_4793,N_4327,N_4482);
nor U4794 (N_4794,N_4473,N_4113);
nor U4795 (N_4795,N_4034,N_4035);
xnor U4796 (N_4796,N_4001,N_4434);
nor U4797 (N_4797,N_4257,N_4324);
and U4798 (N_4798,N_4235,N_4367);
nand U4799 (N_4799,N_4229,N_4444);
or U4800 (N_4800,N_4029,N_4424);
nand U4801 (N_4801,N_4086,N_4372);
nand U4802 (N_4802,N_4334,N_4051);
xor U4803 (N_4803,N_4092,N_4271);
and U4804 (N_4804,N_4214,N_4151);
nand U4805 (N_4805,N_4118,N_4126);
nand U4806 (N_4806,N_4267,N_4013);
or U4807 (N_4807,N_4324,N_4024);
xor U4808 (N_4808,N_4410,N_4061);
or U4809 (N_4809,N_4027,N_4387);
xor U4810 (N_4810,N_4057,N_4302);
or U4811 (N_4811,N_4461,N_4056);
or U4812 (N_4812,N_4149,N_4359);
and U4813 (N_4813,N_4036,N_4438);
nor U4814 (N_4814,N_4286,N_4191);
and U4815 (N_4815,N_4003,N_4075);
nor U4816 (N_4816,N_4191,N_4112);
nand U4817 (N_4817,N_4494,N_4174);
or U4818 (N_4818,N_4377,N_4436);
nand U4819 (N_4819,N_4000,N_4342);
nor U4820 (N_4820,N_4314,N_4130);
nor U4821 (N_4821,N_4351,N_4073);
or U4822 (N_4822,N_4110,N_4130);
nand U4823 (N_4823,N_4338,N_4281);
nand U4824 (N_4824,N_4048,N_4308);
xnor U4825 (N_4825,N_4350,N_4498);
nor U4826 (N_4826,N_4071,N_4383);
and U4827 (N_4827,N_4022,N_4202);
and U4828 (N_4828,N_4459,N_4382);
or U4829 (N_4829,N_4062,N_4448);
or U4830 (N_4830,N_4445,N_4106);
nor U4831 (N_4831,N_4020,N_4149);
xor U4832 (N_4832,N_4166,N_4255);
xnor U4833 (N_4833,N_4333,N_4158);
or U4834 (N_4834,N_4474,N_4298);
nand U4835 (N_4835,N_4322,N_4442);
or U4836 (N_4836,N_4392,N_4263);
nor U4837 (N_4837,N_4184,N_4386);
or U4838 (N_4838,N_4392,N_4023);
or U4839 (N_4839,N_4238,N_4288);
nand U4840 (N_4840,N_4302,N_4012);
nand U4841 (N_4841,N_4433,N_4193);
nand U4842 (N_4842,N_4375,N_4243);
xnor U4843 (N_4843,N_4262,N_4260);
or U4844 (N_4844,N_4059,N_4006);
nor U4845 (N_4845,N_4141,N_4166);
nor U4846 (N_4846,N_4402,N_4002);
nor U4847 (N_4847,N_4334,N_4458);
or U4848 (N_4848,N_4054,N_4152);
or U4849 (N_4849,N_4053,N_4039);
xor U4850 (N_4850,N_4305,N_4466);
nand U4851 (N_4851,N_4039,N_4486);
nand U4852 (N_4852,N_4072,N_4257);
nand U4853 (N_4853,N_4047,N_4050);
and U4854 (N_4854,N_4193,N_4361);
nand U4855 (N_4855,N_4376,N_4313);
xor U4856 (N_4856,N_4160,N_4148);
and U4857 (N_4857,N_4365,N_4248);
or U4858 (N_4858,N_4475,N_4452);
xor U4859 (N_4859,N_4096,N_4285);
and U4860 (N_4860,N_4372,N_4443);
nor U4861 (N_4861,N_4311,N_4401);
and U4862 (N_4862,N_4133,N_4046);
and U4863 (N_4863,N_4273,N_4307);
and U4864 (N_4864,N_4387,N_4487);
xor U4865 (N_4865,N_4440,N_4258);
nand U4866 (N_4866,N_4487,N_4488);
and U4867 (N_4867,N_4243,N_4030);
or U4868 (N_4868,N_4159,N_4179);
nor U4869 (N_4869,N_4192,N_4442);
and U4870 (N_4870,N_4131,N_4324);
nand U4871 (N_4871,N_4487,N_4453);
xor U4872 (N_4872,N_4198,N_4237);
or U4873 (N_4873,N_4074,N_4119);
nor U4874 (N_4874,N_4315,N_4354);
nor U4875 (N_4875,N_4174,N_4312);
nor U4876 (N_4876,N_4064,N_4000);
or U4877 (N_4877,N_4048,N_4044);
nor U4878 (N_4878,N_4070,N_4413);
and U4879 (N_4879,N_4163,N_4499);
or U4880 (N_4880,N_4090,N_4349);
or U4881 (N_4881,N_4226,N_4012);
xor U4882 (N_4882,N_4319,N_4333);
or U4883 (N_4883,N_4314,N_4039);
nor U4884 (N_4884,N_4094,N_4020);
or U4885 (N_4885,N_4035,N_4359);
and U4886 (N_4886,N_4359,N_4394);
and U4887 (N_4887,N_4465,N_4444);
and U4888 (N_4888,N_4085,N_4385);
and U4889 (N_4889,N_4193,N_4150);
xnor U4890 (N_4890,N_4237,N_4377);
and U4891 (N_4891,N_4267,N_4051);
xor U4892 (N_4892,N_4408,N_4201);
nand U4893 (N_4893,N_4056,N_4044);
and U4894 (N_4894,N_4130,N_4157);
nand U4895 (N_4895,N_4350,N_4404);
nand U4896 (N_4896,N_4059,N_4255);
or U4897 (N_4897,N_4171,N_4388);
nor U4898 (N_4898,N_4456,N_4437);
nor U4899 (N_4899,N_4433,N_4468);
nor U4900 (N_4900,N_4192,N_4012);
xnor U4901 (N_4901,N_4118,N_4322);
nor U4902 (N_4902,N_4260,N_4370);
or U4903 (N_4903,N_4463,N_4292);
and U4904 (N_4904,N_4127,N_4286);
nand U4905 (N_4905,N_4405,N_4252);
nand U4906 (N_4906,N_4048,N_4467);
and U4907 (N_4907,N_4062,N_4497);
or U4908 (N_4908,N_4364,N_4373);
or U4909 (N_4909,N_4228,N_4111);
nor U4910 (N_4910,N_4298,N_4047);
nor U4911 (N_4911,N_4015,N_4482);
xnor U4912 (N_4912,N_4265,N_4178);
or U4913 (N_4913,N_4166,N_4216);
or U4914 (N_4914,N_4370,N_4144);
xnor U4915 (N_4915,N_4371,N_4023);
and U4916 (N_4916,N_4176,N_4390);
and U4917 (N_4917,N_4425,N_4170);
nand U4918 (N_4918,N_4364,N_4446);
xor U4919 (N_4919,N_4113,N_4452);
nand U4920 (N_4920,N_4197,N_4441);
and U4921 (N_4921,N_4013,N_4272);
or U4922 (N_4922,N_4197,N_4315);
nand U4923 (N_4923,N_4137,N_4173);
or U4924 (N_4924,N_4494,N_4132);
nand U4925 (N_4925,N_4387,N_4355);
nand U4926 (N_4926,N_4350,N_4104);
and U4927 (N_4927,N_4392,N_4474);
or U4928 (N_4928,N_4471,N_4115);
nor U4929 (N_4929,N_4200,N_4008);
or U4930 (N_4930,N_4342,N_4068);
and U4931 (N_4931,N_4246,N_4353);
or U4932 (N_4932,N_4400,N_4004);
nor U4933 (N_4933,N_4031,N_4410);
and U4934 (N_4934,N_4256,N_4035);
and U4935 (N_4935,N_4032,N_4395);
nand U4936 (N_4936,N_4182,N_4257);
nand U4937 (N_4937,N_4132,N_4498);
xnor U4938 (N_4938,N_4483,N_4414);
and U4939 (N_4939,N_4443,N_4110);
or U4940 (N_4940,N_4078,N_4104);
xnor U4941 (N_4941,N_4279,N_4403);
or U4942 (N_4942,N_4003,N_4073);
or U4943 (N_4943,N_4319,N_4412);
nand U4944 (N_4944,N_4052,N_4206);
and U4945 (N_4945,N_4434,N_4174);
nand U4946 (N_4946,N_4112,N_4483);
nand U4947 (N_4947,N_4414,N_4149);
nand U4948 (N_4948,N_4285,N_4199);
or U4949 (N_4949,N_4239,N_4420);
and U4950 (N_4950,N_4291,N_4411);
or U4951 (N_4951,N_4135,N_4296);
nand U4952 (N_4952,N_4142,N_4158);
nor U4953 (N_4953,N_4451,N_4174);
and U4954 (N_4954,N_4086,N_4442);
nand U4955 (N_4955,N_4329,N_4470);
nand U4956 (N_4956,N_4121,N_4414);
nor U4957 (N_4957,N_4008,N_4315);
or U4958 (N_4958,N_4133,N_4003);
nor U4959 (N_4959,N_4006,N_4236);
and U4960 (N_4960,N_4037,N_4187);
and U4961 (N_4961,N_4218,N_4369);
nor U4962 (N_4962,N_4250,N_4415);
and U4963 (N_4963,N_4201,N_4114);
and U4964 (N_4964,N_4344,N_4065);
or U4965 (N_4965,N_4129,N_4076);
and U4966 (N_4966,N_4159,N_4265);
nor U4967 (N_4967,N_4273,N_4366);
or U4968 (N_4968,N_4006,N_4381);
nand U4969 (N_4969,N_4030,N_4126);
nor U4970 (N_4970,N_4473,N_4240);
nand U4971 (N_4971,N_4395,N_4109);
or U4972 (N_4972,N_4212,N_4000);
nand U4973 (N_4973,N_4106,N_4495);
xor U4974 (N_4974,N_4430,N_4114);
or U4975 (N_4975,N_4214,N_4403);
and U4976 (N_4976,N_4216,N_4108);
nor U4977 (N_4977,N_4266,N_4042);
nor U4978 (N_4978,N_4289,N_4182);
and U4979 (N_4979,N_4205,N_4432);
nand U4980 (N_4980,N_4145,N_4173);
and U4981 (N_4981,N_4120,N_4338);
nor U4982 (N_4982,N_4356,N_4404);
xor U4983 (N_4983,N_4433,N_4013);
nor U4984 (N_4984,N_4282,N_4145);
and U4985 (N_4985,N_4220,N_4047);
nand U4986 (N_4986,N_4302,N_4000);
or U4987 (N_4987,N_4088,N_4045);
xnor U4988 (N_4988,N_4183,N_4174);
nand U4989 (N_4989,N_4423,N_4334);
nand U4990 (N_4990,N_4490,N_4241);
and U4991 (N_4991,N_4397,N_4030);
xor U4992 (N_4992,N_4077,N_4320);
or U4993 (N_4993,N_4039,N_4295);
or U4994 (N_4994,N_4447,N_4463);
or U4995 (N_4995,N_4050,N_4021);
nand U4996 (N_4996,N_4001,N_4278);
or U4997 (N_4997,N_4093,N_4005);
and U4998 (N_4998,N_4250,N_4126);
nand U4999 (N_4999,N_4106,N_4072);
or UO_0 (O_0,N_4510,N_4709);
nand UO_1 (O_1,N_4865,N_4821);
xor UO_2 (O_2,N_4803,N_4917);
nor UO_3 (O_3,N_4848,N_4653);
and UO_4 (O_4,N_4594,N_4868);
or UO_5 (O_5,N_4613,N_4824);
nor UO_6 (O_6,N_4669,N_4684);
and UO_7 (O_7,N_4621,N_4642);
nand UO_8 (O_8,N_4553,N_4651);
nor UO_9 (O_9,N_4729,N_4742);
nor UO_10 (O_10,N_4864,N_4785);
nor UO_11 (O_11,N_4969,N_4750);
nand UO_12 (O_12,N_4609,N_4880);
nor UO_13 (O_13,N_4717,N_4567);
nor UO_14 (O_14,N_4892,N_4850);
or UO_15 (O_15,N_4818,N_4928);
xor UO_16 (O_16,N_4871,N_4507);
nor UO_17 (O_17,N_4731,N_4828);
or UO_18 (O_18,N_4734,N_4679);
or UO_19 (O_19,N_4541,N_4506);
nor UO_20 (O_20,N_4598,N_4988);
nand UO_21 (O_21,N_4820,N_4649);
and UO_22 (O_22,N_4979,N_4667);
nand UO_23 (O_23,N_4557,N_4695);
nor UO_24 (O_24,N_4861,N_4964);
nor UO_25 (O_25,N_4636,N_4602);
or UO_26 (O_26,N_4739,N_4834);
nor UO_27 (O_27,N_4978,N_4758);
nand UO_28 (O_28,N_4652,N_4799);
and UO_29 (O_29,N_4935,N_4592);
or UO_30 (O_30,N_4873,N_4671);
xnor UO_31 (O_31,N_4766,N_4955);
or UO_32 (O_32,N_4989,N_4555);
xnor UO_33 (O_33,N_4833,N_4909);
nor UO_34 (O_34,N_4640,N_4844);
and UO_35 (O_35,N_4749,N_4701);
or UO_36 (O_36,N_4761,N_4681);
nand UO_37 (O_37,N_4804,N_4812);
and UO_38 (O_38,N_4568,N_4891);
nor UO_39 (O_39,N_4948,N_4823);
nor UO_40 (O_40,N_4523,N_4806);
and UO_41 (O_41,N_4554,N_4607);
xnor UO_42 (O_42,N_4784,N_4528);
xnor UO_43 (O_43,N_4614,N_4797);
nand UO_44 (O_44,N_4811,N_4566);
xnor UO_45 (O_45,N_4662,N_4796);
nor UO_46 (O_46,N_4884,N_4882);
nor UO_47 (O_47,N_4929,N_4902);
and UO_48 (O_48,N_4582,N_4793);
or UO_49 (O_49,N_4872,N_4854);
or UO_50 (O_50,N_4942,N_4565);
and UO_51 (O_51,N_4950,N_4561);
and UO_52 (O_52,N_4837,N_4801);
or UO_53 (O_53,N_4774,N_4841);
or UO_54 (O_54,N_4772,N_4617);
or UO_55 (O_55,N_4502,N_4960);
and UO_56 (O_56,N_4623,N_4646);
or UO_57 (O_57,N_4922,N_4580);
nor UO_58 (O_58,N_4672,N_4520);
or UO_59 (O_59,N_4608,N_4515);
or UO_60 (O_60,N_4959,N_4773);
nand UO_61 (O_61,N_4866,N_4511);
nand UO_62 (O_62,N_4665,N_4603);
and UO_63 (O_63,N_4763,N_4753);
and UO_64 (O_64,N_4759,N_4712);
xor UO_65 (O_65,N_4674,N_4707);
and UO_66 (O_66,N_4680,N_4764);
xor UO_67 (O_67,N_4663,N_4659);
nor UO_68 (O_68,N_4536,N_4914);
nand UO_69 (O_69,N_4904,N_4738);
and UO_70 (O_70,N_4626,N_4857);
and UO_71 (O_71,N_4692,N_4666);
xnor UO_72 (O_72,N_4984,N_4588);
nor UO_73 (O_73,N_4503,N_4747);
and UO_74 (O_74,N_4635,N_4877);
and UO_75 (O_75,N_4853,N_4581);
nor UO_76 (O_76,N_4843,N_4593);
and UO_77 (O_77,N_4863,N_4847);
nand UO_78 (O_78,N_4519,N_4965);
nor UO_79 (O_79,N_4745,N_4654);
nor UO_80 (O_80,N_4903,N_4893);
nand UO_81 (O_81,N_4618,N_4562);
nand UO_82 (O_82,N_4631,N_4547);
or UO_83 (O_83,N_4957,N_4549);
or UO_84 (O_84,N_4532,N_4831);
or UO_85 (O_85,N_4619,N_4897);
nor UO_86 (O_86,N_4934,N_4668);
nand UO_87 (O_87,N_4995,N_4779);
or UO_88 (O_88,N_4702,N_4842);
and UO_89 (O_89,N_4725,N_4658);
nor UO_90 (O_90,N_4748,N_4974);
nand UO_91 (O_91,N_4787,N_4870);
or UO_92 (O_92,N_4556,N_4767);
nor UO_93 (O_93,N_4599,N_4878);
and UO_94 (O_94,N_4650,N_4685);
and UO_95 (O_95,N_4505,N_4887);
nand UO_96 (O_96,N_4961,N_4782);
nor UO_97 (O_97,N_4611,N_4776);
and UO_98 (O_98,N_4573,N_4958);
nand UO_99 (O_99,N_4920,N_4867);
and UO_100 (O_100,N_4604,N_4901);
nor UO_101 (O_101,N_4713,N_4938);
nor UO_102 (O_102,N_4587,N_4660);
and UO_103 (O_103,N_4625,N_4544);
nor UO_104 (O_104,N_4673,N_4813);
nand UO_105 (O_105,N_4912,N_4710);
or UO_106 (O_106,N_4876,N_4992);
nor UO_107 (O_107,N_4817,N_4550);
and UO_108 (O_108,N_4762,N_4932);
nand UO_109 (O_109,N_4976,N_4775);
or UO_110 (O_110,N_4634,N_4832);
and UO_111 (O_111,N_4825,N_4620);
and UO_112 (O_112,N_4682,N_4736);
and UO_113 (O_113,N_4805,N_4839);
or UO_114 (O_114,N_4894,N_4540);
and UO_115 (O_115,N_4687,N_4810);
nand UO_116 (O_116,N_4661,N_4786);
nand UO_117 (O_117,N_4918,N_4508);
or UO_118 (O_118,N_4644,N_4951);
or UO_119 (O_119,N_4744,N_4535);
and UO_120 (O_120,N_4728,N_4898);
or UO_121 (O_121,N_4778,N_4755);
or UO_122 (O_122,N_4790,N_4977);
and UO_123 (O_123,N_4916,N_4829);
nand UO_124 (O_124,N_4911,N_4596);
and UO_125 (O_125,N_4648,N_4874);
nor UO_126 (O_126,N_4597,N_4907);
nor UO_127 (O_127,N_4791,N_4963);
and UO_128 (O_128,N_4858,N_4576);
nor UO_129 (O_129,N_4962,N_4983);
nand UO_130 (O_130,N_4639,N_4579);
and UO_131 (O_131,N_4572,N_4973);
or UO_132 (O_132,N_4690,N_4972);
nor UO_133 (O_133,N_4906,N_4723);
and UO_134 (O_134,N_4971,N_4622);
nand UO_135 (O_135,N_4706,N_4548);
nand UO_136 (O_136,N_4678,N_4585);
nor UO_137 (O_137,N_4543,N_4610);
and UO_138 (O_138,N_4638,N_4967);
nand UO_139 (O_139,N_4569,N_4986);
and UO_140 (O_140,N_4531,N_4746);
nor UO_141 (O_141,N_4605,N_4500);
nor UO_142 (O_142,N_4840,N_4838);
nor UO_143 (O_143,N_4693,N_4643);
nor UO_144 (O_144,N_4526,N_4924);
or UO_145 (O_145,N_4601,N_4947);
or UO_146 (O_146,N_4835,N_4931);
nand UO_147 (O_147,N_4885,N_4954);
nor UO_148 (O_148,N_4563,N_4591);
or UO_149 (O_149,N_4637,N_4645);
nor UO_150 (O_150,N_4560,N_4590);
xor UO_151 (O_151,N_4875,N_4883);
and UO_152 (O_152,N_4760,N_4987);
nand UO_153 (O_153,N_4732,N_4985);
nand UO_154 (O_154,N_4752,N_4765);
nor UO_155 (O_155,N_4718,N_4656);
or UO_156 (O_156,N_4552,N_4851);
nand UO_157 (O_157,N_4720,N_4628);
and UO_158 (O_158,N_4941,N_4647);
nand UO_159 (O_159,N_4996,N_4533);
nor UO_160 (O_160,N_4769,N_4538);
xnor UO_161 (O_161,N_4798,N_4937);
nand UO_162 (O_162,N_4991,N_4641);
and UO_163 (O_163,N_4711,N_4952);
and UO_164 (O_164,N_4719,N_4516);
and UO_165 (O_165,N_4923,N_4514);
xnor UO_166 (O_166,N_4993,N_4949);
nor UO_167 (O_167,N_4836,N_4664);
nand UO_168 (O_168,N_4852,N_4694);
nand UO_169 (O_169,N_4808,N_4730);
nor UO_170 (O_170,N_4830,N_4633);
and UO_171 (O_171,N_4819,N_4722);
nand UO_172 (O_172,N_4794,N_4677);
nand UO_173 (O_173,N_4975,N_4615);
or UO_174 (O_174,N_4657,N_4716);
or UO_175 (O_175,N_4869,N_4703);
and UO_176 (O_176,N_4910,N_4956);
nand UO_177 (O_177,N_4529,N_4783);
nand UO_178 (O_178,N_4606,N_4525);
or UO_179 (O_179,N_4899,N_4751);
or UO_180 (O_180,N_4683,N_4913);
xor UO_181 (O_181,N_4822,N_4921);
or UO_182 (O_182,N_4578,N_4925);
or UO_183 (O_183,N_4518,N_4890);
nand UO_184 (O_184,N_4757,N_4688);
nand UO_185 (O_185,N_4564,N_4809);
nand UO_186 (O_186,N_4524,N_4629);
nor UO_187 (O_187,N_4612,N_4999);
or UO_188 (O_188,N_4792,N_4943);
nand UO_189 (O_189,N_4940,N_4849);
nor UO_190 (O_190,N_4704,N_4551);
nand UO_191 (O_191,N_4827,N_4781);
or UO_192 (O_192,N_4737,N_4945);
nand UO_193 (O_193,N_4559,N_4754);
xnor UO_194 (O_194,N_4616,N_4741);
nand UO_195 (O_195,N_4926,N_4727);
xor UO_196 (O_196,N_4517,N_4896);
and UO_197 (O_197,N_4595,N_4530);
nor UO_198 (O_198,N_4708,N_4802);
or UO_199 (O_199,N_4800,N_4527);
and UO_200 (O_200,N_4862,N_4655);
xor UO_201 (O_201,N_4521,N_4994);
or UO_202 (O_202,N_4721,N_4586);
and UO_203 (O_203,N_4879,N_4715);
and UO_204 (O_204,N_4675,N_4600);
nor UO_205 (O_205,N_4905,N_4982);
nor UO_206 (O_206,N_4589,N_4970);
nor UO_207 (O_207,N_4539,N_4933);
nand UO_208 (O_208,N_4768,N_4788);
nand UO_209 (O_209,N_4930,N_4714);
nor UO_210 (O_210,N_4889,N_4733);
nor UO_211 (O_211,N_4845,N_4501);
nand UO_212 (O_212,N_4630,N_4537);
xnor UO_213 (O_213,N_4856,N_4908);
and UO_214 (O_214,N_4670,N_4574);
and UO_215 (O_215,N_4575,N_4504);
xor UO_216 (O_216,N_4946,N_4855);
and UO_217 (O_217,N_4927,N_4583);
or UO_218 (O_218,N_4881,N_4944);
or UO_219 (O_219,N_4522,N_4735);
nand UO_220 (O_220,N_4696,N_4936);
or UO_221 (O_221,N_4698,N_4546);
nand UO_222 (O_222,N_4697,N_4816);
or UO_223 (O_223,N_4826,N_4900);
nand UO_224 (O_224,N_4997,N_4699);
or UO_225 (O_225,N_4571,N_4726);
and UO_226 (O_226,N_4990,N_4570);
or UO_227 (O_227,N_4939,N_4577);
nor UO_228 (O_228,N_4513,N_4686);
xor UO_229 (O_229,N_4743,N_4558);
or UO_230 (O_230,N_4968,N_4886);
and UO_231 (O_231,N_4807,N_4915);
nand UO_232 (O_232,N_4724,N_4700);
nand UO_233 (O_233,N_4691,N_4895);
xnor UO_234 (O_234,N_4814,N_4627);
nand UO_235 (O_235,N_4512,N_4980);
nor UO_236 (O_236,N_4756,N_4676);
xnor UO_237 (O_237,N_4998,N_4888);
nand UO_238 (O_238,N_4689,N_4789);
nor UO_239 (O_239,N_4846,N_4771);
or UO_240 (O_240,N_4542,N_4860);
or UO_241 (O_241,N_4966,N_4545);
and UO_242 (O_242,N_4770,N_4624);
nand UO_243 (O_243,N_4534,N_4740);
nor UO_244 (O_244,N_4953,N_4859);
and UO_245 (O_245,N_4509,N_4795);
nor UO_246 (O_246,N_4919,N_4777);
nor UO_247 (O_247,N_4981,N_4815);
nand UO_248 (O_248,N_4584,N_4780);
and UO_249 (O_249,N_4705,N_4632);
nor UO_250 (O_250,N_4931,N_4506);
and UO_251 (O_251,N_4564,N_4935);
or UO_252 (O_252,N_4676,N_4977);
and UO_253 (O_253,N_4673,N_4561);
xnor UO_254 (O_254,N_4669,N_4567);
nand UO_255 (O_255,N_4800,N_4850);
or UO_256 (O_256,N_4894,N_4763);
nand UO_257 (O_257,N_4565,N_4508);
xnor UO_258 (O_258,N_4881,N_4649);
and UO_259 (O_259,N_4596,N_4877);
nor UO_260 (O_260,N_4966,N_4615);
xor UO_261 (O_261,N_4653,N_4594);
and UO_262 (O_262,N_4797,N_4732);
nand UO_263 (O_263,N_4993,N_4701);
or UO_264 (O_264,N_4969,N_4994);
xor UO_265 (O_265,N_4558,N_4918);
nor UO_266 (O_266,N_4519,N_4725);
nand UO_267 (O_267,N_4988,N_4674);
and UO_268 (O_268,N_4863,N_4643);
or UO_269 (O_269,N_4947,N_4788);
and UO_270 (O_270,N_4974,N_4689);
or UO_271 (O_271,N_4983,N_4824);
and UO_272 (O_272,N_4758,N_4565);
nor UO_273 (O_273,N_4887,N_4936);
or UO_274 (O_274,N_4918,N_4795);
or UO_275 (O_275,N_4553,N_4674);
and UO_276 (O_276,N_4824,N_4607);
nand UO_277 (O_277,N_4793,N_4976);
nand UO_278 (O_278,N_4722,N_4882);
or UO_279 (O_279,N_4695,N_4535);
nor UO_280 (O_280,N_4548,N_4560);
and UO_281 (O_281,N_4914,N_4699);
and UO_282 (O_282,N_4566,N_4942);
nor UO_283 (O_283,N_4978,N_4911);
nand UO_284 (O_284,N_4811,N_4544);
nor UO_285 (O_285,N_4581,N_4623);
nor UO_286 (O_286,N_4782,N_4806);
nor UO_287 (O_287,N_4593,N_4882);
nand UO_288 (O_288,N_4546,N_4704);
xor UO_289 (O_289,N_4531,N_4571);
and UO_290 (O_290,N_4601,N_4578);
and UO_291 (O_291,N_4542,N_4982);
xor UO_292 (O_292,N_4620,N_4616);
nand UO_293 (O_293,N_4735,N_4957);
or UO_294 (O_294,N_4850,N_4986);
and UO_295 (O_295,N_4734,N_4776);
and UO_296 (O_296,N_4950,N_4645);
nor UO_297 (O_297,N_4816,N_4909);
nor UO_298 (O_298,N_4614,N_4665);
nand UO_299 (O_299,N_4555,N_4940);
nand UO_300 (O_300,N_4927,N_4688);
and UO_301 (O_301,N_4609,N_4954);
or UO_302 (O_302,N_4979,N_4759);
or UO_303 (O_303,N_4634,N_4670);
and UO_304 (O_304,N_4530,N_4845);
nor UO_305 (O_305,N_4770,N_4588);
nor UO_306 (O_306,N_4910,N_4648);
or UO_307 (O_307,N_4743,N_4636);
nor UO_308 (O_308,N_4979,N_4893);
and UO_309 (O_309,N_4753,N_4810);
and UO_310 (O_310,N_4998,N_4557);
and UO_311 (O_311,N_4892,N_4593);
or UO_312 (O_312,N_4647,N_4544);
and UO_313 (O_313,N_4829,N_4651);
nor UO_314 (O_314,N_4509,N_4728);
or UO_315 (O_315,N_4631,N_4766);
xnor UO_316 (O_316,N_4944,N_4599);
nor UO_317 (O_317,N_4965,N_4592);
nand UO_318 (O_318,N_4788,N_4883);
nand UO_319 (O_319,N_4882,N_4694);
and UO_320 (O_320,N_4527,N_4677);
nand UO_321 (O_321,N_4647,N_4802);
or UO_322 (O_322,N_4772,N_4621);
nor UO_323 (O_323,N_4934,N_4935);
or UO_324 (O_324,N_4672,N_4794);
and UO_325 (O_325,N_4624,N_4986);
nand UO_326 (O_326,N_4895,N_4765);
or UO_327 (O_327,N_4530,N_4842);
nor UO_328 (O_328,N_4632,N_4619);
nor UO_329 (O_329,N_4884,N_4647);
nor UO_330 (O_330,N_4736,N_4788);
nor UO_331 (O_331,N_4716,N_4915);
or UO_332 (O_332,N_4707,N_4651);
nor UO_333 (O_333,N_4916,N_4528);
nand UO_334 (O_334,N_4529,N_4696);
xnor UO_335 (O_335,N_4931,N_4903);
or UO_336 (O_336,N_4787,N_4927);
nand UO_337 (O_337,N_4645,N_4839);
xnor UO_338 (O_338,N_4630,N_4890);
xnor UO_339 (O_339,N_4905,N_4574);
nor UO_340 (O_340,N_4698,N_4560);
and UO_341 (O_341,N_4666,N_4864);
and UO_342 (O_342,N_4652,N_4718);
nor UO_343 (O_343,N_4948,N_4561);
xor UO_344 (O_344,N_4972,N_4918);
and UO_345 (O_345,N_4821,N_4837);
nor UO_346 (O_346,N_4671,N_4610);
or UO_347 (O_347,N_4841,N_4500);
or UO_348 (O_348,N_4501,N_4627);
and UO_349 (O_349,N_4799,N_4916);
and UO_350 (O_350,N_4753,N_4881);
nand UO_351 (O_351,N_4876,N_4565);
nand UO_352 (O_352,N_4943,N_4512);
xnor UO_353 (O_353,N_4770,N_4578);
nand UO_354 (O_354,N_4663,N_4746);
nor UO_355 (O_355,N_4603,N_4633);
and UO_356 (O_356,N_4784,N_4987);
and UO_357 (O_357,N_4669,N_4929);
or UO_358 (O_358,N_4636,N_4716);
nand UO_359 (O_359,N_4694,N_4896);
and UO_360 (O_360,N_4781,N_4786);
and UO_361 (O_361,N_4846,N_4998);
or UO_362 (O_362,N_4956,N_4836);
nand UO_363 (O_363,N_4904,N_4712);
nor UO_364 (O_364,N_4852,N_4941);
nand UO_365 (O_365,N_4546,N_4995);
or UO_366 (O_366,N_4692,N_4625);
nor UO_367 (O_367,N_4566,N_4658);
nand UO_368 (O_368,N_4507,N_4886);
xnor UO_369 (O_369,N_4695,N_4541);
and UO_370 (O_370,N_4552,N_4537);
and UO_371 (O_371,N_4938,N_4704);
and UO_372 (O_372,N_4694,N_4631);
and UO_373 (O_373,N_4680,N_4731);
nand UO_374 (O_374,N_4842,N_4690);
or UO_375 (O_375,N_4990,N_4666);
and UO_376 (O_376,N_4815,N_4911);
and UO_377 (O_377,N_4569,N_4735);
and UO_378 (O_378,N_4835,N_4640);
and UO_379 (O_379,N_4662,N_4772);
nand UO_380 (O_380,N_4744,N_4739);
nand UO_381 (O_381,N_4766,N_4750);
nor UO_382 (O_382,N_4924,N_4584);
and UO_383 (O_383,N_4595,N_4587);
xnor UO_384 (O_384,N_4943,N_4604);
or UO_385 (O_385,N_4730,N_4641);
or UO_386 (O_386,N_4751,N_4794);
or UO_387 (O_387,N_4650,N_4787);
nor UO_388 (O_388,N_4755,N_4904);
nor UO_389 (O_389,N_4508,N_4728);
nor UO_390 (O_390,N_4676,N_4853);
and UO_391 (O_391,N_4807,N_4842);
nand UO_392 (O_392,N_4685,N_4808);
or UO_393 (O_393,N_4626,N_4816);
or UO_394 (O_394,N_4714,N_4598);
and UO_395 (O_395,N_4743,N_4599);
nor UO_396 (O_396,N_4729,N_4908);
nand UO_397 (O_397,N_4601,N_4964);
nor UO_398 (O_398,N_4660,N_4518);
or UO_399 (O_399,N_4881,N_4723);
nand UO_400 (O_400,N_4754,N_4758);
and UO_401 (O_401,N_4845,N_4542);
nor UO_402 (O_402,N_4783,N_4935);
or UO_403 (O_403,N_4608,N_4840);
nand UO_404 (O_404,N_4570,N_4926);
nand UO_405 (O_405,N_4568,N_4627);
and UO_406 (O_406,N_4574,N_4761);
or UO_407 (O_407,N_4651,N_4713);
nor UO_408 (O_408,N_4849,N_4703);
and UO_409 (O_409,N_4912,N_4532);
nand UO_410 (O_410,N_4637,N_4890);
nand UO_411 (O_411,N_4930,N_4675);
or UO_412 (O_412,N_4602,N_4807);
and UO_413 (O_413,N_4978,N_4647);
and UO_414 (O_414,N_4602,N_4663);
nand UO_415 (O_415,N_4654,N_4538);
and UO_416 (O_416,N_4765,N_4845);
or UO_417 (O_417,N_4577,N_4754);
or UO_418 (O_418,N_4846,N_4514);
and UO_419 (O_419,N_4892,N_4678);
nand UO_420 (O_420,N_4983,N_4651);
nor UO_421 (O_421,N_4743,N_4870);
or UO_422 (O_422,N_4833,N_4968);
nand UO_423 (O_423,N_4681,N_4908);
nand UO_424 (O_424,N_4599,N_4827);
or UO_425 (O_425,N_4539,N_4656);
and UO_426 (O_426,N_4865,N_4593);
or UO_427 (O_427,N_4884,N_4829);
or UO_428 (O_428,N_4798,N_4860);
nor UO_429 (O_429,N_4902,N_4642);
or UO_430 (O_430,N_4739,N_4849);
and UO_431 (O_431,N_4780,N_4572);
nand UO_432 (O_432,N_4717,N_4654);
and UO_433 (O_433,N_4937,N_4861);
xnor UO_434 (O_434,N_4770,N_4798);
or UO_435 (O_435,N_4827,N_4568);
or UO_436 (O_436,N_4874,N_4946);
nand UO_437 (O_437,N_4900,N_4967);
and UO_438 (O_438,N_4731,N_4949);
nor UO_439 (O_439,N_4576,N_4577);
xor UO_440 (O_440,N_4654,N_4697);
nand UO_441 (O_441,N_4762,N_4898);
xnor UO_442 (O_442,N_4662,N_4544);
nor UO_443 (O_443,N_4589,N_4789);
and UO_444 (O_444,N_4743,N_4555);
nand UO_445 (O_445,N_4584,N_4522);
nor UO_446 (O_446,N_4865,N_4794);
nand UO_447 (O_447,N_4838,N_4739);
or UO_448 (O_448,N_4737,N_4500);
nand UO_449 (O_449,N_4521,N_4745);
nand UO_450 (O_450,N_4865,N_4654);
xor UO_451 (O_451,N_4950,N_4870);
and UO_452 (O_452,N_4705,N_4659);
nor UO_453 (O_453,N_4643,N_4804);
nor UO_454 (O_454,N_4991,N_4511);
xnor UO_455 (O_455,N_4924,N_4656);
xnor UO_456 (O_456,N_4857,N_4526);
nand UO_457 (O_457,N_4692,N_4831);
or UO_458 (O_458,N_4804,N_4519);
nand UO_459 (O_459,N_4802,N_4756);
and UO_460 (O_460,N_4774,N_4580);
nor UO_461 (O_461,N_4993,N_4953);
nor UO_462 (O_462,N_4973,N_4949);
nor UO_463 (O_463,N_4630,N_4647);
nand UO_464 (O_464,N_4522,N_4603);
or UO_465 (O_465,N_4556,N_4679);
nor UO_466 (O_466,N_4790,N_4912);
nand UO_467 (O_467,N_4508,N_4684);
nor UO_468 (O_468,N_4673,N_4794);
nand UO_469 (O_469,N_4939,N_4767);
nor UO_470 (O_470,N_4743,N_4580);
nand UO_471 (O_471,N_4561,N_4865);
or UO_472 (O_472,N_4530,N_4513);
or UO_473 (O_473,N_4532,N_4659);
and UO_474 (O_474,N_4735,N_4630);
nor UO_475 (O_475,N_4580,N_4915);
nor UO_476 (O_476,N_4946,N_4627);
nor UO_477 (O_477,N_4810,N_4917);
and UO_478 (O_478,N_4694,N_4600);
and UO_479 (O_479,N_4531,N_4530);
or UO_480 (O_480,N_4934,N_4712);
nand UO_481 (O_481,N_4812,N_4794);
xor UO_482 (O_482,N_4774,N_4788);
and UO_483 (O_483,N_4588,N_4997);
and UO_484 (O_484,N_4688,N_4763);
and UO_485 (O_485,N_4768,N_4892);
nand UO_486 (O_486,N_4637,N_4675);
or UO_487 (O_487,N_4692,N_4507);
nand UO_488 (O_488,N_4791,N_4851);
or UO_489 (O_489,N_4621,N_4856);
or UO_490 (O_490,N_4769,N_4960);
or UO_491 (O_491,N_4521,N_4629);
or UO_492 (O_492,N_4980,N_4912);
nor UO_493 (O_493,N_4534,N_4682);
or UO_494 (O_494,N_4615,N_4518);
and UO_495 (O_495,N_4669,N_4858);
nand UO_496 (O_496,N_4689,N_4538);
nand UO_497 (O_497,N_4616,N_4988);
nor UO_498 (O_498,N_4859,N_4981);
and UO_499 (O_499,N_4858,N_4739);
nand UO_500 (O_500,N_4770,N_4670);
and UO_501 (O_501,N_4703,N_4788);
nor UO_502 (O_502,N_4903,N_4796);
nand UO_503 (O_503,N_4915,N_4823);
nor UO_504 (O_504,N_4585,N_4897);
nor UO_505 (O_505,N_4946,N_4680);
nor UO_506 (O_506,N_4733,N_4571);
xnor UO_507 (O_507,N_4570,N_4902);
nor UO_508 (O_508,N_4799,N_4934);
or UO_509 (O_509,N_4604,N_4915);
nor UO_510 (O_510,N_4739,N_4522);
or UO_511 (O_511,N_4808,N_4828);
or UO_512 (O_512,N_4955,N_4565);
and UO_513 (O_513,N_4583,N_4592);
nor UO_514 (O_514,N_4521,N_4987);
nor UO_515 (O_515,N_4950,N_4988);
nor UO_516 (O_516,N_4891,N_4691);
nor UO_517 (O_517,N_4864,N_4553);
nand UO_518 (O_518,N_4730,N_4939);
xnor UO_519 (O_519,N_4780,N_4744);
nor UO_520 (O_520,N_4978,N_4783);
and UO_521 (O_521,N_4739,N_4854);
or UO_522 (O_522,N_4668,N_4992);
or UO_523 (O_523,N_4916,N_4617);
nor UO_524 (O_524,N_4780,N_4509);
and UO_525 (O_525,N_4590,N_4933);
or UO_526 (O_526,N_4702,N_4943);
and UO_527 (O_527,N_4865,N_4851);
and UO_528 (O_528,N_4625,N_4934);
and UO_529 (O_529,N_4543,N_4994);
and UO_530 (O_530,N_4759,N_4848);
xnor UO_531 (O_531,N_4668,N_4592);
or UO_532 (O_532,N_4729,N_4532);
and UO_533 (O_533,N_4666,N_4897);
xor UO_534 (O_534,N_4779,N_4588);
and UO_535 (O_535,N_4502,N_4925);
or UO_536 (O_536,N_4504,N_4735);
or UO_537 (O_537,N_4647,N_4815);
nand UO_538 (O_538,N_4677,N_4606);
or UO_539 (O_539,N_4990,N_4727);
nor UO_540 (O_540,N_4620,N_4880);
nor UO_541 (O_541,N_4626,N_4759);
or UO_542 (O_542,N_4801,N_4539);
nand UO_543 (O_543,N_4758,N_4908);
nor UO_544 (O_544,N_4668,N_4885);
nor UO_545 (O_545,N_4507,N_4516);
nor UO_546 (O_546,N_4778,N_4946);
and UO_547 (O_547,N_4954,N_4771);
nand UO_548 (O_548,N_4601,N_4647);
nand UO_549 (O_549,N_4992,N_4534);
or UO_550 (O_550,N_4752,N_4561);
or UO_551 (O_551,N_4537,N_4671);
nand UO_552 (O_552,N_4959,N_4898);
nand UO_553 (O_553,N_4772,N_4951);
nand UO_554 (O_554,N_4886,N_4794);
nand UO_555 (O_555,N_4908,N_4935);
nand UO_556 (O_556,N_4896,N_4803);
and UO_557 (O_557,N_4779,N_4750);
or UO_558 (O_558,N_4820,N_4929);
and UO_559 (O_559,N_4976,N_4799);
nor UO_560 (O_560,N_4557,N_4923);
nand UO_561 (O_561,N_4733,N_4888);
nand UO_562 (O_562,N_4835,N_4749);
and UO_563 (O_563,N_4966,N_4878);
nand UO_564 (O_564,N_4748,N_4634);
and UO_565 (O_565,N_4840,N_4567);
nor UO_566 (O_566,N_4609,N_4623);
nand UO_567 (O_567,N_4618,N_4665);
nand UO_568 (O_568,N_4800,N_4609);
nand UO_569 (O_569,N_4919,N_4844);
nor UO_570 (O_570,N_4940,N_4989);
or UO_571 (O_571,N_4561,N_4936);
nand UO_572 (O_572,N_4818,N_4878);
xor UO_573 (O_573,N_4966,N_4525);
nor UO_574 (O_574,N_4879,N_4949);
nor UO_575 (O_575,N_4603,N_4671);
and UO_576 (O_576,N_4745,N_4828);
and UO_577 (O_577,N_4764,N_4718);
or UO_578 (O_578,N_4913,N_4777);
or UO_579 (O_579,N_4940,N_4872);
or UO_580 (O_580,N_4738,N_4980);
nand UO_581 (O_581,N_4629,N_4612);
nand UO_582 (O_582,N_4729,N_4809);
nand UO_583 (O_583,N_4905,N_4597);
nand UO_584 (O_584,N_4528,N_4641);
nor UO_585 (O_585,N_4507,N_4836);
xnor UO_586 (O_586,N_4749,N_4686);
nor UO_587 (O_587,N_4986,N_4696);
or UO_588 (O_588,N_4941,N_4752);
nor UO_589 (O_589,N_4901,N_4842);
and UO_590 (O_590,N_4812,N_4604);
xnor UO_591 (O_591,N_4650,N_4967);
nand UO_592 (O_592,N_4809,N_4619);
nor UO_593 (O_593,N_4972,N_4642);
or UO_594 (O_594,N_4706,N_4895);
xnor UO_595 (O_595,N_4816,N_4908);
nor UO_596 (O_596,N_4552,N_4762);
nor UO_597 (O_597,N_4822,N_4899);
and UO_598 (O_598,N_4574,N_4728);
and UO_599 (O_599,N_4910,N_4674);
nand UO_600 (O_600,N_4618,N_4573);
and UO_601 (O_601,N_4930,N_4998);
xor UO_602 (O_602,N_4899,N_4621);
xnor UO_603 (O_603,N_4815,N_4719);
nor UO_604 (O_604,N_4657,N_4537);
or UO_605 (O_605,N_4960,N_4640);
or UO_606 (O_606,N_4788,N_4964);
nand UO_607 (O_607,N_4687,N_4722);
nor UO_608 (O_608,N_4839,N_4545);
and UO_609 (O_609,N_4742,N_4893);
or UO_610 (O_610,N_4693,N_4569);
or UO_611 (O_611,N_4961,N_4996);
nor UO_612 (O_612,N_4863,N_4591);
and UO_613 (O_613,N_4741,N_4659);
nand UO_614 (O_614,N_4558,N_4747);
or UO_615 (O_615,N_4658,N_4883);
and UO_616 (O_616,N_4915,N_4632);
and UO_617 (O_617,N_4810,N_4650);
or UO_618 (O_618,N_4830,N_4943);
and UO_619 (O_619,N_4551,N_4683);
or UO_620 (O_620,N_4791,N_4908);
and UO_621 (O_621,N_4980,N_4742);
nand UO_622 (O_622,N_4630,N_4562);
or UO_623 (O_623,N_4816,N_4666);
and UO_624 (O_624,N_4732,N_4555);
nor UO_625 (O_625,N_4822,N_4686);
nand UO_626 (O_626,N_4655,N_4660);
and UO_627 (O_627,N_4900,N_4806);
xnor UO_628 (O_628,N_4680,N_4514);
nand UO_629 (O_629,N_4502,N_4820);
or UO_630 (O_630,N_4778,N_4505);
or UO_631 (O_631,N_4644,N_4512);
and UO_632 (O_632,N_4516,N_4533);
and UO_633 (O_633,N_4890,N_4638);
nor UO_634 (O_634,N_4825,N_4681);
and UO_635 (O_635,N_4765,N_4507);
nor UO_636 (O_636,N_4901,N_4766);
nand UO_637 (O_637,N_4697,N_4582);
or UO_638 (O_638,N_4986,N_4605);
or UO_639 (O_639,N_4751,N_4715);
or UO_640 (O_640,N_4740,N_4639);
and UO_641 (O_641,N_4599,N_4874);
nand UO_642 (O_642,N_4641,N_4551);
nor UO_643 (O_643,N_4986,N_4586);
xnor UO_644 (O_644,N_4957,N_4807);
nor UO_645 (O_645,N_4698,N_4757);
and UO_646 (O_646,N_4796,N_4952);
or UO_647 (O_647,N_4548,N_4835);
nand UO_648 (O_648,N_4882,N_4653);
nor UO_649 (O_649,N_4608,N_4905);
or UO_650 (O_650,N_4537,N_4843);
or UO_651 (O_651,N_4610,N_4698);
or UO_652 (O_652,N_4501,N_4664);
nor UO_653 (O_653,N_4753,N_4563);
nor UO_654 (O_654,N_4802,N_4582);
and UO_655 (O_655,N_4938,N_4688);
and UO_656 (O_656,N_4508,N_4588);
and UO_657 (O_657,N_4932,N_4918);
xor UO_658 (O_658,N_4761,N_4897);
and UO_659 (O_659,N_4688,N_4739);
xor UO_660 (O_660,N_4848,N_4607);
or UO_661 (O_661,N_4796,N_4677);
or UO_662 (O_662,N_4562,N_4624);
or UO_663 (O_663,N_4566,N_4889);
nand UO_664 (O_664,N_4790,N_4874);
or UO_665 (O_665,N_4638,N_4573);
and UO_666 (O_666,N_4828,N_4926);
nor UO_667 (O_667,N_4832,N_4662);
and UO_668 (O_668,N_4962,N_4627);
or UO_669 (O_669,N_4684,N_4516);
or UO_670 (O_670,N_4542,N_4799);
nand UO_671 (O_671,N_4717,N_4601);
xor UO_672 (O_672,N_4767,N_4676);
nand UO_673 (O_673,N_4945,N_4601);
or UO_674 (O_674,N_4652,N_4773);
nand UO_675 (O_675,N_4794,N_4731);
or UO_676 (O_676,N_4992,N_4847);
or UO_677 (O_677,N_4525,N_4731);
nor UO_678 (O_678,N_4736,N_4886);
and UO_679 (O_679,N_4985,N_4593);
and UO_680 (O_680,N_4755,N_4589);
or UO_681 (O_681,N_4694,N_4547);
nor UO_682 (O_682,N_4701,N_4844);
nand UO_683 (O_683,N_4703,N_4697);
nand UO_684 (O_684,N_4699,N_4934);
nand UO_685 (O_685,N_4723,N_4724);
nand UO_686 (O_686,N_4582,N_4816);
nor UO_687 (O_687,N_4980,N_4614);
nand UO_688 (O_688,N_4939,N_4544);
nor UO_689 (O_689,N_4998,N_4675);
xnor UO_690 (O_690,N_4608,N_4967);
or UO_691 (O_691,N_4896,N_4596);
or UO_692 (O_692,N_4743,N_4736);
xor UO_693 (O_693,N_4777,N_4810);
xnor UO_694 (O_694,N_4928,N_4745);
and UO_695 (O_695,N_4988,N_4894);
or UO_696 (O_696,N_4648,N_4672);
or UO_697 (O_697,N_4902,N_4805);
xor UO_698 (O_698,N_4992,N_4865);
nand UO_699 (O_699,N_4523,N_4669);
nand UO_700 (O_700,N_4783,N_4545);
nand UO_701 (O_701,N_4911,N_4865);
nand UO_702 (O_702,N_4899,N_4994);
nand UO_703 (O_703,N_4985,N_4571);
nor UO_704 (O_704,N_4781,N_4840);
and UO_705 (O_705,N_4677,N_4716);
nor UO_706 (O_706,N_4805,N_4924);
or UO_707 (O_707,N_4767,N_4982);
nor UO_708 (O_708,N_4526,N_4641);
and UO_709 (O_709,N_4989,N_4795);
nor UO_710 (O_710,N_4682,N_4760);
nor UO_711 (O_711,N_4588,N_4826);
and UO_712 (O_712,N_4774,N_4744);
or UO_713 (O_713,N_4711,N_4626);
and UO_714 (O_714,N_4627,N_4706);
and UO_715 (O_715,N_4533,N_4537);
nor UO_716 (O_716,N_4971,N_4724);
and UO_717 (O_717,N_4907,N_4873);
and UO_718 (O_718,N_4715,N_4938);
xnor UO_719 (O_719,N_4701,N_4850);
xor UO_720 (O_720,N_4578,N_4653);
nand UO_721 (O_721,N_4702,N_4768);
or UO_722 (O_722,N_4763,N_4958);
nand UO_723 (O_723,N_4980,N_4536);
or UO_724 (O_724,N_4893,N_4764);
nand UO_725 (O_725,N_4783,N_4593);
nor UO_726 (O_726,N_4617,N_4610);
nand UO_727 (O_727,N_4782,N_4770);
nand UO_728 (O_728,N_4749,N_4699);
and UO_729 (O_729,N_4850,N_4640);
xor UO_730 (O_730,N_4880,N_4953);
nand UO_731 (O_731,N_4639,N_4875);
and UO_732 (O_732,N_4931,N_4905);
or UO_733 (O_733,N_4534,N_4637);
or UO_734 (O_734,N_4754,N_4759);
nand UO_735 (O_735,N_4933,N_4737);
nor UO_736 (O_736,N_4851,N_4741);
xor UO_737 (O_737,N_4547,N_4647);
nand UO_738 (O_738,N_4861,N_4916);
nor UO_739 (O_739,N_4792,N_4520);
xnor UO_740 (O_740,N_4597,N_4939);
nand UO_741 (O_741,N_4823,N_4944);
nor UO_742 (O_742,N_4968,N_4565);
nand UO_743 (O_743,N_4559,N_4609);
nand UO_744 (O_744,N_4563,N_4820);
and UO_745 (O_745,N_4813,N_4910);
xor UO_746 (O_746,N_4535,N_4864);
or UO_747 (O_747,N_4644,N_4998);
nor UO_748 (O_748,N_4616,N_4955);
or UO_749 (O_749,N_4566,N_4691);
and UO_750 (O_750,N_4639,N_4595);
and UO_751 (O_751,N_4520,N_4596);
and UO_752 (O_752,N_4810,N_4824);
or UO_753 (O_753,N_4564,N_4976);
nor UO_754 (O_754,N_4825,N_4909);
or UO_755 (O_755,N_4905,N_4526);
or UO_756 (O_756,N_4599,N_4558);
nand UO_757 (O_757,N_4627,N_4503);
or UO_758 (O_758,N_4606,N_4599);
and UO_759 (O_759,N_4939,N_4567);
nor UO_760 (O_760,N_4617,N_4547);
nor UO_761 (O_761,N_4808,N_4672);
xnor UO_762 (O_762,N_4681,N_4891);
and UO_763 (O_763,N_4806,N_4638);
nor UO_764 (O_764,N_4900,N_4590);
or UO_765 (O_765,N_4774,N_4566);
nand UO_766 (O_766,N_4807,N_4877);
or UO_767 (O_767,N_4866,N_4878);
or UO_768 (O_768,N_4740,N_4847);
xnor UO_769 (O_769,N_4798,N_4938);
and UO_770 (O_770,N_4606,N_4736);
or UO_771 (O_771,N_4958,N_4813);
xnor UO_772 (O_772,N_4576,N_4870);
nor UO_773 (O_773,N_4561,N_4877);
and UO_774 (O_774,N_4939,N_4614);
nor UO_775 (O_775,N_4711,N_4746);
or UO_776 (O_776,N_4966,N_4640);
or UO_777 (O_777,N_4864,N_4885);
or UO_778 (O_778,N_4512,N_4738);
nand UO_779 (O_779,N_4867,N_4649);
nor UO_780 (O_780,N_4915,N_4670);
xnor UO_781 (O_781,N_4774,N_4782);
or UO_782 (O_782,N_4899,N_4650);
and UO_783 (O_783,N_4565,N_4800);
xor UO_784 (O_784,N_4526,N_4503);
xnor UO_785 (O_785,N_4566,N_4627);
nor UO_786 (O_786,N_4627,N_4912);
nand UO_787 (O_787,N_4847,N_4689);
and UO_788 (O_788,N_4788,N_4709);
nand UO_789 (O_789,N_4657,N_4796);
and UO_790 (O_790,N_4736,N_4644);
and UO_791 (O_791,N_4896,N_4953);
xnor UO_792 (O_792,N_4844,N_4991);
xnor UO_793 (O_793,N_4975,N_4763);
nor UO_794 (O_794,N_4713,N_4761);
nor UO_795 (O_795,N_4574,N_4706);
or UO_796 (O_796,N_4973,N_4666);
nor UO_797 (O_797,N_4566,N_4642);
and UO_798 (O_798,N_4616,N_4537);
and UO_799 (O_799,N_4766,N_4601);
or UO_800 (O_800,N_4666,N_4887);
and UO_801 (O_801,N_4581,N_4844);
or UO_802 (O_802,N_4812,N_4519);
xnor UO_803 (O_803,N_4665,N_4979);
or UO_804 (O_804,N_4837,N_4966);
xnor UO_805 (O_805,N_4694,N_4582);
and UO_806 (O_806,N_4621,N_4875);
nor UO_807 (O_807,N_4922,N_4820);
or UO_808 (O_808,N_4690,N_4664);
nor UO_809 (O_809,N_4934,N_4589);
or UO_810 (O_810,N_4986,N_4723);
and UO_811 (O_811,N_4700,N_4817);
and UO_812 (O_812,N_4854,N_4979);
or UO_813 (O_813,N_4684,N_4899);
nor UO_814 (O_814,N_4676,N_4655);
nor UO_815 (O_815,N_4869,N_4927);
or UO_816 (O_816,N_4989,N_4891);
or UO_817 (O_817,N_4894,N_4774);
or UO_818 (O_818,N_4527,N_4896);
and UO_819 (O_819,N_4906,N_4836);
nand UO_820 (O_820,N_4528,N_4973);
or UO_821 (O_821,N_4968,N_4945);
and UO_822 (O_822,N_4525,N_4991);
nor UO_823 (O_823,N_4852,N_4764);
nand UO_824 (O_824,N_4732,N_4522);
xnor UO_825 (O_825,N_4512,N_4672);
and UO_826 (O_826,N_4547,N_4610);
nand UO_827 (O_827,N_4848,N_4705);
and UO_828 (O_828,N_4538,N_4843);
and UO_829 (O_829,N_4868,N_4790);
and UO_830 (O_830,N_4523,N_4521);
and UO_831 (O_831,N_4651,N_4669);
and UO_832 (O_832,N_4993,N_4848);
nor UO_833 (O_833,N_4853,N_4622);
xnor UO_834 (O_834,N_4956,N_4915);
and UO_835 (O_835,N_4613,N_4734);
or UO_836 (O_836,N_4523,N_4926);
nand UO_837 (O_837,N_4557,N_4890);
nand UO_838 (O_838,N_4573,N_4912);
nand UO_839 (O_839,N_4560,N_4581);
nor UO_840 (O_840,N_4556,N_4965);
nor UO_841 (O_841,N_4618,N_4794);
or UO_842 (O_842,N_4642,N_4999);
and UO_843 (O_843,N_4692,N_4762);
nand UO_844 (O_844,N_4965,N_4951);
nor UO_845 (O_845,N_4526,N_4727);
nand UO_846 (O_846,N_4978,N_4610);
and UO_847 (O_847,N_4629,N_4709);
xor UO_848 (O_848,N_4819,N_4575);
or UO_849 (O_849,N_4551,N_4844);
or UO_850 (O_850,N_4520,N_4950);
nor UO_851 (O_851,N_4934,N_4652);
xnor UO_852 (O_852,N_4547,N_4656);
nor UO_853 (O_853,N_4923,N_4877);
nor UO_854 (O_854,N_4623,N_4603);
nand UO_855 (O_855,N_4525,N_4750);
and UO_856 (O_856,N_4600,N_4673);
nor UO_857 (O_857,N_4974,N_4780);
nor UO_858 (O_858,N_4714,N_4800);
nor UO_859 (O_859,N_4566,N_4713);
nand UO_860 (O_860,N_4851,N_4815);
nand UO_861 (O_861,N_4519,N_4624);
nor UO_862 (O_862,N_4511,N_4813);
or UO_863 (O_863,N_4756,N_4769);
and UO_864 (O_864,N_4816,N_4704);
and UO_865 (O_865,N_4948,N_4981);
or UO_866 (O_866,N_4624,N_4614);
nor UO_867 (O_867,N_4510,N_4633);
nand UO_868 (O_868,N_4569,N_4972);
or UO_869 (O_869,N_4747,N_4841);
or UO_870 (O_870,N_4525,N_4819);
nand UO_871 (O_871,N_4772,N_4529);
and UO_872 (O_872,N_4594,N_4824);
nand UO_873 (O_873,N_4990,N_4758);
nand UO_874 (O_874,N_4543,N_4740);
or UO_875 (O_875,N_4565,N_4996);
or UO_876 (O_876,N_4526,N_4700);
nor UO_877 (O_877,N_4809,N_4907);
nor UO_878 (O_878,N_4686,N_4607);
nor UO_879 (O_879,N_4737,N_4604);
nor UO_880 (O_880,N_4641,N_4575);
or UO_881 (O_881,N_4971,N_4695);
nor UO_882 (O_882,N_4840,N_4547);
xor UO_883 (O_883,N_4921,N_4637);
or UO_884 (O_884,N_4756,N_4623);
and UO_885 (O_885,N_4830,N_4701);
xor UO_886 (O_886,N_4982,N_4985);
nor UO_887 (O_887,N_4510,N_4677);
nand UO_888 (O_888,N_4626,N_4717);
nor UO_889 (O_889,N_4549,N_4845);
nand UO_890 (O_890,N_4600,N_4718);
and UO_891 (O_891,N_4865,N_4515);
and UO_892 (O_892,N_4843,N_4506);
nand UO_893 (O_893,N_4556,N_4721);
nor UO_894 (O_894,N_4936,N_4904);
or UO_895 (O_895,N_4765,N_4544);
nor UO_896 (O_896,N_4554,N_4578);
nor UO_897 (O_897,N_4510,N_4994);
and UO_898 (O_898,N_4530,N_4651);
nor UO_899 (O_899,N_4887,N_4584);
xor UO_900 (O_900,N_4608,N_4628);
nor UO_901 (O_901,N_4641,N_4642);
nor UO_902 (O_902,N_4506,N_4980);
nor UO_903 (O_903,N_4935,N_4723);
and UO_904 (O_904,N_4539,N_4891);
and UO_905 (O_905,N_4672,N_4872);
nor UO_906 (O_906,N_4559,N_4600);
and UO_907 (O_907,N_4817,N_4784);
or UO_908 (O_908,N_4925,N_4857);
or UO_909 (O_909,N_4933,N_4514);
nor UO_910 (O_910,N_4834,N_4566);
nand UO_911 (O_911,N_4592,N_4541);
nand UO_912 (O_912,N_4856,N_4697);
nand UO_913 (O_913,N_4923,N_4677);
and UO_914 (O_914,N_4698,N_4533);
or UO_915 (O_915,N_4533,N_4637);
nand UO_916 (O_916,N_4851,N_4620);
nand UO_917 (O_917,N_4911,N_4775);
nor UO_918 (O_918,N_4719,N_4936);
or UO_919 (O_919,N_4727,N_4547);
nor UO_920 (O_920,N_4777,N_4573);
or UO_921 (O_921,N_4525,N_4685);
or UO_922 (O_922,N_4921,N_4536);
nor UO_923 (O_923,N_4999,N_4721);
nor UO_924 (O_924,N_4695,N_4614);
and UO_925 (O_925,N_4816,N_4885);
nor UO_926 (O_926,N_4524,N_4620);
nand UO_927 (O_927,N_4796,N_4697);
nand UO_928 (O_928,N_4603,N_4704);
nand UO_929 (O_929,N_4899,N_4706);
or UO_930 (O_930,N_4987,N_4813);
xor UO_931 (O_931,N_4864,N_4579);
nor UO_932 (O_932,N_4544,N_4730);
xor UO_933 (O_933,N_4891,N_4629);
nor UO_934 (O_934,N_4877,N_4759);
nor UO_935 (O_935,N_4907,N_4581);
xor UO_936 (O_936,N_4631,N_4716);
nand UO_937 (O_937,N_4604,N_4597);
and UO_938 (O_938,N_4612,N_4665);
nand UO_939 (O_939,N_4968,N_4823);
nor UO_940 (O_940,N_4571,N_4526);
nand UO_941 (O_941,N_4989,N_4863);
nand UO_942 (O_942,N_4659,N_4815);
and UO_943 (O_943,N_4982,N_4562);
and UO_944 (O_944,N_4810,N_4721);
or UO_945 (O_945,N_4628,N_4813);
nand UO_946 (O_946,N_4709,N_4866);
nor UO_947 (O_947,N_4644,N_4873);
nor UO_948 (O_948,N_4789,N_4959);
and UO_949 (O_949,N_4896,N_4797);
or UO_950 (O_950,N_4539,N_4724);
and UO_951 (O_951,N_4873,N_4738);
xor UO_952 (O_952,N_4677,N_4595);
or UO_953 (O_953,N_4552,N_4934);
and UO_954 (O_954,N_4763,N_4841);
nor UO_955 (O_955,N_4592,N_4797);
nor UO_956 (O_956,N_4807,N_4736);
nand UO_957 (O_957,N_4807,N_4539);
and UO_958 (O_958,N_4674,N_4950);
and UO_959 (O_959,N_4645,N_4699);
nor UO_960 (O_960,N_4562,N_4858);
xor UO_961 (O_961,N_4764,N_4581);
nand UO_962 (O_962,N_4798,N_4538);
xor UO_963 (O_963,N_4814,N_4859);
or UO_964 (O_964,N_4788,N_4847);
nand UO_965 (O_965,N_4710,N_4940);
nand UO_966 (O_966,N_4822,N_4736);
xnor UO_967 (O_967,N_4943,N_4866);
and UO_968 (O_968,N_4868,N_4627);
nor UO_969 (O_969,N_4963,N_4896);
or UO_970 (O_970,N_4841,N_4811);
and UO_971 (O_971,N_4687,N_4912);
and UO_972 (O_972,N_4616,N_4551);
or UO_973 (O_973,N_4969,N_4840);
and UO_974 (O_974,N_4653,N_4690);
or UO_975 (O_975,N_4625,N_4974);
nor UO_976 (O_976,N_4741,N_4725);
xnor UO_977 (O_977,N_4652,N_4937);
xnor UO_978 (O_978,N_4780,N_4669);
and UO_979 (O_979,N_4774,N_4869);
or UO_980 (O_980,N_4980,N_4674);
nand UO_981 (O_981,N_4969,N_4824);
nand UO_982 (O_982,N_4544,N_4978);
nand UO_983 (O_983,N_4557,N_4865);
nor UO_984 (O_984,N_4804,N_4722);
or UO_985 (O_985,N_4666,N_4695);
nand UO_986 (O_986,N_4696,N_4566);
nand UO_987 (O_987,N_4539,N_4549);
or UO_988 (O_988,N_4636,N_4540);
nor UO_989 (O_989,N_4638,N_4907);
or UO_990 (O_990,N_4609,N_4588);
nor UO_991 (O_991,N_4569,N_4702);
nor UO_992 (O_992,N_4823,N_4744);
or UO_993 (O_993,N_4509,N_4805);
or UO_994 (O_994,N_4837,N_4539);
nor UO_995 (O_995,N_4830,N_4751);
and UO_996 (O_996,N_4858,N_4744);
nor UO_997 (O_997,N_4508,N_4829);
and UO_998 (O_998,N_4841,N_4973);
nand UO_999 (O_999,N_4871,N_4933);
endmodule