module basic_500_3000_500_30_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_25,In_411);
nand U1 (N_1,In_284,In_405);
and U2 (N_2,In_417,In_15);
or U3 (N_3,In_480,In_76);
or U4 (N_4,In_148,In_344);
and U5 (N_5,In_464,In_376);
nor U6 (N_6,In_277,In_42);
nand U7 (N_7,In_288,In_292);
nand U8 (N_8,In_211,In_300);
and U9 (N_9,In_279,In_106);
nand U10 (N_10,In_466,In_143);
xor U11 (N_11,In_40,In_453);
nand U12 (N_12,In_227,In_334);
nor U13 (N_13,In_141,In_81);
and U14 (N_14,In_339,In_317);
xor U15 (N_15,In_66,In_351);
or U16 (N_16,In_418,In_228);
nand U17 (N_17,In_326,In_77);
xor U18 (N_18,In_73,In_119);
nand U19 (N_19,In_380,In_168);
and U20 (N_20,In_147,In_176);
or U21 (N_21,In_243,In_3);
and U22 (N_22,In_43,In_187);
and U23 (N_23,In_33,In_109);
nor U24 (N_24,In_216,In_375);
or U25 (N_25,In_322,In_205);
nand U26 (N_26,In_154,In_50);
nand U27 (N_27,In_314,In_130);
or U28 (N_28,In_414,In_285);
nor U29 (N_29,In_306,In_84);
and U30 (N_30,In_335,In_220);
or U31 (N_31,In_445,In_366);
nand U32 (N_32,In_398,In_476);
or U33 (N_33,In_194,In_37);
nor U34 (N_34,In_123,In_477);
or U35 (N_35,In_270,In_262);
nor U36 (N_36,In_175,In_49);
nand U37 (N_37,In_470,In_474);
or U38 (N_38,In_161,In_347);
and U39 (N_39,In_295,In_164);
nor U40 (N_40,In_92,In_298);
nand U41 (N_41,In_201,In_421);
or U42 (N_42,In_53,In_210);
and U43 (N_43,In_54,In_431);
or U44 (N_44,In_275,In_6);
and U45 (N_45,In_41,In_308);
nand U46 (N_46,In_125,In_19);
nand U47 (N_47,In_242,In_315);
nand U48 (N_48,In_107,In_425);
and U49 (N_49,In_134,In_459);
xnor U50 (N_50,In_393,In_221);
nand U51 (N_51,In_180,In_72);
and U52 (N_52,In_156,In_35);
or U53 (N_53,In_27,In_213);
or U54 (N_54,In_61,In_248);
nand U55 (N_55,In_124,In_135);
xnor U56 (N_56,In_360,In_118);
nor U57 (N_57,In_424,In_153);
and U58 (N_58,In_138,In_443);
nor U59 (N_59,In_172,In_79);
and U60 (N_60,In_251,In_325);
and U61 (N_61,In_426,In_223);
and U62 (N_62,In_255,In_48);
nor U63 (N_63,In_387,In_203);
nor U64 (N_64,In_450,In_94);
and U65 (N_65,In_39,In_233);
and U66 (N_66,In_30,In_212);
or U67 (N_67,In_454,In_238);
nor U68 (N_68,In_14,In_341);
or U69 (N_69,In_349,In_433);
and U70 (N_70,In_416,In_463);
and U71 (N_71,In_246,In_74);
or U72 (N_72,In_173,In_128);
nand U73 (N_73,In_448,In_139);
nor U74 (N_74,In_80,In_368);
or U75 (N_75,In_394,In_155);
nand U76 (N_76,In_367,In_407);
nor U77 (N_77,In_372,In_268);
and U78 (N_78,In_399,In_457);
and U79 (N_79,In_435,In_171);
nor U80 (N_80,In_362,In_310);
or U81 (N_81,In_202,In_420);
nand U82 (N_82,In_159,In_46);
xor U83 (N_83,In_358,In_69);
nand U84 (N_84,In_116,In_247);
and U85 (N_85,In_432,In_266);
and U86 (N_86,In_467,In_321);
and U87 (N_87,In_149,In_150);
nor U88 (N_88,In_142,In_108);
or U89 (N_89,In_185,In_490);
nor U90 (N_90,In_254,In_353);
nand U91 (N_91,In_396,In_442);
nor U92 (N_92,In_47,In_494);
nand U93 (N_93,In_70,In_458);
nand U94 (N_94,In_38,In_193);
and U95 (N_95,In_302,In_157);
or U96 (N_96,In_265,In_312);
nand U97 (N_97,In_436,In_415);
nand U98 (N_98,In_313,In_361);
nand U99 (N_99,In_191,In_258);
and U100 (N_100,In_388,In_319);
nor U101 (N_101,In_401,In_112);
or U102 (N_102,In_245,In_10);
or U103 (N_103,In_392,In_364);
or U104 (N_104,In_241,In_282);
nand U105 (N_105,In_250,In_13);
nor U106 (N_106,In_311,In_488);
nand U107 (N_107,N_16,In_437);
or U108 (N_108,In_386,N_67);
and U109 (N_109,N_75,In_34);
nor U110 (N_110,In_182,N_65);
nand U111 (N_111,In_32,In_391);
xor U112 (N_112,In_163,In_413);
nor U113 (N_113,N_28,N_29);
nor U114 (N_114,In_338,In_9);
or U115 (N_115,In_440,In_498);
nor U116 (N_116,N_27,In_460);
nand U117 (N_117,N_38,In_115);
and U118 (N_118,In_439,In_110);
or U119 (N_119,N_76,In_271);
and U120 (N_120,N_30,In_198);
nand U121 (N_121,N_3,In_103);
and U122 (N_122,N_5,In_299);
nor U123 (N_123,In_165,N_62);
nand U124 (N_124,In_96,In_309);
or U125 (N_125,In_177,In_354);
nor U126 (N_126,In_447,N_54);
and U127 (N_127,N_74,In_408);
nor U128 (N_128,In_126,In_215);
nor U129 (N_129,In_256,N_24);
and U130 (N_130,In_52,In_479);
nand U131 (N_131,In_499,N_1);
xnor U132 (N_132,In_471,In_8);
nor U133 (N_133,In_59,N_97);
xor U134 (N_134,In_11,N_23);
or U135 (N_135,In_412,N_39);
or U136 (N_136,N_70,In_320);
nand U137 (N_137,In_140,In_287);
nor U138 (N_138,In_296,In_166);
nand U139 (N_139,In_276,In_1);
or U140 (N_140,In_5,In_345);
nand U141 (N_141,N_87,In_356);
and U142 (N_142,In_493,In_289);
or U143 (N_143,In_18,N_48);
and U144 (N_144,In_26,In_224);
and U145 (N_145,In_225,N_69);
and U146 (N_146,In_145,In_465);
or U147 (N_147,In_68,In_133);
or U148 (N_148,In_269,N_46);
nor U149 (N_149,In_263,In_170);
nor U150 (N_150,In_430,N_25);
nand U151 (N_151,In_23,In_350);
nor U152 (N_152,N_47,In_87);
nor U153 (N_153,In_239,In_487);
nand U154 (N_154,In_272,In_62);
or U155 (N_155,In_273,In_146);
and U156 (N_156,In_99,In_200);
or U157 (N_157,In_267,In_117);
nand U158 (N_158,In_348,N_4);
nand U159 (N_159,In_91,N_94);
and U160 (N_160,N_66,In_483);
or U161 (N_161,In_259,N_99);
nor U162 (N_162,In_144,In_136);
or U163 (N_163,In_264,In_88);
or U164 (N_164,N_6,N_59);
nand U165 (N_165,In_304,In_206);
or U166 (N_166,N_8,N_82);
nand U167 (N_167,In_17,In_207);
xnor U168 (N_168,In_281,In_199);
nor U169 (N_169,N_71,In_31);
and U170 (N_170,In_357,In_98);
nand U171 (N_171,In_485,N_53);
nor U172 (N_172,N_21,In_446);
or U173 (N_173,In_363,N_19);
nand U174 (N_174,In_359,In_369);
nand U175 (N_175,In_90,In_340);
nor U176 (N_176,N_33,In_461);
nor U177 (N_177,In_374,In_229);
or U178 (N_178,In_379,N_17);
nand U179 (N_179,In_331,In_86);
nand U180 (N_180,In_137,In_419);
or U181 (N_181,In_462,In_169);
and U182 (N_182,In_378,In_371);
and U183 (N_183,In_236,In_337);
nor U184 (N_184,In_290,N_72);
and U185 (N_185,In_58,In_484);
nand U186 (N_186,N_44,N_51);
and U187 (N_187,N_79,In_4);
nand U188 (N_188,In_129,N_7);
nand U189 (N_189,In_324,N_34);
nor U190 (N_190,In_97,In_283);
nor U191 (N_191,In_218,In_397);
nor U192 (N_192,In_7,N_93);
nand U193 (N_193,N_61,In_410);
and U194 (N_194,In_56,In_162);
nand U195 (N_195,In_252,In_482);
or U196 (N_196,N_88,In_102);
nand U197 (N_197,N_40,In_469);
nor U198 (N_198,In_44,In_196);
or U199 (N_199,N_58,In_131);
nand U200 (N_200,N_184,In_179);
and U201 (N_201,In_83,In_293);
nand U202 (N_202,In_71,N_18);
and U203 (N_203,N_180,In_22);
and U204 (N_204,N_193,N_140);
nand U205 (N_205,N_122,In_342);
nor U206 (N_206,N_121,N_116);
nor U207 (N_207,N_77,In_45);
nand U208 (N_208,N_176,N_114);
and U209 (N_209,N_138,In_231);
nor U210 (N_210,N_183,N_113);
nand U211 (N_211,N_15,In_24);
nor U212 (N_212,In_301,In_55);
xnor U213 (N_213,N_106,N_98);
or U214 (N_214,In_100,In_127);
and U215 (N_215,In_114,N_90);
or U216 (N_216,In_303,In_323);
nor U217 (N_217,In_385,In_189);
and U218 (N_218,In_455,N_56);
or U219 (N_219,N_150,N_172);
and U220 (N_220,In_452,In_332);
nor U221 (N_221,In_261,N_186);
nand U222 (N_222,N_42,In_217);
nor U223 (N_223,N_104,In_473);
and U224 (N_224,In_132,N_152);
nor U225 (N_225,N_12,N_156);
or U226 (N_226,In_370,In_174);
and U227 (N_227,N_117,In_151);
nor U228 (N_228,In_492,N_195);
nand U229 (N_229,N_101,In_355);
and U230 (N_230,In_186,In_65);
nor U231 (N_231,In_104,N_142);
nand U232 (N_232,In_120,N_145);
and U233 (N_233,N_128,N_49);
nand U234 (N_234,N_89,N_153);
or U235 (N_235,N_134,In_409);
or U236 (N_236,In_226,N_95);
nand U237 (N_237,In_330,N_102);
and U238 (N_238,In_346,N_2);
nand U239 (N_239,N_194,In_28);
or U240 (N_240,N_112,In_297);
nand U241 (N_241,In_51,N_32);
and U242 (N_242,N_111,N_73);
or U243 (N_243,N_120,N_115);
xor U244 (N_244,N_100,In_390);
nand U245 (N_245,N_37,N_86);
or U246 (N_246,In_307,In_286);
nand U247 (N_247,N_43,N_9);
nor U248 (N_248,N_173,N_132);
or U249 (N_249,N_14,In_497);
or U250 (N_250,In_152,N_164);
or U251 (N_251,N_36,In_197);
nand U252 (N_252,N_149,N_160);
nor U253 (N_253,In_384,In_456);
nor U254 (N_254,In_101,In_36);
nor U255 (N_255,N_170,In_472);
and U256 (N_256,N_158,In_82);
and U257 (N_257,N_133,In_381);
nand U258 (N_258,N_91,In_428);
or U259 (N_259,N_159,N_192);
or U260 (N_260,N_80,In_328);
nand U261 (N_261,In_204,In_232);
nor U262 (N_262,In_111,In_333);
or U263 (N_263,In_475,In_327);
nor U264 (N_264,N_26,In_160);
nor U265 (N_265,N_126,N_41);
nor U266 (N_266,N_189,In_294);
nand U267 (N_267,In_89,In_373);
or U268 (N_268,In_240,In_318);
or U269 (N_269,N_105,In_316);
and U270 (N_270,N_125,N_130);
and U271 (N_271,In_237,In_395);
or U272 (N_272,N_68,N_139);
xnor U273 (N_273,In_400,N_135);
nand U274 (N_274,N_141,N_78);
nor U275 (N_275,In_21,In_57);
and U276 (N_276,N_161,N_50);
nand U277 (N_277,N_148,In_178);
or U278 (N_278,In_234,In_489);
nor U279 (N_279,In_444,In_244);
or U280 (N_280,In_260,In_190);
and U281 (N_281,In_78,N_157);
nand U282 (N_282,N_109,N_31);
nor U283 (N_283,N_185,N_22);
nor U284 (N_284,N_143,N_196);
or U285 (N_285,N_0,In_377);
and U286 (N_286,In_16,In_222);
nand U287 (N_287,In_122,In_105);
or U288 (N_288,N_103,In_438);
nor U289 (N_289,N_85,N_167);
nand U290 (N_290,In_478,N_124);
or U291 (N_291,N_10,N_147);
or U292 (N_292,N_63,N_197);
nor U293 (N_293,In_280,In_402);
nor U294 (N_294,In_404,N_165);
nor U295 (N_295,N_13,N_182);
nand U296 (N_296,In_491,N_64);
or U297 (N_297,In_208,In_181);
nand U298 (N_298,N_174,In_121);
and U299 (N_299,In_486,In_365);
nor U300 (N_300,N_218,In_257);
nor U301 (N_301,N_212,N_222);
or U302 (N_302,In_60,N_119);
or U303 (N_303,N_276,N_244);
or U304 (N_304,In_441,N_299);
nand U305 (N_305,N_281,N_206);
and U306 (N_306,N_155,N_203);
or U307 (N_307,In_496,N_187);
and U308 (N_308,N_283,N_110);
nor U309 (N_309,N_294,N_209);
or U310 (N_310,In_209,In_468);
xnor U311 (N_311,N_191,N_55);
nand U312 (N_312,N_265,N_293);
nand U313 (N_313,In_427,N_127);
and U314 (N_314,In_167,N_259);
and U315 (N_315,N_228,In_188);
and U316 (N_316,In_219,N_200);
nor U317 (N_317,In_423,N_254);
or U318 (N_318,N_279,N_181);
nand U319 (N_319,N_237,In_2);
nor U320 (N_320,N_96,In_113);
nand U321 (N_321,N_235,N_248);
nor U322 (N_322,N_154,N_256);
or U323 (N_323,N_224,N_163);
nand U324 (N_324,In_383,N_136);
and U325 (N_325,N_213,N_271);
or U326 (N_326,N_108,In_451);
nand U327 (N_327,N_231,N_57);
xnor U328 (N_328,N_190,N_60);
or U329 (N_329,In_305,In_329);
nor U330 (N_330,N_123,N_52);
nand U331 (N_331,N_251,In_192);
nor U332 (N_332,In_29,In_95);
nand U333 (N_333,N_291,In_195);
nand U334 (N_334,N_83,N_286);
or U335 (N_335,N_277,N_284);
or U336 (N_336,N_233,N_211);
and U337 (N_337,In_67,N_177);
and U338 (N_338,N_168,N_246);
and U339 (N_339,N_290,N_296);
nand U340 (N_340,N_226,N_287);
and U341 (N_341,In_481,N_255);
nor U342 (N_342,N_236,N_297);
nor U343 (N_343,N_207,N_260);
and U344 (N_344,N_131,N_266);
or U345 (N_345,In_85,N_229);
or U346 (N_346,N_253,In_389);
nand U347 (N_347,In_336,N_84);
nor U348 (N_348,N_227,N_238);
nor U349 (N_349,N_282,N_234);
nor U350 (N_350,N_241,N_289);
or U351 (N_351,N_81,In_291);
nor U352 (N_352,N_179,N_146);
or U353 (N_353,N_239,N_274);
nor U354 (N_354,N_295,In_235);
and U355 (N_355,N_35,N_270);
and U356 (N_356,In_406,N_166);
nand U357 (N_357,N_245,N_240);
or U358 (N_358,N_217,N_118);
nand U359 (N_359,N_257,In_20);
nor U360 (N_360,N_178,N_129);
and U361 (N_361,N_249,N_201);
and U362 (N_362,In_249,N_285);
nor U363 (N_363,N_247,N_45);
and U364 (N_364,In_495,N_264);
and U365 (N_365,In_93,N_292);
xnor U366 (N_366,In_422,N_263);
or U367 (N_367,N_107,N_220);
nand U368 (N_368,N_92,N_198);
or U369 (N_369,N_204,N_221);
nor U370 (N_370,N_215,N_275);
nand U371 (N_371,In_214,N_225);
nor U372 (N_372,In_278,N_223);
nor U373 (N_373,In_352,In_230);
nor U374 (N_374,N_243,In_0);
nor U375 (N_375,In_403,In_343);
or U376 (N_376,N_216,N_202);
nor U377 (N_377,N_162,N_11);
or U378 (N_378,N_298,N_151);
nor U379 (N_379,N_268,N_175);
nor U380 (N_380,N_169,In_274);
or U381 (N_381,In_429,In_75);
nor U382 (N_382,In_184,In_449);
xor U383 (N_383,N_278,N_261);
nand U384 (N_384,In_434,In_253);
or U385 (N_385,N_252,N_144);
nand U386 (N_386,N_250,In_63);
nand U387 (N_387,N_232,N_219);
nand U388 (N_388,N_214,N_273);
nor U389 (N_389,N_272,N_258);
and U390 (N_390,In_183,N_20);
nand U391 (N_391,N_242,N_210);
and U392 (N_392,N_199,N_137);
nand U393 (N_393,In_64,In_158);
nand U394 (N_394,N_280,N_262);
and U395 (N_395,N_230,N_208);
nand U396 (N_396,In_382,N_267);
and U397 (N_397,N_188,N_269);
nand U398 (N_398,N_205,In_12);
and U399 (N_399,N_171,N_288);
nand U400 (N_400,N_383,N_397);
nor U401 (N_401,N_396,N_309);
nor U402 (N_402,N_315,N_323);
and U403 (N_403,N_357,N_359);
and U404 (N_404,N_342,N_364);
nor U405 (N_405,N_340,N_336);
or U406 (N_406,N_348,N_358);
and U407 (N_407,N_380,N_377);
or U408 (N_408,N_395,N_331);
or U409 (N_409,N_376,N_312);
xor U410 (N_410,N_355,N_369);
nor U411 (N_411,N_346,N_310);
nor U412 (N_412,N_388,N_311);
and U413 (N_413,N_390,N_302);
and U414 (N_414,N_392,N_347);
nand U415 (N_415,N_337,N_371);
nor U416 (N_416,N_363,N_353);
or U417 (N_417,N_366,N_313);
xor U418 (N_418,N_367,N_322);
and U419 (N_419,N_332,N_341);
or U420 (N_420,N_308,N_386);
xnor U421 (N_421,N_385,N_381);
nand U422 (N_422,N_368,N_382);
nor U423 (N_423,N_365,N_345);
nand U424 (N_424,N_306,N_378);
or U425 (N_425,N_325,N_301);
or U426 (N_426,N_370,N_329);
or U427 (N_427,N_351,N_328);
and U428 (N_428,N_374,N_327);
or U429 (N_429,N_389,N_330);
nand U430 (N_430,N_373,N_343);
and U431 (N_431,N_335,N_324);
nor U432 (N_432,N_314,N_344);
nor U433 (N_433,N_321,N_305);
or U434 (N_434,N_304,N_372);
nor U435 (N_435,N_354,N_360);
and U436 (N_436,N_375,N_399);
or U437 (N_437,N_352,N_339);
or U438 (N_438,N_317,N_387);
nor U439 (N_439,N_333,N_338);
or U440 (N_440,N_384,N_303);
and U441 (N_441,N_361,N_356);
and U442 (N_442,N_349,N_316);
nand U443 (N_443,N_307,N_391);
and U444 (N_444,N_326,N_319);
or U445 (N_445,N_320,N_394);
nor U446 (N_446,N_318,N_300);
and U447 (N_447,N_350,N_393);
nor U448 (N_448,N_379,N_334);
and U449 (N_449,N_362,N_398);
and U450 (N_450,N_323,N_387);
xor U451 (N_451,N_357,N_326);
and U452 (N_452,N_314,N_380);
nor U453 (N_453,N_387,N_326);
nand U454 (N_454,N_364,N_302);
and U455 (N_455,N_378,N_399);
or U456 (N_456,N_376,N_392);
nand U457 (N_457,N_300,N_323);
or U458 (N_458,N_391,N_367);
nand U459 (N_459,N_361,N_390);
or U460 (N_460,N_370,N_323);
and U461 (N_461,N_304,N_368);
nor U462 (N_462,N_355,N_324);
and U463 (N_463,N_346,N_398);
or U464 (N_464,N_367,N_389);
nor U465 (N_465,N_372,N_302);
nand U466 (N_466,N_373,N_324);
or U467 (N_467,N_350,N_396);
nand U468 (N_468,N_358,N_328);
or U469 (N_469,N_392,N_390);
nor U470 (N_470,N_313,N_378);
nand U471 (N_471,N_343,N_338);
and U472 (N_472,N_377,N_376);
or U473 (N_473,N_307,N_362);
nor U474 (N_474,N_353,N_306);
and U475 (N_475,N_314,N_373);
and U476 (N_476,N_337,N_312);
nor U477 (N_477,N_306,N_314);
nand U478 (N_478,N_395,N_370);
and U479 (N_479,N_389,N_376);
nand U480 (N_480,N_310,N_305);
and U481 (N_481,N_339,N_312);
nand U482 (N_482,N_302,N_338);
and U483 (N_483,N_383,N_374);
nor U484 (N_484,N_389,N_399);
or U485 (N_485,N_383,N_362);
and U486 (N_486,N_312,N_364);
nor U487 (N_487,N_327,N_378);
nand U488 (N_488,N_334,N_372);
nand U489 (N_489,N_322,N_338);
or U490 (N_490,N_341,N_335);
nand U491 (N_491,N_393,N_342);
and U492 (N_492,N_363,N_355);
and U493 (N_493,N_324,N_345);
and U494 (N_494,N_363,N_321);
and U495 (N_495,N_396,N_348);
nand U496 (N_496,N_370,N_378);
or U497 (N_497,N_307,N_378);
nand U498 (N_498,N_330,N_354);
and U499 (N_499,N_352,N_317);
nor U500 (N_500,N_450,N_424);
nand U501 (N_501,N_423,N_491);
or U502 (N_502,N_411,N_416);
or U503 (N_503,N_428,N_425);
or U504 (N_504,N_488,N_405);
nor U505 (N_505,N_454,N_436);
nor U506 (N_506,N_483,N_460);
or U507 (N_507,N_431,N_400);
nor U508 (N_508,N_496,N_472);
nand U509 (N_509,N_435,N_489);
and U510 (N_510,N_434,N_438);
and U511 (N_511,N_462,N_415);
nor U512 (N_512,N_456,N_401);
nor U513 (N_513,N_480,N_470);
or U514 (N_514,N_441,N_406);
nand U515 (N_515,N_481,N_430);
or U516 (N_516,N_467,N_455);
or U517 (N_517,N_459,N_479);
nor U518 (N_518,N_490,N_494);
and U519 (N_519,N_407,N_477);
nand U520 (N_520,N_484,N_476);
or U521 (N_521,N_427,N_451);
nor U522 (N_522,N_432,N_437);
and U523 (N_523,N_469,N_442);
nand U524 (N_524,N_465,N_497);
or U525 (N_525,N_486,N_449);
nor U526 (N_526,N_446,N_417);
nand U527 (N_527,N_403,N_499);
and U528 (N_528,N_412,N_471);
nand U529 (N_529,N_458,N_429);
nand U530 (N_530,N_478,N_468);
nand U531 (N_531,N_422,N_485);
nor U532 (N_532,N_487,N_495);
or U533 (N_533,N_443,N_448);
or U534 (N_534,N_447,N_492);
nand U535 (N_535,N_482,N_404);
nand U536 (N_536,N_419,N_418);
nand U537 (N_537,N_452,N_402);
and U538 (N_538,N_420,N_426);
nand U539 (N_539,N_457,N_440);
nand U540 (N_540,N_444,N_498);
or U541 (N_541,N_433,N_421);
and U542 (N_542,N_408,N_466);
nand U543 (N_543,N_475,N_463);
nand U544 (N_544,N_473,N_493);
nand U545 (N_545,N_445,N_410);
nand U546 (N_546,N_439,N_461);
and U547 (N_547,N_414,N_413);
nand U548 (N_548,N_409,N_464);
nand U549 (N_549,N_453,N_474);
nor U550 (N_550,N_447,N_434);
or U551 (N_551,N_493,N_483);
nand U552 (N_552,N_491,N_490);
and U553 (N_553,N_416,N_471);
nor U554 (N_554,N_477,N_488);
nand U555 (N_555,N_426,N_435);
or U556 (N_556,N_445,N_451);
nand U557 (N_557,N_404,N_445);
or U558 (N_558,N_476,N_408);
nand U559 (N_559,N_437,N_421);
nand U560 (N_560,N_463,N_441);
or U561 (N_561,N_443,N_430);
or U562 (N_562,N_449,N_415);
nand U563 (N_563,N_472,N_482);
and U564 (N_564,N_461,N_492);
or U565 (N_565,N_421,N_455);
xor U566 (N_566,N_411,N_417);
and U567 (N_567,N_404,N_437);
or U568 (N_568,N_442,N_423);
nand U569 (N_569,N_405,N_485);
or U570 (N_570,N_408,N_419);
or U571 (N_571,N_411,N_492);
and U572 (N_572,N_443,N_422);
or U573 (N_573,N_418,N_411);
nor U574 (N_574,N_478,N_494);
and U575 (N_575,N_434,N_430);
and U576 (N_576,N_465,N_454);
and U577 (N_577,N_481,N_471);
nor U578 (N_578,N_479,N_494);
or U579 (N_579,N_465,N_419);
nand U580 (N_580,N_474,N_429);
or U581 (N_581,N_475,N_415);
nand U582 (N_582,N_458,N_478);
nand U583 (N_583,N_434,N_494);
and U584 (N_584,N_402,N_442);
and U585 (N_585,N_462,N_424);
nor U586 (N_586,N_484,N_494);
or U587 (N_587,N_436,N_464);
and U588 (N_588,N_489,N_428);
and U589 (N_589,N_428,N_465);
nor U590 (N_590,N_489,N_422);
and U591 (N_591,N_463,N_412);
and U592 (N_592,N_405,N_412);
nand U593 (N_593,N_410,N_416);
and U594 (N_594,N_474,N_424);
or U595 (N_595,N_459,N_403);
nand U596 (N_596,N_483,N_418);
nor U597 (N_597,N_410,N_489);
nand U598 (N_598,N_434,N_480);
or U599 (N_599,N_426,N_462);
nand U600 (N_600,N_570,N_533);
nand U601 (N_601,N_501,N_587);
nor U602 (N_602,N_577,N_562);
or U603 (N_603,N_509,N_575);
nor U604 (N_604,N_545,N_552);
nor U605 (N_605,N_596,N_588);
or U606 (N_606,N_544,N_529);
nand U607 (N_607,N_554,N_583);
nor U608 (N_608,N_565,N_578);
and U609 (N_609,N_543,N_566);
or U610 (N_610,N_598,N_556);
nand U611 (N_611,N_503,N_538);
xnor U612 (N_612,N_597,N_548);
nor U613 (N_613,N_582,N_551);
nor U614 (N_614,N_521,N_532);
nand U615 (N_615,N_520,N_557);
or U616 (N_616,N_572,N_531);
nand U617 (N_617,N_567,N_518);
nor U618 (N_618,N_594,N_506);
nor U619 (N_619,N_541,N_510);
or U620 (N_620,N_549,N_500);
nor U621 (N_621,N_580,N_561);
nand U622 (N_622,N_559,N_508);
or U623 (N_623,N_536,N_542);
nor U624 (N_624,N_564,N_517);
nor U625 (N_625,N_526,N_513);
nand U626 (N_626,N_515,N_547);
nand U627 (N_627,N_574,N_571);
xnor U628 (N_628,N_502,N_591);
or U629 (N_629,N_546,N_539);
and U630 (N_630,N_585,N_523);
nor U631 (N_631,N_519,N_568);
nand U632 (N_632,N_555,N_550);
nor U633 (N_633,N_516,N_595);
nor U634 (N_634,N_535,N_573);
xnor U635 (N_635,N_563,N_593);
nand U636 (N_636,N_522,N_569);
nand U637 (N_637,N_590,N_537);
or U638 (N_638,N_560,N_511);
nor U639 (N_639,N_524,N_527);
and U640 (N_640,N_525,N_528);
xor U641 (N_641,N_540,N_553);
nand U642 (N_642,N_534,N_576);
nand U643 (N_643,N_592,N_579);
or U644 (N_644,N_505,N_584);
nor U645 (N_645,N_586,N_530);
nand U646 (N_646,N_507,N_558);
or U647 (N_647,N_581,N_504);
nor U648 (N_648,N_599,N_514);
or U649 (N_649,N_589,N_512);
or U650 (N_650,N_502,N_527);
nand U651 (N_651,N_595,N_575);
and U652 (N_652,N_530,N_584);
nand U653 (N_653,N_564,N_526);
or U654 (N_654,N_501,N_531);
nor U655 (N_655,N_595,N_555);
nand U656 (N_656,N_509,N_561);
or U657 (N_657,N_582,N_505);
xnor U658 (N_658,N_579,N_549);
or U659 (N_659,N_590,N_522);
and U660 (N_660,N_587,N_513);
or U661 (N_661,N_589,N_510);
and U662 (N_662,N_571,N_594);
and U663 (N_663,N_591,N_501);
nor U664 (N_664,N_595,N_530);
nor U665 (N_665,N_566,N_537);
and U666 (N_666,N_545,N_523);
or U667 (N_667,N_556,N_508);
nand U668 (N_668,N_584,N_521);
and U669 (N_669,N_556,N_554);
or U670 (N_670,N_582,N_512);
and U671 (N_671,N_515,N_535);
nor U672 (N_672,N_560,N_581);
and U673 (N_673,N_534,N_556);
and U674 (N_674,N_549,N_532);
nor U675 (N_675,N_526,N_530);
nor U676 (N_676,N_556,N_512);
and U677 (N_677,N_591,N_576);
nand U678 (N_678,N_568,N_543);
or U679 (N_679,N_554,N_567);
nand U680 (N_680,N_533,N_546);
nand U681 (N_681,N_523,N_599);
nor U682 (N_682,N_543,N_597);
or U683 (N_683,N_500,N_508);
and U684 (N_684,N_564,N_506);
and U685 (N_685,N_538,N_548);
and U686 (N_686,N_549,N_570);
or U687 (N_687,N_522,N_528);
xor U688 (N_688,N_531,N_510);
nor U689 (N_689,N_507,N_518);
xnor U690 (N_690,N_505,N_589);
and U691 (N_691,N_578,N_511);
or U692 (N_692,N_515,N_500);
and U693 (N_693,N_575,N_505);
nand U694 (N_694,N_563,N_566);
nand U695 (N_695,N_567,N_571);
and U696 (N_696,N_539,N_564);
and U697 (N_697,N_511,N_592);
nand U698 (N_698,N_531,N_549);
or U699 (N_699,N_512,N_546);
nor U700 (N_700,N_662,N_663);
and U701 (N_701,N_646,N_643);
nand U702 (N_702,N_647,N_629);
nand U703 (N_703,N_678,N_622);
and U704 (N_704,N_645,N_656);
and U705 (N_705,N_610,N_666);
or U706 (N_706,N_636,N_672);
and U707 (N_707,N_657,N_689);
xor U708 (N_708,N_691,N_620);
nand U709 (N_709,N_669,N_698);
or U710 (N_710,N_640,N_632);
or U711 (N_711,N_650,N_612);
nor U712 (N_712,N_677,N_668);
and U713 (N_713,N_693,N_606);
or U714 (N_714,N_664,N_685);
or U715 (N_715,N_680,N_611);
or U716 (N_716,N_655,N_637);
nand U717 (N_717,N_671,N_649);
or U718 (N_718,N_688,N_675);
nor U719 (N_719,N_699,N_631);
nor U720 (N_720,N_648,N_686);
and U721 (N_721,N_604,N_696);
nand U722 (N_722,N_603,N_639);
and U723 (N_723,N_635,N_642);
nor U724 (N_724,N_608,N_695);
or U725 (N_725,N_683,N_697);
nor U726 (N_726,N_651,N_682);
or U727 (N_727,N_630,N_684);
or U728 (N_728,N_623,N_667);
and U729 (N_729,N_607,N_660);
nand U730 (N_730,N_652,N_690);
or U731 (N_731,N_627,N_619);
nand U732 (N_732,N_694,N_615);
nor U733 (N_733,N_628,N_616);
nand U734 (N_734,N_654,N_638);
and U735 (N_735,N_670,N_614);
nand U736 (N_736,N_601,N_665);
and U737 (N_737,N_618,N_600);
or U738 (N_738,N_626,N_602);
nand U739 (N_739,N_609,N_613);
and U740 (N_740,N_658,N_624);
or U741 (N_741,N_625,N_679);
or U742 (N_742,N_617,N_687);
or U743 (N_743,N_692,N_676);
or U744 (N_744,N_674,N_633);
and U745 (N_745,N_653,N_673);
nand U746 (N_746,N_605,N_621);
and U747 (N_747,N_659,N_641);
nand U748 (N_748,N_681,N_644);
or U749 (N_749,N_661,N_634);
nand U750 (N_750,N_600,N_602);
or U751 (N_751,N_692,N_694);
nand U752 (N_752,N_613,N_684);
and U753 (N_753,N_659,N_688);
and U754 (N_754,N_603,N_655);
nor U755 (N_755,N_625,N_692);
nand U756 (N_756,N_670,N_625);
and U757 (N_757,N_680,N_633);
and U758 (N_758,N_655,N_629);
nand U759 (N_759,N_624,N_648);
nor U760 (N_760,N_662,N_649);
nor U761 (N_761,N_636,N_696);
nor U762 (N_762,N_677,N_686);
or U763 (N_763,N_655,N_650);
or U764 (N_764,N_666,N_658);
and U765 (N_765,N_642,N_663);
nor U766 (N_766,N_605,N_679);
and U767 (N_767,N_627,N_667);
nand U768 (N_768,N_635,N_684);
nand U769 (N_769,N_600,N_650);
nand U770 (N_770,N_653,N_606);
or U771 (N_771,N_620,N_608);
nand U772 (N_772,N_676,N_610);
and U773 (N_773,N_604,N_644);
nor U774 (N_774,N_692,N_643);
and U775 (N_775,N_698,N_612);
and U776 (N_776,N_624,N_696);
nor U777 (N_777,N_659,N_699);
and U778 (N_778,N_637,N_668);
xnor U779 (N_779,N_692,N_695);
nand U780 (N_780,N_691,N_626);
nor U781 (N_781,N_651,N_601);
and U782 (N_782,N_679,N_613);
nand U783 (N_783,N_628,N_617);
xnor U784 (N_784,N_695,N_610);
xor U785 (N_785,N_699,N_615);
nor U786 (N_786,N_695,N_699);
and U787 (N_787,N_672,N_699);
nor U788 (N_788,N_605,N_689);
and U789 (N_789,N_651,N_676);
or U790 (N_790,N_691,N_619);
and U791 (N_791,N_624,N_667);
nand U792 (N_792,N_618,N_672);
or U793 (N_793,N_691,N_648);
and U794 (N_794,N_673,N_610);
nor U795 (N_795,N_683,N_694);
nand U796 (N_796,N_643,N_663);
or U797 (N_797,N_673,N_663);
and U798 (N_798,N_606,N_681);
and U799 (N_799,N_639,N_699);
nand U800 (N_800,N_745,N_757);
nand U801 (N_801,N_723,N_797);
and U802 (N_802,N_786,N_711);
and U803 (N_803,N_736,N_734);
or U804 (N_804,N_791,N_766);
and U805 (N_805,N_715,N_775);
or U806 (N_806,N_795,N_751);
and U807 (N_807,N_792,N_724);
nand U808 (N_808,N_740,N_748);
and U809 (N_809,N_778,N_716);
nor U810 (N_810,N_774,N_737);
nor U811 (N_811,N_788,N_755);
or U812 (N_812,N_760,N_764);
and U813 (N_813,N_727,N_752);
or U814 (N_814,N_708,N_758);
nand U815 (N_815,N_728,N_725);
or U816 (N_816,N_798,N_783);
or U817 (N_817,N_731,N_729);
and U818 (N_818,N_741,N_743);
and U819 (N_819,N_789,N_712);
xor U820 (N_820,N_705,N_701);
and U821 (N_821,N_732,N_782);
or U822 (N_822,N_707,N_780);
or U823 (N_823,N_703,N_793);
nor U824 (N_824,N_772,N_738);
and U825 (N_825,N_726,N_767);
nand U826 (N_826,N_776,N_799);
or U827 (N_827,N_753,N_779);
or U828 (N_828,N_749,N_721);
nor U829 (N_829,N_781,N_796);
xnor U830 (N_830,N_761,N_770);
or U831 (N_831,N_717,N_744);
and U832 (N_832,N_784,N_759);
and U833 (N_833,N_790,N_763);
nand U834 (N_834,N_722,N_768);
nand U835 (N_835,N_739,N_769);
and U836 (N_836,N_700,N_746);
nand U837 (N_837,N_765,N_747);
nor U838 (N_838,N_702,N_785);
nor U839 (N_839,N_714,N_710);
or U840 (N_840,N_713,N_706);
nand U841 (N_841,N_773,N_735);
nor U842 (N_842,N_756,N_720);
and U843 (N_843,N_733,N_794);
or U844 (N_844,N_704,N_754);
nor U845 (N_845,N_750,N_771);
nand U846 (N_846,N_787,N_742);
xnor U847 (N_847,N_762,N_709);
or U848 (N_848,N_777,N_719);
nand U849 (N_849,N_730,N_718);
nand U850 (N_850,N_746,N_753);
nor U851 (N_851,N_782,N_703);
and U852 (N_852,N_740,N_790);
and U853 (N_853,N_725,N_714);
or U854 (N_854,N_793,N_752);
or U855 (N_855,N_700,N_747);
and U856 (N_856,N_713,N_732);
nand U857 (N_857,N_771,N_764);
or U858 (N_858,N_725,N_799);
nor U859 (N_859,N_773,N_744);
or U860 (N_860,N_771,N_732);
nand U861 (N_861,N_730,N_795);
nand U862 (N_862,N_770,N_757);
or U863 (N_863,N_798,N_779);
nand U864 (N_864,N_735,N_775);
or U865 (N_865,N_737,N_778);
nand U866 (N_866,N_750,N_720);
nor U867 (N_867,N_709,N_766);
or U868 (N_868,N_705,N_794);
or U869 (N_869,N_750,N_751);
or U870 (N_870,N_755,N_762);
and U871 (N_871,N_783,N_765);
nor U872 (N_872,N_787,N_766);
or U873 (N_873,N_766,N_755);
nand U874 (N_874,N_773,N_706);
or U875 (N_875,N_795,N_763);
nor U876 (N_876,N_703,N_710);
nor U877 (N_877,N_788,N_724);
nand U878 (N_878,N_783,N_712);
nor U879 (N_879,N_721,N_775);
and U880 (N_880,N_759,N_716);
nand U881 (N_881,N_749,N_709);
or U882 (N_882,N_797,N_701);
or U883 (N_883,N_714,N_771);
nor U884 (N_884,N_752,N_765);
nand U885 (N_885,N_734,N_743);
nand U886 (N_886,N_750,N_704);
nor U887 (N_887,N_724,N_760);
nor U888 (N_888,N_715,N_756);
nand U889 (N_889,N_792,N_738);
or U890 (N_890,N_791,N_799);
and U891 (N_891,N_787,N_734);
or U892 (N_892,N_730,N_728);
nor U893 (N_893,N_710,N_732);
nor U894 (N_894,N_784,N_746);
and U895 (N_895,N_785,N_752);
or U896 (N_896,N_776,N_787);
nand U897 (N_897,N_753,N_721);
nor U898 (N_898,N_753,N_751);
and U899 (N_899,N_765,N_758);
nor U900 (N_900,N_881,N_887);
nand U901 (N_901,N_832,N_891);
nor U902 (N_902,N_849,N_861);
nor U903 (N_903,N_896,N_868);
and U904 (N_904,N_855,N_836);
and U905 (N_905,N_844,N_841);
or U906 (N_906,N_898,N_831);
nor U907 (N_907,N_857,N_879);
and U908 (N_908,N_885,N_888);
or U909 (N_909,N_893,N_899);
nand U910 (N_910,N_852,N_864);
and U911 (N_911,N_801,N_895);
or U912 (N_912,N_810,N_871);
nor U913 (N_913,N_823,N_850);
or U914 (N_914,N_867,N_804);
nand U915 (N_915,N_872,N_851);
nor U916 (N_916,N_884,N_890);
nand U917 (N_917,N_856,N_889);
and U918 (N_918,N_821,N_878);
nand U919 (N_919,N_815,N_814);
nand U920 (N_920,N_827,N_894);
nor U921 (N_921,N_842,N_825);
or U922 (N_922,N_876,N_848);
nand U923 (N_923,N_812,N_807);
or U924 (N_924,N_805,N_818);
and U925 (N_925,N_811,N_880);
nand U926 (N_926,N_837,N_886);
or U927 (N_927,N_829,N_826);
nor U928 (N_928,N_854,N_869);
and U929 (N_929,N_846,N_892);
and U930 (N_930,N_875,N_897);
nand U931 (N_931,N_813,N_853);
nand U932 (N_932,N_882,N_830);
nand U933 (N_933,N_809,N_803);
nand U934 (N_934,N_883,N_828);
or U935 (N_935,N_860,N_824);
and U936 (N_936,N_820,N_819);
nor U937 (N_937,N_870,N_859);
nand U938 (N_938,N_822,N_806);
or U939 (N_939,N_843,N_808);
and U940 (N_940,N_816,N_873);
nand U941 (N_941,N_863,N_845);
or U942 (N_942,N_835,N_847);
xnor U943 (N_943,N_840,N_800);
and U944 (N_944,N_838,N_877);
nand U945 (N_945,N_833,N_862);
or U946 (N_946,N_866,N_839);
nand U947 (N_947,N_858,N_834);
and U948 (N_948,N_817,N_865);
nor U949 (N_949,N_802,N_874);
nor U950 (N_950,N_812,N_868);
nor U951 (N_951,N_832,N_863);
and U952 (N_952,N_881,N_848);
or U953 (N_953,N_880,N_822);
and U954 (N_954,N_840,N_891);
and U955 (N_955,N_893,N_855);
xor U956 (N_956,N_805,N_859);
nor U957 (N_957,N_878,N_806);
or U958 (N_958,N_864,N_854);
nand U959 (N_959,N_831,N_856);
nand U960 (N_960,N_840,N_834);
and U961 (N_961,N_873,N_831);
nor U962 (N_962,N_871,N_846);
and U963 (N_963,N_893,N_867);
nand U964 (N_964,N_810,N_823);
and U965 (N_965,N_811,N_896);
or U966 (N_966,N_803,N_827);
nor U967 (N_967,N_890,N_858);
nand U968 (N_968,N_849,N_875);
and U969 (N_969,N_853,N_801);
nand U970 (N_970,N_819,N_852);
nor U971 (N_971,N_841,N_804);
nor U972 (N_972,N_857,N_886);
and U973 (N_973,N_876,N_879);
or U974 (N_974,N_868,N_846);
or U975 (N_975,N_888,N_844);
and U976 (N_976,N_883,N_866);
and U977 (N_977,N_812,N_817);
nand U978 (N_978,N_899,N_878);
nor U979 (N_979,N_899,N_816);
nand U980 (N_980,N_851,N_827);
or U981 (N_981,N_824,N_896);
or U982 (N_982,N_822,N_869);
nor U983 (N_983,N_808,N_874);
nand U984 (N_984,N_877,N_881);
and U985 (N_985,N_896,N_801);
or U986 (N_986,N_881,N_895);
and U987 (N_987,N_828,N_857);
nand U988 (N_988,N_807,N_820);
or U989 (N_989,N_829,N_837);
and U990 (N_990,N_824,N_875);
nor U991 (N_991,N_828,N_814);
and U992 (N_992,N_892,N_800);
and U993 (N_993,N_832,N_833);
nor U994 (N_994,N_877,N_876);
and U995 (N_995,N_853,N_882);
nor U996 (N_996,N_833,N_831);
nand U997 (N_997,N_815,N_862);
nor U998 (N_998,N_833,N_866);
and U999 (N_999,N_883,N_893);
nand U1000 (N_1000,N_920,N_916);
and U1001 (N_1001,N_981,N_934);
and U1002 (N_1002,N_931,N_912);
xnor U1003 (N_1003,N_974,N_952);
and U1004 (N_1004,N_954,N_918);
or U1005 (N_1005,N_970,N_953);
nor U1006 (N_1006,N_988,N_989);
nor U1007 (N_1007,N_992,N_951);
or U1008 (N_1008,N_994,N_959);
and U1009 (N_1009,N_969,N_977);
and U1010 (N_1010,N_911,N_941);
nor U1011 (N_1011,N_938,N_986);
xor U1012 (N_1012,N_967,N_921);
and U1013 (N_1013,N_945,N_955);
and U1014 (N_1014,N_930,N_915);
nor U1015 (N_1015,N_927,N_904);
and U1016 (N_1016,N_906,N_987);
or U1017 (N_1017,N_908,N_972);
nor U1018 (N_1018,N_932,N_925);
nand U1019 (N_1019,N_996,N_935);
or U1020 (N_1020,N_900,N_946);
nand U1021 (N_1021,N_923,N_907);
nand U1022 (N_1022,N_929,N_905);
and U1023 (N_1023,N_922,N_928);
and U1024 (N_1024,N_985,N_983);
and U1025 (N_1025,N_936,N_999);
or U1026 (N_1026,N_933,N_975);
nor U1027 (N_1027,N_937,N_990);
or U1028 (N_1028,N_901,N_980);
or U1029 (N_1029,N_960,N_982);
nand U1030 (N_1030,N_961,N_947);
or U1031 (N_1031,N_965,N_942);
nor U1032 (N_1032,N_909,N_979);
nor U1033 (N_1033,N_910,N_971);
nand U1034 (N_1034,N_949,N_997);
nand U1035 (N_1035,N_948,N_919);
nand U1036 (N_1036,N_940,N_926);
nand U1037 (N_1037,N_958,N_917);
nor U1038 (N_1038,N_993,N_943);
nor U1039 (N_1039,N_939,N_956);
nor U1040 (N_1040,N_963,N_966);
or U1041 (N_1041,N_998,N_962);
nor U1042 (N_1042,N_903,N_902);
nand U1043 (N_1043,N_976,N_914);
nor U1044 (N_1044,N_944,N_913);
nand U1045 (N_1045,N_957,N_984);
nand U1046 (N_1046,N_950,N_991);
and U1047 (N_1047,N_924,N_964);
nor U1048 (N_1048,N_973,N_978);
and U1049 (N_1049,N_968,N_995);
nand U1050 (N_1050,N_903,N_977);
xor U1051 (N_1051,N_938,N_908);
nor U1052 (N_1052,N_985,N_938);
nor U1053 (N_1053,N_997,N_948);
and U1054 (N_1054,N_999,N_933);
nand U1055 (N_1055,N_908,N_980);
xnor U1056 (N_1056,N_973,N_951);
or U1057 (N_1057,N_987,N_972);
or U1058 (N_1058,N_941,N_963);
nand U1059 (N_1059,N_928,N_900);
and U1060 (N_1060,N_986,N_932);
nand U1061 (N_1061,N_991,N_961);
and U1062 (N_1062,N_995,N_959);
nand U1063 (N_1063,N_916,N_976);
nand U1064 (N_1064,N_986,N_971);
or U1065 (N_1065,N_972,N_933);
nand U1066 (N_1066,N_931,N_946);
and U1067 (N_1067,N_976,N_989);
or U1068 (N_1068,N_911,N_976);
nand U1069 (N_1069,N_998,N_900);
nand U1070 (N_1070,N_913,N_954);
and U1071 (N_1071,N_961,N_965);
nor U1072 (N_1072,N_948,N_965);
and U1073 (N_1073,N_941,N_986);
and U1074 (N_1074,N_961,N_912);
or U1075 (N_1075,N_929,N_954);
nor U1076 (N_1076,N_956,N_920);
xnor U1077 (N_1077,N_904,N_951);
or U1078 (N_1078,N_936,N_955);
or U1079 (N_1079,N_961,N_983);
or U1080 (N_1080,N_907,N_927);
nand U1081 (N_1081,N_912,N_996);
nor U1082 (N_1082,N_904,N_934);
or U1083 (N_1083,N_924,N_925);
and U1084 (N_1084,N_967,N_906);
nor U1085 (N_1085,N_950,N_921);
or U1086 (N_1086,N_954,N_999);
or U1087 (N_1087,N_904,N_915);
and U1088 (N_1088,N_946,N_971);
xor U1089 (N_1089,N_906,N_932);
or U1090 (N_1090,N_966,N_967);
xnor U1091 (N_1091,N_934,N_915);
nor U1092 (N_1092,N_902,N_963);
and U1093 (N_1093,N_956,N_935);
or U1094 (N_1094,N_984,N_959);
or U1095 (N_1095,N_939,N_910);
and U1096 (N_1096,N_902,N_913);
nand U1097 (N_1097,N_916,N_949);
or U1098 (N_1098,N_933,N_960);
nor U1099 (N_1099,N_966,N_965);
or U1100 (N_1100,N_1099,N_1037);
nor U1101 (N_1101,N_1017,N_1089);
nand U1102 (N_1102,N_1049,N_1027);
and U1103 (N_1103,N_1033,N_1043);
or U1104 (N_1104,N_1021,N_1077);
or U1105 (N_1105,N_1046,N_1059);
or U1106 (N_1106,N_1002,N_1098);
or U1107 (N_1107,N_1000,N_1079);
nand U1108 (N_1108,N_1020,N_1072);
nand U1109 (N_1109,N_1092,N_1032);
nor U1110 (N_1110,N_1090,N_1042);
and U1111 (N_1111,N_1055,N_1086);
nand U1112 (N_1112,N_1082,N_1084);
nand U1113 (N_1113,N_1029,N_1095);
or U1114 (N_1114,N_1019,N_1070);
nor U1115 (N_1115,N_1035,N_1023);
nor U1116 (N_1116,N_1096,N_1094);
nand U1117 (N_1117,N_1015,N_1064);
or U1118 (N_1118,N_1008,N_1091);
nand U1119 (N_1119,N_1013,N_1093);
or U1120 (N_1120,N_1041,N_1050);
and U1121 (N_1121,N_1034,N_1087);
nor U1122 (N_1122,N_1052,N_1018);
nor U1123 (N_1123,N_1040,N_1026);
or U1124 (N_1124,N_1001,N_1039);
nor U1125 (N_1125,N_1057,N_1047);
nand U1126 (N_1126,N_1031,N_1045);
nand U1127 (N_1127,N_1075,N_1028);
nor U1128 (N_1128,N_1066,N_1030);
and U1129 (N_1129,N_1056,N_1053);
and U1130 (N_1130,N_1016,N_1068);
and U1131 (N_1131,N_1038,N_1080);
nor U1132 (N_1132,N_1025,N_1048);
nor U1133 (N_1133,N_1010,N_1071);
nor U1134 (N_1134,N_1062,N_1069);
nor U1135 (N_1135,N_1076,N_1063);
nor U1136 (N_1136,N_1003,N_1004);
nor U1137 (N_1137,N_1022,N_1054);
and U1138 (N_1138,N_1060,N_1011);
or U1139 (N_1139,N_1007,N_1083);
nor U1140 (N_1140,N_1051,N_1088);
and U1141 (N_1141,N_1065,N_1012);
and U1142 (N_1142,N_1061,N_1097);
nand U1143 (N_1143,N_1005,N_1081);
nand U1144 (N_1144,N_1036,N_1014);
and U1145 (N_1145,N_1009,N_1058);
nand U1146 (N_1146,N_1073,N_1067);
or U1147 (N_1147,N_1044,N_1006);
nand U1148 (N_1148,N_1085,N_1074);
xnor U1149 (N_1149,N_1024,N_1078);
nor U1150 (N_1150,N_1094,N_1088);
and U1151 (N_1151,N_1041,N_1026);
and U1152 (N_1152,N_1000,N_1068);
and U1153 (N_1153,N_1006,N_1007);
nor U1154 (N_1154,N_1061,N_1031);
or U1155 (N_1155,N_1067,N_1063);
nand U1156 (N_1156,N_1050,N_1049);
nor U1157 (N_1157,N_1059,N_1007);
nor U1158 (N_1158,N_1077,N_1049);
and U1159 (N_1159,N_1040,N_1082);
or U1160 (N_1160,N_1059,N_1038);
and U1161 (N_1161,N_1071,N_1062);
nand U1162 (N_1162,N_1023,N_1098);
or U1163 (N_1163,N_1025,N_1078);
and U1164 (N_1164,N_1043,N_1070);
and U1165 (N_1165,N_1092,N_1096);
or U1166 (N_1166,N_1001,N_1044);
or U1167 (N_1167,N_1090,N_1012);
or U1168 (N_1168,N_1069,N_1097);
or U1169 (N_1169,N_1003,N_1028);
nor U1170 (N_1170,N_1030,N_1076);
and U1171 (N_1171,N_1002,N_1054);
nand U1172 (N_1172,N_1031,N_1035);
or U1173 (N_1173,N_1012,N_1083);
or U1174 (N_1174,N_1060,N_1046);
nor U1175 (N_1175,N_1060,N_1056);
nand U1176 (N_1176,N_1092,N_1017);
nor U1177 (N_1177,N_1009,N_1068);
and U1178 (N_1178,N_1037,N_1031);
and U1179 (N_1179,N_1035,N_1071);
or U1180 (N_1180,N_1087,N_1036);
nor U1181 (N_1181,N_1011,N_1021);
and U1182 (N_1182,N_1015,N_1034);
nand U1183 (N_1183,N_1088,N_1007);
nor U1184 (N_1184,N_1081,N_1067);
and U1185 (N_1185,N_1002,N_1090);
or U1186 (N_1186,N_1053,N_1046);
nor U1187 (N_1187,N_1094,N_1040);
and U1188 (N_1188,N_1059,N_1095);
and U1189 (N_1189,N_1054,N_1044);
and U1190 (N_1190,N_1006,N_1089);
or U1191 (N_1191,N_1072,N_1085);
nor U1192 (N_1192,N_1071,N_1042);
nor U1193 (N_1193,N_1050,N_1086);
and U1194 (N_1194,N_1005,N_1045);
or U1195 (N_1195,N_1000,N_1056);
nand U1196 (N_1196,N_1018,N_1036);
nor U1197 (N_1197,N_1048,N_1061);
or U1198 (N_1198,N_1054,N_1008);
nand U1199 (N_1199,N_1005,N_1041);
nand U1200 (N_1200,N_1155,N_1136);
nor U1201 (N_1201,N_1154,N_1147);
nor U1202 (N_1202,N_1184,N_1174);
nor U1203 (N_1203,N_1187,N_1111);
nor U1204 (N_1204,N_1180,N_1140);
nor U1205 (N_1205,N_1151,N_1146);
nand U1206 (N_1206,N_1192,N_1145);
nor U1207 (N_1207,N_1179,N_1109);
nand U1208 (N_1208,N_1130,N_1128);
nand U1209 (N_1209,N_1189,N_1162);
and U1210 (N_1210,N_1120,N_1115);
nand U1211 (N_1211,N_1113,N_1144);
or U1212 (N_1212,N_1188,N_1177);
and U1213 (N_1213,N_1152,N_1186);
or U1214 (N_1214,N_1102,N_1131);
or U1215 (N_1215,N_1166,N_1100);
nor U1216 (N_1216,N_1183,N_1138);
nand U1217 (N_1217,N_1172,N_1178);
and U1218 (N_1218,N_1104,N_1157);
and U1219 (N_1219,N_1193,N_1123);
and U1220 (N_1220,N_1122,N_1121);
or U1221 (N_1221,N_1126,N_1134);
nor U1222 (N_1222,N_1160,N_1112);
and U1223 (N_1223,N_1103,N_1196);
or U1224 (N_1224,N_1118,N_1137);
xnor U1225 (N_1225,N_1168,N_1114);
nand U1226 (N_1226,N_1141,N_1161);
nor U1227 (N_1227,N_1171,N_1199);
or U1228 (N_1228,N_1164,N_1108);
xor U1229 (N_1229,N_1117,N_1150);
and U1230 (N_1230,N_1105,N_1132);
or U1231 (N_1231,N_1181,N_1142);
nand U1232 (N_1232,N_1127,N_1173);
or U1233 (N_1233,N_1110,N_1198);
or U1234 (N_1234,N_1156,N_1148);
xor U1235 (N_1235,N_1116,N_1163);
nor U1236 (N_1236,N_1139,N_1149);
or U1237 (N_1237,N_1125,N_1133);
nand U1238 (N_1238,N_1124,N_1170);
and U1239 (N_1239,N_1159,N_1107);
or U1240 (N_1240,N_1106,N_1129);
nor U1241 (N_1241,N_1194,N_1176);
nor U1242 (N_1242,N_1169,N_1190);
nor U1243 (N_1243,N_1165,N_1158);
nor U1244 (N_1244,N_1185,N_1143);
nor U1245 (N_1245,N_1191,N_1197);
or U1246 (N_1246,N_1175,N_1153);
or U1247 (N_1247,N_1182,N_1101);
nor U1248 (N_1248,N_1135,N_1195);
nor U1249 (N_1249,N_1119,N_1167);
nand U1250 (N_1250,N_1186,N_1191);
or U1251 (N_1251,N_1120,N_1170);
and U1252 (N_1252,N_1122,N_1141);
nor U1253 (N_1253,N_1137,N_1199);
nand U1254 (N_1254,N_1193,N_1181);
and U1255 (N_1255,N_1146,N_1180);
and U1256 (N_1256,N_1142,N_1156);
and U1257 (N_1257,N_1104,N_1179);
nor U1258 (N_1258,N_1154,N_1185);
nor U1259 (N_1259,N_1174,N_1141);
nor U1260 (N_1260,N_1104,N_1154);
or U1261 (N_1261,N_1147,N_1198);
and U1262 (N_1262,N_1124,N_1190);
and U1263 (N_1263,N_1113,N_1142);
nor U1264 (N_1264,N_1145,N_1191);
and U1265 (N_1265,N_1119,N_1190);
nand U1266 (N_1266,N_1151,N_1193);
nor U1267 (N_1267,N_1196,N_1121);
and U1268 (N_1268,N_1137,N_1195);
or U1269 (N_1269,N_1182,N_1158);
nand U1270 (N_1270,N_1183,N_1137);
nor U1271 (N_1271,N_1126,N_1116);
xnor U1272 (N_1272,N_1193,N_1150);
or U1273 (N_1273,N_1148,N_1177);
or U1274 (N_1274,N_1118,N_1131);
nor U1275 (N_1275,N_1146,N_1135);
nand U1276 (N_1276,N_1153,N_1144);
nor U1277 (N_1277,N_1150,N_1147);
nand U1278 (N_1278,N_1183,N_1163);
and U1279 (N_1279,N_1101,N_1119);
and U1280 (N_1280,N_1137,N_1173);
nor U1281 (N_1281,N_1120,N_1141);
nor U1282 (N_1282,N_1120,N_1105);
xnor U1283 (N_1283,N_1157,N_1107);
and U1284 (N_1284,N_1120,N_1180);
and U1285 (N_1285,N_1106,N_1155);
or U1286 (N_1286,N_1152,N_1190);
and U1287 (N_1287,N_1107,N_1127);
and U1288 (N_1288,N_1176,N_1182);
and U1289 (N_1289,N_1124,N_1163);
and U1290 (N_1290,N_1194,N_1117);
or U1291 (N_1291,N_1126,N_1178);
nor U1292 (N_1292,N_1159,N_1154);
nand U1293 (N_1293,N_1197,N_1185);
nor U1294 (N_1294,N_1107,N_1190);
or U1295 (N_1295,N_1146,N_1120);
nor U1296 (N_1296,N_1175,N_1117);
nor U1297 (N_1297,N_1120,N_1188);
xnor U1298 (N_1298,N_1120,N_1123);
or U1299 (N_1299,N_1190,N_1132);
or U1300 (N_1300,N_1200,N_1280);
nor U1301 (N_1301,N_1225,N_1206);
or U1302 (N_1302,N_1230,N_1238);
nor U1303 (N_1303,N_1278,N_1255);
and U1304 (N_1304,N_1263,N_1288);
nand U1305 (N_1305,N_1207,N_1271);
nand U1306 (N_1306,N_1285,N_1213);
nor U1307 (N_1307,N_1268,N_1277);
nand U1308 (N_1308,N_1246,N_1259);
nor U1309 (N_1309,N_1284,N_1218);
nand U1310 (N_1310,N_1294,N_1203);
or U1311 (N_1311,N_1209,N_1286);
or U1312 (N_1312,N_1232,N_1290);
nor U1313 (N_1313,N_1276,N_1235);
and U1314 (N_1314,N_1272,N_1221);
nor U1315 (N_1315,N_1279,N_1264);
and U1316 (N_1316,N_1248,N_1227);
nor U1317 (N_1317,N_1234,N_1295);
nand U1318 (N_1318,N_1243,N_1208);
nor U1319 (N_1319,N_1253,N_1287);
nand U1320 (N_1320,N_1252,N_1273);
and U1321 (N_1321,N_1254,N_1257);
or U1322 (N_1322,N_1293,N_1216);
and U1323 (N_1323,N_1245,N_1215);
or U1324 (N_1324,N_1298,N_1274);
nor U1325 (N_1325,N_1242,N_1291);
or U1326 (N_1326,N_1236,N_1239);
nand U1327 (N_1327,N_1250,N_1237);
xor U1328 (N_1328,N_1219,N_1240);
and U1329 (N_1329,N_1223,N_1260);
and U1330 (N_1330,N_1229,N_1205);
nor U1331 (N_1331,N_1226,N_1210);
nand U1332 (N_1332,N_1292,N_1211);
and U1333 (N_1333,N_1261,N_1217);
nor U1334 (N_1334,N_1201,N_1282);
nand U1335 (N_1335,N_1299,N_1251);
or U1336 (N_1336,N_1233,N_1222);
nor U1337 (N_1337,N_1297,N_1281);
xor U1338 (N_1338,N_1228,N_1296);
and U1339 (N_1339,N_1283,N_1266);
and U1340 (N_1340,N_1241,N_1258);
or U1341 (N_1341,N_1256,N_1224);
or U1342 (N_1342,N_1231,N_1202);
or U1343 (N_1343,N_1270,N_1275);
nor U1344 (N_1344,N_1262,N_1214);
nor U1345 (N_1345,N_1204,N_1244);
or U1346 (N_1346,N_1269,N_1289);
and U1347 (N_1347,N_1212,N_1267);
nand U1348 (N_1348,N_1265,N_1220);
and U1349 (N_1349,N_1247,N_1249);
or U1350 (N_1350,N_1284,N_1266);
nand U1351 (N_1351,N_1248,N_1278);
or U1352 (N_1352,N_1266,N_1274);
and U1353 (N_1353,N_1205,N_1234);
and U1354 (N_1354,N_1225,N_1227);
nor U1355 (N_1355,N_1297,N_1220);
nor U1356 (N_1356,N_1289,N_1263);
and U1357 (N_1357,N_1283,N_1206);
or U1358 (N_1358,N_1212,N_1215);
xnor U1359 (N_1359,N_1295,N_1294);
nand U1360 (N_1360,N_1265,N_1280);
nand U1361 (N_1361,N_1286,N_1258);
nor U1362 (N_1362,N_1231,N_1272);
and U1363 (N_1363,N_1248,N_1282);
and U1364 (N_1364,N_1260,N_1250);
nand U1365 (N_1365,N_1223,N_1296);
nor U1366 (N_1366,N_1269,N_1244);
and U1367 (N_1367,N_1281,N_1274);
and U1368 (N_1368,N_1268,N_1263);
nor U1369 (N_1369,N_1270,N_1262);
nand U1370 (N_1370,N_1295,N_1259);
or U1371 (N_1371,N_1278,N_1237);
and U1372 (N_1372,N_1253,N_1261);
nand U1373 (N_1373,N_1237,N_1248);
or U1374 (N_1374,N_1278,N_1219);
or U1375 (N_1375,N_1238,N_1277);
or U1376 (N_1376,N_1226,N_1214);
nand U1377 (N_1377,N_1257,N_1217);
nor U1378 (N_1378,N_1291,N_1263);
nor U1379 (N_1379,N_1282,N_1210);
or U1380 (N_1380,N_1230,N_1293);
or U1381 (N_1381,N_1283,N_1239);
and U1382 (N_1382,N_1266,N_1240);
nand U1383 (N_1383,N_1213,N_1291);
and U1384 (N_1384,N_1206,N_1203);
nand U1385 (N_1385,N_1201,N_1245);
xor U1386 (N_1386,N_1226,N_1249);
or U1387 (N_1387,N_1247,N_1259);
and U1388 (N_1388,N_1220,N_1242);
and U1389 (N_1389,N_1281,N_1218);
nor U1390 (N_1390,N_1299,N_1202);
nor U1391 (N_1391,N_1204,N_1233);
nor U1392 (N_1392,N_1206,N_1266);
nor U1393 (N_1393,N_1265,N_1216);
and U1394 (N_1394,N_1244,N_1291);
and U1395 (N_1395,N_1284,N_1274);
and U1396 (N_1396,N_1242,N_1230);
nor U1397 (N_1397,N_1212,N_1238);
nor U1398 (N_1398,N_1257,N_1203);
and U1399 (N_1399,N_1265,N_1228);
and U1400 (N_1400,N_1364,N_1394);
and U1401 (N_1401,N_1385,N_1321);
nor U1402 (N_1402,N_1351,N_1341);
nand U1403 (N_1403,N_1309,N_1330);
nand U1404 (N_1404,N_1395,N_1327);
or U1405 (N_1405,N_1342,N_1371);
nand U1406 (N_1406,N_1374,N_1375);
and U1407 (N_1407,N_1310,N_1393);
and U1408 (N_1408,N_1336,N_1312);
nand U1409 (N_1409,N_1356,N_1349);
nand U1410 (N_1410,N_1319,N_1300);
nor U1411 (N_1411,N_1311,N_1302);
and U1412 (N_1412,N_1305,N_1329);
or U1413 (N_1413,N_1359,N_1301);
and U1414 (N_1414,N_1396,N_1387);
nand U1415 (N_1415,N_1365,N_1343);
nand U1416 (N_1416,N_1362,N_1358);
nor U1417 (N_1417,N_1317,N_1368);
or U1418 (N_1418,N_1326,N_1315);
and U1419 (N_1419,N_1308,N_1337);
or U1420 (N_1420,N_1307,N_1383);
and U1421 (N_1421,N_1388,N_1333);
or U1422 (N_1422,N_1370,N_1360);
or U1423 (N_1423,N_1357,N_1340);
nor U1424 (N_1424,N_1314,N_1379);
or U1425 (N_1425,N_1399,N_1372);
nand U1426 (N_1426,N_1334,N_1338);
or U1427 (N_1427,N_1376,N_1304);
and U1428 (N_1428,N_1377,N_1384);
nand U1429 (N_1429,N_1324,N_1318);
xor U1430 (N_1430,N_1344,N_1363);
nor U1431 (N_1431,N_1323,N_1345);
nand U1432 (N_1432,N_1339,N_1354);
nand U1433 (N_1433,N_1378,N_1331);
and U1434 (N_1434,N_1361,N_1347);
and U1435 (N_1435,N_1386,N_1322);
nor U1436 (N_1436,N_1320,N_1381);
and U1437 (N_1437,N_1373,N_1352);
nand U1438 (N_1438,N_1335,N_1390);
nand U1439 (N_1439,N_1353,N_1325);
xor U1440 (N_1440,N_1398,N_1382);
or U1441 (N_1441,N_1350,N_1389);
nor U1442 (N_1442,N_1332,N_1367);
nand U1443 (N_1443,N_1346,N_1306);
and U1444 (N_1444,N_1303,N_1366);
nand U1445 (N_1445,N_1391,N_1369);
or U1446 (N_1446,N_1355,N_1313);
nor U1447 (N_1447,N_1348,N_1316);
xor U1448 (N_1448,N_1392,N_1397);
or U1449 (N_1449,N_1380,N_1328);
and U1450 (N_1450,N_1310,N_1359);
and U1451 (N_1451,N_1363,N_1368);
or U1452 (N_1452,N_1351,N_1311);
nor U1453 (N_1453,N_1393,N_1365);
nor U1454 (N_1454,N_1399,N_1309);
nand U1455 (N_1455,N_1353,N_1340);
xor U1456 (N_1456,N_1363,N_1301);
and U1457 (N_1457,N_1383,N_1319);
and U1458 (N_1458,N_1343,N_1368);
and U1459 (N_1459,N_1366,N_1317);
nor U1460 (N_1460,N_1316,N_1326);
xnor U1461 (N_1461,N_1384,N_1363);
nor U1462 (N_1462,N_1344,N_1316);
and U1463 (N_1463,N_1383,N_1312);
and U1464 (N_1464,N_1349,N_1323);
nand U1465 (N_1465,N_1395,N_1358);
and U1466 (N_1466,N_1338,N_1317);
nor U1467 (N_1467,N_1361,N_1320);
and U1468 (N_1468,N_1316,N_1391);
nand U1469 (N_1469,N_1301,N_1385);
or U1470 (N_1470,N_1348,N_1325);
nand U1471 (N_1471,N_1374,N_1342);
and U1472 (N_1472,N_1317,N_1309);
nor U1473 (N_1473,N_1355,N_1344);
nand U1474 (N_1474,N_1332,N_1390);
or U1475 (N_1475,N_1317,N_1320);
and U1476 (N_1476,N_1322,N_1315);
xnor U1477 (N_1477,N_1353,N_1379);
nand U1478 (N_1478,N_1306,N_1371);
or U1479 (N_1479,N_1365,N_1332);
and U1480 (N_1480,N_1330,N_1306);
and U1481 (N_1481,N_1358,N_1359);
and U1482 (N_1482,N_1330,N_1303);
or U1483 (N_1483,N_1391,N_1393);
xor U1484 (N_1484,N_1301,N_1362);
and U1485 (N_1485,N_1324,N_1310);
and U1486 (N_1486,N_1362,N_1314);
or U1487 (N_1487,N_1321,N_1331);
nand U1488 (N_1488,N_1323,N_1347);
nor U1489 (N_1489,N_1344,N_1331);
and U1490 (N_1490,N_1354,N_1378);
nand U1491 (N_1491,N_1393,N_1345);
xnor U1492 (N_1492,N_1385,N_1343);
or U1493 (N_1493,N_1383,N_1326);
nand U1494 (N_1494,N_1333,N_1319);
and U1495 (N_1495,N_1371,N_1329);
and U1496 (N_1496,N_1360,N_1398);
nand U1497 (N_1497,N_1348,N_1318);
or U1498 (N_1498,N_1310,N_1334);
nand U1499 (N_1499,N_1377,N_1323);
nand U1500 (N_1500,N_1417,N_1437);
or U1501 (N_1501,N_1418,N_1402);
nand U1502 (N_1502,N_1468,N_1461);
nor U1503 (N_1503,N_1441,N_1490);
or U1504 (N_1504,N_1450,N_1413);
nand U1505 (N_1505,N_1470,N_1452);
nor U1506 (N_1506,N_1478,N_1429);
nor U1507 (N_1507,N_1498,N_1479);
nor U1508 (N_1508,N_1444,N_1427);
nand U1509 (N_1509,N_1431,N_1496);
nor U1510 (N_1510,N_1488,N_1474);
and U1511 (N_1511,N_1484,N_1400);
nor U1512 (N_1512,N_1409,N_1458);
and U1513 (N_1513,N_1442,N_1464);
nor U1514 (N_1514,N_1489,N_1414);
xor U1515 (N_1515,N_1411,N_1422);
and U1516 (N_1516,N_1412,N_1473);
and U1517 (N_1517,N_1421,N_1416);
or U1518 (N_1518,N_1471,N_1495);
or U1519 (N_1519,N_1419,N_1405);
nor U1520 (N_1520,N_1447,N_1404);
nand U1521 (N_1521,N_1477,N_1497);
nor U1522 (N_1522,N_1424,N_1481);
or U1523 (N_1523,N_1459,N_1446);
nor U1524 (N_1524,N_1467,N_1439);
or U1525 (N_1525,N_1434,N_1469);
nor U1526 (N_1526,N_1426,N_1423);
nor U1527 (N_1527,N_1487,N_1455);
nor U1528 (N_1528,N_1494,N_1410);
nand U1529 (N_1529,N_1486,N_1425);
and U1530 (N_1530,N_1499,N_1480);
and U1531 (N_1531,N_1440,N_1401);
nand U1532 (N_1532,N_1493,N_1485);
nor U1533 (N_1533,N_1483,N_1449);
and U1534 (N_1534,N_1462,N_1491);
or U1535 (N_1535,N_1448,N_1457);
or U1536 (N_1536,N_1408,N_1407);
nand U1537 (N_1537,N_1472,N_1465);
or U1538 (N_1538,N_1451,N_1415);
nand U1539 (N_1539,N_1430,N_1438);
nor U1540 (N_1540,N_1466,N_1436);
nand U1541 (N_1541,N_1492,N_1460);
or U1542 (N_1542,N_1420,N_1453);
or U1543 (N_1543,N_1406,N_1482);
or U1544 (N_1544,N_1428,N_1443);
nand U1545 (N_1545,N_1432,N_1403);
or U1546 (N_1546,N_1445,N_1454);
and U1547 (N_1547,N_1463,N_1456);
nand U1548 (N_1548,N_1435,N_1475);
nor U1549 (N_1549,N_1433,N_1476);
and U1550 (N_1550,N_1475,N_1455);
nand U1551 (N_1551,N_1402,N_1486);
nor U1552 (N_1552,N_1456,N_1481);
and U1553 (N_1553,N_1450,N_1400);
or U1554 (N_1554,N_1479,N_1487);
nand U1555 (N_1555,N_1439,N_1444);
and U1556 (N_1556,N_1449,N_1439);
or U1557 (N_1557,N_1408,N_1428);
or U1558 (N_1558,N_1443,N_1458);
or U1559 (N_1559,N_1488,N_1461);
nand U1560 (N_1560,N_1449,N_1459);
or U1561 (N_1561,N_1464,N_1445);
and U1562 (N_1562,N_1475,N_1492);
nor U1563 (N_1563,N_1449,N_1466);
and U1564 (N_1564,N_1456,N_1468);
or U1565 (N_1565,N_1491,N_1402);
nand U1566 (N_1566,N_1403,N_1488);
and U1567 (N_1567,N_1416,N_1462);
or U1568 (N_1568,N_1434,N_1462);
nand U1569 (N_1569,N_1466,N_1430);
nand U1570 (N_1570,N_1425,N_1444);
nand U1571 (N_1571,N_1468,N_1494);
nand U1572 (N_1572,N_1457,N_1435);
nand U1573 (N_1573,N_1471,N_1441);
or U1574 (N_1574,N_1442,N_1477);
and U1575 (N_1575,N_1491,N_1498);
and U1576 (N_1576,N_1405,N_1450);
nor U1577 (N_1577,N_1441,N_1410);
and U1578 (N_1578,N_1405,N_1431);
and U1579 (N_1579,N_1417,N_1464);
nand U1580 (N_1580,N_1484,N_1417);
or U1581 (N_1581,N_1403,N_1404);
nand U1582 (N_1582,N_1440,N_1492);
nor U1583 (N_1583,N_1461,N_1425);
or U1584 (N_1584,N_1496,N_1445);
nand U1585 (N_1585,N_1453,N_1431);
or U1586 (N_1586,N_1472,N_1411);
nor U1587 (N_1587,N_1471,N_1406);
nor U1588 (N_1588,N_1470,N_1425);
or U1589 (N_1589,N_1417,N_1491);
nand U1590 (N_1590,N_1429,N_1409);
nand U1591 (N_1591,N_1482,N_1420);
nor U1592 (N_1592,N_1430,N_1477);
or U1593 (N_1593,N_1412,N_1457);
or U1594 (N_1594,N_1440,N_1445);
nand U1595 (N_1595,N_1466,N_1421);
or U1596 (N_1596,N_1456,N_1417);
nor U1597 (N_1597,N_1434,N_1483);
nand U1598 (N_1598,N_1426,N_1414);
nand U1599 (N_1599,N_1465,N_1432);
and U1600 (N_1600,N_1565,N_1522);
nor U1601 (N_1601,N_1540,N_1506);
or U1602 (N_1602,N_1543,N_1520);
nand U1603 (N_1603,N_1571,N_1559);
nor U1604 (N_1604,N_1507,N_1517);
or U1605 (N_1605,N_1588,N_1596);
and U1606 (N_1606,N_1579,N_1508);
and U1607 (N_1607,N_1553,N_1592);
and U1608 (N_1608,N_1511,N_1597);
and U1609 (N_1609,N_1505,N_1510);
nand U1610 (N_1610,N_1555,N_1519);
or U1611 (N_1611,N_1504,N_1561);
and U1612 (N_1612,N_1581,N_1544);
nand U1613 (N_1613,N_1598,N_1590);
xnor U1614 (N_1614,N_1516,N_1568);
and U1615 (N_1615,N_1594,N_1583);
or U1616 (N_1616,N_1535,N_1591);
nand U1617 (N_1617,N_1567,N_1570);
nand U1618 (N_1618,N_1572,N_1552);
nor U1619 (N_1619,N_1500,N_1599);
nor U1620 (N_1620,N_1536,N_1533);
nand U1621 (N_1621,N_1595,N_1503);
nor U1622 (N_1622,N_1525,N_1528);
nand U1623 (N_1623,N_1542,N_1593);
nand U1624 (N_1624,N_1573,N_1512);
and U1625 (N_1625,N_1513,N_1545);
nor U1626 (N_1626,N_1589,N_1501);
nor U1627 (N_1627,N_1539,N_1547);
nor U1628 (N_1628,N_1514,N_1531);
nor U1629 (N_1629,N_1546,N_1576);
and U1630 (N_1630,N_1502,N_1538);
nand U1631 (N_1631,N_1518,N_1586);
and U1632 (N_1632,N_1530,N_1562);
nand U1633 (N_1633,N_1574,N_1532);
or U1634 (N_1634,N_1509,N_1537);
nand U1635 (N_1635,N_1563,N_1582);
xnor U1636 (N_1636,N_1578,N_1575);
or U1637 (N_1637,N_1549,N_1566);
or U1638 (N_1638,N_1526,N_1585);
nand U1639 (N_1639,N_1580,N_1527);
nor U1640 (N_1640,N_1564,N_1558);
nor U1641 (N_1641,N_1523,N_1587);
nand U1642 (N_1642,N_1548,N_1550);
nor U1643 (N_1643,N_1577,N_1557);
nand U1644 (N_1644,N_1541,N_1551);
nor U1645 (N_1645,N_1560,N_1556);
nor U1646 (N_1646,N_1529,N_1521);
and U1647 (N_1647,N_1534,N_1554);
or U1648 (N_1648,N_1515,N_1569);
nor U1649 (N_1649,N_1584,N_1524);
nor U1650 (N_1650,N_1583,N_1507);
nor U1651 (N_1651,N_1598,N_1510);
or U1652 (N_1652,N_1569,N_1502);
nor U1653 (N_1653,N_1543,N_1579);
nor U1654 (N_1654,N_1557,N_1508);
nor U1655 (N_1655,N_1568,N_1513);
or U1656 (N_1656,N_1571,N_1575);
nor U1657 (N_1657,N_1565,N_1595);
or U1658 (N_1658,N_1568,N_1578);
nor U1659 (N_1659,N_1538,N_1541);
nor U1660 (N_1660,N_1518,N_1557);
and U1661 (N_1661,N_1548,N_1537);
nand U1662 (N_1662,N_1524,N_1562);
nor U1663 (N_1663,N_1562,N_1519);
and U1664 (N_1664,N_1565,N_1598);
nor U1665 (N_1665,N_1581,N_1563);
and U1666 (N_1666,N_1547,N_1543);
nand U1667 (N_1667,N_1528,N_1591);
nand U1668 (N_1668,N_1534,N_1515);
or U1669 (N_1669,N_1558,N_1543);
or U1670 (N_1670,N_1559,N_1542);
and U1671 (N_1671,N_1501,N_1591);
nor U1672 (N_1672,N_1536,N_1537);
or U1673 (N_1673,N_1533,N_1520);
nand U1674 (N_1674,N_1549,N_1538);
or U1675 (N_1675,N_1511,N_1502);
or U1676 (N_1676,N_1598,N_1550);
or U1677 (N_1677,N_1556,N_1546);
nand U1678 (N_1678,N_1592,N_1532);
nand U1679 (N_1679,N_1574,N_1518);
nor U1680 (N_1680,N_1554,N_1596);
nor U1681 (N_1681,N_1560,N_1525);
and U1682 (N_1682,N_1545,N_1527);
nor U1683 (N_1683,N_1576,N_1506);
or U1684 (N_1684,N_1504,N_1518);
nand U1685 (N_1685,N_1510,N_1520);
and U1686 (N_1686,N_1521,N_1512);
nor U1687 (N_1687,N_1525,N_1529);
or U1688 (N_1688,N_1589,N_1591);
nand U1689 (N_1689,N_1503,N_1506);
and U1690 (N_1690,N_1537,N_1559);
nor U1691 (N_1691,N_1513,N_1511);
nor U1692 (N_1692,N_1575,N_1589);
and U1693 (N_1693,N_1517,N_1596);
nand U1694 (N_1694,N_1590,N_1546);
and U1695 (N_1695,N_1509,N_1559);
or U1696 (N_1696,N_1521,N_1510);
or U1697 (N_1697,N_1508,N_1592);
or U1698 (N_1698,N_1580,N_1512);
and U1699 (N_1699,N_1518,N_1513);
or U1700 (N_1700,N_1651,N_1643);
nand U1701 (N_1701,N_1639,N_1698);
nand U1702 (N_1702,N_1657,N_1663);
or U1703 (N_1703,N_1614,N_1658);
and U1704 (N_1704,N_1687,N_1638);
nand U1705 (N_1705,N_1670,N_1602);
or U1706 (N_1706,N_1624,N_1684);
or U1707 (N_1707,N_1612,N_1685);
or U1708 (N_1708,N_1634,N_1693);
or U1709 (N_1709,N_1616,N_1696);
and U1710 (N_1710,N_1610,N_1609);
and U1711 (N_1711,N_1622,N_1699);
nand U1712 (N_1712,N_1666,N_1647);
or U1713 (N_1713,N_1617,N_1674);
or U1714 (N_1714,N_1648,N_1686);
or U1715 (N_1715,N_1671,N_1653);
and U1716 (N_1716,N_1681,N_1646);
nand U1717 (N_1717,N_1636,N_1660);
nand U1718 (N_1718,N_1682,N_1601);
xor U1719 (N_1719,N_1652,N_1641);
or U1720 (N_1720,N_1659,N_1662);
and U1721 (N_1721,N_1623,N_1665);
or U1722 (N_1722,N_1697,N_1606);
and U1723 (N_1723,N_1667,N_1688);
and U1724 (N_1724,N_1618,N_1695);
or U1725 (N_1725,N_1604,N_1664);
nand U1726 (N_1726,N_1603,N_1615);
nor U1727 (N_1727,N_1627,N_1640);
and U1728 (N_1728,N_1613,N_1626);
or U1729 (N_1729,N_1644,N_1678);
and U1730 (N_1730,N_1669,N_1680);
nand U1731 (N_1731,N_1611,N_1628);
nor U1732 (N_1732,N_1621,N_1694);
and U1733 (N_1733,N_1654,N_1645);
and U1734 (N_1734,N_1677,N_1679);
and U1735 (N_1735,N_1661,N_1607);
and U1736 (N_1736,N_1675,N_1672);
nor U1737 (N_1737,N_1656,N_1683);
nand U1738 (N_1738,N_1690,N_1619);
and U1739 (N_1739,N_1691,N_1689);
and U1740 (N_1740,N_1673,N_1637);
and U1741 (N_1741,N_1692,N_1600);
or U1742 (N_1742,N_1649,N_1655);
nor U1743 (N_1743,N_1630,N_1629);
and U1744 (N_1744,N_1631,N_1668);
and U1745 (N_1745,N_1620,N_1625);
nor U1746 (N_1746,N_1642,N_1635);
nand U1747 (N_1747,N_1676,N_1633);
and U1748 (N_1748,N_1605,N_1608);
and U1749 (N_1749,N_1650,N_1632);
and U1750 (N_1750,N_1605,N_1613);
and U1751 (N_1751,N_1680,N_1614);
nor U1752 (N_1752,N_1622,N_1656);
nand U1753 (N_1753,N_1669,N_1611);
nor U1754 (N_1754,N_1660,N_1648);
nor U1755 (N_1755,N_1695,N_1676);
nand U1756 (N_1756,N_1674,N_1647);
nand U1757 (N_1757,N_1656,N_1619);
nand U1758 (N_1758,N_1620,N_1642);
nor U1759 (N_1759,N_1621,N_1612);
and U1760 (N_1760,N_1654,N_1688);
and U1761 (N_1761,N_1662,N_1654);
and U1762 (N_1762,N_1665,N_1633);
nor U1763 (N_1763,N_1607,N_1647);
xnor U1764 (N_1764,N_1638,N_1614);
nor U1765 (N_1765,N_1699,N_1633);
or U1766 (N_1766,N_1684,N_1602);
nor U1767 (N_1767,N_1671,N_1611);
nand U1768 (N_1768,N_1647,N_1645);
or U1769 (N_1769,N_1639,N_1605);
or U1770 (N_1770,N_1618,N_1660);
nor U1771 (N_1771,N_1658,N_1612);
or U1772 (N_1772,N_1624,N_1612);
or U1773 (N_1773,N_1643,N_1647);
or U1774 (N_1774,N_1692,N_1607);
nor U1775 (N_1775,N_1658,N_1697);
nand U1776 (N_1776,N_1693,N_1647);
nand U1777 (N_1777,N_1664,N_1639);
nand U1778 (N_1778,N_1669,N_1633);
and U1779 (N_1779,N_1619,N_1616);
and U1780 (N_1780,N_1608,N_1671);
nand U1781 (N_1781,N_1692,N_1667);
and U1782 (N_1782,N_1661,N_1632);
nand U1783 (N_1783,N_1601,N_1674);
and U1784 (N_1784,N_1611,N_1662);
or U1785 (N_1785,N_1656,N_1648);
nand U1786 (N_1786,N_1693,N_1661);
nand U1787 (N_1787,N_1676,N_1612);
or U1788 (N_1788,N_1612,N_1650);
and U1789 (N_1789,N_1605,N_1636);
or U1790 (N_1790,N_1605,N_1647);
and U1791 (N_1791,N_1606,N_1626);
and U1792 (N_1792,N_1651,N_1692);
or U1793 (N_1793,N_1667,N_1653);
and U1794 (N_1794,N_1622,N_1603);
nor U1795 (N_1795,N_1660,N_1650);
and U1796 (N_1796,N_1611,N_1639);
nor U1797 (N_1797,N_1609,N_1677);
nand U1798 (N_1798,N_1660,N_1601);
nand U1799 (N_1799,N_1633,N_1652);
or U1800 (N_1800,N_1774,N_1727);
nand U1801 (N_1801,N_1769,N_1782);
and U1802 (N_1802,N_1703,N_1738);
nand U1803 (N_1803,N_1734,N_1705);
nand U1804 (N_1804,N_1760,N_1779);
or U1805 (N_1805,N_1714,N_1710);
nor U1806 (N_1806,N_1787,N_1716);
nand U1807 (N_1807,N_1797,N_1790);
nor U1808 (N_1808,N_1746,N_1701);
and U1809 (N_1809,N_1742,N_1704);
or U1810 (N_1810,N_1750,N_1763);
nor U1811 (N_1811,N_1767,N_1768);
nand U1812 (N_1812,N_1748,N_1736);
and U1813 (N_1813,N_1783,N_1739);
and U1814 (N_1814,N_1761,N_1747);
and U1815 (N_1815,N_1793,N_1771);
xor U1816 (N_1816,N_1719,N_1786);
nor U1817 (N_1817,N_1702,N_1758);
and U1818 (N_1818,N_1711,N_1721);
nor U1819 (N_1819,N_1794,N_1720);
and U1820 (N_1820,N_1755,N_1775);
nor U1821 (N_1821,N_1780,N_1792);
nand U1822 (N_1822,N_1728,N_1725);
and U1823 (N_1823,N_1723,N_1729);
and U1824 (N_1824,N_1740,N_1752);
nor U1825 (N_1825,N_1743,N_1713);
or U1826 (N_1826,N_1730,N_1754);
and U1827 (N_1827,N_1722,N_1749);
nand U1828 (N_1828,N_1791,N_1766);
or U1829 (N_1829,N_1785,N_1757);
or U1830 (N_1830,N_1717,N_1788);
or U1831 (N_1831,N_1708,N_1715);
nand U1832 (N_1832,N_1765,N_1707);
nand U1833 (N_1833,N_1737,N_1781);
or U1834 (N_1834,N_1744,N_1709);
nand U1835 (N_1835,N_1762,N_1718);
nand U1836 (N_1836,N_1789,N_1773);
nor U1837 (N_1837,N_1776,N_1735);
and U1838 (N_1838,N_1745,N_1772);
and U1839 (N_1839,N_1770,N_1795);
and U1840 (N_1840,N_1753,N_1798);
nand U1841 (N_1841,N_1759,N_1796);
and U1842 (N_1842,N_1706,N_1784);
or U1843 (N_1843,N_1733,N_1732);
and U1844 (N_1844,N_1778,N_1764);
and U1845 (N_1845,N_1724,N_1799);
nor U1846 (N_1846,N_1712,N_1751);
or U1847 (N_1847,N_1700,N_1731);
or U1848 (N_1848,N_1726,N_1756);
nor U1849 (N_1849,N_1741,N_1777);
and U1850 (N_1850,N_1737,N_1713);
and U1851 (N_1851,N_1788,N_1756);
or U1852 (N_1852,N_1744,N_1786);
and U1853 (N_1853,N_1779,N_1793);
and U1854 (N_1854,N_1705,N_1736);
nand U1855 (N_1855,N_1739,N_1793);
nand U1856 (N_1856,N_1711,N_1739);
and U1857 (N_1857,N_1772,N_1730);
nand U1858 (N_1858,N_1758,N_1737);
or U1859 (N_1859,N_1733,N_1714);
and U1860 (N_1860,N_1781,N_1760);
nor U1861 (N_1861,N_1798,N_1731);
nor U1862 (N_1862,N_1745,N_1796);
nand U1863 (N_1863,N_1735,N_1764);
or U1864 (N_1864,N_1770,N_1747);
nand U1865 (N_1865,N_1700,N_1711);
nor U1866 (N_1866,N_1787,N_1734);
nor U1867 (N_1867,N_1746,N_1781);
and U1868 (N_1868,N_1783,N_1702);
or U1869 (N_1869,N_1752,N_1708);
and U1870 (N_1870,N_1723,N_1770);
nand U1871 (N_1871,N_1759,N_1785);
nor U1872 (N_1872,N_1702,N_1776);
nor U1873 (N_1873,N_1795,N_1764);
and U1874 (N_1874,N_1708,N_1726);
and U1875 (N_1875,N_1739,N_1708);
and U1876 (N_1876,N_1782,N_1733);
nor U1877 (N_1877,N_1795,N_1729);
or U1878 (N_1878,N_1763,N_1705);
and U1879 (N_1879,N_1788,N_1743);
xnor U1880 (N_1880,N_1746,N_1776);
nand U1881 (N_1881,N_1793,N_1783);
nand U1882 (N_1882,N_1720,N_1748);
and U1883 (N_1883,N_1775,N_1788);
nor U1884 (N_1884,N_1753,N_1785);
or U1885 (N_1885,N_1706,N_1756);
nor U1886 (N_1886,N_1751,N_1718);
nor U1887 (N_1887,N_1712,N_1792);
nand U1888 (N_1888,N_1784,N_1718);
nand U1889 (N_1889,N_1725,N_1749);
nand U1890 (N_1890,N_1780,N_1706);
nor U1891 (N_1891,N_1741,N_1748);
and U1892 (N_1892,N_1788,N_1757);
nor U1893 (N_1893,N_1782,N_1748);
and U1894 (N_1894,N_1705,N_1706);
and U1895 (N_1895,N_1708,N_1747);
nor U1896 (N_1896,N_1711,N_1709);
nand U1897 (N_1897,N_1758,N_1778);
or U1898 (N_1898,N_1775,N_1722);
nand U1899 (N_1899,N_1722,N_1799);
nand U1900 (N_1900,N_1854,N_1880);
nor U1901 (N_1901,N_1890,N_1878);
xnor U1902 (N_1902,N_1882,N_1851);
nor U1903 (N_1903,N_1828,N_1892);
nand U1904 (N_1904,N_1877,N_1849);
or U1905 (N_1905,N_1894,N_1840);
or U1906 (N_1906,N_1868,N_1856);
nor U1907 (N_1907,N_1887,N_1870);
nand U1908 (N_1908,N_1862,N_1842);
nand U1909 (N_1909,N_1844,N_1825);
xnor U1910 (N_1910,N_1822,N_1897);
nor U1911 (N_1911,N_1864,N_1826);
or U1912 (N_1912,N_1879,N_1865);
nor U1913 (N_1913,N_1835,N_1816);
nand U1914 (N_1914,N_1803,N_1881);
and U1915 (N_1915,N_1812,N_1801);
nor U1916 (N_1916,N_1841,N_1895);
and U1917 (N_1917,N_1839,N_1806);
nand U1918 (N_1918,N_1891,N_1867);
and U1919 (N_1919,N_1871,N_1836);
and U1920 (N_1920,N_1861,N_1809);
and U1921 (N_1921,N_1824,N_1843);
nand U1922 (N_1922,N_1850,N_1811);
or U1923 (N_1923,N_1834,N_1808);
nor U1924 (N_1924,N_1893,N_1875);
nor U1925 (N_1925,N_1860,N_1859);
or U1926 (N_1926,N_1819,N_1838);
nor U1927 (N_1927,N_1872,N_1857);
nor U1928 (N_1928,N_1853,N_1869);
or U1929 (N_1929,N_1896,N_1830);
and U1930 (N_1930,N_1848,N_1888);
or U1931 (N_1931,N_1863,N_1829);
or U1932 (N_1932,N_1813,N_1807);
and U1933 (N_1933,N_1846,N_1866);
nand U1934 (N_1934,N_1898,N_1889);
nand U1935 (N_1935,N_1804,N_1823);
or U1936 (N_1936,N_1820,N_1883);
nand U1937 (N_1937,N_1818,N_1852);
or U1938 (N_1938,N_1845,N_1800);
nand U1939 (N_1939,N_1858,N_1876);
and U1940 (N_1940,N_1847,N_1884);
or U1941 (N_1941,N_1885,N_1899);
and U1942 (N_1942,N_1831,N_1817);
or U1943 (N_1943,N_1821,N_1810);
or U1944 (N_1944,N_1805,N_1832);
nor U1945 (N_1945,N_1855,N_1827);
or U1946 (N_1946,N_1802,N_1873);
nand U1947 (N_1947,N_1814,N_1874);
and U1948 (N_1948,N_1833,N_1815);
nor U1949 (N_1949,N_1886,N_1837);
nor U1950 (N_1950,N_1881,N_1877);
xnor U1951 (N_1951,N_1813,N_1889);
nand U1952 (N_1952,N_1860,N_1821);
nand U1953 (N_1953,N_1816,N_1886);
nand U1954 (N_1954,N_1863,N_1871);
nand U1955 (N_1955,N_1840,N_1825);
nor U1956 (N_1956,N_1894,N_1816);
nand U1957 (N_1957,N_1874,N_1861);
and U1958 (N_1958,N_1893,N_1802);
or U1959 (N_1959,N_1892,N_1833);
nor U1960 (N_1960,N_1849,N_1889);
or U1961 (N_1961,N_1802,N_1833);
and U1962 (N_1962,N_1894,N_1887);
and U1963 (N_1963,N_1813,N_1857);
nor U1964 (N_1964,N_1827,N_1861);
or U1965 (N_1965,N_1879,N_1875);
xnor U1966 (N_1966,N_1881,N_1852);
and U1967 (N_1967,N_1860,N_1884);
and U1968 (N_1968,N_1811,N_1834);
nor U1969 (N_1969,N_1810,N_1899);
and U1970 (N_1970,N_1800,N_1869);
xor U1971 (N_1971,N_1814,N_1888);
nand U1972 (N_1972,N_1869,N_1892);
nor U1973 (N_1973,N_1833,N_1898);
nand U1974 (N_1974,N_1866,N_1887);
nand U1975 (N_1975,N_1807,N_1824);
nor U1976 (N_1976,N_1863,N_1887);
or U1977 (N_1977,N_1853,N_1868);
nand U1978 (N_1978,N_1897,N_1810);
nand U1979 (N_1979,N_1889,N_1830);
or U1980 (N_1980,N_1846,N_1822);
nor U1981 (N_1981,N_1870,N_1878);
nor U1982 (N_1982,N_1822,N_1864);
or U1983 (N_1983,N_1866,N_1854);
nand U1984 (N_1984,N_1884,N_1809);
or U1985 (N_1985,N_1896,N_1857);
nand U1986 (N_1986,N_1823,N_1881);
nor U1987 (N_1987,N_1858,N_1851);
or U1988 (N_1988,N_1836,N_1870);
and U1989 (N_1989,N_1895,N_1889);
nand U1990 (N_1990,N_1814,N_1847);
nand U1991 (N_1991,N_1819,N_1883);
nor U1992 (N_1992,N_1805,N_1808);
and U1993 (N_1993,N_1862,N_1828);
nor U1994 (N_1994,N_1812,N_1830);
nand U1995 (N_1995,N_1802,N_1886);
nand U1996 (N_1996,N_1836,N_1825);
or U1997 (N_1997,N_1893,N_1840);
and U1998 (N_1998,N_1896,N_1828);
xnor U1999 (N_1999,N_1895,N_1839);
nand U2000 (N_2000,N_1970,N_1983);
and U2001 (N_2001,N_1930,N_1936);
and U2002 (N_2002,N_1966,N_1987);
nand U2003 (N_2003,N_1939,N_1937);
and U2004 (N_2004,N_1918,N_1923);
xor U2005 (N_2005,N_1925,N_1948);
nand U2006 (N_2006,N_1932,N_1904);
and U2007 (N_2007,N_1974,N_1999);
nor U2008 (N_2008,N_1909,N_1913);
nor U2009 (N_2009,N_1986,N_1914);
nand U2010 (N_2010,N_1951,N_1993);
nand U2011 (N_2011,N_1997,N_1942);
nor U2012 (N_2012,N_1971,N_1921);
xor U2013 (N_2013,N_1962,N_1996);
nor U2014 (N_2014,N_1955,N_1905);
or U2015 (N_2015,N_1906,N_1958);
nor U2016 (N_2016,N_1928,N_1984);
nor U2017 (N_2017,N_1927,N_1964);
and U2018 (N_2018,N_1941,N_1926);
nor U2019 (N_2019,N_1985,N_1995);
and U2020 (N_2020,N_1929,N_1916);
or U2021 (N_2021,N_1960,N_1907);
nor U2022 (N_2022,N_1945,N_1947);
nor U2023 (N_2023,N_1900,N_1982);
nor U2024 (N_2024,N_1952,N_1963);
or U2025 (N_2025,N_1953,N_1949);
or U2026 (N_2026,N_1944,N_1959);
nand U2027 (N_2027,N_1910,N_1950);
and U2028 (N_2028,N_1917,N_1938);
or U2029 (N_2029,N_1975,N_1922);
nor U2030 (N_2030,N_1979,N_1903);
and U2031 (N_2031,N_1912,N_1943);
and U2032 (N_2032,N_1931,N_1954);
or U2033 (N_2033,N_1994,N_1911);
and U2034 (N_2034,N_1957,N_1969);
nor U2035 (N_2035,N_1977,N_1934);
nor U2036 (N_2036,N_1973,N_1981);
nand U2037 (N_2037,N_1902,N_1961);
and U2038 (N_2038,N_1901,N_1976);
and U2039 (N_2039,N_1980,N_1935);
nand U2040 (N_2040,N_1967,N_1915);
xnor U2041 (N_2041,N_1978,N_1908);
nand U2042 (N_2042,N_1988,N_1920);
and U2043 (N_2043,N_1998,N_1965);
nand U2044 (N_2044,N_1940,N_1956);
nor U2045 (N_2045,N_1946,N_1924);
nand U2046 (N_2046,N_1990,N_1991);
nand U2047 (N_2047,N_1919,N_1968);
nor U2048 (N_2048,N_1972,N_1933);
or U2049 (N_2049,N_1992,N_1989);
and U2050 (N_2050,N_1924,N_1970);
nand U2051 (N_2051,N_1990,N_1926);
and U2052 (N_2052,N_1990,N_1995);
and U2053 (N_2053,N_1974,N_1922);
or U2054 (N_2054,N_1988,N_1998);
xnor U2055 (N_2055,N_1906,N_1984);
nand U2056 (N_2056,N_1934,N_1974);
and U2057 (N_2057,N_1968,N_1999);
or U2058 (N_2058,N_1939,N_1996);
nand U2059 (N_2059,N_1957,N_1986);
nor U2060 (N_2060,N_1989,N_1929);
nor U2061 (N_2061,N_1970,N_1916);
nand U2062 (N_2062,N_1913,N_1929);
nor U2063 (N_2063,N_1983,N_1981);
and U2064 (N_2064,N_1966,N_1910);
xnor U2065 (N_2065,N_1941,N_1988);
nand U2066 (N_2066,N_1926,N_1902);
nand U2067 (N_2067,N_1904,N_1994);
or U2068 (N_2068,N_1993,N_1950);
and U2069 (N_2069,N_1989,N_1914);
and U2070 (N_2070,N_1984,N_1900);
and U2071 (N_2071,N_1956,N_1996);
and U2072 (N_2072,N_1949,N_1910);
and U2073 (N_2073,N_1987,N_1925);
nor U2074 (N_2074,N_1941,N_1962);
nand U2075 (N_2075,N_1973,N_1988);
nand U2076 (N_2076,N_1969,N_1914);
and U2077 (N_2077,N_1989,N_1961);
nand U2078 (N_2078,N_1991,N_1945);
nand U2079 (N_2079,N_1919,N_1963);
or U2080 (N_2080,N_1973,N_1963);
or U2081 (N_2081,N_1991,N_1959);
and U2082 (N_2082,N_1977,N_1920);
nor U2083 (N_2083,N_1942,N_1919);
nor U2084 (N_2084,N_1901,N_1968);
nor U2085 (N_2085,N_1956,N_1972);
nand U2086 (N_2086,N_1929,N_1963);
nor U2087 (N_2087,N_1917,N_1949);
or U2088 (N_2088,N_1906,N_1943);
or U2089 (N_2089,N_1943,N_1900);
or U2090 (N_2090,N_1939,N_1979);
nand U2091 (N_2091,N_1939,N_1944);
and U2092 (N_2092,N_1926,N_1947);
nand U2093 (N_2093,N_1951,N_1911);
and U2094 (N_2094,N_1989,N_1902);
nor U2095 (N_2095,N_1941,N_1978);
nor U2096 (N_2096,N_1944,N_1978);
nand U2097 (N_2097,N_1913,N_1947);
and U2098 (N_2098,N_1966,N_1960);
nor U2099 (N_2099,N_1913,N_1956);
nor U2100 (N_2100,N_2031,N_2097);
nor U2101 (N_2101,N_2079,N_2004);
nand U2102 (N_2102,N_2046,N_2027);
or U2103 (N_2103,N_2082,N_2006);
or U2104 (N_2104,N_2073,N_2072);
nand U2105 (N_2105,N_2066,N_2005);
and U2106 (N_2106,N_2094,N_2009);
or U2107 (N_2107,N_2019,N_2058);
or U2108 (N_2108,N_2098,N_2099);
and U2109 (N_2109,N_2017,N_2076);
xor U2110 (N_2110,N_2010,N_2016);
and U2111 (N_2111,N_2041,N_2096);
xor U2112 (N_2112,N_2008,N_2038);
or U2113 (N_2113,N_2007,N_2028);
nor U2114 (N_2114,N_2000,N_2040);
nor U2115 (N_2115,N_2090,N_2049);
or U2116 (N_2116,N_2035,N_2033);
nand U2117 (N_2117,N_2060,N_2011);
and U2118 (N_2118,N_2020,N_2059);
nand U2119 (N_2119,N_2095,N_2069);
and U2120 (N_2120,N_2071,N_2022);
nor U2121 (N_2121,N_2037,N_2088);
nand U2122 (N_2122,N_2064,N_2055);
or U2123 (N_2123,N_2052,N_2034);
and U2124 (N_2124,N_2061,N_2014);
and U2125 (N_2125,N_2081,N_2070);
and U2126 (N_2126,N_2021,N_2065);
and U2127 (N_2127,N_2089,N_2057);
nand U2128 (N_2128,N_2003,N_2023);
nor U2129 (N_2129,N_2047,N_2043);
nand U2130 (N_2130,N_2056,N_2093);
nand U2131 (N_2131,N_2083,N_2002);
or U2132 (N_2132,N_2045,N_2025);
and U2133 (N_2133,N_2015,N_2091);
or U2134 (N_2134,N_2032,N_2054);
nor U2135 (N_2135,N_2050,N_2030);
nor U2136 (N_2136,N_2024,N_2001);
or U2137 (N_2137,N_2087,N_2026);
xor U2138 (N_2138,N_2086,N_2084);
or U2139 (N_2139,N_2044,N_2077);
nand U2140 (N_2140,N_2051,N_2074);
nand U2141 (N_2141,N_2078,N_2080);
nand U2142 (N_2142,N_2018,N_2036);
nor U2143 (N_2143,N_2068,N_2053);
and U2144 (N_2144,N_2075,N_2067);
nor U2145 (N_2145,N_2012,N_2063);
nor U2146 (N_2146,N_2013,N_2048);
and U2147 (N_2147,N_2029,N_2062);
nand U2148 (N_2148,N_2085,N_2042);
nand U2149 (N_2149,N_2092,N_2039);
and U2150 (N_2150,N_2062,N_2072);
or U2151 (N_2151,N_2072,N_2036);
and U2152 (N_2152,N_2090,N_2059);
or U2153 (N_2153,N_2012,N_2080);
nor U2154 (N_2154,N_2049,N_2095);
nor U2155 (N_2155,N_2004,N_2020);
and U2156 (N_2156,N_2064,N_2080);
nand U2157 (N_2157,N_2062,N_2098);
or U2158 (N_2158,N_2031,N_2070);
nor U2159 (N_2159,N_2027,N_2051);
xor U2160 (N_2160,N_2016,N_2033);
nand U2161 (N_2161,N_2078,N_2074);
and U2162 (N_2162,N_2078,N_2069);
or U2163 (N_2163,N_2061,N_2007);
or U2164 (N_2164,N_2058,N_2002);
nor U2165 (N_2165,N_2003,N_2020);
and U2166 (N_2166,N_2053,N_2056);
nand U2167 (N_2167,N_2028,N_2045);
nor U2168 (N_2168,N_2002,N_2053);
nand U2169 (N_2169,N_2063,N_2046);
nand U2170 (N_2170,N_2018,N_2098);
nand U2171 (N_2171,N_2060,N_2053);
nor U2172 (N_2172,N_2058,N_2098);
nor U2173 (N_2173,N_2028,N_2020);
xor U2174 (N_2174,N_2046,N_2039);
nor U2175 (N_2175,N_2063,N_2061);
and U2176 (N_2176,N_2068,N_2011);
and U2177 (N_2177,N_2032,N_2068);
nor U2178 (N_2178,N_2043,N_2027);
xnor U2179 (N_2179,N_2011,N_2015);
nor U2180 (N_2180,N_2061,N_2001);
or U2181 (N_2181,N_2037,N_2067);
nand U2182 (N_2182,N_2085,N_2026);
xnor U2183 (N_2183,N_2012,N_2033);
nor U2184 (N_2184,N_2021,N_2091);
or U2185 (N_2185,N_2076,N_2086);
and U2186 (N_2186,N_2080,N_2016);
nand U2187 (N_2187,N_2085,N_2044);
or U2188 (N_2188,N_2040,N_2057);
nand U2189 (N_2189,N_2056,N_2085);
nand U2190 (N_2190,N_2018,N_2011);
or U2191 (N_2191,N_2051,N_2083);
nand U2192 (N_2192,N_2024,N_2092);
or U2193 (N_2193,N_2086,N_2003);
and U2194 (N_2194,N_2051,N_2013);
nand U2195 (N_2195,N_2093,N_2014);
nor U2196 (N_2196,N_2033,N_2080);
or U2197 (N_2197,N_2091,N_2058);
and U2198 (N_2198,N_2095,N_2066);
nor U2199 (N_2199,N_2043,N_2037);
or U2200 (N_2200,N_2114,N_2124);
or U2201 (N_2201,N_2168,N_2105);
nor U2202 (N_2202,N_2156,N_2109);
or U2203 (N_2203,N_2133,N_2166);
and U2204 (N_2204,N_2189,N_2120);
and U2205 (N_2205,N_2137,N_2104);
nor U2206 (N_2206,N_2138,N_2106);
nor U2207 (N_2207,N_2140,N_2192);
and U2208 (N_2208,N_2171,N_2194);
nand U2209 (N_2209,N_2110,N_2180);
nor U2210 (N_2210,N_2157,N_2116);
and U2211 (N_2211,N_2103,N_2115);
or U2212 (N_2212,N_2172,N_2163);
and U2213 (N_2213,N_2198,N_2151);
nand U2214 (N_2214,N_2161,N_2149);
or U2215 (N_2215,N_2134,N_2165);
and U2216 (N_2216,N_2148,N_2119);
and U2217 (N_2217,N_2129,N_2178);
nor U2218 (N_2218,N_2136,N_2175);
or U2219 (N_2219,N_2145,N_2170);
nand U2220 (N_2220,N_2185,N_2152);
or U2221 (N_2221,N_2186,N_2108);
and U2222 (N_2222,N_2118,N_2153);
or U2223 (N_2223,N_2167,N_2142);
or U2224 (N_2224,N_2112,N_2121);
nand U2225 (N_2225,N_2130,N_2117);
nand U2226 (N_2226,N_2143,N_2113);
or U2227 (N_2227,N_2164,N_2176);
or U2228 (N_2228,N_2139,N_2193);
or U2229 (N_2229,N_2146,N_2190);
nor U2230 (N_2230,N_2158,N_2101);
or U2231 (N_2231,N_2183,N_2174);
and U2232 (N_2232,N_2126,N_2160);
nand U2233 (N_2233,N_2127,N_2122);
nand U2234 (N_2234,N_2141,N_2154);
or U2235 (N_2235,N_2135,N_2144);
or U2236 (N_2236,N_2182,N_2125);
or U2237 (N_2237,N_2191,N_2188);
or U2238 (N_2238,N_2131,N_2123);
or U2239 (N_2239,N_2169,N_2184);
and U2240 (N_2240,N_2181,N_2102);
or U2241 (N_2241,N_2159,N_2199);
nor U2242 (N_2242,N_2177,N_2179);
nor U2243 (N_2243,N_2100,N_2173);
and U2244 (N_2244,N_2155,N_2128);
and U2245 (N_2245,N_2197,N_2107);
or U2246 (N_2246,N_2147,N_2150);
and U2247 (N_2247,N_2196,N_2111);
nor U2248 (N_2248,N_2132,N_2187);
nor U2249 (N_2249,N_2195,N_2162);
and U2250 (N_2250,N_2160,N_2111);
nor U2251 (N_2251,N_2181,N_2180);
and U2252 (N_2252,N_2189,N_2157);
nor U2253 (N_2253,N_2183,N_2135);
nand U2254 (N_2254,N_2177,N_2154);
nand U2255 (N_2255,N_2108,N_2140);
xnor U2256 (N_2256,N_2129,N_2111);
nand U2257 (N_2257,N_2120,N_2182);
nor U2258 (N_2258,N_2147,N_2130);
nand U2259 (N_2259,N_2149,N_2194);
or U2260 (N_2260,N_2101,N_2193);
and U2261 (N_2261,N_2123,N_2171);
nor U2262 (N_2262,N_2161,N_2166);
or U2263 (N_2263,N_2199,N_2107);
and U2264 (N_2264,N_2151,N_2100);
or U2265 (N_2265,N_2102,N_2106);
and U2266 (N_2266,N_2119,N_2125);
and U2267 (N_2267,N_2146,N_2116);
nand U2268 (N_2268,N_2158,N_2117);
nor U2269 (N_2269,N_2116,N_2123);
nand U2270 (N_2270,N_2198,N_2126);
nor U2271 (N_2271,N_2175,N_2181);
or U2272 (N_2272,N_2181,N_2197);
and U2273 (N_2273,N_2106,N_2175);
and U2274 (N_2274,N_2181,N_2120);
nand U2275 (N_2275,N_2149,N_2129);
and U2276 (N_2276,N_2171,N_2135);
nor U2277 (N_2277,N_2150,N_2187);
and U2278 (N_2278,N_2172,N_2180);
xor U2279 (N_2279,N_2128,N_2164);
nand U2280 (N_2280,N_2161,N_2146);
and U2281 (N_2281,N_2125,N_2146);
or U2282 (N_2282,N_2169,N_2133);
nand U2283 (N_2283,N_2130,N_2151);
nor U2284 (N_2284,N_2117,N_2172);
and U2285 (N_2285,N_2187,N_2179);
and U2286 (N_2286,N_2159,N_2167);
and U2287 (N_2287,N_2103,N_2188);
and U2288 (N_2288,N_2128,N_2178);
nor U2289 (N_2289,N_2145,N_2192);
xor U2290 (N_2290,N_2184,N_2158);
xnor U2291 (N_2291,N_2197,N_2128);
xnor U2292 (N_2292,N_2172,N_2139);
and U2293 (N_2293,N_2167,N_2146);
and U2294 (N_2294,N_2170,N_2127);
and U2295 (N_2295,N_2144,N_2163);
nor U2296 (N_2296,N_2187,N_2145);
or U2297 (N_2297,N_2107,N_2198);
and U2298 (N_2298,N_2131,N_2127);
or U2299 (N_2299,N_2128,N_2123);
or U2300 (N_2300,N_2270,N_2237);
or U2301 (N_2301,N_2289,N_2290);
and U2302 (N_2302,N_2254,N_2216);
or U2303 (N_2303,N_2284,N_2224);
nor U2304 (N_2304,N_2259,N_2213);
and U2305 (N_2305,N_2258,N_2241);
nand U2306 (N_2306,N_2245,N_2280);
or U2307 (N_2307,N_2266,N_2288);
or U2308 (N_2308,N_2243,N_2219);
or U2309 (N_2309,N_2233,N_2293);
or U2310 (N_2310,N_2235,N_2208);
and U2311 (N_2311,N_2274,N_2217);
and U2312 (N_2312,N_2262,N_2287);
nand U2313 (N_2313,N_2220,N_2297);
or U2314 (N_2314,N_2205,N_2294);
or U2315 (N_2315,N_2200,N_2257);
nor U2316 (N_2316,N_2272,N_2283);
and U2317 (N_2317,N_2279,N_2248);
or U2318 (N_2318,N_2201,N_2285);
nor U2319 (N_2319,N_2204,N_2232);
or U2320 (N_2320,N_2207,N_2267);
and U2321 (N_2321,N_2271,N_2227);
or U2322 (N_2322,N_2240,N_2221);
and U2323 (N_2323,N_2228,N_2250);
and U2324 (N_2324,N_2296,N_2281);
and U2325 (N_2325,N_2212,N_2222);
and U2326 (N_2326,N_2242,N_2218);
or U2327 (N_2327,N_2234,N_2278);
nor U2328 (N_2328,N_2295,N_2273);
and U2329 (N_2329,N_2282,N_2268);
nand U2330 (N_2330,N_2256,N_2249);
nor U2331 (N_2331,N_2260,N_2261);
xor U2332 (N_2332,N_2223,N_2202);
nor U2333 (N_2333,N_2229,N_2251);
nand U2334 (N_2334,N_2264,N_2238);
and U2335 (N_2335,N_2230,N_2252);
nand U2336 (N_2336,N_2247,N_2265);
nand U2337 (N_2337,N_2236,N_2209);
or U2338 (N_2338,N_2210,N_2298);
or U2339 (N_2339,N_2214,N_2286);
nor U2340 (N_2340,N_2225,N_2263);
and U2341 (N_2341,N_2299,N_2269);
nand U2342 (N_2342,N_2277,N_2203);
and U2343 (N_2343,N_2255,N_2244);
and U2344 (N_2344,N_2292,N_2231);
nor U2345 (N_2345,N_2211,N_2239);
or U2346 (N_2346,N_2246,N_2253);
nor U2347 (N_2347,N_2291,N_2206);
or U2348 (N_2348,N_2226,N_2215);
or U2349 (N_2349,N_2276,N_2275);
and U2350 (N_2350,N_2289,N_2214);
xnor U2351 (N_2351,N_2296,N_2216);
and U2352 (N_2352,N_2250,N_2209);
and U2353 (N_2353,N_2299,N_2284);
or U2354 (N_2354,N_2212,N_2268);
nand U2355 (N_2355,N_2229,N_2274);
nand U2356 (N_2356,N_2286,N_2283);
nand U2357 (N_2357,N_2261,N_2236);
nor U2358 (N_2358,N_2253,N_2245);
and U2359 (N_2359,N_2276,N_2201);
or U2360 (N_2360,N_2232,N_2212);
or U2361 (N_2361,N_2201,N_2279);
nand U2362 (N_2362,N_2286,N_2274);
nor U2363 (N_2363,N_2222,N_2244);
xor U2364 (N_2364,N_2269,N_2238);
nand U2365 (N_2365,N_2234,N_2292);
or U2366 (N_2366,N_2264,N_2202);
nor U2367 (N_2367,N_2241,N_2267);
and U2368 (N_2368,N_2266,N_2225);
and U2369 (N_2369,N_2288,N_2201);
or U2370 (N_2370,N_2276,N_2243);
or U2371 (N_2371,N_2281,N_2273);
nor U2372 (N_2372,N_2295,N_2205);
or U2373 (N_2373,N_2269,N_2227);
and U2374 (N_2374,N_2206,N_2253);
or U2375 (N_2375,N_2238,N_2217);
and U2376 (N_2376,N_2287,N_2225);
or U2377 (N_2377,N_2213,N_2223);
nor U2378 (N_2378,N_2248,N_2202);
or U2379 (N_2379,N_2291,N_2266);
nor U2380 (N_2380,N_2206,N_2293);
xnor U2381 (N_2381,N_2298,N_2250);
and U2382 (N_2382,N_2201,N_2263);
or U2383 (N_2383,N_2242,N_2216);
nor U2384 (N_2384,N_2267,N_2211);
nor U2385 (N_2385,N_2279,N_2204);
nand U2386 (N_2386,N_2291,N_2239);
nor U2387 (N_2387,N_2223,N_2230);
nand U2388 (N_2388,N_2263,N_2228);
nand U2389 (N_2389,N_2237,N_2288);
nand U2390 (N_2390,N_2286,N_2243);
or U2391 (N_2391,N_2252,N_2281);
nand U2392 (N_2392,N_2218,N_2292);
nor U2393 (N_2393,N_2239,N_2279);
nand U2394 (N_2394,N_2231,N_2275);
and U2395 (N_2395,N_2207,N_2284);
nor U2396 (N_2396,N_2223,N_2299);
nor U2397 (N_2397,N_2234,N_2229);
and U2398 (N_2398,N_2257,N_2248);
or U2399 (N_2399,N_2290,N_2296);
nand U2400 (N_2400,N_2343,N_2394);
and U2401 (N_2401,N_2345,N_2395);
nand U2402 (N_2402,N_2300,N_2338);
or U2403 (N_2403,N_2302,N_2348);
or U2404 (N_2404,N_2362,N_2396);
nor U2405 (N_2405,N_2352,N_2382);
and U2406 (N_2406,N_2399,N_2373);
nor U2407 (N_2407,N_2366,N_2328);
nand U2408 (N_2408,N_2368,N_2379);
or U2409 (N_2409,N_2307,N_2329);
nand U2410 (N_2410,N_2372,N_2390);
or U2411 (N_2411,N_2321,N_2367);
nand U2412 (N_2412,N_2374,N_2391);
nand U2413 (N_2413,N_2375,N_2325);
nor U2414 (N_2414,N_2357,N_2317);
or U2415 (N_2415,N_2380,N_2324);
or U2416 (N_2416,N_2312,N_2347);
nor U2417 (N_2417,N_2330,N_2310);
and U2418 (N_2418,N_2377,N_2322);
and U2419 (N_2419,N_2359,N_2356);
nand U2420 (N_2420,N_2360,N_2311);
nand U2421 (N_2421,N_2384,N_2364);
nand U2422 (N_2422,N_2376,N_2326);
nand U2423 (N_2423,N_2378,N_2354);
or U2424 (N_2424,N_2303,N_2398);
nand U2425 (N_2425,N_2316,N_2351);
and U2426 (N_2426,N_2393,N_2331);
nor U2427 (N_2427,N_2301,N_2385);
nand U2428 (N_2428,N_2386,N_2370);
and U2429 (N_2429,N_2342,N_2340);
nand U2430 (N_2430,N_2349,N_2355);
nor U2431 (N_2431,N_2309,N_2344);
and U2432 (N_2432,N_2335,N_2369);
nand U2433 (N_2433,N_2392,N_2350);
and U2434 (N_2434,N_2320,N_2336);
or U2435 (N_2435,N_2397,N_2339);
or U2436 (N_2436,N_2341,N_2315);
or U2437 (N_2437,N_2365,N_2327);
nor U2438 (N_2438,N_2353,N_2306);
nand U2439 (N_2439,N_2318,N_2388);
or U2440 (N_2440,N_2387,N_2304);
and U2441 (N_2441,N_2319,N_2308);
nand U2442 (N_2442,N_2334,N_2305);
nand U2443 (N_2443,N_2381,N_2361);
nand U2444 (N_2444,N_2314,N_2346);
xor U2445 (N_2445,N_2323,N_2313);
nand U2446 (N_2446,N_2389,N_2333);
or U2447 (N_2447,N_2371,N_2332);
nor U2448 (N_2448,N_2363,N_2337);
and U2449 (N_2449,N_2358,N_2383);
nand U2450 (N_2450,N_2377,N_2391);
nor U2451 (N_2451,N_2304,N_2363);
nor U2452 (N_2452,N_2398,N_2360);
nor U2453 (N_2453,N_2331,N_2371);
or U2454 (N_2454,N_2309,N_2356);
nand U2455 (N_2455,N_2327,N_2335);
nor U2456 (N_2456,N_2323,N_2359);
xor U2457 (N_2457,N_2344,N_2314);
or U2458 (N_2458,N_2373,N_2337);
xnor U2459 (N_2459,N_2387,N_2365);
nand U2460 (N_2460,N_2361,N_2320);
nor U2461 (N_2461,N_2305,N_2348);
or U2462 (N_2462,N_2327,N_2399);
nand U2463 (N_2463,N_2370,N_2395);
nand U2464 (N_2464,N_2309,N_2390);
or U2465 (N_2465,N_2326,N_2380);
nor U2466 (N_2466,N_2399,N_2309);
nand U2467 (N_2467,N_2315,N_2366);
nand U2468 (N_2468,N_2323,N_2398);
or U2469 (N_2469,N_2377,N_2337);
nor U2470 (N_2470,N_2389,N_2388);
nand U2471 (N_2471,N_2333,N_2384);
nand U2472 (N_2472,N_2361,N_2305);
nor U2473 (N_2473,N_2359,N_2340);
nand U2474 (N_2474,N_2396,N_2341);
or U2475 (N_2475,N_2392,N_2351);
nor U2476 (N_2476,N_2385,N_2302);
and U2477 (N_2477,N_2330,N_2375);
nor U2478 (N_2478,N_2350,N_2361);
or U2479 (N_2479,N_2374,N_2381);
nand U2480 (N_2480,N_2354,N_2377);
nand U2481 (N_2481,N_2396,N_2340);
and U2482 (N_2482,N_2395,N_2388);
nor U2483 (N_2483,N_2304,N_2392);
and U2484 (N_2484,N_2352,N_2303);
nand U2485 (N_2485,N_2350,N_2348);
or U2486 (N_2486,N_2396,N_2354);
nor U2487 (N_2487,N_2383,N_2348);
or U2488 (N_2488,N_2322,N_2383);
nand U2489 (N_2489,N_2335,N_2319);
nor U2490 (N_2490,N_2351,N_2326);
and U2491 (N_2491,N_2395,N_2391);
or U2492 (N_2492,N_2319,N_2391);
nor U2493 (N_2493,N_2356,N_2306);
or U2494 (N_2494,N_2301,N_2389);
or U2495 (N_2495,N_2362,N_2369);
nand U2496 (N_2496,N_2327,N_2304);
nor U2497 (N_2497,N_2329,N_2344);
nand U2498 (N_2498,N_2389,N_2366);
or U2499 (N_2499,N_2351,N_2348);
or U2500 (N_2500,N_2447,N_2445);
and U2501 (N_2501,N_2454,N_2426);
or U2502 (N_2502,N_2484,N_2449);
and U2503 (N_2503,N_2451,N_2436);
nand U2504 (N_2504,N_2408,N_2464);
and U2505 (N_2505,N_2425,N_2406);
and U2506 (N_2506,N_2477,N_2486);
nor U2507 (N_2507,N_2429,N_2424);
nand U2508 (N_2508,N_2432,N_2401);
or U2509 (N_2509,N_2440,N_2453);
nor U2510 (N_2510,N_2472,N_2492);
nor U2511 (N_2511,N_2411,N_2413);
or U2512 (N_2512,N_2405,N_2482);
nand U2513 (N_2513,N_2452,N_2473);
nor U2514 (N_2514,N_2459,N_2410);
nor U2515 (N_2515,N_2433,N_2443);
nand U2516 (N_2516,N_2469,N_2437);
nor U2517 (N_2517,N_2499,N_2404);
nor U2518 (N_2518,N_2466,N_2495);
and U2519 (N_2519,N_2418,N_2479);
and U2520 (N_2520,N_2471,N_2434);
nand U2521 (N_2521,N_2483,N_2465);
or U2522 (N_2522,N_2496,N_2497);
nand U2523 (N_2523,N_2430,N_2460);
or U2524 (N_2524,N_2441,N_2403);
nand U2525 (N_2525,N_2455,N_2474);
nand U2526 (N_2526,N_2476,N_2416);
nor U2527 (N_2527,N_2415,N_2463);
nand U2528 (N_2528,N_2450,N_2468);
nand U2529 (N_2529,N_2491,N_2428);
xnor U2530 (N_2530,N_2470,N_2481);
xnor U2531 (N_2531,N_2417,N_2480);
xor U2532 (N_2532,N_2462,N_2427);
nor U2533 (N_2533,N_2412,N_2438);
nand U2534 (N_2534,N_2435,N_2414);
nand U2535 (N_2535,N_2490,N_2488);
nor U2536 (N_2536,N_2494,N_2420);
nand U2537 (N_2537,N_2467,N_2498);
and U2538 (N_2538,N_2475,N_2407);
nor U2539 (N_2539,N_2446,N_2422);
or U2540 (N_2540,N_2457,N_2485);
nor U2541 (N_2541,N_2442,N_2444);
nand U2542 (N_2542,N_2431,N_2409);
and U2543 (N_2543,N_2419,N_2478);
nand U2544 (N_2544,N_2421,N_2423);
nand U2545 (N_2545,N_2487,N_2448);
nor U2546 (N_2546,N_2402,N_2458);
and U2547 (N_2547,N_2493,N_2439);
or U2548 (N_2548,N_2461,N_2400);
or U2549 (N_2549,N_2489,N_2456);
and U2550 (N_2550,N_2487,N_2466);
nor U2551 (N_2551,N_2488,N_2432);
or U2552 (N_2552,N_2460,N_2434);
or U2553 (N_2553,N_2496,N_2474);
nor U2554 (N_2554,N_2445,N_2455);
nand U2555 (N_2555,N_2440,N_2459);
nand U2556 (N_2556,N_2400,N_2458);
and U2557 (N_2557,N_2400,N_2401);
and U2558 (N_2558,N_2452,N_2427);
nand U2559 (N_2559,N_2463,N_2432);
nor U2560 (N_2560,N_2449,N_2473);
and U2561 (N_2561,N_2415,N_2420);
nand U2562 (N_2562,N_2498,N_2471);
or U2563 (N_2563,N_2422,N_2462);
nand U2564 (N_2564,N_2447,N_2442);
nor U2565 (N_2565,N_2411,N_2448);
or U2566 (N_2566,N_2483,N_2496);
and U2567 (N_2567,N_2420,N_2439);
and U2568 (N_2568,N_2475,N_2479);
or U2569 (N_2569,N_2415,N_2466);
or U2570 (N_2570,N_2466,N_2418);
nand U2571 (N_2571,N_2413,N_2462);
nand U2572 (N_2572,N_2469,N_2456);
xnor U2573 (N_2573,N_2407,N_2448);
and U2574 (N_2574,N_2474,N_2414);
and U2575 (N_2575,N_2473,N_2476);
or U2576 (N_2576,N_2426,N_2414);
and U2577 (N_2577,N_2410,N_2421);
or U2578 (N_2578,N_2455,N_2453);
nor U2579 (N_2579,N_2495,N_2481);
xnor U2580 (N_2580,N_2482,N_2467);
or U2581 (N_2581,N_2416,N_2417);
nor U2582 (N_2582,N_2436,N_2455);
and U2583 (N_2583,N_2447,N_2478);
or U2584 (N_2584,N_2444,N_2409);
nand U2585 (N_2585,N_2415,N_2425);
nor U2586 (N_2586,N_2466,N_2455);
or U2587 (N_2587,N_2484,N_2499);
nor U2588 (N_2588,N_2482,N_2492);
or U2589 (N_2589,N_2433,N_2445);
nor U2590 (N_2590,N_2418,N_2430);
nor U2591 (N_2591,N_2414,N_2479);
and U2592 (N_2592,N_2426,N_2455);
or U2593 (N_2593,N_2407,N_2439);
nand U2594 (N_2594,N_2485,N_2448);
nand U2595 (N_2595,N_2434,N_2425);
and U2596 (N_2596,N_2446,N_2483);
or U2597 (N_2597,N_2485,N_2498);
nand U2598 (N_2598,N_2428,N_2418);
nor U2599 (N_2599,N_2426,N_2433);
or U2600 (N_2600,N_2581,N_2534);
or U2601 (N_2601,N_2503,N_2579);
and U2602 (N_2602,N_2561,N_2514);
nand U2603 (N_2603,N_2539,N_2596);
nand U2604 (N_2604,N_2542,N_2516);
or U2605 (N_2605,N_2520,N_2574);
or U2606 (N_2606,N_2583,N_2522);
nand U2607 (N_2607,N_2598,N_2587);
nor U2608 (N_2608,N_2575,N_2535);
nor U2609 (N_2609,N_2549,N_2527);
nand U2610 (N_2610,N_2590,N_2571);
nand U2611 (N_2611,N_2592,N_2588);
nand U2612 (N_2612,N_2566,N_2585);
and U2613 (N_2613,N_2543,N_2524);
and U2614 (N_2614,N_2538,N_2594);
nand U2615 (N_2615,N_2562,N_2544);
nor U2616 (N_2616,N_2504,N_2545);
nor U2617 (N_2617,N_2572,N_2597);
nand U2618 (N_2618,N_2536,N_2576);
xor U2619 (N_2619,N_2565,N_2507);
or U2620 (N_2620,N_2593,N_2586);
or U2621 (N_2621,N_2523,N_2532);
and U2622 (N_2622,N_2553,N_2518);
nand U2623 (N_2623,N_2501,N_2591);
and U2624 (N_2624,N_2556,N_2580);
and U2625 (N_2625,N_2567,N_2506);
and U2626 (N_2626,N_2570,N_2560);
nand U2627 (N_2627,N_2552,N_2533);
or U2628 (N_2628,N_2589,N_2568);
or U2629 (N_2629,N_2564,N_2546);
or U2630 (N_2630,N_2537,N_2577);
nand U2631 (N_2631,N_2510,N_2540);
nor U2632 (N_2632,N_2530,N_2569);
or U2633 (N_2633,N_2551,N_2515);
or U2634 (N_2634,N_2558,N_2595);
and U2635 (N_2635,N_2554,N_2548);
and U2636 (N_2636,N_2526,N_2555);
nand U2637 (N_2637,N_2559,N_2528);
xnor U2638 (N_2638,N_2573,N_2531);
or U2639 (N_2639,N_2547,N_2500);
or U2640 (N_2640,N_2541,N_2599);
nand U2641 (N_2641,N_2511,N_2525);
nor U2642 (N_2642,N_2557,N_2582);
or U2643 (N_2643,N_2519,N_2521);
xor U2644 (N_2644,N_2502,N_2508);
nand U2645 (N_2645,N_2512,N_2517);
or U2646 (N_2646,N_2529,N_2584);
nor U2647 (N_2647,N_2578,N_2509);
and U2648 (N_2648,N_2563,N_2550);
and U2649 (N_2649,N_2505,N_2513);
nor U2650 (N_2650,N_2544,N_2564);
or U2651 (N_2651,N_2502,N_2533);
nand U2652 (N_2652,N_2595,N_2512);
and U2653 (N_2653,N_2588,N_2590);
or U2654 (N_2654,N_2570,N_2595);
or U2655 (N_2655,N_2571,N_2585);
nand U2656 (N_2656,N_2539,N_2514);
or U2657 (N_2657,N_2593,N_2509);
nor U2658 (N_2658,N_2507,N_2524);
nand U2659 (N_2659,N_2558,N_2575);
nor U2660 (N_2660,N_2522,N_2510);
nor U2661 (N_2661,N_2548,N_2599);
or U2662 (N_2662,N_2524,N_2509);
nor U2663 (N_2663,N_2545,N_2544);
and U2664 (N_2664,N_2555,N_2501);
nand U2665 (N_2665,N_2530,N_2562);
nor U2666 (N_2666,N_2522,N_2507);
or U2667 (N_2667,N_2508,N_2559);
or U2668 (N_2668,N_2569,N_2524);
nand U2669 (N_2669,N_2565,N_2545);
nor U2670 (N_2670,N_2535,N_2580);
or U2671 (N_2671,N_2568,N_2573);
and U2672 (N_2672,N_2585,N_2504);
or U2673 (N_2673,N_2597,N_2596);
and U2674 (N_2674,N_2583,N_2523);
and U2675 (N_2675,N_2504,N_2580);
and U2676 (N_2676,N_2561,N_2501);
and U2677 (N_2677,N_2593,N_2566);
nand U2678 (N_2678,N_2597,N_2553);
nor U2679 (N_2679,N_2502,N_2540);
nand U2680 (N_2680,N_2583,N_2519);
or U2681 (N_2681,N_2519,N_2580);
and U2682 (N_2682,N_2583,N_2588);
nand U2683 (N_2683,N_2537,N_2572);
or U2684 (N_2684,N_2563,N_2544);
nand U2685 (N_2685,N_2575,N_2537);
or U2686 (N_2686,N_2540,N_2576);
or U2687 (N_2687,N_2580,N_2569);
or U2688 (N_2688,N_2514,N_2596);
xor U2689 (N_2689,N_2500,N_2593);
nor U2690 (N_2690,N_2542,N_2593);
nand U2691 (N_2691,N_2570,N_2540);
nor U2692 (N_2692,N_2529,N_2508);
nand U2693 (N_2693,N_2584,N_2575);
and U2694 (N_2694,N_2553,N_2512);
nand U2695 (N_2695,N_2566,N_2562);
or U2696 (N_2696,N_2522,N_2552);
or U2697 (N_2697,N_2569,N_2585);
nor U2698 (N_2698,N_2595,N_2543);
nor U2699 (N_2699,N_2592,N_2569);
or U2700 (N_2700,N_2635,N_2691);
nor U2701 (N_2701,N_2690,N_2666);
or U2702 (N_2702,N_2641,N_2643);
and U2703 (N_2703,N_2625,N_2695);
xor U2704 (N_2704,N_2648,N_2610);
and U2705 (N_2705,N_2607,N_2629);
nand U2706 (N_2706,N_2684,N_2636);
or U2707 (N_2707,N_2676,N_2670);
nor U2708 (N_2708,N_2667,N_2689);
and U2709 (N_2709,N_2611,N_2606);
and U2710 (N_2710,N_2668,N_2645);
or U2711 (N_2711,N_2683,N_2680);
nor U2712 (N_2712,N_2608,N_2661);
nor U2713 (N_2713,N_2679,N_2632);
nor U2714 (N_2714,N_2658,N_2687);
nor U2715 (N_2715,N_2631,N_2603);
nand U2716 (N_2716,N_2615,N_2622);
nand U2717 (N_2717,N_2672,N_2677);
and U2718 (N_2718,N_2673,N_2637);
or U2719 (N_2719,N_2646,N_2671);
nand U2720 (N_2720,N_2662,N_2627);
nand U2721 (N_2721,N_2685,N_2656);
and U2722 (N_2722,N_2634,N_2697);
nand U2723 (N_2723,N_2618,N_2654);
or U2724 (N_2724,N_2604,N_2678);
and U2725 (N_2725,N_2620,N_2686);
or U2726 (N_2726,N_2617,N_2630);
xor U2727 (N_2727,N_2605,N_2663);
or U2728 (N_2728,N_2642,N_2601);
nand U2729 (N_2729,N_2614,N_2675);
nor U2730 (N_2730,N_2612,N_2692);
nand U2731 (N_2731,N_2609,N_2621);
or U2732 (N_2732,N_2633,N_2665);
nor U2733 (N_2733,N_2651,N_2600);
nor U2734 (N_2734,N_2694,N_2652);
and U2735 (N_2735,N_2623,N_2688);
or U2736 (N_2736,N_2681,N_2639);
or U2737 (N_2737,N_2619,N_2638);
nand U2738 (N_2738,N_2653,N_2649);
and U2739 (N_2739,N_2650,N_2669);
or U2740 (N_2740,N_2613,N_2602);
nand U2741 (N_2741,N_2657,N_2682);
nand U2742 (N_2742,N_2616,N_2674);
and U2743 (N_2743,N_2696,N_2659);
nand U2744 (N_2744,N_2660,N_2693);
nor U2745 (N_2745,N_2626,N_2655);
nand U2746 (N_2746,N_2664,N_2640);
and U2747 (N_2747,N_2624,N_2628);
nor U2748 (N_2748,N_2698,N_2647);
and U2749 (N_2749,N_2699,N_2644);
nand U2750 (N_2750,N_2617,N_2679);
nand U2751 (N_2751,N_2605,N_2698);
xnor U2752 (N_2752,N_2666,N_2685);
and U2753 (N_2753,N_2655,N_2696);
or U2754 (N_2754,N_2606,N_2672);
and U2755 (N_2755,N_2677,N_2639);
or U2756 (N_2756,N_2685,N_2609);
nand U2757 (N_2757,N_2631,N_2676);
or U2758 (N_2758,N_2603,N_2644);
and U2759 (N_2759,N_2601,N_2668);
nand U2760 (N_2760,N_2662,N_2675);
and U2761 (N_2761,N_2609,N_2633);
nor U2762 (N_2762,N_2623,N_2671);
nor U2763 (N_2763,N_2601,N_2684);
nor U2764 (N_2764,N_2649,N_2682);
nor U2765 (N_2765,N_2601,N_2675);
and U2766 (N_2766,N_2650,N_2657);
nand U2767 (N_2767,N_2667,N_2696);
nor U2768 (N_2768,N_2604,N_2676);
and U2769 (N_2769,N_2671,N_2691);
and U2770 (N_2770,N_2689,N_2692);
and U2771 (N_2771,N_2692,N_2699);
or U2772 (N_2772,N_2660,N_2676);
and U2773 (N_2773,N_2629,N_2675);
and U2774 (N_2774,N_2611,N_2654);
or U2775 (N_2775,N_2653,N_2622);
or U2776 (N_2776,N_2674,N_2692);
and U2777 (N_2777,N_2618,N_2607);
nand U2778 (N_2778,N_2698,N_2665);
nand U2779 (N_2779,N_2694,N_2612);
nor U2780 (N_2780,N_2698,N_2689);
and U2781 (N_2781,N_2670,N_2611);
nand U2782 (N_2782,N_2630,N_2611);
nor U2783 (N_2783,N_2658,N_2602);
nor U2784 (N_2784,N_2698,N_2640);
or U2785 (N_2785,N_2640,N_2692);
or U2786 (N_2786,N_2682,N_2671);
nand U2787 (N_2787,N_2695,N_2676);
nand U2788 (N_2788,N_2638,N_2627);
and U2789 (N_2789,N_2611,N_2691);
and U2790 (N_2790,N_2667,N_2623);
nand U2791 (N_2791,N_2642,N_2691);
nor U2792 (N_2792,N_2628,N_2642);
nand U2793 (N_2793,N_2647,N_2660);
nand U2794 (N_2794,N_2619,N_2656);
and U2795 (N_2795,N_2695,N_2656);
nor U2796 (N_2796,N_2654,N_2667);
nand U2797 (N_2797,N_2625,N_2620);
or U2798 (N_2798,N_2652,N_2645);
nand U2799 (N_2799,N_2694,N_2646);
nor U2800 (N_2800,N_2727,N_2791);
and U2801 (N_2801,N_2752,N_2759);
nor U2802 (N_2802,N_2733,N_2757);
nor U2803 (N_2803,N_2745,N_2735);
and U2804 (N_2804,N_2789,N_2772);
nand U2805 (N_2805,N_2762,N_2718);
nor U2806 (N_2806,N_2744,N_2771);
nand U2807 (N_2807,N_2750,N_2726);
nand U2808 (N_2808,N_2741,N_2793);
and U2809 (N_2809,N_2711,N_2729);
nor U2810 (N_2810,N_2763,N_2767);
or U2811 (N_2811,N_2743,N_2769);
nor U2812 (N_2812,N_2780,N_2760);
nor U2813 (N_2813,N_2749,N_2766);
and U2814 (N_2814,N_2728,N_2702);
nand U2815 (N_2815,N_2754,N_2705);
or U2816 (N_2816,N_2761,N_2747);
or U2817 (N_2817,N_2781,N_2778);
or U2818 (N_2818,N_2776,N_2725);
nand U2819 (N_2819,N_2724,N_2792);
nand U2820 (N_2820,N_2738,N_2786);
or U2821 (N_2821,N_2736,N_2706);
nor U2822 (N_2822,N_2770,N_2740);
nand U2823 (N_2823,N_2707,N_2756);
nor U2824 (N_2824,N_2730,N_2787);
nand U2825 (N_2825,N_2790,N_2746);
or U2826 (N_2826,N_2704,N_2737);
nor U2827 (N_2827,N_2775,N_2714);
nand U2828 (N_2828,N_2797,N_2713);
nor U2829 (N_2829,N_2715,N_2710);
nor U2830 (N_2830,N_2753,N_2734);
nor U2831 (N_2831,N_2773,N_2720);
nor U2832 (N_2832,N_2758,N_2732);
nor U2833 (N_2833,N_2722,N_2788);
and U2834 (N_2834,N_2751,N_2798);
and U2835 (N_2835,N_2703,N_2716);
and U2836 (N_2836,N_2777,N_2748);
and U2837 (N_2837,N_2721,N_2717);
or U2838 (N_2838,N_2700,N_2723);
nand U2839 (N_2839,N_2701,N_2719);
nand U2840 (N_2840,N_2742,N_2795);
nor U2841 (N_2841,N_2785,N_2709);
nand U2842 (N_2842,N_2782,N_2708);
nand U2843 (N_2843,N_2783,N_2765);
nor U2844 (N_2844,N_2794,N_2712);
or U2845 (N_2845,N_2731,N_2739);
and U2846 (N_2846,N_2755,N_2779);
nor U2847 (N_2847,N_2768,N_2774);
and U2848 (N_2848,N_2764,N_2796);
nor U2849 (N_2849,N_2799,N_2784);
and U2850 (N_2850,N_2788,N_2733);
nor U2851 (N_2851,N_2762,N_2765);
nand U2852 (N_2852,N_2787,N_2709);
nor U2853 (N_2853,N_2727,N_2788);
and U2854 (N_2854,N_2787,N_2762);
nand U2855 (N_2855,N_2735,N_2786);
nand U2856 (N_2856,N_2783,N_2731);
or U2857 (N_2857,N_2755,N_2701);
or U2858 (N_2858,N_2726,N_2724);
or U2859 (N_2859,N_2717,N_2794);
and U2860 (N_2860,N_2790,N_2714);
xnor U2861 (N_2861,N_2751,N_2720);
and U2862 (N_2862,N_2740,N_2760);
and U2863 (N_2863,N_2750,N_2747);
nor U2864 (N_2864,N_2719,N_2772);
nor U2865 (N_2865,N_2743,N_2773);
nor U2866 (N_2866,N_2760,N_2738);
and U2867 (N_2867,N_2725,N_2759);
nor U2868 (N_2868,N_2789,N_2729);
nor U2869 (N_2869,N_2713,N_2703);
nand U2870 (N_2870,N_2726,N_2754);
nor U2871 (N_2871,N_2794,N_2778);
or U2872 (N_2872,N_2702,N_2705);
nand U2873 (N_2873,N_2734,N_2785);
nand U2874 (N_2874,N_2776,N_2716);
and U2875 (N_2875,N_2765,N_2714);
and U2876 (N_2876,N_2719,N_2722);
nor U2877 (N_2877,N_2701,N_2764);
and U2878 (N_2878,N_2722,N_2795);
nor U2879 (N_2879,N_2773,N_2726);
and U2880 (N_2880,N_2712,N_2732);
or U2881 (N_2881,N_2779,N_2780);
nor U2882 (N_2882,N_2766,N_2797);
nand U2883 (N_2883,N_2748,N_2701);
nor U2884 (N_2884,N_2756,N_2711);
nand U2885 (N_2885,N_2777,N_2766);
and U2886 (N_2886,N_2784,N_2781);
nand U2887 (N_2887,N_2740,N_2713);
nand U2888 (N_2888,N_2729,N_2762);
nor U2889 (N_2889,N_2738,N_2729);
nand U2890 (N_2890,N_2755,N_2784);
nor U2891 (N_2891,N_2772,N_2778);
and U2892 (N_2892,N_2770,N_2708);
nor U2893 (N_2893,N_2732,N_2766);
and U2894 (N_2894,N_2752,N_2718);
nor U2895 (N_2895,N_2746,N_2700);
or U2896 (N_2896,N_2700,N_2724);
or U2897 (N_2897,N_2766,N_2751);
nor U2898 (N_2898,N_2708,N_2791);
and U2899 (N_2899,N_2725,N_2750);
nor U2900 (N_2900,N_2812,N_2866);
xnor U2901 (N_2901,N_2872,N_2850);
nor U2902 (N_2902,N_2829,N_2894);
nand U2903 (N_2903,N_2825,N_2881);
and U2904 (N_2904,N_2867,N_2864);
nand U2905 (N_2905,N_2834,N_2880);
nand U2906 (N_2906,N_2816,N_2838);
nor U2907 (N_2907,N_2854,N_2831);
nand U2908 (N_2908,N_2828,N_2890);
or U2909 (N_2909,N_2817,N_2874);
nand U2910 (N_2910,N_2809,N_2892);
nand U2911 (N_2911,N_2860,N_2862);
and U2912 (N_2912,N_2876,N_2801);
and U2913 (N_2913,N_2858,N_2803);
or U2914 (N_2914,N_2835,N_2895);
nand U2915 (N_2915,N_2877,N_2885);
and U2916 (N_2916,N_2807,N_2865);
and U2917 (N_2917,N_2839,N_2861);
and U2918 (N_2918,N_2887,N_2806);
nand U2919 (N_2919,N_2802,N_2843);
nand U2920 (N_2920,N_2841,N_2842);
nor U2921 (N_2921,N_2820,N_2814);
nor U2922 (N_2922,N_2873,N_2823);
and U2923 (N_2923,N_2893,N_2852);
and U2924 (N_2924,N_2827,N_2847);
nor U2925 (N_2925,N_2889,N_2856);
nor U2926 (N_2926,N_2853,N_2824);
nand U2927 (N_2927,N_2818,N_2855);
and U2928 (N_2928,N_2898,N_2870);
nor U2929 (N_2929,N_2805,N_2896);
and U2930 (N_2930,N_2883,N_2819);
nand U2931 (N_2931,N_2800,N_2815);
nand U2932 (N_2932,N_2813,N_2884);
nand U2933 (N_2933,N_2888,N_2849);
nand U2934 (N_2934,N_2851,N_2836);
or U2935 (N_2935,N_2821,N_2830);
nor U2936 (N_2936,N_2857,N_2879);
nor U2937 (N_2937,N_2810,N_2899);
or U2938 (N_2938,N_2848,N_2808);
nor U2939 (N_2939,N_2844,N_2868);
nor U2940 (N_2940,N_2840,N_2826);
or U2941 (N_2941,N_2891,N_2897);
or U2942 (N_2942,N_2804,N_2822);
and U2943 (N_2943,N_2846,N_2859);
nor U2944 (N_2944,N_2832,N_2871);
and U2945 (N_2945,N_2886,N_2878);
nand U2946 (N_2946,N_2869,N_2837);
nand U2947 (N_2947,N_2882,N_2833);
or U2948 (N_2948,N_2811,N_2845);
nor U2949 (N_2949,N_2875,N_2863);
nor U2950 (N_2950,N_2822,N_2827);
nand U2951 (N_2951,N_2839,N_2857);
and U2952 (N_2952,N_2834,N_2827);
nor U2953 (N_2953,N_2808,N_2855);
nor U2954 (N_2954,N_2816,N_2872);
or U2955 (N_2955,N_2858,N_2812);
or U2956 (N_2956,N_2896,N_2883);
nand U2957 (N_2957,N_2859,N_2857);
and U2958 (N_2958,N_2876,N_2883);
or U2959 (N_2959,N_2825,N_2834);
nor U2960 (N_2960,N_2841,N_2809);
nor U2961 (N_2961,N_2891,N_2864);
or U2962 (N_2962,N_2868,N_2879);
nand U2963 (N_2963,N_2885,N_2881);
nand U2964 (N_2964,N_2892,N_2891);
or U2965 (N_2965,N_2881,N_2858);
nand U2966 (N_2966,N_2871,N_2875);
or U2967 (N_2967,N_2887,N_2892);
nand U2968 (N_2968,N_2840,N_2896);
and U2969 (N_2969,N_2804,N_2876);
nor U2970 (N_2970,N_2886,N_2842);
and U2971 (N_2971,N_2890,N_2863);
and U2972 (N_2972,N_2845,N_2850);
nand U2973 (N_2973,N_2850,N_2891);
or U2974 (N_2974,N_2865,N_2831);
nor U2975 (N_2975,N_2838,N_2871);
and U2976 (N_2976,N_2803,N_2814);
xor U2977 (N_2977,N_2803,N_2820);
and U2978 (N_2978,N_2888,N_2825);
and U2979 (N_2979,N_2856,N_2854);
nand U2980 (N_2980,N_2868,N_2805);
and U2981 (N_2981,N_2804,N_2853);
nand U2982 (N_2982,N_2892,N_2898);
nand U2983 (N_2983,N_2816,N_2802);
nand U2984 (N_2984,N_2887,N_2805);
and U2985 (N_2985,N_2821,N_2872);
or U2986 (N_2986,N_2804,N_2896);
nor U2987 (N_2987,N_2854,N_2893);
nor U2988 (N_2988,N_2829,N_2858);
nand U2989 (N_2989,N_2887,N_2847);
nor U2990 (N_2990,N_2872,N_2828);
or U2991 (N_2991,N_2886,N_2871);
nand U2992 (N_2992,N_2875,N_2891);
and U2993 (N_2993,N_2858,N_2893);
nor U2994 (N_2994,N_2820,N_2870);
and U2995 (N_2995,N_2825,N_2886);
nand U2996 (N_2996,N_2893,N_2813);
or U2997 (N_2997,N_2896,N_2861);
nor U2998 (N_2998,N_2858,N_2859);
and U2999 (N_2999,N_2889,N_2821);
and UO_0 (O_0,N_2951,N_2900);
nor UO_1 (O_1,N_2998,N_2996);
and UO_2 (O_2,N_2995,N_2907);
nor UO_3 (O_3,N_2931,N_2958);
or UO_4 (O_4,N_2902,N_2956);
nand UO_5 (O_5,N_2912,N_2975);
nand UO_6 (O_6,N_2985,N_2963);
nor UO_7 (O_7,N_2986,N_2945);
or UO_8 (O_8,N_2982,N_2949);
nor UO_9 (O_9,N_2977,N_2999);
xor UO_10 (O_10,N_2934,N_2962);
or UO_11 (O_11,N_2946,N_2959);
nor UO_12 (O_12,N_2965,N_2905);
and UO_13 (O_13,N_2925,N_2937);
nor UO_14 (O_14,N_2923,N_2917);
and UO_15 (O_15,N_2916,N_2929);
nand UO_16 (O_16,N_2981,N_2989);
nand UO_17 (O_17,N_2942,N_2992);
nor UO_18 (O_18,N_2974,N_2909);
and UO_19 (O_19,N_2990,N_2944);
nand UO_20 (O_20,N_2911,N_2940);
nor UO_21 (O_21,N_2997,N_2987);
nand UO_22 (O_22,N_2935,N_2906);
and UO_23 (O_23,N_2918,N_2914);
nor UO_24 (O_24,N_2976,N_2952);
nor UO_25 (O_25,N_2938,N_2943);
or UO_26 (O_26,N_2969,N_2983);
and UO_27 (O_27,N_2954,N_2927);
or UO_28 (O_28,N_2919,N_2941);
nand UO_29 (O_29,N_2968,N_2971);
nor UO_30 (O_30,N_2903,N_2953);
nor UO_31 (O_31,N_2950,N_2948);
and UO_32 (O_32,N_2994,N_2908);
nor UO_33 (O_33,N_2926,N_2901);
and UO_34 (O_34,N_2978,N_2924);
or UO_35 (O_35,N_2964,N_2955);
nand UO_36 (O_36,N_2960,N_2930);
nor UO_37 (O_37,N_2973,N_2993);
or UO_38 (O_38,N_2939,N_2991);
nor UO_39 (O_39,N_2967,N_2961);
nand UO_40 (O_40,N_2920,N_2979);
and UO_41 (O_41,N_2928,N_2922);
or UO_42 (O_42,N_2915,N_2932);
and UO_43 (O_43,N_2972,N_2910);
and UO_44 (O_44,N_2913,N_2947);
or UO_45 (O_45,N_2980,N_2966);
nand UO_46 (O_46,N_2904,N_2936);
nand UO_47 (O_47,N_2988,N_2970);
nor UO_48 (O_48,N_2921,N_2933);
nand UO_49 (O_49,N_2957,N_2984);
or UO_50 (O_50,N_2932,N_2993);
nor UO_51 (O_51,N_2987,N_2930);
nand UO_52 (O_52,N_2921,N_2910);
nand UO_53 (O_53,N_2921,N_2956);
and UO_54 (O_54,N_2922,N_2985);
nand UO_55 (O_55,N_2934,N_2911);
or UO_56 (O_56,N_2931,N_2904);
or UO_57 (O_57,N_2940,N_2936);
nor UO_58 (O_58,N_2983,N_2981);
and UO_59 (O_59,N_2937,N_2958);
nand UO_60 (O_60,N_2946,N_2968);
nor UO_61 (O_61,N_2977,N_2914);
or UO_62 (O_62,N_2953,N_2940);
nand UO_63 (O_63,N_2951,N_2991);
nand UO_64 (O_64,N_2942,N_2925);
or UO_65 (O_65,N_2993,N_2990);
nor UO_66 (O_66,N_2948,N_2935);
and UO_67 (O_67,N_2981,N_2932);
or UO_68 (O_68,N_2954,N_2941);
nor UO_69 (O_69,N_2904,N_2944);
xnor UO_70 (O_70,N_2974,N_2973);
nor UO_71 (O_71,N_2986,N_2971);
nand UO_72 (O_72,N_2972,N_2947);
and UO_73 (O_73,N_2997,N_2948);
or UO_74 (O_74,N_2914,N_2906);
and UO_75 (O_75,N_2945,N_2961);
nand UO_76 (O_76,N_2980,N_2997);
nand UO_77 (O_77,N_2920,N_2987);
nand UO_78 (O_78,N_2931,N_2906);
nor UO_79 (O_79,N_2901,N_2908);
and UO_80 (O_80,N_2979,N_2954);
nand UO_81 (O_81,N_2958,N_2947);
and UO_82 (O_82,N_2979,N_2978);
nand UO_83 (O_83,N_2997,N_2940);
nor UO_84 (O_84,N_2915,N_2910);
xnor UO_85 (O_85,N_2996,N_2909);
and UO_86 (O_86,N_2914,N_2958);
or UO_87 (O_87,N_2946,N_2994);
and UO_88 (O_88,N_2949,N_2983);
nor UO_89 (O_89,N_2944,N_2923);
nand UO_90 (O_90,N_2940,N_2909);
or UO_91 (O_91,N_2909,N_2999);
or UO_92 (O_92,N_2935,N_2929);
and UO_93 (O_93,N_2993,N_2915);
nand UO_94 (O_94,N_2932,N_2999);
or UO_95 (O_95,N_2944,N_2917);
or UO_96 (O_96,N_2935,N_2903);
or UO_97 (O_97,N_2913,N_2953);
nor UO_98 (O_98,N_2936,N_2983);
nor UO_99 (O_99,N_2977,N_2961);
or UO_100 (O_100,N_2912,N_2920);
or UO_101 (O_101,N_2989,N_2953);
and UO_102 (O_102,N_2940,N_2937);
nand UO_103 (O_103,N_2920,N_2957);
nor UO_104 (O_104,N_2964,N_2919);
nand UO_105 (O_105,N_2977,N_2929);
nor UO_106 (O_106,N_2940,N_2907);
nand UO_107 (O_107,N_2989,N_2903);
nand UO_108 (O_108,N_2966,N_2958);
or UO_109 (O_109,N_2931,N_2998);
or UO_110 (O_110,N_2930,N_2939);
nand UO_111 (O_111,N_2991,N_2901);
nand UO_112 (O_112,N_2932,N_2941);
nor UO_113 (O_113,N_2984,N_2911);
or UO_114 (O_114,N_2969,N_2947);
xor UO_115 (O_115,N_2937,N_2971);
nand UO_116 (O_116,N_2957,N_2963);
or UO_117 (O_117,N_2997,N_2958);
nand UO_118 (O_118,N_2965,N_2997);
nor UO_119 (O_119,N_2982,N_2996);
nor UO_120 (O_120,N_2907,N_2970);
nor UO_121 (O_121,N_2977,N_2967);
and UO_122 (O_122,N_2973,N_2966);
nor UO_123 (O_123,N_2986,N_2965);
and UO_124 (O_124,N_2914,N_2959);
and UO_125 (O_125,N_2913,N_2918);
nor UO_126 (O_126,N_2958,N_2999);
and UO_127 (O_127,N_2933,N_2922);
or UO_128 (O_128,N_2913,N_2940);
nor UO_129 (O_129,N_2975,N_2952);
and UO_130 (O_130,N_2921,N_2914);
and UO_131 (O_131,N_2921,N_2943);
and UO_132 (O_132,N_2923,N_2940);
nor UO_133 (O_133,N_2981,N_2904);
or UO_134 (O_134,N_2944,N_2992);
and UO_135 (O_135,N_2964,N_2912);
and UO_136 (O_136,N_2901,N_2997);
nor UO_137 (O_137,N_2978,N_2965);
nor UO_138 (O_138,N_2985,N_2931);
and UO_139 (O_139,N_2957,N_2933);
and UO_140 (O_140,N_2900,N_2904);
and UO_141 (O_141,N_2925,N_2922);
nor UO_142 (O_142,N_2993,N_2967);
nor UO_143 (O_143,N_2919,N_2979);
or UO_144 (O_144,N_2982,N_2925);
and UO_145 (O_145,N_2953,N_2981);
and UO_146 (O_146,N_2908,N_2937);
and UO_147 (O_147,N_2950,N_2994);
xnor UO_148 (O_148,N_2997,N_2985);
and UO_149 (O_149,N_2921,N_2992);
nor UO_150 (O_150,N_2996,N_2903);
and UO_151 (O_151,N_2917,N_2977);
and UO_152 (O_152,N_2937,N_2950);
or UO_153 (O_153,N_2981,N_2913);
nand UO_154 (O_154,N_2996,N_2973);
nor UO_155 (O_155,N_2968,N_2984);
or UO_156 (O_156,N_2919,N_2982);
nand UO_157 (O_157,N_2942,N_2956);
and UO_158 (O_158,N_2977,N_2904);
and UO_159 (O_159,N_2917,N_2973);
nand UO_160 (O_160,N_2998,N_2972);
or UO_161 (O_161,N_2984,N_2992);
and UO_162 (O_162,N_2910,N_2947);
nor UO_163 (O_163,N_2933,N_2915);
nand UO_164 (O_164,N_2920,N_2921);
nand UO_165 (O_165,N_2919,N_2970);
nand UO_166 (O_166,N_2969,N_2953);
and UO_167 (O_167,N_2908,N_2961);
and UO_168 (O_168,N_2922,N_2943);
nand UO_169 (O_169,N_2913,N_2988);
nand UO_170 (O_170,N_2980,N_2994);
and UO_171 (O_171,N_2969,N_2911);
nor UO_172 (O_172,N_2926,N_2903);
and UO_173 (O_173,N_2911,N_2925);
nor UO_174 (O_174,N_2971,N_2984);
and UO_175 (O_175,N_2945,N_2944);
and UO_176 (O_176,N_2936,N_2975);
nor UO_177 (O_177,N_2978,N_2997);
nand UO_178 (O_178,N_2902,N_2927);
nand UO_179 (O_179,N_2937,N_2989);
or UO_180 (O_180,N_2945,N_2953);
nand UO_181 (O_181,N_2922,N_2945);
nand UO_182 (O_182,N_2942,N_2939);
nor UO_183 (O_183,N_2922,N_2951);
nand UO_184 (O_184,N_2962,N_2944);
or UO_185 (O_185,N_2967,N_2930);
or UO_186 (O_186,N_2974,N_2954);
nor UO_187 (O_187,N_2976,N_2979);
nor UO_188 (O_188,N_2994,N_2939);
or UO_189 (O_189,N_2901,N_2995);
or UO_190 (O_190,N_2924,N_2906);
or UO_191 (O_191,N_2919,N_2969);
nor UO_192 (O_192,N_2966,N_2959);
and UO_193 (O_193,N_2990,N_2965);
nand UO_194 (O_194,N_2985,N_2968);
nand UO_195 (O_195,N_2998,N_2911);
nor UO_196 (O_196,N_2934,N_2998);
nand UO_197 (O_197,N_2994,N_2938);
nor UO_198 (O_198,N_2952,N_2961);
and UO_199 (O_199,N_2945,N_2959);
or UO_200 (O_200,N_2967,N_2969);
and UO_201 (O_201,N_2908,N_2911);
or UO_202 (O_202,N_2912,N_2936);
nor UO_203 (O_203,N_2984,N_2939);
nor UO_204 (O_204,N_2951,N_2987);
xor UO_205 (O_205,N_2984,N_2995);
nor UO_206 (O_206,N_2974,N_2975);
or UO_207 (O_207,N_2998,N_2949);
xnor UO_208 (O_208,N_2935,N_2997);
nor UO_209 (O_209,N_2920,N_2965);
and UO_210 (O_210,N_2998,N_2901);
nor UO_211 (O_211,N_2907,N_2945);
nor UO_212 (O_212,N_2993,N_2928);
and UO_213 (O_213,N_2945,N_2934);
or UO_214 (O_214,N_2923,N_2994);
and UO_215 (O_215,N_2935,N_2901);
nand UO_216 (O_216,N_2943,N_2906);
or UO_217 (O_217,N_2957,N_2914);
nor UO_218 (O_218,N_2907,N_2996);
or UO_219 (O_219,N_2996,N_2937);
and UO_220 (O_220,N_2924,N_2991);
and UO_221 (O_221,N_2970,N_2972);
nand UO_222 (O_222,N_2910,N_2991);
or UO_223 (O_223,N_2947,N_2930);
nand UO_224 (O_224,N_2983,N_2944);
nand UO_225 (O_225,N_2922,N_2900);
or UO_226 (O_226,N_2947,N_2923);
or UO_227 (O_227,N_2911,N_2932);
or UO_228 (O_228,N_2976,N_2912);
or UO_229 (O_229,N_2979,N_2999);
or UO_230 (O_230,N_2941,N_2998);
nor UO_231 (O_231,N_2910,N_2970);
nand UO_232 (O_232,N_2937,N_2965);
nor UO_233 (O_233,N_2947,N_2996);
nor UO_234 (O_234,N_2949,N_2913);
nand UO_235 (O_235,N_2940,N_2980);
and UO_236 (O_236,N_2960,N_2902);
or UO_237 (O_237,N_2994,N_2934);
or UO_238 (O_238,N_2959,N_2949);
nand UO_239 (O_239,N_2979,N_2957);
or UO_240 (O_240,N_2989,N_2973);
nand UO_241 (O_241,N_2953,N_2997);
nor UO_242 (O_242,N_2964,N_2985);
nand UO_243 (O_243,N_2949,N_2908);
or UO_244 (O_244,N_2978,N_2967);
xor UO_245 (O_245,N_2960,N_2982);
or UO_246 (O_246,N_2977,N_2987);
nand UO_247 (O_247,N_2960,N_2917);
nand UO_248 (O_248,N_2920,N_2991);
and UO_249 (O_249,N_2940,N_2916);
nand UO_250 (O_250,N_2972,N_2920);
nor UO_251 (O_251,N_2926,N_2904);
and UO_252 (O_252,N_2919,N_2954);
nor UO_253 (O_253,N_2990,N_2920);
nor UO_254 (O_254,N_2902,N_2918);
or UO_255 (O_255,N_2963,N_2911);
or UO_256 (O_256,N_2966,N_2994);
and UO_257 (O_257,N_2985,N_2935);
and UO_258 (O_258,N_2993,N_2930);
nand UO_259 (O_259,N_2927,N_2971);
or UO_260 (O_260,N_2917,N_2965);
nand UO_261 (O_261,N_2952,N_2989);
or UO_262 (O_262,N_2974,N_2922);
and UO_263 (O_263,N_2939,N_2986);
nand UO_264 (O_264,N_2949,N_2924);
and UO_265 (O_265,N_2975,N_2933);
and UO_266 (O_266,N_2933,N_2996);
nor UO_267 (O_267,N_2929,N_2944);
or UO_268 (O_268,N_2939,N_2979);
nor UO_269 (O_269,N_2913,N_2945);
nand UO_270 (O_270,N_2901,N_2969);
nand UO_271 (O_271,N_2958,N_2928);
or UO_272 (O_272,N_2936,N_2953);
nand UO_273 (O_273,N_2980,N_2983);
nor UO_274 (O_274,N_2979,N_2935);
nand UO_275 (O_275,N_2993,N_2984);
nand UO_276 (O_276,N_2902,N_2925);
nand UO_277 (O_277,N_2991,N_2999);
or UO_278 (O_278,N_2920,N_2914);
nor UO_279 (O_279,N_2999,N_2934);
nor UO_280 (O_280,N_2921,N_2988);
or UO_281 (O_281,N_2966,N_2960);
nor UO_282 (O_282,N_2911,N_2901);
or UO_283 (O_283,N_2917,N_2983);
nor UO_284 (O_284,N_2928,N_2906);
nor UO_285 (O_285,N_2946,N_2951);
nor UO_286 (O_286,N_2983,N_2931);
nor UO_287 (O_287,N_2955,N_2969);
xor UO_288 (O_288,N_2953,N_2925);
or UO_289 (O_289,N_2960,N_2918);
nand UO_290 (O_290,N_2909,N_2998);
nand UO_291 (O_291,N_2964,N_2910);
nor UO_292 (O_292,N_2955,N_2963);
nor UO_293 (O_293,N_2977,N_2918);
or UO_294 (O_294,N_2973,N_2988);
or UO_295 (O_295,N_2999,N_2906);
nand UO_296 (O_296,N_2984,N_2941);
nand UO_297 (O_297,N_2962,N_2997);
nor UO_298 (O_298,N_2958,N_2918);
nor UO_299 (O_299,N_2935,N_2975);
nor UO_300 (O_300,N_2933,N_2974);
and UO_301 (O_301,N_2902,N_2939);
nor UO_302 (O_302,N_2940,N_2983);
nor UO_303 (O_303,N_2929,N_2903);
nor UO_304 (O_304,N_2999,N_2937);
or UO_305 (O_305,N_2903,N_2968);
xnor UO_306 (O_306,N_2948,N_2953);
and UO_307 (O_307,N_2904,N_2935);
nand UO_308 (O_308,N_2937,N_2993);
or UO_309 (O_309,N_2997,N_2900);
nor UO_310 (O_310,N_2914,N_2936);
nor UO_311 (O_311,N_2980,N_2959);
nand UO_312 (O_312,N_2911,N_2961);
nor UO_313 (O_313,N_2984,N_2975);
and UO_314 (O_314,N_2995,N_2993);
nand UO_315 (O_315,N_2950,N_2975);
or UO_316 (O_316,N_2996,N_2993);
nand UO_317 (O_317,N_2903,N_2907);
nor UO_318 (O_318,N_2978,N_2994);
nand UO_319 (O_319,N_2914,N_2974);
or UO_320 (O_320,N_2937,N_2921);
nand UO_321 (O_321,N_2989,N_2922);
nand UO_322 (O_322,N_2973,N_2991);
or UO_323 (O_323,N_2912,N_2928);
and UO_324 (O_324,N_2923,N_2963);
nand UO_325 (O_325,N_2929,N_2939);
nand UO_326 (O_326,N_2930,N_2995);
and UO_327 (O_327,N_2931,N_2984);
and UO_328 (O_328,N_2920,N_2984);
nand UO_329 (O_329,N_2975,N_2997);
and UO_330 (O_330,N_2916,N_2991);
or UO_331 (O_331,N_2955,N_2936);
nor UO_332 (O_332,N_2955,N_2913);
nor UO_333 (O_333,N_2944,N_2911);
or UO_334 (O_334,N_2926,N_2999);
or UO_335 (O_335,N_2989,N_2980);
nand UO_336 (O_336,N_2945,N_2958);
nand UO_337 (O_337,N_2992,N_2983);
and UO_338 (O_338,N_2955,N_2979);
nor UO_339 (O_339,N_2947,N_2914);
nand UO_340 (O_340,N_2994,N_2991);
nand UO_341 (O_341,N_2926,N_2965);
or UO_342 (O_342,N_2979,N_2921);
nor UO_343 (O_343,N_2915,N_2976);
and UO_344 (O_344,N_2939,N_2989);
nand UO_345 (O_345,N_2934,N_2955);
or UO_346 (O_346,N_2934,N_2931);
nand UO_347 (O_347,N_2934,N_2949);
nor UO_348 (O_348,N_2947,N_2942);
or UO_349 (O_349,N_2936,N_2926);
or UO_350 (O_350,N_2957,N_2978);
and UO_351 (O_351,N_2981,N_2922);
nor UO_352 (O_352,N_2984,N_2961);
nor UO_353 (O_353,N_2944,N_2922);
or UO_354 (O_354,N_2906,N_2927);
nor UO_355 (O_355,N_2990,N_2960);
and UO_356 (O_356,N_2987,N_2935);
nor UO_357 (O_357,N_2926,N_2921);
nand UO_358 (O_358,N_2931,N_2970);
or UO_359 (O_359,N_2932,N_2929);
or UO_360 (O_360,N_2944,N_2943);
or UO_361 (O_361,N_2931,N_2930);
and UO_362 (O_362,N_2943,N_2965);
nor UO_363 (O_363,N_2973,N_2981);
nand UO_364 (O_364,N_2914,N_2905);
nand UO_365 (O_365,N_2924,N_2919);
nor UO_366 (O_366,N_2917,N_2912);
nand UO_367 (O_367,N_2983,N_2994);
or UO_368 (O_368,N_2996,N_2963);
and UO_369 (O_369,N_2955,N_2908);
nor UO_370 (O_370,N_2997,N_2929);
and UO_371 (O_371,N_2904,N_2932);
nor UO_372 (O_372,N_2931,N_2915);
or UO_373 (O_373,N_2962,N_2961);
nor UO_374 (O_374,N_2965,N_2960);
nand UO_375 (O_375,N_2942,N_2901);
nand UO_376 (O_376,N_2968,N_2987);
nor UO_377 (O_377,N_2991,N_2954);
xnor UO_378 (O_378,N_2995,N_2918);
and UO_379 (O_379,N_2905,N_2949);
or UO_380 (O_380,N_2935,N_2938);
nor UO_381 (O_381,N_2926,N_2930);
and UO_382 (O_382,N_2991,N_2932);
or UO_383 (O_383,N_2917,N_2954);
nand UO_384 (O_384,N_2912,N_2973);
or UO_385 (O_385,N_2969,N_2962);
nor UO_386 (O_386,N_2951,N_2954);
and UO_387 (O_387,N_2929,N_2967);
nor UO_388 (O_388,N_2901,N_2902);
nor UO_389 (O_389,N_2987,N_2975);
or UO_390 (O_390,N_2989,N_2993);
and UO_391 (O_391,N_2938,N_2922);
nor UO_392 (O_392,N_2978,N_2940);
nor UO_393 (O_393,N_2956,N_2976);
and UO_394 (O_394,N_2980,N_2948);
nand UO_395 (O_395,N_2915,N_2988);
nor UO_396 (O_396,N_2962,N_2957);
and UO_397 (O_397,N_2954,N_2968);
nand UO_398 (O_398,N_2910,N_2902);
and UO_399 (O_399,N_2967,N_2936);
and UO_400 (O_400,N_2925,N_2957);
and UO_401 (O_401,N_2987,N_2976);
and UO_402 (O_402,N_2946,N_2931);
and UO_403 (O_403,N_2991,N_2906);
and UO_404 (O_404,N_2914,N_2946);
nand UO_405 (O_405,N_2928,N_2931);
nand UO_406 (O_406,N_2990,N_2935);
nand UO_407 (O_407,N_2925,N_2901);
and UO_408 (O_408,N_2957,N_2990);
and UO_409 (O_409,N_2929,N_2911);
and UO_410 (O_410,N_2973,N_2983);
nor UO_411 (O_411,N_2915,N_2900);
or UO_412 (O_412,N_2901,N_2950);
nor UO_413 (O_413,N_2911,N_2907);
or UO_414 (O_414,N_2997,N_2950);
nor UO_415 (O_415,N_2945,N_2971);
nand UO_416 (O_416,N_2912,N_2965);
or UO_417 (O_417,N_2922,N_2906);
or UO_418 (O_418,N_2930,N_2922);
and UO_419 (O_419,N_2926,N_2945);
and UO_420 (O_420,N_2933,N_2958);
nand UO_421 (O_421,N_2955,N_2907);
nand UO_422 (O_422,N_2915,N_2979);
xnor UO_423 (O_423,N_2928,N_2955);
or UO_424 (O_424,N_2911,N_2983);
nand UO_425 (O_425,N_2925,N_2918);
and UO_426 (O_426,N_2999,N_2960);
nand UO_427 (O_427,N_2990,N_2961);
nor UO_428 (O_428,N_2926,N_2994);
and UO_429 (O_429,N_2981,N_2945);
nand UO_430 (O_430,N_2994,N_2972);
nand UO_431 (O_431,N_2990,N_2945);
and UO_432 (O_432,N_2908,N_2924);
nand UO_433 (O_433,N_2934,N_2981);
or UO_434 (O_434,N_2904,N_2959);
or UO_435 (O_435,N_2987,N_2999);
nor UO_436 (O_436,N_2954,N_2962);
nand UO_437 (O_437,N_2938,N_2945);
and UO_438 (O_438,N_2997,N_2920);
nor UO_439 (O_439,N_2945,N_2996);
nand UO_440 (O_440,N_2928,N_2905);
or UO_441 (O_441,N_2919,N_2944);
and UO_442 (O_442,N_2981,N_2966);
nor UO_443 (O_443,N_2905,N_2932);
or UO_444 (O_444,N_2950,N_2949);
and UO_445 (O_445,N_2999,N_2902);
or UO_446 (O_446,N_2908,N_2951);
nor UO_447 (O_447,N_2927,N_2936);
nand UO_448 (O_448,N_2984,N_2908);
nand UO_449 (O_449,N_2971,N_2959);
or UO_450 (O_450,N_2996,N_2983);
nor UO_451 (O_451,N_2915,N_2940);
nor UO_452 (O_452,N_2957,N_2940);
nand UO_453 (O_453,N_2973,N_2916);
nor UO_454 (O_454,N_2977,N_2965);
nor UO_455 (O_455,N_2952,N_2900);
nand UO_456 (O_456,N_2930,N_2951);
or UO_457 (O_457,N_2934,N_2990);
xor UO_458 (O_458,N_2966,N_2975);
and UO_459 (O_459,N_2933,N_2973);
and UO_460 (O_460,N_2966,N_2935);
or UO_461 (O_461,N_2912,N_2903);
and UO_462 (O_462,N_2919,N_2936);
and UO_463 (O_463,N_2931,N_2957);
and UO_464 (O_464,N_2977,N_2974);
nand UO_465 (O_465,N_2922,N_2986);
nand UO_466 (O_466,N_2932,N_2982);
nand UO_467 (O_467,N_2985,N_2952);
and UO_468 (O_468,N_2958,N_2968);
nor UO_469 (O_469,N_2927,N_2914);
or UO_470 (O_470,N_2982,N_2910);
and UO_471 (O_471,N_2968,N_2921);
and UO_472 (O_472,N_2974,N_2980);
xor UO_473 (O_473,N_2990,N_2908);
nand UO_474 (O_474,N_2906,N_2970);
or UO_475 (O_475,N_2925,N_2963);
nand UO_476 (O_476,N_2930,N_2980);
xor UO_477 (O_477,N_2976,N_2925);
nand UO_478 (O_478,N_2939,N_2938);
or UO_479 (O_479,N_2924,N_2927);
nor UO_480 (O_480,N_2909,N_2922);
and UO_481 (O_481,N_2934,N_2929);
or UO_482 (O_482,N_2926,N_2949);
nand UO_483 (O_483,N_2936,N_2979);
nand UO_484 (O_484,N_2996,N_2961);
and UO_485 (O_485,N_2955,N_2941);
or UO_486 (O_486,N_2982,N_2957);
nand UO_487 (O_487,N_2988,N_2920);
nand UO_488 (O_488,N_2965,N_2927);
nand UO_489 (O_489,N_2926,N_2950);
or UO_490 (O_490,N_2987,N_2927);
nor UO_491 (O_491,N_2937,N_2988);
nand UO_492 (O_492,N_2987,N_2949);
nand UO_493 (O_493,N_2920,N_2916);
or UO_494 (O_494,N_2988,N_2912);
or UO_495 (O_495,N_2906,N_2918);
and UO_496 (O_496,N_2954,N_2996);
or UO_497 (O_497,N_2933,N_2938);
and UO_498 (O_498,N_2926,N_2943);
nor UO_499 (O_499,N_2955,N_2945);
endmodule