module basic_1500_15000_2000_15_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_815,In_614);
or U1 (N_1,In_339,In_707);
and U2 (N_2,In_493,In_397);
or U3 (N_3,In_1457,In_681);
nand U4 (N_4,In_1211,In_340);
or U5 (N_5,In_218,In_41);
nor U6 (N_6,In_302,In_1112);
xor U7 (N_7,In_1417,In_1159);
nor U8 (N_8,In_229,In_828);
or U9 (N_9,In_305,In_1143);
nand U10 (N_10,In_425,In_474);
nor U11 (N_11,In_1221,In_285);
nand U12 (N_12,In_889,In_416);
or U13 (N_13,In_668,In_1069);
nand U14 (N_14,In_1066,In_1032);
and U15 (N_15,In_1123,In_867);
nand U16 (N_16,In_312,In_823);
nand U17 (N_17,In_851,In_619);
or U18 (N_18,In_445,In_814);
nor U19 (N_19,In_993,In_1480);
and U20 (N_20,In_361,In_1477);
nor U21 (N_21,In_1286,In_783);
xor U22 (N_22,In_1384,In_1149);
nand U23 (N_23,In_1333,In_478);
nor U24 (N_24,In_1138,In_646);
nand U25 (N_25,In_740,In_1453);
nor U26 (N_26,In_831,In_852);
nor U27 (N_27,In_435,In_468);
nand U28 (N_28,In_654,In_1022);
nor U29 (N_29,In_1188,In_1014);
and U30 (N_30,In_1376,In_1442);
nand U31 (N_31,In_1420,In_535);
nor U32 (N_32,In_824,In_1358);
or U33 (N_33,In_669,In_1258);
or U34 (N_34,In_221,In_438);
nor U35 (N_35,In_684,In_934);
nand U36 (N_36,In_816,In_219);
nor U37 (N_37,In_933,In_1409);
or U38 (N_38,In_286,In_723);
and U39 (N_39,In_835,In_1312);
nor U40 (N_40,In_807,In_631);
nand U41 (N_41,In_1083,In_829);
nand U42 (N_42,In_539,In_1397);
or U43 (N_43,In_1257,In_247);
and U44 (N_44,In_738,In_848);
nor U45 (N_45,In_1184,In_201);
or U46 (N_46,In_57,In_1445);
nand U47 (N_47,In_153,In_1183);
nor U48 (N_48,In_1297,In_1178);
or U49 (N_49,In_885,In_1317);
nand U50 (N_50,In_357,In_1227);
and U51 (N_51,In_273,In_21);
nor U52 (N_52,In_1475,In_1266);
xor U53 (N_53,In_639,In_659);
or U54 (N_54,In_1130,In_709);
or U55 (N_55,In_336,In_134);
or U56 (N_56,In_1119,In_941);
or U57 (N_57,In_653,In_618);
and U58 (N_58,In_315,In_132);
xor U59 (N_59,In_891,In_935);
or U60 (N_60,In_382,In_109);
and U61 (N_61,In_513,In_560);
nor U62 (N_62,In_197,In_91);
and U63 (N_63,In_1137,In_75);
nor U64 (N_64,In_368,In_1351);
and U65 (N_65,In_702,In_259);
or U66 (N_66,In_245,In_180);
nor U67 (N_67,In_1401,In_1155);
nand U68 (N_68,In_78,In_144);
xor U69 (N_69,In_367,In_264);
and U70 (N_70,In_1412,In_101);
and U71 (N_71,In_862,In_688);
nor U72 (N_72,In_1443,In_342);
nor U73 (N_73,In_248,In_353);
nand U74 (N_74,In_1287,In_534);
or U75 (N_75,In_411,In_591);
or U76 (N_76,In_656,In_1365);
and U77 (N_77,In_817,In_274);
and U78 (N_78,In_0,In_770);
nand U79 (N_79,In_626,In_1111);
nor U80 (N_80,In_296,In_1470);
nor U81 (N_81,In_1395,In_211);
nor U82 (N_82,In_613,In_1060);
xnor U83 (N_83,In_1386,In_925);
and U84 (N_84,In_426,In_721);
nor U85 (N_85,In_433,In_1424);
nand U86 (N_86,In_304,In_175);
nand U87 (N_87,In_524,In_152);
nor U88 (N_88,In_223,In_1447);
nor U89 (N_89,In_676,In_1306);
or U90 (N_90,In_1251,In_773);
nor U91 (N_91,In_1262,In_948);
nor U92 (N_92,In_151,In_1175);
and U93 (N_93,In_896,In_333);
and U94 (N_94,In_769,In_252);
xnor U95 (N_95,In_1415,In_737);
xnor U96 (N_96,In_784,In_951);
and U97 (N_97,In_365,In_750);
nand U98 (N_98,In_508,In_563);
or U99 (N_99,In_25,In_1281);
or U100 (N_100,In_103,In_1205);
nor U101 (N_101,In_892,In_297);
and U102 (N_102,In_1013,In_359);
nand U103 (N_103,In_1139,In_1483);
nand U104 (N_104,In_202,In_1244);
nand U105 (N_105,In_39,In_94);
xnor U106 (N_106,In_1464,In_1146);
or U107 (N_107,In_225,In_520);
or U108 (N_108,In_371,In_905);
nor U109 (N_109,In_1154,In_160);
and U110 (N_110,In_1356,In_808);
nand U111 (N_111,In_840,In_548);
nor U112 (N_112,In_240,In_827);
nor U113 (N_113,In_1168,In_545);
or U114 (N_114,In_422,In_847);
nand U115 (N_115,In_1054,In_251);
nand U116 (N_116,In_332,In_11);
and U117 (N_117,In_70,In_1327);
nor U118 (N_118,In_429,In_1302);
or U119 (N_119,In_1355,In_1132);
or U120 (N_120,In_624,In_980);
nand U121 (N_121,In_1448,In_1209);
nor U122 (N_122,In_1191,In_962);
nand U123 (N_123,In_1202,In_1434);
or U124 (N_124,In_992,In_1097);
and U125 (N_125,In_1190,In_573);
or U126 (N_126,In_237,In_698);
nand U127 (N_127,In_826,In_1031);
and U128 (N_128,In_494,In_1224);
nand U129 (N_129,In_1016,In_1003);
or U130 (N_130,In_177,In_1337);
xor U131 (N_131,In_466,In_1291);
or U132 (N_132,In_1182,In_1163);
nor U133 (N_133,In_1379,In_1493);
and U134 (N_134,In_1238,In_913);
or U135 (N_135,In_562,In_1289);
nand U136 (N_136,In_483,In_984);
nor U137 (N_137,In_1240,In_334);
nor U138 (N_138,In_637,In_489);
nand U139 (N_139,In_526,In_685);
and U140 (N_140,In_1400,In_1360);
xnor U141 (N_141,In_756,In_1428);
xor U142 (N_142,In_125,In_766);
xnor U143 (N_143,In_155,In_116);
nor U144 (N_144,In_1394,In_704);
and U145 (N_145,In_1098,In_401);
nor U146 (N_146,In_1167,In_35);
or U147 (N_147,In_779,In_1418);
nand U148 (N_148,In_89,In_323);
nand U149 (N_149,In_945,In_481);
or U150 (N_150,In_1374,In_348);
nor U151 (N_151,In_419,In_1487);
nor U152 (N_152,In_1080,In_909);
or U153 (N_153,In_1044,In_644);
nor U154 (N_154,In_162,In_987);
nand U155 (N_155,In_20,In_1288);
or U156 (N_156,In_1279,In_1268);
nor U157 (N_157,In_679,In_1348);
and U158 (N_158,In_127,In_1164);
or U159 (N_159,In_1450,In_574);
and U160 (N_160,In_71,In_1491);
and U161 (N_161,In_174,In_551);
and U162 (N_162,In_597,In_841);
or U163 (N_163,In_795,In_215);
nor U164 (N_164,In_739,In_448);
and U165 (N_165,In_161,In_275);
nor U166 (N_166,In_781,In_128);
and U167 (N_167,In_897,In_436);
or U168 (N_168,In_585,In_1335);
nor U169 (N_169,In_308,In_1070);
nor U170 (N_170,In_1040,In_431);
and U171 (N_171,In_977,In_236);
and U172 (N_172,In_1092,In_204);
xnor U173 (N_173,In_726,In_1116);
nor U174 (N_174,In_576,In_188);
and U175 (N_175,In_1438,In_895);
nor U176 (N_176,In_1332,In_281);
xnor U177 (N_177,In_1263,In_65);
nand U178 (N_178,In_1380,In_1313);
or U179 (N_179,In_1090,In_380);
nand U180 (N_180,In_486,In_966);
or U181 (N_181,In_212,In_752);
or U182 (N_182,In_724,In_875);
and U183 (N_183,In_250,In_1241);
and U184 (N_184,In_327,In_374);
nand U185 (N_185,In_34,In_865);
xnor U186 (N_186,In_146,In_156);
nor U187 (N_187,In_772,In_460);
nand U188 (N_188,In_1458,In_179);
and U189 (N_189,In_1037,In_1057);
nor U190 (N_190,In_882,In_695);
nor U191 (N_191,In_864,In_697);
xor U192 (N_192,In_51,In_12);
or U193 (N_193,In_1490,In_923);
xnor U194 (N_194,In_1282,In_810);
xor U195 (N_195,In_423,In_1398);
nand U196 (N_196,In_44,In_1153);
and U197 (N_197,In_131,In_1285);
and U198 (N_198,In_1315,In_1436);
nand U199 (N_199,In_475,In_1405);
nor U200 (N_200,In_1466,In_56);
and U201 (N_201,In_813,In_1077);
and U202 (N_202,In_1005,In_803);
nor U203 (N_203,In_981,In_791);
nor U204 (N_204,In_860,In_662);
and U205 (N_205,In_825,In_949);
xnor U206 (N_206,In_1231,In_410);
and U207 (N_207,In_461,In_1304);
nor U208 (N_208,In_1185,In_767);
or U209 (N_209,In_1200,In_506);
or U210 (N_210,In_257,In_846);
and U211 (N_211,In_115,In_344);
nand U212 (N_212,In_1203,In_249);
or U213 (N_213,In_1310,In_288);
or U214 (N_214,In_1048,In_836);
or U215 (N_215,In_625,In_964);
xnor U216 (N_216,In_1102,In_720);
or U217 (N_217,In_893,In_324);
and U218 (N_218,In_372,In_1296);
nand U219 (N_219,In_652,In_501);
nand U220 (N_220,In_108,In_496);
nor U221 (N_221,In_96,In_1273);
nand U222 (N_222,In_942,In_412);
and U223 (N_223,In_914,In_552);
nand U224 (N_224,In_1246,In_1017);
or U225 (N_225,In_504,In_46);
nor U226 (N_226,In_728,In_183);
nand U227 (N_227,In_122,In_787);
and U228 (N_228,In_121,In_965);
nand U229 (N_229,In_459,In_606);
or U230 (N_230,In_953,In_1148);
and U231 (N_231,In_1468,In_612);
nand U232 (N_232,In_1125,In_1218);
nor U233 (N_233,In_1195,In_337);
and U234 (N_234,In_629,In_1391);
xnor U235 (N_235,In_74,In_651);
nand U236 (N_236,In_66,In_581);
nor U237 (N_237,In_1027,In_1382);
and U238 (N_238,In_178,In_976);
nor U239 (N_239,In_734,In_565);
or U240 (N_240,In_262,In_838);
xor U241 (N_241,In_266,In_870);
or U242 (N_242,In_1423,In_119);
nand U243 (N_243,In_241,In_1301);
nor U244 (N_244,In_1187,In_1024);
or U245 (N_245,In_1068,In_1318);
xnor U246 (N_246,In_1026,In_1215);
or U247 (N_247,In_1117,In_561);
nand U248 (N_248,In_97,In_671);
nand U249 (N_249,In_370,In_1330);
or U250 (N_250,In_1147,In_716);
nand U251 (N_251,In_157,In_1481);
and U252 (N_252,In_804,In_64);
or U253 (N_253,In_499,In_620);
nor U254 (N_254,In_1440,In_531);
or U255 (N_255,In_924,In_341);
or U256 (N_256,In_871,In_173);
or U257 (N_257,In_647,In_997);
nand U258 (N_258,In_443,In_1316);
nand U259 (N_259,In_670,In_441);
or U260 (N_260,In_572,In_900);
and U261 (N_261,In_1081,In_18);
or U262 (N_262,In_1088,In_1454);
or U263 (N_263,In_1019,In_420);
nor U264 (N_264,In_1496,In_839);
nand U265 (N_265,In_802,In_158);
and U266 (N_266,In_446,In_170);
or U267 (N_267,In_788,In_49);
and U268 (N_268,In_917,In_150);
or U269 (N_269,In_261,In_373);
or U270 (N_270,In_604,In_636);
or U271 (N_271,In_605,In_1103);
nor U272 (N_272,In_1298,In_1091);
nand U273 (N_273,In_32,In_1414);
or U274 (N_274,In_1213,In_564);
and U275 (N_275,In_450,In_138);
or U276 (N_276,In_616,In_495);
nor U277 (N_277,In_1311,In_269);
nor U278 (N_278,In_1219,In_1115);
nor U279 (N_279,In_1011,In_746);
nor U280 (N_280,In_1074,In_1290);
or U281 (N_281,In_1237,In_471);
xor U282 (N_282,In_1035,In_1180);
or U283 (N_283,In_37,In_90);
and U284 (N_284,In_350,In_1383);
xor U285 (N_285,In_1134,In_1413);
nor U286 (N_286,In_389,In_352);
or U287 (N_287,In_5,In_1193);
nor U288 (N_288,In_806,In_511);
and U289 (N_289,In_329,In_351);
or U290 (N_290,In_1425,In_797);
and U291 (N_291,In_1267,In_1194);
nor U292 (N_292,In_1441,In_23);
xor U293 (N_293,In_936,In_529);
or U294 (N_294,In_849,In_298);
and U295 (N_295,In_1126,In_316);
xor U296 (N_296,In_9,In_47);
and U297 (N_297,In_745,In_226);
and U298 (N_298,In_710,In_477);
xnor U299 (N_299,In_1176,In_1431);
nor U300 (N_300,In_335,In_171);
nand U301 (N_301,In_322,In_550);
or U302 (N_302,In_915,In_113);
nor U303 (N_303,In_955,In_785);
and U304 (N_304,In_887,In_768);
nand U305 (N_305,In_714,In_593);
or U306 (N_306,In_1484,In_1094);
and U307 (N_307,In_880,In_658);
nand U308 (N_308,In_575,In_479);
xnor U309 (N_309,In_195,In_538);
and U310 (N_310,In_1086,In_107);
xnor U311 (N_311,In_983,In_1377);
nand U312 (N_312,In_40,In_1328);
nor U313 (N_313,In_759,In_314);
and U314 (N_314,In_580,In_117);
nand U315 (N_315,In_922,In_1270);
nand U316 (N_316,In_908,In_990);
nand U317 (N_317,In_973,In_154);
nor U318 (N_318,In_655,In_1127);
nor U319 (N_319,In_363,In_786);
nand U320 (N_320,In_272,In_693);
nand U321 (N_321,In_1122,In_400);
xnor U322 (N_322,In_1172,In_907);
nor U323 (N_323,In_124,In_208);
nor U324 (N_324,In_1249,In_845);
nand U325 (N_325,In_1364,In_776);
xnor U326 (N_326,In_543,In_856);
or U327 (N_327,In_366,In_1252);
nor U328 (N_328,In_1082,In_1233);
and U329 (N_329,In_837,In_541);
nor U330 (N_330,In_338,In_1004);
nand U331 (N_331,In_80,In_449);
and U332 (N_332,In_99,In_633);
or U333 (N_333,In_279,In_735);
nand U334 (N_334,In_17,In_635);
nand U335 (N_335,In_1388,In_729);
and U336 (N_336,In_1245,In_457);
nand U337 (N_337,In_509,In_1140);
nand U338 (N_338,In_528,In_1248);
nand U339 (N_339,In_883,In_570);
or U340 (N_340,In_969,In_510);
nor U341 (N_341,In_790,In_617);
nor U342 (N_342,In_55,In_863);
and U343 (N_343,In_800,In_694);
and U344 (N_344,In_1214,In_940);
or U345 (N_345,In_1259,In_1095);
nor U346 (N_346,In_569,In_1078);
nand U347 (N_347,In_1427,In_518);
xnor U348 (N_348,In_660,In_1023);
and U349 (N_349,In_163,In_1229);
xor U350 (N_350,In_855,In_730);
and U351 (N_351,In_77,In_164);
xnor U352 (N_352,In_715,In_1444);
or U353 (N_353,In_456,In_1407);
xor U354 (N_354,In_1071,In_703);
nor U355 (N_355,In_1096,In_1001);
or U356 (N_356,In_749,In_638);
xor U357 (N_357,In_1157,In_417);
and U358 (N_358,In_199,In_1265);
nand U359 (N_359,In_85,In_198);
nand U360 (N_360,In_1170,In_282);
nand U361 (N_361,In_1120,In_1150);
nand U362 (N_362,In_399,In_396);
and U363 (N_363,In_86,In_857);
or U364 (N_364,In_1275,In_243);
or U365 (N_365,In_26,In_1207);
or U366 (N_366,In_52,In_943);
or U367 (N_367,In_1135,In_1456);
nand U368 (N_368,In_683,In_191);
and U369 (N_369,In_927,In_611);
or U370 (N_370,In_379,In_1223);
nor U371 (N_371,In_63,In_514);
nand U372 (N_372,In_1276,In_1124);
nand U373 (N_373,In_415,In_1101);
and U374 (N_374,In_203,In_485);
nand U375 (N_375,In_1410,In_982);
or U376 (N_376,In_437,In_888);
nor U377 (N_377,In_1321,In_289);
nand U378 (N_378,In_622,In_490);
or U379 (N_379,In_931,In_588);
nor U380 (N_380,In_1010,In_301);
or U381 (N_381,In_995,In_453);
nor U382 (N_382,In_24,In_884);
nand U383 (N_383,In_1058,In_794);
and U384 (N_384,In_1152,In_780);
nand U385 (N_385,In_1280,In_196);
nand U386 (N_386,In_452,In_2);
nor U387 (N_387,In_525,In_821);
or U388 (N_388,In_858,In_1253);
or U389 (N_389,In_1220,In_553);
and U390 (N_390,In_1160,In_1106);
or U391 (N_391,In_1354,In_761);
xor U392 (N_392,In_187,In_1344);
nor U393 (N_393,In_873,In_182);
xor U394 (N_394,In_165,In_516);
nand U395 (N_395,In_29,In_392);
or U396 (N_396,In_126,In_623);
or U397 (N_397,In_13,In_1369);
or U398 (N_398,In_645,In_1136);
nand U399 (N_399,In_1000,In_978);
nand U400 (N_400,In_1338,In_1085);
or U401 (N_401,In_385,In_105);
and U402 (N_402,In_328,In_610);
nand U403 (N_403,In_1465,In_1271);
and U404 (N_404,In_280,In_1034);
or U405 (N_405,In_809,In_267);
nor U406 (N_406,In_691,In_38);
or U407 (N_407,In_300,In_1210);
nor U408 (N_408,In_258,In_1021);
nand U409 (N_409,In_53,In_246);
or U410 (N_410,In_507,In_1197);
and U411 (N_411,In_1411,In_112);
nor U412 (N_412,In_775,In_375);
xor U413 (N_413,In_994,In_1208);
nor U414 (N_414,In_1368,In_1072);
xnor U415 (N_415,In_1,In_255);
xor U416 (N_416,In_764,In_985);
xnor U417 (N_417,In_6,In_1269);
nand U418 (N_418,In_1459,In_584);
nor U419 (N_419,In_699,In_515);
nand U420 (N_420,In_522,In_952);
xnor U421 (N_421,In_220,In_307);
nand U422 (N_422,In_207,In_868);
or U423 (N_423,In_1173,In_320);
nand U424 (N_424,In_1067,In_1056);
nor U425 (N_425,In_1437,In_1087);
or U426 (N_426,In_100,In_254);
xnor U427 (N_427,In_185,In_1389);
nor U428 (N_428,In_583,In_242);
xor U429 (N_429,In_901,In_505);
nand U430 (N_430,In_22,In_799);
and U431 (N_431,In_1256,In_230);
or U432 (N_432,In_231,In_1341);
or U433 (N_433,In_330,In_384);
and U434 (N_434,In_1378,In_388);
nor U435 (N_435,In_1357,In_760);
nand U436 (N_436,In_599,In_488);
or U437 (N_437,In_722,In_1006);
nor U438 (N_438,In_595,In_1347);
xor U439 (N_439,In_566,In_532);
nand U440 (N_440,In_556,In_467);
nor U441 (N_441,In_1495,In_239);
and U442 (N_442,In_447,In_1232);
nand U443 (N_443,In_1045,In_1174);
nand U444 (N_444,In_454,In_717);
or U445 (N_445,In_184,In_1373);
and U446 (N_446,In_1179,In_975);
nand U447 (N_447,In_500,In_1186);
xnor U448 (N_448,In_503,In_1349);
nor U449 (N_449,In_428,In_277);
xor U450 (N_450,In_7,In_930);
and U451 (N_451,In_832,In_615);
nand U452 (N_452,In_675,In_678);
nand U453 (N_453,In_98,In_944);
or U454 (N_454,In_79,In_427);
and U455 (N_455,In_906,In_1303);
nand U456 (N_456,In_58,In_557);
or U457 (N_457,In_213,In_1469);
or U458 (N_458,In_1162,In_916);
nor U459 (N_459,In_1230,In_1029);
xnor U460 (N_460,In_946,In_598);
or U461 (N_461,In_912,In_1051);
nand U462 (N_462,In_833,In_1226);
or U463 (N_463,In_1002,In_1308);
or U464 (N_464,In_120,In_1254);
or U465 (N_465,In_1189,In_487);
xor U466 (N_466,In_899,In_706);
or U467 (N_467,In_172,In_349);
nand U468 (N_468,In_114,In_558);
or U469 (N_469,In_1359,In_309);
nor U470 (N_470,In_643,In_42);
nor U471 (N_471,In_1361,In_744);
or U472 (N_472,In_876,In_210);
or U473 (N_473,In_1079,In_8);
xor U474 (N_474,In_1049,In_88);
nor U475 (N_475,In_387,In_886);
nand U476 (N_476,In_232,In_577);
or U477 (N_477,In_1295,In_1322);
and U478 (N_478,In_1065,In_512);
nor U479 (N_479,In_533,In_465);
nand U480 (N_480,In_782,In_421);
and U481 (N_481,In_60,In_1104);
nand U482 (N_482,In_956,In_665);
nor U483 (N_483,In_104,In_303);
nor U484 (N_484,In_1419,In_771);
nor U485 (N_485,In_1314,In_798);
nand U486 (N_486,In_920,In_793);
nor U487 (N_487,In_866,In_1055);
or U488 (N_488,In_1225,In_758);
nand U489 (N_489,In_1261,In_148);
and U490 (N_490,In_1050,In_1375);
and U491 (N_491,In_1482,In_186);
and U492 (N_492,In_291,In_1433);
nand U493 (N_493,In_530,In_319);
and U494 (N_494,In_233,In_642);
nor U495 (N_495,In_902,In_527);
or U496 (N_496,In_834,In_1293);
or U497 (N_497,In_1043,In_1371);
xnor U498 (N_498,In_48,In_455);
and U499 (N_499,In_967,In_1346);
or U500 (N_500,In_1449,In_1008);
or U501 (N_501,In_440,In_1250);
nand U502 (N_502,In_1272,In_1396);
or U503 (N_503,In_413,In_812);
or U504 (N_504,In_169,In_1039);
nand U505 (N_505,In_345,In_843);
or U506 (N_506,In_1201,In_974);
or U507 (N_507,In_1292,In_1118);
and U508 (N_508,In_747,In_1393);
or U509 (N_509,In_292,In_1461);
nand U510 (N_510,In_1025,In_238);
nor U511 (N_511,In_696,In_1422);
and U512 (N_512,In_1260,In_318);
or U513 (N_513,In_674,In_1114);
nand U514 (N_514,In_1216,In_1047);
and U515 (N_515,In_168,In_872);
or U516 (N_516,In_476,In_1429);
nand U517 (N_517,In_473,In_1326);
nand U518 (N_518,In_850,In_1093);
or U519 (N_519,In_36,In_1052);
and U520 (N_520,In_579,In_227);
xor U521 (N_521,In_1463,In_283);
nor U522 (N_522,In_407,In_555);
or U523 (N_523,In_362,In_711);
and U524 (N_524,In_1331,In_140);
nand U525 (N_525,In_1063,In_713);
xnor U526 (N_526,In_554,In_1156);
nor U527 (N_527,In_110,In_284);
nor U528 (N_528,In_1370,In_311);
or U529 (N_529,In_762,In_763);
or U530 (N_530,In_765,In_1432);
nor U531 (N_531,In_1479,In_1020);
or U532 (N_532,In_657,In_536);
xnor U533 (N_533,In_742,In_76);
xnor U534 (N_534,In_181,In_1129);
nand U535 (N_535,In_708,In_664);
or U536 (N_536,In_1007,In_3);
nand U537 (N_537,In_621,In_792);
nor U538 (N_538,In_381,In_1452);
and U539 (N_539,In_1430,In_778);
nor U540 (N_540,In_1402,In_957);
nor U541 (N_541,In_1062,In_159);
xnor U542 (N_542,In_263,In_937);
nor U543 (N_543,In_686,In_540);
and U544 (N_544,In_497,In_43);
and U545 (N_545,In_1145,In_567);
and U546 (N_546,In_1061,In_214);
nor U547 (N_547,In_484,In_1309);
nand U548 (N_548,In_1345,In_1499);
or U549 (N_549,In_1451,In_1416);
xnor U550 (N_550,In_692,In_1121);
nor U551 (N_551,In_390,In_861);
nor U552 (N_552,In_313,In_287);
or U553 (N_553,In_1177,In_135);
xor U554 (N_554,In_1399,In_1462);
nand U555 (N_555,In_960,In_194);
and U556 (N_556,In_627,In_1196);
xnor U557 (N_557,In_680,In_463);
nor U558 (N_558,In_601,In_234);
or U559 (N_559,In_462,In_959);
xnor U560 (N_560,In_141,In_1350);
nor U561 (N_561,In_1372,In_491);
xnor U562 (N_562,In_634,In_1305);
nor U563 (N_563,In_130,In_1206);
nor U564 (N_564,In_682,In_641);
and U565 (N_565,In_911,In_395);
and U566 (N_566,In_1274,In_732);
nor U567 (N_567,In_853,In_354);
nand U568 (N_568,In_1133,In_1075);
or U569 (N_569,In_4,In_632);
xnor U570 (N_570,In_592,In_1144);
or U571 (N_571,In_751,In_61);
and U572 (N_572,In_268,In_403);
and U573 (N_573,In_1277,In_1204);
nand U574 (N_574,In_216,In_822);
nand U575 (N_575,In_898,In_1015);
or U576 (N_576,In_1319,In_1033);
nand U577 (N_577,In_919,In_193);
nand U578 (N_578,In_1492,In_1476);
and U579 (N_579,In_1041,In_894);
or U580 (N_580,In_72,In_1455);
nand U581 (N_581,In_589,In_346);
and U582 (N_582,In_1234,In_295);
nand U583 (N_583,In_377,In_1105);
nor U584 (N_584,In_271,In_470);
nor U585 (N_585,In_1494,In_986);
or U586 (N_586,In_1235,In_1192);
nand U587 (N_587,In_1199,In_299);
and U588 (N_588,In_1404,In_903);
nand U589 (N_589,In_859,In_378);
or U590 (N_590,In_1042,In_648);
and U591 (N_591,In_1323,In_123);
and U592 (N_592,In_1336,In_700);
nor U593 (N_593,In_1478,In_82);
or U594 (N_594,In_492,In_1161);
nand U595 (N_595,In_190,In_559);
or U596 (N_596,In_958,In_31);
nor U597 (N_597,In_133,In_590);
or U598 (N_598,In_1131,In_1342);
or U599 (N_599,In_265,In_928);
or U600 (N_600,In_939,In_1181);
and U601 (N_601,In_1497,In_712);
nor U602 (N_602,In_442,In_938);
nor U603 (N_603,In_968,In_1100);
nor U604 (N_604,In_1486,In_310);
and U605 (N_605,In_439,In_306);
nand U606 (N_606,In_1366,In_256);
nand U607 (N_607,In_736,In_727);
and U608 (N_608,In_149,In_731);
nor U609 (N_609,In_544,In_1171);
nor U610 (N_610,In_1099,In_129);
nor U611 (N_611,In_480,In_69);
nand U612 (N_612,In_877,In_1264);
or U613 (N_613,In_432,In_1198);
nand U614 (N_614,In_364,In_347);
or U615 (N_615,In_1169,In_406);
or U616 (N_616,In_1009,In_1406);
and U617 (N_617,In_321,In_325);
nor U618 (N_618,In_988,In_517);
xor U619 (N_619,In_1343,In_81);
nor U620 (N_620,In_842,In_630);
or U621 (N_621,In_1242,In_879);
and U622 (N_622,In_424,In_918);
and U623 (N_623,In_818,In_1334);
nand U624 (N_624,In_92,In_1076);
or U625 (N_625,In_755,In_1294);
nand U626 (N_626,In_587,In_881);
and U627 (N_627,In_93,In_1408);
or U628 (N_628,In_1329,In_73);
nand U629 (N_629,In_1236,In_68);
nand U630 (N_630,In_801,In_1158);
and U631 (N_631,In_434,In_878);
nor U632 (N_632,In_192,In_603);
nand U633 (N_633,In_1028,In_356);
or U634 (N_634,In_50,In_498);
xor U635 (N_635,In_1473,In_1381);
and U636 (N_636,In_1283,In_444);
xnor U637 (N_637,In_521,In_1352);
or U638 (N_638,In_244,In_519);
nor U639 (N_639,In_176,In_95);
or U640 (N_640,In_1324,In_929);
nor U641 (N_641,In_217,In_398);
and U642 (N_642,In_1460,In_458);
nand U643 (N_643,In_1089,In_1472);
and U644 (N_644,In_578,In_369);
and U645 (N_645,In_147,In_469);
or U646 (N_646,In_1217,In_999);
nand U647 (N_647,In_1467,In_1325);
nor U648 (N_648,In_947,In_394);
and U649 (N_649,In_482,In_1488);
and U650 (N_650,In_757,In_854);
nor U651 (N_651,In_996,In_1108);
nor U652 (N_652,In_542,In_673);
nor U653 (N_653,In_1367,In_409);
xnor U654 (N_654,In_143,In_464);
nand U655 (N_655,In_360,In_294);
nor U656 (N_656,In_950,In_1387);
or U657 (N_657,In_1363,In_718);
nor U658 (N_658,In_502,In_1498);
and U659 (N_659,In_1390,In_405);
nand U660 (N_660,In_1239,In_687);
nor U661 (N_661,In_1421,In_393);
nand U662 (N_662,In_27,In_404);
xor U663 (N_663,In_753,In_1059);
or U664 (N_664,In_1109,In_594);
nor U665 (N_665,In_15,In_139);
nand U666 (N_666,In_1128,In_1362);
or U667 (N_667,In_14,In_16);
nand U668 (N_668,In_206,In_1255);
or U669 (N_669,In_62,In_430);
and U670 (N_670,In_1339,In_705);
or U671 (N_671,In_111,In_30);
nor U672 (N_672,In_830,In_971);
and U673 (N_673,In_1018,In_874);
nand U674 (N_674,In_1247,In_253);
nor U675 (N_675,In_167,In_1307);
and U676 (N_676,In_1110,In_145);
nor U677 (N_677,In_719,In_991);
nor U678 (N_678,In_970,In_628);
nor U679 (N_679,In_166,In_200);
or U680 (N_680,In_1036,In_963);
or U681 (N_681,In_689,In_932);
nor U682 (N_682,In_28,In_1030);
and U683 (N_683,In_1435,In_1228);
or U684 (N_684,In_820,In_45);
or U685 (N_685,In_260,In_1320);
and U686 (N_686,In_189,In_205);
nand U687 (N_687,In_1107,In_819);
nor U688 (N_688,In_869,In_290);
nor U689 (N_689,In_1141,In_600);
xor U690 (N_690,In_805,In_649);
xor U691 (N_691,In_355,In_1392);
nand U692 (N_692,In_83,In_844);
nand U693 (N_693,In_640,In_278);
nand U694 (N_694,In_1278,In_666);
or U695 (N_695,In_921,In_270);
nor U696 (N_696,In_568,In_596);
nor U697 (N_697,In_1113,In_743);
and U698 (N_698,In_1300,In_741);
or U699 (N_699,In_391,In_137);
and U700 (N_700,In_331,In_67);
nand U701 (N_701,In_451,In_972);
xor U702 (N_702,In_383,In_228);
xor U703 (N_703,In_690,In_571);
nand U704 (N_704,In_1212,In_33);
or U705 (N_705,In_725,In_989);
nand U706 (N_706,In_1053,In_317);
nand U707 (N_707,In_102,In_677);
or U708 (N_708,In_1165,In_386);
xor U709 (N_709,In_890,In_1073);
nor U710 (N_710,In_326,In_663);
or U711 (N_711,In_926,In_608);
or U712 (N_712,In_547,In_1064);
nor U713 (N_713,In_1012,In_1084);
nand U714 (N_714,In_402,In_748);
and U715 (N_715,In_904,In_1142);
nor U716 (N_716,In_1299,In_789);
nand U717 (N_717,In_1046,In_1284);
xnor U718 (N_718,In_954,In_222);
and U719 (N_719,In_418,In_586);
nand U720 (N_720,In_796,In_733);
and U721 (N_721,In_672,In_1403);
or U722 (N_722,In_1243,In_546);
nand U723 (N_723,In_84,In_979);
nor U724 (N_724,In_87,In_1474);
nand U725 (N_725,In_408,In_701);
or U726 (N_726,In_106,In_1485);
nand U727 (N_727,In_650,In_376);
or U728 (N_728,In_1439,In_1426);
and U729 (N_729,In_472,In_667);
nor U730 (N_730,In_777,In_59);
or U731 (N_731,In_19,In_607);
or U732 (N_732,In_549,In_537);
xor U733 (N_733,In_235,In_998);
or U734 (N_734,In_293,In_1471);
and U735 (N_735,In_1340,In_910);
and U736 (N_736,In_209,In_1038);
nand U737 (N_737,In_811,In_1166);
and U738 (N_738,In_1151,In_343);
and U739 (N_739,In_118,In_10);
or U740 (N_740,In_1222,In_1385);
or U741 (N_741,In_276,In_754);
xnor U742 (N_742,In_54,In_1489);
nor U743 (N_743,In_414,In_1353);
and U744 (N_744,In_1446,In_961);
nand U745 (N_745,In_136,In_602);
nand U746 (N_746,In_582,In_358);
nand U747 (N_747,In_774,In_661);
and U748 (N_748,In_224,In_142);
nand U749 (N_749,In_609,In_523);
nand U750 (N_750,In_1339,In_647);
nand U751 (N_751,In_345,In_318);
or U752 (N_752,In_1140,In_1040);
and U753 (N_753,In_1141,In_1476);
or U754 (N_754,In_1294,In_553);
or U755 (N_755,In_1017,In_523);
or U756 (N_756,In_692,In_26);
nand U757 (N_757,In_661,In_1290);
nor U758 (N_758,In_462,In_808);
nor U759 (N_759,In_1203,In_124);
nand U760 (N_760,In_539,In_1389);
and U761 (N_761,In_357,In_606);
and U762 (N_762,In_215,In_456);
nor U763 (N_763,In_1079,In_1336);
and U764 (N_764,In_1102,In_804);
and U765 (N_765,In_1443,In_1473);
and U766 (N_766,In_855,In_321);
and U767 (N_767,In_797,In_81);
and U768 (N_768,In_697,In_35);
or U769 (N_769,In_1283,In_1344);
nand U770 (N_770,In_446,In_685);
or U771 (N_771,In_344,In_884);
and U772 (N_772,In_265,In_524);
nor U773 (N_773,In_854,In_870);
nand U774 (N_774,In_395,In_802);
or U775 (N_775,In_880,In_1250);
nor U776 (N_776,In_1248,In_666);
and U777 (N_777,In_1277,In_1255);
and U778 (N_778,In_1374,In_101);
xnor U779 (N_779,In_386,In_1276);
or U780 (N_780,In_380,In_1223);
and U781 (N_781,In_652,In_733);
or U782 (N_782,In_236,In_540);
nor U783 (N_783,In_170,In_161);
nand U784 (N_784,In_1318,In_38);
and U785 (N_785,In_1398,In_1184);
nor U786 (N_786,In_28,In_1155);
or U787 (N_787,In_1379,In_478);
nor U788 (N_788,In_283,In_1408);
nand U789 (N_789,In_1443,In_653);
xnor U790 (N_790,In_671,In_128);
or U791 (N_791,In_343,In_1403);
nor U792 (N_792,In_1429,In_742);
nand U793 (N_793,In_1430,In_337);
or U794 (N_794,In_347,In_772);
nor U795 (N_795,In_705,In_78);
and U796 (N_796,In_1184,In_772);
and U797 (N_797,In_123,In_1018);
nand U798 (N_798,In_1399,In_1465);
nor U799 (N_799,In_1228,In_1026);
nor U800 (N_800,In_833,In_650);
and U801 (N_801,In_356,In_993);
nor U802 (N_802,In_1106,In_150);
xnor U803 (N_803,In_13,In_892);
nor U804 (N_804,In_577,In_1063);
nor U805 (N_805,In_1032,In_322);
nand U806 (N_806,In_635,In_952);
and U807 (N_807,In_525,In_1412);
or U808 (N_808,In_8,In_823);
or U809 (N_809,In_105,In_1257);
nor U810 (N_810,In_177,In_957);
nand U811 (N_811,In_430,In_956);
nand U812 (N_812,In_499,In_698);
and U813 (N_813,In_687,In_1191);
and U814 (N_814,In_262,In_117);
nor U815 (N_815,In_58,In_5);
nor U816 (N_816,In_462,In_1394);
nand U817 (N_817,In_1465,In_1217);
and U818 (N_818,In_618,In_673);
and U819 (N_819,In_1201,In_607);
and U820 (N_820,In_1331,In_592);
or U821 (N_821,In_320,In_1364);
nand U822 (N_822,In_1286,In_1284);
nand U823 (N_823,In_814,In_3);
nor U824 (N_824,In_10,In_1128);
nand U825 (N_825,In_1038,In_51);
and U826 (N_826,In_302,In_787);
nand U827 (N_827,In_262,In_1181);
xnor U828 (N_828,In_1069,In_441);
or U829 (N_829,In_213,In_952);
and U830 (N_830,In_369,In_573);
and U831 (N_831,In_926,In_389);
and U832 (N_832,In_830,In_1458);
nand U833 (N_833,In_796,In_978);
nor U834 (N_834,In_271,In_1292);
nor U835 (N_835,In_473,In_734);
nor U836 (N_836,In_411,In_346);
and U837 (N_837,In_293,In_453);
nor U838 (N_838,In_1226,In_465);
or U839 (N_839,In_738,In_411);
nor U840 (N_840,In_121,In_725);
or U841 (N_841,In_547,In_1220);
nor U842 (N_842,In_984,In_649);
nor U843 (N_843,In_510,In_1286);
or U844 (N_844,In_1034,In_918);
nand U845 (N_845,In_1236,In_1057);
xor U846 (N_846,In_105,In_1138);
nand U847 (N_847,In_828,In_80);
and U848 (N_848,In_94,In_683);
nor U849 (N_849,In_1069,In_72);
nand U850 (N_850,In_550,In_1383);
or U851 (N_851,In_1374,In_1498);
or U852 (N_852,In_796,In_186);
nor U853 (N_853,In_112,In_82);
nand U854 (N_854,In_1212,In_393);
or U855 (N_855,In_340,In_655);
nor U856 (N_856,In_1141,In_697);
nand U857 (N_857,In_201,In_178);
and U858 (N_858,In_737,In_211);
xnor U859 (N_859,In_41,In_154);
nand U860 (N_860,In_989,In_357);
nand U861 (N_861,In_615,In_833);
xor U862 (N_862,In_881,In_664);
nor U863 (N_863,In_502,In_730);
or U864 (N_864,In_849,In_453);
or U865 (N_865,In_1328,In_900);
nand U866 (N_866,In_1083,In_852);
nor U867 (N_867,In_429,In_935);
xnor U868 (N_868,In_736,In_1149);
and U869 (N_869,In_1006,In_732);
nand U870 (N_870,In_1406,In_811);
nor U871 (N_871,In_853,In_1357);
nand U872 (N_872,In_1485,In_1463);
nor U873 (N_873,In_126,In_1108);
nor U874 (N_874,In_673,In_291);
or U875 (N_875,In_1486,In_900);
and U876 (N_876,In_1356,In_274);
nor U877 (N_877,In_439,In_105);
xnor U878 (N_878,In_1115,In_1435);
or U879 (N_879,In_136,In_786);
or U880 (N_880,In_1460,In_1034);
or U881 (N_881,In_531,In_319);
or U882 (N_882,In_217,In_176);
nor U883 (N_883,In_491,In_989);
nor U884 (N_884,In_190,In_88);
nand U885 (N_885,In_557,In_1451);
xnor U886 (N_886,In_1308,In_402);
nand U887 (N_887,In_923,In_317);
and U888 (N_888,In_418,In_1207);
nor U889 (N_889,In_1240,In_342);
nor U890 (N_890,In_737,In_1380);
and U891 (N_891,In_173,In_540);
nand U892 (N_892,In_648,In_1006);
and U893 (N_893,In_1406,In_507);
nor U894 (N_894,In_1178,In_794);
nand U895 (N_895,In_141,In_1397);
or U896 (N_896,In_373,In_556);
and U897 (N_897,In_208,In_1325);
nand U898 (N_898,In_757,In_1238);
xnor U899 (N_899,In_653,In_1008);
and U900 (N_900,In_768,In_530);
or U901 (N_901,In_204,In_993);
xor U902 (N_902,In_1183,In_145);
nand U903 (N_903,In_358,In_639);
nor U904 (N_904,In_307,In_256);
nand U905 (N_905,In_917,In_978);
nor U906 (N_906,In_28,In_861);
nor U907 (N_907,In_226,In_954);
or U908 (N_908,In_394,In_80);
or U909 (N_909,In_904,In_1224);
and U910 (N_910,In_394,In_1137);
nor U911 (N_911,In_851,In_365);
and U912 (N_912,In_497,In_955);
nand U913 (N_913,In_35,In_659);
and U914 (N_914,In_185,In_580);
nor U915 (N_915,In_540,In_45);
nor U916 (N_916,In_1382,In_157);
nand U917 (N_917,In_1142,In_448);
and U918 (N_918,In_1057,In_155);
or U919 (N_919,In_1360,In_1256);
or U920 (N_920,In_60,In_610);
xor U921 (N_921,In_308,In_483);
and U922 (N_922,In_1143,In_96);
and U923 (N_923,In_342,In_1324);
nand U924 (N_924,In_1356,In_347);
nand U925 (N_925,In_1237,In_1277);
nand U926 (N_926,In_972,In_1486);
or U927 (N_927,In_879,In_594);
or U928 (N_928,In_260,In_1031);
or U929 (N_929,In_1347,In_65);
and U930 (N_930,In_596,In_45);
nor U931 (N_931,In_611,In_1382);
nand U932 (N_932,In_67,In_543);
nand U933 (N_933,In_351,In_605);
and U934 (N_934,In_105,In_1105);
nand U935 (N_935,In_1353,In_638);
or U936 (N_936,In_792,In_1166);
and U937 (N_937,In_1450,In_741);
or U938 (N_938,In_1070,In_371);
or U939 (N_939,In_505,In_1230);
nand U940 (N_940,In_564,In_407);
nand U941 (N_941,In_1080,In_367);
nor U942 (N_942,In_671,In_1048);
nor U943 (N_943,In_926,In_121);
nand U944 (N_944,In_1330,In_399);
xnor U945 (N_945,In_1069,In_288);
nand U946 (N_946,In_479,In_1162);
nor U947 (N_947,In_82,In_1212);
or U948 (N_948,In_969,In_1143);
and U949 (N_949,In_1320,In_1417);
nand U950 (N_950,In_1336,In_632);
nand U951 (N_951,In_105,In_229);
nor U952 (N_952,In_970,In_842);
or U953 (N_953,In_958,In_640);
nand U954 (N_954,In_898,In_746);
nand U955 (N_955,In_251,In_304);
or U956 (N_956,In_698,In_869);
nand U957 (N_957,In_801,In_1041);
or U958 (N_958,In_216,In_709);
nand U959 (N_959,In_276,In_1302);
nor U960 (N_960,In_943,In_354);
and U961 (N_961,In_1079,In_1016);
nor U962 (N_962,In_980,In_763);
and U963 (N_963,In_1094,In_1022);
xnor U964 (N_964,In_1452,In_695);
nor U965 (N_965,In_1459,In_383);
nor U966 (N_966,In_27,In_97);
nand U967 (N_967,In_241,In_1222);
nor U968 (N_968,In_657,In_1484);
nand U969 (N_969,In_665,In_1458);
nor U970 (N_970,In_899,In_362);
nand U971 (N_971,In_714,In_1035);
nand U972 (N_972,In_1453,In_231);
nor U973 (N_973,In_358,In_1053);
nand U974 (N_974,In_866,In_59);
xnor U975 (N_975,In_951,In_758);
and U976 (N_976,In_1176,In_146);
or U977 (N_977,In_269,In_1108);
and U978 (N_978,In_173,In_764);
or U979 (N_979,In_1473,In_61);
xnor U980 (N_980,In_1143,In_200);
nor U981 (N_981,In_1284,In_291);
and U982 (N_982,In_785,In_290);
nor U983 (N_983,In_1022,In_890);
nand U984 (N_984,In_452,In_576);
xor U985 (N_985,In_1047,In_100);
and U986 (N_986,In_871,In_793);
nand U987 (N_987,In_1347,In_130);
nor U988 (N_988,In_1239,In_158);
and U989 (N_989,In_945,In_1135);
and U990 (N_990,In_1355,In_599);
nor U991 (N_991,In_340,In_334);
xnor U992 (N_992,In_348,In_1160);
nand U993 (N_993,In_724,In_1373);
nand U994 (N_994,In_633,In_406);
nor U995 (N_995,In_1165,In_35);
and U996 (N_996,In_1010,In_824);
and U997 (N_997,In_1402,In_566);
and U998 (N_998,In_347,In_421);
or U999 (N_999,In_669,In_1179);
or U1000 (N_1000,N_106,N_433);
nor U1001 (N_1001,N_154,N_972);
or U1002 (N_1002,N_490,N_137);
and U1003 (N_1003,N_666,N_928);
and U1004 (N_1004,N_477,N_424);
and U1005 (N_1005,N_686,N_521);
xnor U1006 (N_1006,N_634,N_791);
nand U1007 (N_1007,N_60,N_245);
nor U1008 (N_1008,N_779,N_39);
and U1009 (N_1009,N_738,N_565);
nand U1010 (N_1010,N_994,N_488);
nand U1011 (N_1011,N_407,N_473);
or U1012 (N_1012,N_96,N_760);
or U1013 (N_1013,N_489,N_648);
or U1014 (N_1014,N_415,N_107);
or U1015 (N_1015,N_177,N_935);
and U1016 (N_1016,N_331,N_194);
nand U1017 (N_1017,N_764,N_729);
nand U1018 (N_1018,N_139,N_581);
nor U1019 (N_1019,N_924,N_386);
or U1020 (N_1020,N_468,N_753);
nand U1021 (N_1021,N_66,N_153);
and U1022 (N_1022,N_905,N_838);
nand U1023 (N_1023,N_512,N_885);
or U1024 (N_1024,N_731,N_541);
or U1025 (N_1025,N_495,N_48);
nand U1026 (N_1026,N_151,N_175);
nor U1027 (N_1027,N_528,N_134);
nor U1028 (N_1028,N_500,N_567);
and U1029 (N_1029,N_882,N_769);
or U1030 (N_1030,N_78,N_827);
and U1031 (N_1031,N_171,N_448);
xor U1032 (N_1032,N_94,N_683);
and U1033 (N_1033,N_427,N_915);
nor U1034 (N_1034,N_985,N_259);
xnor U1035 (N_1035,N_75,N_74);
nor U1036 (N_1036,N_966,N_146);
nand U1037 (N_1037,N_609,N_166);
xnor U1038 (N_1038,N_923,N_384);
nor U1039 (N_1039,N_230,N_102);
xor U1040 (N_1040,N_796,N_510);
or U1041 (N_1041,N_92,N_933);
and U1042 (N_1042,N_740,N_774);
nor U1043 (N_1043,N_709,N_948);
or U1044 (N_1044,N_294,N_958);
or U1045 (N_1045,N_292,N_271);
nand U1046 (N_1046,N_221,N_76);
and U1047 (N_1047,N_464,N_345);
nor U1048 (N_1048,N_17,N_700);
and U1049 (N_1049,N_636,N_785);
nor U1050 (N_1050,N_472,N_428);
or U1051 (N_1051,N_998,N_670);
and U1052 (N_1052,N_291,N_243);
nor U1053 (N_1053,N_635,N_531);
nor U1054 (N_1054,N_632,N_560);
nand U1055 (N_1055,N_550,N_114);
or U1056 (N_1056,N_737,N_72);
nor U1057 (N_1057,N_867,N_274);
and U1058 (N_1058,N_982,N_810);
xnor U1059 (N_1059,N_147,N_113);
xor U1060 (N_1060,N_398,N_319);
nand U1061 (N_1061,N_617,N_685);
and U1062 (N_1062,N_936,N_820);
and U1063 (N_1063,N_318,N_711);
or U1064 (N_1064,N_367,N_187);
or U1065 (N_1065,N_359,N_226);
or U1066 (N_1066,N_911,N_695);
or U1067 (N_1067,N_903,N_725);
xnor U1068 (N_1068,N_880,N_423);
nor U1069 (N_1069,N_556,N_614);
and U1070 (N_1070,N_437,N_397);
nand U1071 (N_1071,N_688,N_976);
nand U1072 (N_1072,N_492,N_482);
or U1073 (N_1073,N_912,N_138);
xnor U1074 (N_1074,N_582,N_45);
or U1075 (N_1075,N_620,N_741);
nor U1076 (N_1076,N_768,N_209);
xor U1077 (N_1077,N_507,N_111);
and U1078 (N_1078,N_651,N_947);
or U1079 (N_1079,N_354,N_261);
and U1080 (N_1080,N_6,N_623);
and U1081 (N_1081,N_411,N_952);
or U1082 (N_1082,N_997,N_401);
or U1083 (N_1083,N_414,N_619);
xnor U1084 (N_1084,N_536,N_157);
and U1085 (N_1085,N_256,N_506);
or U1086 (N_1086,N_937,N_594);
xnor U1087 (N_1087,N_290,N_461);
or U1088 (N_1088,N_100,N_26);
nand U1089 (N_1089,N_302,N_999);
or U1090 (N_1090,N_744,N_578);
or U1091 (N_1091,N_719,N_450);
or U1092 (N_1092,N_108,N_38);
nor U1093 (N_1093,N_965,N_773);
nor U1094 (N_1094,N_534,N_913);
xor U1095 (N_1095,N_28,N_844);
nand U1096 (N_1096,N_54,N_178);
or U1097 (N_1097,N_15,N_983);
or U1098 (N_1098,N_210,N_69);
nor U1099 (N_1099,N_877,N_723);
and U1100 (N_1100,N_504,N_950);
or U1101 (N_1101,N_373,N_203);
nor U1102 (N_1102,N_745,N_81);
nand U1103 (N_1103,N_197,N_961);
nor U1104 (N_1104,N_44,N_992);
or U1105 (N_1105,N_35,N_172);
or U1106 (N_1106,N_806,N_347);
nand U1107 (N_1107,N_861,N_771);
xnor U1108 (N_1108,N_758,N_416);
and U1109 (N_1109,N_342,N_25);
nor U1110 (N_1110,N_809,N_975);
nand U1111 (N_1111,N_660,N_142);
xor U1112 (N_1112,N_988,N_590);
or U1113 (N_1113,N_244,N_351);
and U1114 (N_1114,N_756,N_735);
nor U1115 (N_1115,N_353,N_665);
nor U1116 (N_1116,N_165,N_377);
and U1117 (N_1117,N_324,N_370);
or U1118 (N_1118,N_963,N_730);
nand U1119 (N_1119,N_276,N_846);
nand U1120 (N_1120,N_339,N_253);
and U1121 (N_1121,N_555,N_859);
xor U1122 (N_1122,N_97,N_974);
nand U1123 (N_1123,N_224,N_158);
or U1124 (N_1124,N_707,N_368);
or U1125 (N_1125,N_229,N_549);
or U1126 (N_1126,N_195,N_479);
or U1127 (N_1127,N_518,N_393);
and U1128 (N_1128,N_257,N_691);
and U1129 (N_1129,N_727,N_445);
nor U1130 (N_1130,N_340,N_193);
xor U1131 (N_1131,N_40,N_798);
and U1132 (N_1132,N_833,N_890);
nand U1133 (N_1133,N_501,N_484);
or U1134 (N_1134,N_973,N_687);
nand U1135 (N_1135,N_854,N_625);
nor U1136 (N_1136,N_326,N_442);
nand U1137 (N_1137,N_465,N_509);
nand U1138 (N_1138,N_65,N_979);
or U1139 (N_1139,N_770,N_250);
and U1140 (N_1140,N_378,N_749);
nand U1141 (N_1141,N_466,N_304);
and U1142 (N_1142,N_894,N_438);
or U1143 (N_1143,N_120,N_830);
or U1144 (N_1144,N_184,N_851);
or U1145 (N_1145,N_904,N_321);
or U1146 (N_1146,N_786,N_382);
or U1147 (N_1147,N_778,N_191);
nor U1148 (N_1148,N_128,N_18);
nor U1149 (N_1149,N_82,N_824);
nand U1150 (N_1150,N_951,N_538);
or U1151 (N_1151,N_369,N_646);
nand U1152 (N_1152,N_641,N_588);
or U1153 (N_1153,N_713,N_576);
and U1154 (N_1154,N_944,N_611);
or U1155 (N_1155,N_858,N_739);
xor U1156 (N_1156,N_306,N_322);
nand U1157 (N_1157,N_355,N_19);
or U1158 (N_1158,N_70,N_957);
xnor U1159 (N_1159,N_170,N_669);
xnor U1160 (N_1160,N_516,N_412);
nand U1161 (N_1161,N_458,N_857);
xor U1162 (N_1162,N_453,N_562);
nand U1163 (N_1163,N_33,N_606);
nand U1164 (N_1164,N_527,N_467);
and U1165 (N_1165,N_199,N_405);
nor U1166 (N_1166,N_246,N_9);
or U1167 (N_1167,N_227,N_540);
nand U1168 (N_1168,N_255,N_312);
and U1169 (N_1169,N_551,N_471);
and U1170 (N_1170,N_907,N_742);
or U1171 (N_1171,N_47,N_986);
nor U1172 (N_1172,N_396,N_273);
and U1173 (N_1173,N_736,N_2);
nor U1174 (N_1174,N_494,N_637);
or U1175 (N_1175,N_116,N_365);
nand U1176 (N_1176,N_788,N_478);
and U1177 (N_1177,N_547,N_176);
or U1178 (N_1178,N_808,N_649);
nand U1179 (N_1179,N_394,N_168);
nand U1180 (N_1180,N_657,N_743);
xnor U1181 (N_1181,N_161,N_557);
and U1182 (N_1182,N_252,N_895);
or U1183 (N_1183,N_505,N_891);
nand U1184 (N_1184,N_887,N_628);
nor U1185 (N_1185,N_647,N_835);
xor U1186 (N_1186,N_457,N_863);
and U1187 (N_1187,N_520,N_783);
or U1188 (N_1188,N_941,N_497);
nor U1189 (N_1189,N_874,N_62);
nor U1190 (N_1190,N_127,N_43);
and U1191 (N_1191,N_260,N_926);
and U1192 (N_1192,N_480,N_109);
xnor U1193 (N_1193,N_186,N_240);
nand U1194 (N_1194,N_288,N_645);
and U1195 (N_1195,N_362,N_802);
nand U1196 (N_1196,N_971,N_52);
nand U1197 (N_1197,N_539,N_558);
nor U1198 (N_1198,N_277,N_295);
and U1199 (N_1199,N_722,N_279);
and U1200 (N_1200,N_875,N_222);
and U1201 (N_1201,N_409,N_4);
nor U1202 (N_1202,N_462,N_441);
xor U1203 (N_1203,N_608,N_853);
and U1204 (N_1204,N_254,N_852);
nand U1205 (N_1205,N_297,N_36);
nor U1206 (N_1206,N_63,N_389);
nand U1207 (N_1207,N_570,N_275);
xor U1208 (N_1208,N_443,N_855);
nor U1209 (N_1209,N_383,N_548);
xnor U1210 (N_1210,N_860,N_233);
and U1211 (N_1211,N_434,N_671);
nand U1212 (N_1212,N_826,N_598);
or U1213 (N_1213,N_865,N_41);
nand U1214 (N_1214,N_699,N_970);
or U1215 (N_1215,N_643,N_893);
and U1216 (N_1216,N_262,N_470);
and U1217 (N_1217,N_511,N_589);
nand U1218 (N_1218,N_385,N_990);
and U1219 (N_1219,N_150,N_420);
nand U1220 (N_1220,N_638,N_610);
or U1221 (N_1221,N_718,N_902);
nor U1222 (N_1222,N_626,N_217);
nand U1223 (N_1223,N_658,N_751);
nand U1224 (N_1224,N_403,N_429);
nor U1225 (N_1225,N_118,N_16);
or U1226 (N_1226,N_231,N_781);
nor U1227 (N_1227,N_616,N_164);
nor U1228 (N_1228,N_301,N_836);
nand U1229 (N_1229,N_303,N_964);
and U1230 (N_1230,N_159,N_757);
xnor U1231 (N_1231,N_5,N_661);
or U1232 (N_1232,N_12,N_934);
and U1233 (N_1233,N_573,N_604);
xnor U1234 (N_1234,N_870,N_659);
nand U1235 (N_1235,N_375,N_56);
nor U1236 (N_1236,N_358,N_721);
or U1237 (N_1237,N_705,N_234);
nand U1238 (N_1238,N_901,N_90);
nor U1239 (N_1239,N_91,N_77);
nand U1240 (N_1240,N_432,N_816);
nand U1241 (N_1241,N_122,N_828);
and U1242 (N_1242,N_336,N_247);
and U1243 (N_1243,N_676,N_525);
nand U1244 (N_1244,N_121,N_395);
or U1245 (N_1245,N_921,N_694);
nand U1246 (N_1246,N_64,N_529);
nand U1247 (N_1247,N_829,N_612);
or U1248 (N_1248,N_115,N_602);
nor U1249 (N_1249,N_207,N_272);
and U1250 (N_1250,N_591,N_282);
nor U1251 (N_1251,N_190,N_130);
and U1252 (N_1252,N_883,N_156);
or U1253 (N_1253,N_960,N_3);
or U1254 (N_1254,N_328,N_330);
and U1255 (N_1255,N_714,N_821);
and U1256 (N_1256,N_878,N_919);
nand U1257 (N_1257,N_579,N_173);
or U1258 (N_1258,N_55,N_697);
nand U1259 (N_1259,N_334,N_668);
nand U1260 (N_1260,N_248,N_129);
xnor U1261 (N_1261,N_496,N_922);
nand U1262 (N_1262,N_677,N_126);
and U1263 (N_1263,N_814,N_580);
nand U1264 (N_1264,N_103,N_640);
nor U1265 (N_1265,N_662,N_864);
xnor U1266 (N_1266,N_624,N_644);
xnor U1267 (N_1267,N_402,N_514);
or U1268 (N_1268,N_879,N_361);
or U1269 (N_1269,N_568,N_469);
nor U1270 (N_1270,N_553,N_117);
nand U1271 (N_1271,N_325,N_93);
nand U1272 (N_1272,N_376,N_728);
nor U1273 (N_1273,N_241,N_296);
nand U1274 (N_1274,N_873,N_452);
and U1275 (N_1275,N_703,N_439);
nor U1276 (N_1276,N_68,N_815);
nor U1277 (N_1277,N_112,N_978);
and U1278 (N_1278,N_889,N_654);
and U1279 (N_1279,N_615,N_782);
nor U1280 (N_1280,N_991,N_818);
nor U1281 (N_1281,N_430,N_344);
and U1282 (N_1282,N_898,N_185);
nand U1283 (N_1283,N_704,N_475);
xor U1284 (N_1284,N_653,N_696);
and U1285 (N_1285,N_338,N_236);
or U1286 (N_1286,N_198,N_455);
and U1287 (N_1287,N_583,N_67);
nor U1288 (N_1288,N_357,N_84);
xor U1289 (N_1289,N_140,N_599);
and U1290 (N_1290,N_216,N_350);
and U1291 (N_1291,N_546,N_503);
and U1292 (N_1292,N_425,N_715);
nand U1293 (N_1293,N_881,N_208);
or U1294 (N_1294,N_679,N_87);
nor U1295 (N_1295,N_223,N_352);
nor U1296 (N_1296,N_840,N_752);
nor U1297 (N_1297,N_968,N_99);
nor U1298 (N_1298,N_20,N_278);
nand U1299 (N_1299,N_487,N_285);
and U1300 (N_1300,N_46,N_967);
nand U1301 (N_1301,N_772,N_535);
nand U1302 (N_1302,N_513,N_459);
and U1303 (N_1303,N_832,N_733);
xnor U1304 (N_1304,N_849,N_572);
nor U1305 (N_1305,N_410,N_141);
nor U1306 (N_1306,N_613,N_329);
nor U1307 (N_1307,N_213,N_673);
nand U1308 (N_1308,N_10,N_57);
nand U1309 (N_1309,N_61,N_238);
and U1310 (N_1310,N_940,N_413);
and U1311 (N_1311,N_119,N_789);
nor U1312 (N_1312,N_943,N_268);
nand U1313 (N_1313,N_766,N_419);
nor U1314 (N_1314,N_431,N_989);
or U1315 (N_1315,N_239,N_460);
and U1316 (N_1316,N_508,N_848);
nand U1317 (N_1317,N_908,N_220);
and U1318 (N_1318,N_58,N_435);
or U1319 (N_1319,N_201,N_311);
nand U1320 (N_1320,N_53,N_537);
and U1321 (N_1321,N_135,N_862);
nand U1322 (N_1322,N_123,N_436);
xnor U1323 (N_1323,N_110,N_313);
or U1324 (N_1324,N_680,N_42);
or U1325 (N_1325,N_163,N_561);
xnor U1326 (N_1326,N_88,N_249);
and U1327 (N_1327,N_211,N_633);
nand U1328 (N_1328,N_346,N_639);
and U1329 (N_1329,N_754,N_984);
or U1330 (N_1330,N_200,N_544);
nor U1331 (N_1331,N_242,N_869);
nand U1332 (N_1332,N_600,N_759);
or U1333 (N_1333,N_499,N_631);
nor U1334 (N_1334,N_552,N_732);
or U1335 (N_1335,N_51,N_834);
nand U1336 (N_1336,N_235,N_954);
and U1337 (N_1337,N_196,N_839);
or U1338 (N_1338,N_945,N_916);
or U1339 (N_1339,N_283,N_763);
nand U1340 (N_1340,N_392,N_664);
nor U1341 (N_1341,N_144,N_517);
xor U1342 (N_1342,N_627,N_847);
nand U1343 (N_1343,N_794,N_426);
or U1344 (N_1344,N_674,N_189);
nand U1345 (N_1345,N_765,N_896);
or U1346 (N_1346,N_298,N_927);
or U1347 (N_1347,N_577,N_474);
xnor U1348 (N_1348,N_86,N_388);
nor U1349 (N_1349,N_803,N_335);
or U1350 (N_1350,N_603,N_932);
or U1351 (N_1351,N_183,N_83);
or U1352 (N_1352,N_162,N_287);
and U1353 (N_1353,N_485,N_149);
and U1354 (N_1354,N_486,N_899);
nand U1355 (N_1355,N_85,N_931);
and U1356 (N_1356,N_289,N_218);
and U1357 (N_1357,N_897,N_845);
nor U1358 (N_1358,N_314,N_710);
and U1359 (N_1359,N_205,N_996);
nand U1360 (N_1360,N_981,N_799);
and U1361 (N_1361,N_366,N_206);
or U1362 (N_1362,N_569,N_575);
or U1363 (N_1363,N_237,N_349);
and U1364 (N_1364,N_447,N_136);
nor U1365 (N_1365,N_571,N_21);
or U1366 (N_1366,N_400,N_792);
xor U1367 (N_1367,N_73,N_790);
and U1368 (N_1368,N_8,N_27);
nor U1369 (N_1369,N_596,N_800);
xnor U1370 (N_1370,N_251,N_956);
nand U1371 (N_1371,N_762,N_805);
nand U1372 (N_1372,N_31,N_502);
or U1373 (N_1373,N_71,N_174);
or U1374 (N_1374,N_160,N_925);
or U1375 (N_1375,N_585,N_124);
nand U1376 (N_1376,N_219,N_315);
nor U1377 (N_1377,N_797,N_299);
nand U1378 (N_1378,N_724,N_446);
or U1379 (N_1379,N_871,N_24);
or U1380 (N_1380,N_152,N_374);
nand U1381 (N_1381,N_59,N_281);
and U1382 (N_1382,N_483,N_748);
and U1383 (N_1383,N_258,N_148);
and U1384 (N_1384,N_906,N_418);
or U1385 (N_1385,N_980,N_49);
nand U1386 (N_1386,N_390,N_716);
and U1387 (N_1387,N_702,N_656);
nand U1388 (N_1388,N_309,N_761);
and U1389 (N_1389,N_812,N_391);
and U1390 (N_1390,N_689,N_892);
or U1391 (N_1391,N_13,N_678);
nor U1392 (N_1392,N_684,N_543);
and U1393 (N_1393,N_995,N_920);
and U1394 (N_1394,N_607,N_372);
and U1395 (N_1395,N_532,N_0);
xor U1396 (N_1396,N_942,N_95);
nor U1397 (N_1397,N_655,N_300);
nor U1398 (N_1398,N_650,N_690);
and U1399 (N_1399,N_566,N_232);
or U1400 (N_1400,N_712,N_652);
and U1401 (N_1401,N_337,N_167);
nand U1402 (N_1402,N_630,N_182);
nor U1403 (N_1403,N_850,N_180);
xnor U1404 (N_1404,N_316,N_969);
nor U1405 (N_1405,N_593,N_962);
and U1406 (N_1406,N_456,N_381);
nand U1407 (N_1407,N_533,N_422);
nor U1408 (N_1408,N_542,N_842);
nor U1409 (N_1409,N_701,N_519);
or U1410 (N_1410,N_597,N_179);
xor U1411 (N_1411,N_987,N_399);
nor U1412 (N_1412,N_1,N_563);
or U1413 (N_1413,N_32,N_214);
or U1414 (N_1414,N_938,N_79);
nand U1415 (N_1415,N_305,N_621);
nand U1416 (N_1416,N_793,N_837);
nand U1417 (N_1417,N_204,N_498);
and U1418 (N_1418,N_601,N_310);
and U1419 (N_1419,N_841,N_417);
and U1420 (N_1420,N_605,N_586);
xor U1421 (N_1421,N_269,N_667);
and U1422 (N_1422,N_900,N_155);
nor U1423 (N_1423,N_22,N_672);
nand U1424 (N_1424,N_132,N_918);
nor U1425 (N_1425,N_34,N_408);
or U1426 (N_1426,N_584,N_522);
and U1427 (N_1427,N_681,N_284);
nor U1428 (N_1428,N_622,N_192);
nor U1429 (N_1429,N_360,N_949);
or U1430 (N_1430,N_491,N_663);
nor U1431 (N_1431,N_267,N_775);
nand U1432 (N_1432,N_831,N_286);
nand U1433 (N_1433,N_866,N_145);
and U1434 (N_1434,N_526,N_265);
nor U1435 (N_1435,N_341,N_888);
nand U1436 (N_1436,N_440,N_706);
or U1437 (N_1437,N_225,N_993);
nand U1438 (N_1438,N_188,N_101);
or U1439 (N_1439,N_228,N_293);
and U1440 (N_1440,N_574,N_787);
nor U1441 (N_1441,N_939,N_872);
or U1442 (N_1442,N_7,N_317);
nand U1443 (N_1443,N_953,N_30);
or U1444 (N_1444,N_332,N_776);
and U1445 (N_1445,N_618,N_817);
nor U1446 (N_1446,N_955,N_559);
or U1447 (N_1447,N_929,N_780);
nor U1448 (N_1448,N_29,N_50);
xor U1449 (N_1449,N_777,N_451);
and U1450 (N_1450,N_587,N_554);
and U1451 (N_1451,N_530,N_977);
nand U1452 (N_1452,N_454,N_327);
or U1453 (N_1453,N_343,N_524);
xnor U1454 (N_1454,N_734,N_682);
or U1455 (N_1455,N_37,N_876);
nand U1456 (N_1456,N_80,N_14);
or U1457 (N_1457,N_592,N_421);
and U1458 (N_1458,N_819,N_856);
xnor U1459 (N_1459,N_755,N_125);
nor U1460 (N_1460,N_804,N_181);
nor U1461 (N_1461,N_169,N_105);
or U1462 (N_1462,N_463,N_811);
or U1463 (N_1463,N_215,N_476);
or U1464 (N_1464,N_323,N_212);
nand U1465 (N_1465,N_692,N_917);
nor U1466 (N_1466,N_909,N_822);
and U1467 (N_1467,N_364,N_406);
and U1468 (N_1468,N_801,N_843);
and U1469 (N_1469,N_143,N_98);
nor U1470 (N_1470,N_642,N_750);
nor U1471 (N_1471,N_449,N_444);
or U1472 (N_1472,N_868,N_356);
nor U1473 (N_1473,N_266,N_675);
nor U1474 (N_1474,N_348,N_308);
nand U1475 (N_1475,N_795,N_333);
xnor U1476 (N_1476,N_363,N_930);
or U1477 (N_1477,N_11,N_823);
and U1478 (N_1478,N_629,N_280);
nand U1479 (N_1479,N_914,N_131);
nand U1480 (N_1480,N_813,N_545);
nand U1481 (N_1481,N_264,N_380);
and U1482 (N_1482,N_784,N_89);
nand U1483 (N_1483,N_133,N_746);
xnor U1484 (N_1484,N_886,N_693);
and U1485 (N_1485,N_884,N_726);
xnor U1486 (N_1486,N_595,N_910);
or U1487 (N_1487,N_263,N_404);
or U1488 (N_1488,N_320,N_23);
or U1489 (N_1489,N_720,N_202);
xnor U1490 (N_1490,N_767,N_523);
nor U1491 (N_1491,N_708,N_387);
nor U1492 (N_1492,N_481,N_515);
nor U1493 (N_1493,N_825,N_946);
and U1494 (N_1494,N_564,N_959);
xor U1495 (N_1495,N_717,N_747);
xnor U1496 (N_1496,N_307,N_371);
or U1497 (N_1497,N_807,N_270);
nor U1498 (N_1498,N_104,N_698);
or U1499 (N_1499,N_493,N_379);
nor U1500 (N_1500,N_566,N_188);
and U1501 (N_1501,N_60,N_604);
and U1502 (N_1502,N_539,N_158);
and U1503 (N_1503,N_868,N_307);
nor U1504 (N_1504,N_704,N_758);
or U1505 (N_1505,N_730,N_718);
nand U1506 (N_1506,N_875,N_645);
nor U1507 (N_1507,N_81,N_274);
and U1508 (N_1508,N_40,N_759);
and U1509 (N_1509,N_6,N_28);
xor U1510 (N_1510,N_342,N_561);
nand U1511 (N_1511,N_199,N_306);
or U1512 (N_1512,N_251,N_518);
or U1513 (N_1513,N_330,N_484);
and U1514 (N_1514,N_459,N_674);
and U1515 (N_1515,N_222,N_897);
or U1516 (N_1516,N_521,N_605);
or U1517 (N_1517,N_994,N_152);
and U1518 (N_1518,N_527,N_702);
nor U1519 (N_1519,N_589,N_470);
nand U1520 (N_1520,N_973,N_396);
and U1521 (N_1521,N_784,N_653);
nor U1522 (N_1522,N_889,N_446);
and U1523 (N_1523,N_582,N_757);
nor U1524 (N_1524,N_740,N_647);
or U1525 (N_1525,N_627,N_718);
nand U1526 (N_1526,N_195,N_409);
and U1527 (N_1527,N_394,N_999);
nand U1528 (N_1528,N_487,N_207);
nand U1529 (N_1529,N_60,N_893);
nor U1530 (N_1530,N_89,N_447);
nor U1531 (N_1531,N_659,N_250);
or U1532 (N_1532,N_943,N_296);
nand U1533 (N_1533,N_528,N_125);
nor U1534 (N_1534,N_523,N_585);
and U1535 (N_1535,N_113,N_236);
and U1536 (N_1536,N_447,N_40);
or U1537 (N_1537,N_942,N_678);
nor U1538 (N_1538,N_120,N_704);
or U1539 (N_1539,N_763,N_709);
nand U1540 (N_1540,N_928,N_365);
nand U1541 (N_1541,N_725,N_548);
nand U1542 (N_1542,N_296,N_162);
or U1543 (N_1543,N_139,N_240);
nand U1544 (N_1544,N_780,N_18);
or U1545 (N_1545,N_304,N_837);
or U1546 (N_1546,N_454,N_510);
and U1547 (N_1547,N_64,N_700);
nand U1548 (N_1548,N_750,N_499);
nand U1549 (N_1549,N_664,N_366);
or U1550 (N_1550,N_514,N_245);
nand U1551 (N_1551,N_404,N_882);
or U1552 (N_1552,N_645,N_741);
or U1553 (N_1553,N_838,N_39);
nand U1554 (N_1554,N_698,N_348);
nand U1555 (N_1555,N_719,N_215);
or U1556 (N_1556,N_689,N_809);
or U1557 (N_1557,N_247,N_727);
xnor U1558 (N_1558,N_36,N_660);
nand U1559 (N_1559,N_777,N_536);
or U1560 (N_1560,N_833,N_939);
or U1561 (N_1561,N_297,N_410);
xor U1562 (N_1562,N_474,N_557);
nand U1563 (N_1563,N_35,N_951);
and U1564 (N_1564,N_314,N_621);
nand U1565 (N_1565,N_779,N_390);
and U1566 (N_1566,N_712,N_541);
or U1567 (N_1567,N_287,N_820);
nor U1568 (N_1568,N_726,N_494);
nand U1569 (N_1569,N_528,N_435);
nand U1570 (N_1570,N_618,N_954);
and U1571 (N_1571,N_116,N_525);
and U1572 (N_1572,N_626,N_530);
nand U1573 (N_1573,N_503,N_568);
nor U1574 (N_1574,N_409,N_281);
nand U1575 (N_1575,N_262,N_736);
and U1576 (N_1576,N_928,N_706);
nor U1577 (N_1577,N_747,N_173);
or U1578 (N_1578,N_361,N_569);
or U1579 (N_1579,N_173,N_602);
and U1580 (N_1580,N_299,N_143);
nor U1581 (N_1581,N_358,N_980);
xnor U1582 (N_1582,N_917,N_808);
nor U1583 (N_1583,N_734,N_687);
nor U1584 (N_1584,N_705,N_473);
nor U1585 (N_1585,N_389,N_116);
and U1586 (N_1586,N_351,N_280);
nand U1587 (N_1587,N_233,N_730);
or U1588 (N_1588,N_141,N_614);
nor U1589 (N_1589,N_6,N_670);
nand U1590 (N_1590,N_166,N_472);
nand U1591 (N_1591,N_592,N_747);
xor U1592 (N_1592,N_236,N_310);
xor U1593 (N_1593,N_409,N_31);
nand U1594 (N_1594,N_423,N_612);
nor U1595 (N_1595,N_458,N_721);
nand U1596 (N_1596,N_412,N_595);
and U1597 (N_1597,N_466,N_836);
or U1598 (N_1598,N_672,N_637);
xnor U1599 (N_1599,N_41,N_494);
or U1600 (N_1600,N_409,N_292);
or U1601 (N_1601,N_528,N_57);
nand U1602 (N_1602,N_481,N_19);
or U1603 (N_1603,N_248,N_221);
or U1604 (N_1604,N_483,N_686);
nand U1605 (N_1605,N_556,N_737);
nor U1606 (N_1606,N_76,N_41);
xor U1607 (N_1607,N_261,N_229);
nand U1608 (N_1608,N_653,N_594);
or U1609 (N_1609,N_769,N_606);
xnor U1610 (N_1610,N_297,N_488);
nor U1611 (N_1611,N_38,N_27);
nor U1612 (N_1612,N_966,N_575);
nor U1613 (N_1613,N_413,N_145);
and U1614 (N_1614,N_526,N_432);
nand U1615 (N_1615,N_407,N_307);
or U1616 (N_1616,N_50,N_511);
and U1617 (N_1617,N_225,N_735);
nand U1618 (N_1618,N_726,N_624);
or U1619 (N_1619,N_317,N_807);
nand U1620 (N_1620,N_499,N_984);
and U1621 (N_1621,N_498,N_742);
and U1622 (N_1622,N_467,N_157);
xor U1623 (N_1623,N_617,N_373);
nand U1624 (N_1624,N_172,N_292);
nor U1625 (N_1625,N_566,N_311);
nor U1626 (N_1626,N_86,N_138);
or U1627 (N_1627,N_333,N_197);
or U1628 (N_1628,N_860,N_141);
nor U1629 (N_1629,N_900,N_424);
and U1630 (N_1630,N_882,N_959);
nor U1631 (N_1631,N_784,N_573);
nand U1632 (N_1632,N_748,N_310);
and U1633 (N_1633,N_130,N_820);
or U1634 (N_1634,N_549,N_585);
xor U1635 (N_1635,N_361,N_669);
nand U1636 (N_1636,N_923,N_107);
nand U1637 (N_1637,N_442,N_230);
and U1638 (N_1638,N_211,N_105);
or U1639 (N_1639,N_558,N_326);
nand U1640 (N_1640,N_930,N_574);
nor U1641 (N_1641,N_93,N_131);
and U1642 (N_1642,N_755,N_346);
nor U1643 (N_1643,N_503,N_213);
and U1644 (N_1644,N_185,N_548);
nand U1645 (N_1645,N_174,N_704);
nand U1646 (N_1646,N_804,N_801);
or U1647 (N_1647,N_523,N_483);
and U1648 (N_1648,N_211,N_323);
or U1649 (N_1649,N_812,N_333);
nor U1650 (N_1650,N_751,N_142);
nand U1651 (N_1651,N_416,N_805);
nor U1652 (N_1652,N_218,N_767);
and U1653 (N_1653,N_295,N_311);
or U1654 (N_1654,N_535,N_199);
and U1655 (N_1655,N_152,N_587);
nor U1656 (N_1656,N_632,N_416);
nand U1657 (N_1657,N_978,N_812);
and U1658 (N_1658,N_464,N_90);
or U1659 (N_1659,N_719,N_138);
and U1660 (N_1660,N_350,N_604);
or U1661 (N_1661,N_402,N_378);
nor U1662 (N_1662,N_76,N_908);
or U1663 (N_1663,N_563,N_366);
and U1664 (N_1664,N_558,N_332);
and U1665 (N_1665,N_961,N_358);
or U1666 (N_1666,N_921,N_209);
or U1667 (N_1667,N_855,N_316);
and U1668 (N_1668,N_391,N_167);
nand U1669 (N_1669,N_798,N_214);
and U1670 (N_1670,N_741,N_836);
nand U1671 (N_1671,N_222,N_11);
nand U1672 (N_1672,N_968,N_955);
or U1673 (N_1673,N_16,N_244);
and U1674 (N_1674,N_240,N_967);
nor U1675 (N_1675,N_229,N_746);
nor U1676 (N_1676,N_37,N_377);
nor U1677 (N_1677,N_970,N_145);
nor U1678 (N_1678,N_583,N_116);
nand U1679 (N_1679,N_59,N_943);
or U1680 (N_1680,N_921,N_562);
nor U1681 (N_1681,N_704,N_175);
nand U1682 (N_1682,N_443,N_226);
nand U1683 (N_1683,N_417,N_613);
nor U1684 (N_1684,N_657,N_885);
or U1685 (N_1685,N_364,N_941);
xor U1686 (N_1686,N_712,N_726);
and U1687 (N_1687,N_622,N_607);
xor U1688 (N_1688,N_71,N_17);
nand U1689 (N_1689,N_13,N_204);
or U1690 (N_1690,N_989,N_586);
and U1691 (N_1691,N_697,N_642);
or U1692 (N_1692,N_337,N_577);
nor U1693 (N_1693,N_780,N_582);
or U1694 (N_1694,N_924,N_318);
xor U1695 (N_1695,N_827,N_184);
xor U1696 (N_1696,N_642,N_791);
nor U1697 (N_1697,N_925,N_614);
nor U1698 (N_1698,N_759,N_746);
and U1699 (N_1699,N_468,N_82);
nand U1700 (N_1700,N_46,N_823);
or U1701 (N_1701,N_125,N_147);
or U1702 (N_1702,N_691,N_414);
xor U1703 (N_1703,N_924,N_524);
or U1704 (N_1704,N_923,N_221);
and U1705 (N_1705,N_263,N_708);
nand U1706 (N_1706,N_724,N_784);
nand U1707 (N_1707,N_553,N_451);
nand U1708 (N_1708,N_939,N_377);
or U1709 (N_1709,N_867,N_789);
nor U1710 (N_1710,N_89,N_584);
or U1711 (N_1711,N_589,N_406);
or U1712 (N_1712,N_260,N_296);
and U1713 (N_1713,N_256,N_821);
and U1714 (N_1714,N_466,N_954);
nor U1715 (N_1715,N_455,N_748);
nand U1716 (N_1716,N_508,N_803);
xnor U1717 (N_1717,N_307,N_56);
nor U1718 (N_1718,N_535,N_908);
nor U1719 (N_1719,N_598,N_576);
nand U1720 (N_1720,N_942,N_576);
or U1721 (N_1721,N_360,N_791);
xnor U1722 (N_1722,N_211,N_72);
or U1723 (N_1723,N_684,N_856);
nand U1724 (N_1724,N_554,N_233);
xor U1725 (N_1725,N_143,N_973);
nand U1726 (N_1726,N_949,N_525);
and U1727 (N_1727,N_748,N_12);
or U1728 (N_1728,N_893,N_249);
xor U1729 (N_1729,N_196,N_66);
or U1730 (N_1730,N_729,N_652);
and U1731 (N_1731,N_769,N_353);
and U1732 (N_1732,N_980,N_468);
xor U1733 (N_1733,N_356,N_957);
nand U1734 (N_1734,N_550,N_891);
and U1735 (N_1735,N_834,N_126);
nor U1736 (N_1736,N_147,N_993);
nand U1737 (N_1737,N_15,N_956);
nor U1738 (N_1738,N_885,N_712);
nor U1739 (N_1739,N_794,N_992);
nor U1740 (N_1740,N_243,N_738);
nor U1741 (N_1741,N_763,N_510);
nand U1742 (N_1742,N_401,N_948);
nand U1743 (N_1743,N_515,N_924);
and U1744 (N_1744,N_258,N_888);
nand U1745 (N_1745,N_788,N_496);
and U1746 (N_1746,N_304,N_811);
nand U1747 (N_1747,N_982,N_219);
or U1748 (N_1748,N_253,N_123);
xnor U1749 (N_1749,N_553,N_696);
or U1750 (N_1750,N_109,N_300);
or U1751 (N_1751,N_3,N_758);
and U1752 (N_1752,N_739,N_937);
xnor U1753 (N_1753,N_318,N_678);
and U1754 (N_1754,N_5,N_645);
and U1755 (N_1755,N_589,N_178);
nor U1756 (N_1756,N_210,N_8);
xor U1757 (N_1757,N_40,N_698);
nand U1758 (N_1758,N_77,N_335);
or U1759 (N_1759,N_375,N_211);
nand U1760 (N_1760,N_120,N_714);
or U1761 (N_1761,N_985,N_24);
nor U1762 (N_1762,N_298,N_569);
nor U1763 (N_1763,N_306,N_895);
nor U1764 (N_1764,N_582,N_670);
and U1765 (N_1765,N_672,N_337);
and U1766 (N_1766,N_754,N_473);
and U1767 (N_1767,N_800,N_812);
and U1768 (N_1768,N_37,N_950);
nand U1769 (N_1769,N_156,N_429);
or U1770 (N_1770,N_986,N_865);
or U1771 (N_1771,N_188,N_730);
and U1772 (N_1772,N_815,N_245);
and U1773 (N_1773,N_622,N_982);
and U1774 (N_1774,N_66,N_958);
nand U1775 (N_1775,N_781,N_23);
nor U1776 (N_1776,N_426,N_34);
nor U1777 (N_1777,N_400,N_227);
or U1778 (N_1778,N_319,N_853);
xnor U1779 (N_1779,N_165,N_938);
and U1780 (N_1780,N_302,N_837);
or U1781 (N_1781,N_499,N_998);
nor U1782 (N_1782,N_198,N_166);
nand U1783 (N_1783,N_508,N_981);
nand U1784 (N_1784,N_246,N_941);
and U1785 (N_1785,N_777,N_293);
nand U1786 (N_1786,N_971,N_695);
nand U1787 (N_1787,N_831,N_763);
nor U1788 (N_1788,N_725,N_269);
and U1789 (N_1789,N_525,N_940);
and U1790 (N_1790,N_40,N_848);
xnor U1791 (N_1791,N_215,N_489);
xor U1792 (N_1792,N_712,N_956);
or U1793 (N_1793,N_844,N_69);
or U1794 (N_1794,N_362,N_950);
and U1795 (N_1795,N_953,N_459);
nor U1796 (N_1796,N_261,N_51);
and U1797 (N_1797,N_888,N_639);
nor U1798 (N_1798,N_589,N_190);
nor U1799 (N_1799,N_432,N_390);
or U1800 (N_1800,N_517,N_495);
xor U1801 (N_1801,N_423,N_530);
or U1802 (N_1802,N_498,N_845);
or U1803 (N_1803,N_798,N_300);
nand U1804 (N_1804,N_548,N_118);
or U1805 (N_1805,N_556,N_48);
or U1806 (N_1806,N_155,N_630);
nor U1807 (N_1807,N_936,N_812);
nand U1808 (N_1808,N_453,N_757);
nand U1809 (N_1809,N_193,N_891);
nor U1810 (N_1810,N_279,N_533);
or U1811 (N_1811,N_195,N_670);
or U1812 (N_1812,N_665,N_469);
nand U1813 (N_1813,N_854,N_820);
and U1814 (N_1814,N_26,N_895);
and U1815 (N_1815,N_930,N_998);
xnor U1816 (N_1816,N_847,N_307);
or U1817 (N_1817,N_741,N_155);
xor U1818 (N_1818,N_574,N_971);
and U1819 (N_1819,N_417,N_245);
or U1820 (N_1820,N_226,N_0);
or U1821 (N_1821,N_994,N_917);
and U1822 (N_1822,N_689,N_726);
and U1823 (N_1823,N_498,N_746);
or U1824 (N_1824,N_896,N_689);
or U1825 (N_1825,N_121,N_577);
nor U1826 (N_1826,N_864,N_690);
or U1827 (N_1827,N_923,N_452);
nand U1828 (N_1828,N_110,N_940);
nor U1829 (N_1829,N_422,N_725);
and U1830 (N_1830,N_418,N_734);
nor U1831 (N_1831,N_73,N_138);
nand U1832 (N_1832,N_999,N_91);
or U1833 (N_1833,N_510,N_394);
nor U1834 (N_1834,N_679,N_214);
and U1835 (N_1835,N_322,N_18);
nand U1836 (N_1836,N_707,N_4);
nand U1837 (N_1837,N_670,N_126);
nand U1838 (N_1838,N_216,N_9);
xor U1839 (N_1839,N_8,N_242);
nand U1840 (N_1840,N_225,N_41);
nor U1841 (N_1841,N_232,N_150);
nor U1842 (N_1842,N_294,N_385);
nor U1843 (N_1843,N_52,N_203);
nor U1844 (N_1844,N_87,N_6);
nor U1845 (N_1845,N_462,N_768);
or U1846 (N_1846,N_516,N_36);
nand U1847 (N_1847,N_357,N_796);
or U1848 (N_1848,N_871,N_976);
nor U1849 (N_1849,N_436,N_373);
nand U1850 (N_1850,N_748,N_336);
nand U1851 (N_1851,N_616,N_954);
xor U1852 (N_1852,N_768,N_629);
nor U1853 (N_1853,N_395,N_249);
nor U1854 (N_1854,N_810,N_875);
and U1855 (N_1855,N_486,N_914);
nor U1856 (N_1856,N_252,N_501);
and U1857 (N_1857,N_663,N_997);
and U1858 (N_1858,N_553,N_106);
or U1859 (N_1859,N_192,N_416);
and U1860 (N_1860,N_183,N_398);
and U1861 (N_1861,N_167,N_330);
nand U1862 (N_1862,N_839,N_657);
or U1863 (N_1863,N_205,N_708);
and U1864 (N_1864,N_389,N_977);
nand U1865 (N_1865,N_892,N_620);
and U1866 (N_1866,N_192,N_489);
xnor U1867 (N_1867,N_216,N_346);
nor U1868 (N_1868,N_331,N_468);
and U1869 (N_1869,N_590,N_971);
or U1870 (N_1870,N_149,N_723);
nor U1871 (N_1871,N_851,N_545);
nor U1872 (N_1872,N_722,N_524);
and U1873 (N_1873,N_26,N_187);
or U1874 (N_1874,N_597,N_827);
nand U1875 (N_1875,N_739,N_437);
nor U1876 (N_1876,N_78,N_592);
nor U1877 (N_1877,N_621,N_987);
nand U1878 (N_1878,N_733,N_23);
xor U1879 (N_1879,N_874,N_128);
nand U1880 (N_1880,N_407,N_421);
and U1881 (N_1881,N_892,N_863);
or U1882 (N_1882,N_438,N_492);
nand U1883 (N_1883,N_520,N_889);
nand U1884 (N_1884,N_370,N_50);
nor U1885 (N_1885,N_521,N_563);
nand U1886 (N_1886,N_984,N_859);
nor U1887 (N_1887,N_152,N_85);
or U1888 (N_1888,N_338,N_990);
and U1889 (N_1889,N_733,N_67);
nor U1890 (N_1890,N_375,N_493);
nor U1891 (N_1891,N_940,N_759);
nor U1892 (N_1892,N_297,N_4);
nor U1893 (N_1893,N_430,N_809);
nor U1894 (N_1894,N_711,N_579);
nand U1895 (N_1895,N_937,N_161);
nand U1896 (N_1896,N_886,N_343);
nor U1897 (N_1897,N_830,N_975);
or U1898 (N_1898,N_374,N_682);
xor U1899 (N_1899,N_252,N_783);
or U1900 (N_1900,N_127,N_405);
nor U1901 (N_1901,N_431,N_246);
or U1902 (N_1902,N_377,N_554);
and U1903 (N_1903,N_658,N_590);
or U1904 (N_1904,N_879,N_714);
xnor U1905 (N_1905,N_560,N_559);
nand U1906 (N_1906,N_35,N_939);
or U1907 (N_1907,N_318,N_559);
and U1908 (N_1908,N_365,N_596);
nand U1909 (N_1909,N_575,N_930);
nor U1910 (N_1910,N_925,N_495);
and U1911 (N_1911,N_562,N_604);
nand U1912 (N_1912,N_803,N_496);
nor U1913 (N_1913,N_585,N_396);
and U1914 (N_1914,N_979,N_314);
nor U1915 (N_1915,N_454,N_208);
nor U1916 (N_1916,N_681,N_450);
and U1917 (N_1917,N_995,N_466);
and U1918 (N_1918,N_262,N_817);
nor U1919 (N_1919,N_171,N_684);
nand U1920 (N_1920,N_510,N_39);
nor U1921 (N_1921,N_470,N_563);
and U1922 (N_1922,N_583,N_228);
and U1923 (N_1923,N_860,N_69);
and U1924 (N_1924,N_652,N_740);
or U1925 (N_1925,N_566,N_938);
nor U1926 (N_1926,N_583,N_786);
nor U1927 (N_1927,N_584,N_740);
nand U1928 (N_1928,N_653,N_880);
or U1929 (N_1929,N_714,N_607);
and U1930 (N_1930,N_782,N_184);
xor U1931 (N_1931,N_870,N_797);
and U1932 (N_1932,N_556,N_583);
or U1933 (N_1933,N_80,N_155);
and U1934 (N_1934,N_681,N_479);
or U1935 (N_1935,N_635,N_6);
nor U1936 (N_1936,N_836,N_460);
nor U1937 (N_1937,N_759,N_686);
or U1938 (N_1938,N_698,N_466);
and U1939 (N_1939,N_253,N_503);
xor U1940 (N_1940,N_266,N_375);
nor U1941 (N_1941,N_523,N_818);
or U1942 (N_1942,N_965,N_434);
and U1943 (N_1943,N_404,N_827);
or U1944 (N_1944,N_947,N_218);
or U1945 (N_1945,N_21,N_278);
or U1946 (N_1946,N_393,N_838);
nand U1947 (N_1947,N_522,N_556);
nand U1948 (N_1948,N_409,N_921);
nand U1949 (N_1949,N_522,N_114);
and U1950 (N_1950,N_157,N_342);
or U1951 (N_1951,N_987,N_846);
or U1952 (N_1952,N_386,N_470);
nand U1953 (N_1953,N_969,N_45);
nand U1954 (N_1954,N_489,N_336);
nand U1955 (N_1955,N_691,N_518);
or U1956 (N_1956,N_955,N_190);
or U1957 (N_1957,N_751,N_113);
and U1958 (N_1958,N_551,N_115);
xnor U1959 (N_1959,N_406,N_755);
xor U1960 (N_1960,N_112,N_144);
nand U1961 (N_1961,N_753,N_460);
nor U1962 (N_1962,N_880,N_884);
or U1963 (N_1963,N_136,N_926);
nor U1964 (N_1964,N_659,N_177);
xor U1965 (N_1965,N_612,N_734);
nand U1966 (N_1966,N_870,N_578);
or U1967 (N_1967,N_568,N_544);
xnor U1968 (N_1968,N_758,N_343);
nor U1969 (N_1969,N_727,N_25);
nand U1970 (N_1970,N_832,N_533);
and U1971 (N_1971,N_264,N_779);
or U1972 (N_1972,N_809,N_192);
xnor U1973 (N_1973,N_429,N_708);
or U1974 (N_1974,N_120,N_418);
nor U1975 (N_1975,N_70,N_772);
nor U1976 (N_1976,N_71,N_392);
and U1977 (N_1977,N_765,N_443);
and U1978 (N_1978,N_617,N_921);
or U1979 (N_1979,N_906,N_649);
nor U1980 (N_1980,N_772,N_14);
nand U1981 (N_1981,N_423,N_625);
or U1982 (N_1982,N_85,N_31);
nand U1983 (N_1983,N_970,N_360);
nor U1984 (N_1984,N_218,N_906);
xnor U1985 (N_1985,N_975,N_231);
or U1986 (N_1986,N_343,N_447);
or U1987 (N_1987,N_13,N_19);
and U1988 (N_1988,N_19,N_799);
or U1989 (N_1989,N_11,N_20);
or U1990 (N_1990,N_152,N_867);
and U1991 (N_1991,N_627,N_977);
nand U1992 (N_1992,N_361,N_680);
nand U1993 (N_1993,N_207,N_861);
xnor U1994 (N_1994,N_321,N_56);
nor U1995 (N_1995,N_262,N_273);
xor U1996 (N_1996,N_79,N_877);
or U1997 (N_1997,N_636,N_195);
nand U1998 (N_1998,N_697,N_91);
and U1999 (N_1999,N_70,N_939);
nor U2000 (N_2000,N_1390,N_1282);
and U2001 (N_2001,N_1264,N_1425);
nor U2002 (N_2002,N_1608,N_1977);
nor U2003 (N_2003,N_1424,N_1045);
and U2004 (N_2004,N_1937,N_1662);
or U2005 (N_2005,N_1094,N_1435);
or U2006 (N_2006,N_1923,N_1947);
nor U2007 (N_2007,N_1628,N_1349);
or U2008 (N_2008,N_1790,N_1604);
and U2009 (N_2009,N_1399,N_1489);
xor U2010 (N_2010,N_1456,N_1611);
and U2011 (N_2011,N_1183,N_1479);
and U2012 (N_2012,N_1524,N_1253);
nor U2013 (N_2013,N_1029,N_1108);
nor U2014 (N_2014,N_1088,N_1493);
nand U2015 (N_2015,N_1231,N_1246);
nor U2016 (N_2016,N_1685,N_1063);
or U2017 (N_2017,N_1076,N_1280);
nand U2018 (N_2018,N_1721,N_1695);
xnor U2019 (N_2019,N_1558,N_1196);
xnor U2020 (N_2020,N_1749,N_1211);
and U2021 (N_2021,N_1309,N_1383);
nand U2022 (N_2022,N_1776,N_1346);
or U2023 (N_2023,N_1237,N_1434);
xnor U2024 (N_2024,N_1563,N_1751);
nor U2025 (N_2025,N_1601,N_1925);
or U2026 (N_2026,N_1012,N_1199);
xnor U2027 (N_2027,N_1665,N_1117);
nor U2028 (N_2028,N_1921,N_1120);
or U2029 (N_2029,N_1321,N_1566);
nand U2030 (N_2030,N_1955,N_1328);
and U2031 (N_2031,N_1292,N_1711);
or U2032 (N_2032,N_1984,N_1463);
nand U2033 (N_2033,N_1946,N_1759);
xnor U2034 (N_2034,N_1418,N_1053);
and U2035 (N_2035,N_1836,N_1723);
nand U2036 (N_2036,N_1146,N_1016);
and U2037 (N_2037,N_1382,N_1296);
or U2038 (N_2038,N_1743,N_1506);
and U2039 (N_2039,N_1889,N_1103);
xor U2040 (N_2040,N_1884,N_1326);
nand U2041 (N_2041,N_1518,N_1672);
nor U2042 (N_2042,N_1366,N_1896);
and U2043 (N_2043,N_1763,N_1397);
and U2044 (N_2044,N_1811,N_1165);
and U2045 (N_2045,N_1444,N_1141);
nor U2046 (N_2046,N_1930,N_1359);
nand U2047 (N_2047,N_1861,N_1215);
nand U2048 (N_2048,N_1090,N_1993);
nor U2049 (N_2049,N_1394,N_1371);
nand U2050 (N_2050,N_1426,N_1293);
nor U2051 (N_2051,N_1143,N_1501);
nand U2052 (N_2052,N_1013,N_1275);
and U2053 (N_2053,N_1976,N_1970);
nor U2054 (N_2054,N_1138,N_1148);
and U2055 (N_2055,N_1529,N_1269);
nor U2056 (N_2056,N_1173,N_1107);
xor U2057 (N_2057,N_1065,N_1846);
nand U2058 (N_2058,N_1755,N_1786);
or U2059 (N_2059,N_1168,N_1335);
or U2060 (N_2060,N_1431,N_1548);
xor U2061 (N_2061,N_1803,N_1830);
nor U2062 (N_2062,N_1322,N_1297);
or U2063 (N_2063,N_1163,N_1824);
nor U2064 (N_2064,N_1879,N_1208);
or U2065 (N_2065,N_1017,N_1433);
xnor U2066 (N_2066,N_1066,N_1051);
nor U2067 (N_2067,N_1754,N_1391);
nand U2068 (N_2068,N_1762,N_1298);
nor U2069 (N_2069,N_1202,N_1974);
nor U2070 (N_2070,N_1235,N_1500);
nor U2071 (N_2071,N_1182,N_1184);
xnor U2072 (N_2072,N_1841,N_1942);
nor U2073 (N_2073,N_1207,N_1798);
xor U2074 (N_2074,N_1064,N_1758);
or U2075 (N_2075,N_1516,N_1174);
nor U2076 (N_2076,N_1089,N_1586);
nand U2077 (N_2077,N_1416,N_1134);
or U2078 (N_2078,N_1155,N_1238);
and U2079 (N_2079,N_1589,N_1847);
nand U2080 (N_2080,N_1071,N_1839);
or U2081 (N_2081,N_1655,N_1689);
and U2082 (N_2082,N_1048,N_1052);
and U2083 (N_2083,N_1285,N_1927);
and U2084 (N_2084,N_1592,N_1599);
nand U2085 (N_2085,N_1475,N_1440);
or U2086 (N_2086,N_1062,N_1580);
nor U2087 (N_2087,N_1307,N_1883);
and U2088 (N_2088,N_1800,N_1964);
nand U2089 (N_2089,N_1512,N_1791);
nand U2090 (N_2090,N_1818,N_1538);
nand U2091 (N_2091,N_1209,N_1018);
or U2092 (N_2092,N_1697,N_1423);
and U2093 (N_2093,N_1442,N_1405);
nor U2094 (N_2094,N_1775,N_1810);
xnor U2095 (N_2095,N_1644,N_1642);
and U2096 (N_2096,N_1498,N_1272);
and U2097 (N_2097,N_1669,N_1733);
xor U2098 (N_2098,N_1649,N_1631);
nor U2099 (N_2099,N_1746,N_1240);
or U2100 (N_2100,N_1428,N_1951);
nor U2101 (N_2101,N_1850,N_1877);
xor U2102 (N_2102,N_1083,N_1505);
nor U2103 (N_2103,N_1038,N_1792);
nor U2104 (N_2104,N_1948,N_1194);
or U2105 (N_2105,N_1645,N_1115);
or U2106 (N_2106,N_1230,N_1190);
or U2107 (N_2107,N_1429,N_1907);
nand U2108 (N_2108,N_1187,N_1136);
nand U2109 (N_2109,N_1975,N_1254);
and U2110 (N_2110,N_1369,N_1717);
xnor U2111 (N_2111,N_1300,N_1871);
nor U2112 (N_2112,N_1157,N_1815);
nand U2113 (N_2113,N_1351,N_1314);
xor U2114 (N_2114,N_1806,N_1073);
nor U2115 (N_2115,N_1583,N_1849);
nand U2116 (N_2116,N_1398,N_1514);
and U2117 (N_2117,N_1989,N_1992);
nand U2118 (N_2118,N_1794,N_1259);
and U2119 (N_2119,N_1195,N_1125);
and U2120 (N_2120,N_1893,N_1613);
nor U2121 (N_2121,N_1482,N_1284);
nor U2122 (N_2122,N_1354,N_1761);
and U2123 (N_2123,N_1510,N_1378);
or U2124 (N_2124,N_1783,N_1778);
or U2125 (N_2125,N_1149,N_1327);
and U2126 (N_2126,N_1216,N_1312);
and U2127 (N_2127,N_1342,N_1526);
xor U2128 (N_2128,N_1823,N_1166);
nand U2129 (N_2129,N_1439,N_1311);
and U2130 (N_2130,N_1279,N_1922);
nand U2131 (N_2131,N_1971,N_1099);
and U2132 (N_2132,N_1543,N_1600);
and U2133 (N_2133,N_1480,N_1820);
nand U2134 (N_2134,N_1213,N_1039);
xnor U2135 (N_2135,N_1318,N_1863);
nand U2136 (N_2136,N_1987,N_1736);
nand U2137 (N_2137,N_1283,N_1528);
nand U2138 (N_2138,N_1161,N_1044);
and U2139 (N_2139,N_1464,N_1109);
or U2140 (N_2140,N_1513,N_1263);
nand U2141 (N_2141,N_1688,N_1453);
and U2142 (N_2142,N_1966,N_1504);
xnor U2143 (N_2143,N_1097,N_1178);
nor U2144 (N_2144,N_1034,N_1875);
xor U2145 (N_2145,N_1236,N_1119);
nand U2146 (N_2146,N_1005,N_1793);
or U2147 (N_2147,N_1324,N_1706);
or U2148 (N_2148,N_1415,N_1188);
xor U2149 (N_2149,N_1028,N_1882);
and U2150 (N_2150,N_1919,N_1805);
nand U2151 (N_2151,N_1363,N_1986);
nand U2152 (N_2152,N_1549,N_1234);
and U2153 (N_2153,N_1021,N_1782);
xor U2154 (N_2154,N_1625,N_1539);
nand U2155 (N_2155,N_1481,N_1059);
and U2156 (N_2156,N_1734,N_1286);
nand U2157 (N_2157,N_1694,N_1200);
and U2158 (N_2158,N_1036,N_1486);
and U2159 (N_2159,N_1870,N_1671);
nor U2160 (N_2160,N_1308,N_1130);
or U2161 (N_2161,N_1602,N_1931);
nand U2162 (N_2162,N_1040,N_1670);
nor U2163 (N_2163,N_1509,N_1079);
nand U2164 (N_2164,N_1336,N_1057);
or U2165 (N_2165,N_1080,N_1816);
nand U2166 (N_2166,N_1630,N_1325);
and U2167 (N_2167,N_1700,N_1864);
nor U2168 (N_2168,N_1680,N_1522);
nor U2169 (N_2169,N_1068,N_1180);
nor U2170 (N_2170,N_1595,N_1361);
or U2171 (N_2171,N_1027,N_1340);
nand U2172 (N_2172,N_1641,N_1111);
or U2173 (N_2173,N_1449,N_1347);
or U2174 (N_2174,N_1997,N_1807);
and U2175 (N_2175,N_1020,N_1888);
nand U2176 (N_2176,N_1570,N_1619);
xnor U2177 (N_2177,N_1056,N_1606);
nor U2178 (N_2178,N_1446,N_1898);
or U2179 (N_2179,N_1709,N_1329);
nor U2180 (N_2180,N_1193,N_1467);
nor U2181 (N_2181,N_1705,N_1210);
nor U2182 (N_2182,N_1677,N_1637);
nand U2183 (N_2183,N_1627,N_1544);
nand U2184 (N_2184,N_1960,N_1724);
or U2185 (N_2185,N_1855,N_1095);
nand U2186 (N_2186,N_1781,N_1904);
and U2187 (N_2187,N_1462,N_1160);
nand U2188 (N_2188,N_1962,N_1487);
and U2189 (N_2189,N_1978,N_1353);
and U2190 (N_2190,N_1164,N_1069);
nand U2191 (N_2191,N_1963,N_1437);
and U2192 (N_2192,N_1281,N_1933);
xnor U2193 (N_2193,N_1100,N_1750);
and U2194 (N_2194,N_1273,N_1058);
or U2195 (N_2195,N_1646,N_1972);
and U2196 (N_2196,N_1114,N_1417);
nand U2197 (N_2197,N_1535,N_1935);
xnor U2198 (N_2198,N_1133,N_1873);
nand U2199 (N_2199,N_1204,N_1660);
or U2200 (N_2200,N_1511,N_1084);
or U2201 (N_2201,N_1690,N_1085);
nand U2202 (N_2202,N_1448,N_1014);
nand U2203 (N_2203,N_1317,N_1176);
nand U2204 (N_2204,N_1345,N_1490);
nor U2205 (N_2205,N_1373,N_1222);
or U2206 (N_2206,N_1961,N_1306);
nand U2207 (N_2207,N_1334,N_1332);
or U2208 (N_2208,N_1362,N_1344);
nor U2209 (N_2209,N_1075,N_1077);
or U2210 (N_2210,N_1086,N_1722);
nor U2211 (N_2211,N_1192,N_1268);
xnor U2212 (N_2212,N_1607,N_1980);
nand U2213 (N_2213,N_1954,N_1031);
and U2214 (N_2214,N_1965,N_1532);
nor U2215 (N_2215,N_1145,N_1559);
nor U2216 (N_2216,N_1620,N_1092);
xnor U2217 (N_2217,N_1742,N_1945);
nor U2218 (N_2218,N_1692,N_1507);
nand U2219 (N_2219,N_1226,N_1828);
nand U2220 (N_2220,N_1414,N_1981);
or U2221 (N_2221,N_1147,N_1007);
nand U2222 (N_2222,N_1170,N_1227);
and U2223 (N_2223,N_1900,N_1957);
and U2224 (N_2224,N_1205,N_1728);
and U2225 (N_2225,N_1305,N_1666);
xnor U2226 (N_2226,N_1768,N_1396);
xor U2227 (N_2227,N_1508,N_1973);
nor U2228 (N_2228,N_1153,N_1001);
or U2229 (N_2229,N_1203,N_1358);
and U2230 (N_2230,N_1116,N_1523);
and U2231 (N_2231,N_1386,N_1869);
or U2232 (N_2232,N_1410,N_1406);
nand U2233 (N_2233,N_1003,N_1185);
nand U2234 (N_2234,N_1780,N_1659);
and U2235 (N_2235,N_1616,N_1653);
and U2236 (N_2236,N_1252,N_1047);
and U2237 (N_2237,N_1740,N_1719);
and U2238 (N_2238,N_1458,N_1531);
and U2239 (N_2239,N_1880,N_1579);
or U2240 (N_2240,N_1872,N_1530);
nand U2241 (N_2241,N_1679,N_1663);
and U2242 (N_2242,N_1181,N_1023);
or U2243 (N_2243,N_1537,N_1339);
nand U2244 (N_2244,N_1113,N_1019);
nand U2245 (N_2245,N_1212,N_1476);
nor U2246 (N_2246,N_1419,N_1137);
and U2247 (N_2247,N_1995,N_1858);
or U2248 (N_2248,N_1123,N_1255);
or U2249 (N_2249,N_1802,N_1998);
or U2250 (N_2250,N_1096,N_1191);
xor U2251 (N_2251,N_1771,N_1162);
nor U2252 (N_2252,N_1796,N_1647);
or U2253 (N_2253,N_1030,N_1129);
or U2254 (N_2254,N_1367,N_1867);
or U2255 (N_2255,N_1443,N_1310);
and U2256 (N_2256,N_1067,N_1242);
nor U2257 (N_2257,N_1699,N_1233);
nor U2258 (N_2258,N_1801,N_1936);
xor U2259 (N_2259,N_1395,N_1035);
xor U2260 (N_2260,N_1996,N_1049);
and U2261 (N_2261,N_1959,N_1503);
and U2262 (N_2262,N_1704,N_1009);
xor U2263 (N_2263,N_1590,N_1206);
nand U2264 (N_2264,N_1172,N_1375);
nor U2265 (N_2265,N_1767,N_1251);
or U2266 (N_2266,N_1897,N_1041);
nor U2267 (N_2267,N_1929,N_1545);
and U2268 (N_2268,N_1152,N_1906);
nor U2269 (N_2269,N_1288,N_1569);
nand U2270 (N_2270,N_1257,N_1320);
or U2271 (N_2271,N_1471,N_1054);
nor U2272 (N_2272,N_1261,N_1266);
or U2273 (N_2273,N_1624,N_1789);
or U2274 (N_2274,N_1638,N_1409);
or U2275 (N_2275,N_1495,N_1577);
or U2276 (N_2276,N_1000,N_1492);
or U2277 (N_2277,N_1720,N_1105);
and U2278 (N_2278,N_1228,N_1832);
and U2279 (N_2279,N_1276,N_1814);
nand U2280 (N_2280,N_1400,N_1248);
and U2281 (N_2281,N_1004,N_1142);
xor U2282 (N_2282,N_1756,N_1333);
nor U2283 (N_2283,N_1393,N_1729);
or U2284 (N_2284,N_1716,N_1725);
nor U2285 (N_2285,N_1247,N_1702);
nand U2286 (N_2286,N_1676,N_1681);
or U2287 (N_2287,N_1483,N_1411);
nor U2288 (N_2288,N_1615,N_1967);
or U2289 (N_2289,N_1744,N_1301);
nand U2290 (N_2290,N_1278,N_1784);
nand U2291 (N_2291,N_1478,N_1675);
nand U2292 (N_2292,N_1407,N_1737);
xor U2293 (N_2293,N_1330,N_1703);
nor U2294 (N_2294,N_1696,N_1932);
or U2295 (N_2295,N_1988,N_1732);
nor U2296 (N_2296,N_1905,N_1886);
or U2297 (N_2297,N_1427,N_1229);
nor U2298 (N_2298,N_1150,N_1909);
or U2299 (N_2299,N_1132,N_1348);
xnor U2300 (N_2300,N_1691,N_1106);
xor U2301 (N_2301,N_1256,N_1916);
nand U2302 (N_2302,N_1693,N_1555);
nand U2303 (N_2303,N_1868,N_1316);
nand U2304 (N_2304,N_1885,N_1926);
and U2305 (N_2305,N_1037,N_1707);
nor U2306 (N_2306,N_1892,N_1451);
or U2307 (N_2307,N_1454,N_1837);
nand U2308 (N_2308,N_1629,N_1878);
or U2309 (N_2309,N_1668,N_1384);
or U2310 (N_2310,N_1623,N_1661);
xor U2311 (N_2311,N_1343,N_1422);
and U2312 (N_2312,N_1682,N_1924);
and U2313 (N_2313,N_1060,N_1730);
nand U2314 (N_2314,N_1969,N_1785);
nand U2315 (N_2315,N_1745,N_1573);
and U2316 (N_2316,N_1860,N_1817);
and U2317 (N_2317,N_1812,N_1835);
and U2318 (N_2318,N_1777,N_1774);
or U2319 (N_2319,N_1943,N_1757);
nand U2320 (N_2320,N_1990,N_1770);
or U2321 (N_2321,N_1122,N_1154);
and U2322 (N_2322,N_1657,N_1773);
and U2323 (N_2323,N_1968,N_1502);
xor U2324 (N_2324,N_1712,N_1603);
nor U2325 (N_2325,N_1683,N_1748);
or U2326 (N_2326,N_1026,N_1684);
nand U2327 (N_2327,N_1982,N_1686);
or U2328 (N_2328,N_1587,N_1144);
or U2329 (N_2329,N_1169,N_1739);
or U2330 (N_2330,N_1295,N_1852);
nor U2331 (N_2331,N_1714,N_1118);
and U2332 (N_2332,N_1460,N_1357);
and U2333 (N_2333,N_1760,N_1825);
and U2334 (N_2334,N_1158,N_1258);
nor U2335 (N_2335,N_1956,N_1618);
and U2336 (N_2336,N_1547,N_1643);
and U2337 (N_2337,N_1940,N_1403);
xnor U2338 (N_2338,N_1465,N_1626);
xnor U2339 (N_2339,N_1379,N_1331);
nor U2340 (N_2340,N_1614,N_1302);
nand U2341 (N_2341,N_1452,N_1766);
and U2342 (N_2342,N_1635,N_1186);
nand U2343 (N_2343,N_1198,N_1387);
and U2344 (N_2344,N_1466,N_1214);
or U2345 (N_2345,N_1651,N_1859);
nor U2346 (N_2346,N_1389,N_1177);
nand U2347 (N_2347,N_1159,N_1833);
and U2348 (N_2348,N_1043,N_1572);
or U2349 (N_2349,N_1584,N_1912);
and U2350 (N_2350,N_1673,N_1370);
xnor U2351 (N_2351,N_1491,N_1474);
nand U2352 (N_2352,N_1350,N_1365);
or U2353 (N_2353,N_1779,N_1441);
and U2354 (N_2354,N_1032,N_1609);
or U2355 (N_2355,N_1552,N_1102);
or U2356 (N_2356,N_1376,N_1827);
or U2357 (N_2357,N_1715,N_1808);
nor U2358 (N_2358,N_1593,N_1854);
or U2359 (N_2359,N_1313,N_1455);
and U2360 (N_2360,N_1461,N_1135);
nor U2361 (N_2361,N_1845,N_1171);
xor U2362 (N_2362,N_1112,N_1110);
nand U2363 (N_2363,N_1804,N_1050);
nand U2364 (N_2364,N_1542,N_1950);
or U2365 (N_2365,N_1033,N_1006);
and U2366 (N_2366,N_1352,N_1388);
and U2367 (N_2367,N_1949,N_1450);
nor U2368 (N_2368,N_1477,N_1617);
or U2369 (N_2369,N_1323,N_1941);
nand U2370 (N_2370,N_1876,N_1903);
nor U2371 (N_2371,N_1179,N_1223);
nand U2372 (N_2372,N_1519,N_1560);
or U2373 (N_2373,N_1843,N_1219);
nand U2374 (N_2374,N_1561,N_1087);
xnor U2375 (N_2375,N_1291,N_1999);
nor U2376 (N_2376,N_1726,N_1844);
and U2377 (N_2377,N_1011,N_1622);
or U2378 (N_2378,N_1913,N_1533);
xor U2379 (N_2379,N_1656,N_1727);
nor U2380 (N_2380,N_1612,N_1874);
nor U2381 (N_2381,N_1738,N_1380);
or U2382 (N_2382,N_1866,N_1022);
or U2383 (N_2383,N_1270,N_1408);
nand U2384 (N_2384,N_1232,N_1081);
nand U2385 (N_2385,N_1404,N_1632);
nor U2386 (N_2386,N_1597,N_1652);
nor U2387 (N_2387,N_1472,N_1834);
nand U2388 (N_2388,N_1224,N_1731);
or U2389 (N_2389,N_1862,N_1819);
xor U2390 (N_2390,N_1008,N_1315);
nand U2391 (N_2391,N_1540,N_1356);
or U2392 (N_2392,N_1797,N_1848);
nor U2393 (N_2393,N_1753,N_1290);
or U2394 (N_2394,N_1708,N_1564);
nand U2395 (N_2395,N_1024,N_1851);
nand U2396 (N_2396,N_1459,N_1582);
xnor U2397 (N_2397,N_1091,N_1918);
and U2398 (N_2398,N_1430,N_1260);
nand U2399 (N_2399,N_1287,N_1074);
and U2400 (N_2400,N_1574,N_1127);
xnor U2401 (N_2401,N_1250,N_1217);
nor U2402 (N_2402,N_1241,N_1497);
nand U2403 (N_2403,N_1636,N_1894);
and U2404 (N_2404,N_1496,N_1055);
or U2405 (N_2405,N_1197,N_1289);
or U2406 (N_2406,N_1741,N_1294);
nor U2407 (N_2407,N_1985,N_1385);
or U2408 (N_2408,N_1994,N_1550);
and U2409 (N_2409,N_1436,N_1902);
nor U2410 (N_2410,N_1591,N_1713);
nand U2411 (N_2411,N_1674,N_1856);
nor U2412 (N_2412,N_1557,N_1262);
xor U2413 (N_2413,N_1765,N_1402);
nand U2414 (N_2414,N_1881,N_1840);
and U2415 (N_2415,N_1917,N_1274);
nand U2416 (N_2416,N_1447,N_1072);
nor U2417 (N_2417,N_1788,N_1101);
or U2418 (N_2418,N_1887,N_1596);
xor U2419 (N_2419,N_1920,N_1139);
and U2420 (N_2420,N_1381,N_1556);
nand U2421 (N_2421,N_1319,N_1244);
xor U2422 (N_2422,N_1710,N_1928);
and U2423 (N_2423,N_1664,N_1910);
nor U2424 (N_2424,N_1245,N_1438);
and U2425 (N_2425,N_1658,N_1842);
nand U2426 (N_2426,N_1140,N_1991);
xnor U2427 (N_2427,N_1372,N_1243);
and U2428 (N_2428,N_1764,N_1831);
and U2429 (N_2429,N_1915,N_1594);
xor U2430 (N_2430,N_1585,N_1128);
or U2431 (N_2431,N_1747,N_1412);
and U2432 (N_2432,N_1581,N_1553);
nor U2433 (N_2433,N_1121,N_1979);
or U2434 (N_2434,N_1271,N_1473);
xor U2435 (N_2435,N_1265,N_1799);
and U2436 (N_2436,N_1826,N_1953);
and U2437 (N_2437,N_1485,N_1249);
and U2438 (N_2438,N_1795,N_1061);
nand U2439 (N_2439,N_1025,N_1838);
nand U2440 (N_2440,N_1401,N_1698);
nor U2441 (N_2441,N_1654,N_1648);
nand U2442 (N_2442,N_1634,N_1901);
or U2443 (N_2443,N_1908,N_1527);
nor U2444 (N_2444,N_1070,N_1639);
and U2445 (N_2445,N_1914,N_1131);
or U2446 (N_2446,N_1221,N_1650);
nor U2447 (N_2447,N_1857,N_1568);
nor U2448 (N_2448,N_1678,N_1534);
or U2449 (N_2449,N_1126,N_1718);
or U2450 (N_2450,N_1983,N_1470);
xnor U2451 (N_2451,N_1239,N_1341);
and U2452 (N_2452,N_1640,N_1360);
and U2453 (N_2453,N_1822,N_1277);
or U2454 (N_2454,N_1633,N_1218);
xnor U2455 (N_2455,N_1899,N_1010);
and U2456 (N_2456,N_1167,N_1895);
nor U2457 (N_2457,N_1042,N_1488);
nand U2458 (N_2458,N_1605,N_1787);
nand U2459 (N_2459,N_1220,N_1078);
xnor U2460 (N_2460,N_1338,N_1104);
or U2461 (N_2461,N_1562,N_1494);
or U2462 (N_2462,N_1201,N_1457);
nand U2463 (N_2463,N_1934,N_1364);
and U2464 (N_2464,N_1469,N_1420);
and U2465 (N_2465,N_1701,N_1355);
nand U2466 (N_2466,N_1575,N_1939);
xor U2467 (N_2467,N_1829,N_1541);
or U2468 (N_2468,N_1156,N_1952);
nor U2469 (N_2469,N_1944,N_1865);
or U2470 (N_2470,N_1304,N_1392);
and U2471 (N_2471,N_1938,N_1890);
nor U2472 (N_2472,N_1571,N_1175);
nand U2473 (N_2473,N_1082,N_1413);
nor U2474 (N_2474,N_1588,N_1267);
and U2475 (N_2475,N_1667,N_1567);
or U2476 (N_2476,N_1621,N_1551);
nand U2477 (N_2477,N_1520,N_1687);
nand U2478 (N_2478,N_1735,N_1445);
nor U2479 (N_2479,N_1772,N_1525);
and U2480 (N_2480,N_1303,N_1752);
nor U2481 (N_2481,N_1377,N_1521);
nand U2482 (N_2482,N_1093,N_1546);
nand U2483 (N_2483,N_1610,N_1911);
xnor U2484 (N_2484,N_1299,N_1499);
nor U2485 (N_2485,N_1536,N_1225);
nor U2486 (N_2486,N_1515,N_1432);
and U2487 (N_2487,N_1554,N_1598);
xnor U2488 (N_2488,N_1368,N_1769);
nor U2489 (N_2489,N_1002,N_1813);
and U2490 (N_2490,N_1337,N_1484);
nand U2491 (N_2491,N_1189,N_1468);
xnor U2492 (N_2492,N_1421,N_1046);
and U2493 (N_2493,N_1374,N_1576);
nand U2494 (N_2494,N_1891,N_1853);
or U2495 (N_2495,N_1565,N_1821);
xor U2496 (N_2496,N_1151,N_1015);
nand U2497 (N_2497,N_1124,N_1809);
xor U2498 (N_2498,N_1098,N_1958);
xor U2499 (N_2499,N_1578,N_1517);
or U2500 (N_2500,N_1147,N_1246);
nand U2501 (N_2501,N_1730,N_1843);
and U2502 (N_2502,N_1010,N_1122);
and U2503 (N_2503,N_1371,N_1021);
xnor U2504 (N_2504,N_1866,N_1798);
xor U2505 (N_2505,N_1873,N_1307);
and U2506 (N_2506,N_1607,N_1149);
and U2507 (N_2507,N_1204,N_1189);
nand U2508 (N_2508,N_1828,N_1935);
nand U2509 (N_2509,N_1609,N_1488);
and U2510 (N_2510,N_1908,N_1409);
nand U2511 (N_2511,N_1208,N_1735);
xnor U2512 (N_2512,N_1139,N_1668);
or U2513 (N_2513,N_1216,N_1840);
or U2514 (N_2514,N_1622,N_1157);
nor U2515 (N_2515,N_1848,N_1416);
nand U2516 (N_2516,N_1547,N_1015);
or U2517 (N_2517,N_1543,N_1910);
or U2518 (N_2518,N_1705,N_1632);
nand U2519 (N_2519,N_1217,N_1152);
nand U2520 (N_2520,N_1763,N_1062);
and U2521 (N_2521,N_1575,N_1665);
and U2522 (N_2522,N_1846,N_1223);
nand U2523 (N_2523,N_1411,N_1547);
and U2524 (N_2524,N_1266,N_1115);
nor U2525 (N_2525,N_1178,N_1355);
nand U2526 (N_2526,N_1185,N_1863);
and U2527 (N_2527,N_1719,N_1417);
or U2528 (N_2528,N_1901,N_1418);
or U2529 (N_2529,N_1911,N_1284);
or U2530 (N_2530,N_1545,N_1028);
nand U2531 (N_2531,N_1622,N_1252);
and U2532 (N_2532,N_1049,N_1221);
and U2533 (N_2533,N_1498,N_1722);
and U2534 (N_2534,N_1748,N_1068);
nand U2535 (N_2535,N_1185,N_1290);
nand U2536 (N_2536,N_1378,N_1415);
and U2537 (N_2537,N_1237,N_1347);
nand U2538 (N_2538,N_1018,N_1914);
or U2539 (N_2539,N_1167,N_1956);
or U2540 (N_2540,N_1812,N_1731);
nor U2541 (N_2541,N_1700,N_1292);
nor U2542 (N_2542,N_1626,N_1705);
or U2543 (N_2543,N_1033,N_1212);
nor U2544 (N_2544,N_1392,N_1855);
nand U2545 (N_2545,N_1117,N_1014);
nor U2546 (N_2546,N_1074,N_1122);
xor U2547 (N_2547,N_1360,N_1470);
and U2548 (N_2548,N_1067,N_1406);
and U2549 (N_2549,N_1681,N_1227);
and U2550 (N_2550,N_1776,N_1351);
or U2551 (N_2551,N_1465,N_1533);
nor U2552 (N_2552,N_1353,N_1473);
nor U2553 (N_2553,N_1728,N_1845);
xor U2554 (N_2554,N_1662,N_1154);
nand U2555 (N_2555,N_1442,N_1321);
and U2556 (N_2556,N_1606,N_1146);
and U2557 (N_2557,N_1215,N_1968);
and U2558 (N_2558,N_1185,N_1774);
and U2559 (N_2559,N_1545,N_1621);
nand U2560 (N_2560,N_1418,N_1373);
nor U2561 (N_2561,N_1674,N_1980);
and U2562 (N_2562,N_1426,N_1748);
nor U2563 (N_2563,N_1984,N_1080);
nor U2564 (N_2564,N_1893,N_1709);
or U2565 (N_2565,N_1012,N_1594);
or U2566 (N_2566,N_1003,N_1285);
nand U2567 (N_2567,N_1273,N_1559);
and U2568 (N_2568,N_1916,N_1701);
and U2569 (N_2569,N_1463,N_1302);
or U2570 (N_2570,N_1001,N_1454);
and U2571 (N_2571,N_1787,N_1437);
and U2572 (N_2572,N_1177,N_1344);
nor U2573 (N_2573,N_1176,N_1510);
or U2574 (N_2574,N_1469,N_1551);
xnor U2575 (N_2575,N_1823,N_1107);
xor U2576 (N_2576,N_1468,N_1497);
or U2577 (N_2577,N_1622,N_1682);
nor U2578 (N_2578,N_1141,N_1655);
and U2579 (N_2579,N_1050,N_1473);
and U2580 (N_2580,N_1948,N_1432);
nor U2581 (N_2581,N_1117,N_1196);
or U2582 (N_2582,N_1706,N_1208);
and U2583 (N_2583,N_1113,N_1923);
nor U2584 (N_2584,N_1057,N_1200);
nand U2585 (N_2585,N_1857,N_1082);
or U2586 (N_2586,N_1154,N_1617);
nand U2587 (N_2587,N_1830,N_1905);
nand U2588 (N_2588,N_1269,N_1263);
nor U2589 (N_2589,N_1463,N_1499);
nor U2590 (N_2590,N_1382,N_1039);
or U2591 (N_2591,N_1834,N_1955);
and U2592 (N_2592,N_1156,N_1846);
or U2593 (N_2593,N_1414,N_1253);
or U2594 (N_2594,N_1337,N_1189);
or U2595 (N_2595,N_1147,N_1238);
or U2596 (N_2596,N_1643,N_1541);
and U2597 (N_2597,N_1363,N_1435);
nand U2598 (N_2598,N_1987,N_1357);
and U2599 (N_2599,N_1605,N_1407);
nand U2600 (N_2600,N_1193,N_1572);
nand U2601 (N_2601,N_1992,N_1240);
and U2602 (N_2602,N_1815,N_1656);
xor U2603 (N_2603,N_1101,N_1413);
nand U2604 (N_2604,N_1076,N_1488);
and U2605 (N_2605,N_1050,N_1824);
nand U2606 (N_2606,N_1250,N_1602);
and U2607 (N_2607,N_1546,N_1191);
xor U2608 (N_2608,N_1336,N_1478);
nand U2609 (N_2609,N_1191,N_1468);
nand U2610 (N_2610,N_1534,N_1061);
and U2611 (N_2611,N_1609,N_1886);
nor U2612 (N_2612,N_1661,N_1553);
and U2613 (N_2613,N_1466,N_1699);
xnor U2614 (N_2614,N_1091,N_1627);
nor U2615 (N_2615,N_1484,N_1004);
and U2616 (N_2616,N_1574,N_1722);
or U2617 (N_2617,N_1679,N_1434);
nor U2618 (N_2618,N_1120,N_1272);
nand U2619 (N_2619,N_1781,N_1248);
nand U2620 (N_2620,N_1070,N_1493);
xnor U2621 (N_2621,N_1296,N_1115);
nand U2622 (N_2622,N_1864,N_1654);
nand U2623 (N_2623,N_1835,N_1958);
nor U2624 (N_2624,N_1102,N_1441);
nor U2625 (N_2625,N_1738,N_1378);
and U2626 (N_2626,N_1316,N_1413);
and U2627 (N_2627,N_1571,N_1337);
and U2628 (N_2628,N_1591,N_1071);
nor U2629 (N_2629,N_1229,N_1934);
nand U2630 (N_2630,N_1343,N_1880);
nand U2631 (N_2631,N_1280,N_1418);
and U2632 (N_2632,N_1079,N_1382);
xnor U2633 (N_2633,N_1521,N_1321);
xor U2634 (N_2634,N_1151,N_1741);
nor U2635 (N_2635,N_1605,N_1537);
nor U2636 (N_2636,N_1237,N_1896);
or U2637 (N_2637,N_1007,N_1314);
xnor U2638 (N_2638,N_1929,N_1254);
nand U2639 (N_2639,N_1122,N_1515);
nand U2640 (N_2640,N_1249,N_1975);
and U2641 (N_2641,N_1648,N_1139);
or U2642 (N_2642,N_1328,N_1930);
nand U2643 (N_2643,N_1404,N_1715);
xnor U2644 (N_2644,N_1936,N_1397);
or U2645 (N_2645,N_1783,N_1498);
xor U2646 (N_2646,N_1692,N_1107);
or U2647 (N_2647,N_1230,N_1687);
and U2648 (N_2648,N_1735,N_1632);
nor U2649 (N_2649,N_1010,N_1057);
or U2650 (N_2650,N_1173,N_1720);
nor U2651 (N_2651,N_1452,N_1239);
xnor U2652 (N_2652,N_1472,N_1722);
and U2653 (N_2653,N_1450,N_1854);
or U2654 (N_2654,N_1272,N_1001);
xnor U2655 (N_2655,N_1914,N_1383);
and U2656 (N_2656,N_1615,N_1498);
nand U2657 (N_2657,N_1755,N_1586);
and U2658 (N_2658,N_1751,N_1664);
xnor U2659 (N_2659,N_1289,N_1296);
nand U2660 (N_2660,N_1156,N_1622);
and U2661 (N_2661,N_1534,N_1844);
and U2662 (N_2662,N_1304,N_1131);
or U2663 (N_2663,N_1893,N_1240);
and U2664 (N_2664,N_1316,N_1595);
xor U2665 (N_2665,N_1652,N_1844);
nor U2666 (N_2666,N_1239,N_1276);
xor U2667 (N_2667,N_1759,N_1281);
nand U2668 (N_2668,N_1676,N_1863);
and U2669 (N_2669,N_1533,N_1170);
nand U2670 (N_2670,N_1172,N_1043);
and U2671 (N_2671,N_1913,N_1179);
and U2672 (N_2672,N_1830,N_1896);
and U2673 (N_2673,N_1406,N_1988);
nor U2674 (N_2674,N_1624,N_1412);
nor U2675 (N_2675,N_1444,N_1760);
nand U2676 (N_2676,N_1245,N_1440);
or U2677 (N_2677,N_1109,N_1206);
nor U2678 (N_2678,N_1814,N_1859);
or U2679 (N_2679,N_1421,N_1840);
nand U2680 (N_2680,N_1767,N_1202);
and U2681 (N_2681,N_1811,N_1897);
xnor U2682 (N_2682,N_1304,N_1809);
nor U2683 (N_2683,N_1757,N_1125);
xor U2684 (N_2684,N_1670,N_1068);
and U2685 (N_2685,N_1545,N_1626);
nand U2686 (N_2686,N_1486,N_1880);
nand U2687 (N_2687,N_1308,N_1030);
or U2688 (N_2688,N_1759,N_1943);
nor U2689 (N_2689,N_1317,N_1424);
and U2690 (N_2690,N_1766,N_1969);
nand U2691 (N_2691,N_1230,N_1314);
or U2692 (N_2692,N_1280,N_1568);
nand U2693 (N_2693,N_1857,N_1978);
nand U2694 (N_2694,N_1976,N_1193);
nor U2695 (N_2695,N_1013,N_1327);
nand U2696 (N_2696,N_1957,N_1585);
and U2697 (N_2697,N_1155,N_1325);
and U2698 (N_2698,N_1572,N_1276);
nand U2699 (N_2699,N_1581,N_1613);
nor U2700 (N_2700,N_1363,N_1035);
and U2701 (N_2701,N_1719,N_1704);
nand U2702 (N_2702,N_1288,N_1740);
nand U2703 (N_2703,N_1508,N_1071);
or U2704 (N_2704,N_1838,N_1628);
or U2705 (N_2705,N_1385,N_1749);
nor U2706 (N_2706,N_1722,N_1006);
and U2707 (N_2707,N_1126,N_1757);
and U2708 (N_2708,N_1095,N_1699);
or U2709 (N_2709,N_1864,N_1194);
or U2710 (N_2710,N_1195,N_1165);
or U2711 (N_2711,N_1922,N_1014);
and U2712 (N_2712,N_1903,N_1036);
or U2713 (N_2713,N_1736,N_1490);
or U2714 (N_2714,N_1777,N_1902);
and U2715 (N_2715,N_1622,N_1858);
nor U2716 (N_2716,N_1579,N_1416);
or U2717 (N_2717,N_1845,N_1957);
nand U2718 (N_2718,N_1979,N_1940);
or U2719 (N_2719,N_1468,N_1528);
or U2720 (N_2720,N_1961,N_1363);
nor U2721 (N_2721,N_1428,N_1031);
nor U2722 (N_2722,N_1832,N_1209);
nor U2723 (N_2723,N_1962,N_1888);
or U2724 (N_2724,N_1706,N_1107);
xnor U2725 (N_2725,N_1970,N_1786);
and U2726 (N_2726,N_1257,N_1972);
or U2727 (N_2727,N_1821,N_1978);
and U2728 (N_2728,N_1733,N_1113);
and U2729 (N_2729,N_1081,N_1013);
nand U2730 (N_2730,N_1529,N_1892);
xor U2731 (N_2731,N_1066,N_1028);
nand U2732 (N_2732,N_1976,N_1015);
nand U2733 (N_2733,N_1785,N_1763);
or U2734 (N_2734,N_1397,N_1930);
nor U2735 (N_2735,N_1355,N_1134);
nand U2736 (N_2736,N_1487,N_1529);
nand U2737 (N_2737,N_1590,N_1686);
and U2738 (N_2738,N_1475,N_1007);
and U2739 (N_2739,N_1921,N_1059);
nand U2740 (N_2740,N_1062,N_1315);
nand U2741 (N_2741,N_1925,N_1215);
or U2742 (N_2742,N_1611,N_1140);
nor U2743 (N_2743,N_1976,N_1608);
nand U2744 (N_2744,N_1811,N_1022);
or U2745 (N_2745,N_1910,N_1969);
nor U2746 (N_2746,N_1263,N_1239);
or U2747 (N_2747,N_1070,N_1736);
nor U2748 (N_2748,N_1429,N_1644);
and U2749 (N_2749,N_1762,N_1423);
and U2750 (N_2750,N_1606,N_1012);
nand U2751 (N_2751,N_1989,N_1302);
nor U2752 (N_2752,N_1473,N_1386);
nand U2753 (N_2753,N_1536,N_1572);
and U2754 (N_2754,N_1121,N_1004);
and U2755 (N_2755,N_1622,N_1330);
or U2756 (N_2756,N_1977,N_1810);
nor U2757 (N_2757,N_1179,N_1055);
nor U2758 (N_2758,N_1379,N_1480);
nor U2759 (N_2759,N_1242,N_1462);
and U2760 (N_2760,N_1238,N_1898);
and U2761 (N_2761,N_1617,N_1058);
and U2762 (N_2762,N_1540,N_1045);
nor U2763 (N_2763,N_1114,N_1191);
or U2764 (N_2764,N_1067,N_1624);
and U2765 (N_2765,N_1741,N_1098);
nand U2766 (N_2766,N_1746,N_1758);
nand U2767 (N_2767,N_1895,N_1000);
or U2768 (N_2768,N_1031,N_1943);
xor U2769 (N_2769,N_1753,N_1014);
or U2770 (N_2770,N_1127,N_1535);
nor U2771 (N_2771,N_1973,N_1850);
and U2772 (N_2772,N_1535,N_1814);
or U2773 (N_2773,N_1088,N_1416);
nand U2774 (N_2774,N_1292,N_1737);
nor U2775 (N_2775,N_1159,N_1967);
nand U2776 (N_2776,N_1148,N_1899);
nand U2777 (N_2777,N_1117,N_1477);
or U2778 (N_2778,N_1364,N_1269);
nor U2779 (N_2779,N_1149,N_1312);
and U2780 (N_2780,N_1251,N_1959);
nor U2781 (N_2781,N_1194,N_1718);
nand U2782 (N_2782,N_1376,N_1723);
nor U2783 (N_2783,N_1971,N_1298);
or U2784 (N_2784,N_1334,N_1631);
and U2785 (N_2785,N_1866,N_1686);
or U2786 (N_2786,N_1358,N_1752);
xnor U2787 (N_2787,N_1144,N_1157);
and U2788 (N_2788,N_1759,N_1918);
nor U2789 (N_2789,N_1867,N_1362);
nand U2790 (N_2790,N_1555,N_1489);
or U2791 (N_2791,N_1281,N_1665);
nand U2792 (N_2792,N_1412,N_1129);
or U2793 (N_2793,N_1570,N_1013);
nor U2794 (N_2794,N_1195,N_1484);
xnor U2795 (N_2795,N_1488,N_1224);
and U2796 (N_2796,N_1659,N_1786);
xor U2797 (N_2797,N_1285,N_1747);
and U2798 (N_2798,N_1982,N_1225);
or U2799 (N_2799,N_1431,N_1200);
and U2800 (N_2800,N_1631,N_1372);
nor U2801 (N_2801,N_1549,N_1119);
or U2802 (N_2802,N_1221,N_1191);
or U2803 (N_2803,N_1196,N_1815);
nand U2804 (N_2804,N_1729,N_1281);
nand U2805 (N_2805,N_1273,N_1639);
and U2806 (N_2806,N_1084,N_1447);
nand U2807 (N_2807,N_1616,N_1762);
and U2808 (N_2808,N_1035,N_1374);
and U2809 (N_2809,N_1275,N_1207);
or U2810 (N_2810,N_1823,N_1335);
and U2811 (N_2811,N_1608,N_1071);
and U2812 (N_2812,N_1796,N_1007);
nand U2813 (N_2813,N_1275,N_1582);
and U2814 (N_2814,N_1106,N_1816);
or U2815 (N_2815,N_1499,N_1943);
and U2816 (N_2816,N_1738,N_1121);
nor U2817 (N_2817,N_1741,N_1037);
and U2818 (N_2818,N_1717,N_1529);
nand U2819 (N_2819,N_1061,N_1267);
xor U2820 (N_2820,N_1251,N_1064);
nor U2821 (N_2821,N_1270,N_1876);
nand U2822 (N_2822,N_1103,N_1024);
xor U2823 (N_2823,N_1858,N_1651);
nor U2824 (N_2824,N_1251,N_1053);
and U2825 (N_2825,N_1205,N_1593);
or U2826 (N_2826,N_1110,N_1164);
nand U2827 (N_2827,N_1066,N_1659);
or U2828 (N_2828,N_1829,N_1226);
and U2829 (N_2829,N_1146,N_1350);
or U2830 (N_2830,N_1117,N_1161);
nor U2831 (N_2831,N_1295,N_1624);
nand U2832 (N_2832,N_1704,N_1254);
or U2833 (N_2833,N_1824,N_1451);
and U2834 (N_2834,N_1683,N_1823);
nor U2835 (N_2835,N_1169,N_1003);
xor U2836 (N_2836,N_1814,N_1274);
and U2837 (N_2837,N_1869,N_1640);
or U2838 (N_2838,N_1608,N_1885);
or U2839 (N_2839,N_1963,N_1474);
or U2840 (N_2840,N_1117,N_1254);
nor U2841 (N_2841,N_1626,N_1947);
nor U2842 (N_2842,N_1220,N_1905);
and U2843 (N_2843,N_1773,N_1912);
nor U2844 (N_2844,N_1221,N_1931);
nor U2845 (N_2845,N_1202,N_1070);
or U2846 (N_2846,N_1864,N_1134);
and U2847 (N_2847,N_1324,N_1143);
nor U2848 (N_2848,N_1527,N_1389);
or U2849 (N_2849,N_1638,N_1479);
and U2850 (N_2850,N_1177,N_1835);
and U2851 (N_2851,N_1908,N_1768);
nand U2852 (N_2852,N_1157,N_1697);
nor U2853 (N_2853,N_1795,N_1008);
nand U2854 (N_2854,N_1199,N_1783);
or U2855 (N_2855,N_1360,N_1612);
or U2856 (N_2856,N_1734,N_1328);
nand U2857 (N_2857,N_1782,N_1965);
or U2858 (N_2858,N_1100,N_1405);
nor U2859 (N_2859,N_1793,N_1769);
xor U2860 (N_2860,N_1077,N_1108);
or U2861 (N_2861,N_1394,N_1133);
and U2862 (N_2862,N_1925,N_1401);
nor U2863 (N_2863,N_1416,N_1182);
nand U2864 (N_2864,N_1237,N_1606);
or U2865 (N_2865,N_1257,N_1188);
and U2866 (N_2866,N_1122,N_1445);
and U2867 (N_2867,N_1286,N_1722);
nand U2868 (N_2868,N_1099,N_1982);
xnor U2869 (N_2869,N_1382,N_1795);
xor U2870 (N_2870,N_1805,N_1488);
nand U2871 (N_2871,N_1945,N_1036);
and U2872 (N_2872,N_1150,N_1473);
and U2873 (N_2873,N_1849,N_1295);
nand U2874 (N_2874,N_1457,N_1666);
nand U2875 (N_2875,N_1978,N_1296);
or U2876 (N_2876,N_1837,N_1372);
nand U2877 (N_2877,N_1532,N_1671);
nor U2878 (N_2878,N_1638,N_1567);
or U2879 (N_2879,N_1194,N_1856);
and U2880 (N_2880,N_1837,N_1171);
nand U2881 (N_2881,N_1270,N_1967);
and U2882 (N_2882,N_1430,N_1654);
nand U2883 (N_2883,N_1641,N_1793);
and U2884 (N_2884,N_1421,N_1627);
nor U2885 (N_2885,N_1324,N_1246);
or U2886 (N_2886,N_1698,N_1932);
nand U2887 (N_2887,N_1165,N_1695);
nand U2888 (N_2888,N_1659,N_1750);
nor U2889 (N_2889,N_1393,N_1193);
nor U2890 (N_2890,N_1035,N_1111);
nand U2891 (N_2891,N_1156,N_1640);
or U2892 (N_2892,N_1860,N_1606);
nand U2893 (N_2893,N_1083,N_1907);
nand U2894 (N_2894,N_1283,N_1767);
nor U2895 (N_2895,N_1851,N_1801);
nand U2896 (N_2896,N_1123,N_1318);
nand U2897 (N_2897,N_1801,N_1272);
nand U2898 (N_2898,N_1928,N_1012);
or U2899 (N_2899,N_1315,N_1474);
nor U2900 (N_2900,N_1084,N_1555);
and U2901 (N_2901,N_1485,N_1473);
and U2902 (N_2902,N_1518,N_1788);
or U2903 (N_2903,N_1521,N_1682);
and U2904 (N_2904,N_1660,N_1025);
nand U2905 (N_2905,N_1309,N_1999);
or U2906 (N_2906,N_1835,N_1847);
and U2907 (N_2907,N_1465,N_1287);
or U2908 (N_2908,N_1864,N_1802);
nor U2909 (N_2909,N_1555,N_1050);
and U2910 (N_2910,N_1306,N_1067);
nor U2911 (N_2911,N_1132,N_1095);
nand U2912 (N_2912,N_1462,N_1914);
nand U2913 (N_2913,N_1326,N_1797);
nor U2914 (N_2914,N_1884,N_1253);
or U2915 (N_2915,N_1396,N_1996);
nor U2916 (N_2916,N_1221,N_1066);
nand U2917 (N_2917,N_1382,N_1443);
and U2918 (N_2918,N_1204,N_1564);
nor U2919 (N_2919,N_1436,N_1334);
nand U2920 (N_2920,N_1553,N_1262);
nand U2921 (N_2921,N_1495,N_1838);
nand U2922 (N_2922,N_1590,N_1881);
or U2923 (N_2923,N_1206,N_1056);
nor U2924 (N_2924,N_1502,N_1770);
nand U2925 (N_2925,N_1986,N_1401);
or U2926 (N_2926,N_1396,N_1408);
nor U2927 (N_2927,N_1039,N_1858);
and U2928 (N_2928,N_1099,N_1798);
and U2929 (N_2929,N_1538,N_1498);
or U2930 (N_2930,N_1967,N_1739);
nand U2931 (N_2931,N_1268,N_1941);
nor U2932 (N_2932,N_1090,N_1702);
nor U2933 (N_2933,N_1921,N_1180);
or U2934 (N_2934,N_1744,N_1046);
and U2935 (N_2935,N_1846,N_1393);
nor U2936 (N_2936,N_1483,N_1329);
and U2937 (N_2937,N_1899,N_1777);
nor U2938 (N_2938,N_1046,N_1232);
or U2939 (N_2939,N_1512,N_1725);
xor U2940 (N_2940,N_1712,N_1042);
xor U2941 (N_2941,N_1427,N_1361);
nand U2942 (N_2942,N_1372,N_1951);
and U2943 (N_2943,N_1735,N_1112);
or U2944 (N_2944,N_1399,N_1708);
nand U2945 (N_2945,N_1276,N_1359);
or U2946 (N_2946,N_1627,N_1990);
and U2947 (N_2947,N_1046,N_1835);
xor U2948 (N_2948,N_1410,N_1720);
and U2949 (N_2949,N_1479,N_1186);
nor U2950 (N_2950,N_1114,N_1851);
xnor U2951 (N_2951,N_1481,N_1718);
nand U2952 (N_2952,N_1828,N_1791);
nor U2953 (N_2953,N_1265,N_1819);
or U2954 (N_2954,N_1521,N_1591);
nor U2955 (N_2955,N_1134,N_1925);
nor U2956 (N_2956,N_1198,N_1878);
or U2957 (N_2957,N_1627,N_1356);
xnor U2958 (N_2958,N_1218,N_1361);
and U2959 (N_2959,N_1739,N_1216);
nor U2960 (N_2960,N_1254,N_1802);
nand U2961 (N_2961,N_1054,N_1467);
and U2962 (N_2962,N_1021,N_1717);
or U2963 (N_2963,N_1593,N_1250);
and U2964 (N_2964,N_1427,N_1782);
and U2965 (N_2965,N_1458,N_1573);
and U2966 (N_2966,N_1352,N_1575);
and U2967 (N_2967,N_1135,N_1549);
nand U2968 (N_2968,N_1870,N_1990);
nand U2969 (N_2969,N_1228,N_1695);
nor U2970 (N_2970,N_1746,N_1431);
nand U2971 (N_2971,N_1417,N_1132);
and U2972 (N_2972,N_1449,N_1922);
nor U2973 (N_2973,N_1369,N_1555);
and U2974 (N_2974,N_1386,N_1523);
or U2975 (N_2975,N_1522,N_1486);
nor U2976 (N_2976,N_1139,N_1307);
and U2977 (N_2977,N_1489,N_1660);
or U2978 (N_2978,N_1159,N_1295);
nand U2979 (N_2979,N_1916,N_1848);
or U2980 (N_2980,N_1016,N_1596);
or U2981 (N_2981,N_1049,N_1326);
or U2982 (N_2982,N_1546,N_1434);
nand U2983 (N_2983,N_1372,N_1675);
or U2984 (N_2984,N_1065,N_1369);
and U2985 (N_2985,N_1182,N_1094);
nor U2986 (N_2986,N_1755,N_1926);
xnor U2987 (N_2987,N_1860,N_1273);
nor U2988 (N_2988,N_1877,N_1078);
or U2989 (N_2989,N_1219,N_1610);
nor U2990 (N_2990,N_1654,N_1458);
and U2991 (N_2991,N_1029,N_1060);
or U2992 (N_2992,N_1590,N_1144);
or U2993 (N_2993,N_1947,N_1518);
and U2994 (N_2994,N_1541,N_1660);
nor U2995 (N_2995,N_1975,N_1670);
or U2996 (N_2996,N_1395,N_1143);
and U2997 (N_2997,N_1446,N_1908);
and U2998 (N_2998,N_1786,N_1741);
nor U2999 (N_2999,N_1052,N_1440);
nor U3000 (N_3000,N_2198,N_2683);
nand U3001 (N_3001,N_2040,N_2521);
nand U3002 (N_3002,N_2454,N_2249);
nand U3003 (N_3003,N_2897,N_2688);
nand U3004 (N_3004,N_2921,N_2136);
xnor U3005 (N_3005,N_2226,N_2647);
nand U3006 (N_3006,N_2819,N_2134);
nor U3007 (N_3007,N_2391,N_2724);
and U3008 (N_3008,N_2761,N_2477);
xor U3009 (N_3009,N_2227,N_2809);
or U3010 (N_3010,N_2919,N_2772);
or U3011 (N_3011,N_2931,N_2725);
nor U3012 (N_3012,N_2052,N_2442);
nand U3013 (N_3013,N_2902,N_2885);
or U3014 (N_3014,N_2230,N_2263);
and U3015 (N_3015,N_2039,N_2103);
nand U3016 (N_3016,N_2755,N_2355);
nor U3017 (N_3017,N_2232,N_2085);
nand U3018 (N_3018,N_2543,N_2874);
and U3019 (N_3019,N_2468,N_2238);
nand U3020 (N_3020,N_2455,N_2222);
nand U3021 (N_3021,N_2267,N_2182);
or U3022 (N_3022,N_2627,N_2786);
or U3023 (N_3023,N_2090,N_2169);
or U3024 (N_3024,N_2882,N_2953);
xnor U3025 (N_3025,N_2569,N_2705);
nor U3026 (N_3026,N_2423,N_2638);
nor U3027 (N_3027,N_2504,N_2250);
xor U3028 (N_3028,N_2133,N_2609);
xnor U3029 (N_3029,N_2219,N_2907);
nand U3030 (N_3030,N_2000,N_2561);
and U3031 (N_3031,N_2694,N_2354);
and U3032 (N_3032,N_2181,N_2390);
nor U3033 (N_3033,N_2110,N_2572);
and U3034 (N_3034,N_2971,N_2240);
xor U3035 (N_3035,N_2139,N_2838);
nand U3036 (N_3036,N_2845,N_2371);
nand U3037 (N_3037,N_2324,N_2239);
and U3038 (N_3038,N_2526,N_2422);
nand U3039 (N_3039,N_2474,N_2911);
xnor U3040 (N_3040,N_2899,N_2787);
nor U3041 (N_3041,N_2886,N_2369);
xnor U3042 (N_3042,N_2934,N_2395);
nand U3043 (N_3043,N_2550,N_2475);
or U3044 (N_3044,N_2042,N_2245);
nand U3045 (N_3045,N_2457,N_2863);
nand U3046 (N_3046,N_2187,N_2614);
nand U3047 (N_3047,N_2758,N_2428);
nor U3048 (N_3048,N_2447,N_2165);
nand U3049 (N_3049,N_2028,N_2364);
and U3050 (N_3050,N_2545,N_2008);
xor U3051 (N_3051,N_2681,N_2795);
and U3052 (N_3052,N_2098,N_2484);
xnor U3053 (N_3053,N_2106,N_2376);
or U3054 (N_3054,N_2556,N_2692);
nor U3055 (N_3055,N_2224,N_2962);
nor U3056 (N_3056,N_2112,N_2316);
nand U3057 (N_3057,N_2487,N_2126);
nor U3058 (N_3058,N_2602,N_2933);
and U3059 (N_3059,N_2818,N_2483);
and U3060 (N_3060,N_2436,N_2805);
nand U3061 (N_3061,N_2349,N_2438);
and U3062 (N_3062,N_2288,N_2412);
nand U3063 (N_3063,N_2651,N_2381);
nor U3064 (N_3064,N_2485,N_2065);
nor U3065 (N_3065,N_2678,N_2220);
nand U3066 (N_3066,N_2603,N_2654);
xnor U3067 (N_3067,N_2033,N_2858);
and U3068 (N_3068,N_2401,N_2168);
nand U3069 (N_3069,N_2489,N_2690);
or U3070 (N_3070,N_2014,N_2900);
or U3071 (N_3071,N_2473,N_2307);
or U3072 (N_3072,N_2597,N_2036);
nor U3073 (N_3073,N_2937,N_2659);
nand U3074 (N_3074,N_2520,N_2914);
nand U3075 (N_3075,N_2820,N_2979);
nor U3076 (N_3076,N_2549,N_2162);
nand U3077 (N_3077,N_2124,N_2613);
or U3078 (N_3078,N_2070,N_2723);
and U3079 (N_3079,N_2164,N_2233);
xor U3080 (N_3080,N_2975,N_2687);
nor U3081 (N_3081,N_2693,N_2793);
xnor U3082 (N_3082,N_2655,N_2924);
or U3083 (N_3083,N_2199,N_2857);
and U3084 (N_3084,N_2449,N_2297);
and U3085 (N_3085,N_2575,N_2825);
nand U3086 (N_3086,N_2301,N_2741);
or U3087 (N_3087,N_2987,N_2606);
nor U3088 (N_3088,N_2947,N_2887);
nand U3089 (N_3089,N_2289,N_2174);
nand U3090 (N_3090,N_2822,N_2275);
and U3091 (N_3091,N_2806,N_2406);
and U3092 (N_3092,N_2470,N_2508);
and U3093 (N_3093,N_2045,N_2326);
nor U3094 (N_3094,N_2754,N_2257);
xnor U3095 (N_3095,N_2643,N_2298);
or U3096 (N_3096,N_2127,N_2202);
nand U3097 (N_3097,N_2954,N_2993);
or U3098 (N_3098,N_2519,N_2766);
or U3099 (N_3099,N_2185,N_2328);
nor U3100 (N_3100,N_2350,N_2961);
or U3101 (N_3101,N_2781,N_2721);
nand U3102 (N_3102,N_2827,N_2808);
nor U3103 (N_3103,N_2667,N_2679);
or U3104 (N_3104,N_2970,N_2459);
nand U3105 (N_3105,N_2161,N_2178);
xor U3106 (N_3106,N_2498,N_2300);
or U3107 (N_3107,N_2749,N_2022);
and U3108 (N_3108,N_2216,N_2205);
or U3109 (N_3109,N_2278,N_2864);
and U3110 (N_3110,N_2372,N_2906);
nand U3111 (N_3111,N_2844,N_2190);
nor U3112 (N_3112,N_2876,N_2195);
and U3113 (N_3113,N_2591,N_2756);
nor U3114 (N_3114,N_2676,N_2061);
or U3115 (N_3115,N_2285,N_2035);
nand U3116 (N_3116,N_2730,N_2941);
or U3117 (N_3117,N_2336,N_2833);
xnor U3118 (N_3118,N_2433,N_2612);
or U3119 (N_3119,N_2317,N_2523);
xnor U3120 (N_3120,N_2091,N_2341);
or U3121 (N_3121,N_2744,N_2983);
nand U3122 (N_3122,N_2020,N_2742);
nor U3123 (N_3123,N_2658,N_2567);
xnor U3124 (N_3124,N_2813,N_2560);
and U3125 (N_3125,N_2728,N_2765);
nand U3126 (N_3126,N_2367,N_2034);
xnor U3127 (N_3127,N_2430,N_2751);
nand U3128 (N_3128,N_2154,N_2172);
nor U3129 (N_3129,N_2850,N_2163);
and U3130 (N_3130,N_2479,N_2048);
nor U3131 (N_3131,N_2878,N_2529);
nor U3132 (N_3132,N_2284,N_2365);
or U3133 (N_3133,N_2616,N_2265);
nor U3134 (N_3134,N_2571,N_2225);
nor U3135 (N_3135,N_2720,N_2566);
nand U3136 (N_3136,N_2645,N_2060);
nor U3137 (N_3137,N_2290,N_2269);
or U3138 (N_3138,N_2596,N_2246);
or U3139 (N_3139,N_2434,N_2228);
nand U3140 (N_3140,N_2502,N_2122);
and U3141 (N_3141,N_2244,N_2166);
xnor U3142 (N_3142,N_2535,N_2757);
nand U3143 (N_3143,N_2105,N_2204);
and U3144 (N_3144,N_2778,N_2404);
or U3145 (N_3145,N_2461,N_2894);
nor U3146 (N_3146,N_2506,N_2294);
nor U3147 (N_3147,N_2149,N_2836);
or U3148 (N_3148,N_2623,N_2665);
or U3149 (N_3149,N_2991,N_2184);
nor U3150 (N_3150,N_2366,N_2160);
and U3151 (N_3151,N_2088,N_2837);
nor U3152 (N_3152,N_2405,N_2243);
and U3153 (N_3153,N_2291,N_2703);
nor U3154 (N_3154,N_2069,N_2792);
nand U3155 (N_3155,N_2802,N_2699);
xor U3156 (N_3156,N_2025,N_2064);
or U3157 (N_3157,N_2377,N_2305);
nand U3158 (N_3158,N_2829,N_2223);
or U3159 (N_3159,N_2096,N_2598);
xnor U3160 (N_3160,N_2399,N_2691);
or U3161 (N_3161,N_2717,N_2200);
or U3162 (N_3162,N_2628,N_2488);
xnor U3163 (N_3163,N_2839,N_2218);
and U3164 (N_3164,N_2943,N_2242);
nor U3165 (N_3165,N_2080,N_2023);
or U3166 (N_3166,N_2932,N_2056);
xnor U3167 (N_3167,N_2775,N_2279);
and U3168 (N_3168,N_2800,N_2729);
nand U3169 (N_3169,N_2558,N_2344);
or U3170 (N_3170,N_2002,N_2856);
nand U3171 (N_3171,N_2977,N_2453);
or U3172 (N_3172,N_2854,N_2905);
and U3173 (N_3173,N_2736,N_2109);
xor U3174 (N_3174,N_2649,N_2472);
nand U3175 (N_3175,N_2686,N_2790);
and U3176 (N_3176,N_2896,N_2142);
and U3177 (N_3177,N_2562,N_2570);
nand U3178 (N_3178,N_2582,N_2868);
and U3179 (N_3179,N_2817,N_2051);
nand U3180 (N_3180,N_2481,N_2927);
nand U3181 (N_3181,N_2304,N_2147);
nor U3182 (N_3182,N_2115,N_2893);
nor U3183 (N_3183,N_2965,N_2116);
nand U3184 (N_3184,N_2215,N_2752);
nand U3185 (N_3185,N_2746,N_2611);
nand U3186 (N_3186,N_2770,N_2462);
or U3187 (N_3187,N_2068,N_2231);
nand U3188 (N_3188,N_2458,N_2338);
and U3189 (N_3189,N_2939,N_2392);
nor U3190 (N_3190,N_2276,N_2092);
nor U3191 (N_3191,N_2875,N_2985);
and U3192 (N_3192,N_2062,N_2855);
nand U3193 (N_3193,N_2920,N_2883);
xnor U3194 (N_3194,N_2511,N_2674);
nand U3195 (N_3195,N_2415,N_2016);
or U3196 (N_3196,N_2049,N_2201);
xnor U3197 (N_3197,N_2083,N_2140);
or U3198 (N_3198,N_2210,N_2236);
and U3199 (N_3199,N_2492,N_2329);
xnor U3200 (N_3200,N_2776,N_2135);
nand U3201 (N_3201,N_2918,N_2644);
and U3202 (N_3202,N_2880,N_2797);
nor U3203 (N_3203,N_2258,N_2617);
nor U3204 (N_3204,N_2928,N_2141);
xnor U3205 (N_3205,N_2500,N_2830);
nand U3206 (N_3206,N_2066,N_2534);
nand U3207 (N_3207,N_2302,N_2007);
or U3208 (N_3208,N_2960,N_2144);
nand U3209 (N_3209,N_2642,N_2347);
or U3210 (N_3210,N_2320,N_2196);
nand U3211 (N_3211,N_2234,N_2537);
nand U3212 (N_3212,N_2451,N_2248);
nor U3213 (N_3213,N_2807,N_2622);
and U3214 (N_3214,N_2426,N_2277);
and U3215 (N_3215,N_2408,N_2132);
nand U3216 (N_3216,N_2113,N_2386);
or U3217 (N_3217,N_2966,N_2890);
or U3218 (N_3218,N_2726,N_2359);
nor U3219 (N_3219,N_2945,N_2539);
xnor U3220 (N_3220,N_2476,N_2959);
nand U3221 (N_3221,N_2058,N_2176);
and U3222 (N_3222,N_2646,N_2211);
nor U3223 (N_3223,N_2926,N_2074);
and U3224 (N_3224,N_2026,N_2564);
nand U3225 (N_3225,N_2385,N_2716);
and U3226 (N_3226,N_2400,N_2949);
nor U3227 (N_3227,N_2273,N_2374);
nand U3228 (N_3228,N_2173,N_2138);
and U3229 (N_3229,N_2771,N_2794);
nor U3230 (N_3230,N_2929,N_2394);
and U3231 (N_3231,N_2525,N_2727);
nor U3232 (N_3232,N_2626,N_2984);
xor U3233 (N_3233,N_2997,N_2750);
nor U3234 (N_3234,N_2318,N_2397);
and U3235 (N_3235,N_2266,N_2873);
nand U3236 (N_3236,N_2403,N_2621);
and U3237 (N_3237,N_2860,N_2774);
nand U3238 (N_3238,N_2710,N_2013);
nand U3239 (N_3239,N_2573,N_2235);
nor U3240 (N_3240,N_2541,N_2956);
nor U3241 (N_3241,N_2313,N_2432);
nor U3242 (N_3242,N_2043,N_2670);
nand U3243 (N_3243,N_2206,N_2824);
and U3244 (N_3244,N_2912,N_2292);
or U3245 (N_3245,N_2557,N_2588);
nand U3246 (N_3246,N_2634,N_2847);
and U3247 (N_3247,N_2865,N_2624);
and U3248 (N_3248,N_2321,N_2779);
and U3249 (N_3249,N_2396,N_2763);
nor U3250 (N_3250,N_2047,N_2437);
nor U3251 (N_3251,N_2950,N_2996);
and U3252 (N_3252,N_2895,N_2063);
nand U3253 (N_3253,N_2496,N_2466);
nand U3254 (N_3254,N_2524,N_2375);
nand U3255 (N_3255,N_2361,N_2517);
or U3256 (N_3256,N_2274,N_2107);
nor U3257 (N_3257,N_2203,N_2981);
and U3258 (N_3258,N_2814,N_2170);
and U3259 (N_3259,N_2417,N_2859);
xor U3260 (N_3260,N_2700,N_2828);
nand U3261 (N_3261,N_2425,N_2031);
nand U3262 (N_3262,N_2348,N_2711);
and U3263 (N_3263,N_2785,N_2652);
nor U3264 (N_3264,N_2282,N_2853);
nand U3265 (N_3265,N_2054,N_2281);
and U3266 (N_3266,N_2323,N_2363);
nor U3267 (N_3267,N_2186,N_2935);
nand U3268 (N_3268,N_2682,N_2333);
or U3269 (N_3269,N_2759,N_2578);
nor U3270 (N_3270,N_2146,N_2259);
nand U3271 (N_3271,N_2995,N_2393);
nand U3272 (N_3272,N_2082,N_2576);
nor U3273 (N_3273,N_2528,N_2641);
nor U3274 (N_3274,N_2384,N_2099);
nor U3275 (N_3275,N_2252,N_2019);
or U3276 (N_3276,N_2118,N_2293);
nor U3277 (N_3277,N_2695,N_2590);
nor U3278 (N_3278,N_2319,N_2743);
xor U3279 (N_3279,N_2762,N_2867);
nand U3280 (N_3280,N_2669,N_2509);
or U3281 (N_3281,N_2119,N_2131);
or U3282 (N_3282,N_2471,N_2811);
or U3283 (N_3283,N_2898,N_2680);
nand U3284 (N_3284,N_2256,N_2214);
xnor U3285 (N_3285,N_2071,N_2130);
and U3286 (N_3286,N_2769,N_2101);
xnor U3287 (N_3287,N_2358,N_2418);
nand U3288 (N_3288,N_2078,N_2413);
and U3289 (N_3289,N_2387,N_2490);
or U3290 (N_3290,N_2055,N_2701);
nor U3291 (N_3291,N_2656,N_2512);
or U3292 (N_3292,N_2870,N_2798);
or U3293 (N_3293,N_2137,N_2102);
nor U3294 (N_3294,N_2255,N_2183);
nand U3295 (N_3295,N_2123,N_2310);
xor U3296 (N_3296,N_2563,N_2908);
nand U3297 (N_3297,N_2969,N_2677);
nor U3298 (N_3298,N_2610,N_2788);
or U3299 (N_3299,N_2901,N_2012);
nor U3300 (N_3300,N_2330,N_2823);
or U3301 (N_3301,N_2673,N_2346);
nand U3302 (N_3302,N_2017,N_2153);
nor U3303 (N_3303,N_2041,N_2536);
nand U3304 (N_3304,N_2922,N_2826);
and U3305 (N_3305,N_2579,N_2930);
and U3306 (N_3306,N_2117,N_2988);
or U3307 (N_3307,N_2456,N_2059);
nor U3308 (N_3308,N_2286,N_2664);
or U3309 (N_3309,N_2668,N_2378);
and U3310 (N_3310,N_2208,N_2532);
nor U3311 (N_3311,N_2650,N_2325);
and U3312 (N_3312,N_2555,N_2663);
nand U3313 (N_3313,N_2948,N_2803);
nor U3314 (N_3314,N_2848,N_2915);
or U3315 (N_3315,N_2832,N_2018);
nor U3316 (N_3316,N_2862,N_2072);
nand U3317 (N_3317,N_2424,N_2849);
and U3318 (N_3318,N_2871,N_2601);
nand U3319 (N_3319,N_2760,N_2067);
nand U3320 (N_3320,N_2335,N_2379);
or U3321 (N_3321,N_2768,N_2270);
nor U3322 (N_3322,N_2212,N_2799);
or U3323 (N_3323,N_2815,N_2308);
xor U3324 (N_3324,N_2331,N_2731);
and U3325 (N_3325,N_2145,N_2493);
and U3326 (N_3326,N_2167,N_2129);
xnor U3327 (N_3327,N_2005,N_2619);
and U3328 (N_3328,N_2574,N_2639);
or U3329 (N_3329,N_2660,N_2618);
or U3330 (N_3330,N_2419,N_2531);
and U3331 (N_3331,N_2514,N_2306);
and U3332 (N_3332,N_2260,N_2990);
nand U3333 (N_3333,N_2152,N_2209);
and U3334 (N_3334,N_2748,N_2625);
or U3335 (N_3335,N_2075,N_2356);
and U3336 (N_3336,N_2444,N_2565);
and U3337 (N_3337,N_2095,N_2734);
xor U3338 (N_3338,N_2188,N_2151);
and U3339 (N_3339,N_2967,N_2339);
and U3340 (N_3340,N_2719,N_2009);
nor U3341 (N_3341,N_2380,N_2604);
nor U3342 (N_3342,N_2093,N_2001);
nand U3343 (N_3343,N_2450,N_2046);
or U3344 (N_3344,N_2964,N_2630);
or U3345 (N_3345,N_2121,N_2334);
or U3346 (N_3346,N_2373,N_2615);
or U3347 (N_3347,N_2010,N_2552);
nand U3348 (N_3348,N_2207,N_2309);
nor U3349 (N_3349,N_2636,N_2006);
nor U3350 (N_3350,N_2992,N_2503);
nor U3351 (N_3351,N_2904,N_2360);
nor U3352 (N_3352,N_2241,N_2972);
and U3353 (N_3353,N_2280,N_2559);
or U3354 (N_3354,N_2217,N_2675);
or U3355 (N_3355,N_2494,N_2159);
nand U3356 (N_3356,N_2702,N_2327);
or U3357 (N_3357,N_2831,N_2733);
and U3358 (N_3358,N_2938,N_2577);
or U3359 (N_3359,N_2689,N_2707);
or U3360 (N_3360,N_2251,N_2445);
and U3361 (N_3361,N_2100,N_2592);
xnor U3362 (N_3362,N_2816,N_2986);
and U3363 (N_3363,N_2024,N_2653);
nor U3364 (N_3364,N_2037,N_2084);
nor U3365 (N_3365,N_2957,N_2551);
nand U3366 (N_3366,N_2580,N_2889);
nand U3367 (N_3367,N_2057,N_2633);
or U3368 (N_3368,N_2029,N_2311);
nor U3369 (N_3369,N_2662,N_2343);
and U3370 (N_3370,N_2314,N_2732);
nor U3371 (N_3371,N_2465,N_2843);
nor U3372 (N_3372,N_2852,N_2715);
or U3373 (N_3373,N_2411,N_2073);
nand U3374 (N_3374,N_2158,N_2801);
and U3375 (N_3375,N_2632,N_2478);
nor U3376 (N_3376,N_2076,N_2157);
and U3377 (N_3377,N_2999,N_2342);
nor U3378 (N_3378,N_2104,N_2607);
or U3379 (N_3379,N_2989,N_2722);
nand U3380 (N_3380,N_2388,N_2357);
nand U3381 (N_3381,N_2782,N_2974);
nor U3382 (N_3382,N_2629,N_2299);
or U3383 (N_3383,N_2542,N_2540);
nand U3384 (N_3384,N_2946,N_2963);
or U3385 (N_3385,N_2398,N_2796);
nor U3386 (N_3386,N_2467,N_2955);
and U3387 (N_3387,N_2495,N_2463);
and U3388 (N_3388,N_2546,N_2175);
and U3389 (N_3389,N_2353,N_2745);
nand U3390 (N_3390,N_2261,N_2709);
nor U3391 (N_3391,N_2586,N_2410);
nor U3392 (N_3392,N_2156,N_2268);
nand U3393 (N_3393,N_2704,N_2253);
or U3394 (N_3394,N_2708,N_2108);
nand U3395 (N_3395,N_2114,N_2735);
nand U3396 (N_3396,N_2595,N_2620);
and U3397 (N_3397,N_2522,N_2978);
nand U3398 (N_3398,N_2877,N_2368);
or U3399 (N_3399,N_2530,N_2737);
or U3400 (N_3400,N_2697,N_2581);
nand U3401 (N_3401,N_2671,N_2407);
nor U3402 (N_3402,N_2191,N_2976);
nand U3403 (N_3403,N_2337,N_2443);
nor U3404 (N_3404,N_2194,N_2402);
nand U3405 (N_3405,N_2420,N_2891);
or U3406 (N_3406,N_2583,N_2777);
nand U3407 (N_3407,N_2180,N_2648);
xor U3408 (N_3408,N_2189,N_2544);
or U3409 (N_3409,N_2125,N_2527);
nand U3410 (N_3410,N_2605,N_2846);
or U3411 (N_3411,N_2295,N_2910);
and U3412 (N_3412,N_2370,N_2916);
xnor U3413 (N_3413,N_2128,N_2315);
xor U3414 (N_3414,N_2942,N_2784);
and U3415 (N_3415,N_2143,N_2851);
and U3416 (N_3416,N_2427,N_2739);
and U3417 (N_3417,N_2821,N_2296);
nand U3418 (N_3418,N_2038,N_2952);
nor U3419 (N_3419,N_2482,N_2486);
and U3420 (N_3420,N_2764,N_2177);
or U3421 (N_3421,N_2698,N_2553);
and U3422 (N_3422,N_2448,N_2460);
nand U3423 (N_3423,N_2740,N_2272);
or U3424 (N_3424,N_2980,N_2672);
and U3425 (N_3425,N_2469,N_2909);
or U3426 (N_3426,N_2712,N_2303);
or U3427 (N_3427,N_2538,N_2050);
or U3428 (N_3428,N_2213,N_2841);
xnor U3429 (N_3429,N_2352,N_2738);
nor U3430 (N_3430,N_2507,N_2869);
or U3431 (N_3431,N_2600,N_2666);
or U3432 (N_3432,N_2155,N_2322);
and U3433 (N_3433,N_2593,N_2086);
or U3434 (N_3434,N_2568,N_2081);
nor U3435 (N_3435,N_2747,N_2441);
xor U3436 (N_3436,N_2903,N_2079);
nand U3437 (N_3437,N_2513,N_2015);
nor U3438 (N_3438,N_2554,N_2030);
xor U3439 (N_3439,N_2192,N_2497);
xnor U3440 (N_3440,N_2684,N_2362);
and U3441 (N_3441,N_2608,N_2003);
nand U3442 (N_3442,N_2594,N_2925);
nand U3443 (N_3443,N_2958,N_2637);
and U3444 (N_3444,N_2714,N_2416);
nand U3445 (N_3445,N_2812,N_2271);
nand U3446 (N_3446,N_2789,N_2247);
or U3447 (N_3447,N_2439,N_2718);
nand U3448 (N_3448,N_2657,N_2501);
nor U3449 (N_3449,N_2835,N_2810);
or U3450 (N_3450,N_2077,N_2094);
or U3451 (N_3451,N_2446,N_2409);
xnor U3452 (N_3452,N_2791,N_2193);
xnor U3453 (N_3453,N_2968,N_2340);
nor U3454 (N_3454,N_2510,N_2685);
nand U3455 (N_3455,N_2533,N_2753);
and U3456 (N_3456,N_2936,N_2767);
nor U3457 (N_3457,N_2599,N_2585);
and U3458 (N_3458,N_2262,N_2713);
or U3459 (N_3459,N_2383,N_2923);
or U3460 (N_3460,N_2435,N_2089);
nor U3461 (N_3461,N_2773,N_2881);
and U3462 (N_3462,N_2884,N_2097);
nand U3463 (N_3463,N_2515,N_2548);
or U3464 (N_3464,N_2706,N_2345);
nand U3465 (N_3465,N_2229,N_2998);
or U3466 (N_3466,N_2021,N_2892);
or U3467 (N_3467,N_2452,N_2429);
nand U3468 (N_3468,N_2505,N_2414);
xnor U3469 (N_3469,N_2032,N_2237);
and U3470 (N_3470,N_2351,N_2834);
or U3471 (N_3471,N_2547,N_2491);
xor U3472 (N_3472,N_2879,N_2004);
nor U3473 (N_3473,N_2866,N_2940);
nor U3474 (N_3474,N_2888,N_2872);
xor U3475 (N_3475,N_2421,N_2780);
or U3476 (N_3476,N_2332,N_2661);
xor U3477 (N_3477,N_2516,N_2842);
or U3478 (N_3478,N_2587,N_2861);
and U3479 (N_3479,N_2221,N_2640);
xnor U3480 (N_3480,N_2464,N_2382);
nand U3481 (N_3481,N_2171,N_2584);
nand U3482 (N_3482,N_2783,N_2804);
nor U3483 (N_3483,N_2011,N_2053);
nand U3484 (N_3484,N_2389,N_2148);
nor U3485 (N_3485,N_2044,N_2480);
and U3486 (N_3486,N_2518,N_2913);
and U3487 (N_3487,N_2264,N_2087);
xor U3488 (N_3488,N_2287,N_2917);
nor U3489 (N_3489,N_2973,N_2944);
nor U3490 (N_3490,N_2197,N_2431);
or U3491 (N_3491,N_2312,N_2150);
or U3492 (N_3492,N_2982,N_2179);
or U3493 (N_3493,N_2120,N_2951);
nand U3494 (N_3494,N_2027,N_2589);
and U3495 (N_3495,N_2111,N_2840);
nor U3496 (N_3496,N_2994,N_2696);
nor U3497 (N_3497,N_2440,N_2254);
nand U3498 (N_3498,N_2635,N_2499);
and U3499 (N_3499,N_2283,N_2631);
or U3500 (N_3500,N_2732,N_2286);
nor U3501 (N_3501,N_2372,N_2259);
and U3502 (N_3502,N_2051,N_2337);
or U3503 (N_3503,N_2037,N_2266);
and U3504 (N_3504,N_2548,N_2614);
and U3505 (N_3505,N_2822,N_2459);
and U3506 (N_3506,N_2851,N_2229);
nand U3507 (N_3507,N_2091,N_2514);
nor U3508 (N_3508,N_2549,N_2541);
nor U3509 (N_3509,N_2132,N_2723);
nor U3510 (N_3510,N_2197,N_2740);
or U3511 (N_3511,N_2630,N_2842);
or U3512 (N_3512,N_2594,N_2212);
or U3513 (N_3513,N_2260,N_2437);
nand U3514 (N_3514,N_2898,N_2788);
xnor U3515 (N_3515,N_2120,N_2678);
xor U3516 (N_3516,N_2339,N_2869);
or U3517 (N_3517,N_2249,N_2334);
or U3518 (N_3518,N_2468,N_2832);
nand U3519 (N_3519,N_2669,N_2706);
and U3520 (N_3520,N_2980,N_2180);
nor U3521 (N_3521,N_2357,N_2556);
or U3522 (N_3522,N_2326,N_2495);
xnor U3523 (N_3523,N_2763,N_2973);
xnor U3524 (N_3524,N_2335,N_2640);
nand U3525 (N_3525,N_2491,N_2687);
and U3526 (N_3526,N_2905,N_2211);
nand U3527 (N_3527,N_2527,N_2921);
or U3528 (N_3528,N_2265,N_2559);
nand U3529 (N_3529,N_2039,N_2916);
nor U3530 (N_3530,N_2896,N_2631);
or U3531 (N_3531,N_2320,N_2717);
xnor U3532 (N_3532,N_2920,N_2142);
or U3533 (N_3533,N_2792,N_2650);
nand U3534 (N_3534,N_2044,N_2051);
and U3535 (N_3535,N_2860,N_2410);
nand U3536 (N_3536,N_2712,N_2480);
or U3537 (N_3537,N_2069,N_2070);
and U3538 (N_3538,N_2365,N_2183);
or U3539 (N_3539,N_2733,N_2703);
or U3540 (N_3540,N_2586,N_2692);
and U3541 (N_3541,N_2167,N_2923);
nand U3542 (N_3542,N_2967,N_2935);
and U3543 (N_3543,N_2758,N_2295);
nor U3544 (N_3544,N_2415,N_2803);
or U3545 (N_3545,N_2248,N_2828);
nand U3546 (N_3546,N_2690,N_2240);
xor U3547 (N_3547,N_2689,N_2040);
nor U3548 (N_3548,N_2610,N_2336);
or U3549 (N_3549,N_2533,N_2662);
nor U3550 (N_3550,N_2309,N_2624);
nor U3551 (N_3551,N_2647,N_2591);
nand U3552 (N_3552,N_2524,N_2838);
and U3553 (N_3553,N_2772,N_2493);
nor U3554 (N_3554,N_2479,N_2656);
or U3555 (N_3555,N_2505,N_2834);
and U3556 (N_3556,N_2777,N_2247);
or U3557 (N_3557,N_2554,N_2343);
or U3558 (N_3558,N_2209,N_2153);
nand U3559 (N_3559,N_2967,N_2293);
nor U3560 (N_3560,N_2411,N_2272);
or U3561 (N_3561,N_2084,N_2530);
nor U3562 (N_3562,N_2078,N_2284);
xor U3563 (N_3563,N_2570,N_2876);
or U3564 (N_3564,N_2762,N_2976);
nor U3565 (N_3565,N_2231,N_2710);
and U3566 (N_3566,N_2642,N_2059);
and U3567 (N_3567,N_2377,N_2425);
xnor U3568 (N_3568,N_2363,N_2707);
nor U3569 (N_3569,N_2190,N_2816);
nor U3570 (N_3570,N_2353,N_2205);
xor U3571 (N_3571,N_2118,N_2783);
xor U3572 (N_3572,N_2012,N_2423);
or U3573 (N_3573,N_2573,N_2996);
or U3574 (N_3574,N_2695,N_2454);
or U3575 (N_3575,N_2543,N_2301);
nor U3576 (N_3576,N_2648,N_2172);
or U3577 (N_3577,N_2883,N_2639);
nand U3578 (N_3578,N_2941,N_2093);
or U3579 (N_3579,N_2046,N_2827);
nand U3580 (N_3580,N_2925,N_2627);
nand U3581 (N_3581,N_2784,N_2609);
or U3582 (N_3582,N_2857,N_2790);
nand U3583 (N_3583,N_2553,N_2104);
nand U3584 (N_3584,N_2740,N_2923);
and U3585 (N_3585,N_2196,N_2015);
and U3586 (N_3586,N_2218,N_2539);
or U3587 (N_3587,N_2017,N_2007);
or U3588 (N_3588,N_2076,N_2530);
nor U3589 (N_3589,N_2677,N_2159);
or U3590 (N_3590,N_2803,N_2352);
and U3591 (N_3591,N_2298,N_2037);
nand U3592 (N_3592,N_2202,N_2349);
nor U3593 (N_3593,N_2155,N_2909);
or U3594 (N_3594,N_2038,N_2257);
xnor U3595 (N_3595,N_2219,N_2530);
nor U3596 (N_3596,N_2062,N_2439);
nand U3597 (N_3597,N_2813,N_2304);
xor U3598 (N_3598,N_2673,N_2433);
xnor U3599 (N_3599,N_2481,N_2673);
or U3600 (N_3600,N_2941,N_2649);
nand U3601 (N_3601,N_2103,N_2622);
nand U3602 (N_3602,N_2334,N_2551);
nand U3603 (N_3603,N_2304,N_2743);
nor U3604 (N_3604,N_2103,N_2066);
nand U3605 (N_3605,N_2031,N_2067);
nor U3606 (N_3606,N_2011,N_2808);
or U3607 (N_3607,N_2526,N_2402);
or U3608 (N_3608,N_2255,N_2773);
and U3609 (N_3609,N_2828,N_2960);
and U3610 (N_3610,N_2394,N_2739);
or U3611 (N_3611,N_2841,N_2198);
and U3612 (N_3612,N_2990,N_2500);
nand U3613 (N_3613,N_2784,N_2728);
xor U3614 (N_3614,N_2547,N_2407);
nand U3615 (N_3615,N_2380,N_2865);
xor U3616 (N_3616,N_2263,N_2622);
nand U3617 (N_3617,N_2060,N_2962);
and U3618 (N_3618,N_2384,N_2228);
xnor U3619 (N_3619,N_2025,N_2700);
and U3620 (N_3620,N_2201,N_2702);
xor U3621 (N_3621,N_2231,N_2714);
and U3622 (N_3622,N_2063,N_2014);
nor U3623 (N_3623,N_2726,N_2147);
xnor U3624 (N_3624,N_2461,N_2498);
and U3625 (N_3625,N_2571,N_2391);
nor U3626 (N_3626,N_2460,N_2768);
nor U3627 (N_3627,N_2416,N_2570);
or U3628 (N_3628,N_2554,N_2842);
nand U3629 (N_3629,N_2695,N_2836);
xor U3630 (N_3630,N_2648,N_2545);
nor U3631 (N_3631,N_2449,N_2751);
nand U3632 (N_3632,N_2406,N_2733);
nor U3633 (N_3633,N_2475,N_2154);
nor U3634 (N_3634,N_2606,N_2372);
nand U3635 (N_3635,N_2872,N_2344);
nand U3636 (N_3636,N_2657,N_2426);
nand U3637 (N_3637,N_2398,N_2222);
and U3638 (N_3638,N_2645,N_2169);
and U3639 (N_3639,N_2972,N_2948);
nand U3640 (N_3640,N_2050,N_2574);
or U3641 (N_3641,N_2256,N_2236);
and U3642 (N_3642,N_2756,N_2690);
and U3643 (N_3643,N_2397,N_2704);
nor U3644 (N_3644,N_2736,N_2045);
nand U3645 (N_3645,N_2585,N_2249);
xnor U3646 (N_3646,N_2799,N_2695);
nand U3647 (N_3647,N_2362,N_2067);
nand U3648 (N_3648,N_2696,N_2243);
xnor U3649 (N_3649,N_2351,N_2570);
nor U3650 (N_3650,N_2712,N_2262);
nor U3651 (N_3651,N_2028,N_2603);
nor U3652 (N_3652,N_2295,N_2162);
or U3653 (N_3653,N_2259,N_2147);
and U3654 (N_3654,N_2361,N_2073);
and U3655 (N_3655,N_2219,N_2270);
or U3656 (N_3656,N_2237,N_2383);
or U3657 (N_3657,N_2735,N_2529);
nand U3658 (N_3658,N_2033,N_2247);
nor U3659 (N_3659,N_2827,N_2081);
nor U3660 (N_3660,N_2691,N_2733);
nor U3661 (N_3661,N_2392,N_2329);
nor U3662 (N_3662,N_2846,N_2229);
and U3663 (N_3663,N_2898,N_2464);
nand U3664 (N_3664,N_2796,N_2047);
nand U3665 (N_3665,N_2447,N_2113);
and U3666 (N_3666,N_2792,N_2395);
xnor U3667 (N_3667,N_2118,N_2495);
or U3668 (N_3668,N_2346,N_2549);
and U3669 (N_3669,N_2617,N_2915);
nand U3670 (N_3670,N_2642,N_2516);
nor U3671 (N_3671,N_2081,N_2134);
nor U3672 (N_3672,N_2477,N_2348);
xor U3673 (N_3673,N_2053,N_2925);
or U3674 (N_3674,N_2082,N_2902);
nor U3675 (N_3675,N_2107,N_2956);
or U3676 (N_3676,N_2655,N_2487);
and U3677 (N_3677,N_2873,N_2885);
or U3678 (N_3678,N_2127,N_2869);
nand U3679 (N_3679,N_2747,N_2563);
nand U3680 (N_3680,N_2478,N_2707);
and U3681 (N_3681,N_2847,N_2625);
or U3682 (N_3682,N_2571,N_2512);
and U3683 (N_3683,N_2566,N_2005);
nor U3684 (N_3684,N_2999,N_2000);
and U3685 (N_3685,N_2718,N_2873);
or U3686 (N_3686,N_2791,N_2157);
and U3687 (N_3687,N_2731,N_2287);
or U3688 (N_3688,N_2958,N_2551);
nand U3689 (N_3689,N_2378,N_2422);
nor U3690 (N_3690,N_2438,N_2509);
and U3691 (N_3691,N_2486,N_2256);
and U3692 (N_3692,N_2568,N_2463);
nor U3693 (N_3693,N_2789,N_2089);
nand U3694 (N_3694,N_2159,N_2570);
nand U3695 (N_3695,N_2576,N_2797);
nand U3696 (N_3696,N_2269,N_2859);
and U3697 (N_3697,N_2002,N_2212);
and U3698 (N_3698,N_2784,N_2559);
xor U3699 (N_3699,N_2682,N_2216);
or U3700 (N_3700,N_2173,N_2388);
or U3701 (N_3701,N_2799,N_2257);
and U3702 (N_3702,N_2621,N_2634);
nand U3703 (N_3703,N_2655,N_2065);
nand U3704 (N_3704,N_2651,N_2969);
and U3705 (N_3705,N_2743,N_2025);
nand U3706 (N_3706,N_2756,N_2769);
nor U3707 (N_3707,N_2095,N_2984);
or U3708 (N_3708,N_2151,N_2507);
and U3709 (N_3709,N_2819,N_2874);
or U3710 (N_3710,N_2934,N_2634);
nand U3711 (N_3711,N_2907,N_2299);
xnor U3712 (N_3712,N_2227,N_2596);
nand U3713 (N_3713,N_2539,N_2785);
and U3714 (N_3714,N_2334,N_2095);
xnor U3715 (N_3715,N_2751,N_2115);
nor U3716 (N_3716,N_2359,N_2819);
nor U3717 (N_3717,N_2564,N_2641);
nand U3718 (N_3718,N_2249,N_2030);
and U3719 (N_3719,N_2461,N_2514);
nor U3720 (N_3720,N_2982,N_2541);
nand U3721 (N_3721,N_2466,N_2299);
xnor U3722 (N_3722,N_2197,N_2170);
nor U3723 (N_3723,N_2523,N_2594);
or U3724 (N_3724,N_2267,N_2764);
and U3725 (N_3725,N_2545,N_2774);
nand U3726 (N_3726,N_2423,N_2917);
nand U3727 (N_3727,N_2736,N_2494);
and U3728 (N_3728,N_2770,N_2666);
and U3729 (N_3729,N_2093,N_2597);
xnor U3730 (N_3730,N_2705,N_2766);
nor U3731 (N_3731,N_2517,N_2314);
nor U3732 (N_3732,N_2153,N_2219);
and U3733 (N_3733,N_2019,N_2680);
nand U3734 (N_3734,N_2080,N_2382);
or U3735 (N_3735,N_2288,N_2248);
nor U3736 (N_3736,N_2045,N_2754);
nand U3737 (N_3737,N_2483,N_2650);
and U3738 (N_3738,N_2682,N_2028);
nor U3739 (N_3739,N_2399,N_2946);
nand U3740 (N_3740,N_2645,N_2498);
nand U3741 (N_3741,N_2911,N_2284);
nand U3742 (N_3742,N_2893,N_2261);
and U3743 (N_3743,N_2227,N_2499);
and U3744 (N_3744,N_2086,N_2766);
and U3745 (N_3745,N_2638,N_2446);
nand U3746 (N_3746,N_2735,N_2158);
or U3747 (N_3747,N_2899,N_2422);
and U3748 (N_3748,N_2655,N_2680);
or U3749 (N_3749,N_2671,N_2356);
and U3750 (N_3750,N_2094,N_2607);
nor U3751 (N_3751,N_2839,N_2895);
or U3752 (N_3752,N_2645,N_2187);
and U3753 (N_3753,N_2277,N_2969);
nor U3754 (N_3754,N_2937,N_2264);
nor U3755 (N_3755,N_2393,N_2905);
nand U3756 (N_3756,N_2532,N_2865);
nand U3757 (N_3757,N_2750,N_2080);
nor U3758 (N_3758,N_2729,N_2968);
and U3759 (N_3759,N_2622,N_2176);
nand U3760 (N_3760,N_2497,N_2549);
nor U3761 (N_3761,N_2883,N_2002);
and U3762 (N_3762,N_2634,N_2017);
and U3763 (N_3763,N_2363,N_2883);
or U3764 (N_3764,N_2168,N_2148);
nand U3765 (N_3765,N_2393,N_2910);
nor U3766 (N_3766,N_2035,N_2316);
or U3767 (N_3767,N_2398,N_2665);
or U3768 (N_3768,N_2659,N_2222);
nand U3769 (N_3769,N_2026,N_2555);
nor U3770 (N_3770,N_2996,N_2474);
and U3771 (N_3771,N_2978,N_2821);
and U3772 (N_3772,N_2875,N_2269);
nor U3773 (N_3773,N_2476,N_2378);
nor U3774 (N_3774,N_2661,N_2118);
xor U3775 (N_3775,N_2802,N_2390);
and U3776 (N_3776,N_2523,N_2956);
and U3777 (N_3777,N_2605,N_2396);
or U3778 (N_3778,N_2011,N_2208);
nand U3779 (N_3779,N_2062,N_2948);
and U3780 (N_3780,N_2233,N_2239);
and U3781 (N_3781,N_2072,N_2348);
xor U3782 (N_3782,N_2881,N_2978);
or U3783 (N_3783,N_2088,N_2136);
and U3784 (N_3784,N_2215,N_2515);
or U3785 (N_3785,N_2605,N_2637);
xor U3786 (N_3786,N_2220,N_2829);
or U3787 (N_3787,N_2458,N_2494);
or U3788 (N_3788,N_2138,N_2531);
nand U3789 (N_3789,N_2819,N_2917);
or U3790 (N_3790,N_2188,N_2079);
nand U3791 (N_3791,N_2054,N_2656);
nand U3792 (N_3792,N_2650,N_2964);
nand U3793 (N_3793,N_2721,N_2292);
and U3794 (N_3794,N_2048,N_2584);
or U3795 (N_3795,N_2865,N_2447);
and U3796 (N_3796,N_2323,N_2193);
nand U3797 (N_3797,N_2053,N_2451);
nand U3798 (N_3798,N_2497,N_2125);
and U3799 (N_3799,N_2228,N_2006);
nor U3800 (N_3800,N_2710,N_2743);
and U3801 (N_3801,N_2176,N_2026);
nor U3802 (N_3802,N_2447,N_2074);
and U3803 (N_3803,N_2086,N_2275);
nand U3804 (N_3804,N_2737,N_2146);
and U3805 (N_3805,N_2580,N_2691);
or U3806 (N_3806,N_2986,N_2108);
or U3807 (N_3807,N_2471,N_2060);
and U3808 (N_3808,N_2070,N_2905);
and U3809 (N_3809,N_2370,N_2929);
and U3810 (N_3810,N_2009,N_2624);
xnor U3811 (N_3811,N_2630,N_2368);
or U3812 (N_3812,N_2001,N_2855);
and U3813 (N_3813,N_2794,N_2695);
xnor U3814 (N_3814,N_2935,N_2276);
and U3815 (N_3815,N_2704,N_2104);
nor U3816 (N_3816,N_2172,N_2205);
nand U3817 (N_3817,N_2959,N_2383);
and U3818 (N_3818,N_2777,N_2119);
xnor U3819 (N_3819,N_2354,N_2209);
or U3820 (N_3820,N_2750,N_2655);
or U3821 (N_3821,N_2533,N_2885);
and U3822 (N_3822,N_2420,N_2720);
and U3823 (N_3823,N_2271,N_2341);
nor U3824 (N_3824,N_2820,N_2660);
nor U3825 (N_3825,N_2208,N_2445);
or U3826 (N_3826,N_2372,N_2708);
and U3827 (N_3827,N_2187,N_2827);
or U3828 (N_3828,N_2705,N_2648);
nor U3829 (N_3829,N_2658,N_2179);
or U3830 (N_3830,N_2844,N_2550);
nand U3831 (N_3831,N_2124,N_2091);
nand U3832 (N_3832,N_2368,N_2504);
and U3833 (N_3833,N_2009,N_2247);
nand U3834 (N_3834,N_2388,N_2679);
xnor U3835 (N_3835,N_2667,N_2801);
nor U3836 (N_3836,N_2171,N_2383);
nand U3837 (N_3837,N_2498,N_2545);
nor U3838 (N_3838,N_2387,N_2398);
xnor U3839 (N_3839,N_2239,N_2278);
and U3840 (N_3840,N_2997,N_2249);
nor U3841 (N_3841,N_2281,N_2862);
and U3842 (N_3842,N_2668,N_2478);
and U3843 (N_3843,N_2249,N_2932);
or U3844 (N_3844,N_2096,N_2256);
and U3845 (N_3845,N_2300,N_2081);
nor U3846 (N_3846,N_2035,N_2326);
nor U3847 (N_3847,N_2311,N_2424);
nand U3848 (N_3848,N_2648,N_2451);
nor U3849 (N_3849,N_2033,N_2044);
nor U3850 (N_3850,N_2541,N_2339);
nand U3851 (N_3851,N_2333,N_2979);
nor U3852 (N_3852,N_2963,N_2488);
nor U3853 (N_3853,N_2184,N_2798);
nand U3854 (N_3854,N_2462,N_2289);
nand U3855 (N_3855,N_2820,N_2893);
nand U3856 (N_3856,N_2930,N_2998);
and U3857 (N_3857,N_2533,N_2056);
and U3858 (N_3858,N_2232,N_2899);
or U3859 (N_3859,N_2693,N_2440);
xnor U3860 (N_3860,N_2976,N_2717);
or U3861 (N_3861,N_2610,N_2480);
xnor U3862 (N_3862,N_2337,N_2219);
nand U3863 (N_3863,N_2289,N_2071);
and U3864 (N_3864,N_2415,N_2019);
xnor U3865 (N_3865,N_2580,N_2027);
nor U3866 (N_3866,N_2909,N_2308);
nand U3867 (N_3867,N_2307,N_2474);
xor U3868 (N_3868,N_2101,N_2794);
nand U3869 (N_3869,N_2188,N_2660);
or U3870 (N_3870,N_2803,N_2185);
or U3871 (N_3871,N_2457,N_2426);
and U3872 (N_3872,N_2551,N_2221);
and U3873 (N_3873,N_2845,N_2514);
and U3874 (N_3874,N_2542,N_2556);
nand U3875 (N_3875,N_2329,N_2937);
or U3876 (N_3876,N_2963,N_2521);
nand U3877 (N_3877,N_2965,N_2056);
or U3878 (N_3878,N_2072,N_2313);
or U3879 (N_3879,N_2062,N_2908);
and U3880 (N_3880,N_2999,N_2528);
or U3881 (N_3881,N_2273,N_2903);
xor U3882 (N_3882,N_2566,N_2739);
or U3883 (N_3883,N_2172,N_2649);
or U3884 (N_3884,N_2613,N_2048);
nand U3885 (N_3885,N_2839,N_2719);
or U3886 (N_3886,N_2229,N_2759);
nand U3887 (N_3887,N_2962,N_2330);
or U3888 (N_3888,N_2042,N_2284);
and U3889 (N_3889,N_2931,N_2259);
and U3890 (N_3890,N_2535,N_2091);
or U3891 (N_3891,N_2450,N_2876);
or U3892 (N_3892,N_2065,N_2193);
xor U3893 (N_3893,N_2309,N_2306);
or U3894 (N_3894,N_2327,N_2794);
nor U3895 (N_3895,N_2336,N_2968);
nand U3896 (N_3896,N_2474,N_2730);
nor U3897 (N_3897,N_2357,N_2410);
xnor U3898 (N_3898,N_2245,N_2833);
and U3899 (N_3899,N_2318,N_2954);
nor U3900 (N_3900,N_2757,N_2629);
nor U3901 (N_3901,N_2369,N_2314);
xor U3902 (N_3902,N_2396,N_2010);
and U3903 (N_3903,N_2213,N_2151);
nand U3904 (N_3904,N_2967,N_2614);
and U3905 (N_3905,N_2424,N_2702);
or U3906 (N_3906,N_2268,N_2796);
nor U3907 (N_3907,N_2154,N_2231);
nand U3908 (N_3908,N_2207,N_2180);
or U3909 (N_3909,N_2925,N_2534);
and U3910 (N_3910,N_2500,N_2864);
nand U3911 (N_3911,N_2432,N_2291);
nand U3912 (N_3912,N_2133,N_2276);
nand U3913 (N_3913,N_2720,N_2476);
or U3914 (N_3914,N_2854,N_2927);
nor U3915 (N_3915,N_2644,N_2618);
and U3916 (N_3916,N_2823,N_2388);
nor U3917 (N_3917,N_2318,N_2806);
nor U3918 (N_3918,N_2851,N_2544);
and U3919 (N_3919,N_2255,N_2850);
nand U3920 (N_3920,N_2101,N_2076);
and U3921 (N_3921,N_2440,N_2102);
and U3922 (N_3922,N_2489,N_2905);
nand U3923 (N_3923,N_2158,N_2298);
nor U3924 (N_3924,N_2122,N_2405);
nor U3925 (N_3925,N_2362,N_2259);
xor U3926 (N_3926,N_2772,N_2323);
nor U3927 (N_3927,N_2713,N_2463);
nand U3928 (N_3928,N_2404,N_2661);
nand U3929 (N_3929,N_2929,N_2978);
nand U3930 (N_3930,N_2733,N_2584);
xor U3931 (N_3931,N_2066,N_2293);
or U3932 (N_3932,N_2965,N_2951);
nor U3933 (N_3933,N_2621,N_2137);
nand U3934 (N_3934,N_2458,N_2712);
nand U3935 (N_3935,N_2643,N_2988);
nand U3936 (N_3936,N_2120,N_2254);
or U3937 (N_3937,N_2350,N_2234);
nand U3938 (N_3938,N_2993,N_2052);
xor U3939 (N_3939,N_2148,N_2987);
nor U3940 (N_3940,N_2917,N_2651);
xnor U3941 (N_3941,N_2114,N_2213);
nor U3942 (N_3942,N_2843,N_2188);
and U3943 (N_3943,N_2798,N_2324);
nand U3944 (N_3944,N_2249,N_2342);
nor U3945 (N_3945,N_2957,N_2633);
xor U3946 (N_3946,N_2119,N_2859);
and U3947 (N_3947,N_2117,N_2166);
or U3948 (N_3948,N_2731,N_2146);
or U3949 (N_3949,N_2080,N_2050);
and U3950 (N_3950,N_2896,N_2894);
nand U3951 (N_3951,N_2835,N_2263);
and U3952 (N_3952,N_2679,N_2727);
and U3953 (N_3953,N_2074,N_2472);
and U3954 (N_3954,N_2206,N_2091);
nand U3955 (N_3955,N_2832,N_2427);
nor U3956 (N_3956,N_2679,N_2084);
and U3957 (N_3957,N_2473,N_2839);
nand U3958 (N_3958,N_2244,N_2900);
and U3959 (N_3959,N_2732,N_2098);
or U3960 (N_3960,N_2998,N_2008);
and U3961 (N_3961,N_2938,N_2979);
nor U3962 (N_3962,N_2067,N_2141);
nor U3963 (N_3963,N_2737,N_2841);
nor U3964 (N_3964,N_2376,N_2433);
or U3965 (N_3965,N_2706,N_2220);
nand U3966 (N_3966,N_2560,N_2294);
and U3967 (N_3967,N_2719,N_2251);
nand U3968 (N_3968,N_2285,N_2196);
or U3969 (N_3969,N_2855,N_2472);
or U3970 (N_3970,N_2508,N_2910);
nor U3971 (N_3971,N_2963,N_2160);
or U3972 (N_3972,N_2706,N_2683);
nor U3973 (N_3973,N_2402,N_2569);
and U3974 (N_3974,N_2712,N_2512);
or U3975 (N_3975,N_2430,N_2526);
nand U3976 (N_3976,N_2454,N_2935);
and U3977 (N_3977,N_2197,N_2054);
nor U3978 (N_3978,N_2079,N_2722);
nand U3979 (N_3979,N_2257,N_2327);
nor U3980 (N_3980,N_2542,N_2847);
or U3981 (N_3981,N_2539,N_2856);
and U3982 (N_3982,N_2229,N_2385);
nand U3983 (N_3983,N_2680,N_2170);
nand U3984 (N_3984,N_2054,N_2328);
and U3985 (N_3985,N_2900,N_2890);
or U3986 (N_3986,N_2523,N_2512);
and U3987 (N_3987,N_2716,N_2165);
and U3988 (N_3988,N_2674,N_2633);
or U3989 (N_3989,N_2841,N_2576);
nand U3990 (N_3990,N_2908,N_2564);
nand U3991 (N_3991,N_2383,N_2567);
or U3992 (N_3992,N_2987,N_2109);
nor U3993 (N_3993,N_2422,N_2224);
and U3994 (N_3994,N_2912,N_2376);
nor U3995 (N_3995,N_2058,N_2322);
or U3996 (N_3996,N_2339,N_2537);
nand U3997 (N_3997,N_2941,N_2402);
xor U3998 (N_3998,N_2263,N_2597);
nor U3999 (N_3999,N_2159,N_2834);
nand U4000 (N_4000,N_3680,N_3091);
nor U4001 (N_4001,N_3872,N_3499);
nor U4002 (N_4002,N_3697,N_3899);
nor U4003 (N_4003,N_3967,N_3730);
or U4004 (N_4004,N_3287,N_3609);
nand U4005 (N_4005,N_3992,N_3192);
and U4006 (N_4006,N_3475,N_3310);
nor U4007 (N_4007,N_3957,N_3322);
or U4008 (N_4008,N_3031,N_3525);
nor U4009 (N_4009,N_3465,N_3646);
nor U4010 (N_4010,N_3043,N_3877);
or U4011 (N_4011,N_3921,N_3330);
and U4012 (N_4012,N_3253,N_3364);
xnor U4013 (N_4013,N_3267,N_3035);
xnor U4014 (N_4014,N_3559,N_3344);
xor U4015 (N_4015,N_3599,N_3666);
and U4016 (N_4016,N_3954,N_3760);
nor U4017 (N_4017,N_3911,N_3889);
xnor U4018 (N_4018,N_3713,N_3504);
nor U4019 (N_4019,N_3434,N_3359);
nand U4020 (N_4020,N_3819,N_3397);
nand U4021 (N_4021,N_3928,N_3789);
nand U4022 (N_4022,N_3802,N_3386);
or U4023 (N_4023,N_3486,N_3809);
xor U4024 (N_4024,N_3065,N_3903);
nor U4025 (N_4025,N_3976,N_3729);
nor U4026 (N_4026,N_3027,N_3966);
or U4027 (N_4027,N_3868,N_3707);
nand U4028 (N_4028,N_3356,N_3949);
or U4029 (N_4029,N_3279,N_3180);
or U4030 (N_4030,N_3781,N_3573);
xnor U4031 (N_4031,N_3764,N_3214);
nor U4032 (N_4032,N_3178,N_3564);
or U4033 (N_4033,N_3830,N_3661);
or U4034 (N_4034,N_3672,N_3053);
nor U4035 (N_4035,N_3880,N_3400);
nand U4036 (N_4036,N_3191,N_3312);
or U4037 (N_4037,N_3775,N_3745);
or U4038 (N_4038,N_3807,N_3329);
nor U4039 (N_4039,N_3207,N_3102);
nor U4040 (N_4040,N_3469,N_3510);
xnor U4041 (N_4041,N_3528,N_3358);
nand U4042 (N_4042,N_3700,N_3141);
nand U4043 (N_4043,N_3530,N_3398);
or U4044 (N_4044,N_3686,N_3962);
nor U4045 (N_4045,N_3032,N_3020);
nor U4046 (N_4046,N_3431,N_3218);
nand U4047 (N_4047,N_3624,N_3127);
and U4048 (N_4048,N_3704,N_3139);
nor U4049 (N_4049,N_3580,N_3822);
nand U4050 (N_4050,N_3457,N_3814);
or U4051 (N_4051,N_3154,N_3313);
or U4052 (N_4052,N_3806,N_3343);
and U4053 (N_4053,N_3682,N_3912);
xor U4054 (N_4054,N_3447,N_3059);
nor U4055 (N_4055,N_3800,N_3701);
xnor U4056 (N_4056,N_3754,N_3288);
nor U4057 (N_4057,N_3289,N_3519);
and U4058 (N_4058,N_3346,N_3078);
nor U4059 (N_4059,N_3402,N_3524);
and U4060 (N_4060,N_3710,N_3569);
and U4061 (N_4061,N_3222,N_3349);
or U4062 (N_4062,N_3621,N_3792);
and U4063 (N_4063,N_3847,N_3454);
nand U4064 (N_4064,N_3058,N_3732);
nor U4065 (N_4065,N_3805,N_3037);
or U4066 (N_4066,N_3523,N_3147);
xnor U4067 (N_4067,N_3747,N_3614);
nand U4068 (N_4068,N_3981,N_3296);
nand U4069 (N_4069,N_3015,N_3901);
or U4070 (N_4070,N_3369,N_3810);
or U4071 (N_4071,N_3379,N_3837);
nand U4072 (N_4072,N_3136,N_3227);
and U4073 (N_4073,N_3278,N_3190);
or U4074 (N_4074,N_3104,N_3458);
and U4075 (N_4075,N_3452,N_3739);
nor U4076 (N_4076,N_3615,N_3488);
or U4077 (N_4077,N_3874,N_3639);
and U4078 (N_4078,N_3994,N_3224);
nand U4079 (N_4079,N_3892,N_3007);
or U4080 (N_4080,N_3759,N_3772);
nand U4081 (N_4081,N_3121,N_3202);
and U4082 (N_4082,N_3778,N_3385);
nand U4083 (N_4083,N_3768,N_3156);
or U4084 (N_4084,N_3886,N_3719);
or U4085 (N_4085,N_3572,N_3155);
or U4086 (N_4086,N_3665,N_3753);
xor U4087 (N_4087,N_3861,N_3327);
or U4088 (N_4088,N_3542,N_3252);
nand U4089 (N_4089,N_3758,N_3446);
and U4090 (N_4090,N_3917,N_3036);
or U4091 (N_4091,N_3087,N_3437);
and U4092 (N_4092,N_3675,N_3604);
and U4093 (N_4093,N_3487,N_3770);
nor U4094 (N_4094,N_3424,N_3555);
xor U4095 (N_4095,N_3384,N_3211);
nor U4096 (N_4096,N_3898,N_3855);
and U4097 (N_4097,N_3471,N_3265);
and U4098 (N_4098,N_3698,N_3926);
nor U4099 (N_4099,N_3652,N_3984);
and U4100 (N_4100,N_3688,N_3785);
and U4101 (N_4101,N_3750,N_3858);
and U4102 (N_4102,N_3380,N_3915);
nor U4103 (N_4103,N_3137,N_3435);
nor U4104 (N_4104,N_3683,N_3902);
nand U4105 (N_4105,N_3163,N_3071);
nand U4106 (N_4106,N_3206,N_3244);
and U4107 (N_4107,N_3923,N_3009);
nor U4108 (N_4108,N_3060,N_3250);
or U4109 (N_4109,N_3410,N_3010);
and U4110 (N_4110,N_3149,N_3423);
nand U4111 (N_4111,N_3134,N_3570);
nor U4112 (N_4112,N_3742,N_3464);
nor U4113 (N_4113,N_3674,N_3721);
or U4114 (N_4114,N_3838,N_3221);
nor U4115 (N_4115,N_3692,N_3044);
nand U4116 (N_4116,N_3520,N_3272);
nand U4117 (N_4117,N_3895,N_3997);
and U4118 (N_4118,N_3918,N_3930);
and U4119 (N_4119,N_3425,N_3537);
nand U4120 (N_4120,N_3762,N_3378);
and U4121 (N_4121,N_3647,N_3000);
xor U4122 (N_4122,N_3394,N_3268);
or U4123 (N_4123,N_3187,N_3611);
and U4124 (N_4124,N_3333,N_3427);
nor U4125 (N_4125,N_3245,N_3170);
and U4126 (N_4126,N_3428,N_3029);
and U4127 (N_4127,N_3399,N_3413);
or U4128 (N_4128,N_3687,N_3374);
or U4129 (N_4129,N_3406,N_3857);
nor U4130 (N_4130,N_3421,N_3888);
nand U4131 (N_4131,N_3086,N_3633);
xnor U4132 (N_4132,N_3130,N_3973);
xnor U4133 (N_4133,N_3543,N_3936);
nand U4134 (N_4134,N_3718,N_3634);
and U4135 (N_4135,N_3303,N_3812);
nand U4136 (N_4136,N_3547,N_3073);
or U4137 (N_4137,N_3390,N_3168);
nor U4138 (N_4138,N_3376,N_3144);
xor U4139 (N_4139,N_3350,N_3238);
or U4140 (N_4140,N_3587,N_3642);
or U4141 (N_4141,N_3117,N_3695);
and U4142 (N_4142,N_3392,N_3175);
nand U4143 (N_4143,N_3567,N_3324);
or U4144 (N_4144,N_3591,N_3975);
or U4145 (N_4145,N_3255,N_3140);
or U4146 (N_4146,N_3685,N_3019);
nor U4147 (N_4147,N_3012,N_3022);
and U4148 (N_4148,N_3630,N_3625);
or U4149 (N_4149,N_3662,N_3260);
nor U4150 (N_4150,N_3028,N_3408);
and U4151 (N_4151,N_3950,N_3948);
nand U4152 (N_4152,N_3212,N_3516);
xnor U4153 (N_4153,N_3724,N_3450);
or U4154 (N_4154,N_3182,N_3919);
nand U4155 (N_4155,N_3723,N_3199);
nand U4156 (N_4156,N_3321,N_3714);
nor U4157 (N_4157,N_3635,N_3365);
or U4158 (N_4158,N_3002,N_3595);
xor U4159 (N_4159,N_3722,N_3920);
nand U4160 (N_4160,N_3944,N_3460);
nand U4161 (N_4161,N_3148,N_3033);
and U4162 (N_4162,N_3852,N_3859);
xor U4163 (N_4163,N_3512,N_3231);
nor U4164 (N_4164,N_3645,N_3856);
or U4165 (N_4165,N_3051,N_3257);
and U4166 (N_4166,N_3203,N_3699);
xor U4167 (N_4167,N_3799,N_3362);
nor U4168 (N_4168,N_3924,N_3042);
or U4169 (N_4169,N_3644,N_3720);
xor U4170 (N_4170,N_3293,N_3318);
nor U4171 (N_4171,N_3054,N_3101);
nand U4172 (N_4172,N_3617,N_3913);
and U4173 (N_4173,N_3068,N_3968);
nand U4174 (N_4174,N_3473,N_3081);
nor U4175 (N_4175,N_3125,N_3334);
or U4176 (N_4176,N_3932,N_3395);
nand U4177 (N_4177,N_3416,N_3643);
nand U4178 (N_4178,N_3440,N_3709);
nand U4179 (N_4179,N_3072,N_3097);
and U4180 (N_4180,N_3828,N_3654);
nor U4181 (N_4181,N_3790,N_3640);
nand U4182 (N_4182,N_3582,N_3368);
or U4183 (N_4183,N_3039,N_3439);
nand U4184 (N_4184,N_3773,N_3438);
and U4185 (N_4185,N_3167,N_3574);
or U4186 (N_4186,N_3561,N_3734);
nand U4187 (N_4187,N_3453,N_3953);
and U4188 (N_4188,N_3534,N_3109);
nand U4189 (N_4189,N_3174,N_3468);
and U4190 (N_4190,N_3933,N_3788);
or U4191 (N_4191,N_3660,N_3993);
nand U4192 (N_4192,N_3301,N_3114);
xor U4193 (N_4193,N_3251,N_3879);
and U4194 (N_4194,N_3355,N_3648);
nand U4195 (N_4195,N_3526,N_3793);
nor U4196 (N_4196,N_3726,N_3490);
nand U4197 (N_4197,N_3162,N_3223);
and U4198 (N_4198,N_3177,N_3825);
and U4199 (N_4199,N_3636,N_3878);
nand U4200 (N_4200,N_3340,N_3196);
nand U4201 (N_4201,N_3655,N_3373);
xor U4202 (N_4202,N_3588,N_3205);
and U4203 (N_4203,N_3215,N_3483);
nand U4204 (N_4204,N_3011,N_3885);
nor U4205 (N_4205,N_3779,N_3466);
and U4206 (N_4206,N_3910,N_3744);
nand U4207 (N_4207,N_3405,N_3098);
xor U4208 (N_4208,N_3835,N_3099);
nand U4209 (N_4209,N_3094,N_3583);
nor U4210 (N_4210,N_3864,N_3095);
or U4211 (N_4211,N_3733,N_3232);
xnor U4212 (N_4212,N_3315,N_3332);
nand U4213 (N_4213,N_3598,N_3089);
nand U4214 (N_4214,N_3618,N_3706);
nand U4215 (N_4215,N_3083,N_3943);
or U4216 (N_4216,N_3725,N_3608);
or U4217 (N_4217,N_3767,N_3908);
or U4218 (N_4218,N_3791,N_3357);
and U4219 (N_4219,N_3103,N_3023);
and U4220 (N_4220,N_3143,N_3090);
or U4221 (N_4221,N_3290,N_3703);
or U4222 (N_4222,N_3563,N_3348);
nand U4223 (N_4223,N_3045,N_3782);
and U4224 (N_4224,N_3834,N_3851);
or U4225 (N_4225,N_3463,N_3233);
xor U4226 (N_4226,N_3396,N_3401);
and U4227 (N_4227,N_3605,N_3508);
or U4228 (N_4228,N_3527,N_3470);
or U4229 (N_4229,N_3216,N_3195);
nand U4230 (N_4230,N_3627,N_3727);
and U4231 (N_4231,N_3063,N_3455);
and U4232 (N_4232,N_3030,N_3974);
and U4233 (N_4233,N_3286,N_3546);
nand U4234 (N_4234,N_3776,N_3676);
and U4235 (N_4235,N_3184,N_3496);
and U4236 (N_4236,N_3014,N_3247);
nor U4237 (N_4237,N_3940,N_3389);
nand U4238 (N_4238,N_3189,N_3076);
nand U4239 (N_4239,N_3562,N_3026);
xor U4240 (N_4240,N_3711,N_3169);
and U4241 (N_4241,N_3995,N_3153);
or U4242 (N_4242,N_3291,N_3517);
nand U4243 (N_4243,N_3339,N_3075);
nand U4244 (N_4244,N_3987,N_3442);
or U4245 (N_4245,N_3836,N_3057);
nor U4246 (N_4246,N_3217,N_3467);
or U4247 (N_4247,N_3817,N_3066);
nor U4248 (N_4248,N_3533,N_3818);
nor U4249 (N_4249,N_3659,N_3208);
nor U4250 (N_4250,N_3897,N_3213);
and U4251 (N_4251,N_3484,N_3619);
nor U4252 (N_4252,N_3575,N_3668);
nor U4253 (N_4253,N_3985,N_3941);
or U4254 (N_4254,N_3585,N_3938);
nor U4255 (N_4255,N_3774,N_3521);
nor U4256 (N_4256,N_3448,N_3084);
nor U4257 (N_4257,N_3055,N_3197);
and U4258 (N_4258,N_3444,N_3613);
or U4259 (N_4259,N_3578,N_3480);
xor U4260 (N_4260,N_3873,N_3108);
nor U4261 (N_4261,N_3816,N_3341);
nor U4262 (N_4262,N_3629,N_3445);
nor U4263 (N_4263,N_3518,N_3568);
and U4264 (N_4264,N_3607,N_3069);
xor U4265 (N_4265,N_3338,N_3079);
nand U4266 (N_4266,N_3074,N_3352);
or U4267 (N_4267,N_3544,N_3557);
or U4268 (N_4268,N_3146,N_3371);
nor U4269 (N_4269,N_3005,N_3963);
or U4270 (N_4270,N_3041,N_3495);
nor U4271 (N_4271,N_3869,N_3986);
nand U4272 (N_4272,N_3276,N_3240);
and U4273 (N_4273,N_3942,N_3783);
xor U4274 (N_4274,N_3381,N_3284);
and U4275 (N_4275,N_3294,N_3536);
nand U4276 (N_4276,N_3326,N_3375);
nor U4277 (N_4277,N_3656,N_3166);
and U4278 (N_4278,N_3937,N_3787);
and U4279 (N_4279,N_3377,N_3651);
nor U4280 (N_4280,N_3909,N_3922);
and U4281 (N_4281,N_3712,N_3833);
or U4282 (N_4282,N_3979,N_3337);
and U4283 (N_4283,N_3161,N_3843);
nor U4284 (N_4284,N_3300,N_3539);
nand U4285 (N_4285,N_3887,N_3417);
and U4286 (N_4286,N_3669,N_3307);
nor U4287 (N_4287,N_3980,N_3637);
nand U4288 (N_4288,N_3958,N_3248);
or U4289 (N_4289,N_3596,N_3696);
xnor U4290 (N_4290,N_3436,N_3193);
nor U4291 (N_4291,N_3200,N_3970);
or U4292 (N_4292,N_3638,N_3441);
xnor U4293 (N_4293,N_3363,N_3821);
and U4294 (N_4294,N_3840,N_3653);
nand U4295 (N_4295,N_3280,N_3173);
and U4296 (N_4296,N_3763,N_3871);
or U4297 (N_4297,N_3716,N_3275);
nor U4298 (N_4298,N_3946,N_3305);
nor U4299 (N_4299,N_3632,N_3308);
xor U4300 (N_4300,N_3849,N_3025);
nand U4301 (N_4301,N_3803,N_3304);
and U4302 (N_4302,N_3641,N_3977);
and U4303 (N_4303,N_3412,N_3925);
nor U4304 (N_4304,N_3875,N_3505);
and U4305 (N_4305,N_3477,N_3336);
nor U4306 (N_4306,N_3106,N_3535);
or U4307 (N_4307,N_3115,N_3786);
nand U4308 (N_4308,N_3319,N_3854);
and U4309 (N_4309,N_3961,N_3893);
xor U4310 (N_4310,N_3292,N_3274);
and U4311 (N_4311,N_3209,N_3996);
or U4312 (N_4312,N_3616,N_3241);
nor U4313 (N_4313,N_3449,N_3111);
nor U4314 (N_4314,N_3320,N_3485);
nand U4315 (N_4315,N_3929,N_3663);
nor U4316 (N_4316,N_3931,N_3132);
or U4317 (N_4317,N_3080,N_3658);
and U4318 (N_4318,N_3482,N_3430);
and U4319 (N_4319,N_3258,N_3540);
nor U4320 (N_4320,N_3354,N_3511);
nor U4321 (N_4321,N_3808,N_3050);
xor U4322 (N_4322,N_3263,N_3052);
xnor U4323 (N_4323,N_3008,N_3311);
xor U4324 (N_4324,N_3151,N_3694);
or U4325 (N_4325,N_3361,N_3024);
nand U4326 (N_4326,N_3387,N_3419);
nand U4327 (N_4327,N_3201,N_3670);
nand U4328 (N_4328,N_3164,N_3479);
nor U4329 (N_4329,N_3415,N_3982);
nor U4330 (N_4330,N_3914,N_3277);
nand U4331 (N_4331,N_3264,N_3229);
and U4332 (N_4332,N_3664,N_3335);
or U4333 (N_4333,N_3935,N_3876);
xor U4334 (N_4334,N_3798,N_3093);
and U4335 (N_4335,N_3813,N_3531);
and U4336 (N_4336,N_3422,N_3082);
and U4337 (N_4337,N_3804,N_3593);
and U4338 (N_4338,N_3309,N_3597);
nor U4339 (N_4339,N_3502,N_3566);
or U4340 (N_4340,N_3728,N_3497);
or U4341 (N_4341,N_3780,N_3118);
or U4342 (N_4342,N_3594,N_3185);
or U4343 (N_4343,N_3736,N_3135);
and U4344 (N_4344,N_3393,N_3493);
and U4345 (N_4345,N_3702,N_3503);
nand U4346 (N_4346,N_3955,N_3690);
xor U4347 (N_4347,N_3756,N_3577);
and U4348 (N_4348,N_3541,N_3269);
and U4349 (N_4349,N_3766,N_3951);
or U4350 (N_4350,N_3628,N_3239);
nor U4351 (N_4351,N_3171,N_3242);
nor U4352 (N_4352,N_3004,N_3602);
and U4353 (N_4353,N_3684,N_3771);
and U4354 (N_4354,N_3299,N_3498);
or U4355 (N_4355,N_3679,N_3571);
and U4356 (N_4356,N_3945,N_3983);
nand U4357 (N_4357,N_3345,N_3603);
or U4358 (N_4358,N_3867,N_3681);
or U4359 (N_4359,N_3494,N_3298);
or U4360 (N_4360,N_3420,N_3579);
xor U4361 (N_4361,N_3225,N_3959);
xor U4362 (N_4362,N_3172,N_3048);
and U4363 (N_4363,N_3194,N_3403);
nand U4364 (N_4364,N_3620,N_3705);
xnor U4365 (N_4365,N_3295,N_3249);
nor U4366 (N_4366,N_3509,N_3092);
nand U4367 (N_4367,N_3126,N_3906);
and U4368 (N_4368,N_3956,N_3491);
xor U4369 (N_4369,N_3991,N_3501);
or U4370 (N_4370,N_3123,N_3746);
or U4371 (N_4371,N_3158,N_3259);
or U4372 (N_4372,N_3243,N_3096);
or U4373 (N_4373,N_3283,N_3894);
nor U4374 (N_4374,N_3749,N_3492);
nor U4375 (N_4375,N_3998,N_3418);
and U4376 (N_4376,N_3560,N_3198);
nand U4377 (N_4377,N_3478,N_3230);
and U4378 (N_4378,N_3088,N_3565);
nand U4379 (N_4379,N_3891,N_3451);
nand U4380 (N_4380,N_3219,N_3234);
or U4381 (N_4381,N_3297,N_3677);
or U4382 (N_4382,N_3481,N_3794);
nand U4383 (N_4383,N_3316,N_3743);
and U4384 (N_4384,N_3863,N_3735);
nand U4385 (N_4385,N_3965,N_3317);
nor U4386 (N_4386,N_3757,N_3765);
or U4387 (N_4387,N_3456,N_3314);
or U4388 (N_4388,N_3969,N_3657);
xnor U4389 (N_4389,N_3815,N_3673);
nor U4390 (N_4390,N_3328,N_3323);
or U4391 (N_4391,N_3179,N_3119);
nand U4392 (N_4392,N_3831,N_3513);
nand U4393 (N_4393,N_3500,N_3034);
xor U4394 (N_4394,N_3529,N_3631);
nand U4395 (N_4395,N_3407,N_3353);
nand U4396 (N_4396,N_3124,N_3989);
nand U4397 (N_4397,N_3254,N_3186);
nor U4398 (N_4398,N_3285,N_3761);
xnor U4399 (N_4399,N_3882,N_3235);
and U4400 (N_4400,N_3848,N_3839);
or U4401 (N_4401,N_3853,N_3841);
or U4402 (N_4402,N_3347,N_3586);
nand U4403 (N_4403,N_3755,N_3270);
and U4404 (N_4404,N_3370,N_3476);
and U4405 (N_4405,N_3741,N_3112);
or U4406 (N_4406,N_3228,N_3827);
xnor U4407 (N_4407,N_3592,N_3650);
nor U4408 (N_4408,N_3040,N_3623);
xor U4409 (N_4409,N_3105,N_3751);
and U4410 (N_4410,N_3784,N_3047);
nor U4411 (N_4411,N_3777,N_3122);
or U4412 (N_4412,N_3554,N_3138);
and U4413 (N_4413,N_3832,N_3999);
nor U4414 (N_4414,N_3691,N_3883);
nand U4415 (N_4415,N_3934,N_3905);
nor U4416 (N_4416,N_3964,N_3801);
and U4417 (N_4417,N_3331,N_3157);
and U4418 (N_4418,N_3689,N_3866);
nand U4419 (N_4419,N_3988,N_3367);
nor U4420 (N_4420,N_3046,N_3013);
nor U4421 (N_4421,N_3971,N_3693);
nor U4422 (N_4422,N_3273,N_3717);
nand U4423 (N_4423,N_3145,N_3522);
or U4424 (N_4424,N_3845,N_3952);
or U4425 (N_4425,N_3266,N_3429);
and U4426 (N_4426,N_3738,N_3960);
nand U4427 (N_4427,N_3237,N_3432);
and U4428 (N_4428,N_3667,N_3409);
and U4429 (N_4429,N_3056,N_3506);
nand U4430 (N_4430,N_3862,N_3133);
nand U4431 (N_4431,N_3939,N_3826);
nand U4432 (N_4432,N_3550,N_3796);
and U4433 (N_4433,N_3433,N_3204);
xor U4434 (N_4434,N_3246,N_3110);
nand U4435 (N_4435,N_3870,N_3538);
xnor U4436 (N_4436,N_3850,N_3459);
nand U4437 (N_4437,N_3606,N_3820);
xor U4438 (N_4438,N_3708,N_3116);
or U4439 (N_4439,N_3584,N_3342);
nand U4440 (N_4440,N_3558,N_3576);
and U4441 (N_4441,N_3165,N_3085);
and U4442 (N_4442,N_3282,N_3210);
xnor U4443 (N_4443,N_3545,N_3601);
nor U4444 (N_4444,N_3552,N_3107);
xnor U4445 (N_4445,N_3077,N_3006);
nor U4446 (N_4446,N_3001,N_3612);
and U4447 (N_4447,N_3062,N_3404);
and U4448 (N_4448,N_3515,N_3797);
and U4449 (N_4449,N_3462,N_3426);
and U4450 (N_4450,N_3391,N_3070);
nand U4451 (N_4451,N_3947,N_3150);
nand U4452 (N_4452,N_3600,N_3553);
and U4453 (N_4453,N_3900,N_3183);
or U4454 (N_4454,N_3881,N_3306);
xnor U4455 (N_4455,N_3927,N_3769);
and U4456 (N_4456,N_3067,N_3049);
nor U4457 (N_4457,N_3100,N_3302);
nand U4458 (N_4458,N_3896,N_3884);
nand U4459 (N_4459,N_3748,N_3532);
and U4460 (N_4460,N_3366,N_3626);
and U4461 (N_4461,N_3907,N_3678);
nor U4462 (N_4462,N_3383,N_3474);
nand U4463 (N_4463,N_3740,N_3795);
nand U4464 (N_4464,N_3860,N_3351);
and U4465 (N_4465,N_3671,N_3472);
or U4466 (N_4466,N_3281,N_3551);
or U4467 (N_4467,N_3113,N_3842);
nor U4468 (N_4468,N_3017,N_3414);
and U4469 (N_4469,N_3360,N_3256);
nand U4470 (N_4470,N_3622,N_3811);
nor U4471 (N_4471,N_3489,N_3176);
nor U4472 (N_4472,N_3865,N_3731);
nand U4473 (N_4473,N_3904,N_3443);
and U4474 (N_4474,N_3589,N_3978);
or U4475 (N_4475,N_3131,N_3021);
xnor U4476 (N_4476,N_3824,N_3844);
xnor U4477 (N_4477,N_3382,N_3507);
or U4478 (N_4478,N_3715,N_3737);
or U4479 (N_4479,N_3016,N_3590);
nand U4480 (N_4480,N_3226,N_3548);
or U4481 (N_4481,N_3372,N_3061);
nor U4482 (N_4482,N_3181,N_3846);
and U4483 (N_4483,N_3018,N_3823);
xor U4484 (N_4484,N_3271,N_3411);
xnor U4485 (N_4485,N_3829,N_3972);
nand U4486 (N_4486,N_3142,N_3128);
or U4487 (N_4487,N_3514,N_3916);
or U4488 (N_4488,N_3159,N_3220);
nand U4489 (N_4489,N_3752,N_3556);
or U4490 (N_4490,N_3325,N_3188);
nand U4491 (N_4491,N_3890,N_3649);
or U4492 (N_4492,N_3038,N_3388);
and U4493 (N_4493,N_3129,N_3581);
nand U4494 (N_4494,N_3003,N_3064);
and U4495 (N_4495,N_3120,N_3990);
nand U4496 (N_4496,N_3461,N_3160);
nand U4497 (N_4497,N_3610,N_3261);
nor U4498 (N_4498,N_3549,N_3152);
xnor U4499 (N_4499,N_3262,N_3236);
nor U4500 (N_4500,N_3302,N_3377);
or U4501 (N_4501,N_3875,N_3428);
and U4502 (N_4502,N_3238,N_3449);
or U4503 (N_4503,N_3437,N_3703);
and U4504 (N_4504,N_3741,N_3968);
or U4505 (N_4505,N_3226,N_3199);
nand U4506 (N_4506,N_3960,N_3035);
and U4507 (N_4507,N_3290,N_3016);
or U4508 (N_4508,N_3781,N_3542);
nand U4509 (N_4509,N_3171,N_3857);
and U4510 (N_4510,N_3761,N_3875);
nor U4511 (N_4511,N_3011,N_3777);
nand U4512 (N_4512,N_3348,N_3822);
and U4513 (N_4513,N_3210,N_3442);
nand U4514 (N_4514,N_3936,N_3754);
xor U4515 (N_4515,N_3472,N_3428);
nor U4516 (N_4516,N_3780,N_3655);
and U4517 (N_4517,N_3548,N_3054);
and U4518 (N_4518,N_3561,N_3344);
nor U4519 (N_4519,N_3319,N_3024);
nand U4520 (N_4520,N_3496,N_3852);
nand U4521 (N_4521,N_3064,N_3347);
or U4522 (N_4522,N_3042,N_3850);
nand U4523 (N_4523,N_3800,N_3265);
and U4524 (N_4524,N_3963,N_3769);
xor U4525 (N_4525,N_3445,N_3734);
nor U4526 (N_4526,N_3247,N_3975);
or U4527 (N_4527,N_3309,N_3515);
xnor U4528 (N_4528,N_3399,N_3702);
nor U4529 (N_4529,N_3330,N_3270);
and U4530 (N_4530,N_3022,N_3958);
nor U4531 (N_4531,N_3948,N_3661);
nand U4532 (N_4532,N_3633,N_3022);
and U4533 (N_4533,N_3861,N_3635);
nor U4534 (N_4534,N_3839,N_3348);
nor U4535 (N_4535,N_3895,N_3501);
nor U4536 (N_4536,N_3245,N_3664);
and U4537 (N_4537,N_3385,N_3785);
nand U4538 (N_4538,N_3702,N_3083);
and U4539 (N_4539,N_3160,N_3821);
or U4540 (N_4540,N_3476,N_3295);
nor U4541 (N_4541,N_3291,N_3623);
nand U4542 (N_4542,N_3512,N_3279);
or U4543 (N_4543,N_3568,N_3127);
or U4544 (N_4544,N_3798,N_3848);
nor U4545 (N_4545,N_3924,N_3177);
nand U4546 (N_4546,N_3311,N_3699);
and U4547 (N_4547,N_3862,N_3547);
and U4548 (N_4548,N_3907,N_3922);
nand U4549 (N_4549,N_3572,N_3686);
nand U4550 (N_4550,N_3391,N_3811);
nand U4551 (N_4551,N_3198,N_3358);
xor U4552 (N_4552,N_3223,N_3915);
xnor U4553 (N_4553,N_3891,N_3253);
and U4554 (N_4554,N_3018,N_3805);
nand U4555 (N_4555,N_3342,N_3225);
nand U4556 (N_4556,N_3095,N_3527);
nor U4557 (N_4557,N_3512,N_3418);
nand U4558 (N_4558,N_3169,N_3577);
or U4559 (N_4559,N_3649,N_3960);
and U4560 (N_4560,N_3739,N_3701);
and U4561 (N_4561,N_3867,N_3701);
and U4562 (N_4562,N_3236,N_3229);
and U4563 (N_4563,N_3272,N_3067);
nand U4564 (N_4564,N_3181,N_3147);
xor U4565 (N_4565,N_3227,N_3521);
nor U4566 (N_4566,N_3460,N_3962);
and U4567 (N_4567,N_3192,N_3684);
or U4568 (N_4568,N_3335,N_3976);
nand U4569 (N_4569,N_3533,N_3027);
xor U4570 (N_4570,N_3442,N_3350);
or U4571 (N_4571,N_3314,N_3678);
nand U4572 (N_4572,N_3971,N_3491);
nor U4573 (N_4573,N_3344,N_3686);
or U4574 (N_4574,N_3955,N_3626);
nor U4575 (N_4575,N_3148,N_3609);
or U4576 (N_4576,N_3903,N_3217);
or U4577 (N_4577,N_3506,N_3101);
nor U4578 (N_4578,N_3697,N_3496);
or U4579 (N_4579,N_3512,N_3763);
nand U4580 (N_4580,N_3600,N_3405);
or U4581 (N_4581,N_3174,N_3992);
nand U4582 (N_4582,N_3455,N_3296);
or U4583 (N_4583,N_3338,N_3931);
or U4584 (N_4584,N_3288,N_3352);
nand U4585 (N_4585,N_3061,N_3787);
and U4586 (N_4586,N_3695,N_3339);
and U4587 (N_4587,N_3260,N_3063);
xnor U4588 (N_4588,N_3859,N_3127);
or U4589 (N_4589,N_3789,N_3932);
or U4590 (N_4590,N_3614,N_3715);
and U4591 (N_4591,N_3611,N_3516);
nand U4592 (N_4592,N_3741,N_3154);
and U4593 (N_4593,N_3117,N_3827);
xor U4594 (N_4594,N_3440,N_3810);
nor U4595 (N_4595,N_3442,N_3900);
nand U4596 (N_4596,N_3883,N_3742);
or U4597 (N_4597,N_3318,N_3922);
nor U4598 (N_4598,N_3037,N_3640);
nor U4599 (N_4599,N_3098,N_3188);
xnor U4600 (N_4600,N_3165,N_3338);
and U4601 (N_4601,N_3828,N_3033);
nand U4602 (N_4602,N_3228,N_3455);
xor U4603 (N_4603,N_3693,N_3176);
nor U4604 (N_4604,N_3662,N_3425);
nand U4605 (N_4605,N_3134,N_3578);
nor U4606 (N_4606,N_3749,N_3124);
nor U4607 (N_4607,N_3177,N_3933);
nor U4608 (N_4608,N_3792,N_3844);
nand U4609 (N_4609,N_3423,N_3226);
or U4610 (N_4610,N_3166,N_3995);
nor U4611 (N_4611,N_3144,N_3706);
and U4612 (N_4612,N_3830,N_3831);
nand U4613 (N_4613,N_3616,N_3371);
or U4614 (N_4614,N_3840,N_3118);
nor U4615 (N_4615,N_3304,N_3482);
xnor U4616 (N_4616,N_3247,N_3333);
or U4617 (N_4617,N_3073,N_3047);
nor U4618 (N_4618,N_3694,N_3479);
nor U4619 (N_4619,N_3511,N_3013);
nand U4620 (N_4620,N_3044,N_3576);
or U4621 (N_4621,N_3194,N_3848);
nand U4622 (N_4622,N_3306,N_3185);
xor U4623 (N_4623,N_3781,N_3750);
nor U4624 (N_4624,N_3169,N_3037);
nand U4625 (N_4625,N_3792,N_3049);
or U4626 (N_4626,N_3703,N_3676);
and U4627 (N_4627,N_3362,N_3648);
or U4628 (N_4628,N_3262,N_3394);
xor U4629 (N_4629,N_3700,N_3727);
nor U4630 (N_4630,N_3587,N_3143);
or U4631 (N_4631,N_3521,N_3909);
and U4632 (N_4632,N_3184,N_3068);
and U4633 (N_4633,N_3267,N_3608);
nor U4634 (N_4634,N_3758,N_3022);
and U4635 (N_4635,N_3557,N_3551);
nand U4636 (N_4636,N_3693,N_3797);
or U4637 (N_4637,N_3056,N_3945);
or U4638 (N_4638,N_3869,N_3969);
nand U4639 (N_4639,N_3446,N_3993);
and U4640 (N_4640,N_3768,N_3577);
or U4641 (N_4641,N_3245,N_3115);
or U4642 (N_4642,N_3951,N_3378);
nand U4643 (N_4643,N_3800,N_3649);
or U4644 (N_4644,N_3064,N_3426);
nor U4645 (N_4645,N_3847,N_3793);
nor U4646 (N_4646,N_3816,N_3575);
or U4647 (N_4647,N_3074,N_3636);
nand U4648 (N_4648,N_3498,N_3252);
xnor U4649 (N_4649,N_3289,N_3168);
or U4650 (N_4650,N_3022,N_3561);
nand U4651 (N_4651,N_3177,N_3191);
nand U4652 (N_4652,N_3866,N_3128);
nor U4653 (N_4653,N_3220,N_3877);
or U4654 (N_4654,N_3876,N_3863);
nor U4655 (N_4655,N_3823,N_3481);
and U4656 (N_4656,N_3849,N_3194);
nand U4657 (N_4657,N_3578,N_3005);
or U4658 (N_4658,N_3415,N_3712);
or U4659 (N_4659,N_3495,N_3403);
nand U4660 (N_4660,N_3153,N_3879);
or U4661 (N_4661,N_3528,N_3719);
and U4662 (N_4662,N_3988,N_3817);
nand U4663 (N_4663,N_3551,N_3392);
xor U4664 (N_4664,N_3977,N_3240);
and U4665 (N_4665,N_3711,N_3403);
nor U4666 (N_4666,N_3576,N_3345);
xnor U4667 (N_4667,N_3440,N_3617);
or U4668 (N_4668,N_3583,N_3123);
nor U4669 (N_4669,N_3070,N_3639);
or U4670 (N_4670,N_3693,N_3859);
nand U4671 (N_4671,N_3703,N_3365);
nor U4672 (N_4672,N_3909,N_3953);
nor U4673 (N_4673,N_3861,N_3951);
or U4674 (N_4674,N_3203,N_3472);
or U4675 (N_4675,N_3769,N_3117);
or U4676 (N_4676,N_3880,N_3836);
or U4677 (N_4677,N_3750,N_3163);
and U4678 (N_4678,N_3144,N_3712);
nand U4679 (N_4679,N_3571,N_3731);
and U4680 (N_4680,N_3830,N_3300);
nand U4681 (N_4681,N_3959,N_3195);
and U4682 (N_4682,N_3455,N_3522);
nor U4683 (N_4683,N_3731,N_3604);
or U4684 (N_4684,N_3450,N_3233);
and U4685 (N_4685,N_3987,N_3193);
and U4686 (N_4686,N_3732,N_3784);
nor U4687 (N_4687,N_3982,N_3602);
nand U4688 (N_4688,N_3385,N_3598);
or U4689 (N_4689,N_3804,N_3573);
xor U4690 (N_4690,N_3597,N_3300);
nand U4691 (N_4691,N_3734,N_3303);
or U4692 (N_4692,N_3103,N_3733);
nand U4693 (N_4693,N_3834,N_3552);
and U4694 (N_4694,N_3978,N_3904);
or U4695 (N_4695,N_3334,N_3888);
xor U4696 (N_4696,N_3165,N_3294);
nor U4697 (N_4697,N_3447,N_3176);
or U4698 (N_4698,N_3332,N_3998);
nand U4699 (N_4699,N_3858,N_3170);
nor U4700 (N_4700,N_3573,N_3147);
and U4701 (N_4701,N_3603,N_3469);
nand U4702 (N_4702,N_3930,N_3171);
nand U4703 (N_4703,N_3114,N_3975);
nand U4704 (N_4704,N_3747,N_3864);
and U4705 (N_4705,N_3117,N_3998);
and U4706 (N_4706,N_3296,N_3311);
nor U4707 (N_4707,N_3533,N_3392);
or U4708 (N_4708,N_3017,N_3357);
or U4709 (N_4709,N_3134,N_3673);
nor U4710 (N_4710,N_3487,N_3620);
and U4711 (N_4711,N_3913,N_3733);
and U4712 (N_4712,N_3522,N_3621);
and U4713 (N_4713,N_3774,N_3563);
or U4714 (N_4714,N_3631,N_3866);
and U4715 (N_4715,N_3772,N_3273);
nand U4716 (N_4716,N_3763,N_3032);
or U4717 (N_4717,N_3766,N_3601);
nor U4718 (N_4718,N_3134,N_3704);
or U4719 (N_4719,N_3835,N_3719);
xor U4720 (N_4720,N_3230,N_3411);
nand U4721 (N_4721,N_3568,N_3768);
xor U4722 (N_4722,N_3532,N_3950);
and U4723 (N_4723,N_3245,N_3700);
or U4724 (N_4724,N_3636,N_3053);
and U4725 (N_4725,N_3256,N_3698);
xnor U4726 (N_4726,N_3944,N_3617);
and U4727 (N_4727,N_3218,N_3752);
or U4728 (N_4728,N_3853,N_3150);
or U4729 (N_4729,N_3747,N_3942);
nor U4730 (N_4730,N_3742,N_3888);
nand U4731 (N_4731,N_3507,N_3569);
nor U4732 (N_4732,N_3374,N_3339);
nand U4733 (N_4733,N_3517,N_3094);
or U4734 (N_4734,N_3607,N_3310);
or U4735 (N_4735,N_3068,N_3056);
nand U4736 (N_4736,N_3213,N_3461);
and U4737 (N_4737,N_3085,N_3588);
nor U4738 (N_4738,N_3421,N_3402);
and U4739 (N_4739,N_3697,N_3261);
nor U4740 (N_4740,N_3611,N_3923);
nand U4741 (N_4741,N_3677,N_3398);
nor U4742 (N_4742,N_3023,N_3262);
and U4743 (N_4743,N_3831,N_3089);
nor U4744 (N_4744,N_3435,N_3246);
or U4745 (N_4745,N_3405,N_3412);
nand U4746 (N_4746,N_3095,N_3009);
nand U4747 (N_4747,N_3492,N_3771);
xnor U4748 (N_4748,N_3136,N_3040);
or U4749 (N_4749,N_3161,N_3673);
and U4750 (N_4750,N_3257,N_3794);
and U4751 (N_4751,N_3617,N_3095);
nor U4752 (N_4752,N_3127,N_3805);
and U4753 (N_4753,N_3036,N_3763);
or U4754 (N_4754,N_3934,N_3434);
or U4755 (N_4755,N_3748,N_3217);
nand U4756 (N_4756,N_3858,N_3787);
nand U4757 (N_4757,N_3274,N_3394);
nor U4758 (N_4758,N_3394,N_3487);
or U4759 (N_4759,N_3593,N_3519);
nand U4760 (N_4760,N_3952,N_3060);
nand U4761 (N_4761,N_3206,N_3271);
or U4762 (N_4762,N_3914,N_3673);
or U4763 (N_4763,N_3250,N_3581);
or U4764 (N_4764,N_3055,N_3832);
nor U4765 (N_4765,N_3123,N_3375);
nor U4766 (N_4766,N_3826,N_3790);
and U4767 (N_4767,N_3694,N_3370);
and U4768 (N_4768,N_3339,N_3640);
nand U4769 (N_4769,N_3464,N_3709);
or U4770 (N_4770,N_3951,N_3259);
and U4771 (N_4771,N_3400,N_3312);
or U4772 (N_4772,N_3405,N_3212);
nor U4773 (N_4773,N_3030,N_3477);
and U4774 (N_4774,N_3438,N_3520);
nand U4775 (N_4775,N_3662,N_3042);
nand U4776 (N_4776,N_3655,N_3498);
or U4777 (N_4777,N_3307,N_3319);
nor U4778 (N_4778,N_3480,N_3420);
nand U4779 (N_4779,N_3600,N_3529);
nand U4780 (N_4780,N_3084,N_3414);
and U4781 (N_4781,N_3325,N_3990);
nand U4782 (N_4782,N_3341,N_3588);
or U4783 (N_4783,N_3081,N_3117);
and U4784 (N_4784,N_3243,N_3831);
and U4785 (N_4785,N_3058,N_3522);
nor U4786 (N_4786,N_3592,N_3499);
nand U4787 (N_4787,N_3107,N_3372);
or U4788 (N_4788,N_3685,N_3073);
xnor U4789 (N_4789,N_3668,N_3059);
xor U4790 (N_4790,N_3585,N_3989);
nand U4791 (N_4791,N_3075,N_3048);
or U4792 (N_4792,N_3646,N_3382);
nand U4793 (N_4793,N_3322,N_3618);
nor U4794 (N_4794,N_3997,N_3007);
nor U4795 (N_4795,N_3865,N_3575);
nor U4796 (N_4796,N_3615,N_3262);
nor U4797 (N_4797,N_3890,N_3600);
nor U4798 (N_4798,N_3310,N_3100);
or U4799 (N_4799,N_3673,N_3644);
nor U4800 (N_4800,N_3418,N_3617);
nand U4801 (N_4801,N_3849,N_3117);
nor U4802 (N_4802,N_3267,N_3939);
and U4803 (N_4803,N_3379,N_3463);
and U4804 (N_4804,N_3898,N_3476);
nand U4805 (N_4805,N_3193,N_3040);
nand U4806 (N_4806,N_3763,N_3910);
and U4807 (N_4807,N_3820,N_3612);
nand U4808 (N_4808,N_3716,N_3616);
nand U4809 (N_4809,N_3849,N_3540);
nand U4810 (N_4810,N_3700,N_3026);
xnor U4811 (N_4811,N_3682,N_3039);
nor U4812 (N_4812,N_3261,N_3445);
or U4813 (N_4813,N_3257,N_3687);
or U4814 (N_4814,N_3927,N_3860);
xor U4815 (N_4815,N_3500,N_3715);
and U4816 (N_4816,N_3563,N_3726);
or U4817 (N_4817,N_3446,N_3318);
nor U4818 (N_4818,N_3843,N_3909);
or U4819 (N_4819,N_3858,N_3611);
xnor U4820 (N_4820,N_3319,N_3333);
and U4821 (N_4821,N_3684,N_3060);
nor U4822 (N_4822,N_3048,N_3818);
nor U4823 (N_4823,N_3121,N_3401);
or U4824 (N_4824,N_3542,N_3818);
nor U4825 (N_4825,N_3347,N_3274);
xor U4826 (N_4826,N_3264,N_3789);
and U4827 (N_4827,N_3842,N_3374);
and U4828 (N_4828,N_3253,N_3226);
and U4829 (N_4829,N_3822,N_3137);
xor U4830 (N_4830,N_3967,N_3020);
or U4831 (N_4831,N_3860,N_3619);
or U4832 (N_4832,N_3085,N_3479);
nand U4833 (N_4833,N_3287,N_3893);
and U4834 (N_4834,N_3820,N_3714);
nor U4835 (N_4835,N_3079,N_3470);
or U4836 (N_4836,N_3791,N_3821);
and U4837 (N_4837,N_3571,N_3072);
nor U4838 (N_4838,N_3111,N_3656);
xnor U4839 (N_4839,N_3642,N_3990);
nand U4840 (N_4840,N_3375,N_3817);
nand U4841 (N_4841,N_3337,N_3854);
and U4842 (N_4842,N_3614,N_3231);
and U4843 (N_4843,N_3080,N_3778);
xnor U4844 (N_4844,N_3951,N_3552);
nand U4845 (N_4845,N_3844,N_3407);
or U4846 (N_4846,N_3629,N_3708);
and U4847 (N_4847,N_3353,N_3280);
nand U4848 (N_4848,N_3905,N_3779);
or U4849 (N_4849,N_3766,N_3886);
nor U4850 (N_4850,N_3809,N_3911);
nor U4851 (N_4851,N_3328,N_3877);
nor U4852 (N_4852,N_3351,N_3788);
or U4853 (N_4853,N_3945,N_3648);
or U4854 (N_4854,N_3467,N_3900);
or U4855 (N_4855,N_3010,N_3941);
nand U4856 (N_4856,N_3637,N_3391);
or U4857 (N_4857,N_3817,N_3221);
xnor U4858 (N_4858,N_3847,N_3835);
nand U4859 (N_4859,N_3043,N_3256);
xor U4860 (N_4860,N_3333,N_3514);
nor U4861 (N_4861,N_3141,N_3889);
or U4862 (N_4862,N_3513,N_3560);
and U4863 (N_4863,N_3572,N_3236);
nand U4864 (N_4864,N_3786,N_3881);
nor U4865 (N_4865,N_3752,N_3489);
or U4866 (N_4866,N_3146,N_3224);
or U4867 (N_4867,N_3937,N_3159);
xor U4868 (N_4868,N_3423,N_3494);
nor U4869 (N_4869,N_3910,N_3552);
xor U4870 (N_4870,N_3897,N_3076);
or U4871 (N_4871,N_3773,N_3954);
nor U4872 (N_4872,N_3264,N_3846);
or U4873 (N_4873,N_3118,N_3045);
or U4874 (N_4874,N_3114,N_3270);
nor U4875 (N_4875,N_3985,N_3768);
nand U4876 (N_4876,N_3307,N_3918);
xnor U4877 (N_4877,N_3372,N_3324);
and U4878 (N_4878,N_3299,N_3501);
nand U4879 (N_4879,N_3531,N_3789);
xor U4880 (N_4880,N_3317,N_3477);
nand U4881 (N_4881,N_3704,N_3364);
nor U4882 (N_4882,N_3896,N_3628);
or U4883 (N_4883,N_3567,N_3634);
and U4884 (N_4884,N_3805,N_3515);
and U4885 (N_4885,N_3521,N_3982);
nand U4886 (N_4886,N_3443,N_3771);
nand U4887 (N_4887,N_3712,N_3452);
xnor U4888 (N_4888,N_3510,N_3089);
nand U4889 (N_4889,N_3097,N_3647);
or U4890 (N_4890,N_3614,N_3973);
nand U4891 (N_4891,N_3026,N_3860);
nand U4892 (N_4892,N_3615,N_3785);
and U4893 (N_4893,N_3992,N_3036);
nand U4894 (N_4894,N_3075,N_3466);
nor U4895 (N_4895,N_3861,N_3404);
nor U4896 (N_4896,N_3204,N_3734);
nand U4897 (N_4897,N_3371,N_3015);
nor U4898 (N_4898,N_3818,N_3858);
and U4899 (N_4899,N_3674,N_3140);
or U4900 (N_4900,N_3462,N_3903);
and U4901 (N_4901,N_3357,N_3821);
or U4902 (N_4902,N_3902,N_3443);
nand U4903 (N_4903,N_3322,N_3805);
and U4904 (N_4904,N_3148,N_3770);
nand U4905 (N_4905,N_3404,N_3800);
nand U4906 (N_4906,N_3626,N_3964);
nor U4907 (N_4907,N_3996,N_3504);
xnor U4908 (N_4908,N_3926,N_3098);
nor U4909 (N_4909,N_3585,N_3705);
nand U4910 (N_4910,N_3409,N_3092);
and U4911 (N_4911,N_3737,N_3192);
and U4912 (N_4912,N_3856,N_3042);
and U4913 (N_4913,N_3894,N_3693);
xnor U4914 (N_4914,N_3764,N_3648);
nor U4915 (N_4915,N_3450,N_3749);
xor U4916 (N_4916,N_3791,N_3044);
or U4917 (N_4917,N_3470,N_3092);
nor U4918 (N_4918,N_3779,N_3911);
xor U4919 (N_4919,N_3881,N_3897);
and U4920 (N_4920,N_3118,N_3754);
or U4921 (N_4921,N_3333,N_3827);
nand U4922 (N_4922,N_3532,N_3503);
or U4923 (N_4923,N_3180,N_3559);
or U4924 (N_4924,N_3632,N_3094);
and U4925 (N_4925,N_3878,N_3619);
nor U4926 (N_4926,N_3518,N_3821);
or U4927 (N_4927,N_3712,N_3610);
nor U4928 (N_4928,N_3191,N_3224);
nor U4929 (N_4929,N_3850,N_3126);
nor U4930 (N_4930,N_3912,N_3778);
and U4931 (N_4931,N_3723,N_3102);
nand U4932 (N_4932,N_3025,N_3264);
nand U4933 (N_4933,N_3688,N_3301);
or U4934 (N_4934,N_3628,N_3593);
nor U4935 (N_4935,N_3501,N_3519);
and U4936 (N_4936,N_3816,N_3510);
nor U4937 (N_4937,N_3759,N_3942);
nor U4938 (N_4938,N_3350,N_3701);
and U4939 (N_4939,N_3203,N_3503);
nand U4940 (N_4940,N_3638,N_3692);
nand U4941 (N_4941,N_3596,N_3466);
or U4942 (N_4942,N_3788,N_3041);
xor U4943 (N_4943,N_3001,N_3642);
nor U4944 (N_4944,N_3691,N_3473);
nor U4945 (N_4945,N_3822,N_3119);
nand U4946 (N_4946,N_3132,N_3151);
nor U4947 (N_4947,N_3484,N_3927);
nor U4948 (N_4948,N_3989,N_3138);
xnor U4949 (N_4949,N_3784,N_3066);
or U4950 (N_4950,N_3342,N_3170);
and U4951 (N_4951,N_3279,N_3255);
nor U4952 (N_4952,N_3179,N_3794);
nor U4953 (N_4953,N_3557,N_3849);
nor U4954 (N_4954,N_3986,N_3990);
nand U4955 (N_4955,N_3059,N_3412);
and U4956 (N_4956,N_3498,N_3196);
or U4957 (N_4957,N_3694,N_3824);
nor U4958 (N_4958,N_3815,N_3167);
and U4959 (N_4959,N_3965,N_3192);
nand U4960 (N_4960,N_3642,N_3251);
nor U4961 (N_4961,N_3953,N_3293);
or U4962 (N_4962,N_3101,N_3776);
nor U4963 (N_4963,N_3197,N_3845);
nor U4964 (N_4964,N_3946,N_3414);
nand U4965 (N_4965,N_3120,N_3620);
and U4966 (N_4966,N_3683,N_3639);
or U4967 (N_4967,N_3043,N_3614);
nand U4968 (N_4968,N_3825,N_3106);
nand U4969 (N_4969,N_3334,N_3233);
nand U4970 (N_4970,N_3644,N_3580);
nor U4971 (N_4971,N_3656,N_3620);
or U4972 (N_4972,N_3782,N_3007);
and U4973 (N_4973,N_3243,N_3826);
nand U4974 (N_4974,N_3369,N_3632);
and U4975 (N_4975,N_3727,N_3657);
and U4976 (N_4976,N_3361,N_3624);
xor U4977 (N_4977,N_3205,N_3822);
xnor U4978 (N_4978,N_3691,N_3201);
or U4979 (N_4979,N_3115,N_3881);
or U4980 (N_4980,N_3122,N_3559);
nand U4981 (N_4981,N_3745,N_3341);
and U4982 (N_4982,N_3210,N_3343);
or U4983 (N_4983,N_3506,N_3612);
nand U4984 (N_4984,N_3935,N_3160);
nand U4985 (N_4985,N_3989,N_3007);
and U4986 (N_4986,N_3633,N_3549);
nand U4987 (N_4987,N_3817,N_3426);
nand U4988 (N_4988,N_3931,N_3334);
nand U4989 (N_4989,N_3718,N_3778);
and U4990 (N_4990,N_3138,N_3254);
or U4991 (N_4991,N_3773,N_3566);
or U4992 (N_4992,N_3823,N_3618);
nor U4993 (N_4993,N_3712,N_3204);
nor U4994 (N_4994,N_3711,N_3863);
nor U4995 (N_4995,N_3914,N_3526);
nand U4996 (N_4996,N_3648,N_3285);
nor U4997 (N_4997,N_3499,N_3218);
and U4998 (N_4998,N_3762,N_3247);
xor U4999 (N_4999,N_3334,N_3508);
nor U5000 (N_5000,N_4504,N_4799);
or U5001 (N_5001,N_4171,N_4222);
nor U5002 (N_5002,N_4165,N_4653);
nor U5003 (N_5003,N_4281,N_4709);
or U5004 (N_5004,N_4532,N_4478);
or U5005 (N_5005,N_4746,N_4017);
xnor U5006 (N_5006,N_4909,N_4649);
nor U5007 (N_5007,N_4263,N_4160);
nor U5008 (N_5008,N_4033,N_4391);
and U5009 (N_5009,N_4704,N_4250);
and U5010 (N_5010,N_4121,N_4659);
nand U5011 (N_5011,N_4351,N_4661);
nor U5012 (N_5012,N_4777,N_4278);
nand U5013 (N_5013,N_4436,N_4955);
xnor U5014 (N_5014,N_4758,N_4334);
and U5015 (N_5015,N_4193,N_4242);
or U5016 (N_5016,N_4969,N_4498);
xor U5017 (N_5017,N_4695,N_4755);
nor U5018 (N_5018,N_4198,N_4534);
nor U5019 (N_5019,N_4823,N_4308);
nor U5020 (N_5020,N_4817,N_4535);
nand U5021 (N_5021,N_4690,N_4793);
or U5022 (N_5022,N_4139,N_4177);
nor U5023 (N_5023,N_4830,N_4781);
or U5024 (N_5024,N_4975,N_4540);
or U5025 (N_5025,N_4025,N_4673);
or U5026 (N_5026,N_4031,N_4905);
xnor U5027 (N_5027,N_4063,N_4923);
nand U5028 (N_5028,N_4618,N_4306);
and U5029 (N_5029,N_4378,N_4485);
xor U5030 (N_5030,N_4617,N_4983);
or U5031 (N_5031,N_4068,N_4287);
nand U5032 (N_5032,N_4769,N_4097);
and U5033 (N_5033,N_4325,N_4006);
nor U5034 (N_5034,N_4414,N_4232);
or U5035 (N_5035,N_4884,N_4275);
or U5036 (N_5036,N_4609,N_4127);
nor U5037 (N_5037,N_4226,N_4423);
or U5038 (N_5038,N_4217,N_4066);
and U5039 (N_5039,N_4277,N_4965);
xor U5040 (N_5040,N_4625,N_4772);
nor U5041 (N_5041,N_4502,N_4529);
nor U5042 (N_5042,N_4548,N_4851);
nand U5043 (N_5043,N_4922,N_4749);
nor U5044 (N_5044,N_4071,N_4013);
nor U5045 (N_5045,N_4811,N_4435);
and U5046 (N_5046,N_4113,N_4696);
nor U5047 (N_5047,N_4432,N_4734);
or U5048 (N_5048,N_4952,N_4701);
or U5049 (N_5049,N_4740,N_4579);
nor U5050 (N_5050,N_4258,N_4296);
or U5051 (N_5051,N_4018,N_4512);
nand U5052 (N_5052,N_4642,N_4824);
xor U5053 (N_5053,N_4350,N_4474);
nor U5054 (N_5054,N_4570,N_4587);
nand U5055 (N_5055,N_4519,N_4981);
and U5056 (N_5056,N_4228,N_4191);
or U5057 (N_5057,N_4327,N_4770);
and U5058 (N_5058,N_4312,N_4329);
or U5059 (N_5059,N_4976,N_4132);
nor U5060 (N_5060,N_4784,N_4493);
and U5061 (N_5061,N_4883,N_4118);
or U5062 (N_5062,N_4463,N_4731);
nand U5063 (N_5063,N_4645,N_4856);
and U5064 (N_5064,N_4594,N_4789);
and U5065 (N_5065,N_4314,N_4814);
xor U5066 (N_5066,N_4773,N_4487);
and U5067 (N_5067,N_4410,N_4767);
nand U5068 (N_5068,N_4220,N_4804);
and U5069 (N_5069,N_4488,N_4933);
xor U5070 (N_5070,N_4073,N_4465);
nand U5071 (N_5071,N_4517,N_4868);
and U5072 (N_5072,N_4251,N_4227);
xnor U5073 (N_5073,N_4212,N_4954);
or U5074 (N_5074,N_4169,N_4866);
or U5075 (N_5075,N_4751,N_4706);
nand U5076 (N_5076,N_4224,N_4108);
nor U5077 (N_5077,N_4748,N_4691);
nand U5078 (N_5078,N_4128,N_4982);
or U5079 (N_5079,N_4028,N_4211);
nand U5080 (N_5080,N_4900,N_4276);
xnor U5081 (N_5081,N_4766,N_4871);
or U5082 (N_5082,N_4754,N_4371);
or U5083 (N_5083,N_4274,N_4084);
or U5084 (N_5084,N_4328,N_4189);
nor U5085 (N_5085,N_4421,N_4362);
or U5086 (N_5086,N_4455,N_4882);
and U5087 (N_5087,N_4925,N_4492);
nand U5088 (N_5088,N_4243,N_4176);
nor U5089 (N_5089,N_4660,N_4168);
and U5090 (N_5090,N_4787,N_4928);
nor U5091 (N_5091,N_4141,N_4626);
or U5092 (N_5092,N_4522,N_4458);
nor U5093 (N_5093,N_4462,N_4292);
and U5094 (N_5094,N_4857,N_4307);
and U5095 (N_5095,N_4873,N_4639);
or U5096 (N_5096,N_4855,N_4663);
and U5097 (N_5097,N_4914,N_4903);
and U5098 (N_5098,N_4852,N_4651);
or U5099 (N_5099,N_4468,N_4947);
and U5100 (N_5100,N_4916,N_4449);
xor U5101 (N_5101,N_4072,N_4581);
nand U5102 (N_5102,N_4816,N_4967);
nand U5103 (N_5103,N_4786,N_4346);
and U5104 (N_5104,N_4942,N_4050);
and U5105 (N_5105,N_4144,N_4398);
or U5106 (N_5106,N_4820,N_4082);
or U5107 (N_5107,N_4714,N_4496);
xor U5108 (N_5108,N_4537,N_4298);
nor U5109 (N_5109,N_4472,N_4842);
or U5110 (N_5110,N_4231,N_4099);
and U5111 (N_5111,N_4005,N_4111);
nor U5112 (N_5112,N_4284,N_4333);
or U5113 (N_5113,N_4322,N_4524);
nor U5114 (N_5114,N_4098,N_4646);
nand U5115 (N_5115,N_4388,N_4592);
nor U5116 (N_5116,N_4297,N_4878);
and U5117 (N_5117,N_4405,N_4505);
and U5118 (N_5118,N_4439,N_4602);
nand U5119 (N_5119,N_4178,N_4509);
nand U5120 (N_5120,N_4170,N_4630);
nand U5121 (N_5121,N_4611,N_4620);
nand U5122 (N_5122,N_4917,N_4107);
nor U5123 (N_5123,N_4513,N_4727);
nor U5124 (N_5124,N_4588,N_4778);
and U5125 (N_5125,N_4683,N_4939);
xnor U5126 (N_5126,N_4647,N_4945);
or U5127 (N_5127,N_4153,N_4416);
xnor U5128 (N_5128,N_4486,N_4270);
or U5129 (N_5129,N_4154,N_4273);
nand U5130 (N_5130,N_4407,N_4853);
or U5131 (N_5131,N_4996,N_4070);
nor U5132 (N_5132,N_4359,N_4818);
or U5133 (N_5133,N_4302,N_4632);
xor U5134 (N_5134,N_4460,N_4424);
or U5135 (N_5135,N_4149,N_4244);
or U5136 (N_5136,N_4563,N_4815);
nand U5137 (N_5137,N_4155,N_4138);
xor U5138 (N_5138,N_4961,N_4538);
and U5139 (N_5139,N_4790,N_4973);
or U5140 (N_5140,N_4791,N_4940);
or U5141 (N_5141,N_4461,N_4763);
nor U5142 (N_5142,N_4397,N_4725);
nor U5143 (N_5143,N_4356,N_4822);
nand U5144 (N_5144,N_4195,N_4571);
nor U5145 (N_5145,N_4627,N_4007);
nand U5146 (N_5146,N_4729,N_4849);
and U5147 (N_5147,N_4698,N_4023);
and U5148 (N_5148,N_4860,N_4010);
and U5149 (N_5149,N_4089,N_4349);
nand U5150 (N_5150,N_4466,N_4774);
or U5151 (N_5151,N_4958,N_4655);
and U5152 (N_5152,N_4283,N_4213);
nand U5153 (N_5153,N_4608,N_4511);
or U5154 (N_5154,N_4289,N_4825);
and U5155 (N_5155,N_4357,N_4876);
and U5156 (N_5156,N_4420,N_4959);
nor U5157 (N_5157,N_4009,N_4235);
or U5158 (N_5158,N_4848,N_4812);
nor U5159 (N_5159,N_4321,N_4190);
or U5160 (N_5160,N_4544,N_4204);
nor U5161 (N_5161,N_4590,N_4172);
nor U5162 (N_5162,N_4209,N_4951);
nand U5163 (N_5163,N_4831,N_4591);
nor U5164 (N_5164,N_4484,N_4305);
and U5165 (N_5165,N_4182,N_4313);
and U5166 (N_5166,N_4862,N_4207);
nand U5167 (N_5167,N_4992,N_4676);
nand U5168 (N_5168,N_4719,N_4366);
nor U5169 (N_5169,N_4384,N_4990);
and U5170 (N_5170,N_4722,N_4944);
nand U5171 (N_5171,N_4348,N_4562);
nor U5172 (N_5172,N_4389,N_4913);
nor U5173 (N_5173,N_4123,N_4881);
nor U5174 (N_5174,N_4158,N_4636);
xor U5175 (N_5175,N_4495,N_4723);
or U5176 (N_5176,N_4995,N_4672);
and U5177 (N_5177,N_4643,N_4827);
nand U5178 (N_5178,N_4867,N_4352);
nor U5179 (N_5179,N_4467,N_4670);
nand U5180 (N_5180,N_4026,N_4180);
nand U5181 (N_5181,N_4819,N_4614);
nor U5182 (N_5182,N_4078,N_4606);
xor U5183 (N_5183,N_4794,N_4797);
and U5184 (N_5184,N_4055,N_4151);
nand U5185 (N_5185,N_4607,N_4788);
xor U5186 (N_5186,N_4264,N_4253);
nand U5187 (N_5187,N_4092,N_4635);
or U5188 (N_5188,N_4454,N_4518);
and U5189 (N_5189,N_4104,N_4022);
and U5190 (N_5190,N_4971,N_4716);
nand U5191 (N_5191,N_4442,N_4057);
and U5192 (N_5192,N_4680,N_4911);
or U5193 (N_5193,N_4252,N_4064);
nand U5194 (N_5194,N_4150,N_4931);
or U5195 (N_5195,N_4906,N_4126);
nand U5196 (N_5196,N_4700,N_4146);
xor U5197 (N_5197,N_4280,N_4316);
nand U5198 (N_5198,N_4717,N_4662);
nor U5199 (N_5199,N_4796,N_4689);
nand U5200 (N_5200,N_4527,N_4393);
and U5201 (N_5201,N_4890,N_4575);
nand U5202 (N_5202,N_4623,N_4805);
nor U5203 (N_5203,N_4234,N_4425);
or U5204 (N_5204,N_4214,N_4051);
and U5205 (N_5205,N_4644,N_4765);
nor U5206 (N_5206,N_4225,N_4230);
and U5207 (N_5207,N_4186,N_4894);
nor U5208 (N_5208,N_4648,N_4666);
and U5209 (N_5209,N_4879,N_4932);
nor U5210 (N_5210,N_4125,N_4102);
xor U5211 (N_5211,N_4688,N_4757);
nand U5212 (N_5212,N_4012,N_4324);
or U5213 (N_5213,N_4943,N_4516);
or U5214 (N_5214,N_4674,N_4434);
or U5215 (N_5215,N_4194,N_4236);
nor U5216 (N_5216,N_4323,N_4382);
nor U5217 (N_5217,N_4374,N_4802);
nand U5218 (N_5218,N_4265,N_4556);
xnor U5219 (N_5219,N_4373,N_4558);
nand U5220 (N_5220,N_4979,N_4596);
or U5221 (N_5221,N_4412,N_4394);
and U5222 (N_5222,N_4039,N_4589);
and U5223 (N_5223,N_4285,N_4196);
nor U5224 (N_5224,N_4390,N_4946);
and U5225 (N_5225,N_4929,N_4795);
or U5226 (N_5226,N_4500,N_4266);
or U5227 (N_5227,N_4525,N_4987);
nor U5228 (N_5228,N_4259,N_4885);
nor U5229 (N_5229,N_4238,N_4785);
xor U5230 (N_5230,N_4046,N_4865);
nand U5231 (N_5231,N_4119,N_4874);
nor U5232 (N_5232,N_4507,N_4237);
and U5233 (N_5233,N_4376,N_4573);
nor U5234 (N_5234,N_4326,N_4464);
and U5235 (N_5235,N_4963,N_4197);
or U5236 (N_5236,N_4678,N_4404);
or U5237 (N_5237,N_4241,N_4761);
or U5238 (N_5238,N_4567,N_4930);
nor U5239 (N_5239,N_4960,N_4030);
nor U5240 (N_5240,N_4541,N_4664);
nand U5241 (N_5241,N_4730,N_4320);
and U5242 (N_5242,N_4372,N_4910);
or U5243 (N_5243,N_4137,N_4347);
and U5244 (N_5244,N_4510,N_4985);
nor U5245 (N_5245,N_4409,N_4713);
nand U5246 (N_5246,N_4120,N_4984);
and U5247 (N_5247,N_4304,N_4187);
xor U5248 (N_5248,N_4294,N_4049);
nor U5249 (N_5249,N_4248,N_4353);
xor U5250 (N_5250,N_4872,N_4949);
or U5251 (N_5251,N_4041,N_4724);
nor U5252 (N_5252,N_4744,N_4330);
nand U5253 (N_5253,N_4919,N_4065);
and U5254 (N_5254,N_4654,N_4290);
and U5255 (N_5255,N_4735,N_4553);
nor U5256 (N_5256,N_4994,N_4311);
nor U5257 (N_5257,N_4218,N_4219);
xor U5258 (N_5258,N_4363,N_4047);
nand U5259 (N_5259,N_4574,N_4048);
and U5260 (N_5260,N_4896,N_4800);
or U5261 (N_5261,N_4667,N_4058);
or U5262 (N_5262,N_4637,N_4315);
nor U5263 (N_5263,N_4164,N_4288);
nor U5264 (N_5264,N_4891,N_4085);
nor U5265 (N_5265,N_4934,N_4038);
nand U5266 (N_5266,N_4506,N_4400);
or U5267 (N_5267,N_4711,N_4838);
nand U5268 (N_5268,N_4560,N_4448);
or U5269 (N_5269,N_4019,N_4001);
nor U5270 (N_5270,N_4403,N_4972);
xnor U5271 (N_5271,N_4957,N_4081);
nor U5272 (N_5272,N_4615,N_4583);
nor U5273 (N_5273,N_4451,N_4568);
nor U5274 (N_5274,N_4803,N_4418);
nor U5275 (N_5275,N_4843,N_4752);
and U5276 (N_5276,N_4427,N_4612);
nand U5277 (N_5277,N_4956,N_4134);
and U5278 (N_5278,N_4122,N_4024);
nand U5279 (N_5279,N_4888,N_4042);
xor U5280 (N_5280,N_4970,N_4336);
and U5281 (N_5281,N_4665,N_4114);
or U5282 (N_5282,N_4743,N_4858);
and U5283 (N_5283,N_4927,N_4783);
nand U5284 (N_5284,N_4091,N_4806);
nor U5285 (N_5285,N_4142,N_4014);
nand U5286 (N_5286,N_4015,N_4991);
nand U5287 (N_5287,N_4768,N_4383);
nand U5288 (N_5288,N_4052,N_4210);
and U5289 (N_5289,N_4441,N_4301);
and U5290 (N_5290,N_4741,N_4585);
nor U5291 (N_5291,N_4053,N_4836);
and U5292 (N_5292,N_4572,N_4159);
and U5293 (N_5293,N_4503,N_4950);
and U5294 (N_5294,N_4686,N_4968);
nor U5295 (N_5295,N_4986,N_4798);
nor U5296 (N_5296,N_4738,N_4728);
and U5297 (N_5297,N_4835,N_4989);
nor U5298 (N_5298,N_4337,N_4056);
or U5299 (N_5299,N_4610,N_4669);
xnor U5300 (N_5300,N_4813,N_4999);
and U5301 (N_5301,N_4859,N_4396);
nor U5302 (N_5302,N_4687,N_4216);
and U5303 (N_5303,N_4408,N_4300);
nand U5304 (N_5304,N_4726,N_4489);
nor U5305 (N_5305,N_4339,N_4175);
and U5306 (N_5306,N_4286,N_4401);
or U5307 (N_5307,N_4721,N_4497);
xor U5308 (N_5308,N_4115,N_4753);
or U5309 (N_5309,N_4693,N_4707);
xnor U5310 (N_5310,N_4453,N_4392);
or U5311 (N_5311,N_4745,N_4941);
nor U5312 (N_5312,N_4034,N_4656);
nor U5313 (N_5313,N_4907,N_4966);
and U5314 (N_5314,N_4246,N_4948);
and U5315 (N_5315,N_4597,N_4331);
or U5316 (N_5316,N_4898,N_4832);
or U5317 (N_5317,N_4720,N_4029);
nand U5318 (N_5318,N_4157,N_4840);
or U5319 (N_5319,N_4240,N_4437);
or U5320 (N_5320,N_4559,N_4846);
nand U5321 (N_5321,N_4112,N_4718);
or U5322 (N_5322,N_4760,N_4577);
xnor U5323 (N_5323,N_4199,N_4430);
nor U5324 (N_5324,N_4096,N_4545);
and U5325 (N_5325,N_4482,N_4578);
nand U5326 (N_5326,N_4043,N_4710);
nand U5327 (N_5327,N_4087,N_4978);
or U5328 (N_5328,N_4200,N_4652);
or U5329 (N_5329,N_4077,N_4433);
nor U5330 (N_5330,N_4379,N_4546);
or U5331 (N_5331,N_4060,N_4054);
nor U5332 (N_5332,N_4552,N_4679);
nor U5333 (N_5333,N_4974,N_4309);
nand U5334 (N_5334,N_4776,N_4844);
and U5335 (N_5335,N_4699,N_4501);
nand U5336 (N_5336,N_4549,N_4547);
and U5337 (N_5337,N_4551,N_4417);
and U5338 (N_5338,N_4531,N_4100);
nand U5339 (N_5339,N_4828,N_4143);
nor U5340 (N_5340,N_4845,N_4036);
and U5341 (N_5341,N_4685,N_4083);
and U5342 (N_5342,N_4477,N_4452);
xnor U5343 (N_5343,N_4045,N_4936);
nand U5344 (N_5344,N_4365,N_4775);
nor U5345 (N_5345,N_4254,N_4550);
nand U5346 (N_5346,N_4937,N_4479);
and U5347 (N_5347,N_4600,N_4364);
and U5348 (N_5348,N_4106,N_4147);
xnor U5349 (N_5349,N_4450,N_4779);
nand U5350 (N_5350,N_4032,N_4456);
nand U5351 (N_5351,N_4619,N_4762);
or U5352 (N_5352,N_4640,N_4631);
nand U5353 (N_5353,N_4415,N_4367);
or U5354 (N_5354,N_4332,N_4542);
or U5355 (N_5355,N_4249,N_4117);
nand U5356 (N_5356,N_4912,N_4953);
nor U5357 (N_5357,N_4834,N_4129);
nor U5358 (N_5358,N_4514,N_4402);
or U5359 (N_5359,N_4893,N_4901);
nor U5360 (N_5360,N_4657,N_4554);
and U5361 (N_5361,N_4103,N_4443);
xnor U5362 (N_5362,N_4343,N_4037);
nor U5363 (N_5363,N_4136,N_4515);
and U5364 (N_5364,N_4998,N_4580);
nand U5365 (N_5365,N_4291,N_4335);
or U5366 (N_5366,N_4490,N_4183);
and U5367 (N_5367,N_4692,N_4921);
or U5368 (N_5368,N_4557,N_4526);
xnor U5369 (N_5369,N_4926,N_4257);
nand U5370 (N_5370,N_4438,N_4475);
or U5371 (N_5371,N_4377,N_4847);
or U5372 (N_5372,N_4295,N_4148);
and U5373 (N_5373,N_4299,N_4003);
nor U5374 (N_5374,N_4564,N_4020);
xnor U5375 (N_5375,N_4703,N_4267);
and U5376 (N_5376,N_4145,N_4062);
xor U5377 (N_5377,N_4413,N_4074);
and U5378 (N_5378,N_4705,N_4271);
xor U5379 (N_5379,N_4863,N_4833);
nand U5380 (N_5380,N_4869,N_4569);
nand U5381 (N_5381,N_4156,N_4469);
nor U5382 (N_5382,N_4188,N_4124);
nor U5383 (N_5383,N_4093,N_4539);
and U5384 (N_5384,N_4215,N_4536);
nand U5385 (N_5385,N_4245,N_4476);
nand U5386 (N_5386,N_4809,N_4110);
and U5387 (N_5387,N_4543,N_4715);
nand U5388 (N_5388,N_4622,N_4262);
and U5389 (N_5389,N_4962,N_4810);
nor U5390 (N_5390,N_4341,N_4361);
nand U5391 (N_5391,N_4837,N_4915);
nand U5392 (N_5392,N_4008,N_4279);
nor U5393 (N_5393,N_4877,N_4445);
and U5394 (N_5394,N_4161,N_4595);
xnor U5395 (N_5395,N_4864,N_4861);
or U5396 (N_5396,N_4821,N_4059);
or U5397 (N_5397,N_4255,N_4629);
nor U5398 (N_5398,N_4533,N_4854);
or U5399 (N_5399,N_4239,N_4422);
or U5400 (N_5400,N_4131,N_4261);
nand U5401 (N_5401,N_4889,N_4399);
or U5402 (N_5402,N_4736,N_4997);
xor U5403 (N_5403,N_4338,N_4920);
nor U5404 (N_5404,N_4340,N_4895);
xnor U5405 (N_5405,N_4528,N_4202);
or U5406 (N_5406,N_4875,N_4116);
nor U5407 (N_5407,N_4918,N_4841);
or U5408 (N_5408,N_4395,N_4650);
or U5409 (N_5409,N_4483,N_4268);
or U5410 (N_5410,N_4344,N_4004);
or U5411 (N_5411,N_4586,N_4801);
nand U5412 (N_5412,N_4105,N_4908);
xor U5413 (N_5413,N_4681,N_4782);
nand U5414 (N_5414,N_4561,N_4582);
nor U5415 (N_5415,N_4426,N_4203);
nor U5416 (N_5416,N_4675,N_4576);
or U5417 (N_5417,N_4850,N_4494);
nor U5418 (N_5418,N_4499,N_4163);
and U5419 (N_5419,N_4369,N_4079);
and U5420 (N_5420,N_4358,N_4613);
nand U5421 (N_5421,N_4694,N_4319);
or U5422 (N_5422,N_4095,N_4130);
nor U5423 (N_5423,N_4604,N_4584);
nor U5424 (N_5424,N_4601,N_4621);
nand U5425 (N_5425,N_4040,N_4523);
or U5426 (N_5426,N_4808,N_4342);
or U5427 (N_5427,N_4088,N_4457);
nor U5428 (N_5428,N_4924,N_4428);
nand U5429 (N_5429,N_4229,N_4385);
nand U5430 (N_5430,N_4759,N_4223);
xnor U5431 (N_5431,N_4192,N_4094);
and U5432 (N_5432,N_4387,N_4269);
xor U5433 (N_5433,N_4076,N_4899);
and U5434 (N_5434,N_4303,N_4807);
nand U5435 (N_5435,N_4221,N_4712);
and U5436 (N_5436,N_4419,N_4902);
and U5437 (N_5437,N_4829,N_4166);
or U5438 (N_5438,N_4598,N_4742);
and U5439 (N_5439,N_4090,N_4247);
nor U5440 (N_5440,N_4109,N_4892);
nor U5441 (N_5441,N_4521,N_4599);
nand U5442 (N_5442,N_4035,N_4764);
and U5443 (N_5443,N_4839,N_4152);
and U5444 (N_5444,N_4061,N_4792);
and U5445 (N_5445,N_4206,N_4381);
and U5446 (N_5446,N_4826,N_4075);
nand U5447 (N_5447,N_4444,N_4880);
and U5448 (N_5448,N_4002,N_4605);
and U5449 (N_5449,N_4668,N_4697);
and U5450 (N_5450,N_4386,N_4897);
or U5451 (N_5451,N_4555,N_4684);
nand U5452 (N_5452,N_4733,N_4446);
nor U5453 (N_5453,N_4440,N_4508);
or U5454 (N_5454,N_4272,N_4411);
nand U5455 (N_5455,N_4677,N_4016);
xnor U5456 (N_5456,N_4739,N_4317);
xnor U5457 (N_5457,N_4603,N_4011);
nand U5458 (N_5458,N_4355,N_4293);
nor U5459 (N_5459,N_4565,N_4633);
or U5460 (N_5460,N_4641,N_4162);
nand U5461 (N_5461,N_4520,N_4368);
and U5462 (N_5462,N_4375,N_4988);
xor U5463 (N_5463,N_4000,N_4964);
nand U5464 (N_5464,N_4135,N_4935);
and U5465 (N_5465,N_4682,N_4282);
nor U5466 (N_5466,N_4260,N_4167);
nand U5467 (N_5467,N_4360,N_4201);
nor U5468 (N_5468,N_4737,N_4471);
xnor U5469 (N_5469,N_4233,N_4634);
or U5470 (N_5470,N_4780,N_4616);
or U5471 (N_5471,N_4140,N_4887);
and U5472 (N_5472,N_4491,N_4470);
nand U5473 (N_5473,N_4354,N_4101);
nor U5474 (N_5474,N_4530,N_4993);
nor U5475 (N_5475,N_4756,N_4027);
xor U5476 (N_5476,N_4370,N_4181);
or U5477 (N_5477,N_4406,N_4069);
nand U5478 (N_5478,N_4429,N_4459);
or U5479 (N_5479,N_4380,N_4480);
nand U5480 (N_5480,N_4750,N_4624);
xnor U5481 (N_5481,N_4658,N_4256);
nor U5482 (N_5482,N_4086,N_4481);
or U5483 (N_5483,N_4886,N_4310);
nand U5484 (N_5484,N_4870,N_4566);
or U5485 (N_5485,N_4980,N_4747);
and U5486 (N_5486,N_4208,N_4593);
nor U5487 (N_5487,N_4671,N_4904);
and U5488 (N_5488,N_4174,N_4977);
or U5489 (N_5489,N_4702,N_4067);
nand U5490 (N_5490,N_4638,N_4080);
and U5491 (N_5491,N_4185,N_4173);
nor U5492 (N_5492,N_4044,N_4771);
and U5493 (N_5493,N_4133,N_4431);
or U5494 (N_5494,N_4708,N_4732);
and U5495 (N_5495,N_4345,N_4447);
or U5496 (N_5496,N_4205,N_4628);
nor U5497 (N_5497,N_4473,N_4318);
or U5498 (N_5498,N_4021,N_4179);
nor U5499 (N_5499,N_4184,N_4938);
nor U5500 (N_5500,N_4094,N_4058);
nor U5501 (N_5501,N_4200,N_4830);
nor U5502 (N_5502,N_4000,N_4751);
nand U5503 (N_5503,N_4972,N_4292);
or U5504 (N_5504,N_4991,N_4629);
or U5505 (N_5505,N_4422,N_4671);
and U5506 (N_5506,N_4122,N_4924);
nor U5507 (N_5507,N_4751,N_4770);
nand U5508 (N_5508,N_4892,N_4677);
and U5509 (N_5509,N_4219,N_4489);
xnor U5510 (N_5510,N_4699,N_4194);
nor U5511 (N_5511,N_4297,N_4777);
nor U5512 (N_5512,N_4262,N_4684);
or U5513 (N_5513,N_4093,N_4508);
or U5514 (N_5514,N_4811,N_4538);
nor U5515 (N_5515,N_4995,N_4144);
nand U5516 (N_5516,N_4284,N_4554);
nor U5517 (N_5517,N_4797,N_4996);
and U5518 (N_5518,N_4183,N_4838);
nor U5519 (N_5519,N_4904,N_4609);
or U5520 (N_5520,N_4191,N_4505);
nand U5521 (N_5521,N_4541,N_4095);
or U5522 (N_5522,N_4831,N_4466);
or U5523 (N_5523,N_4505,N_4103);
and U5524 (N_5524,N_4318,N_4706);
nor U5525 (N_5525,N_4561,N_4931);
xor U5526 (N_5526,N_4409,N_4210);
nor U5527 (N_5527,N_4313,N_4018);
nor U5528 (N_5528,N_4708,N_4145);
and U5529 (N_5529,N_4138,N_4211);
or U5530 (N_5530,N_4278,N_4769);
or U5531 (N_5531,N_4807,N_4453);
or U5532 (N_5532,N_4198,N_4712);
nor U5533 (N_5533,N_4212,N_4981);
or U5534 (N_5534,N_4497,N_4856);
nor U5535 (N_5535,N_4833,N_4376);
and U5536 (N_5536,N_4308,N_4345);
and U5537 (N_5537,N_4853,N_4186);
nor U5538 (N_5538,N_4122,N_4145);
nor U5539 (N_5539,N_4298,N_4539);
nor U5540 (N_5540,N_4761,N_4680);
nand U5541 (N_5541,N_4302,N_4962);
and U5542 (N_5542,N_4030,N_4152);
nand U5543 (N_5543,N_4647,N_4274);
or U5544 (N_5544,N_4366,N_4396);
or U5545 (N_5545,N_4742,N_4727);
or U5546 (N_5546,N_4377,N_4457);
xnor U5547 (N_5547,N_4712,N_4959);
xor U5548 (N_5548,N_4880,N_4509);
nand U5549 (N_5549,N_4885,N_4920);
or U5550 (N_5550,N_4433,N_4409);
or U5551 (N_5551,N_4968,N_4561);
and U5552 (N_5552,N_4428,N_4990);
or U5553 (N_5553,N_4997,N_4075);
and U5554 (N_5554,N_4864,N_4357);
and U5555 (N_5555,N_4198,N_4917);
xnor U5556 (N_5556,N_4638,N_4033);
xnor U5557 (N_5557,N_4826,N_4922);
and U5558 (N_5558,N_4593,N_4034);
and U5559 (N_5559,N_4597,N_4258);
and U5560 (N_5560,N_4213,N_4537);
or U5561 (N_5561,N_4082,N_4959);
or U5562 (N_5562,N_4851,N_4496);
nand U5563 (N_5563,N_4296,N_4919);
nand U5564 (N_5564,N_4115,N_4869);
and U5565 (N_5565,N_4478,N_4544);
and U5566 (N_5566,N_4230,N_4312);
and U5567 (N_5567,N_4852,N_4410);
or U5568 (N_5568,N_4888,N_4521);
nor U5569 (N_5569,N_4347,N_4151);
nand U5570 (N_5570,N_4466,N_4032);
xnor U5571 (N_5571,N_4584,N_4911);
or U5572 (N_5572,N_4625,N_4236);
nand U5573 (N_5573,N_4841,N_4464);
nand U5574 (N_5574,N_4102,N_4457);
or U5575 (N_5575,N_4948,N_4260);
and U5576 (N_5576,N_4606,N_4320);
nand U5577 (N_5577,N_4045,N_4726);
or U5578 (N_5578,N_4121,N_4449);
nand U5579 (N_5579,N_4851,N_4417);
nor U5580 (N_5580,N_4659,N_4332);
or U5581 (N_5581,N_4176,N_4168);
nand U5582 (N_5582,N_4718,N_4372);
nor U5583 (N_5583,N_4314,N_4934);
nand U5584 (N_5584,N_4211,N_4371);
nand U5585 (N_5585,N_4411,N_4312);
nor U5586 (N_5586,N_4083,N_4570);
and U5587 (N_5587,N_4779,N_4009);
nand U5588 (N_5588,N_4104,N_4873);
nor U5589 (N_5589,N_4119,N_4696);
nand U5590 (N_5590,N_4739,N_4721);
nand U5591 (N_5591,N_4904,N_4570);
or U5592 (N_5592,N_4247,N_4153);
and U5593 (N_5593,N_4826,N_4705);
nand U5594 (N_5594,N_4965,N_4238);
or U5595 (N_5595,N_4520,N_4786);
or U5596 (N_5596,N_4444,N_4832);
xor U5597 (N_5597,N_4584,N_4246);
nor U5598 (N_5598,N_4891,N_4953);
and U5599 (N_5599,N_4138,N_4743);
nor U5600 (N_5600,N_4971,N_4674);
nand U5601 (N_5601,N_4565,N_4033);
and U5602 (N_5602,N_4444,N_4626);
and U5603 (N_5603,N_4128,N_4300);
or U5604 (N_5604,N_4065,N_4015);
or U5605 (N_5605,N_4888,N_4190);
xor U5606 (N_5606,N_4456,N_4685);
and U5607 (N_5607,N_4249,N_4870);
or U5608 (N_5608,N_4478,N_4584);
nand U5609 (N_5609,N_4352,N_4340);
nand U5610 (N_5610,N_4068,N_4269);
or U5611 (N_5611,N_4754,N_4272);
or U5612 (N_5612,N_4711,N_4745);
nor U5613 (N_5613,N_4252,N_4144);
nor U5614 (N_5614,N_4382,N_4857);
nand U5615 (N_5615,N_4407,N_4007);
nand U5616 (N_5616,N_4662,N_4740);
or U5617 (N_5617,N_4047,N_4596);
or U5618 (N_5618,N_4224,N_4656);
nand U5619 (N_5619,N_4380,N_4164);
nor U5620 (N_5620,N_4675,N_4057);
nand U5621 (N_5621,N_4395,N_4233);
nand U5622 (N_5622,N_4135,N_4482);
and U5623 (N_5623,N_4661,N_4423);
or U5624 (N_5624,N_4075,N_4514);
nor U5625 (N_5625,N_4444,N_4904);
or U5626 (N_5626,N_4122,N_4840);
xnor U5627 (N_5627,N_4965,N_4432);
nor U5628 (N_5628,N_4701,N_4284);
or U5629 (N_5629,N_4682,N_4089);
xor U5630 (N_5630,N_4176,N_4924);
or U5631 (N_5631,N_4140,N_4298);
nor U5632 (N_5632,N_4340,N_4355);
xnor U5633 (N_5633,N_4837,N_4397);
and U5634 (N_5634,N_4545,N_4768);
or U5635 (N_5635,N_4000,N_4326);
nand U5636 (N_5636,N_4155,N_4078);
and U5637 (N_5637,N_4736,N_4407);
nand U5638 (N_5638,N_4983,N_4596);
nand U5639 (N_5639,N_4505,N_4782);
and U5640 (N_5640,N_4434,N_4018);
nor U5641 (N_5641,N_4220,N_4491);
xor U5642 (N_5642,N_4103,N_4345);
and U5643 (N_5643,N_4748,N_4091);
nor U5644 (N_5644,N_4170,N_4066);
nor U5645 (N_5645,N_4288,N_4294);
or U5646 (N_5646,N_4318,N_4484);
nor U5647 (N_5647,N_4393,N_4003);
xnor U5648 (N_5648,N_4637,N_4137);
or U5649 (N_5649,N_4473,N_4404);
or U5650 (N_5650,N_4617,N_4710);
or U5651 (N_5651,N_4128,N_4490);
and U5652 (N_5652,N_4970,N_4980);
or U5653 (N_5653,N_4421,N_4498);
or U5654 (N_5654,N_4186,N_4338);
xnor U5655 (N_5655,N_4607,N_4289);
xor U5656 (N_5656,N_4476,N_4444);
and U5657 (N_5657,N_4299,N_4064);
or U5658 (N_5658,N_4535,N_4376);
nor U5659 (N_5659,N_4034,N_4209);
or U5660 (N_5660,N_4558,N_4177);
nor U5661 (N_5661,N_4236,N_4265);
or U5662 (N_5662,N_4390,N_4603);
nor U5663 (N_5663,N_4167,N_4168);
nand U5664 (N_5664,N_4581,N_4901);
and U5665 (N_5665,N_4932,N_4709);
and U5666 (N_5666,N_4114,N_4377);
nor U5667 (N_5667,N_4466,N_4315);
nand U5668 (N_5668,N_4209,N_4510);
and U5669 (N_5669,N_4850,N_4978);
nor U5670 (N_5670,N_4907,N_4204);
or U5671 (N_5671,N_4913,N_4888);
nand U5672 (N_5672,N_4860,N_4757);
nand U5673 (N_5673,N_4439,N_4657);
nand U5674 (N_5674,N_4378,N_4441);
nand U5675 (N_5675,N_4767,N_4922);
xor U5676 (N_5676,N_4236,N_4604);
or U5677 (N_5677,N_4973,N_4076);
nor U5678 (N_5678,N_4823,N_4878);
and U5679 (N_5679,N_4563,N_4810);
xnor U5680 (N_5680,N_4325,N_4927);
and U5681 (N_5681,N_4918,N_4458);
xnor U5682 (N_5682,N_4939,N_4866);
or U5683 (N_5683,N_4146,N_4811);
nor U5684 (N_5684,N_4678,N_4778);
or U5685 (N_5685,N_4902,N_4206);
and U5686 (N_5686,N_4985,N_4122);
and U5687 (N_5687,N_4411,N_4721);
xor U5688 (N_5688,N_4630,N_4016);
or U5689 (N_5689,N_4217,N_4759);
nand U5690 (N_5690,N_4729,N_4490);
nand U5691 (N_5691,N_4497,N_4640);
and U5692 (N_5692,N_4825,N_4112);
nand U5693 (N_5693,N_4060,N_4986);
xor U5694 (N_5694,N_4150,N_4596);
nor U5695 (N_5695,N_4510,N_4674);
nor U5696 (N_5696,N_4305,N_4392);
nand U5697 (N_5697,N_4441,N_4055);
and U5698 (N_5698,N_4045,N_4789);
or U5699 (N_5699,N_4107,N_4839);
or U5700 (N_5700,N_4137,N_4851);
and U5701 (N_5701,N_4685,N_4300);
or U5702 (N_5702,N_4016,N_4100);
nand U5703 (N_5703,N_4334,N_4669);
or U5704 (N_5704,N_4198,N_4683);
nor U5705 (N_5705,N_4338,N_4240);
or U5706 (N_5706,N_4484,N_4501);
or U5707 (N_5707,N_4684,N_4729);
nand U5708 (N_5708,N_4336,N_4219);
nand U5709 (N_5709,N_4969,N_4787);
nand U5710 (N_5710,N_4943,N_4561);
nor U5711 (N_5711,N_4826,N_4185);
xor U5712 (N_5712,N_4151,N_4499);
xor U5713 (N_5713,N_4186,N_4485);
nor U5714 (N_5714,N_4211,N_4787);
or U5715 (N_5715,N_4780,N_4271);
nor U5716 (N_5716,N_4730,N_4814);
nand U5717 (N_5717,N_4624,N_4039);
and U5718 (N_5718,N_4997,N_4350);
nand U5719 (N_5719,N_4171,N_4281);
nor U5720 (N_5720,N_4897,N_4791);
nor U5721 (N_5721,N_4708,N_4974);
and U5722 (N_5722,N_4136,N_4360);
nor U5723 (N_5723,N_4594,N_4531);
or U5724 (N_5724,N_4288,N_4880);
and U5725 (N_5725,N_4469,N_4031);
nand U5726 (N_5726,N_4122,N_4811);
or U5727 (N_5727,N_4852,N_4451);
or U5728 (N_5728,N_4850,N_4277);
nor U5729 (N_5729,N_4704,N_4021);
and U5730 (N_5730,N_4437,N_4930);
nor U5731 (N_5731,N_4514,N_4836);
xnor U5732 (N_5732,N_4734,N_4666);
and U5733 (N_5733,N_4924,N_4242);
nand U5734 (N_5734,N_4834,N_4671);
nor U5735 (N_5735,N_4669,N_4799);
xnor U5736 (N_5736,N_4324,N_4676);
nand U5737 (N_5737,N_4883,N_4175);
and U5738 (N_5738,N_4132,N_4916);
or U5739 (N_5739,N_4682,N_4604);
and U5740 (N_5740,N_4520,N_4718);
xnor U5741 (N_5741,N_4335,N_4617);
nand U5742 (N_5742,N_4977,N_4861);
and U5743 (N_5743,N_4442,N_4400);
xnor U5744 (N_5744,N_4115,N_4382);
xnor U5745 (N_5745,N_4391,N_4138);
or U5746 (N_5746,N_4620,N_4065);
or U5747 (N_5747,N_4436,N_4356);
nand U5748 (N_5748,N_4795,N_4434);
and U5749 (N_5749,N_4366,N_4865);
xnor U5750 (N_5750,N_4712,N_4347);
nor U5751 (N_5751,N_4653,N_4143);
nand U5752 (N_5752,N_4052,N_4874);
or U5753 (N_5753,N_4414,N_4562);
or U5754 (N_5754,N_4530,N_4027);
xnor U5755 (N_5755,N_4610,N_4933);
or U5756 (N_5756,N_4059,N_4881);
and U5757 (N_5757,N_4191,N_4957);
nand U5758 (N_5758,N_4264,N_4289);
and U5759 (N_5759,N_4445,N_4549);
nor U5760 (N_5760,N_4890,N_4665);
and U5761 (N_5761,N_4877,N_4734);
nand U5762 (N_5762,N_4030,N_4679);
or U5763 (N_5763,N_4775,N_4097);
and U5764 (N_5764,N_4593,N_4512);
nor U5765 (N_5765,N_4011,N_4273);
nor U5766 (N_5766,N_4289,N_4584);
nor U5767 (N_5767,N_4510,N_4863);
nand U5768 (N_5768,N_4331,N_4534);
nor U5769 (N_5769,N_4661,N_4035);
and U5770 (N_5770,N_4146,N_4025);
or U5771 (N_5771,N_4300,N_4063);
nand U5772 (N_5772,N_4508,N_4652);
nand U5773 (N_5773,N_4123,N_4651);
or U5774 (N_5774,N_4576,N_4534);
and U5775 (N_5775,N_4851,N_4450);
nor U5776 (N_5776,N_4774,N_4600);
nor U5777 (N_5777,N_4576,N_4075);
nand U5778 (N_5778,N_4756,N_4985);
and U5779 (N_5779,N_4356,N_4814);
nand U5780 (N_5780,N_4960,N_4753);
or U5781 (N_5781,N_4964,N_4090);
nand U5782 (N_5782,N_4807,N_4590);
nand U5783 (N_5783,N_4101,N_4530);
nor U5784 (N_5784,N_4174,N_4501);
nor U5785 (N_5785,N_4293,N_4307);
and U5786 (N_5786,N_4323,N_4318);
and U5787 (N_5787,N_4407,N_4439);
and U5788 (N_5788,N_4298,N_4483);
nand U5789 (N_5789,N_4502,N_4441);
or U5790 (N_5790,N_4001,N_4003);
or U5791 (N_5791,N_4908,N_4317);
nand U5792 (N_5792,N_4305,N_4301);
or U5793 (N_5793,N_4957,N_4385);
or U5794 (N_5794,N_4154,N_4041);
nor U5795 (N_5795,N_4487,N_4514);
and U5796 (N_5796,N_4429,N_4730);
or U5797 (N_5797,N_4779,N_4801);
nand U5798 (N_5798,N_4957,N_4526);
nand U5799 (N_5799,N_4574,N_4402);
and U5800 (N_5800,N_4727,N_4200);
xor U5801 (N_5801,N_4276,N_4631);
and U5802 (N_5802,N_4951,N_4541);
and U5803 (N_5803,N_4941,N_4761);
nor U5804 (N_5804,N_4268,N_4646);
or U5805 (N_5805,N_4527,N_4920);
nand U5806 (N_5806,N_4859,N_4673);
nand U5807 (N_5807,N_4155,N_4665);
nand U5808 (N_5808,N_4625,N_4090);
and U5809 (N_5809,N_4172,N_4844);
or U5810 (N_5810,N_4959,N_4830);
nor U5811 (N_5811,N_4374,N_4914);
nor U5812 (N_5812,N_4497,N_4929);
nor U5813 (N_5813,N_4175,N_4108);
nor U5814 (N_5814,N_4352,N_4259);
and U5815 (N_5815,N_4365,N_4134);
or U5816 (N_5816,N_4223,N_4063);
and U5817 (N_5817,N_4946,N_4979);
nand U5818 (N_5818,N_4019,N_4190);
or U5819 (N_5819,N_4684,N_4274);
and U5820 (N_5820,N_4347,N_4439);
or U5821 (N_5821,N_4054,N_4680);
nor U5822 (N_5822,N_4608,N_4578);
and U5823 (N_5823,N_4647,N_4817);
nor U5824 (N_5824,N_4532,N_4294);
or U5825 (N_5825,N_4007,N_4753);
nand U5826 (N_5826,N_4280,N_4502);
nor U5827 (N_5827,N_4645,N_4781);
or U5828 (N_5828,N_4247,N_4087);
or U5829 (N_5829,N_4222,N_4370);
nor U5830 (N_5830,N_4129,N_4534);
nand U5831 (N_5831,N_4666,N_4414);
nor U5832 (N_5832,N_4008,N_4268);
and U5833 (N_5833,N_4130,N_4552);
nand U5834 (N_5834,N_4953,N_4265);
and U5835 (N_5835,N_4665,N_4658);
nand U5836 (N_5836,N_4598,N_4019);
or U5837 (N_5837,N_4351,N_4134);
nor U5838 (N_5838,N_4520,N_4194);
xnor U5839 (N_5839,N_4235,N_4748);
and U5840 (N_5840,N_4240,N_4996);
nand U5841 (N_5841,N_4697,N_4452);
or U5842 (N_5842,N_4412,N_4603);
nand U5843 (N_5843,N_4274,N_4999);
nor U5844 (N_5844,N_4393,N_4753);
or U5845 (N_5845,N_4097,N_4423);
nor U5846 (N_5846,N_4278,N_4599);
and U5847 (N_5847,N_4583,N_4864);
and U5848 (N_5848,N_4263,N_4697);
nor U5849 (N_5849,N_4346,N_4387);
nor U5850 (N_5850,N_4655,N_4477);
and U5851 (N_5851,N_4977,N_4947);
or U5852 (N_5852,N_4450,N_4261);
nor U5853 (N_5853,N_4188,N_4013);
nor U5854 (N_5854,N_4780,N_4497);
or U5855 (N_5855,N_4736,N_4112);
nand U5856 (N_5856,N_4182,N_4114);
and U5857 (N_5857,N_4299,N_4725);
xnor U5858 (N_5858,N_4901,N_4716);
and U5859 (N_5859,N_4780,N_4381);
xnor U5860 (N_5860,N_4510,N_4215);
xnor U5861 (N_5861,N_4916,N_4510);
or U5862 (N_5862,N_4848,N_4431);
and U5863 (N_5863,N_4391,N_4100);
nor U5864 (N_5864,N_4296,N_4584);
nor U5865 (N_5865,N_4226,N_4983);
xnor U5866 (N_5866,N_4539,N_4188);
nand U5867 (N_5867,N_4578,N_4412);
and U5868 (N_5868,N_4854,N_4782);
nand U5869 (N_5869,N_4899,N_4060);
or U5870 (N_5870,N_4247,N_4755);
and U5871 (N_5871,N_4811,N_4975);
nor U5872 (N_5872,N_4704,N_4692);
nand U5873 (N_5873,N_4408,N_4916);
nor U5874 (N_5874,N_4086,N_4387);
nand U5875 (N_5875,N_4560,N_4796);
and U5876 (N_5876,N_4118,N_4930);
xnor U5877 (N_5877,N_4474,N_4284);
nand U5878 (N_5878,N_4910,N_4524);
and U5879 (N_5879,N_4063,N_4058);
and U5880 (N_5880,N_4026,N_4953);
or U5881 (N_5881,N_4627,N_4448);
nor U5882 (N_5882,N_4689,N_4941);
and U5883 (N_5883,N_4847,N_4611);
xor U5884 (N_5884,N_4442,N_4093);
nand U5885 (N_5885,N_4626,N_4807);
and U5886 (N_5886,N_4654,N_4108);
nand U5887 (N_5887,N_4264,N_4328);
nor U5888 (N_5888,N_4573,N_4219);
xnor U5889 (N_5889,N_4320,N_4162);
nand U5890 (N_5890,N_4122,N_4257);
nor U5891 (N_5891,N_4671,N_4052);
or U5892 (N_5892,N_4962,N_4352);
nor U5893 (N_5893,N_4880,N_4631);
or U5894 (N_5894,N_4475,N_4890);
or U5895 (N_5895,N_4984,N_4336);
and U5896 (N_5896,N_4955,N_4715);
xnor U5897 (N_5897,N_4286,N_4690);
nand U5898 (N_5898,N_4799,N_4240);
or U5899 (N_5899,N_4961,N_4091);
nand U5900 (N_5900,N_4385,N_4855);
nor U5901 (N_5901,N_4705,N_4827);
or U5902 (N_5902,N_4663,N_4281);
and U5903 (N_5903,N_4318,N_4697);
or U5904 (N_5904,N_4106,N_4803);
and U5905 (N_5905,N_4148,N_4048);
or U5906 (N_5906,N_4134,N_4308);
or U5907 (N_5907,N_4478,N_4060);
nand U5908 (N_5908,N_4728,N_4105);
xor U5909 (N_5909,N_4313,N_4689);
and U5910 (N_5910,N_4425,N_4101);
and U5911 (N_5911,N_4570,N_4364);
xor U5912 (N_5912,N_4472,N_4638);
nand U5913 (N_5913,N_4912,N_4355);
and U5914 (N_5914,N_4277,N_4703);
and U5915 (N_5915,N_4601,N_4038);
and U5916 (N_5916,N_4195,N_4918);
nand U5917 (N_5917,N_4433,N_4845);
nand U5918 (N_5918,N_4802,N_4616);
nand U5919 (N_5919,N_4617,N_4901);
or U5920 (N_5920,N_4925,N_4596);
and U5921 (N_5921,N_4729,N_4949);
nand U5922 (N_5922,N_4822,N_4063);
and U5923 (N_5923,N_4621,N_4877);
and U5924 (N_5924,N_4625,N_4819);
nand U5925 (N_5925,N_4222,N_4290);
nor U5926 (N_5926,N_4856,N_4523);
and U5927 (N_5927,N_4979,N_4333);
nor U5928 (N_5928,N_4431,N_4663);
nor U5929 (N_5929,N_4190,N_4168);
or U5930 (N_5930,N_4149,N_4003);
or U5931 (N_5931,N_4254,N_4572);
nor U5932 (N_5932,N_4671,N_4782);
nor U5933 (N_5933,N_4881,N_4113);
nand U5934 (N_5934,N_4766,N_4202);
nand U5935 (N_5935,N_4667,N_4513);
or U5936 (N_5936,N_4632,N_4828);
or U5937 (N_5937,N_4737,N_4599);
and U5938 (N_5938,N_4128,N_4380);
and U5939 (N_5939,N_4674,N_4259);
nor U5940 (N_5940,N_4707,N_4151);
nand U5941 (N_5941,N_4471,N_4402);
or U5942 (N_5942,N_4812,N_4392);
or U5943 (N_5943,N_4839,N_4037);
or U5944 (N_5944,N_4282,N_4865);
nor U5945 (N_5945,N_4311,N_4705);
nand U5946 (N_5946,N_4534,N_4242);
nor U5947 (N_5947,N_4919,N_4014);
and U5948 (N_5948,N_4828,N_4282);
nor U5949 (N_5949,N_4716,N_4717);
and U5950 (N_5950,N_4503,N_4142);
nand U5951 (N_5951,N_4273,N_4390);
nand U5952 (N_5952,N_4647,N_4225);
nand U5953 (N_5953,N_4638,N_4451);
or U5954 (N_5954,N_4902,N_4639);
nand U5955 (N_5955,N_4326,N_4060);
and U5956 (N_5956,N_4809,N_4933);
xor U5957 (N_5957,N_4854,N_4773);
nand U5958 (N_5958,N_4731,N_4368);
nand U5959 (N_5959,N_4706,N_4552);
nand U5960 (N_5960,N_4844,N_4165);
nand U5961 (N_5961,N_4355,N_4595);
and U5962 (N_5962,N_4587,N_4130);
or U5963 (N_5963,N_4664,N_4312);
nand U5964 (N_5964,N_4659,N_4001);
or U5965 (N_5965,N_4073,N_4533);
or U5966 (N_5966,N_4352,N_4767);
or U5967 (N_5967,N_4715,N_4572);
nor U5968 (N_5968,N_4192,N_4485);
and U5969 (N_5969,N_4979,N_4036);
nand U5970 (N_5970,N_4243,N_4751);
or U5971 (N_5971,N_4144,N_4800);
and U5972 (N_5972,N_4429,N_4191);
nor U5973 (N_5973,N_4503,N_4833);
and U5974 (N_5974,N_4495,N_4535);
or U5975 (N_5975,N_4464,N_4973);
nand U5976 (N_5976,N_4611,N_4979);
nor U5977 (N_5977,N_4683,N_4619);
or U5978 (N_5978,N_4170,N_4899);
nand U5979 (N_5979,N_4428,N_4906);
nor U5980 (N_5980,N_4557,N_4853);
or U5981 (N_5981,N_4062,N_4125);
or U5982 (N_5982,N_4997,N_4080);
and U5983 (N_5983,N_4137,N_4522);
or U5984 (N_5984,N_4466,N_4330);
and U5985 (N_5985,N_4027,N_4290);
nor U5986 (N_5986,N_4913,N_4137);
or U5987 (N_5987,N_4925,N_4939);
or U5988 (N_5988,N_4380,N_4140);
nand U5989 (N_5989,N_4380,N_4570);
nand U5990 (N_5990,N_4671,N_4364);
and U5991 (N_5991,N_4001,N_4704);
nor U5992 (N_5992,N_4849,N_4356);
nand U5993 (N_5993,N_4529,N_4780);
and U5994 (N_5994,N_4935,N_4892);
nand U5995 (N_5995,N_4563,N_4104);
nor U5996 (N_5996,N_4424,N_4061);
nor U5997 (N_5997,N_4847,N_4800);
and U5998 (N_5998,N_4802,N_4207);
xnor U5999 (N_5999,N_4396,N_4662);
and U6000 (N_6000,N_5121,N_5116);
nor U6001 (N_6001,N_5696,N_5286);
nand U6002 (N_6002,N_5647,N_5228);
and U6003 (N_6003,N_5347,N_5072);
and U6004 (N_6004,N_5161,N_5520);
and U6005 (N_6005,N_5113,N_5603);
and U6006 (N_6006,N_5948,N_5595);
or U6007 (N_6007,N_5170,N_5109);
nor U6008 (N_6008,N_5041,N_5049);
and U6009 (N_6009,N_5571,N_5877);
nor U6010 (N_6010,N_5568,N_5995);
nand U6011 (N_6011,N_5043,N_5446);
or U6012 (N_6012,N_5433,N_5269);
nor U6013 (N_6013,N_5962,N_5781);
and U6014 (N_6014,N_5892,N_5127);
and U6015 (N_6015,N_5429,N_5076);
nor U6016 (N_6016,N_5117,N_5312);
nand U6017 (N_6017,N_5472,N_5190);
or U6018 (N_6018,N_5832,N_5600);
and U6019 (N_6019,N_5066,N_5914);
nand U6020 (N_6020,N_5434,N_5275);
and U6021 (N_6021,N_5368,N_5421);
nand U6022 (N_6022,N_5662,N_5985);
nand U6023 (N_6023,N_5719,N_5863);
xnor U6024 (N_6024,N_5266,N_5592);
nand U6025 (N_6025,N_5742,N_5423);
or U6026 (N_6026,N_5739,N_5871);
xnor U6027 (N_6027,N_5375,N_5726);
and U6028 (N_6028,N_5240,N_5959);
nand U6029 (N_6029,N_5847,N_5417);
and U6030 (N_6030,N_5796,N_5627);
and U6031 (N_6031,N_5765,N_5015);
nor U6032 (N_6032,N_5316,N_5694);
nor U6033 (N_6033,N_5924,N_5654);
and U6034 (N_6034,N_5242,N_5083);
nor U6035 (N_6035,N_5912,N_5993);
nand U6036 (N_6036,N_5252,N_5369);
xnor U6037 (N_6037,N_5588,N_5510);
nor U6038 (N_6038,N_5887,N_5780);
or U6039 (N_6039,N_5606,N_5574);
nor U6040 (N_6040,N_5189,N_5343);
or U6041 (N_6041,N_5427,N_5966);
nand U6042 (N_6042,N_5063,N_5014);
nor U6043 (N_6043,N_5619,N_5178);
nand U6044 (N_6044,N_5512,N_5108);
or U6045 (N_6045,N_5837,N_5929);
or U6046 (N_6046,N_5990,N_5208);
or U6047 (N_6047,N_5907,N_5388);
or U6048 (N_6048,N_5750,N_5953);
and U6049 (N_6049,N_5707,N_5748);
or U6050 (N_6050,N_5743,N_5874);
nand U6051 (N_6051,N_5209,N_5261);
and U6052 (N_6052,N_5448,N_5068);
nor U6053 (N_6053,N_5257,N_5523);
and U6054 (N_6054,N_5771,N_5495);
and U6055 (N_6055,N_5975,N_5310);
nor U6056 (N_6056,N_5688,N_5908);
xnor U6057 (N_6057,N_5671,N_5853);
and U6058 (N_6058,N_5483,N_5809);
nor U6059 (N_6059,N_5082,N_5454);
and U6060 (N_6060,N_5415,N_5441);
nor U6061 (N_6061,N_5905,N_5033);
xnor U6062 (N_6062,N_5885,N_5406);
or U6063 (N_6063,N_5638,N_5136);
xor U6064 (N_6064,N_5509,N_5879);
or U6065 (N_6065,N_5770,N_5493);
nand U6066 (N_6066,N_5609,N_5449);
and U6067 (N_6067,N_5569,N_5143);
nor U6068 (N_6068,N_5410,N_5790);
or U6069 (N_6069,N_5235,N_5808);
nor U6070 (N_6070,N_5420,N_5535);
nand U6071 (N_6071,N_5515,N_5119);
nand U6072 (N_6072,N_5296,N_5154);
nor U6073 (N_6073,N_5830,N_5684);
and U6074 (N_6074,N_5802,N_5494);
nand U6075 (N_6075,N_5295,N_5164);
or U6076 (N_6076,N_5271,N_5792);
nand U6077 (N_6077,N_5691,N_5760);
or U6078 (N_6078,N_5020,N_5452);
nor U6079 (N_6079,N_5221,N_5336);
or U6080 (N_6080,N_5193,N_5361);
or U6081 (N_6081,N_5087,N_5156);
and U6082 (N_6082,N_5826,N_5645);
or U6083 (N_6083,N_5820,N_5047);
and U6084 (N_6084,N_5073,N_5777);
and U6085 (N_6085,N_5301,N_5868);
or U6086 (N_6086,N_5559,N_5167);
xor U6087 (N_6087,N_5475,N_5653);
nor U6088 (N_6088,N_5195,N_5218);
or U6089 (N_6089,N_5800,N_5002);
nor U6090 (N_6090,N_5498,N_5884);
nor U6091 (N_6091,N_5814,N_5216);
xor U6092 (N_6092,N_5931,N_5348);
nand U6093 (N_6093,N_5032,N_5057);
and U6094 (N_6094,N_5810,N_5008);
or U6095 (N_6095,N_5858,N_5545);
or U6096 (N_6096,N_5166,N_5185);
nand U6097 (N_6097,N_5560,N_5173);
and U6098 (N_6098,N_5786,N_5668);
nand U6099 (N_6099,N_5112,N_5430);
and U6100 (N_6100,N_5608,N_5612);
xor U6101 (N_6101,N_5815,N_5724);
and U6102 (N_6102,N_5673,N_5141);
xnor U6103 (N_6103,N_5764,N_5318);
and U6104 (N_6104,N_5327,N_5618);
nand U6105 (N_6105,N_5404,N_5756);
nand U6106 (N_6106,N_5980,N_5089);
xnor U6107 (N_6107,N_5539,N_5276);
or U6108 (N_6108,N_5284,N_5659);
xnor U6109 (N_6109,N_5122,N_5747);
nand U6110 (N_6110,N_5891,N_5660);
nor U6111 (N_6111,N_5181,N_5398);
nor U6112 (N_6112,N_5939,N_5784);
and U6113 (N_6113,N_5789,N_5075);
or U6114 (N_6114,N_5570,N_5675);
nor U6115 (N_6115,N_5320,N_5424);
and U6116 (N_6116,N_5442,N_5935);
and U6117 (N_6117,N_5744,N_5718);
nand U6118 (N_6118,N_5249,N_5870);
nand U6119 (N_6119,N_5947,N_5330);
nand U6120 (N_6120,N_5986,N_5150);
xor U6121 (N_6121,N_5840,N_5629);
and U6122 (N_6122,N_5299,N_5053);
nand U6123 (N_6123,N_5666,N_5944);
nand U6124 (N_6124,N_5363,N_5591);
nand U6125 (N_6125,N_5731,N_5182);
nand U6126 (N_6126,N_5146,N_5360);
or U6127 (N_6127,N_5613,N_5904);
xnor U6128 (N_6128,N_5147,N_5357);
nor U6129 (N_6129,N_5701,N_5699);
and U6130 (N_6130,N_5478,N_5517);
or U6131 (N_6131,N_5172,N_5321);
or U6132 (N_6132,N_5798,N_5951);
and U6133 (N_6133,N_5910,N_5359);
nand U6134 (N_6134,N_5916,N_5486);
or U6135 (N_6135,N_5665,N_5054);
nor U6136 (N_6136,N_5397,N_5833);
nand U6137 (N_6137,N_5855,N_5605);
nor U6138 (N_6138,N_5524,N_5381);
or U6139 (N_6139,N_5872,N_5499);
nand U6140 (N_6140,N_5395,N_5846);
nand U6141 (N_6141,N_5017,N_5695);
nand U6142 (N_6142,N_5546,N_5028);
nor U6143 (N_6143,N_5580,N_5497);
and U6144 (N_6144,N_5307,N_5945);
nand U6145 (N_6145,N_5680,N_5925);
xnor U6146 (N_6146,N_5543,N_5457);
and U6147 (N_6147,N_5233,N_5374);
or U6148 (N_6148,N_5186,N_5393);
xor U6149 (N_6149,N_5367,N_5344);
nor U6150 (N_6150,N_5576,N_5358);
nand U6151 (N_6151,N_5288,N_5090);
xnor U6152 (N_6152,N_5206,N_5729);
nand U6153 (N_6153,N_5268,N_5950);
nor U6154 (N_6154,N_5585,N_5056);
or U6155 (N_6155,N_5824,N_5354);
nor U6156 (N_6156,N_5876,N_5958);
nand U6157 (N_6157,N_5617,N_5835);
nand U6158 (N_6158,N_5414,N_5599);
or U6159 (N_6159,N_5079,N_5501);
nor U6160 (N_6160,N_5697,N_5260);
and U6161 (N_6161,N_5304,N_5010);
or U6162 (N_6162,N_5909,N_5283);
nand U6163 (N_6163,N_5727,N_5752);
nor U6164 (N_6164,N_5270,N_5487);
nand U6165 (N_6165,N_5812,N_5303);
nand U6166 (N_6166,N_5467,N_5223);
nor U6167 (N_6167,N_5065,N_5378);
nand U6168 (N_6168,N_5011,N_5519);
nor U6169 (N_6169,N_5992,N_5297);
nand U6170 (N_6170,N_5841,N_5251);
or U6171 (N_6171,N_5362,N_5540);
or U6172 (N_6172,N_5794,N_5708);
nor U6173 (N_6173,N_5716,N_5970);
xor U6174 (N_6174,N_5941,N_5715);
or U6175 (N_6175,N_5775,N_5596);
or U6176 (N_6176,N_5313,N_5031);
or U6177 (N_6177,N_5530,N_5394);
nor U6178 (N_6178,N_5086,N_5435);
and U6179 (N_6179,N_5881,N_5827);
and U6180 (N_6180,N_5412,N_5293);
nor U6181 (N_6181,N_5018,N_5633);
nand U6182 (N_6182,N_5721,N_5714);
nor U6183 (N_6183,N_5188,N_5019);
and U6184 (N_6184,N_5469,N_5215);
nand U6185 (N_6185,N_5758,N_5070);
nor U6186 (N_6186,N_5484,N_5507);
nor U6187 (N_6187,N_5176,N_5825);
and U6188 (N_6188,N_5438,N_5376);
and U6189 (N_6189,N_5128,N_5409);
or U6190 (N_6190,N_5542,N_5094);
nor U6191 (N_6191,N_5774,N_5131);
nor U6192 (N_6192,N_5883,N_5278);
xnor U6193 (N_6193,N_5844,N_5329);
xnor U6194 (N_6194,N_5803,N_5920);
nor U6195 (N_6195,N_5256,N_5700);
nor U6196 (N_6196,N_5839,N_5566);
or U6197 (N_6197,N_5021,N_5641);
or U6198 (N_6198,N_5811,N_5007);
nand U6199 (N_6199,N_5965,N_5254);
and U6200 (N_6200,N_5664,N_5772);
nor U6201 (N_6201,N_5594,N_5650);
or U6202 (N_6202,N_5500,N_5728);
and U6203 (N_6203,N_5804,N_5300);
nor U6204 (N_6204,N_5335,N_5503);
nor U6205 (N_6205,N_5624,N_5439);
and U6206 (N_6206,N_5287,N_5443);
nor U6207 (N_6207,N_5851,N_5149);
or U6208 (N_6208,N_5573,N_5042);
or U6209 (N_6209,N_5558,N_5129);
and U6210 (N_6210,N_5101,N_5759);
and U6211 (N_6211,N_5411,N_5528);
or U6212 (N_6212,N_5511,N_5746);
and U6213 (N_6213,N_5848,N_5705);
or U6214 (N_6214,N_5106,N_5140);
nand U6215 (N_6215,N_5198,N_5055);
nor U6216 (N_6216,N_5201,N_5064);
nand U6217 (N_6217,N_5207,N_5508);
or U6218 (N_6218,N_5126,N_5977);
nor U6219 (N_6219,N_5037,N_5999);
nor U6220 (N_6220,N_5898,N_5027);
xnor U6221 (N_6221,N_5972,N_5901);
or U6222 (N_6222,N_5952,N_5735);
xor U6223 (N_6223,N_5490,N_5960);
or U6224 (N_6224,N_5308,N_5567);
or U6225 (N_6225,N_5681,N_5949);
and U6226 (N_6226,N_5698,N_5579);
and U6227 (N_6227,N_5956,N_5187);
and U6228 (N_6228,N_5610,N_5139);
nand U6229 (N_6229,N_5946,N_5819);
or U6230 (N_6230,N_5290,N_5713);
or U6231 (N_6231,N_5062,N_5934);
nor U6232 (N_6232,N_5889,N_5482);
nand U6233 (N_6233,N_5620,N_5416);
nand U6234 (N_6234,N_5937,N_5074);
and U6235 (N_6235,N_5184,N_5604);
and U6236 (N_6236,N_5365,N_5776);
or U6237 (N_6237,N_5006,N_5737);
nor U6238 (N_6238,N_5936,N_5849);
nor U6239 (N_6239,N_5636,N_5036);
nand U6240 (N_6240,N_5103,N_5899);
nand U6241 (N_6241,N_5229,N_5882);
xor U6242 (N_6242,N_5547,N_5640);
and U6243 (N_6243,N_5954,N_5918);
nor U6244 (N_6244,N_5538,N_5403);
or U6245 (N_6245,N_5635,N_5125);
or U6246 (N_6246,N_5900,N_5943);
and U6247 (N_6247,N_5693,N_5464);
nor U6248 (N_6248,N_5687,N_5392);
nand U6249 (N_6249,N_5518,N_5413);
or U6250 (N_6250,N_5625,N_5023);
or U6251 (N_6251,N_5437,N_5529);
and U6252 (N_6252,N_5631,N_5473);
and U6253 (N_6253,N_5982,N_5720);
nand U6254 (N_6254,N_5204,N_5305);
nor U6255 (N_6255,N_5179,N_5130);
nor U6256 (N_6256,N_5753,N_5553);
nand U6257 (N_6257,N_5258,N_5259);
and U6258 (N_6258,N_5341,N_5401);
and U6259 (N_6259,N_5273,N_5351);
nor U6260 (N_6260,N_5667,N_5602);
xor U6261 (N_6261,N_5180,N_5340);
nor U6262 (N_6262,N_5194,N_5581);
and U6263 (N_6263,N_5859,N_5890);
or U6264 (N_6264,N_5525,N_5557);
nand U6265 (N_6265,N_5502,N_5440);
and U6266 (N_6266,N_5183,N_5092);
and U6267 (N_6267,N_5471,N_5552);
nand U6268 (N_6268,N_5339,N_5038);
or U6269 (N_6269,N_5657,N_5197);
nand U6270 (N_6270,N_5616,N_5102);
nand U6271 (N_6271,N_5372,N_5767);
nand U6272 (N_6272,N_5202,N_5292);
nand U6273 (N_6273,N_5024,N_5807);
nand U6274 (N_6274,N_5211,N_5455);
or U6275 (N_6275,N_5039,N_5245);
or U6276 (N_6276,N_5644,N_5768);
xor U6277 (N_6277,N_5477,N_5704);
and U6278 (N_6278,N_5740,N_5788);
nor U6279 (N_6279,N_5370,N_5799);
and U6280 (N_6280,N_5496,N_5782);
nor U6281 (N_6281,N_5199,N_5458);
and U6282 (N_6282,N_5264,N_5801);
xnor U6283 (N_6283,N_5058,N_5408);
nand U6284 (N_6284,N_5238,N_5778);
nand U6285 (N_6285,N_5445,N_5733);
nor U6286 (N_6286,N_5761,N_5717);
nor U6287 (N_6287,N_5096,N_5219);
or U6288 (N_6288,N_5793,N_5865);
or U6289 (N_6289,N_5513,N_5168);
and U6290 (N_6290,N_5867,N_5461);
or U6291 (N_6291,N_5725,N_5927);
nand U6292 (N_6292,N_5544,N_5669);
nor U6293 (N_6293,N_5224,N_5231);
and U6294 (N_6294,N_5142,N_5035);
and U6295 (N_6295,N_5353,N_5399);
nor U6296 (N_6296,N_5345,N_5896);
or U6297 (N_6297,N_5003,N_5137);
nand U6298 (N_6298,N_5236,N_5917);
nor U6299 (N_6299,N_5983,N_5279);
and U6300 (N_6300,N_5422,N_5026);
nor U6301 (N_6301,N_5730,N_5060);
and U6302 (N_6302,N_5813,N_5911);
nor U6303 (N_6303,N_5565,N_5895);
or U6304 (N_6304,N_5852,N_5674);
nor U6305 (N_6305,N_5751,N_5762);
nor U6306 (N_6306,N_5615,N_5611);
and U6307 (N_6307,N_5016,N_5506);
nand U6308 (N_6308,N_5856,N_5806);
nor U6309 (N_6309,N_5226,N_5391);
and U6310 (N_6310,N_5628,N_5466);
and U6311 (N_6311,N_5196,N_5536);
nor U6312 (N_6312,N_5658,N_5159);
and U6313 (N_6313,N_5816,N_5880);
and U6314 (N_6314,N_5621,N_5045);
nor U6315 (N_6315,N_5034,N_5319);
or U6316 (N_6316,N_5317,N_5785);
or U6317 (N_6317,N_5988,N_5243);
nand U6318 (N_6318,N_5325,N_5677);
or U6319 (N_6319,N_5736,N_5685);
and U6320 (N_6320,N_5648,N_5000);
and U6321 (N_6321,N_5474,N_5419);
nor U6322 (N_6322,N_5582,N_5373);
nand U6323 (N_6323,N_5331,N_5145);
nand U6324 (N_6324,N_5078,N_5652);
and U6325 (N_6325,N_5875,N_5428);
nand U6326 (N_6326,N_5583,N_5135);
nor U6327 (N_6327,N_5818,N_5151);
xor U6328 (N_6328,N_5564,N_5514);
nor U6329 (N_6329,N_5732,N_5124);
nor U6330 (N_6330,N_5886,N_5821);
and U6331 (N_6331,N_5174,N_5175);
xnor U6332 (N_6332,N_5133,N_5138);
nor U6333 (N_6333,N_5843,N_5459);
xnor U6334 (N_6334,N_5230,N_5144);
and U6335 (N_6335,N_5548,N_5250);
nand U6336 (N_6336,N_5930,N_5384);
or U6337 (N_6337,N_5614,N_5153);
and U6338 (N_6338,N_5479,N_5850);
and U6339 (N_6339,N_5118,N_5842);
nor U6340 (N_6340,N_5309,N_5333);
nor U6341 (N_6341,N_5971,N_5822);
xor U6342 (N_6342,N_5672,N_5551);
and U6343 (N_6343,N_5157,N_5649);
nand U6344 (N_6344,N_5248,N_5382);
nor U6345 (N_6345,N_5597,N_5561);
nor U6346 (N_6346,N_5212,N_5400);
or U6347 (N_6347,N_5244,N_5030);
and U6348 (N_6348,N_5622,N_5831);
nor U6349 (N_6349,N_5922,N_5091);
and U6350 (N_6350,N_5787,N_5081);
or U6351 (N_6351,N_5589,N_5389);
or U6352 (N_6352,N_5387,N_5294);
nor U6353 (N_6353,N_5526,N_5823);
xor U6354 (N_6354,N_5302,N_5040);
and U6355 (N_6355,N_5436,N_5556);
and U6356 (N_6356,N_5407,N_5104);
and U6357 (N_6357,N_5655,N_5749);
nor U6358 (N_6358,N_5763,N_5634);
or U6359 (N_6359,N_5134,N_5828);
or U6360 (N_6360,N_5338,N_5860);
xor U6361 (N_6361,N_5607,N_5969);
nor U6362 (N_6362,N_5651,N_5379);
xor U6363 (N_6363,N_5285,N_5791);
or U6364 (N_6364,N_5110,N_5342);
nor U6365 (N_6365,N_5637,N_5232);
and U6366 (N_6366,N_5915,N_5460);
nor U6367 (N_6367,N_5541,N_5861);
nand U6368 (N_6368,N_5085,N_5987);
nand U6369 (N_6369,N_5386,N_5456);
nor U6370 (N_6370,N_5396,N_5100);
nand U6371 (N_6371,N_5098,N_5690);
nor U6372 (N_6372,N_5095,N_5741);
or U6373 (N_6373,N_5205,N_5323);
or U6374 (N_6374,N_5451,N_5902);
and U6375 (N_6375,N_5111,N_5418);
or U6376 (N_6376,N_5702,N_5795);
nand U6377 (N_6377,N_5578,N_5996);
and U6378 (N_6378,N_5678,N_5431);
and U6379 (N_6379,N_5356,N_5994);
nand U6380 (N_6380,N_5575,N_5214);
or U6381 (N_6381,N_5324,N_5926);
and U6382 (N_6382,N_5314,N_5928);
and U6383 (N_6383,N_5754,N_5077);
and U6384 (N_6384,N_5080,N_5974);
and U6385 (N_6385,N_5282,N_5022);
xor U6386 (N_6386,N_5632,N_5405);
and U6387 (N_6387,N_5012,N_5377);
xor U6388 (N_6388,N_5864,N_5572);
nor U6389 (N_6389,N_5531,N_5274);
xnor U6390 (N_6390,N_5169,N_5380);
nor U6391 (N_6391,N_5088,N_5587);
or U6392 (N_6392,N_5964,N_5485);
or U6393 (N_6393,N_5402,N_5311);
nand U6394 (N_6394,N_5838,N_5371);
or U6395 (N_6395,N_5061,N_5998);
xnor U6396 (N_6396,N_5630,N_5586);
or U6397 (N_6397,N_5679,N_5955);
and U6398 (N_6398,N_5834,N_5326);
nand U6399 (N_6399,N_5683,N_5906);
or U6400 (N_6400,N_5480,N_5722);
and U6401 (N_6401,N_5048,N_5577);
or U6402 (N_6402,N_5470,N_5845);
and U6403 (N_6403,N_5527,N_5656);
nand U6404 (N_6404,N_5247,N_5554);
nor U6405 (N_6405,N_5281,N_5504);
and U6406 (N_6406,N_5967,N_5979);
and U6407 (N_6407,N_5385,N_5670);
nand U6408 (N_6408,N_5973,N_5352);
xnor U6409 (N_6409,N_5921,N_5981);
and U6410 (N_6410,N_5769,N_5562);
and U6411 (N_6411,N_5052,N_5105);
nand U6412 (N_6412,N_5488,N_5532);
nand U6413 (N_6413,N_5366,N_5069);
nand U6414 (N_6414,N_5328,N_5120);
nand U6415 (N_6415,N_5961,N_5267);
nor U6416 (N_6416,N_5155,N_5706);
and U6417 (N_6417,N_5099,N_5940);
nor U6418 (N_6418,N_5255,N_5593);
nor U6419 (N_6419,N_5162,N_5521);
and U6420 (N_6420,N_5160,N_5465);
or U6421 (N_6421,N_5280,N_5888);
nand U6422 (N_6422,N_5709,N_5976);
and U6423 (N_6423,N_5355,N_5676);
and U6424 (N_6424,N_5757,N_5783);
nand U6425 (N_6425,N_5067,N_5623);
nor U6426 (N_6426,N_5210,N_5710);
and U6427 (N_6427,N_5913,N_5097);
and U6428 (N_6428,N_5334,N_5584);
or U6429 (N_6429,N_5289,N_5059);
nand U6430 (N_6430,N_5265,N_5878);
nand U6431 (N_6431,N_5332,N_5234);
nor U6432 (N_6432,N_5723,N_5766);
xor U6433 (N_6433,N_5009,N_5453);
nand U6434 (N_6434,N_5817,N_5555);
nor U6435 (N_6435,N_5426,N_5491);
or U6436 (N_6436,N_5989,N_5114);
nor U6437 (N_6437,N_5854,N_5192);
xor U6438 (N_6438,N_5857,N_5692);
xnor U6439 (N_6439,N_5869,N_5163);
xor U6440 (N_6440,N_5225,N_5779);
nor U6441 (N_6441,N_5350,N_5957);
or U6442 (N_6442,N_5262,N_5712);
nor U6443 (N_6443,N_5963,N_5237);
nor U6444 (N_6444,N_5873,N_5991);
or U6445 (N_6445,N_5866,N_5123);
or U6446 (N_6446,N_5533,N_5703);
and U6447 (N_6447,N_5646,N_5191);
nand U6448 (N_6448,N_5601,N_5383);
xor U6449 (N_6449,N_5661,N_5829);
and U6450 (N_6450,N_5220,N_5932);
and U6451 (N_6451,N_5246,N_5241);
or U6452 (N_6452,N_5263,N_5462);
and U6453 (N_6453,N_5203,N_5306);
and U6454 (N_6454,N_5029,N_5450);
and U6455 (N_6455,N_5590,N_5938);
nand U6456 (N_6456,N_5227,N_5158);
xor U6457 (N_6457,N_5537,N_5978);
or U6458 (N_6458,N_5682,N_5004);
nor U6459 (N_6459,N_5346,N_5534);
nand U6460 (N_6460,N_5836,N_5797);
nor U6461 (N_6461,N_5689,N_5468);
and U6462 (N_6462,N_5492,N_5919);
nand U6463 (N_6463,N_5171,N_5046);
and U6464 (N_6464,N_5277,N_5432);
and U6465 (N_6465,N_5711,N_5071);
and U6466 (N_6466,N_5298,N_5148);
nor U6467 (N_6467,N_5755,N_5050);
nand U6468 (N_6468,N_5745,N_5115);
nand U6469 (N_6469,N_5903,N_5337);
and U6470 (N_6470,N_5177,N_5476);
and U6471 (N_6471,N_5322,N_5505);
and U6472 (N_6472,N_5222,N_5984);
or U6473 (N_6473,N_5862,N_5663);
or U6474 (N_6474,N_5349,N_5522);
nor U6475 (N_6475,N_5626,N_5643);
nor U6476 (N_6476,N_5942,N_5213);
or U6477 (N_6477,N_5217,N_5425);
nor U6478 (N_6478,N_5107,N_5894);
or U6479 (N_6479,N_5013,N_5390);
nand U6480 (N_6480,N_5549,N_5132);
xnor U6481 (N_6481,N_5550,N_5897);
and U6482 (N_6482,N_5093,N_5933);
xor U6483 (N_6483,N_5315,N_5152);
xnor U6484 (N_6484,N_5686,N_5165);
and U6485 (N_6485,N_5773,N_5001);
or U6486 (N_6486,N_5563,N_5444);
or U6487 (N_6487,N_5734,N_5291);
nor U6488 (N_6488,N_5200,N_5516);
and U6489 (N_6489,N_5044,N_5253);
and U6490 (N_6490,N_5051,N_5463);
nand U6491 (N_6491,N_5481,N_5005);
or U6492 (N_6492,N_5642,N_5923);
nand U6493 (N_6493,N_5489,N_5447);
and U6494 (N_6494,N_5738,N_5805);
nand U6495 (N_6495,N_5364,N_5272);
nand U6496 (N_6496,N_5997,N_5239);
nand U6497 (N_6497,N_5084,N_5598);
or U6498 (N_6498,N_5639,N_5025);
nand U6499 (N_6499,N_5893,N_5968);
nand U6500 (N_6500,N_5478,N_5157);
or U6501 (N_6501,N_5204,N_5373);
or U6502 (N_6502,N_5261,N_5057);
and U6503 (N_6503,N_5491,N_5231);
and U6504 (N_6504,N_5579,N_5228);
nand U6505 (N_6505,N_5651,N_5070);
and U6506 (N_6506,N_5001,N_5454);
nand U6507 (N_6507,N_5381,N_5049);
and U6508 (N_6508,N_5548,N_5205);
or U6509 (N_6509,N_5805,N_5264);
or U6510 (N_6510,N_5616,N_5582);
and U6511 (N_6511,N_5561,N_5200);
and U6512 (N_6512,N_5963,N_5645);
or U6513 (N_6513,N_5027,N_5114);
and U6514 (N_6514,N_5375,N_5539);
or U6515 (N_6515,N_5664,N_5351);
or U6516 (N_6516,N_5811,N_5307);
nand U6517 (N_6517,N_5049,N_5895);
or U6518 (N_6518,N_5567,N_5756);
or U6519 (N_6519,N_5658,N_5271);
xor U6520 (N_6520,N_5360,N_5514);
nor U6521 (N_6521,N_5249,N_5900);
nor U6522 (N_6522,N_5348,N_5799);
and U6523 (N_6523,N_5313,N_5906);
nand U6524 (N_6524,N_5894,N_5071);
and U6525 (N_6525,N_5012,N_5766);
nand U6526 (N_6526,N_5370,N_5242);
nor U6527 (N_6527,N_5887,N_5747);
nor U6528 (N_6528,N_5156,N_5441);
xor U6529 (N_6529,N_5919,N_5222);
nand U6530 (N_6530,N_5777,N_5084);
nand U6531 (N_6531,N_5916,N_5984);
or U6532 (N_6532,N_5478,N_5025);
nand U6533 (N_6533,N_5973,N_5516);
or U6534 (N_6534,N_5669,N_5401);
nor U6535 (N_6535,N_5548,N_5460);
nand U6536 (N_6536,N_5486,N_5409);
and U6537 (N_6537,N_5710,N_5245);
or U6538 (N_6538,N_5808,N_5993);
nor U6539 (N_6539,N_5571,N_5118);
nand U6540 (N_6540,N_5554,N_5991);
nor U6541 (N_6541,N_5848,N_5258);
nand U6542 (N_6542,N_5505,N_5295);
or U6543 (N_6543,N_5207,N_5068);
nand U6544 (N_6544,N_5723,N_5466);
nand U6545 (N_6545,N_5674,N_5760);
nor U6546 (N_6546,N_5081,N_5834);
or U6547 (N_6547,N_5983,N_5727);
xnor U6548 (N_6548,N_5401,N_5698);
nand U6549 (N_6549,N_5203,N_5778);
nor U6550 (N_6550,N_5225,N_5228);
xor U6551 (N_6551,N_5967,N_5152);
xor U6552 (N_6552,N_5374,N_5751);
xor U6553 (N_6553,N_5818,N_5213);
nand U6554 (N_6554,N_5817,N_5362);
or U6555 (N_6555,N_5700,N_5612);
xnor U6556 (N_6556,N_5534,N_5401);
or U6557 (N_6557,N_5970,N_5567);
nand U6558 (N_6558,N_5698,N_5306);
nor U6559 (N_6559,N_5387,N_5025);
nor U6560 (N_6560,N_5433,N_5704);
xnor U6561 (N_6561,N_5165,N_5024);
nor U6562 (N_6562,N_5339,N_5604);
nor U6563 (N_6563,N_5522,N_5176);
xnor U6564 (N_6564,N_5788,N_5742);
and U6565 (N_6565,N_5126,N_5329);
nand U6566 (N_6566,N_5786,N_5556);
or U6567 (N_6567,N_5633,N_5042);
nor U6568 (N_6568,N_5993,N_5859);
or U6569 (N_6569,N_5958,N_5561);
xnor U6570 (N_6570,N_5295,N_5714);
nand U6571 (N_6571,N_5444,N_5393);
nand U6572 (N_6572,N_5585,N_5985);
and U6573 (N_6573,N_5924,N_5081);
nand U6574 (N_6574,N_5752,N_5835);
or U6575 (N_6575,N_5103,N_5925);
or U6576 (N_6576,N_5344,N_5516);
and U6577 (N_6577,N_5476,N_5817);
and U6578 (N_6578,N_5511,N_5637);
nand U6579 (N_6579,N_5610,N_5576);
nor U6580 (N_6580,N_5550,N_5640);
and U6581 (N_6581,N_5524,N_5039);
and U6582 (N_6582,N_5591,N_5476);
nor U6583 (N_6583,N_5717,N_5501);
nand U6584 (N_6584,N_5512,N_5278);
or U6585 (N_6585,N_5843,N_5022);
and U6586 (N_6586,N_5660,N_5255);
nand U6587 (N_6587,N_5193,N_5240);
or U6588 (N_6588,N_5285,N_5702);
xor U6589 (N_6589,N_5964,N_5158);
nand U6590 (N_6590,N_5873,N_5626);
and U6591 (N_6591,N_5062,N_5536);
nand U6592 (N_6592,N_5447,N_5529);
and U6593 (N_6593,N_5525,N_5933);
or U6594 (N_6594,N_5160,N_5462);
and U6595 (N_6595,N_5283,N_5936);
nand U6596 (N_6596,N_5997,N_5096);
nor U6597 (N_6597,N_5816,N_5038);
nor U6598 (N_6598,N_5203,N_5775);
or U6599 (N_6599,N_5775,N_5473);
and U6600 (N_6600,N_5490,N_5174);
nand U6601 (N_6601,N_5954,N_5304);
or U6602 (N_6602,N_5394,N_5757);
xor U6603 (N_6603,N_5702,N_5108);
nor U6604 (N_6604,N_5362,N_5176);
nand U6605 (N_6605,N_5631,N_5397);
or U6606 (N_6606,N_5738,N_5046);
or U6607 (N_6607,N_5726,N_5903);
or U6608 (N_6608,N_5018,N_5482);
and U6609 (N_6609,N_5038,N_5993);
and U6610 (N_6610,N_5201,N_5996);
nor U6611 (N_6611,N_5659,N_5620);
and U6612 (N_6612,N_5074,N_5214);
or U6613 (N_6613,N_5078,N_5650);
and U6614 (N_6614,N_5474,N_5063);
nand U6615 (N_6615,N_5609,N_5242);
nand U6616 (N_6616,N_5275,N_5018);
nand U6617 (N_6617,N_5608,N_5951);
nand U6618 (N_6618,N_5552,N_5551);
nor U6619 (N_6619,N_5157,N_5724);
and U6620 (N_6620,N_5489,N_5108);
and U6621 (N_6621,N_5821,N_5672);
nor U6622 (N_6622,N_5053,N_5778);
and U6623 (N_6623,N_5880,N_5060);
or U6624 (N_6624,N_5134,N_5385);
or U6625 (N_6625,N_5624,N_5833);
nand U6626 (N_6626,N_5844,N_5316);
nand U6627 (N_6627,N_5504,N_5933);
or U6628 (N_6628,N_5868,N_5641);
or U6629 (N_6629,N_5364,N_5095);
xor U6630 (N_6630,N_5778,N_5932);
nand U6631 (N_6631,N_5135,N_5464);
nand U6632 (N_6632,N_5322,N_5369);
nor U6633 (N_6633,N_5869,N_5691);
or U6634 (N_6634,N_5774,N_5217);
or U6635 (N_6635,N_5424,N_5717);
xor U6636 (N_6636,N_5866,N_5211);
or U6637 (N_6637,N_5784,N_5158);
and U6638 (N_6638,N_5352,N_5983);
and U6639 (N_6639,N_5538,N_5143);
nor U6640 (N_6640,N_5058,N_5590);
or U6641 (N_6641,N_5252,N_5032);
and U6642 (N_6642,N_5089,N_5339);
nand U6643 (N_6643,N_5491,N_5008);
and U6644 (N_6644,N_5428,N_5743);
and U6645 (N_6645,N_5907,N_5024);
nand U6646 (N_6646,N_5942,N_5238);
nor U6647 (N_6647,N_5352,N_5936);
or U6648 (N_6648,N_5997,N_5726);
or U6649 (N_6649,N_5187,N_5858);
xor U6650 (N_6650,N_5653,N_5637);
nor U6651 (N_6651,N_5224,N_5821);
or U6652 (N_6652,N_5152,N_5159);
and U6653 (N_6653,N_5639,N_5412);
and U6654 (N_6654,N_5760,N_5949);
nand U6655 (N_6655,N_5807,N_5161);
and U6656 (N_6656,N_5531,N_5564);
or U6657 (N_6657,N_5716,N_5446);
nor U6658 (N_6658,N_5740,N_5441);
nor U6659 (N_6659,N_5105,N_5921);
or U6660 (N_6660,N_5498,N_5723);
or U6661 (N_6661,N_5309,N_5738);
nor U6662 (N_6662,N_5197,N_5607);
and U6663 (N_6663,N_5883,N_5144);
nor U6664 (N_6664,N_5088,N_5883);
or U6665 (N_6665,N_5372,N_5632);
nor U6666 (N_6666,N_5616,N_5924);
nand U6667 (N_6667,N_5212,N_5048);
nand U6668 (N_6668,N_5146,N_5911);
nand U6669 (N_6669,N_5399,N_5876);
and U6670 (N_6670,N_5993,N_5719);
nor U6671 (N_6671,N_5106,N_5575);
nor U6672 (N_6672,N_5492,N_5789);
nand U6673 (N_6673,N_5969,N_5250);
nor U6674 (N_6674,N_5565,N_5064);
and U6675 (N_6675,N_5881,N_5604);
nor U6676 (N_6676,N_5494,N_5756);
and U6677 (N_6677,N_5542,N_5028);
nand U6678 (N_6678,N_5723,N_5107);
nor U6679 (N_6679,N_5019,N_5636);
nand U6680 (N_6680,N_5157,N_5431);
or U6681 (N_6681,N_5185,N_5662);
xor U6682 (N_6682,N_5665,N_5017);
and U6683 (N_6683,N_5406,N_5369);
and U6684 (N_6684,N_5153,N_5967);
nor U6685 (N_6685,N_5185,N_5049);
and U6686 (N_6686,N_5057,N_5616);
nand U6687 (N_6687,N_5713,N_5351);
xor U6688 (N_6688,N_5198,N_5075);
and U6689 (N_6689,N_5738,N_5205);
nor U6690 (N_6690,N_5224,N_5566);
nand U6691 (N_6691,N_5633,N_5761);
nand U6692 (N_6692,N_5994,N_5136);
nor U6693 (N_6693,N_5671,N_5305);
xnor U6694 (N_6694,N_5194,N_5163);
or U6695 (N_6695,N_5197,N_5072);
and U6696 (N_6696,N_5276,N_5142);
xnor U6697 (N_6697,N_5742,N_5975);
nand U6698 (N_6698,N_5683,N_5681);
nand U6699 (N_6699,N_5596,N_5740);
and U6700 (N_6700,N_5904,N_5992);
nand U6701 (N_6701,N_5182,N_5531);
or U6702 (N_6702,N_5804,N_5085);
nand U6703 (N_6703,N_5206,N_5784);
xnor U6704 (N_6704,N_5022,N_5786);
nor U6705 (N_6705,N_5816,N_5114);
or U6706 (N_6706,N_5554,N_5240);
nand U6707 (N_6707,N_5128,N_5966);
nor U6708 (N_6708,N_5034,N_5663);
or U6709 (N_6709,N_5398,N_5682);
xor U6710 (N_6710,N_5376,N_5621);
and U6711 (N_6711,N_5689,N_5370);
xnor U6712 (N_6712,N_5901,N_5540);
and U6713 (N_6713,N_5849,N_5716);
xnor U6714 (N_6714,N_5105,N_5897);
nor U6715 (N_6715,N_5462,N_5020);
xnor U6716 (N_6716,N_5926,N_5140);
or U6717 (N_6717,N_5586,N_5575);
nor U6718 (N_6718,N_5342,N_5315);
nand U6719 (N_6719,N_5371,N_5205);
nand U6720 (N_6720,N_5374,N_5881);
and U6721 (N_6721,N_5607,N_5286);
and U6722 (N_6722,N_5182,N_5423);
nand U6723 (N_6723,N_5786,N_5819);
xnor U6724 (N_6724,N_5821,N_5774);
or U6725 (N_6725,N_5546,N_5014);
or U6726 (N_6726,N_5405,N_5440);
nand U6727 (N_6727,N_5747,N_5142);
and U6728 (N_6728,N_5823,N_5460);
xnor U6729 (N_6729,N_5525,N_5977);
or U6730 (N_6730,N_5602,N_5446);
nand U6731 (N_6731,N_5031,N_5918);
and U6732 (N_6732,N_5692,N_5082);
nor U6733 (N_6733,N_5245,N_5363);
nand U6734 (N_6734,N_5210,N_5035);
or U6735 (N_6735,N_5686,N_5572);
and U6736 (N_6736,N_5721,N_5039);
and U6737 (N_6737,N_5651,N_5425);
and U6738 (N_6738,N_5072,N_5152);
or U6739 (N_6739,N_5350,N_5476);
nor U6740 (N_6740,N_5462,N_5365);
and U6741 (N_6741,N_5626,N_5455);
nor U6742 (N_6742,N_5971,N_5771);
or U6743 (N_6743,N_5718,N_5655);
and U6744 (N_6744,N_5911,N_5999);
nand U6745 (N_6745,N_5356,N_5870);
or U6746 (N_6746,N_5479,N_5870);
nand U6747 (N_6747,N_5140,N_5321);
nand U6748 (N_6748,N_5952,N_5145);
nor U6749 (N_6749,N_5971,N_5353);
or U6750 (N_6750,N_5195,N_5401);
or U6751 (N_6751,N_5726,N_5277);
nand U6752 (N_6752,N_5649,N_5588);
nand U6753 (N_6753,N_5557,N_5610);
nor U6754 (N_6754,N_5735,N_5769);
or U6755 (N_6755,N_5873,N_5795);
and U6756 (N_6756,N_5565,N_5305);
or U6757 (N_6757,N_5422,N_5697);
nor U6758 (N_6758,N_5482,N_5067);
nand U6759 (N_6759,N_5870,N_5168);
nand U6760 (N_6760,N_5996,N_5336);
and U6761 (N_6761,N_5985,N_5827);
nor U6762 (N_6762,N_5012,N_5108);
nor U6763 (N_6763,N_5832,N_5164);
xnor U6764 (N_6764,N_5773,N_5753);
nor U6765 (N_6765,N_5867,N_5184);
xnor U6766 (N_6766,N_5318,N_5437);
xor U6767 (N_6767,N_5041,N_5577);
or U6768 (N_6768,N_5638,N_5397);
nand U6769 (N_6769,N_5106,N_5655);
and U6770 (N_6770,N_5001,N_5968);
and U6771 (N_6771,N_5184,N_5387);
nor U6772 (N_6772,N_5978,N_5067);
and U6773 (N_6773,N_5772,N_5036);
or U6774 (N_6774,N_5690,N_5395);
xor U6775 (N_6775,N_5989,N_5677);
or U6776 (N_6776,N_5679,N_5016);
nand U6777 (N_6777,N_5228,N_5687);
and U6778 (N_6778,N_5424,N_5621);
nor U6779 (N_6779,N_5093,N_5868);
nand U6780 (N_6780,N_5014,N_5656);
xor U6781 (N_6781,N_5218,N_5754);
nor U6782 (N_6782,N_5649,N_5604);
nor U6783 (N_6783,N_5127,N_5158);
nand U6784 (N_6784,N_5228,N_5940);
nor U6785 (N_6785,N_5252,N_5191);
and U6786 (N_6786,N_5145,N_5622);
xor U6787 (N_6787,N_5818,N_5575);
nand U6788 (N_6788,N_5866,N_5579);
nand U6789 (N_6789,N_5274,N_5680);
nand U6790 (N_6790,N_5987,N_5310);
or U6791 (N_6791,N_5984,N_5507);
nor U6792 (N_6792,N_5413,N_5847);
nand U6793 (N_6793,N_5952,N_5678);
nand U6794 (N_6794,N_5851,N_5360);
xor U6795 (N_6795,N_5093,N_5998);
and U6796 (N_6796,N_5922,N_5134);
or U6797 (N_6797,N_5997,N_5642);
nor U6798 (N_6798,N_5734,N_5270);
or U6799 (N_6799,N_5052,N_5659);
and U6800 (N_6800,N_5931,N_5030);
xnor U6801 (N_6801,N_5690,N_5484);
nand U6802 (N_6802,N_5991,N_5999);
nor U6803 (N_6803,N_5204,N_5864);
xnor U6804 (N_6804,N_5173,N_5381);
or U6805 (N_6805,N_5873,N_5416);
nor U6806 (N_6806,N_5732,N_5653);
nor U6807 (N_6807,N_5852,N_5547);
or U6808 (N_6808,N_5464,N_5772);
or U6809 (N_6809,N_5877,N_5783);
nor U6810 (N_6810,N_5065,N_5079);
or U6811 (N_6811,N_5013,N_5469);
nor U6812 (N_6812,N_5987,N_5565);
nor U6813 (N_6813,N_5802,N_5705);
or U6814 (N_6814,N_5122,N_5102);
nor U6815 (N_6815,N_5410,N_5392);
or U6816 (N_6816,N_5185,N_5507);
or U6817 (N_6817,N_5451,N_5378);
and U6818 (N_6818,N_5736,N_5466);
or U6819 (N_6819,N_5242,N_5633);
nand U6820 (N_6820,N_5296,N_5538);
nor U6821 (N_6821,N_5850,N_5163);
nor U6822 (N_6822,N_5604,N_5152);
nand U6823 (N_6823,N_5104,N_5714);
nor U6824 (N_6824,N_5893,N_5567);
or U6825 (N_6825,N_5414,N_5097);
and U6826 (N_6826,N_5694,N_5438);
and U6827 (N_6827,N_5294,N_5568);
or U6828 (N_6828,N_5047,N_5055);
and U6829 (N_6829,N_5824,N_5011);
nand U6830 (N_6830,N_5509,N_5019);
xor U6831 (N_6831,N_5247,N_5913);
or U6832 (N_6832,N_5407,N_5344);
nand U6833 (N_6833,N_5973,N_5641);
nand U6834 (N_6834,N_5273,N_5480);
or U6835 (N_6835,N_5604,N_5911);
nand U6836 (N_6836,N_5911,N_5924);
or U6837 (N_6837,N_5638,N_5403);
or U6838 (N_6838,N_5351,N_5233);
and U6839 (N_6839,N_5196,N_5892);
xor U6840 (N_6840,N_5865,N_5738);
and U6841 (N_6841,N_5139,N_5256);
nor U6842 (N_6842,N_5283,N_5313);
or U6843 (N_6843,N_5420,N_5057);
nor U6844 (N_6844,N_5938,N_5415);
xor U6845 (N_6845,N_5167,N_5629);
and U6846 (N_6846,N_5226,N_5230);
nand U6847 (N_6847,N_5871,N_5507);
and U6848 (N_6848,N_5652,N_5360);
or U6849 (N_6849,N_5100,N_5015);
or U6850 (N_6850,N_5905,N_5293);
or U6851 (N_6851,N_5026,N_5086);
or U6852 (N_6852,N_5256,N_5376);
or U6853 (N_6853,N_5953,N_5109);
or U6854 (N_6854,N_5116,N_5231);
nand U6855 (N_6855,N_5185,N_5945);
nand U6856 (N_6856,N_5878,N_5959);
nor U6857 (N_6857,N_5809,N_5860);
nor U6858 (N_6858,N_5610,N_5771);
or U6859 (N_6859,N_5743,N_5293);
nand U6860 (N_6860,N_5600,N_5164);
and U6861 (N_6861,N_5807,N_5788);
and U6862 (N_6862,N_5909,N_5348);
xor U6863 (N_6863,N_5971,N_5829);
xor U6864 (N_6864,N_5736,N_5338);
or U6865 (N_6865,N_5119,N_5985);
and U6866 (N_6866,N_5316,N_5901);
xnor U6867 (N_6867,N_5574,N_5095);
or U6868 (N_6868,N_5866,N_5147);
or U6869 (N_6869,N_5815,N_5446);
nand U6870 (N_6870,N_5794,N_5792);
nor U6871 (N_6871,N_5320,N_5363);
xor U6872 (N_6872,N_5731,N_5704);
and U6873 (N_6873,N_5169,N_5894);
nor U6874 (N_6874,N_5313,N_5737);
nor U6875 (N_6875,N_5019,N_5167);
and U6876 (N_6876,N_5478,N_5524);
and U6877 (N_6877,N_5035,N_5291);
and U6878 (N_6878,N_5619,N_5890);
nor U6879 (N_6879,N_5896,N_5396);
and U6880 (N_6880,N_5838,N_5285);
nor U6881 (N_6881,N_5139,N_5668);
xnor U6882 (N_6882,N_5653,N_5663);
nor U6883 (N_6883,N_5331,N_5784);
nor U6884 (N_6884,N_5601,N_5095);
and U6885 (N_6885,N_5728,N_5048);
and U6886 (N_6886,N_5173,N_5883);
nand U6887 (N_6887,N_5377,N_5642);
nor U6888 (N_6888,N_5648,N_5676);
and U6889 (N_6889,N_5002,N_5082);
and U6890 (N_6890,N_5843,N_5485);
nor U6891 (N_6891,N_5027,N_5906);
nor U6892 (N_6892,N_5028,N_5221);
nor U6893 (N_6893,N_5323,N_5872);
or U6894 (N_6894,N_5715,N_5059);
nor U6895 (N_6895,N_5238,N_5843);
or U6896 (N_6896,N_5662,N_5467);
nand U6897 (N_6897,N_5940,N_5292);
and U6898 (N_6898,N_5480,N_5184);
nand U6899 (N_6899,N_5009,N_5884);
or U6900 (N_6900,N_5953,N_5780);
nand U6901 (N_6901,N_5041,N_5937);
nand U6902 (N_6902,N_5303,N_5173);
and U6903 (N_6903,N_5612,N_5065);
nand U6904 (N_6904,N_5895,N_5504);
or U6905 (N_6905,N_5426,N_5457);
and U6906 (N_6906,N_5054,N_5589);
xor U6907 (N_6907,N_5713,N_5416);
and U6908 (N_6908,N_5488,N_5078);
nand U6909 (N_6909,N_5688,N_5733);
or U6910 (N_6910,N_5636,N_5632);
xor U6911 (N_6911,N_5148,N_5609);
and U6912 (N_6912,N_5071,N_5858);
and U6913 (N_6913,N_5261,N_5942);
nor U6914 (N_6914,N_5010,N_5861);
nand U6915 (N_6915,N_5207,N_5415);
nor U6916 (N_6916,N_5707,N_5050);
and U6917 (N_6917,N_5335,N_5843);
or U6918 (N_6918,N_5706,N_5739);
nand U6919 (N_6919,N_5738,N_5919);
nand U6920 (N_6920,N_5141,N_5204);
or U6921 (N_6921,N_5271,N_5519);
nor U6922 (N_6922,N_5967,N_5156);
nand U6923 (N_6923,N_5017,N_5061);
nand U6924 (N_6924,N_5874,N_5047);
nor U6925 (N_6925,N_5084,N_5797);
or U6926 (N_6926,N_5514,N_5201);
and U6927 (N_6927,N_5425,N_5900);
nor U6928 (N_6928,N_5797,N_5689);
nand U6929 (N_6929,N_5588,N_5800);
or U6930 (N_6930,N_5959,N_5904);
nor U6931 (N_6931,N_5957,N_5820);
nand U6932 (N_6932,N_5082,N_5577);
nor U6933 (N_6933,N_5407,N_5897);
nor U6934 (N_6934,N_5562,N_5230);
nor U6935 (N_6935,N_5711,N_5963);
and U6936 (N_6936,N_5857,N_5789);
or U6937 (N_6937,N_5671,N_5280);
or U6938 (N_6938,N_5807,N_5418);
nand U6939 (N_6939,N_5239,N_5637);
nand U6940 (N_6940,N_5094,N_5242);
and U6941 (N_6941,N_5613,N_5427);
nand U6942 (N_6942,N_5556,N_5512);
or U6943 (N_6943,N_5587,N_5637);
or U6944 (N_6944,N_5672,N_5081);
xor U6945 (N_6945,N_5032,N_5021);
and U6946 (N_6946,N_5401,N_5607);
nor U6947 (N_6947,N_5968,N_5555);
xor U6948 (N_6948,N_5759,N_5597);
nand U6949 (N_6949,N_5419,N_5252);
or U6950 (N_6950,N_5226,N_5583);
or U6951 (N_6951,N_5937,N_5734);
nor U6952 (N_6952,N_5126,N_5841);
xor U6953 (N_6953,N_5488,N_5184);
or U6954 (N_6954,N_5383,N_5186);
nor U6955 (N_6955,N_5568,N_5864);
nor U6956 (N_6956,N_5763,N_5209);
xor U6957 (N_6957,N_5436,N_5494);
nor U6958 (N_6958,N_5558,N_5522);
nor U6959 (N_6959,N_5622,N_5244);
and U6960 (N_6960,N_5803,N_5608);
nand U6961 (N_6961,N_5083,N_5121);
or U6962 (N_6962,N_5209,N_5520);
or U6963 (N_6963,N_5209,N_5369);
nor U6964 (N_6964,N_5396,N_5600);
or U6965 (N_6965,N_5526,N_5511);
and U6966 (N_6966,N_5310,N_5554);
or U6967 (N_6967,N_5664,N_5844);
xnor U6968 (N_6968,N_5158,N_5590);
and U6969 (N_6969,N_5459,N_5124);
nor U6970 (N_6970,N_5718,N_5547);
nor U6971 (N_6971,N_5955,N_5907);
nand U6972 (N_6972,N_5126,N_5550);
nand U6973 (N_6973,N_5364,N_5424);
or U6974 (N_6974,N_5617,N_5776);
nand U6975 (N_6975,N_5869,N_5408);
nand U6976 (N_6976,N_5020,N_5904);
or U6977 (N_6977,N_5684,N_5163);
or U6978 (N_6978,N_5704,N_5687);
nand U6979 (N_6979,N_5300,N_5265);
or U6980 (N_6980,N_5329,N_5438);
nand U6981 (N_6981,N_5041,N_5273);
or U6982 (N_6982,N_5151,N_5672);
xor U6983 (N_6983,N_5981,N_5881);
nor U6984 (N_6984,N_5047,N_5570);
and U6985 (N_6985,N_5694,N_5277);
and U6986 (N_6986,N_5686,N_5701);
nor U6987 (N_6987,N_5769,N_5215);
nor U6988 (N_6988,N_5314,N_5590);
and U6989 (N_6989,N_5504,N_5202);
nor U6990 (N_6990,N_5451,N_5694);
nor U6991 (N_6991,N_5572,N_5368);
xor U6992 (N_6992,N_5498,N_5629);
nand U6993 (N_6993,N_5822,N_5118);
or U6994 (N_6994,N_5327,N_5278);
and U6995 (N_6995,N_5608,N_5671);
or U6996 (N_6996,N_5408,N_5041);
nor U6997 (N_6997,N_5009,N_5915);
nand U6998 (N_6998,N_5629,N_5067);
and U6999 (N_6999,N_5950,N_5414);
xnor U7000 (N_7000,N_6184,N_6359);
nand U7001 (N_7001,N_6876,N_6998);
or U7002 (N_7002,N_6809,N_6954);
nor U7003 (N_7003,N_6315,N_6860);
or U7004 (N_7004,N_6419,N_6991);
nand U7005 (N_7005,N_6476,N_6721);
nor U7006 (N_7006,N_6239,N_6942);
nand U7007 (N_7007,N_6678,N_6278);
xor U7008 (N_7008,N_6081,N_6387);
nor U7009 (N_7009,N_6852,N_6715);
or U7010 (N_7010,N_6693,N_6139);
nor U7011 (N_7011,N_6204,N_6245);
or U7012 (N_7012,N_6968,N_6875);
and U7013 (N_7013,N_6085,N_6172);
xor U7014 (N_7014,N_6485,N_6066);
or U7015 (N_7015,N_6530,N_6189);
nor U7016 (N_7016,N_6163,N_6389);
nand U7017 (N_7017,N_6486,N_6620);
xnor U7018 (N_7018,N_6347,N_6123);
or U7019 (N_7019,N_6258,N_6298);
nand U7020 (N_7020,N_6576,N_6345);
nand U7021 (N_7021,N_6899,N_6031);
or U7022 (N_7022,N_6124,N_6197);
and U7023 (N_7023,N_6279,N_6846);
nand U7024 (N_7024,N_6282,N_6767);
and U7025 (N_7025,N_6810,N_6736);
or U7026 (N_7026,N_6836,N_6540);
or U7027 (N_7027,N_6341,N_6803);
and U7028 (N_7028,N_6548,N_6330);
and U7029 (N_7029,N_6076,N_6395);
or U7030 (N_7030,N_6270,N_6946);
and U7031 (N_7031,N_6498,N_6331);
nand U7032 (N_7032,N_6499,N_6006);
nor U7033 (N_7033,N_6152,N_6661);
and U7034 (N_7034,N_6324,N_6391);
nand U7035 (N_7035,N_6786,N_6764);
or U7036 (N_7036,N_6554,N_6658);
and U7037 (N_7037,N_6884,N_6725);
nand U7038 (N_7038,N_6089,N_6606);
nor U7039 (N_7039,N_6779,N_6717);
xnor U7040 (N_7040,N_6585,N_6597);
nor U7041 (N_7041,N_6343,N_6862);
nor U7042 (N_7042,N_6325,N_6513);
or U7043 (N_7043,N_6101,N_6667);
nand U7044 (N_7044,N_6837,N_6003);
or U7045 (N_7045,N_6580,N_6980);
nand U7046 (N_7046,N_6417,N_6794);
or U7047 (N_7047,N_6571,N_6115);
nor U7048 (N_7048,N_6007,N_6989);
or U7049 (N_7049,N_6246,N_6569);
nand U7050 (N_7050,N_6255,N_6562);
nor U7051 (N_7051,N_6553,N_6136);
nor U7052 (N_7052,N_6542,N_6782);
nor U7053 (N_7053,N_6493,N_6844);
and U7054 (N_7054,N_6581,N_6900);
nor U7055 (N_7055,N_6393,N_6097);
nand U7056 (N_7056,N_6484,N_6156);
or U7057 (N_7057,N_6262,N_6240);
nor U7058 (N_7058,N_6549,N_6543);
nand U7059 (N_7059,N_6538,N_6168);
nor U7060 (N_7060,N_6413,N_6170);
or U7061 (N_7061,N_6222,N_6425);
nand U7062 (N_7062,N_6774,N_6941);
and U7063 (N_7063,N_6473,N_6853);
or U7064 (N_7064,N_6212,N_6028);
nand U7065 (N_7065,N_6988,N_6171);
or U7066 (N_7066,N_6025,N_6877);
or U7067 (N_7067,N_6679,N_6149);
nor U7068 (N_7068,N_6924,N_6649);
and U7069 (N_7069,N_6456,N_6971);
xnor U7070 (N_7070,N_6444,N_6688);
nor U7071 (N_7071,N_6645,N_6958);
or U7072 (N_7072,N_6348,N_6407);
or U7073 (N_7073,N_6630,N_6592);
and U7074 (N_7074,N_6314,N_6800);
nor U7075 (N_7075,N_6607,N_6323);
and U7076 (N_7076,N_6272,N_6362);
or U7077 (N_7077,N_6823,N_6832);
and U7078 (N_7078,N_6052,N_6372);
and U7079 (N_7079,N_6628,N_6472);
nand U7080 (N_7080,N_6510,N_6833);
or U7081 (N_7081,N_6882,N_6889);
or U7082 (N_7082,N_6281,N_6340);
nand U7083 (N_7083,N_6728,N_6627);
nor U7084 (N_7084,N_6927,N_6121);
nor U7085 (N_7085,N_6509,N_6237);
and U7086 (N_7086,N_6730,N_6408);
xor U7087 (N_7087,N_6365,N_6586);
nor U7088 (N_7088,N_6894,N_6455);
or U7089 (N_7089,N_6026,N_6870);
and U7090 (N_7090,N_6429,N_6888);
nor U7091 (N_7091,N_6344,N_6880);
nor U7092 (N_7092,N_6225,N_6634);
xnor U7093 (N_7093,N_6221,N_6826);
and U7094 (N_7094,N_6394,N_6653);
and U7095 (N_7095,N_6093,N_6249);
nor U7096 (N_7096,N_6854,N_6609);
and U7097 (N_7097,N_6415,N_6175);
nand U7098 (N_7098,N_6652,N_6605);
nor U7099 (N_7099,N_6783,N_6944);
nor U7100 (N_7100,N_6896,N_6082);
or U7101 (N_7101,N_6707,N_6705);
or U7102 (N_7102,N_6883,N_6985);
nor U7103 (N_7103,N_6271,N_6040);
or U7104 (N_7104,N_6914,N_6874);
or U7105 (N_7105,N_6088,N_6032);
nand U7106 (N_7106,N_6179,N_6771);
and U7107 (N_7107,N_6412,N_6447);
nor U7108 (N_7108,N_6441,N_6719);
nand U7109 (N_7109,N_6952,N_6073);
nand U7110 (N_7110,N_6435,N_6500);
or U7111 (N_7111,N_6062,N_6937);
and U7112 (N_7112,N_6740,N_6213);
nand U7113 (N_7113,N_6935,N_6129);
and U7114 (N_7114,N_6648,N_6778);
nor U7115 (N_7115,N_6898,N_6697);
xor U7116 (N_7116,N_6892,N_6147);
nand U7117 (N_7117,N_6828,N_6915);
and U7118 (N_7118,N_6113,N_6694);
and U7119 (N_7119,N_6600,N_6296);
nand U7120 (N_7120,N_6611,N_6403);
nor U7121 (N_7121,N_6573,N_6247);
and U7122 (N_7122,N_6064,N_6722);
nand U7123 (N_7123,N_6893,N_6077);
xor U7124 (N_7124,N_6005,N_6502);
xnor U7125 (N_7125,N_6838,N_6020);
nand U7126 (N_7126,N_6729,N_6636);
nor U7127 (N_7127,N_6598,N_6938);
nand U7128 (N_7128,N_6680,N_6069);
or U7129 (N_7129,N_6329,N_6057);
xnor U7130 (N_7130,N_6406,N_6478);
or U7131 (N_7131,N_6690,N_6112);
and U7132 (N_7132,N_6030,N_6370);
or U7133 (N_7133,N_6462,N_6303);
or U7134 (N_7134,N_6201,N_6483);
and U7135 (N_7135,N_6831,N_6046);
or U7136 (N_7136,N_6651,N_6067);
xnor U7137 (N_7137,N_6735,N_6326);
or U7138 (N_7138,N_6834,N_6792);
nor U7139 (N_7139,N_6858,N_6308);
nor U7140 (N_7140,N_6199,N_6922);
and U7141 (N_7141,N_6550,N_6866);
or U7142 (N_7142,N_6961,N_6770);
nand U7143 (N_7143,N_6511,N_6855);
or U7144 (N_7144,N_6777,N_6228);
nor U7145 (N_7145,N_6100,N_6364);
nand U7146 (N_7146,N_6471,N_6529);
xnor U7147 (N_7147,N_6632,N_6912);
nor U7148 (N_7148,N_6733,N_6891);
and U7149 (N_7149,N_6805,N_6675);
nand U7150 (N_7150,N_6063,N_6321);
nor U7151 (N_7151,N_6037,N_6144);
nand U7152 (N_7152,N_6781,N_6928);
nor U7153 (N_7153,N_6098,N_6078);
nand U7154 (N_7154,N_6790,N_6458);
nand U7155 (N_7155,N_6134,N_6383);
nor U7156 (N_7156,N_6254,N_6619);
or U7157 (N_7157,N_6993,N_6428);
nand U7158 (N_7158,N_6293,N_6290);
and U7159 (N_7159,N_6738,N_6399);
nor U7160 (N_7160,N_6351,N_6061);
and U7161 (N_7161,N_6582,N_6566);
and U7162 (N_7162,N_6801,N_6772);
and U7163 (N_7163,N_6984,N_6754);
xor U7164 (N_7164,N_6501,N_6557);
and U7165 (N_7165,N_6038,N_6295);
and U7166 (N_7166,N_6635,N_6186);
and U7167 (N_7167,N_6518,N_6737);
or U7168 (N_7168,N_6034,N_6158);
nor U7169 (N_7169,N_6018,N_6533);
or U7170 (N_7170,N_6842,N_6224);
xor U7171 (N_7171,N_6319,N_6327);
xor U7172 (N_7172,N_6027,N_6107);
nor U7173 (N_7173,N_6521,N_6773);
nand U7174 (N_7174,N_6440,N_6130);
xor U7175 (N_7175,N_6350,N_6301);
and U7176 (N_7176,N_6559,N_6263);
nor U7177 (N_7177,N_6102,N_6616);
and U7178 (N_7178,N_6741,N_6925);
nor U7179 (N_7179,N_6074,N_6957);
and U7180 (N_7180,N_6438,N_6167);
nor U7181 (N_7181,N_6071,N_6223);
nand U7182 (N_7182,N_6033,N_6241);
or U7183 (N_7183,N_6380,N_6570);
nand U7184 (N_7184,N_6516,N_6604);
nor U7185 (N_7185,N_6595,N_6904);
nand U7186 (N_7186,N_6353,N_6042);
or U7187 (N_7187,N_6475,N_6299);
and U7188 (N_7188,N_6119,N_6704);
nor U7189 (N_7189,N_6614,N_6994);
nor U7190 (N_7190,N_6219,N_6140);
or U7191 (N_7191,N_6494,N_6804);
and U7192 (N_7192,N_6227,N_6701);
nor U7193 (N_7193,N_6215,N_6662);
nand U7194 (N_7194,N_6517,N_6229);
nand U7195 (N_7195,N_6996,N_6318);
nor U7196 (N_7196,N_6808,N_6879);
nor U7197 (N_7197,N_6713,N_6474);
xor U7198 (N_7198,N_6449,N_6011);
nand U7199 (N_7199,N_6709,N_6871);
and U7200 (N_7200,N_6205,N_6748);
and U7201 (N_7201,N_6143,N_6274);
nor U7202 (N_7202,N_6931,N_6712);
nand U7203 (N_7203,N_6349,N_6235);
and U7204 (N_7204,N_6572,N_6742);
and U7205 (N_7205,N_6584,N_6336);
and U7206 (N_7206,N_6048,N_6819);
nand U7207 (N_7207,N_6257,N_6374);
nand U7208 (N_7208,N_6430,N_6014);
nor U7209 (N_7209,N_6226,N_6194);
and U7210 (N_7210,N_6234,N_6575);
nand U7211 (N_7211,N_6162,N_6747);
and U7212 (N_7212,N_6791,N_6930);
nand U7213 (N_7213,N_6962,N_6176);
and U7214 (N_7214,N_6165,N_6655);
or U7215 (N_7215,N_6676,N_6666);
nand U7216 (N_7216,N_6945,N_6285);
xnor U7217 (N_7217,N_6997,N_6090);
nor U7218 (N_7218,N_6216,N_6872);
nor U7219 (N_7219,N_6718,N_6758);
and U7220 (N_7220,N_6625,N_6811);
or U7221 (N_7221,N_6190,N_6505);
xor U7222 (N_7222,N_6587,N_6789);
and U7223 (N_7223,N_6198,N_6354);
nor U7224 (N_7224,N_6490,N_6813);
nor U7225 (N_7225,N_6467,N_6544);
or U7226 (N_7226,N_6681,N_6951);
and U7227 (N_7227,N_6388,N_6133);
and U7228 (N_7228,N_6835,N_6452);
nand U7229 (N_7229,N_6322,N_6200);
nand U7230 (N_7230,N_6659,N_6703);
nor U7231 (N_7231,N_6768,N_6016);
xnor U7232 (N_7232,N_6250,N_6141);
nor U7233 (N_7233,N_6480,N_6035);
nor U7234 (N_7234,N_6489,N_6049);
xnor U7235 (N_7235,N_6799,N_6881);
and U7236 (N_7236,N_6264,N_6563);
nand U7237 (N_7237,N_6695,N_6639);
nand U7238 (N_7238,N_6907,N_6964);
or U7239 (N_7239,N_6268,N_6137);
and U7240 (N_7240,N_6917,N_6131);
nor U7241 (N_7241,N_6337,N_6091);
nand U7242 (N_7242,N_6459,N_6045);
nor U7243 (N_7243,N_6379,N_6385);
nand U7244 (N_7244,N_6381,N_6041);
nand U7245 (N_7245,N_6677,N_6919);
xnor U7246 (N_7246,N_6432,N_6716);
or U7247 (N_7247,N_6105,N_6276);
and U7248 (N_7248,N_6373,N_6304);
nor U7249 (N_7249,N_6291,N_6650);
nor U7250 (N_7250,N_6863,N_6785);
nand U7251 (N_7251,N_6103,N_6470);
and U7252 (N_7252,N_6411,N_6055);
xor U7253 (N_7253,N_6079,N_6434);
xnor U7254 (N_7254,N_6450,N_6943);
nor U7255 (N_7255,N_6684,N_6665);
nor U7256 (N_7256,N_6457,N_6236);
and U7257 (N_7257,N_6185,N_6671);
and U7258 (N_7258,N_6206,N_6885);
xnor U7259 (N_7259,N_6092,N_6948);
or U7260 (N_7260,N_6851,N_6638);
nand U7261 (N_7261,N_6682,N_6183);
and U7262 (N_7262,N_6702,N_6940);
and U7263 (N_7263,N_6259,N_6512);
and U7264 (N_7264,N_6454,N_6699);
xnor U7265 (N_7265,N_6626,N_6547);
and U7266 (N_7266,N_6905,N_6802);
nand U7267 (N_7267,N_6536,N_6643);
or U7268 (N_7268,N_6002,N_6384);
nor U7269 (N_7269,N_6416,N_6352);
and U7270 (N_7270,N_6177,N_6292);
and U7271 (N_7271,N_6850,N_6193);
or U7272 (N_7272,N_6155,N_6277);
nand U7273 (N_7273,N_6160,N_6135);
and U7274 (N_7274,N_6132,N_6979);
or U7275 (N_7275,N_6686,N_6775);
nand U7276 (N_7276,N_6451,N_6356);
or U7277 (N_7277,N_6094,N_6685);
nor U7278 (N_7278,N_6106,N_6443);
nand U7279 (N_7279,N_6487,N_6496);
and U7280 (N_7280,N_6442,N_6065);
and U7281 (N_7281,N_6251,N_6378);
or U7282 (N_7282,N_6843,N_6567);
or U7283 (N_7283,N_6044,N_6903);
nand U7284 (N_7284,N_6873,N_6286);
or U7285 (N_7285,N_6358,N_6756);
nor U7286 (N_7286,N_6947,N_6009);
xor U7287 (N_7287,N_6418,N_6766);
or U7288 (N_7288,N_6817,N_6551);
and U7289 (N_7289,N_6939,N_6910);
nand U7290 (N_7290,N_6188,N_6845);
and U7291 (N_7291,N_6099,N_6217);
nand U7292 (N_7292,N_6956,N_6750);
nand U7293 (N_7293,N_6982,N_6692);
nand U7294 (N_7294,N_6153,N_6732);
nor U7295 (N_7295,N_6955,N_6840);
or U7296 (N_7296,N_6820,N_6829);
and U7297 (N_7297,N_6448,N_6966);
or U7298 (N_7298,N_6749,N_6392);
or U7299 (N_7299,N_6355,N_6926);
and U7300 (N_7300,N_6054,N_6793);
or U7301 (N_7301,N_6981,N_6531);
xnor U7302 (N_7302,N_6753,N_6302);
and U7303 (N_7303,N_6895,N_6402);
or U7304 (N_7304,N_6950,N_6537);
and U7305 (N_7305,N_6111,N_6477);
nor U7306 (N_7306,N_6723,N_6492);
or U7307 (N_7307,N_6488,N_6368);
nor U7308 (N_7308,N_6861,N_6466);
xnor U7309 (N_7309,N_6503,N_6528);
nand U7310 (N_7310,N_6618,N_6977);
nor U7311 (N_7311,N_6433,N_6796);
nor U7312 (N_7312,N_6109,N_6967);
nand U7313 (N_7313,N_6495,N_6633);
nand U7314 (N_7314,N_6424,N_6687);
or U7315 (N_7315,N_6288,N_6409);
xor U7316 (N_7316,N_6734,N_6560);
nor U7317 (N_7317,N_6269,N_6987);
nand U7318 (N_7318,N_6328,N_6519);
nor U7319 (N_7319,N_6960,N_6248);
and U7320 (N_7320,N_6593,N_6776);
or U7321 (N_7321,N_6689,N_6357);
nand U7322 (N_7322,N_6589,N_6959);
nor U7323 (N_7323,N_6847,N_6640);
or U7324 (N_7324,N_6398,N_6588);
or U7325 (N_7325,N_6646,N_6827);
nor U7326 (N_7326,N_6594,N_6283);
or U7327 (N_7327,N_6230,N_6624);
or U7328 (N_7328,N_6210,N_6615);
or U7329 (N_7329,N_6673,N_6744);
nand U7330 (N_7330,N_6086,N_6053);
and U7331 (N_7331,N_6859,N_6751);
xor U7332 (N_7332,N_6706,N_6514);
and U7333 (N_7333,N_6612,N_6508);
xnor U7334 (N_7334,N_6507,N_6075);
nand U7335 (N_7335,N_6672,N_6181);
nor U7336 (N_7336,N_6526,N_6669);
or U7337 (N_7337,N_6752,N_6390);
or U7338 (N_7338,N_6375,N_6642);
and U7339 (N_7339,N_6127,N_6668);
xnor U7340 (N_7340,N_6739,N_6965);
or U7341 (N_7341,N_6506,N_6126);
and U7342 (N_7342,N_6108,N_6414);
nor U7343 (N_7343,N_6869,N_6469);
nor U7344 (N_7344,N_6305,N_6504);
xor U7345 (N_7345,N_6608,N_6660);
nand U7346 (N_7346,N_6761,N_6004);
and U7347 (N_7347,N_6436,N_6759);
xor U7348 (N_7348,N_6720,N_6564);
xor U7349 (N_7349,N_6294,N_6339);
nand U7350 (N_7350,N_6267,N_6700);
nor U7351 (N_7351,N_6481,N_6024);
nor U7352 (N_7352,N_6929,N_6312);
and U7353 (N_7353,N_6050,N_6901);
nor U7354 (N_7354,N_6724,N_6934);
nand U7355 (N_7355,N_6887,N_6120);
nand U7356 (N_7356,N_6360,N_6769);
nand U7357 (N_7357,N_6203,N_6807);
and U7358 (N_7358,N_6110,N_6405);
nor U7359 (N_7359,N_6664,N_6051);
or U7360 (N_7360,N_6986,N_6856);
nor U7361 (N_7361,N_6902,N_6310);
nand U7362 (N_7362,N_6253,N_6696);
nand U7363 (N_7363,N_6555,N_6975);
xnor U7364 (N_7364,N_6599,N_6404);
and U7365 (N_7365,N_6117,N_6663);
xnor U7366 (N_7366,N_6656,N_6287);
nor U7367 (N_7367,N_6118,N_6577);
nor U7368 (N_7368,N_6070,N_6784);
or U7369 (N_7369,N_6932,N_6146);
and U7370 (N_7370,N_6397,N_6963);
nand U7371 (N_7371,N_6579,N_6261);
nor U7372 (N_7372,N_6825,N_6814);
nor U7373 (N_7373,N_6479,N_6461);
xor U7374 (N_7374,N_6252,N_6243);
and U7375 (N_7375,N_6161,N_6265);
nor U7376 (N_7376,N_6897,N_6332);
or U7377 (N_7377,N_6218,N_6333);
or U7378 (N_7378,N_6710,N_6220);
xor U7379 (N_7379,N_6148,N_6166);
and U7380 (N_7380,N_6174,N_6909);
xor U7381 (N_7381,N_6936,N_6012);
nor U7382 (N_7382,N_6953,N_6561);
nor U7383 (N_7383,N_6320,N_6008);
nand U7384 (N_7384,N_6039,N_6056);
or U7385 (N_7385,N_6596,N_6180);
nand U7386 (N_7386,N_6568,N_6795);
or U7387 (N_7387,N_6195,N_6990);
nor U7388 (N_7388,N_6464,N_6164);
nor U7389 (N_7389,N_6421,N_6232);
or U7390 (N_7390,N_6868,N_6017);
and U7391 (N_7391,N_6812,N_6995);
xor U7392 (N_7392,N_6746,N_6244);
xor U7393 (N_7393,N_6157,N_6921);
nor U7394 (N_7394,N_6545,N_6116);
and U7395 (N_7395,N_6797,N_6242);
nor U7396 (N_7396,N_6182,N_6209);
nor U7397 (N_7397,N_6439,N_6306);
or U7398 (N_7398,N_6029,N_6765);
and U7399 (N_7399,N_6266,N_6969);
nor U7400 (N_7400,N_6491,N_6151);
xor U7401 (N_7401,N_6520,N_6202);
nand U7402 (N_7402,N_6238,N_6437);
nand U7403 (N_7403,N_6371,N_6192);
and U7404 (N_7404,N_6787,N_6601);
nor U7405 (N_7405,N_6482,N_6708);
and U7406 (N_7406,N_6644,N_6886);
or U7407 (N_7407,N_6000,N_6463);
or U7408 (N_7408,N_6974,N_6552);
nor U7409 (N_7409,N_6617,N_6556);
and U7410 (N_7410,N_6015,N_6565);
nand U7411 (N_7411,N_6821,N_6857);
nor U7412 (N_7412,N_6822,N_6818);
or U7413 (N_7413,N_6023,N_6401);
or U7414 (N_7414,N_6714,N_6933);
nor U7415 (N_7415,N_6497,N_6603);
or U7416 (N_7416,N_6527,N_6431);
or U7417 (N_7417,N_6726,N_6231);
nand U7418 (N_7418,N_6317,N_6068);
and U7419 (N_7419,N_6623,N_6036);
nor U7420 (N_7420,N_6522,N_6072);
nand U7421 (N_7421,N_6260,N_6114);
or U7422 (N_7422,N_6515,N_6363);
nor U7423 (N_7423,N_6637,N_6546);
or U7424 (N_7424,N_6446,N_6711);
and U7425 (N_7425,N_6335,N_6670);
and U7426 (N_7426,N_6763,N_6154);
or U7427 (N_7427,N_6369,N_6001);
and U7428 (N_7428,N_6824,N_6890);
xor U7429 (N_7429,N_6342,N_6013);
xnor U7430 (N_7430,N_6613,N_6641);
nor U7431 (N_7431,N_6908,N_6084);
nand U7432 (N_7432,N_6420,N_6083);
and U7433 (N_7433,N_6095,N_6460);
nand U7434 (N_7434,N_6839,N_6346);
and U7435 (N_7435,N_6972,N_6830);
nor U7436 (N_7436,N_6970,N_6534);
and U7437 (N_7437,N_6558,N_6629);
or U7438 (N_7438,N_6523,N_6973);
nand U7439 (N_7439,N_6532,N_6142);
or U7440 (N_7440,N_6080,N_6465);
and U7441 (N_7441,N_6191,N_6674);
and U7442 (N_7442,N_6361,N_6920);
nor U7443 (N_7443,N_6280,N_6196);
nand U7444 (N_7444,N_6622,N_6574);
nor U7445 (N_7445,N_6426,N_6731);
and U7446 (N_7446,N_6583,N_6541);
nor U7447 (N_7447,N_6918,N_6757);
nor U7448 (N_7448,N_6976,N_6410);
nor U7449 (N_7449,N_6524,N_6590);
and U7450 (N_7450,N_6647,N_6949);
or U7451 (N_7451,N_6760,N_6683);
or U7452 (N_7452,N_6021,N_6535);
xnor U7453 (N_7453,N_6311,N_6816);
or U7454 (N_7454,N_6019,N_6762);
xnor U7455 (N_7455,N_6211,N_6864);
or U7456 (N_7456,N_6386,N_6376);
and U7457 (N_7457,N_6525,N_6104);
xnor U7458 (N_7458,N_6591,N_6841);
nand U7459 (N_7459,N_6788,N_6159);
and U7460 (N_7460,N_6128,N_6780);
xnor U7461 (N_7461,N_6422,N_6297);
xor U7462 (N_7462,N_6207,N_6289);
xor U7463 (N_7463,N_6631,N_6275);
nand U7464 (N_7464,N_6755,N_6233);
or U7465 (N_7465,N_6145,N_6906);
and U7466 (N_7466,N_6691,N_6923);
xor U7467 (N_7467,N_6468,N_6169);
nor U7468 (N_7468,N_6983,N_6913);
or U7469 (N_7469,N_6423,N_6539);
or U7470 (N_7470,N_6377,N_6125);
nor U7471 (N_7471,N_6334,N_6911);
and U7472 (N_7472,N_6743,N_6060);
and U7473 (N_7473,N_6396,N_6214);
and U7474 (N_7474,N_6043,N_6878);
nor U7475 (N_7475,N_6256,N_6745);
nor U7476 (N_7476,N_6427,N_6307);
nand U7477 (N_7477,N_6367,N_6453);
or U7478 (N_7478,N_6727,N_6122);
nand U7479 (N_7479,N_6610,N_6698);
nor U7480 (N_7480,N_6178,N_6806);
xnor U7481 (N_7481,N_6400,N_6173);
nand U7482 (N_7482,N_6445,N_6978);
xnor U7483 (N_7483,N_6058,N_6654);
nor U7484 (N_7484,N_6059,N_6187);
nand U7485 (N_7485,N_6150,N_6284);
or U7486 (N_7486,N_6047,N_6096);
xor U7487 (N_7487,N_6992,N_6382);
nor U7488 (N_7488,N_6798,N_6366);
or U7489 (N_7489,N_6087,N_6022);
nand U7490 (N_7490,N_6815,N_6999);
and U7491 (N_7491,N_6273,N_6316);
nor U7492 (N_7492,N_6138,N_6309);
nor U7493 (N_7493,N_6602,N_6313);
or U7494 (N_7494,N_6621,N_6849);
xnor U7495 (N_7495,N_6208,N_6578);
or U7496 (N_7496,N_6916,N_6848);
and U7497 (N_7497,N_6865,N_6300);
nor U7498 (N_7498,N_6867,N_6338);
nor U7499 (N_7499,N_6010,N_6657);
nand U7500 (N_7500,N_6284,N_6959);
nor U7501 (N_7501,N_6594,N_6019);
and U7502 (N_7502,N_6717,N_6944);
or U7503 (N_7503,N_6350,N_6095);
and U7504 (N_7504,N_6830,N_6956);
and U7505 (N_7505,N_6291,N_6238);
and U7506 (N_7506,N_6568,N_6021);
and U7507 (N_7507,N_6921,N_6623);
nand U7508 (N_7508,N_6992,N_6331);
nor U7509 (N_7509,N_6425,N_6288);
or U7510 (N_7510,N_6240,N_6779);
nor U7511 (N_7511,N_6418,N_6026);
and U7512 (N_7512,N_6187,N_6922);
nand U7513 (N_7513,N_6749,N_6190);
xor U7514 (N_7514,N_6797,N_6328);
nand U7515 (N_7515,N_6773,N_6441);
nand U7516 (N_7516,N_6966,N_6012);
and U7517 (N_7517,N_6058,N_6851);
nor U7518 (N_7518,N_6211,N_6217);
nor U7519 (N_7519,N_6679,N_6499);
nor U7520 (N_7520,N_6733,N_6159);
nand U7521 (N_7521,N_6527,N_6821);
xor U7522 (N_7522,N_6748,N_6184);
and U7523 (N_7523,N_6142,N_6678);
and U7524 (N_7524,N_6526,N_6662);
nor U7525 (N_7525,N_6678,N_6654);
nand U7526 (N_7526,N_6039,N_6083);
nor U7527 (N_7527,N_6120,N_6464);
nor U7528 (N_7528,N_6612,N_6384);
nor U7529 (N_7529,N_6232,N_6532);
nand U7530 (N_7530,N_6805,N_6174);
nand U7531 (N_7531,N_6037,N_6094);
nor U7532 (N_7532,N_6972,N_6579);
or U7533 (N_7533,N_6338,N_6987);
nor U7534 (N_7534,N_6740,N_6876);
nor U7535 (N_7535,N_6770,N_6838);
nand U7536 (N_7536,N_6389,N_6589);
nand U7537 (N_7537,N_6676,N_6929);
nor U7538 (N_7538,N_6711,N_6733);
nand U7539 (N_7539,N_6035,N_6791);
xnor U7540 (N_7540,N_6441,N_6955);
nand U7541 (N_7541,N_6495,N_6835);
nand U7542 (N_7542,N_6116,N_6130);
or U7543 (N_7543,N_6607,N_6415);
nand U7544 (N_7544,N_6607,N_6121);
nor U7545 (N_7545,N_6138,N_6914);
nor U7546 (N_7546,N_6118,N_6084);
xor U7547 (N_7547,N_6009,N_6216);
and U7548 (N_7548,N_6986,N_6526);
nor U7549 (N_7549,N_6551,N_6092);
nor U7550 (N_7550,N_6888,N_6029);
or U7551 (N_7551,N_6945,N_6148);
nand U7552 (N_7552,N_6834,N_6816);
and U7553 (N_7553,N_6528,N_6416);
or U7554 (N_7554,N_6713,N_6535);
nand U7555 (N_7555,N_6933,N_6561);
and U7556 (N_7556,N_6982,N_6822);
or U7557 (N_7557,N_6837,N_6271);
nand U7558 (N_7558,N_6818,N_6642);
nand U7559 (N_7559,N_6488,N_6316);
nand U7560 (N_7560,N_6354,N_6461);
nor U7561 (N_7561,N_6212,N_6378);
and U7562 (N_7562,N_6094,N_6137);
nand U7563 (N_7563,N_6066,N_6658);
xnor U7564 (N_7564,N_6856,N_6923);
or U7565 (N_7565,N_6163,N_6839);
nor U7566 (N_7566,N_6985,N_6756);
xnor U7567 (N_7567,N_6588,N_6327);
or U7568 (N_7568,N_6049,N_6231);
nor U7569 (N_7569,N_6349,N_6366);
nand U7570 (N_7570,N_6349,N_6150);
and U7571 (N_7571,N_6813,N_6189);
and U7572 (N_7572,N_6761,N_6325);
or U7573 (N_7573,N_6555,N_6964);
nand U7574 (N_7574,N_6574,N_6382);
nor U7575 (N_7575,N_6878,N_6261);
nand U7576 (N_7576,N_6267,N_6428);
and U7577 (N_7577,N_6235,N_6598);
or U7578 (N_7578,N_6843,N_6399);
nor U7579 (N_7579,N_6783,N_6269);
or U7580 (N_7580,N_6608,N_6375);
nand U7581 (N_7581,N_6750,N_6244);
nand U7582 (N_7582,N_6573,N_6774);
nor U7583 (N_7583,N_6052,N_6963);
nand U7584 (N_7584,N_6032,N_6098);
nor U7585 (N_7585,N_6338,N_6978);
nand U7586 (N_7586,N_6782,N_6333);
xnor U7587 (N_7587,N_6395,N_6004);
nand U7588 (N_7588,N_6712,N_6109);
or U7589 (N_7589,N_6337,N_6404);
nand U7590 (N_7590,N_6373,N_6970);
or U7591 (N_7591,N_6575,N_6330);
and U7592 (N_7592,N_6330,N_6034);
nand U7593 (N_7593,N_6149,N_6276);
nand U7594 (N_7594,N_6251,N_6094);
and U7595 (N_7595,N_6319,N_6982);
xnor U7596 (N_7596,N_6558,N_6693);
or U7597 (N_7597,N_6634,N_6623);
nand U7598 (N_7598,N_6166,N_6955);
and U7599 (N_7599,N_6450,N_6485);
and U7600 (N_7600,N_6949,N_6734);
nand U7601 (N_7601,N_6078,N_6681);
nand U7602 (N_7602,N_6378,N_6298);
nand U7603 (N_7603,N_6162,N_6079);
and U7604 (N_7604,N_6976,N_6552);
nor U7605 (N_7605,N_6097,N_6141);
and U7606 (N_7606,N_6461,N_6016);
or U7607 (N_7607,N_6737,N_6150);
nor U7608 (N_7608,N_6944,N_6107);
or U7609 (N_7609,N_6549,N_6663);
or U7610 (N_7610,N_6659,N_6820);
xnor U7611 (N_7611,N_6994,N_6401);
nor U7612 (N_7612,N_6284,N_6356);
or U7613 (N_7613,N_6959,N_6949);
or U7614 (N_7614,N_6881,N_6055);
nand U7615 (N_7615,N_6594,N_6235);
xnor U7616 (N_7616,N_6353,N_6348);
nor U7617 (N_7617,N_6617,N_6070);
nor U7618 (N_7618,N_6416,N_6190);
and U7619 (N_7619,N_6195,N_6042);
nor U7620 (N_7620,N_6113,N_6859);
and U7621 (N_7621,N_6836,N_6244);
and U7622 (N_7622,N_6720,N_6994);
nand U7623 (N_7623,N_6714,N_6560);
nor U7624 (N_7624,N_6603,N_6290);
and U7625 (N_7625,N_6016,N_6004);
or U7626 (N_7626,N_6896,N_6248);
xor U7627 (N_7627,N_6357,N_6962);
nand U7628 (N_7628,N_6000,N_6933);
and U7629 (N_7629,N_6417,N_6654);
xnor U7630 (N_7630,N_6480,N_6653);
and U7631 (N_7631,N_6428,N_6899);
or U7632 (N_7632,N_6199,N_6649);
xnor U7633 (N_7633,N_6891,N_6879);
nand U7634 (N_7634,N_6288,N_6266);
xnor U7635 (N_7635,N_6837,N_6736);
nand U7636 (N_7636,N_6941,N_6742);
nand U7637 (N_7637,N_6830,N_6640);
and U7638 (N_7638,N_6381,N_6644);
or U7639 (N_7639,N_6852,N_6163);
nand U7640 (N_7640,N_6484,N_6701);
nand U7641 (N_7641,N_6150,N_6851);
nand U7642 (N_7642,N_6138,N_6353);
and U7643 (N_7643,N_6840,N_6514);
or U7644 (N_7644,N_6778,N_6116);
and U7645 (N_7645,N_6824,N_6465);
or U7646 (N_7646,N_6415,N_6978);
or U7647 (N_7647,N_6156,N_6326);
or U7648 (N_7648,N_6085,N_6849);
and U7649 (N_7649,N_6721,N_6973);
and U7650 (N_7650,N_6995,N_6761);
nand U7651 (N_7651,N_6776,N_6280);
or U7652 (N_7652,N_6417,N_6128);
or U7653 (N_7653,N_6113,N_6926);
and U7654 (N_7654,N_6298,N_6713);
or U7655 (N_7655,N_6565,N_6122);
and U7656 (N_7656,N_6920,N_6804);
nand U7657 (N_7657,N_6425,N_6974);
xnor U7658 (N_7658,N_6155,N_6934);
xor U7659 (N_7659,N_6698,N_6761);
or U7660 (N_7660,N_6182,N_6315);
or U7661 (N_7661,N_6385,N_6312);
nand U7662 (N_7662,N_6526,N_6083);
or U7663 (N_7663,N_6523,N_6607);
or U7664 (N_7664,N_6641,N_6611);
and U7665 (N_7665,N_6488,N_6313);
and U7666 (N_7666,N_6400,N_6405);
nor U7667 (N_7667,N_6077,N_6670);
and U7668 (N_7668,N_6041,N_6427);
nor U7669 (N_7669,N_6784,N_6984);
and U7670 (N_7670,N_6236,N_6770);
nand U7671 (N_7671,N_6780,N_6323);
and U7672 (N_7672,N_6684,N_6347);
nand U7673 (N_7673,N_6958,N_6073);
and U7674 (N_7674,N_6298,N_6413);
nand U7675 (N_7675,N_6203,N_6845);
nor U7676 (N_7676,N_6216,N_6950);
and U7677 (N_7677,N_6436,N_6570);
xnor U7678 (N_7678,N_6531,N_6200);
and U7679 (N_7679,N_6452,N_6464);
and U7680 (N_7680,N_6355,N_6685);
and U7681 (N_7681,N_6454,N_6414);
and U7682 (N_7682,N_6238,N_6830);
nor U7683 (N_7683,N_6141,N_6242);
xnor U7684 (N_7684,N_6191,N_6141);
and U7685 (N_7685,N_6331,N_6622);
nor U7686 (N_7686,N_6933,N_6441);
xnor U7687 (N_7687,N_6585,N_6293);
xor U7688 (N_7688,N_6603,N_6933);
xnor U7689 (N_7689,N_6066,N_6446);
and U7690 (N_7690,N_6862,N_6320);
or U7691 (N_7691,N_6922,N_6096);
and U7692 (N_7692,N_6320,N_6106);
nand U7693 (N_7693,N_6105,N_6212);
and U7694 (N_7694,N_6846,N_6634);
nor U7695 (N_7695,N_6023,N_6841);
nor U7696 (N_7696,N_6629,N_6499);
and U7697 (N_7697,N_6742,N_6529);
or U7698 (N_7698,N_6842,N_6012);
nand U7699 (N_7699,N_6671,N_6976);
and U7700 (N_7700,N_6977,N_6214);
nor U7701 (N_7701,N_6804,N_6140);
and U7702 (N_7702,N_6640,N_6096);
nand U7703 (N_7703,N_6968,N_6341);
xnor U7704 (N_7704,N_6730,N_6355);
and U7705 (N_7705,N_6722,N_6970);
nand U7706 (N_7706,N_6998,N_6443);
or U7707 (N_7707,N_6838,N_6473);
nor U7708 (N_7708,N_6829,N_6824);
and U7709 (N_7709,N_6209,N_6123);
nor U7710 (N_7710,N_6058,N_6908);
and U7711 (N_7711,N_6202,N_6771);
nor U7712 (N_7712,N_6813,N_6472);
nor U7713 (N_7713,N_6501,N_6567);
nand U7714 (N_7714,N_6388,N_6683);
or U7715 (N_7715,N_6503,N_6943);
and U7716 (N_7716,N_6447,N_6030);
nor U7717 (N_7717,N_6854,N_6541);
xor U7718 (N_7718,N_6264,N_6578);
nor U7719 (N_7719,N_6736,N_6089);
nor U7720 (N_7720,N_6715,N_6180);
or U7721 (N_7721,N_6960,N_6032);
xnor U7722 (N_7722,N_6894,N_6508);
nand U7723 (N_7723,N_6083,N_6344);
nor U7724 (N_7724,N_6176,N_6201);
or U7725 (N_7725,N_6365,N_6887);
nand U7726 (N_7726,N_6904,N_6821);
and U7727 (N_7727,N_6236,N_6348);
and U7728 (N_7728,N_6178,N_6275);
or U7729 (N_7729,N_6103,N_6573);
and U7730 (N_7730,N_6884,N_6874);
and U7731 (N_7731,N_6907,N_6871);
and U7732 (N_7732,N_6939,N_6169);
and U7733 (N_7733,N_6984,N_6753);
nor U7734 (N_7734,N_6213,N_6944);
nor U7735 (N_7735,N_6590,N_6519);
nor U7736 (N_7736,N_6950,N_6231);
nor U7737 (N_7737,N_6340,N_6841);
and U7738 (N_7738,N_6846,N_6107);
nor U7739 (N_7739,N_6382,N_6568);
nand U7740 (N_7740,N_6995,N_6862);
or U7741 (N_7741,N_6460,N_6097);
nor U7742 (N_7742,N_6036,N_6640);
nand U7743 (N_7743,N_6325,N_6614);
nor U7744 (N_7744,N_6042,N_6462);
or U7745 (N_7745,N_6778,N_6354);
or U7746 (N_7746,N_6313,N_6659);
or U7747 (N_7747,N_6790,N_6976);
and U7748 (N_7748,N_6836,N_6431);
or U7749 (N_7749,N_6651,N_6211);
nor U7750 (N_7750,N_6543,N_6721);
nor U7751 (N_7751,N_6114,N_6385);
or U7752 (N_7752,N_6963,N_6388);
nand U7753 (N_7753,N_6860,N_6212);
and U7754 (N_7754,N_6468,N_6708);
xnor U7755 (N_7755,N_6610,N_6014);
and U7756 (N_7756,N_6538,N_6160);
or U7757 (N_7757,N_6559,N_6768);
xor U7758 (N_7758,N_6541,N_6275);
and U7759 (N_7759,N_6233,N_6690);
and U7760 (N_7760,N_6484,N_6466);
xor U7761 (N_7761,N_6592,N_6162);
nand U7762 (N_7762,N_6666,N_6020);
and U7763 (N_7763,N_6093,N_6079);
or U7764 (N_7764,N_6164,N_6791);
nand U7765 (N_7765,N_6511,N_6679);
nor U7766 (N_7766,N_6855,N_6714);
nand U7767 (N_7767,N_6172,N_6642);
nor U7768 (N_7768,N_6126,N_6611);
nand U7769 (N_7769,N_6417,N_6326);
and U7770 (N_7770,N_6637,N_6774);
and U7771 (N_7771,N_6514,N_6421);
nor U7772 (N_7772,N_6637,N_6933);
nand U7773 (N_7773,N_6424,N_6420);
and U7774 (N_7774,N_6848,N_6033);
or U7775 (N_7775,N_6258,N_6035);
nand U7776 (N_7776,N_6439,N_6882);
nor U7777 (N_7777,N_6998,N_6036);
or U7778 (N_7778,N_6712,N_6143);
nor U7779 (N_7779,N_6253,N_6365);
xor U7780 (N_7780,N_6995,N_6407);
nor U7781 (N_7781,N_6091,N_6968);
nand U7782 (N_7782,N_6870,N_6695);
and U7783 (N_7783,N_6699,N_6858);
or U7784 (N_7784,N_6758,N_6299);
and U7785 (N_7785,N_6171,N_6457);
nor U7786 (N_7786,N_6109,N_6089);
nor U7787 (N_7787,N_6663,N_6091);
and U7788 (N_7788,N_6096,N_6690);
nor U7789 (N_7789,N_6456,N_6268);
nand U7790 (N_7790,N_6908,N_6086);
nand U7791 (N_7791,N_6834,N_6629);
or U7792 (N_7792,N_6123,N_6504);
nor U7793 (N_7793,N_6017,N_6039);
or U7794 (N_7794,N_6904,N_6468);
nor U7795 (N_7795,N_6106,N_6588);
nor U7796 (N_7796,N_6652,N_6199);
or U7797 (N_7797,N_6863,N_6361);
and U7798 (N_7798,N_6278,N_6200);
xor U7799 (N_7799,N_6783,N_6627);
or U7800 (N_7800,N_6061,N_6807);
nand U7801 (N_7801,N_6669,N_6675);
nand U7802 (N_7802,N_6851,N_6176);
nand U7803 (N_7803,N_6357,N_6576);
nor U7804 (N_7804,N_6429,N_6800);
nor U7805 (N_7805,N_6977,N_6850);
nand U7806 (N_7806,N_6923,N_6514);
nor U7807 (N_7807,N_6502,N_6139);
nand U7808 (N_7808,N_6485,N_6553);
nand U7809 (N_7809,N_6490,N_6036);
nand U7810 (N_7810,N_6365,N_6132);
and U7811 (N_7811,N_6523,N_6561);
or U7812 (N_7812,N_6004,N_6980);
or U7813 (N_7813,N_6920,N_6666);
or U7814 (N_7814,N_6477,N_6170);
nor U7815 (N_7815,N_6331,N_6289);
nand U7816 (N_7816,N_6019,N_6763);
nor U7817 (N_7817,N_6039,N_6203);
and U7818 (N_7818,N_6907,N_6356);
nand U7819 (N_7819,N_6246,N_6265);
nor U7820 (N_7820,N_6965,N_6576);
or U7821 (N_7821,N_6136,N_6039);
and U7822 (N_7822,N_6928,N_6722);
and U7823 (N_7823,N_6336,N_6225);
nand U7824 (N_7824,N_6529,N_6597);
nand U7825 (N_7825,N_6474,N_6408);
nand U7826 (N_7826,N_6770,N_6495);
nand U7827 (N_7827,N_6143,N_6763);
and U7828 (N_7828,N_6357,N_6716);
or U7829 (N_7829,N_6865,N_6092);
and U7830 (N_7830,N_6044,N_6628);
and U7831 (N_7831,N_6366,N_6970);
or U7832 (N_7832,N_6127,N_6305);
nand U7833 (N_7833,N_6107,N_6171);
or U7834 (N_7834,N_6972,N_6593);
nor U7835 (N_7835,N_6478,N_6642);
nor U7836 (N_7836,N_6369,N_6641);
xnor U7837 (N_7837,N_6053,N_6713);
or U7838 (N_7838,N_6551,N_6626);
nand U7839 (N_7839,N_6814,N_6800);
and U7840 (N_7840,N_6950,N_6975);
or U7841 (N_7841,N_6130,N_6102);
xnor U7842 (N_7842,N_6114,N_6762);
nor U7843 (N_7843,N_6997,N_6011);
and U7844 (N_7844,N_6871,N_6123);
nand U7845 (N_7845,N_6676,N_6132);
or U7846 (N_7846,N_6058,N_6752);
nor U7847 (N_7847,N_6444,N_6531);
nand U7848 (N_7848,N_6698,N_6593);
nor U7849 (N_7849,N_6594,N_6669);
nand U7850 (N_7850,N_6057,N_6607);
nor U7851 (N_7851,N_6227,N_6987);
xnor U7852 (N_7852,N_6660,N_6932);
or U7853 (N_7853,N_6161,N_6372);
nor U7854 (N_7854,N_6578,N_6945);
nand U7855 (N_7855,N_6870,N_6156);
and U7856 (N_7856,N_6494,N_6876);
or U7857 (N_7857,N_6552,N_6731);
xor U7858 (N_7858,N_6994,N_6310);
nand U7859 (N_7859,N_6456,N_6751);
and U7860 (N_7860,N_6420,N_6761);
and U7861 (N_7861,N_6477,N_6599);
or U7862 (N_7862,N_6298,N_6758);
or U7863 (N_7863,N_6335,N_6135);
or U7864 (N_7864,N_6997,N_6939);
nand U7865 (N_7865,N_6595,N_6137);
nand U7866 (N_7866,N_6429,N_6453);
and U7867 (N_7867,N_6040,N_6713);
or U7868 (N_7868,N_6628,N_6411);
xnor U7869 (N_7869,N_6433,N_6659);
xor U7870 (N_7870,N_6614,N_6735);
nand U7871 (N_7871,N_6574,N_6216);
or U7872 (N_7872,N_6979,N_6578);
and U7873 (N_7873,N_6543,N_6628);
nand U7874 (N_7874,N_6730,N_6616);
nor U7875 (N_7875,N_6516,N_6623);
nand U7876 (N_7876,N_6422,N_6152);
xor U7877 (N_7877,N_6786,N_6622);
or U7878 (N_7878,N_6776,N_6066);
xnor U7879 (N_7879,N_6920,N_6860);
nand U7880 (N_7880,N_6338,N_6811);
or U7881 (N_7881,N_6096,N_6583);
xnor U7882 (N_7882,N_6925,N_6813);
nand U7883 (N_7883,N_6245,N_6892);
nand U7884 (N_7884,N_6591,N_6440);
and U7885 (N_7885,N_6576,N_6593);
nor U7886 (N_7886,N_6123,N_6713);
and U7887 (N_7887,N_6340,N_6196);
and U7888 (N_7888,N_6322,N_6514);
nand U7889 (N_7889,N_6815,N_6632);
and U7890 (N_7890,N_6414,N_6856);
nor U7891 (N_7891,N_6871,N_6446);
nand U7892 (N_7892,N_6373,N_6297);
nor U7893 (N_7893,N_6617,N_6339);
nand U7894 (N_7894,N_6081,N_6023);
and U7895 (N_7895,N_6301,N_6314);
or U7896 (N_7896,N_6654,N_6526);
or U7897 (N_7897,N_6404,N_6760);
and U7898 (N_7898,N_6764,N_6698);
nand U7899 (N_7899,N_6714,N_6125);
or U7900 (N_7900,N_6547,N_6147);
nor U7901 (N_7901,N_6671,N_6805);
nor U7902 (N_7902,N_6837,N_6105);
nor U7903 (N_7903,N_6917,N_6845);
and U7904 (N_7904,N_6406,N_6846);
and U7905 (N_7905,N_6128,N_6424);
xnor U7906 (N_7906,N_6084,N_6060);
nor U7907 (N_7907,N_6448,N_6700);
or U7908 (N_7908,N_6554,N_6085);
and U7909 (N_7909,N_6361,N_6917);
nor U7910 (N_7910,N_6606,N_6289);
xnor U7911 (N_7911,N_6665,N_6397);
nor U7912 (N_7912,N_6119,N_6443);
or U7913 (N_7913,N_6116,N_6118);
or U7914 (N_7914,N_6721,N_6335);
xnor U7915 (N_7915,N_6548,N_6294);
or U7916 (N_7916,N_6267,N_6283);
and U7917 (N_7917,N_6980,N_6870);
nand U7918 (N_7918,N_6716,N_6968);
or U7919 (N_7919,N_6230,N_6448);
or U7920 (N_7920,N_6394,N_6228);
nor U7921 (N_7921,N_6239,N_6383);
or U7922 (N_7922,N_6994,N_6413);
nor U7923 (N_7923,N_6413,N_6677);
xor U7924 (N_7924,N_6990,N_6363);
or U7925 (N_7925,N_6529,N_6526);
and U7926 (N_7926,N_6971,N_6811);
or U7927 (N_7927,N_6776,N_6131);
and U7928 (N_7928,N_6605,N_6354);
or U7929 (N_7929,N_6091,N_6401);
nor U7930 (N_7930,N_6368,N_6175);
and U7931 (N_7931,N_6384,N_6656);
and U7932 (N_7932,N_6803,N_6554);
nand U7933 (N_7933,N_6872,N_6826);
nand U7934 (N_7934,N_6417,N_6437);
nor U7935 (N_7935,N_6982,N_6861);
xnor U7936 (N_7936,N_6396,N_6094);
nor U7937 (N_7937,N_6807,N_6612);
or U7938 (N_7938,N_6649,N_6354);
nand U7939 (N_7939,N_6936,N_6921);
nor U7940 (N_7940,N_6188,N_6280);
nand U7941 (N_7941,N_6212,N_6538);
nor U7942 (N_7942,N_6567,N_6775);
nor U7943 (N_7943,N_6190,N_6223);
nor U7944 (N_7944,N_6186,N_6039);
and U7945 (N_7945,N_6398,N_6818);
nand U7946 (N_7946,N_6053,N_6478);
nand U7947 (N_7947,N_6228,N_6113);
and U7948 (N_7948,N_6512,N_6712);
or U7949 (N_7949,N_6861,N_6606);
or U7950 (N_7950,N_6832,N_6939);
and U7951 (N_7951,N_6070,N_6559);
or U7952 (N_7952,N_6805,N_6551);
and U7953 (N_7953,N_6027,N_6765);
nor U7954 (N_7954,N_6371,N_6974);
or U7955 (N_7955,N_6631,N_6726);
and U7956 (N_7956,N_6775,N_6121);
xnor U7957 (N_7957,N_6676,N_6772);
nand U7958 (N_7958,N_6633,N_6472);
or U7959 (N_7959,N_6621,N_6934);
nand U7960 (N_7960,N_6924,N_6666);
nand U7961 (N_7961,N_6681,N_6858);
or U7962 (N_7962,N_6128,N_6917);
and U7963 (N_7963,N_6895,N_6428);
nand U7964 (N_7964,N_6333,N_6291);
xor U7965 (N_7965,N_6931,N_6327);
nand U7966 (N_7966,N_6736,N_6056);
or U7967 (N_7967,N_6352,N_6594);
and U7968 (N_7968,N_6952,N_6429);
and U7969 (N_7969,N_6286,N_6231);
nand U7970 (N_7970,N_6631,N_6639);
nor U7971 (N_7971,N_6466,N_6872);
nand U7972 (N_7972,N_6124,N_6671);
or U7973 (N_7973,N_6355,N_6514);
nor U7974 (N_7974,N_6732,N_6178);
nor U7975 (N_7975,N_6115,N_6251);
nand U7976 (N_7976,N_6566,N_6082);
nand U7977 (N_7977,N_6601,N_6638);
and U7978 (N_7978,N_6903,N_6145);
or U7979 (N_7979,N_6189,N_6009);
and U7980 (N_7980,N_6251,N_6419);
nor U7981 (N_7981,N_6207,N_6762);
and U7982 (N_7982,N_6020,N_6600);
nand U7983 (N_7983,N_6304,N_6252);
nor U7984 (N_7984,N_6690,N_6299);
or U7985 (N_7985,N_6865,N_6692);
or U7986 (N_7986,N_6066,N_6103);
and U7987 (N_7987,N_6475,N_6266);
or U7988 (N_7988,N_6366,N_6207);
or U7989 (N_7989,N_6940,N_6441);
and U7990 (N_7990,N_6045,N_6823);
nand U7991 (N_7991,N_6915,N_6457);
and U7992 (N_7992,N_6454,N_6468);
nor U7993 (N_7993,N_6869,N_6241);
and U7994 (N_7994,N_6231,N_6303);
nand U7995 (N_7995,N_6245,N_6748);
and U7996 (N_7996,N_6472,N_6502);
or U7997 (N_7997,N_6950,N_6714);
nand U7998 (N_7998,N_6710,N_6260);
and U7999 (N_7999,N_6472,N_6037);
nand U8000 (N_8000,N_7830,N_7740);
and U8001 (N_8001,N_7037,N_7812);
or U8002 (N_8002,N_7182,N_7527);
nor U8003 (N_8003,N_7891,N_7264);
or U8004 (N_8004,N_7026,N_7315);
or U8005 (N_8005,N_7077,N_7146);
nor U8006 (N_8006,N_7250,N_7633);
nand U8007 (N_8007,N_7177,N_7660);
nor U8008 (N_8008,N_7137,N_7242);
or U8009 (N_8009,N_7678,N_7130);
nand U8010 (N_8010,N_7961,N_7796);
and U8011 (N_8011,N_7430,N_7200);
and U8012 (N_8012,N_7846,N_7156);
or U8013 (N_8013,N_7931,N_7682);
nand U8014 (N_8014,N_7958,N_7576);
or U8015 (N_8015,N_7963,N_7174);
nor U8016 (N_8016,N_7870,N_7067);
nand U8017 (N_8017,N_7967,N_7916);
nand U8018 (N_8018,N_7380,N_7256);
and U8019 (N_8019,N_7120,N_7694);
and U8020 (N_8020,N_7378,N_7737);
xor U8021 (N_8021,N_7586,N_7573);
nor U8022 (N_8022,N_7897,N_7868);
and U8023 (N_8023,N_7747,N_7018);
nand U8024 (N_8024,N_7447,N_7934);
and U8025 (N_8025,N_7939,N_7493);
nand U8026 (N_8026,N_7713,N_7483);
nand U8027 (N_8027,N_7331,N_7986);
or U8028 (N_8028,N_7650,N_7236);
or U8029 (N_8029,N_7635,N_7983);
nand U8030 (N_8030,N_7571,N_7754);
and U8031 (N_8031,N_7270,N_7498);
and U8032 (N_8032,N_7759,N_7941);
and U8033 (N_8033,N_7071,N_7136);
and U8034 (N_8034,N_7770,N_7122);
nand U8035 (N_8035,N_7887,N_7959);
or U8036 (N_8036,N_7422,N_7040);
and U8037 (N_8037,N_7679,N_7881);
or U8038 (N_8038,N_7393,N_7502);
or U8039 (N_8039,N_7508,N_7415);
and U8040 (N_8040,N_7839,N_7632);
and U8041 (N_8041,N_7160,N_7003);
or U8042 (N_8042,N_7534,N_7608);
and U8043 (N_8043,N_7738,N_7423);
xor U8044 (N_8044,N_7662,N_7952);
and U8045 (N_8045,N_7712,N_7186);
xnor U8046 (N_8046,N_7278,N_7735);
and U8047 (N_8047,N_7700,N_7723);
and U8048 (N_8048,N_7869,N_7115);
nand U8049 (N_8049,N_7057,N_7074);
or U8050 (N_8050,N_7613,N_7239);
or U8051 (N_8051,N_7305,N_7257);
nor U8052 (N_8052,N_7478,N_7756);
nor U8053 (N_8053,N_7020,N_7129);
xor U8054 (N_8054,N_7228,N_7676);
or U8055 (N_8055,N_7143,N_7794);
or U8056 (N_8056,N_7299,N_7234);
or U8057 (N_8057,N_7776,N_7086);
xnor U8058 (N_8058,N_7989,N_7968);
or U8059 (N_8059,N_7368,N_7933);
nand U8060 (N_8060,N_7164,N_7334);
or U8061 (N_8061,N_7545,N_7243);
or U8062 (N_8062,N_7010,N_7094);
or U8063 (N_8063,N_7029,N_7926);
nand U8064 (N_8064,N_7157,N_7212);
nand U8065 (N_8065,N_7117,N_7511);
nand U8066 (N_8066,N_7826,N_7799);
nor U8067 (N_8067,N_7861,N_7021);
and U8068 (N_8068,N_7189,N_7286);
and U8069 (N_8069,N_7804,N_7567);
and U8070 (N_8070,N_7978,N_7943);
nor U8071 (N_8071,N_7731,N_7283);
or U8072 (N_8072,N_7784,N_7128);
and U8073 (N_8073,N_7798,N_7932);
nor U8074 (N_8074,N_7199,N_7670);
nor U8075 (N_8075,N_7039,N_7742);
and U8076 (N_8076,N_7051,N_7760);
nand U8077 (N_8077,N_7894,N_7795);
nor U8078 (N_8078,N_7452,N_7644);
or U8079 (N_8079,N_7848,N_7651);
xor U8080 (N_8080,N_7639,N_7762);
nor U8081 (N_8081,N_7523,N_7123);
xor U8082 (N_8082,N_7597,N_7956);
or U8083 (N_8083,N_7641,N_7488);
and U8084 (N_8084,N_7079,N_7110);
nor U8085 (N_8085,N_7703,N_7522);
or U8086 (N_8086,N_7335,N_7268);
and U8087 (N_8087,N_7339,N_7974);
xnor U8088 (N_8088,N_7169,N_7455);
nand U8089 (N_8089,N_7363,N_7290);
or U8090 (N_8090,N_7387,N_7945);
nand U8091 (N_8091,N_7697,N_7813);
nor U8092 (N_8092,N_7882,N_7831);
and U8093 (N_8093,N_7828,N_7995);
or U8094 (N_8094,N_7457,N_7246);
nand U8095 (N_8095,N_7458,N_7816);
xnor U8096 (N_8096,N_7574,N_7255);
nor U8097 (N_8097,N_7092,N_7991);
nor U8098 (N_8098,N_7500,N_7377);
nand U8099 (N_8099,N_7992,N_7004);
and U8100 (N_8100,N_7180,N_7016);
nand U8101 (N_8101,N_7902,N_7272);
or U8102 (N_8102,N_7207,N_7789);
nor U8103 (N_8103,N_7960,N_7862);
or U8104 (N_8104,N_7125,N_7658);
nand U8105 (N_8105,N_7203,N_7287);
and U8106 (N_8106,N_7540,N_7181);
and U8107 (N_8107,N_7605,N_7197);
nand U8108 (N_8108,N_7350,N_7011);
or U8109 (N_8109,N_7060,N_7345);
and U8110 (N_8110,N_7076,N_7819);
nand U8111 (N_8111,N_7313,N_7744);
nor U8112 (N_8112,N_7898,N_7730);
xnor U8113 (N_8113,N_7844,N_7957);
or U8114 (N_8114,N_7520,N_7426);
or U8115 (N_8115,N_7318,N_7022);
nor U8116 (N_8116,N_7303,N_7410);
nand U8117 (N_8117,N_7329,N_7873);
or U8118 (N_8118,N_7854,N_7507);
or U8119 (N_8119,N_7672,N_7253);
xnor U8120 (N_8120,N_7494,N_7505);
and U8121 (N_8121,N_7400,N_7656);
xnor U8122 (N_8122,N_7757,N_7519);
nor U8123 (N_8123,N_7954,N_7971);
or U8124 (N_8124,N_7667,N_7791);
or U8125 (N_8125,N_7215,N_7102);
nor U8126 (N_8126,N_7763,N_7080);
or U8127 (N_8127,N_7401,N_7402);
or U8128 (N_8128,N_7793,N_7803);
nand U8129 (N_8129,N_7416,N_7726);
nor U8130 (N_8130,N_7893,N_7013);
nand U8131 (N_8131,N_7973,N_7688);
nand U8132 (N_8132,N_7225,N_7462);
nand U8133 (N_8133,N_7440,N_7443);
nor U8134 (N_8134,N_7563,N_7372);
and U8135 (N_8135,N_7147,N_7418);
or U8136 (N_8136,N_7301,N_7965);
nand U8137 (N_8137,N_7056,N_7063);
nor U8138 (N_8138,N_7994,N_7309);
or U8139 (N_8139,N_7254,N_7914);
nor U8140 (N_8140,N_7346,N_7370);
nand U8141 (N_8141,N_7161,N_7909);
and U8142 (N_8142,N_7775,N_7850);
nand U8143 (N_8143,N_7005,N_7023);
nand U8144 (N_8144,N_7944,N_7646);
and U8145 (N_8145,N_7665,N_7612);
or U8146 (N_8146,N_7513,N_7925);
and U8147 (N_8147,N_7714,N_7461);
nand U8148 (N_8148,N_7442,N_7319);
nand U8149 (N_8149,N_7361,N_7431);
or U8150 (N_8150,N_7090,N_7012);
nand U8151 (N_8151,N_7981,N_7222);
or U8152 (N_8152,N_7541,N_7787);
nor U8153 (N_8153,N_7104,N_7988);
nand U8154 (N_8154,N_7620,N_7293);
and U8155 (N_8155,N_7155,N_7942);
nand U8156 (N_8156,N_7546,N_7477);
nor U8157 (N_8157,N_7214,N_7836);
xor U8158 (N_8158,N_7360,N_7645);
nand U8159 (N_8159,N_7950,N_7817);
nand U8160 (N_8160,N_7908,N_7069);
or U8161 (N_8161,N_7411,N_7030);
nor U8162 (N_8162,N_7053,N_7216);
nor U8163 (N_8163,N_7751,N_7584);
and U8164 (N_8164,N_7716,N_7187);
nor U8165 (N_8165,N_7248,N_7677);
nor U8166 (N_8166,N_7226,N_7824);
nand U8167 (N_8167,N_7434,N_7093);
or U8168 (N_8168,N_7877,N_7445);
or U8169 (N_8169,N_7525,N_7111);
or U8170 (N_8170,N_7482,N_7112);
xor U8171 (N_8171,N_7711,N_7055);
or U8172 (N_8172,N_7395,N_7915);
or U8173 (N_8173,N_7581,N_7427);
and U8174 (N_8174,N_7918,N_7359);
nand U8175 (N_8175,N_7347,N_7785);
nor U8176 (N_8176,N_7885,N_7000);
nand U8177 (N_8177,N_7634,N_7383);
nand U8178 (N_8178,N_7900,N_7481);
nor U8179 (N_8179,N_7348,N_7603);
nor U8180 (N_8180,N_7772,N_7209);
or U8181 (N_8181,N_7341,N_7962);
nor U8182 (N_8182,N_7453,N_7947);
and U8183 (N_8183,N_7859,N_7970);
nand U8184 (N_8184,N_7321,N_7134);
or U8185 (N_8185,N_7038,N_7154);
nand U8186 (N_8186,N_7072,N_7999);
xnor U8187 (N_8187,N_7116,N_7251);
or U8188 (N_8188,N_7152,N_7923);
or U8189 (N_8189,N_7183,N_7903);
nor U8190 (N_8190,N_7940,N_7718);
nand U8191 (N_8191,N_7876,N_7252);
or U8192 (N_8192,N_7066,N_7237);
or U8193 (N_8193,N_7556,N_7185);
xor U8194 (N_8194,N_7463,N_7704);
nor U8195 (N_8195,N_7668,N_7460);
and U8196 (N_8196,N_7514,N_7244);
xor U8197 (N_8197,N_7001,N_7166);
nand U8198 (N_8198,N_7337,N_7698);
nor U8199 (N_8199,N_7886,N_7165);
or U8200 (N_8200,N_7807,N_7459);
nor U8201 (N_8201,N_7298,N_7946);
nand U8202 (N_8202,N_7930,N_7213);
xnor U8203 (N_8203,N_7366,N_7709);
xor U8204 (N_8204,N_7087,N_7376);
nand U8205 (N_8205,N_7008,N_7899);
and U8206 (N_8206,N_7764,N_7669);
or U8207 (N_8207,N_7564,N_7230);
xnor U8208 (N_8208,N_7542,N_7657);
and U8209 (N_8209,N_7465,N_7352);
nor U8210 (N_8210,N_7035,N_7538);
nor U8211 (N_8211,N_7739,N_7889);
nor U8212 (N_8212,N_7977,N_7241);
nand U8213 (N_8213,N_7727,N_7162);
nor U8214 (N_8214,N_7768,N_7951);
and U8215 (N_8215,N_7607,N_7953);
xnor U8216 (N_8216,N_7625,N_7671);
and U8217 (N_8217,N_7195,N_7972);
nand U8218 (N_8218,N_7654,N_7158);
nor U8219 (N_8219,N_7385,N_7725);
nand U8220 (N_8220,N_7687,N_7064);
nand U8221 (N_8221,N_7690,N_7238);
or U8222 (N_8222,N_7843,N_7466);
nor U8223 (N_8223,N_7872,N_7476);
xnor U8224 (N_8224,N_7998,N_7856);
or U8225 (N_8225,N_7528,N_7598);
nor U8226 (N_8226,N_7708,N_7548);
or U8227 (N_8227,N_7838,N_7446);
or U8228 (N_8228,N_7083,N_7219);
nand U8229 (N_8229,N_7314,N_7405);
or U8230 (N_8230,N_7680,N_7097);
nand U8231 (N_8231,N_7509,N_7913);
nor U8232 (N_8232,N_7379,N_7451);
nand U8233 (N_8233,N_7503,N_7444);
nand U8234 (N_8234,N_7653,N_7622);
nand U8235 (N_8235,N_7719,N_7306);
nor U8236 (N_8236,N_7617,N_7629);
nor U8237 (N_8237,N_7765,N_7788);
or U8238 (N_8238,N_7752,N_7232);
and U8239 (N_8239,N_7937,N_7472);
nand U8240 (N_8240,N_7865,N_7096);
nor U8241 (N_8241,N_7261,N_7663);
xnor U8242 (N_8242,N_7533,N_7374);
or U8243 (N_8243,N_7874,N_7135);
or U8244 (N_8244,N_7295,N_7621);
or U8245 (N_8245,N_7208,N_7474);
nand U8246 (N_8246,N_7172,N_7741);
nor U8247 (N_8247,N_7652,N_7845);
nor U8248 (N_8248,N_7602,N_7570);
nand U8249 (N_8249,N_7088,N_7420);
nand U8250 (N_8250,N_7371,N_7437);
nor U8251 (N_8251,N_7267,N_7818);
and U8252 (N_8252,N_7375,N_7070);
nand U8253 (N_8253,N_7275,N_7666);
nand U8254 (N_8254,N_7766,N_7864);
nand U8255 (N_8255,N_7468,N_7099);
nor U8256 (N_8256,N_7260,N_7851);
xor U8257 (N_8257,N_7928,N_7578);
xnor U8258 (N_8258,N_7492,N_7684);
nand U8259 (N_8259,N_7041,N_7743);
nand U8260 (N_8260,N_7204,N_7028);
and U8261 (N_8261,N_7414,N_7132);
or U8262 (N_8262,N_7810,N_7769);
and U8263 (N_8263,N_7312,N_7349);
nor U8264 (N_8264,N_7484,N_7288);
and U8265 (N_8265,N_7042,N_7240);
nor U8266 (N_8266,N_7618,N_7495);
or U8267 (N_8267,N_7131,N_7342);
xnor U8268 (N_8268,N_7210,N_7580);
xnor U8269 (N_8269,N_7211,N_7497);
or U8270 (N_8270,N_7728,N_7373);
or U8271 (N_8271,N_7336,N_7606);
nand U8272 (N_8272,N_7328,N_7823);
xor U8273 (N_8273,N_7114,N_7834);
xnor U8274 (N_8274,N_7343,N_7340);
xor U8275 (N_8275,N_7168,N_7875);
nor U8276 (N_8276,N_7192,N_7761);
nor U8277 (N_8277,N_7516,N_7753);
xnor U8278 (N_8278,N_7085,N_7058);
or U8279 (N_8279,N_7594,N_7565);
nand U8280 (N_8280,N_7140,N_7002);
or U8281 (N_8281,N_7691,N_7351);
nor U8282 (N_8282,N_7681,N_7802);
and U8283 (N_8283,N_7296,N_7424);
or U8284 (N_8284,N_7686,N_7307);
and U8285 (N_8285,N_7901,N_7867);
and U8286 (N_8286,N_7386,N_7223);
nor U8287 (N_8287,N_7229,N_7358);
and U8288 (N_8288,N_7979,N_7715);
or U8289 (N_8289,N_7403,N_7218);
or U8290 (N_8290,N_7732,N_7389);
nand U8291 (N_8291,N_7569,N_7938);
or U8292 (N_8292,N_7510,N_7126);
and U8293 (N_8293,N_7638,N_7227);
and U8294 (N_8294,N_7025,N_7544);
nand U8295 (N_8295,N_7078,N_7600);
nor U8296 (N_8296,N_7279,N_7014);
nor U8297 (N_8297,N_7664,N_7863);
or U8298 (N_8298,N_7579,N_7936);
or U8299 (N_8299,N_7593,N_7693);
or U8300 (N_8300,N_7475,N_7982);
nand U8301 (N_8301,N_7758,N_7969);
xnor U8302 (N_8302,N_7746,N_7138);
and U8303 (N_8303,N_7683,N_7878);
nand U8304 (N_8304,N_7549,N_7630);
or U8305 (N_8305,N_7109,N_7193);
xnor U8306 (N_8306,N_7551,N_7024);
nor U8307 (N_8307,N_7550,N_7710);
and U8308 (N_8308,N_7141,N_7432);
and U8309 (N_8309,N_7610,N_7280);
or U8310 (N_8310,N_7249,N_7486);
nand U8311 (N_8311,N_7557,N_7043);
nor U8312 (N_8312,N_7879,N_7044);
nor U8313 (N_8313,N_7852,N_7748);
nand U8314 (N_8314,N_7188,N_7499);
and U8315 (N_8315,N_7696,N_7771);
or U8316 (N_8316,N_7045,N_7450);
xnor U8317 (N_8317,N_7205,N_7628);
nand U8318 (N_8318,N_7515,N_7398);
or U8319 (N_8319,N_7105,N_7033);
or U8320 (N_8320,N_7643,N_7419);
and U8321 (N_8321,N_7521,N_7289);
nor U8322 (N_8322,N_7006,N_7572);
xnor U8323 (N_8323,N_7456,N_7441);
and U8324 (N_8324,N_7435,N_7566);
nor U8325 (N_8325,N_7479,N_7101);
or U8326 (N_8326,N_7036,N_7220);
xor U8327 (N_8327,N_7404,N_7027);
nand U8328 (N_8328,N_7847,N_7291);
nand U8329 (N_8329,N_7190,N_7439);
nand U8330 (N_8330,N_7536,N_7855);
or U8331 (N_8331,N_7031,N_7568);
nand U8332 (N_8332,N_7655,N_7783);
nor U8333 (N_8333,N_7118,N_7692);
xnor U8334 (N_8334,N_7052,N_7050);
or U8335 (N_8335,N_7489,N_7326);
nand U8336 (N_8336,N_7706,N_7107);
or U8337 (N_8337,N_7317,N_7320);
xor U8338 (N_8338,N_7394,N_7091);
or U8339 (N_8339,N_7562,N_7391);
and U8340 (N_8340,N_7535,N_7592);
xnor U8341 (N_8341,N_7832,N_7811);
or U8342 (N_8342,N_7661,N_7619);
nor U8343 (N_8343,N_7469,N_7098);
nand U8344 (N_8344,N_7695,N_7993);
xor U8345 (N_8345,N_7647,N_7559);
and U8346 (N_8346,N_7631,N_7364);
and U8347 (N_8347,N_7191,N_7532);
or U8348 (N_8348,N_7552,N_7736);
or U8349 (N_8349,N_7139,N_7009);
or U8350 (N_8350,N_7833,N_7159);
and U8351 (N_8351,N_7061,N_7108);
or U8352 (N_8352,N_7910,N_7384);
nor U8353 (N_8353,N_7263,N_7642);
nand U8354 (N_8354,N_7805,N_7302);
or U8355 (N_8355,N_7310,N_7984);
and U8356 (N_8356,N_7919,N_7124);
nand U8357 (N_8357,N_7381,N_7448);
xnor U8358 (N_8358,N_7113,N_7178);
or U8359 (N_8359,N_7777,N_7814);
and U8360 (N_8360,N_7582,N_7007);
nor U8361 (N_8361,N_7106,N_7575);
nor U8362 (N_8362,N_7614,N_7840);
or U8363 (N_8363,N_7888,N_7705);
nand U8364 (N_8364,N_7323,N_7827);
nor U8365 (N_8365,N_7526,N_7369);
and U8366 (N_8366,N_7425,N_7906);
and U8367 (N_8367,N_7196,N_7734);
nand U8368 (N_8368,N_7356,N_7412);
or U8369 (N_8369,N_7858,N_7912);
or U8370 (N_8370,N_7322,N_7924);
nor U8371 (N_8371,N_7217,N_7773);
nor U8372 (N_8372,N_7717,N_7194);
nor U8373 (N_8373,N_7673,N_7512);
xnor U8374 (N_8374,N_7648,N_7324);
or U8375 (N_8375,N_7853,N_7911);
and U8376 (N_8376,N_7413,N_7184);
or U8377 (N_8377,N_7964,N_7547);
nor U8378 (N_8378,N_7553,N_7997);
and U8379 (N_8379,N_7539,N_7095);
nand U8380 (N_8380,N_7274,N_7357);
nor U8381 (N_8381,N_7860,N_7955);
nand U8382 (N_8382,N_7059,N_7046);
nand U8383 (N_8383,N_7948,N_7429);
nand U8384 (N_8384,N_7201,N_7801);
nor U8385 (N_8385,N_7733,N_7577);
nand U8386 (N_8386,N_7782,N_7390);
nand U8387 (N_8387,N_7406,N_7311);
or U8388 (N_8388,N_7224,N_7015);
nand U8389 (N_8389,N_7327,N_7808);
nand U8390 (N_8390,N_7890,N_7585);
or U8391 (N_8391,N_7127,N_7929);
or U8392 (N_8392,N_7543,N_7599);
or U8393 (N_8393,N_7588,N_7722);
nor U8394 (N_8394,N_7332,N_7778);
or U8395 (N_8395,N_7835,N_7221);
or U8396 (N_8396,N_7917,N_7049);
nor U8397 (N_8397,N_7464,N_7985);
nand U8398 (N_8398,N_7245,N_7467);
xor U8399 (N_8399,N_7659,N_7153);
xor U8400 (N_8400,N_7707,N_7880);
and U8401 (N_8401,N_7454,N_7407);
nand U8402 (N_8402,N_7428,N_7518);
and U8403 (N_8403,N_7627,N_7685);
or U8404 (N_8404,N_7081,N_7167);
nor U8405 (N_8405,N_7780,N_7176);
or U8406 (N_8406,N_7702,N_7297);
and U8407 (N_8407,N_7636,N_7750);
or U8408 (N_8408,N_7304,N_7857);
or U8409 (N_8409,N_7841,N_7048);
nor U8410 (N_8410,N_7388,N_7701);
nor U8411 (N_8411,N_7517,N_7333);
nor U8412 (N_8412,N_7017,N_7921);
or U8413 (N_8413,N_7103,N_7075);
or U8414 (N_8414,N_7171,N_7344);
or U8415 (N_8415,N_7300,N_7524);
nor U8416 (N_8416,N_7609,N_7206);
and U8417 (N_8417,N_7179,N_7531);
nand U8418 (N_8418,N_7259,N_7145);
nand U8419 (N_8419,N_7905,N_7119);
nor U8420 (N_8420,N_7285,N_7640);
xor U8421 (N_8421,N_7815,N_7792);
nor U8422 (N_8422,N_7354,N_7842);
nand U8423 (N_8423,N_7271,N_7142);
nor U8424 (N_8424,N_7896,N_7996);
nand U8425 (N_8425,N_7724,N_7365);
xnor U8426 (N_8426,N_7047,N_7235);
and U8427 (N_8427,N_7721,N_7073);
nor U8428 (N_8428,N_7884,N_7537);
and U8429 (N_8429,N_7806,N_7247);
nor U8430 (N_8430,N_7871,N_7907);
and U8431 (N_8431,N_7809,N_7825);
nor U8432 (N_8432,N_7262,N_7892);
nor U8433 (N_8433,N_7487,N_7822);
and U8434 (N_8434,N_7399,N_7821);
nand U8435 (N_8435,N_7675,N_7471);
nand U8436 (N_8436,N_7749,N_7560);
and U8437 (N_8437,N_7904,N_7774);
or U8438 (N_8438,N_7362,N_7353);
nand U8439 (N_8439,N_7504,N_7922);
and U8440 (N_8440,N_7820,N_7699);
nand U8441 (N_8441,N_7121,N_7990);
and U8442 (N_8442,N_7438,N_7276);
or U8443 (N_8443,N_7175,N_7367);
nor U8444 (N_8444,N_7409,N_7449);
or U8445 (N_8445,N_7019,N_7587);
and U8446 (N_8446,N_7355,N_7595);
xor U8447 (N_8447,N_7555,N_7408);
and U8448 (N_8448,N_7554,N_7797);
and U8449 (N_8449,N_7720,N_7089);
or U8450 (N_8450,N_7616,N_7148);
and U8451 (N_8451,N_7281,N_7202);
or U8452 (N_8452,N_7269,N_7173);
nor U8453 (N_8453,N_7150,N_7436);
nor U8454 (N_8454,N_7800,N_7980);
nor U8455 (N_8455,N_7491,N_7265);
or U8456 (N_8456,N_7604,N_7781);
xor U8457 (N_8457,N_7485,N_7849);
and U8458 (N_8458,N_7325,N_7266);
and U8459 (N_8459,N_7065,N_7790);
or U8460 (N_8460,N_7624,N_7949);
and U8461 (N_8461,N_7976,N_7198);
xnor U8462 (N_8462,N_7966,N_7062);
nand U8463 (N_8463,N_7433,N_7231);
and U8464 (N_8464,N_7558,N_7927);
or U8465 (N_8465,N_7397,N_7590);
or U8466 (N_8466,N_7054,N_7233);
and U8467 (N_8467,N_7649,N_7417);
xnor U8468 (N_8468,N_7674,N_7895);
xor U8469 (N_8469,N_7529,N_7496);
nor U8470 (N_8470,N_7829,N_7615);
nand U8471 (N_8471,N_7591,N_7133);
nand U8472 (N_8472,N_7920,N_7032);
or U8473 (N_8473,N_7729,N_7987);
nand U8474 (N_8474,N_7382,N_7596);
and U8475 (N_8475,N_7601,N_7837);
or U8476 (N_8476,N_7068,N_7755);
xor U8477 (N_8477,N_7294,N_7626);
or U8478 (N_8478,N_7082,N_7779);
xnor U8479 (N_8479,N_7277,N_7316);
and U8480 (N_8480,N_7149,N_7767);
and U8481 (N_8481,N_7490,N_7084);
nor U8482 (N_8482,N_7866,N_7258);
and U8483 (N_8483,N_7163,N_7473);
or U8484 (N_8484,N_7689,N_7392);
and U8485 (N_8485,N_7530,N_7561);
nand U8486 (N_8486,N_7506,N_7100);
nand U8487 (N_8487,N_7589,N_7480);
xnor U8488 (N_8488,N_7501,N_7151);
or U8489 (N_8489,N_7396,N_7330);
nand U8490 (N_8490,N_7935,N_7144);
and U8491 (N_8491,N_7611,N_7292);
nor U8492 (N_8492,N_7282,N_7786);
or U8493 (N_8493,N_7470,N_7623);
or U8494 (N_8494,N_7975,N_7284);
nand U8495 (N_8495,N_7170,N_7308);
or U8496 (N_8496,N_7338,N_7034);
and U8497 (N_8497,N_7883,N_7583);
or U8498 (N_8498,N_7273,N_7745);
nand U8499 (N_8499,N_7637,N_7421);
nand U8500 (N_8500,N_7156,N_7675);
or U8501 (N_8501,N_7674,N_7736);
nor U8502 (N_8502,N_7519,N_7342);
xor U8503 (N_8503,N_7003,N_7736);
nand U8504 (N_8504,N_7960,N_7086);
xor U8505 (N_8505,N_7367,N_7977);
nor U8506 (N_8506,N_7788,N_7137);
nor U8507 (N_8507,N_7616,N_7433);
nor U8508 (N_8508,N_7905,N_7305);
nand U8509 (N_8509,N_7027,N_7973);
or U8510 (N_8510,N_7326,N_7524);
nand U8511 (N_8511,N_7292,N_7178);
nor U8512 (N_8512,N_7060,N_7988);
and U8513 (N_8513,N_7989,N_7933);
and U8514 (N_8514,N_7983,N_7217);
nand U8515 (N_8515,N_7174,N_7575);
and U8516 (N_8516,N_7939,N_7728);
nand U8517 (N_8517,N_7305,N_7475);
nand U8518 (N_8518,N_7241,N_7739);
nor U8519 (N_8519,N_7640,N_7171);
xnor U8520 (N_8520,N_7385,N_7280);
nor U8521 (N_8521,N_7145,N_7012);
and U8522 (N_8522,N_7703,N_7828);
xnor U8523 (N_8523,N_7332,N_7261);
nand U8524 (N_8524,N_7205,N_7618);
or U8525 (N_8525,N_7082,N_7961);
nor U8526 (N_8526,N_7084,N_7252);
nand U8527 (N_8527,N_7561,N_7302);
xor U8528 (N_8528,N_7391,N_7579);
nand U8529 (N_8529,N_7706,N_7245);
and U8530 (N_8530,N_7685,N_7000);
xnor U8531 (N_8531,N_7774,N_7913);
nand U8532 (N_8532,N_7187,N_7200);
and U8533 (N_8533,N_7284,N_7620);
xnor U8534 (N_8534,N_7832,N_7553);
nor U8535 (N_8535,N_7950,N_7810);
and U8536 (N_8536,N_7902,N_7781);
and U8537 (N_8537,N_7418,N_7956);
or U8538 (N_8538,N_7550,N_7093);
nand U8539 (N_8539,N_7611,N_7963);
nor U8540 (N_8540,N_7224,N_7104);
nand U8541 (N_8541,N_7848,N_7078);
nand U8542 (N_8542,N_7788,N_7697);
nand U8543 (N_8543,N_7641,N_7194);
or U8544 (N_8544,N_7806,N_7574);
nor U8545 (N_8545,N_7280,N_7473);
and U8546 (N_8546,N_7689,N_7740);
nand U8547 (N_8547,N_7018,N_7332);
xnor U8548 (N_8548,N_7143,N_7192);
nor U8549 (N_8549,N_7455,N_7938);
nor U8550 (N_8550,N_7577,N_7963);
and U8551 (N_8551,N_7572,N_7480);
nand U8552 (N_8552,N_7052,N_7873);
or U8553 (N_8553,N_7791,N_7442);
nand U8554 (N_8554,N_7141,N_7953);
or U8555 (N_8555,N_7190,N_7010);
and U8556 (N_8556,N_7784,N_7283);
or U8557 (N_8557,N_7864,N_7247);
nand U8558 (N_8558,N_7919,N_7098);
nor U8559 (N_8559,N_7293,N_7405);
nor U8560 (N_8560,N_7040,N_7194);
xor U8561 (N_8561,N_7563,N_7738);
and U8562 (N_8562,N_7737,N_7085);
nor U8563 (N_8563,N_7672,N_7063);
nand U8564 (N_8564,N_7305,N_7295);
and U8565 (N_8565,N_7784,N_7191);
nor U8566 (N_8566,N_7865,N_7217);
xor U8567 (N_8567,N_7060,N_7927);
xor U8568 (N_8568,N_7102,N_7169);
or U8569 (N_8569,N_7611,N_7219);
xnor U8570 (N_8570,N_7399,N_7126);
nand U8571 (N_8571,N_7477,N_7290);
nor U8572 (N_8572,N_7220,N_7027);
and U8573 (N_8573,N_7510,N_7707);
nor U8574 (N_8574,N_7283,N_7191);
or U8575 (N_8575,N_7410,N_7764);
xor U8576 (N_8576,N_7066,N_7185);
or U8577 (N_8577,N_7501,N_7569);
and U8578 (N_8578,N_7210,N_7259);
xnor U8579 (N_8579,N_7542,N_7760);
nor U8580 (N_8580,N_7479,N_7329);
and U8581 (N_8581,N_7991,N_7175);
nor U8582 (N_8582,N_7716,N_7560);
nor U8583 (N_8583,N_7039,N_7605);
or U8584 (N_8584,N_7375,N_7010);
and U8585 (N_8585,N_7843,N_7162);
or U8586 (N_8586,N_7308,N_7607);
or U8587 (N_8587,N_7895,N_7133);
and U8588 (N_8588,N_7991,N_7204);
nand U8589 (N_8589,N_7349,N_7324);
nor U8590 (N_8590,N_7346,N_7826);
nand U8591 (N_8591,N_7606,N_7714);
or U8592 (N_8592,N_7800,N_7601);
and U8593 (N_8593,N_7608,N_7620);
nand U8594 (N_8594,N_7463,N_7365);
xor U8595 (N_8595,N_7931,N_7675);
nand U8596 (N_8596,N_7904,N_7290);
and U8597 (N_8597,N_7839,N_7709);
and U8598 (N_8598,N_7209,N_7083);
and U8599 (N_8599,N_7474,N_7138);
nand U8600 (N_8600,N_7277,N_7847);
nor U8601 (N_8601,N_7766,N_7122);
nand U8602 (N_8602,N_7035,N_7133);
nor U8603 (N_8603,N_7709,N_7174);
and U8604 (N_8604,N_7596,N_7388);
and U8605 (N_8605,N_7512,N_7122);
or U8606 (N_8606,N_7271,N_7928);
nor U8607 (N_8607,N_7682,N_7523);
xnor U8608 (N_8608,N_7962,N_7932);
nor U8609 (N_8609,N_7109,N_7788);
nor U8610 (N_8610,N_7921,N_7501);
nand U8611 (N_8611,N_7268,N_7989);
and U8612 (N_8612,N_7517,N_7040);
nor U8613 (N_8613,N_7323,N_7705);
and U8614 (N_8614,N_7955,N_7086);
nand U8615 (N_8615,N_7496,N_7761);
nand U8616 (N_8616,N_7329,N_7974);
or U8617 (N_8617,N_7864,N_7976);
and U8618 (N_8618,N_7091,N_7243);
xor U8619 (N_8619,N_7687,N_7285);
nand U8620 (N_8620,N_7436,N_7356);
or U8621 (N_8621,N_7533,N_7476);
xnor U8622 (N_8622,N_7143,N_7895);
nand U8623 (N_8623,N_7165,N_7423);
nand U8624 (N_8624,N_7405,N_7831);
or U8625 (N_8625,N_7257,N_7689);
and U8626 (N_8626,N_7368,N_7196);
nor U8627 (N_8627,N_7826,N_7815);
and U8628 (N_8628,N_7193,N_7357);
and U8629 (N_8629,N_7734,N_7582);
nor U8630 (N_8630,N_7398,N_7736);
or U8631 (N_8631,N_7716,N_7131);
nand U8632 (N_8632,N_7375,N_7344);
xor U8633 (N_8633,N_7110,N_7067);
and U8634 (N_8634,N_7616,N_7546);
xnor U8635 (N_8635,N_7891,N_7227);
nor U8636 (N_8636,N_7783,N_7383);
or U8637 (N_8637,N_7893,N_7253);
and U8638 (N_8638,N_7424,N_7319);
and U8639 (N_8639,N_7160,N_7078);
nor U8640 (N_8640,N_7232,N_7972);
nand U8641 (N_8641,N_7282,N_7318);
and U8642 (N_8642,N_7261,N_7323);
or U8643 (N_8643,N_7229,N_7898);
nor U8644 (N_8644,N_7877,N_7750);
nand U8645 (N_8645,N_7837,N_7926);
nor U8646 (N_8646,N_7723,N_7860);
xor U8647 (N_8647,N_7944,N_7469);
and U8648 (N_8648,N_7367,N_7097);
or U8649 (N_8649,N_7182,N_7860);
and U8650 (N_8650,N_7012,N_7449);
nor U8651 (N_8651,N_7195,N_7479);
and U8652 (N_8652,N_7782,N_7983);
nor U8653 (N_8653,N_7209,N_7667);
or U8654 (N_8654,N_7305,N_7411);
and U8655 (N_8655,N_7405,N_7066);
nor U8656 (N_8656,N_7841,N_7451);
or U8657 (N_8657,N_7516,N_7500);
or U8658 (N_8658,N_7277,N_7801);
xor U8659 (N_8659,N_7046,N_7029);
or U8660 (N_8660,N_7259,N_7323);
nand U8661 (N_8661,N_7329,N_7138);
or U8662 (N_8662,N_7058,N_7269);
xor U8663 (N_8663,N_7969,N_7415);
nand U8664 (N_8664,N_7646,N_7186);
or U8665 (N_8665,N_7783,N_7603);
and U8666 (N_8666,N_7042,N_7069);
and U8667 (N_8667,N_7519,N_7299);
nor U8668 (N_8668,N_7462,N_7849);
and U8669 (N_8669,N_7317,N_7279);
or U8670 (N_8670,N_7786,N_7413);
or U8671 (N_8671,N_7937,N_7523);
and U8672 (N_8672,N_7757,N_7346);
nor U8673 (N_8673,N_7486,N_7807);
nor U8674 (N_8674,N_7941,N_7619);
and U8675 (N_8675,N_7170,N_7552);
and U8676 (N_8676,N_7860,N_7229);
and U8677 (N_8677,N_7434,N_7834);
xnor U8678 (N_8678,N_7422,N_7524);
xnor U8679 (N_8679,N_7208,N_7466);
or U8680 (N_8680,N_7720,N_7668);
nor U8681 (N_8681,N_7792,N_7951);
and U8682 (N_8682,N_7506,N_7201);
or U8683 (N_8683,N_7904,N_7995);
nor U8684 (N_8684,N_7275,N_7829);
nor U8685 (N_8685,N_7012,N_7771);
or U8686 (N_8686,N_7782,N_7221);
and U8687 (N_8687,N_7268,N_7914);
or U8688 (N_8688,N_7791,N_7725);
and U8689 (N_8689,N_7642,N_7829);
nand U8690 (N_8690,N_7249,N_7524);
xnor U8691 (N_8691,N_7254,N_7015);
or U8692 (N_8692,N_7164,N_7917);
nor U8693 (N_8693,N_7930,N_7768);
or U8694 (N_8694,N_7544,N_7463);
nand U8695 (N_8695,N_7999,N_7115);
nand U8696 (N_8696,N_7537,N_7327);
or U8697 (N_8697,N_7208,N_7515);
or U8698 (N_8698,N_7927,N_7687);
nor U8699 (N_8699,N_7510,N_7465);
nand U8700 (N_8700,N_7551,N_7577);
or U8701 (N_8701,N_7320,N_7359);
nand U8702 (N_8702,N_7843,N_7082);
and U8703 (N_8703,N_7225,N_7074);
and U8704 (N_8704,N_7250,N_7367);
nand U8705 (N_8705,N_7373,N_7544);
or U8706 (N_8706,N_7546,N_7470);
nand U8707 (N_8707,N_7459,N_7503);
nor U8708 (N_8708,N_7556,N_7342);
nand U8709 (N_8709,N_7408,N_7789);
nor U8710 (N_8710,N_7737,N_7072);
nor U8711 (N_8711,N_7844,N_7653);
and U8712 (N_8712,N_7782,N_7020);
nand U8713 (N_8713,N_7736,N_7453);
nor U8714 (N_8714,N_7558,N_7594);
and U8715 (N_8715,N_7391,N_7016);
xnor U8716 (N_8716,N_7492,N_7054);
nand U8717 (N_8717,N_7175,N_7951);
nand U8718 (N_8718,N_7317,N_7060);
and U8719 (N_8719,N_7055,N_7874);
nand U8720 (N_8720,N_7870,N_7003);
nand U8721 (N_8721,N_7915,N_7050);
or U8722 (N_8722,N_7762,N_7406);
nand U8723 (N_8723,N_7441,N_7257);
and U8724 (N_8724,N_7793,N_7105);
nor U8725 (N_8725,N_7264,N_7276);
nand U8726 (N_8726,N_7126,N_7505);
nand U8727 (N_8727,N_7516,N_7028);
nand U8728 (N_8728,N_7459,N_7980);
or U8729 (N_8729,N_7565,N_7980);
nand U8730 (N_8730,N_7917,N_7316);
nor U8731 (N_8731,N_7556,N_7089);
xor U8732 (N_8732,N_7523,N_7218);
nor U8733 (N_8733,N_7193,N_7158);
xor U8734 (N_8734,N_7217,N_7995);
and U8735 (N_8735,N_7344,N_7024);
or U8736 (N_8736,N_7281,N_7337);
xnor U8737 (N_8737,N_7146,N_7652);
or U8738 (N_8738,N_7589,N_7603);
nand U8739 (N_8739,N_7869,N_7360);
or U8740 (N_8740,N_7783,N_7968);
or U8741 (N_8741,N_7680,N_7106);
nand U8742 (N_8742,N_7677,N_7804);
nor U8743 (N_8743,N_7255,N_7522);
nor U8744 (N_8744,N_7016,N_7484);
xor U8745 (N_8745,N_7442,N_7934);
and U8746 (N_8746,N_7091,N_7005);
and U8747 (N_8747,N_7466,N_7845);
or U8748 (N_8748,N_7946,N_7604);
nor U8749 (N_8749,N_7696,N_7693);
and U8750 (N_8750,N_7113,N_7739);
xnor U8751 (N_8751,N_7653,N_7073);
nand U8752 (N_8752,N_7831,N_7724);
nand U8753 (N_8753,N_7388,N_7896);
nand U8754 (N_8754,N_7475,N_7684);
nor U8755 (N_8755,N_7202,N_7758);
or U8756 (N_8756,N_7145,N_7905);
nand U8757 (N_8757,N_7695,N_7024);
or U8758 (N_8758,N_7696,N_7422);
and U8759 (N_8759,N_7517,N_7142);
nor U8760 (N_8760,N_7480,N_7189);
and U8761 (N_8761,N_7053,N_7345);
nor U8762 (N_8762,N_7486,N_7653);
nor U8763 (N_8763,N_7745,N_7888);
xnor U8764 (N_8764,N_7144,N_7401);
or U8765 (N_8765,N_7416,N_7351);
xor U8766 (N_8766,N_7106,N_7485);
or U8767 (N_8767,N_7795,N_7516);
nand U8768 (N_8768,N_7630,N_7598);
or U8769 (N_8769,N_7705,N_7802);
or U8770 (N_8770,N_7961,N_7603);
xor U8771 (N_8771,N_7060,N_7511);
nand U8772 (N_8772,N_7675,N_7710);
or U8773 (N_8773,N_7747,N_7724);
nor U8774 (N_8774,N_7460,N_7687);
or U8775 (N_8775,N_7278,N_7075);
or U8776 (N_8776,N_7142,N_7683);
or U8777 (N_8777,N_7304,N_7702);
and U8778 (N_8778,N_7545,N_7346);
nor U8779 (N_8779,N_7585,N_7468);
or U8780 (N_8780,N_7570,N_7549);
or U8781 (N_8781,N_7205,N_7638);
nor U8782 (N_8782,N_7382,N_7591);
and U8783 (N_8783,N_7482,N_7126);
nor U8784 (N_8784,N_7355,N_7006);
or U8785 (N_8785,N_7078,N_7900);
and U8786 (N_8786,N_7807,N_7041);
or U8787 (N_8787,N_7848,N_7147);
and U8788 (N_8788,N_7155,N_7615);
nand U8789 (N_8789,N_7219,N_7729);
nand U8790 (N_8790,N_7370,N_7654);
nand U8791 (N_8791,N_7264,N_7844);
xnor U8792 (N_8792,N_7758,N_7323);
and U8793 (N_8793,N_7887,N_7298);
nor U8794 (N_8794,N_7015,N_7248);
nor U8795 (N_8795,N_7471,N_7008);
nor U8796 (N_8796,N_7332,N_7674);
or U8797 (N_8797,N_7277,N_7172);
and U8798 (N_8798,N_7329,N_7259);
xnor U8799 (N_8799,N_7931,N_7715);
or U8800 (N_8800,N_7307,N_7636);
and U8801 (N_8801,N_7348,N_7167);
or U8802 (N_8802,N_7488,N_7716);
nor U8803 (N_8803,N_7876,N_7041);
and U8804 (N_8804,N_7096,N_7210);
and U8805 (N_8805,N_7770,N_7097);
xor U8806 (N_8806,N_7273,N_7526);
and U8807 (N_8807,N_7150,N_7455);
nand U8808 (N_8808,N_7265,N_7267);
nor U8809 (N_8809,N_7365,N_7347);
xor U8810 (N_8810,N_7073,N_7011);
nor U8811 (N_8811,N_7351,N_7448);
nand U8812 (N_8812,N_7058,N_7770);
nand U8813 (N_8813,N_7755,N_7355);
or U8814 (N_8814,N_7696,N_7299);
nor U8815 (N_8815,N_7376,N_7232);
and U8816 (N_8816,N_7558,N_7385);
nand U8817 (N_8817,N_7896,N_7958);
and U8818 (N_8818,N_7518,N_7564);
nor U8819 (N_8819,N_7601,N_7373);
or U8820 (N_8820,N_7797,N_7673);
nor U8821 (N_8821,N_7386,N_7488);
nand U8822 (N_8822,N_7503,N_7864);
and U8823 (N_8823,N_7933,N_7155);
and U8824 (N_8824,N_7256,N_7410);
xor U8825 (N_8825,N_7534,N_7708);
nor U8826 (N_8826,N_7399,N_7200);
nor U8827 (N_8827,N_7041,N_7515);
or U8828 (N_8828,N_7688,N_7438);
and U8829 (N_8829,N_7607,N_7939);
nor U8830 (N_8830,N_7191,N_7105);
and U8831 (N_8831,N_7291,N_7063);
nand U8832 (N_8832,N_7559,N_7243);
nand U8833 (N_8833,N_7238,N_7432);
and U8834 (N_8834,N_7786,N_7621);
nand U8835 (N_8835,N_7256,N_7529);
nor U8836 (N_8836,N_7101,N_7394);
and U8837 (N_8837,N_7698,N_7507);
or U8838 (N_8838,N_7835,N_7114);
nor U8839 (N_8839,N_7400,N_7162);
or U8840 (N_8840,N_7174,N_7930);
nand U8841 (N_8841,N_7858,N_7992);
nor U8842 (N_8842,N_7355,N_7032);
nor U8843 (N_8843,N_7365,N_7606);
or U8844 (N_8844,N_7777,N_7157);
and U8845 (N_8845,N_7525,N_7075);
nand U8846 (N_8846,N_7091,N_7143);
nor U8847 (N_8847,N_7024,N_7902);
nand U8848 (N_8848,N_7357,N_7235);
xnor U8849 (N_8849,N_7000,N_7756);
and U8850 (N_8850,N_7396,N_7008);
nor U8851 (N_8851,N_7833,N_7290);
nor U8852 (N_8852,N_7126,N_7907);
nor U8853 (N_8853,N_7572,N_7524);
and U8854 (N_8854,N_7407,N_7100);
and U8855 (N_8855,N_7632,N_7513);
nor U8856 (N_8856,N_7511,N_7786);
nor U8857 (N_8857,N_7255,N_7450);
nand U8858 (N_8858,N_7403,N_7127);
nand U8859 (N_8859,N_7928,N_7550);
and U8860 (N_8860,N_7175,N_7100);
nor U8861 (N_8861,N_7160,N_7569);
nand U8862 (N_8862,N_7087,N_7078);
nand U8863 (N_8863,N_7068,N_7524);
and U8864 (N_8864,N_7994,N_7001);
or U8865 (N_8865,N_7359,N_7647);
nand U8866 (N_8866,N_7303,N_7117);
or U8867 (N_8867,N_7536,N_7681);
xnor U8868 (N_8868,N_7726,N_7348);
and U8869 (N_8869,N_7287,N_7475);
and U8870 (N_8870,N_7853,N_7624);
xnor U8871 (N_8871,N_7168,N_7836);
or U8872 (N_8872,N_7849,N_7222);
or U8873 (N_8873,N_7398,N_7135);
and U8874 (N_8874,N_7296,N_7022);
or U8875 (N_8875,N_7258,N_7679);
or U8876 (N_8876,N_7852,N_7648);
and U8877 (N_8877,N_7350,N_7283);
and U8878 (N_8878,N_7053,N_7237);
nor U8879 (N_8879,N_7793,N_7468);
xnor U8880 (N_8880,N_7006,N_7328);
nand U8881 (N_8881,N_7943,N_7176);
and U8882 (N_8882,N_7557,N_7942);
nand U8883 (N_8883,N_7301,N_7072);
nor U8884 (N_8884,N_7541,N_7707);
xor U8885 (N_8885,N_7249,N_7750);
or U8886 (N_8886,N_7641,N_7452);
nor U8887 (N_8887,N_7716,N_7542);
nand U8888 (N_8888,N_7562,N_7649);
and U8889 (N_8889,N_7466,N_7936);
nand U8890 (N_8890,N_7987,N_7993);
nand U8891 (N_8891,N_7618,N_7711);
nand U8892 (N_8892,N_7192,N_7075);
and U8893 (N_8893,N_7326,N_7804);
nand U8894 (N_8894,N_7162,N_7255);
and U8895 (N_8895,N_7422,N_7023);
or U8896 (N_8896,N_7364,N_7194);
nand U8897 (N_8897,N_7232,N_7843);
nand U8898 (N_8898,N_7745,N_7170);
and U8899 (N_8899,N_7193,N_7461);
nor U8900 (N_8900,N_7167,N_7306);
and U8901 (N_8901,N_7985,N_7651);
xnor U8902 (N_8902,N_7246,N_7734);
or U8903 (N_8903,N_7390,N_7617);
and U8904 (N_8904,N_7876,N_7207);
or U8905 (N_8905,N_7907,N_7471);
or U8906 (N_8906,N_7074,N_7748);
and U8907 (N_8907,N_7536,N_7144);
xor U8908 (N_8908,N_7681,N_7788);
xnor U8909 (N_8909,N_7184,N_7822);
and U8910 (N_8910,N_7448,N_7470);
nand U8911 (N_8911,N_7692,N_7894);
xor U8912 (N_8912,N_7942,N_7859);
and U8913 (N_8913,N_7324,N_7610);
or U8914 (N_8914,N_7538,N_7290);
nand U8915 (N_8915,N_7908,N_7304);
nand U8916 (N_8916,N_7955,N_7810);
nand U8917 (N_8917,N_7035,N_7310);
nand U8918 (N_8918,N_7466,N_7894);
xor U8919 (N_8919,N_7175,N_7998);
or U8920 (N_8920,N_7484,N_7651);
xnor U8921 (N_8921,N_7501,N_7829);
and U8922 (N_8922,N_7839,N_7716);
and U8923 (N_8923,N_7355,N_7579);
or U8924 (N_8924,N_7543,N_7003);
and U8925 (N_8925,N_7224,N_7809);
nor U8926 (N_8926,N_7456,N_7021);
or U8927 (N_8927,N_7760,N_7304);
nor U8928 (N_8928,N_7277,N_7100);
and U8929 (N_8929,N_7626,N_7008);
nand U8930 (N_8930,N_7333,N_7477);
nand U8931 (N_8931,N_7117,N_7036);
or U8932 (N_8932,N_7201,N_7267);
or U8933 (N_8933,N_7497,N_7470);
or U8934 (N_8934,N_7300,N_7502);
nand U8935 (N_8935,N_7245,N_7765);
or U8936 (N_8936,N_7819,N_7042);
nand U8937 (N_8937,N_7610,N_7579);
and U8938 (N_8938,N_7025,N_7116);
or U8939 (N_8939,N_7703,N_7058);
and U8940 (N_8940,N_7397,N_7293);
or U8941 (N_8941,N_7125,N_7405);
xnor U8942 (N_8942,N_7464,N_7762);
and U8943 (N_8943,N_7653,N_7227);
or U8944 (N_8944,N_7076,N_7394);
or U8945 (N_8945,N_7075,N_7357);
xnor U8946 (N_8946,N_7077,N_7198);
nand U8947 (N_8947,N_7917,N_7247);
xnor U8948 (N_8948,N_7348,N_7749);
nand U8949 (N_8949,N_7491,N_7017);
and U8950 (N_8950,N_7086,N_7071);
or U8951 (N_8951,N_7298,N_7535);
nand U8952 (N_8952,N_7804,N_7178);
nand U8953 (N_8953,N_7085,N_7619);
nor U8954 (N_8954,N_7514,N_7655);
and U8955 (N_8955,N_7266,N_7803);
nand U8956 (N_8956,N_7690,N_7104);
nand U8957 (N_8957,N_7396,N_7201);
and U8958 (N_8958,N_7691,N_7131);
nand U8959 (N_8959,N_7677,N_7835);
and U8960 (N_8960,N_7934,N_7498);
and U8961 (N_8961,N_7422,N_7027);
nand U8962 (N_8962,N_7287,N_7658);
nor U8963 (N_8963,N_7626,N_7982);
nor U8964 (N_8964,N_7589,N_7126);
nor U8965 (N_8965,N_7083,N_7316);
xnor U8966 (N_8966,N_7863,N_7912);
or U8967 (N_8967,N_7206,N_7762);
nand U8968 (N_8968,N_7989,N_7779);
nor U8969 (N_8969,N_7818,N_7641);
nand U8970 (N_8970,N_7619,N_7716);
nor U8971 (N_8971,N_7700,N_7290);
and U8972 (N_8972,N_7442,N_7414);
xnor U8973 (N_8973,N_7447,N_7642);
nor U8974 (N_8974,N_7350,N_7857);
nand U8975 (N_8975,N_7173,N_7505);
and U8976 (N_8976,N_7257,N_7605);
nand U8977 (N_8977,N_7031,N_7762);
and U8978 (N_8978,N_7569,N_7206);
nand U8979 (N_8979,N_7060,N_7004);
xnor U8980 (N_8980,N_7575,N_7579);
nor U8981 (N_8981,N_7510,N_7191);
or U8982 (N_8982,N_7257,N_7345);
or U8983 (N_8983,N_7964,N_7036);
nor U8984 (N_8984,N_7639,N_7287);
nor U8985 (N_8985,N_7474,N_7166);
xnor U8986 (N_8986,N_7726,N_7203);
or U8987 (N_8987,N_7672,N_7154);
and U8988 (N_8988,N_7384,N_7640);
and U8989 (N_8989,N_7015,N_7463);
or U8990 (N_8990,N_7837,N_7813);
or U8991 (N_8991,N_7622,N_7430);
nand U8992 (N_8992,N_7165,N_7753);
nor U8993 (N_8993,N_7792,N_7444);
and U8994 (N_8994,N_7342,N_7520);
nor U8995 (N_8995,N_7565,N_7363);
nand U8996 (N_8996,N_7581,N_7074);
and U8997 (N_8997,N_7983,N_7106);
or U8998 (N_8998,N_7862,N_7414);
and U8999 (N_8999,N_7405,N_7096);
nor U9000 (N_9000,N_8900,N_8455);
nor U9001 (N_9001,N_8906,N_8006);
and U9002 (N_9002,N_8484,N_8185);
and U9003 (N_9003,N_8251,N_8406);
xor U9004 (N_9004,N_8654,N_8687);
or U9005 (N_9005,N_8367,N_8511);
nor U9006 (N_9006,N_8239,N_8273);
or U9007 (N_9007,N_8005,N_8163);
nor U9008 (N_9008,N_8076,N_8816);
nand U9009 (N_9009,N_8299,N_8690);
xnor U9010 (N_9010,N_8675,N_8033);
nand U9011 (N_9011,N_8392,N_8446);
nand U9012 (N_9012,N_8674,N_8193);
or U9013 (N_9013,N_8361,N_8994);
and U9014 (N_9014,N_8398,N_8089);
nor U9015 (N_9015,N_8716,N_8826);
and U9016 (N_9016,N_8257,N_8054);
and U9017 (N_9017,N_8757,N_8551);
and U9018 (N_9018,N_8669,N_8042);
or U9019 (N_9019,N_8466,N_8195);
or U9020 (N_9020,N_8104,N_8268);
and U9021 (N_9021,N_8187,N_8979);
or U9022 (N_9022,N_8748,N_8682);
nand U9023 (N_9023,N_8937,N_8001);
nand U9024 (N_9024,N_8055,N_8323);
and U9025 (N_9025,N_8493,N_8920);
or U9026 (N_9026,N_8766,N_8798);
nand U9027 (N_9027,N_8604,N_8307);
or U9028 (N_9028,N_8987,N_8708);
or U9029 (N_9029,N_8717,N_8694);
nor U9030 (N_9030,N_8837,N_8784);
or U9031 (N_9031,N_8772,N_8767);
and U9032 (N_9032,N_8890,N_8732);
nand U9033 (N_9033,N_8123,N_8616);
or U9034 (N_9034,N_8939,N_8754);
or U9035 (N_9035,N_8894,N_8197);
or U9036 (N_9036,N_8934,N_8714);
nand U9037 (N_9037,N_8243,N_8339);
or U9038 (N_9038,N_8968,N_8643);
nand U9039 (N_9039,N_8014,N_8788);
xnor U9040 (N_9040,N_8603,N_8085);
nand U9041 (N_9041,N_8366,N_8018);
xnor U9042 (N_9042,N_8561,N_8067);
and U9043 (N_9043,N_8293,N_8094);
xnor U9044 (N_9044,N_8335,N_8061);
nor U9045 (N_9045,N_8636,N_8324);
or U9046 (N_9046,N_8809,N_8501);
nand U9047 (N_9047,N_8030,N_8091);
nor U9048 (N_9048,N_8681,N_8962);
and U9049 (N_9049,N_8560,N_8581);
nand U9050 (N_9050,N_8262,N_8146);
or U9051 (N_9051,N_8918,N_8200);
nand U9052 (N_9052,N_8778,N_8993);
or U9053 (N_9053,N_8388,N_8519);
nor U9054 (N_9054,N_8700,N_8638);
and U9055 (N_9055,N_8562,N_8420);
nand U9056 (N_9056,N_8469,N_8238);
nor U9057 (N_9057,N_8723,N_8851);
nor U9058 (N_9058,N_8095,N_8384);
and U9059 (N_9059,N_8096,N_8743);
and U9060 (N_9060,N_8342,N_8397);
nor U9061 (N_9061,N_8641,N_8426);
nand U9062 (N_9062,N_8995,N_8556);
nor U9063 (N_9063,N_8491,N_8627);
and U9064 (N_9064,N_8751,N_8242);
nor U9065 (N_9065,N_8044,N_8752);
nand U9066 (N_9066,N_8790,N_8269);
and U9067 (N_9067,N_8571,N_8023);
and U9068 (N_9068,N_8407,N_8348);
and U9069 (N_9069,N_8969,N_8341);
nor U9070 (N_9070,N_8494,N_8222);
or U9071 (N_9071,N_8924,N_8564);
or U9072 (N_9072,N_8905,N_8136);
nand U9073 (N_9073,N_8530,N_8219);
nor U9074 (N_9074,N_8908,N_8212);
nor U9075 (N_9075,N_8000,N_8797);
nor U9076 (N_9076,N_8165,N_8977);
nand U9077 (N_9077,N_8590,N_8775);
and U9078 (N_9078,N_8457,N_8836);
nand U9079 (N_9079,N_8409,N_8835);
and U9080 (N_9080,N_8637,N_8550);
nand U9081 (N_9081,N_8725,N_8207);
nand U9082 (N_9082,N_8921,N_8624);
and U9083 (N_9083,N_8387,N_8733);
nor U9084 (N_9084,N_8970,N_8202);
or U9085 (N_9085,N_8782,N_8761);
nor U9086 (N_9086,N_8280,N_8504);
or U9087 (N_9087,N_8133,N_8275);
nand U9088 (N_9088,N_8728,N_8451);
and U9089 (N_9089,N_8092,N_8686);
and U9090 (N_9090,N_8507,N_8959);
or U9091 (N_9091,N_8629,N_8442);
nor U9092 (N_9092,N_8319,N_8777);
or U9093 (N_9093,N_8952,N_8443);
nand U9094 (N_9094,N_8283,N_8138);
nor U9095 (N_9095,N_8325,N_8002);
nand U9096 (N_9096,N_8350,N_8810);
nor U9097 (N_9097,N_8320,N_8801);
nand U9098 (N_9098,N_8377,N_8196);
nor U9099 (N_9099,N_8660,N_8266);
or U9100 (N_9100,N_8263,N_8673);
xor U9101 (N_9101,N_8972,N_8817);
nor U9102 (N_9102,N_8763,N_8399);
nand U9103 (N_9103,N_8058,N_8218);
xnor U9104 (N_9104,N_8842,N_8359);
nand U9105 (N_9105,N_8631,N_8662);
nor U9106 (N_9106,N_8157,N_8705);
nand U9107 (N_9107,N_8247,N_8883);
or U9108 (N_9108,N_8578,N_8567);
nor U9109 (N_9109,N_8791,N_8475);
nor U9110 (N_9110,N_8227,N_8448);
or U9111 (N_9111,N_8779,N_8818);
nor U9112 (N_9112,N_8804,N_8396);
nand U9113 (N_9113,N_8431,N_8453);
and U9114 (N_9114,N_8462,N_8034);
nand U9115 (N_9115,N_8106,N_8704);
or U9116 (N_9116,N_8539,N_8346);
nand U9117 (N_9117,N_8543,N_8427);
nor U9118 (N_9118,N_8771,N_8870);
or U9119 (N_9119,N_8516,N_8614);
nor U9120 (N_9120,N_8830,N_8368);
and U9121 (N_9121,N_8984,N_8330);
and U9122 (N_9122,N_8666,N_8363);
and U9123 (N_9123,N_8711,N_8792);
or U9124 (N_9124,N_8943,N_8632);
or U9125 (N_9125,N_8486,N_8699);
nor U9126 (N_9126,N_8724,N_8132);
and U9127 (N_9127,N_8881,N_8594);
and U9128 (N_9128,N_8866,N_8355);
xor U9129 (N_9129,N_8464,N_8436);
xnor U9130 (N_9130,N_8800,N_8946);
nand U9131 (N_9131,N_8848,N_8043);
or U9132 (N_9132,N_8889,N_8070);
and U9133 (N_9133,N_8858,N_8220);
nor U9134 (N_9134,N_8011,N_8912);
nand U9135 (N_9135,N_8344,N_8620);
xnor U9136 (N_9136,N_8385,N_8260);
and U9137 (N_9137,N_8524,N_8531);
or U9138 (N_9138,N_8986,N_8031);
and U9139 (N_9139,N_8537,N_8932);
nor U9140 (N_9140,N_8973,N_8131);
nor U9141 (N_9141,N_8261,N_8615);
and U9142 (N_9142,N_8793,N_8211);
or U9143 (N_9143,N_8877,N_8819);
or U9144 (N_9144,N_8941,N_8610);
nand U9145 (N_9145,N_8608,N_8672);
xnor U9146 (N_9146,N_8419,N_8823);
and U9147 (N_9147,N_8035,N_8016);
nand U9148 (N_9148,N_8857,N_8463);
nand U9149 (N_9149,N_8843,N_8568);
or U9150 (N_9150,N_8735,N_8048);
and U9151 (N_9151,N_8471,N_8479);
and U9152 (N_9152,N_8379,N_8141);
or U9153 (N_9153,N_8671,N_8618);
or U9154 (N_9154,N_8591,N_8532);
or U9155 (N_9155,N_8100,N_8898);
nor U9156 (N_9156,N_8458,N_8508);
and U9157 (N_9157,N_8954,N_8170);
nor U9158 (N_9158,N_8529,N_8270);
or U9159 (N_9159,N_8485,N_8712);
or U9160 (N_9160,N_8884,N_8496);
and U9161 (N_9161,N_8333,N_8997);
nor U9162 (N_9162,N_8281,N_8976);
or U9163 (N_9163,N_8512,N_8116);
nor U9164 (N_9164,N_8190,N_8720);
nand U9165 (N_9165,N_8391,N_8855);
nor U9166 (N_9166,N_8580,N_8267);
and U9167 (N_9167,N_8722,N_8376);
nor U9168 (N_9168,N_8204,N_8098);
and U9169 (N_9169,N_8066,N_8520);
nand U9170 (N_9170,N_8282,N_8559);
and U9171 (N_9171,N_8421,N_8873);
nor U9172 (N_9172,N_8393,N_8037);
nor U9173 (N_9173,N_8789,N_8249);
or U9174 (N_9174,N_8923,N_8434);
xnor U9175 (N_9175,N_8910,N_8410);
xor U9176 (N_9176,N_8354,N_8670);
nand U9177 (N_9177,N_8691,N_8745);
or U9178 (N_9178,N_8533,N_8750);
xor U9179 (N_9179,N_8435,N_8483);
and U9180 (N_9180,N_8768,N_8661);
and U9181 (N_9181,N_8774,N_8130);
or U9182 (N_9182,N_8558,N_8412);
and U9183 (N_9183,N_8606,N_8360);
or U9184 (N_9184,N_8476,N_8358);
nor U9185 (N_9185,N_8780,N_8825);
and U9186 (N_9186,N_8039,N_8065);
xor U9187 (N_9187,N_8209,N_8137);
nand U9188 (N_9188,N_8981,N_8785);
and U9189 (N_9189,N_8740,N_8613);
nand U9190 (N_9190,N_8097,N_8191);
and U9191 (N_9191,N_8680,N_8689);
or U9192 (N_9192,N_8731,N_8776);
or U9193 (N_9193,N_8506,N_8549);
or U9194 (N_9194,N_8961,N_8115);
nor U9195 (N_9195,N_8080,N_8229);
or U9196 (N_9196,N_8860,N_8888);
or U9197 (N_9197,N_8237,N_8331);
or U9198 (N_9198,N_8276,N_8063);
and U9199 (N_9199,N_8235,N_8878);
nor U9200 (N_9200,N_8683,N_8566);
nand U9201 (N_9201,N_8232,N_8459);
nand U9202 (N_9202,N_8996,N_8955);
nor U9203 (N_9203,N_8916,N_8314);
or U9204 (N_9204,N_8832,N_8250);
nor U9205 (N_9205,N_8922,N_8929);
nor U9206 (N_9206,N_8153,N_8726);
and U9207 (N_9207,N_8875,N_8940);
and U9208 (N_9208,N_8022,N_8576);
and U9209 (N_9209,N_8555,N_8846);
nand U9210 (N_9210,N_8164,N_8536);
nand U9211 (N_9211,N_8893,N_8473);
and U9212 (N_9212,N_8432,N_8492);
nand U9213 (N_9213,N_8684,N_8915);
and U9214 (N_9214,N_8773,N_8667);
nor U9215 (N_9215,N_8974,N_8874);
or U9216 (N_9216,N_8167,N_8844);
nor U9217 (N_9217,N_8978,N_8381);
or U9218 (N_9218,N_8297,N_8935);
and U9219 (N_9219,N_8075,N_8862);
nand U9220 (N_9220,N_8989,N_8545);
xnor U9221 (N_9221,N_8692,N_8886);
and U9222 (N_9222,N_8659,N_8394);
nand U9223 (N_9223,N_8265,N_8600);
and U9224 (N_9224,N_8288,N_8291);
nor U9225 (N_9225,N_8872,N_8114);
nand U9226 (N_9226,N_8389,N_8719);
xor U9227 (N_9227,N_8069,N_8225);
nand U9228 (N_9228,N_8992,N_8828);
nand U9229 (N_9229,N_8272,N_8619);
nor U9230 (N_9230,N_8813,N_8152);
or U9231 (N_9231,N_8799,N_8199);
nor U9232 (N_9232,N_8839,N_8375);
or U9233 (N_9233,N_8697,N_8214);
and U9234 (N_9234,N_8327,N_8628);
nand U9235 (N_9235,N_8072,N_8701);
and U9236 (N_9236,N_8271,N_8764);
and U9237 (N_9237,N_8640,N_8944);
or U9238 (N_9238,N_8953,N_8461);
and U9239 (N_9239,N_8626,N_8605);
or U9240 (N_9240,N_8585,N_8695);
nor U9241 (N_9241,N_8621,N_8895);
nand U9242 (N_9242,N_8161,N_8885);
and U9243 (N_9243,N_8803,N_8221);
nor U9244 (N_9244,N_8429,N_8201);
or U9245 (N_9245,N_8255,N_8490);
nor U9246 (N_9246,N_8302,N_8440);
nand U9247 (N_9247,N_8447,N_8090);
nand U9248 (N_9248,N_8513,N_8181);
nand U9249 (N_9249,N_8216,N_8574);
nor U9250 (N_9250,N_8470,N_8509);
nor U9251 (N_9251,N_8706,N_8311);
nand U9252 (N_9252,N_8329,N_8166);
xor U9253 (N_9253,N_8480,N_8078);
nand U9254 (N_9254,N_8150,N_8413);
nand U9255 (N_9255,N_8967,N_8142);
nor U9256 (N_9256,N_8548,N_8821);
and U9257 (N_9257,N_8449,N_8592);
and U9258 (N_9258,N_8956,N_8403);
nand U9259 (N_9259,N_8256,N_8926);
and U9260 (N_9260,N_8254,N_8652);
or U9261 (N_9261,N_8038,N_8749);
nor U9262 (N_9262,N_8315,N_8294);
nand U9263 (N_9263,N_8059,N_8345);
xor U9264 (N_9264,N_8515,N_8685);
or U9265 (N_9265,N_8965,N_8349);
nor U9266 (N_9266,N_8032,N_8328);
or U9267 (N_9267,N_8514,N_8400);
nand U9268 (N_9268,N_8177,N_8184);
nor U9269 (N_9269,N_8815,N_8351);
nand U9270 (N_9270,N_8739,N_8373);
xnor U9271 (N_9271,N_8625,N_8126);
nand U9272 (N_9272,N_8914,N_8897);
xor U9273 (N_9273,N_8891,N_8122);
and U9274 (N_9274,N_8071,N_8084);
and U9275 (N_9275,N_8309,N_8642);
or U9276 (N_9276,N_8102,N_8390);
and U9277 (N_9277,N_8301,N_8575);
nand U9278 (N_9278,N_8964,N_8593);
nor U9279 (N_9279,N_8991,N_8057);
nor U9280 (N_9280,N_8865,N_8194);
nor U9281 (N_9281,N_8264,N_8960);
nand U9282 (N_9282,N_8430,N_8180);
and U9283 (N_9283,N_8093,N_8310);
nand U9284 (N_9284,N_8452,N_8356);
nand U9285 (N_9285,N_8824,N_8244);
nand U9286 (N_9286,N_8074,N_8240);
or U9287 (N_9287,N_8121,N_8119);
nor U9288 (N_9288,N_8178,N_8087);
or U9289 (N_9289,N_8445,N_8917);
or U9290 (N_9290,N_8868,N_8588);
or U9291 (N_9291,N_8975,N_8882);
nand U9292 (N_9292,N_8497,N_8522);
or U9293 (N_9293,N_8665,N_8337);
nand U9294 (N_9294,N_8101,N_8113);
nand U9295 (N_9295,N_8854,N_8664);
nor U9296 (N_9296,N_8786,N_8077);
nand U9297 (N_9297,N_8488,N_8428);
nand U9298 (N_9298,N_8611,N_8759);
and U9299 (N_9299,N_8911,N_8481);
and U9300 (N_9300,N_8644,N_8334);
nor U9301 (N_9301,N_8338,N_8017);
or U9302 (N_9302,N_8736,N_8456);
or U9303 (N_9303,N_8781,N_8124);
and U9304 (N_9304,N_8983,N_8296);
or U9305 (N_9305,N_8174,N_8159);
and U9306 (N_9306,N_8007,N_8521);
and U9307 (N_9307,N_8274,N_8902);
and U9308 (N_9308,N_8709,N_8582);
or U9309 (N_9309,N_8317,N_8127);
nor U9310 (N_9310,N_8727,N_8050);
xnor U9311 (N_9311,N_8770,N_8730);
and U9312 (N_9312,N_8099,N_8760);
nand U9313 (N_9313,N_8942,N_8907);
nand U9314 (N_9314,N_8156,N_8226);
and U9315 (N_9315,N_8160,N_8586);
and U9316 (N_9316,N_8012,N_8051);
nand U9317 (N_9317,N_8829,N_8655);
and U9318 (N_9318,N_8583,N_8904);
and U9319 (N_9319,N_8847,N_8290);
or U9320 (N_9320,N_8863,N_8252);
nand U9321 (N_9321,N_8584,N_8405);
nor U9322 (N_9322,N_8026,N_8950);
and U9323 (N_9323,N_8111,N_8850);
nor U9324 (N_9324,N_8707,N_8563);
nand U9325 (N_9325,N_8738,N_8171);
or U9326 (N_9326,N_8742,N_8696);
and U9327 (N_9327,N_8149,N_8175);
or U9328 (N_9328,N_8477,N_8292);
and U9329 (N_9329,N_8702,N_8298);
or U9330 (N_9330,N_8688,N_8049);
and U9331 (N_9331,N_8423,N_8552);
xor U9332 (N_9332,N_8498,N_8896);
or U9333 (N_9333,N_8321,N_8899);
or U9334 (N_9334,N_8762,N_8217);
or U9335 (N_9335,N_8489,N_8721);
nor U9336 (N_9336,N_8487,N_8340);
nand U9337 (N_9337,N_8408,N_8831);
nand U9338 (N_9338,N_8852,N_8892);
and U9339 (N_9339,N_8849,N_8472);
nor U9340 (N_9340,N_8980,N_8378);
nor U9341 (N_9341,N_8248,N_8318);
nand U9342 (N_9342,N_8756,N_8999);
nor U9343 (N_9343,N_8734,N_8554);
nor U9344 (N_9344,N_8253,N_8679);
nor U9345 (N_9345,N_8668,N_8144);
and U9346 (N_9346,N_8758,N_8502);
nor U9347 (N_9347,N_8370,N_8794);
xor U9348 (N_9348,N_8024,N_8103);
xnor U9349 (N_9349,N_8417,N_8052);
nor U9350 (N_9350,N_8008,N_8186);
nand U9351 (N_9351,N_8747,N_8172);
nand U9352 (N_9352,N_8909,N_8919);
nor U9353 (N_9353,N_8347,N_8930);
nor U9354 (N_9354,N_8966,N_8439);
and U9355 (N_9355,N_8401,N_8025);
and U9356 (N_9356,N_8258,N_8278);
and U9357 (N_9357,N_8465,N_8598);
nand U9358 (N_9358,N_8303,N_8158);
nor U9359 (N_9359,N_8901,N_8577);
nor U9360 (N_9360,N_8173,N_8542);
or U9361 (N_9361,N_8633,N_8424);
and U9362 (N_9362,N_8518,N_8651);
nor U9363 (N_9363,N_8802,N_8467);
and U9364 (N_9364,N_8805,N_8343);
nor U9365 (N_9365,N_8230,N_8646);
nor U9366 (N_9366,N_8231,N_8082);
nand U9367 (N_9367,N_8003,N_8041);
or U9368 (N_9368,N_8538,N_8474);
or U9369 (N_9369,N_8279,N_8415);
and U9370 (N_9370,N_8595,N_8125);
nand U9371 (N_9371,N_8414,N_8362);
and U9372 (N_9372,N_8383,N_8154);
xor U9373 (N_9373,N_8210,N_8086);
nor U9374 (N_9374,N_8312,N_8045);
nand U9375 (N_9375,N_8653,N_8369);
nand U9376 (N_9376,N_8192,N_8259);
and U9377 (N_9377,N_8812,N_8988);
and U9378 (N_9378,N_8246,N_8105);
and U9379 (N_9379,N_8162,N_8769);
and U9380 (N_9380,N_8450,N_8845);
nor U9381 (N_9381,N_8046,N_8645);
nand U9382 (N_9382,N_8546,N_8109);
nor U9383 (N_9383,N_8236,N_8188);
nand U9384 (N_9384,N_8169,N_8557);
nor U9385 (N_9385,N_8634,N_8223);
nor U9386 (N_9386,N_8525,N_8411);
and U9387 (N_9387,N_8234,N_8083);
nor U9388 (N_9388,N_8056,N_8808);
and U9389 (N_9389,N_8198,N_8635);
nor U9390 (N_9390,N_8963,N_8482);
or U9391 (N_9391,N_8553,N_8938);
nand U9392 (N_9392,N_8676,N_8599);
nor U9393 (N_9393,N_8155,N_8503);
nor U9394 (N_9394,N_8336,N_8925);
nand U9395 (N_9395,N_8316,N_8112);
and U9396 (N_9396,N_8047,N_8304);
nand U9397 (N_9397,N_8565,N_8206);
or U9398 (N_9398,N_8755,N_8208);
nand U9399 (N_9399,N_8928,N_8019);
or U9400 (N_9400,N_8985,N_8936);
xnor U9401 (N_9401,N_8814,N_8510);
or U9402 (N_9402,N_8820,N_8650);
nand U9403 (N_9403,N_8374,N_8737);
nand U9404 (N_9404,N_8744,N_8718);
and U9405 (N_9405,N_8148,N_8079);
xnor U9406 (N_9406,N_8787,N_8617);
and U9407 (N_9407,N_8478,N_8179);
nand U9408 (N_9408,N_8028,N_8460);
xor U9409 (N_9409,N_8416,N_8887);
xor U9410 (N_9410,N_8371,N_8437);
and U9411 (N_9411,N_8286,N_8534);
nand U9412 (N_9412,N_8713,N_8505);
xnor U9413 (N_9413,N_8027,N_8677);
nor U9414 (N_9414,N_8541,N_8958);
nand U9415 (N_9415,N_8404,N_8495);
and U9416 (N_9416,N_8657,N_8833);
xnor U9417 (N_9417,N_8658,N_8570);
and U9418 (N_9418,N_8945,N_8649);
or U9419 (N_9419,N_8295,N_8129);
or U9420 (N_9420,N_8678,N_8998);
nand U9421 (N_9421,N_8607,N_8053);
or U9422 (N_9422,N_8703,N_8168);
nor U9423 (N_9423,N_8622,N_8500);
nor U9424 (N_9424,N_8139,N_8840);
or U9425 (N_9425,N_8205,N_8648);
nor U9426 (N_9426,N_8134,N_8118);
and U9427 (N_9427,N_8357,N_8535);
or U9428 (N_9428,N_8971,N_8796);
or U9429 (N_9429,N_8300,N_8064);
nand U9430 (N_9430,N_8425,N_8871);
and U9431 (N_9431,N_8110,N_8589);
xnor U9432 (N_9432,N_8903,N_8765);
or U9433 (N_9433,N_8395,N_8364);
and U9434 (N_9434,N_8656,N_8795);
and U9435 (N_9435,N_8528,N_8284);
or U9436 (N_9436,N_8203,N_8352);
or U9437 (N_9437,N_8746,N_8062);
or U9438 (N_9438,N_8151,N_8068);
nand U9439 (N_9439,N_8927,N_8107);
xor U9440 (N_9440,N_8876,N_8880);
and U9441 (N_9441,N_8841,N_8741);
nand U9442 (N_9442,N_8468,N_8630);
or U9443 (N_9443,N_8010,N_8380);
xor U9444 (N_9444,N_8596,N_8004);
nand U9445 (N_9445,N_8020,N_8879);
and U9446 (N_9446,N_8579,N_8444);
or U9447 (N_9447,N_8609,N_8332);
and U9448 (N_9448,N_8856,N_8982);
nand U9449 (N_9449,N_8601,N_8305);
or U9450 (N_9450,N_8933,N_8827);
xnor U9451 (N_9451,N_8569,N_8612);
and U9452 (N_9452,N_8313,N_8710);
nor U9453 (N_9453,N_8499,N_8753);
or U9454 (N_9454,N_8108,N_8233);
and U9455 (N_9455,N_8869,N_8224);
and U9456 (N_9456,N_8402,N_8544);
or U9457 (N_9457,N_8382,N_8811);
and U9458 (N_9458,N_8693,N_8572);
nand U9459 (N_9459,N_8215,N_8289);
nand U9460 (N_9460,N_8285,N_8009);
and U9461 (N_9461,N_8931,N_8322);
nand U9462 (N_9462,N_8128,N_8949);
nand U9463 (N_9463,N_8602,N_8143);
xnor U9464 (N_9464,N_8015,N_8523);
nand U9465 (N_9465,N_8698,N_8081);
or U9466 (N_9466,N_8036,N_8326);
nand U9467 (N_9467,N_8287,N_8040);
nor U9468 (N_9468,N_8029,N_8913);
nor U9469 (N_9469,N_8947,N_8864);
nand U9470 (N_9470,N_8990,N_8353);
or U9471 (N_9471,N_8140,N_8365);
xnor U9472 (N_9472,N_8454,N_8951);
nor U9473 (N_9473,N_8441,N_8135);
and U9474 (N_9474,N_8867,N_8526);
and U9475 (N_9475,N_8386,N_8540);
nor U9476 (N_9476,N_8088,N_8822);
or U9477 (N_9477,N_8729,N_8418);
nor U9478 (N_9478,N_8663,N_8573);
nor U9479 (N_9479,N_8807,N_8853);
nand U9480 (N_9480,N_8647,N_8117);
nor U9481 (N_9481,N_8623,N_8245);
nand U9482 (N_9482,N_8241,N_8120);
nor U9483 (N_9483,N_8183,N_8021);
nor U9484 (N_9484,N_8073,N_8834);
and U9485 (N_9485,N_8147,N_8639);
and U9486 (N_9486,N_8859,N_8783);
xnor U9487 (N_9487,N_8372,N_8145);
nor U9488 (N_9488,N_8189,N_8838);
and U9489 (N_9489,N_8213,N_8176);
nor U9490 (N_9490,N_8806,N_8948);
and U9491 (N_9491,N_8306,N_8013);
nor U9492 (N_9492,N_8433,N_8060);
or U9493 (N_9493,N_8277,N_8308);
nand U9494 (N_9494,N_8597,N_8422);
nand U9495 (N_9495,N_8587,N_8547);
and U9496 (N_9496,N_8957,N_8527);
or U9497 (N_9497,N_8861,N_8517);
nor U9498 (N_9498,N_8228,N_8715);
and U9499 (N_9499,N_8182,N_8438);
nor U9500 (N_9500,N_8797,N_8619);
and U9501 (N_9501,N_8520,N_8496);
nor U9502 (N_9502,N_8443,N_8929);
nand U9503 (N_9503,N_8897,N_8268);
nand U9504 (N_9504,N_8380,N_8573);
nor U9505 (N_9505,N_8342,N_8173);
nor U9506 (N_9506,N_8625,N_8190);
nand U9507 (N_9507,N_8566,N_8008);
nand U9508 (N_9508,N_8578,N_8640);
or U9509 (N_9509,N_8848,N_8975);
nor U9510 (N_9510,N_8755,N_8547);
and U9511 (N_9511,N_8708,N_8481);
nand U9512 (N_9512,N_8223,N_8102);
or U9513 (N_9513,N_8562,N_8151);
xor U9514 (N_9514,N_8486,N_8558);
and U9515 (N_9515,N_8206,N_8318);
and U9516 (N_9516,N_8176,N_8856);
nand U9517 (N_9517,N_8840,N_8806);
and U9518 (N_9518,N_8371,N_8762);
nor U9519 (N_9519,N_8031,N_8832);
nand U9520 (N_9520,N_8402,N_8931);
nand U9521 (N_9521,N_8696,N_8731);
nand U9522 (N_9522,N_8895,N_8474);
xnor U9523 (N_9523,N_8936,N_8002);
or U9524 (N_9524,N_8139,N_8456);
xor U9525 (N_9525,N_8448,N_8807);
nand U9526 (N_9526,N_8547,N_8478);
or U9527 (N_9527,N_8206,N_8619);
nor U9528 (N_9528,N_8940,N_8876);
or U9529 (N_9529,N_8317,N_8895);
and U9530 (N_9530,N_8767,N_8597);
nor U9531 (N_9531,N_8159,N_8307);
or U9532 (N_9532,N_8072,N_8822);
or U9533 (N_9533,N_8136,N_8007);
nand U9534 (N_9534,N_8265,N_8931);
nand U9535 (N_9535,N_8122,N_8866);
xor U9536 (N_9536,N_8789,N_8133);
nand U9537 (N_9537,N_8900,N_8155);
nand U9538 (N_9538,N_8071,N_8642);
nand U9539 (N_9539,N_8400,N_8594);
or U9540 (N_9540,N_8660,N_8899);
nand U9541 (N_9541,N_8155,N_8096);
and U9542 (N_9542,N_8379,N_8084);
nand U9543 (N_9543,N_8969,N_8931);
nor U9544 (N_9544,N_8085,N_8745);
and U9545 (N_9545,N_8335,N_8184);
nand U9546 (N_9546,N_8834,N_8840);
nor U9547 (N_9547,N_8809,N_8476);
nor U9548 (N_9548,N_8600,N_8545);
nand U9549 (N_9549,N_8603,N_8936);
nand U9550 (N_9550,N_8985,N_8269);
or U9551 (N_9551,N_8034,N_8488);
and U9552 (N_9552,N_8243,N_8316);
or U9553 (N_9553,N_8077,N_8108);
xor U9554 (N_9554,N_8019,N_8776);
or U9555 (N_9555,N_8637,N_8221);
nand U9556 (N_9556,N_8405,N_8214);
and U9557 (N_9557,N_8958,N_8802);
nor U9558 (N_9558,N_8069,N_8337);
and U9559 (N_9559,N_8468,N_8570);
nand U9560 (N_9560,N_8198,N_8874);
and U9561 (N_9561,N_8229,N_8993);
nand U9562 (N_9562,N_8047,N_8927);
or U9563 (N_9563,N_8340,N_8952);
and U9564 (N_9564,N_8635,N_8299);
and U9565 (N_9565,N_8505,N_8195);
nor U9566 (N_9566,N_8315,N_8465);
nand U9567 (N_9567,N_8458,N_8066);
xor U9568 (N_9568,N_8901,N_8752);
or U9569 (N_9569,N_8936,N_8129);
or U9570 (N_9570,N_8725,N_8336);
nand U9571 (N_9571,N_8364,N_8385);
nor U9572 (N_9572,N_8795,N_8600);
xor U9573 (N_9573,N_8841,N_8944);
nand U9574 (N_9574,N_8892,N_8510);
or U9575 (N_9575,N_8887,N_8132);
or U9576 (N_9576,N_8929,N_8638);
xor U9577 (N_9577,N_8421,N_8554);
and U9578 (N_9578,N_8350,N_8218);
nand U9579 (N_9579,N_8273,N_8413);
and U9580 (N_9580,N_8501,N_8682);
or U9581 (N_9581,N_8934,N_8373);
and U9582 (N_9582,N_8857,N_8976);
and U9583 (N_9583,N_8580,N_8366);
or U9584 (N_9584,N_8261,N_8880);
or U9585 (N_9585,N_8974,N_8562);
or U9586 (N_9586,N_8422,N_8793);
and U9587 (N_9587,N_8499,N_8351);
and U9588 (N_9588,N_8222,N_8623);
or U9589 (N_9589,N_8520,N_8438);
and U9590 (N_9590,N_8603,N_8887);
nor U9591 (N_9591,N_8677,N_8866);
or U9592 (N_9592,N_8707,N_8131);
nand U9593 (N_9593,N_8650,N_8012);
nor U9594 (N_9594,N_8999,N_8197);
and U9595 (N_9595,N_8947,N_8611);
or U9596 (N_9596,N_8594,N_8248);
nand U9597 (N_9597,N_8229,N_8536);
nand U9598 (N_9598,N_8155,N_8729);
nand U9599 (N_9599,N_8937,N_8923);
and U9600 (N_9600,N_8229,N_8691);
nor U9601 (N_9601,N_8957,N_8504);
and U9602 (N_9602,N_8209,N_8121);
xor U9603 (N_9603,N_8733,N_8465);
and U9604 (N_9604,N_8587,N_8228);
nor U9605 (N_9605,N_8865,N_8690);
and U9606 (N_9606,N_8285,N_8134);
and U9607 (N_9607,N_8362,N_8852);
nor U9608 (N_9608,N_8744,N_8921);
and U9609 (N_9609,N_8279,N_8889);
nand U9610 (N_9610,N_8589,N_8239);
xor U9611 (N_9611,N_8830,N_8231);
nor U9612 (N_9612,N_8465,N_8243);
or U9613 (N_9613,N_8537,N_8176);
nor U9614 (N_9614,N_8253,N_8676);
or U9615 (N_9615,N_8312,N_8697);
nand U9616 (N_9616,N_8288,N_8312);
nor U9617 (N_9617,N_8685,N_8888);
or U9618 (N_9618,N_8511,N_8082);
nor U9619 (N_9619,N_8086,N_8878);
and U9620 (N_9620,N_8280,N_8551);
and U9621 (N_9621,N_8344,N_8904);
nand U9622 (N_9622,N_8941,N_8691);
or U9623 (N_9623,N_8313,N_8171);
nand U9624 (N_9624,N_8529,N_8783);
or U9625 (N_9625,N_8040,N_8242);
nor U9626 (N_9626,N_8268,N_8968);
nor U9627 (N_9627,N_8775,N_8564);
and U9628 (N_9628,N_8713,N_8726);
or U9629 (N_9629,N_8822,N_8641);
nor U9630 (N_9630,N_8783,N_8547);
or U9631 (N_9631,N_8709,N_8342);
or U9632 (N_9632,N_8093,N_8437);
xor U9633 (N_9633,N_8547,N_8256);
nand U9634 (N_9634,N_8486,N_8720);
nor U9635 (N_9635,N_8213,N_8444);
nor U9636 (N_9636,N_8516,N_8316);
nor U9637 (N_9637,N_8458,N_8797);
or U9638 (N_9638,N_8251,N_8351);
nand U9639 (N_9639,N_8748,N_8855);
nand U9640 (N_9640,N_8379,N_8020);
nor U9641 (N_9641,N_8027,N_8055);
nor U9642 (N_9642,N_8052,N_8019);
nor U9643 (N_9643,N_8234,N_8763);
or U9644 (N_9644,N_8930,N_8725);
and U9645 (N_9645,N_8863,N_8471);
nor U9646 (N_9646,N_8074,N_8902);
or U9647 (N_9647,N_8335,N_8758);
nand U9648 (N_9648,N_8564,N_8593);
and U9649 (N_9649,N_8104,N_8775);
nand U9650 (N_9650,N_8543,N_8053);
nand U9651 (N_9651,N_8934,N_8286);
nand U9652 (N_9652,N_8811,N_8672);
nand U9653 (N_9653,N_8082,N_8739);
nor U9654 (N_9654,N_8274,N_8034);
and U9655 (N_9655,N_8556,N_8951);
xor U9656 (N_9656,N_8053,N_8965);
nand U9657 (N_9657,N_8456,N_8440);
and U9658 (N_9658,N_8858,N_8754);
and U9659 (N_9659,N_8966,N_8029);
nor U9660 (N_9660,N_8069,N_8049);
or U9661 (N_9661,N_8996,N_8305);
and U9662 (N_9662,N_8382,N_8485);
nand U9663 (N_9663,N_8633,N_8945);
or U9664 (N_9664,N_8014,N_8932);
or U9665 (N_9665,N_8600,N_8115);
or U9666 (N_9666,N_8267,N_8191);
nand U9667 (N_9667,N_8316,N_8534);
nor U9668 (N_9668,N_8605,N_8127);
nand U9669 (N_9669,N_8535,N_8170);
or U9670 (N_9670,N_8105,N_8979);
and U9671 (N_9671,N_8572,N_8069);
or U9672 (N_9672,N_8493,N_8325);
xor U9673 (N_9673,N_8912,N_8842);
nor U9674 (N_9674,N_8036,N_8519);
and U9675 (N_9675,N_8170,N_8942);
and U9676 (N_9676,N_8970,N_8053);
and U9677 (N_9677,N_8311,N_8021);
nor U9678 (N_9678,N_8308,N_8774);
nand U9679 (N_9679,N_8332,N_8640);
nand U9680 (N_9680,N_8938,N_8417);
nand U9681 (N_9681,N_8437,N_8240);
nor U9682 (N_9682,N_8184,N_8461);
nand U9683 (N_9683,N_8859,N_8815);
nand U9684 (N_9684,N_8448,N_8750);
nor U9685 (N_9685,N_8199,N_8267);
nor U9686 (N_9686,N_8252,N_8164);
or U9687 (N_9687,N_8438,N_8373);
and U9688 (N_9688,N_8297,N_8230);
nand U9689 (N_9689,N_8684,N_8785);
and U9690 (N_9690,N_8464,N_8151);
nand U9691 (N_9691,N_8622,N_8787);
xnor U9692 (N_9692,N_8609,N_8045);
xnor U9693 (N_9693,N_8407,N_8370);
and U9694 (N_9694,N_8616,N_8799);
and U9695 (N_9695,N_8858,N_8596);
nand U9696 (N_9696,N_8717,N_8175);
nand U9697 (N_9697,N_8555,N_8397);
nand U9698 (N_9698,N_8268,N_8442);
nor U9699 (N_9699,N_8742,N_8586);
nand U9700 (N_9700,N_8922,N_8294);
and U9701 (N_9701,N_8697,N_8013);
nor U9702 (N_9702,N_8092,N_8605);
or U9703 (N_9703,N_8386,N_8311);
nand U9704 (N_9704,N_8941,N_8009);
nand U9705 (N_9705,N_8178,N_8730);
nand U9706 (N_9706,N_8407,N_8030);
or U9707 (N_9707,N_8549,N_8432);
nand U9708 (N_9708,N_8423,N_8190);
nand U9709 (N_9709,N_8768,N_8900);
and U9710 (N_9710,N_8471,N_8230);
xnor U9711 (N_9711,N_8094,N_8062);
and U9712 (N_9712,N_8683,N_8412);
nor U9713 (N_9713,N_8972,N_8984);
nand U9714 (N_9714,N_8706,N_8875);
and U9715 (N_9715,N_8005,N_8190);
nand U9716 (N_9716,N_8368,N_8211);
or U9717 (N_9717,N_8661,N_8667);
and U9718 (N_9718,N_8134,N_8262);
nand U9719 (N_9719,N_8094,N_8769);
nor U9720 (N_9720,N_8175,N_8965);
xor U9721 (N_9721,N_8093,N_8809);
xnor U9722 (N_9722,N_8812,N_8291);
xor U9723 (N_9723,N_8476,N_8953);
nand U9724 (N_9724,N_8584,N_8005);
or U9725 (N_9725,N_8820,N_8980);
nor U9726 (N_9726,N_8581,N_8609);
or U9727 (N_9727,N_8545,N_8409);
or U9728 (N_9728,N_8584,N_8677);
xnor U9729 (N_9729,N_8578,N_8861);
nor U9730 (N_9730,N_8068,N_8072);
or U9731 (N_9731,N_8331,N_8626);
nand U9732 (N_9732,N_8483,N_8543);
and U9733 (N_9733,N_8734,N_8853);
nor U9734 (N_9734,N_8909,N_8715);
nand U9735 (N_9735,N_8578,N_8327);
nand U9736 (N_9736,N_8401,N_8423);
or U9737 (N_9737,N_8107,N_8397);
and U9738 (N_9738,N_8287,N_8365);
nor U9739 (N_9739,N_8434,N_8104);
nor U9740 (N_9740,N_8228,N_8786);
and U9741 (N_9741,N_8068,N_8905);
nor U9742 (N_9742,N_8465,N_8318);
nand U9743 (N_9743,N_8618,N_8662);
nand U9744 (N_9744,N_8466,N_8912);
nand U9745 (N_9745,N_8195,N_8711);
nor U9746 (N_9746,N_8043,N_8594);
xnor U9747 (N_9747,N_8964,N_8646);
and U9748 (N_9748,N_8247,N_8158);
nand U9749 (N_9749,N_8959,N_8700);
nor U9750 (N_9750,N_8989,N_8606);
or U9751 (N_9751,N_8461,N_8305);
nor U9752 (N_9752,N_8232,N_8505);
and U9753 (N_9753,N_8734,N_8681);
or U9754 (N_9754,N_8422,N_8495);
and U9755 (N_9755,N_8350,N_8657);
nand U9756 (N_9756,N_8862,N_8455);
and U9757 (N_9757,N_8153,N_8934);
or U9758 (N_9758,N_8026,N_8414);
and U9759 (N_9759,N_8366,N_8604);
and U9760 (N_9760,N_8092,N_8430);
nor U9761 (N_9761,N_8357,N_8473);
or U9762 (N_9762,N_8356,N_8330);
and U9763 (N_9763,N_8743,N_8703);
and U9764 (N_9764,N_8423,N_8229);
nand U9765 (N_9765,N_8320,N_8959);
nand U9766 (N_9766,N_8761,N_8317);
nor U9767 (N_9767,N_8207,N_8138);
and U9768 (N_9768,N_8421,N_8566);
nor U9769 (N_9769,N_8126,N_8950);
nand U9770 (N_9770,N_8619,N_8689);
nor U9771 (N_9771,N_8238,N_8830);
or U9772 (N_9772,N_8335,N_8126);
nand U9773 (N_9773,N_8115,N_8581);
nor U9774 (N_9774,N_8706,N_8083);
nand U9775 (N_9775,N_8051,N_8695);
or U9776 (N_9776,N_8475,N_8646);
nor U9777 (N_9777,N_8022,N_8003);
and U9778 (N_9778,N_8450,N_8722);
or U9779 (N_9779,N_8765,N_8184);
and U9780 (N_9780,N_8660,N_8088);
or U9781 (N_9781,N_8581,N_8501);
nor U9782 (N_9782,N_8024,N_8641);
nand U9783 (N_9783,N_8313,N_8633);
or U9784 (N_9784,N_8803,N_8814);
nand U9785 (N_9785,N_8435,N_8526);
nor U9786 (N_9786,N_8649,N_8936);
nand U9787 (N_9787,N_8155,N_8274);
or U9788 (N_9788,N_8574,N_8830);
or U9789 (N_9789,N_8239,N_8181);
xor U9790 (N_9790,N_8287,N_8164);
or U9791 (N_9791,N_8075,N_8984);
nand U9792 (N_9792,N_8671,N_8159);
nand U9793 (N_9793,N_8305,N_8014);
xor U9794 (N_9794,N_8731,N_8993);
and U9795 (N_9795,N_8930,N_8524);
nand U9796 (N_9796,N_8035,N_8868);
nor U9797 (N_9797,N_8929,N_8362);
and U9798 (N_9798,N_8612,N_8645);
nand U9799 (N_9799,N_8605,N_8818);
nor U9800 (N_9800,N_8807,N_8851);
or U9801 (N_9801,N_8261,N_8451);
nor U9802 (N_9802,N_8694,N_8418);
or U9803 (N_9803,N_8097,N_8940);
nor U9804 (N_9804,N_8444,N_8581);
and U9805 (N_9805,N_8978,N_8617);
xnor U9806 (N_9806,N_8436,N_8873);
or U9807 (N_9807,N_8831,N_8481);
xor U9808 (N_9808,N_8089,N_8821);
nor U9809 (N_9809,N_8576,N_8911);
nor U9810 (N_9810,N_8422,N_8759);
nand U9811 (N_9811,N_8653,N_8270);
nor U9812 (N_9812,N_8421,N_8015);
and U9813 (N_9813,N_8046,N_8997);
and U9814 (N_9814,N_8724,N_8849);
or U9815 (N_9815,N_8509,N_8639);
xnor U9816 (N_9816,N_8542,N_8750);
xor U9817 (N_9817,N_8178,N_8638);
or U9818 (N_9818,N_8218,N_8002);
or U9819 (N_9819,N_8330,N_8816);
nand U9820 (N_9820,N_8966,N_8615);
nand U9821 (N_9821,N_8018,N_8999);
nor U9822 (N_9822,N_8210,N_8127);
xnor U9823 (N_9823,N_8452,N_8084);
or U9824 (N_9824,N_8196,N_8412);
and U9825 (N_9825,N_8190,N_8312);
or U9826 (N_9826,N_8072,N_8499);
or U9827 (N_9827,N_8591,N_8849);
nor U9828 (N_9828,N_8724,N_8020);
nor U9829 (N_9829,N_8760,N_8069);
nand U9830 (N_9830,N_8168,N_8112);
or U9831 (N_9831,N_8062,N_8456);
nor U9832 (N_9832,N_8456,N_8714);
nor U9833 (N_9833,N_8600,N_8427);
nand U9834 (N_9834,N_8350,N_8536);
nor U9835 (N_9835,N_8026,N_8872);
nor U9836 (N_9836,N_8289,N_8334);
and U9837 (N_9837,N_8146,N_8004);
nor U9838 (N_9838,N_8199,N_8015);
nor U9839 (N_9839,N_8389,N_8768);
xnor U9840 (N_9840,N_8881,N_8260);
nand U9841 (N_9841,N_8150,N_8523);
xnor U9842 (N_9842,N_8981,N_8420);
xor U9843 (N_9843,N_8435,N_8801);
or U9844 (N_9844,N_8675,N_8830);
nand U9845 (N_9845,N_8084,N_8228);
nand U9846 (N_9846,N_8555,N_8559);
or U9847 (N_9847,N_8625,N_8981);
or U9848 (N_9848,N_8734,N_8659);
or U9849 (N_9849,N_8936,N_8778);
or U9850 (N_9850,N_8929,N_8904);
xnor U9851 (N_9851,N_8690,N_8544);
nand U9852 (N_9852,N_8442,N_8446);
xor U9853 (N_9853,N_8554,N_8517);
nor U9854 (N_9854,N_8099,N_8542);
or U9855 (N_9855,N_8239,N_8369);
or U9856 (N_9856,N_8629,N_8642);
nand U9857 (N_9857,N_8949,N_8523);
or U9858 (N_9858,N_8329,N_8467);
nor U9859 (N_9859,N_8521,N_8511);
nor U9860 (N_9860,N_8952,N_8871);
nor U9861 (N_9861,N_8127,N_8433);
and U9862 (N_9862,N_8298,N_8119);
and U9863 (N_9863,N_8426,N_8343);
nand U9864 (N_9864,N_8831,N_8388);
or U9865 (N_9865,N_8375,N_8166);
xor U9866 (N_9866,N_8211,N_8371);
and U9867 (N_9867,N_8023,N_8553);
nand U9868 (N_9868,N_8841,N_8069);
and U9869 (N_9869,N_8274,N_8855);
nand U9870 (N_9870,N_8269,N_8323);
or U9871 (N_9871,N_8215,N_8031);
and U9872 (N_9872,N_8480,N_8830);
nand U9873 (N_9873,N_8054,N_8981);
and U9874 (N_9874,N_8103,N_8367);
and U9875 (N_9875,N_8951,N_8196);
nand U9876 (N_9876,N_8492,N_8527);
nor U9877 (N_9877,N_8009,N_8027);
xor U9878 (N_9878,N_8231,N_8843);
and U9879 (N_9879,N_8643,N_8575);
nor U9880 (N_9880,N_8705,N_8123);
or U9881 (N_9881,N_8871,N_8627);
and U9882 (N_9882,N_8325,N_8737);
and U9883 (N_9883,N_8494,N_8403);
nand U9884 (N_9884,N_8441,N_8840);
nor U9885 (N_9885,N_8269,N_8897);
nand U9886 (N_9886,N_8331,N_8196);
nand U9887 (N_9887,N_8085,N_8088);
nor U9888 (N_9888,N_8960,N_8147);
nor U9889 (N_9889,N_8098,N_8302);
and U9890 (N_9890,N_8720,N_8993);
nand U9891 (N_9891,N_8277,N_8088);
nor U9892 (N_9892,N_8801,N_8866);
or U9893 (N_9893,N_8995,N_8967);
nor U9894 (N_9894,N_8410,N_8594);
nand U9895 (N_9895,N_8771,N_8930);
and U9896 (N_9896,N_8110,N_8784);
nand U9897 (N_9897,N_8039,N_8214);
or U9898 (N_9898,N_8477,N_8878);
xor U9899 (N_9899,N_8538,N_8784);
nor U9900 (N_9900,N_8857,N_8538);
or U9901 (N_9901,N_8019,N_8818);
nor U9902 (N_9902,N_8320,N_8742);
nor U9903 (N_9903,N_8227,N_8688);
nor U9904 (N_9904,N_8804,N_8918);
nor U9905 (N_9905,N_8398,N_8522);
nand U9906 (N_9906,N_8980,N_8073);
nor U9907 (N_9907,N_8311,N_8338);
and U9908 (N_9908,N_8549,N_8773);
nor U9909 (N_9909,N_8434,N_8471);
or U9910 (N_9910,N_8109,N_8449);
nor U9911 (N_9911,N_8236,N_8795);
nand U9912 (N_9912,N_8611,N_8941);
nor U9913 (N_9913,N_8157,N_8851);
nand U9914 (N_9914,N_8426,N_8336);
or U9915 (N_9915,N_8880,N_8872);
nand U9916 (N_9916,N_8012,N_8004);
or U9917 (N_9917,N_8857,N_8386);
nand U9918 (N_9918,N_8460,N_8250);
nand U9919 (N_9919,N_8760,N_8165);
nor U9920 (N_9920,N_8672,N_8787);
nor U9921 (N_9921,N_8830,N_8825);
nor U9922 (N_9922,N_8946,N_8790);
nand U9923 (N_9923,N_8859,N_8210);
nor U9924 (N_9924,N_8438,N_8230);
and U9925 (N_9925,N_8001,N_8231);
and U9926 (N_9926,N_8531,N_8841);
and U9927 (N_9927,N_8372,N_8326);
or U9928 (N_9928,N_8636,N_8336);
nand U9929 (N_9929,N_8518,N_8244);
nor U9930 (N_9930,N_8950,N_8179);
nor U9931 (N_9931,N_8046,N_8806);
and U9932 (N_9932,N_8960,N_8796);
or U9933 (N_9933,N_8872,N_8377);
or U9934 (N_9934,N_8027,N_8144);
or U9935 (N_9935,N_8429,N_8929);
or U9936 (N_9936,N_8315,N_8641);
nor U9937 (N_9937,N_8670,N_8167);
and U9938 (N_9938,N_8754,N_8843);
nor U9939 (N_9939,N_8145,N_8476);
and U9940 (N_9940,N_8797,N_8669);
nand U9941 (N_9941,N_8066,N_8271);
nand U9942 (N_9942,N_8784,N_8649);
and U9943 (N_9943,N_8310,N_8979);
nand U9944 (N_9944,N_8741,N_8997);
or U9945 (N_9945,N_8641,N_8182);
nor U9946 (N_9946,N_8914,N_8391);
or U9947 (N_9947,N_8402,N_8586);
xor U9948 (N_9948,N_8296,N_8956);
or U9949 (N_9949,N_8172,N_8095);
xnor U9950 (N_9950,N_8741,N_8943);
xnor U9951 (N_9951,N_8855,N_8949);
and U9952 (N_9952,N_8916,N_8056);
and U9953 (N_9953,N_8601,N_8631);
nand U9954 (N_9954,N_8006,N_8387);
and U9955 (N_9955,N_8488,N_8983);
or U9956 (N_9956,N_8459,N_8278);
nand U9957 (N_9957,N_8807,N_8588);
nor U9958 (N_9958,N_8117,N_8001);
or U9959 (N_9959,N_8465,N_8050);
and U9960 (N_9960,N_8486,N_8468);
xnor U9961 (N_9961,N_8352,N_8044);
or U9962 (N_9962,N_8360,N_8700);
or U9963 (N_9963,N_8791,N_8645);
nand U9964 (N_9964,N_8468,N_8368);
xor U9965 (N_9965,N_8386,N_8609);
and U9966 (N_9966,N_8482,N_8115);
nand U9967 (N_9967,N_8350,N_8906);
or U9968 (N_9968,N_8152,N_8692);
nand U9969 (N_9969,N_8197,N_8057);
nor U9970 (N_9970,N_8668,N_8041);
or U9971 (N_9971,N_8239,N_8219);
and U9972 (N_9972,N_8790,N_8323);
or U9973 (N_9973,N_8501,N_8106);
nand U9974 (N_9974,N_8143,N_8814);
or U9975 (N_9975,N_8310,N_8602);
and U9976 (N_9976,N_8213,N_8910);
nor U9977 (N_9977,N_8036,N_8369);
and U9978 (N_9978,N_8565,N_8984);
and U9979 (N_9979,N_8430,N_8053);
or U9980 (N_9980,N_8128,N_8728);
nand U9981 (N_9981,N_8005,N_8837);
and U9982 (N_9982,N_8183,N_8586);
or U9983 (N_9983,N_8074,N_8557);
nor U9984 (N_9984,N_8630,N_8462);
nor U9985 (N_9985,N_8150,N_8730);
and U9986 (N_9986,N_8691,N_8316);
xnor U9987 (N_9987,N_8330,N_8044);
nand U9988 (N_9988,N_8741,N_8343);
or U9989 (N_9989,N_8577,N_8607);
nand U9990 (N_9990,N_8634,N_8953);
and U9991 (N_9991,N_8594,N_8758);
and U9992 (N_9992,N_8517,N_8540);
or U9993 (N_9993,N_8148,N_8437);
or U9994 (N_9994,N_8644,N_8567);
and U9995 (N_9995,N_8468,N_8218);
and U9996 (N_9996,N_8579,N_8550);
and U9997 (N_9997,N_8427,N_8504);
and U9998 (N_9998,N_8343,N_8556);
and U9999 (N_9999,N_8460,N_8103);
or U10000 (N_10000,N_9154,N_9119);
nor U10001 (N_10001,N_9310,N_9749);
and U10002 (N_10002,N_9207,N_9343);
xor U10003 (N_10003,N_9495,N_9179);
nand U10004 (N_10004,N_9445,N_9585);
nor U10005 (N_10005,N_9663,N_9852);
and U10006 (N_10006,N_9622,N_9210);
nand U10007 (N_10007,N_9231,N_9840);
and U10008 (N_10008,N_9972,N_9188);
nor U10009 (N_10009,N_9912,N_9669);
and U10010 (N_10010,N_9047,N_9787);
nor U10011 (N_10011,N_9220,N_9412);
xor U10012 (N_10012,N_9494,N_9111);
nand U10013 (N_10013,N_9628,N_9291);
or U10014 (N_10014,N_9809,N_9515);
and U10015 (N_10015,N_9355,N_9392);
or U10016 (N_10016,N_9872,N_9710);
and U10017 (N_10017,N_9136,N_9238);
and U10018 (N_10018,N_9617,N_9689);
nand U10019 (N_10019,N_9435,N_9977);
or U10020 (N_10020,N_9399,N_9090);
or U10021 (N_10021,N_9096,N_9714);
or U10022 (N_10022,N_9151,N_9288);
nand U10023 (N_10023,N_9674,N_9402);
nor U10024 (N_10024,N_9043,N_9795);
or U10025 (N_10025,N_9286,N_9223);
nor U10026 (N_10026,N_9409,N_9061);
or U10027 (N_10027,N_9479,N_9724);
or U10028 (N_10028,N_9771,N_9906);
nand U10029 (N_10029,N_9611,N_9229);
and U10030 (N_10030,N_9228,N_9967);
and U10031 (N_10031,N_9497,N_9401);
and U10032 (N_10032,N_9793,N_9051);
nand U10033 (N_10033,N_9106,N_9785);
or U10034 (N_10034,N_9079,N_9193);
nand U10035 (N_10035,N_9224,N_9375);
nand U10036 (N_10036,N_9461,N_9650);
and U10037 (N_10037,N_9137,N_9150);
and U10038 (N_10038,N_9128,N_9425);
xor U10039 (N_10039,N_9541,N_9751);
or U10040 (N_10040,N_9177,N_9635);
nand U10041 (N_10041,N_9115,N_9857);
and U10042 (N_10042,N_9518,N_9567);
xor U10043 (N_10043,N_9152,N_9083);
and U10044 (N_10044,N_9510,N_9102);
xnor U10045 (N_10045,N_9995,N_9529);
and U10046 (N_10046,N_9187,N_9269);
or U10047 (N_10047,N_9917,N_9900);
nand U10048 (N_10048,N_9595,N_9608);
and U10049 (N_10049,N_9742,N_9465);
nor U10050 (N_10050,N_9736,N_9033);
nand U10051 (N_10051,N_9904,N_9341);
or U10052 (N_10052,N_9830,N_9261);
nor U10053 (N_10053,N_9557,N_9593);
and U10054 (N_10054,N_9538,N_9705);
nand U10055 (N_10055,N_9773,N_9748);
and U10056 (N_10056,N_9300,N_9896);
or U10057 (N_10057,N_9262,N_9271);
nor U10058 (N_10058,N_9376,N_9321);
nor U10059 (N_10059,N_9373,N_9958);
nor U10060 (N_10060,N_9816,N_9537);
nor U10061 (N_10061,N_9219,N_9333);
or U10062 (N_10062,N_9755,N_9860);
or U10063 (N_10063,N_9670,N_9827);
or U10064 (N_10064,N_9075,N_9189);
or U10065 (N_10065,N_9643,N_9122);
nand U10066 (N_10066,N_9024,N_9902);
nor U10067 (N_10067,N_9569,N_9073);
xor U10068 (N_10068,N_9209,N_9991);
nand U10069 (N_10069,N_9626,N_9535);
or U10070 (N_10070,N_9359,N_9532);
nor U10071 (N_10071,N_9730,N_9947);
nand U10072 (N_10072,N_9215,N_9147);
xor U10073 (N_10073,N_9053,N_9149);
nand U10074 (N_10074,N_9881,N_9020);
and U10075 (N_10075,N_9824,N_9843);
and U10076 (N_10076,N_9839,N_9503);
xnor U10077 (N_10077,N_9492,N_9416);
nand U10078 (N_10078,N_9973,N_9350);
and U10079 (N_10079,N_9031,N_9299);
xnor U10080 (N_10080,N_9968,N_9417);
nand U10081 (N_10081,N_9536,N_9531);
or U10082 (N_10082,N_9358,N_9754);
or U10083 (N_10083,N_9313,N_9138);
xnor U10084 (N_10084,N_9324,N_9411);
and U10085 (N_10085,N_9985,N_9264);
nand U10086 (N_10086,N_9954,N_9914);
nor U10087 (N_10087,N_9928,N_9588);
nand U10088 (N_10088,N_9630,N_9268);
nor U10089 (N_10089,N_9429,N_9239);
nor U10090 (N_10090,N_9513,N_9870);
or U10091 (N_10091,N_9555,N_9481);
and U10092 (N_10092,N_9242,N_9428);
or U10093 (N_10093,N_9794,N_9564);
nand U10094 (N_10094,N_9318,N_9370);
xnor U10095 (N_10095,N_9104,N_9606);
or U10096 (N_10096,N_9576,N_9103);
and U10097 (N_10097,N_9565,N_9533);
nand U10098 (N_10098,N_9380,N_9197);
or U10099 (N_10099,N_9213,N_9680);
or U10100 (N_10100,N_9562,N_9591);
nand U10101 (N_10101,N_9661,N_9191);
and U10102 (N_10102,N_9278,N_9050);
or U10103 (N_10103,N_9303,N_9715);
nand U10104 (N_10104,N_9884,N_9056);
and U10105 (N_10105,N_9903,N_9009);
or U10106 (N_10106,N_9587,N_9552);
and U10107 (N_10107,N_9941,N_9700);
or U10108 (N_10108,N_9022,N_9471);
xnor U10109 (N_10109,N_9498,N_9920);
or U10110 (N_10110,N_9041,N_9062);
nor U10111 (N_10111,N_9944,N_9157);
nor U10112 (N_10112,N_9665,N_9943);
and U10113 (N_10113,N_9989,N_9558);
nor U10114 (N_10114,N_9963,N_9984);
nand U10115 (N_10115,N_9717,N_9257);
xnor U10116 (N_10116,N_9249,N_9232);
nand U10117 (N_10117,N_9378,N_9691);
nand U10118 (N_10118,N_9706,N_9406);
nor U10119 (N_10119,N_9899,N_9699);
nand U10120 (N_10120,N_9357,N_9619);
nor U10121 (N_10121,N_9618,N_9988);
xor U10122 (N_10122,N_9331,N_9776);
and U10123 (N_10123,N_9627,N_9999);
and U10124 (N_10124,N_9256,N_9281);
nand U10125 (N_10125,N_9267,N_9673);
and U10126 (N_10126,N_9400,N_9686);
nor U10127 (N_10127,N_9733,N_9522);
or U10128 (N_10128,N_9372,N_9817);
xnor U10129 (N_10129,N_9616,N_9277);
nand U10130 (N_10130,N_9756,N_9164);
and U10131 (N_10131,N_9089,N_9638);
and U10132 (N_10132,N_9329,N_9875);
and U10133 (N_10133,N_9486,N_9969);
or U10134 (N_10134,N_9194,N_9589);
and U10135 (N_10135,N_9646,N_9226);
nand U10136 (N_10136,N_9470,N_9117);
nand U10137 (N_10137,N_9205,N_9933);
or U10138 (N_10138,N_9764,N_9812);
nor U10139 (N_10139,N_9237,N_9559);
or U10140 (N_10140,N_9605,N_9624);
xor U10141 (N_10141,N_9013,N_9039);
nand U10142 (N_10142,N_9474,N_9678);
xor U10143 (N_10143,N_9453,N_9489);
or U10144 (N_10144,N_9016,N_9444);
and U10145 (N_10145,N_9731,N_9405);
nor U10146 (N_10146,N_9540,N_9586);
nand U10147 (N_10147,N_9332,N_9314);
nor U10148 (N_10148,N_9876,N_9592);
or U10149 (N_10149,N_9190,N_9996);
nor U10150 (N_10150,N_9369,N_9385);
and U10151 (N_10151,N_9085,N_9389);
nor U10152 (N_10152,N_9011,N_9741);
nor U10153 (N_10153,N_9720,N_9603);
xor U10154 (N_10154,N_9502,N_9820);
nor U10155 (N_10155,N_9709,N_9679);
and U10156 (N_10156,N_9055,N_9792);
nor U10157 (N_10157,N_9460,N_9818);
and U10158 (N_10158,N_9544,N_9227);
xor U10159 (N_10159,N_9750,N_9921);
and U10160 (N_10160,N_9295,N_9955);
nor U10161 (N_10161,N_9038,N_9601);
xnor U10162 (N_10162,N_9883,N_9032);
nor U10163 (N_10163,N_9517,N_9124);
or U10164 (N_10164,N_9382,N_9074);
or U10165 (N_10165,N_9415,N_9655);
nor U10166 (N_10166,N_9721,N_9992);
nor U10167 (N_10167,N_9161,N_9484);
nor U10168 (N_10168,N_9446,N_9393);
and U10169 (N_10169,N_9092,N_9637);
and U10170 (N_10170,N_9782,N_9200);
and U10171 (N_10171,N_9671,N_9965);
nand U10172 (N_10172,N_9865,N_9814);
xnor U10173 (N_10173,N_9347,N_9718);
xnor U10174 (N_10174,N_9805,N_9183);
or U10175 (N_10175,N_9916,N_9072);
or U10176 (N_10176,N_9905,N_9110);
and U10177 (N_10177,N_9296,N_9362);
nand U10178 (N_10178,N_9178,N_9482);
or U10179 (N_10179,N_9035,N_9712);
and U10180 (N_10180,N_9897,N_9289);
or U10181 (N_10181,N_9285,N_9107);
nand U10182 (N_10182,N_9521,N_9214);
and U10183 (N_10183,N_9026,N_9174);
nand U10184 (N_10184,N_9182,N_9097);
nand U10185 (N_10185,N_9054,N_9040);
nor U10186 (N_10186,N_9728,N_9675);
nand U10187 (N_10187,N_9560,N_9432);
or U10188 (N_10188,N_9774,N_9911);
or U10189 (N_10189,N_9863,N_9683);
and U10190 (N_10190,N_9623,N_9255);
xnor U10191 (N_10191,N_9848,N_9711);
and U10192 (N_10192,N_9338,N_9422);
nand U10193 (N_10193,N_9767,N_9000);
and U10194 (N_10194,N_9530,N_9993);
nand U10195 (N_10195,N_9468,N_9625);
and U10196 (N_10196,N_9579,N_9994);
xnor U10197 (N_10197,N_9688,N_9936);
nor U10198 (N_10198,N_9088,N_9383);
and U10199 (N_10199,N_9005,N_9421);
or U10200 (N_10200,N_9859,N_9241);
and U10201 (N_10201,N_9456,N_9930);
and U10202 (N_10202,N_9306,N_9156);
and U10203 (N_10203,N_9582,N_9781);
and U10204 (N_10204,N_9997,N_9654);
nand U10205 (N_10205,N_9769,N_9270);
nor U10206 (N_10206,N_9274,N_9835);
nor U10207 (N_10207,N_9173,N_9546);
or U10208 (N_10208,N_9858,N_9121);
nand U10209 (N_10209,N_9808,N_9120);
nand U10210 (N_10210,N_9398,N_9452);
nor U10211 (N_10211,N_9929,N_9135);
nand U10212 (N_10212,N_9263,N_9826);
and U10213 (N_10213,N_9970,N_9259);
nor U10214 (N_10214,N_9974,N_9065);
and U10215 (N_10215,N_9507,N_9685);
nand U10216 (N_10216,N_9790,N_9134);
or U10217 (N_10217,N_9363,N_9339);
nor U10218 (N_10218,N_9433,N_9570);
and U10219 (N_10219,N_9165,N_9240);
and U10220 (N_10220,N_9114,N_9308);
nor U10221 (N_10221,N_9327,N_9312);
or U10222 (N_10222,N_9325,N_9922);
nand U10223 (N_10223,N_9757,N_9634);
xor U10224 (N_10224,N_9353,N_9485);
or U10225 (N_10225,N_9765,N_9801);
nor U10226 (N_10226,N_9804,N_9866);
and U10227 (N_10227,N_9823,N_9130);
xor U10228 (N_10228,N_9335,N_9172);
or U10229 (N_10229,N_9580,N_9366);
or U10230 (N_10230,N_9512,N_9841);
nand U10231 (N_10231,N_9247,N_9059);
or U10232 (N_10232,N_9607,N_9713);
nor U10233 (N_10233,N_9919,N_9046);
and U10234 (N_10234,N_9186,N_9690);
nor U10235 (N_10235,N_9108,N_9519);
and U10236 (N_10236,N_9836,N_9575);
nand U10237 (N_10237,N_9140,N_9923);
and U10238 (N_10238,N_9001,N_9893);
and U10239 (N_10239,N_9282,N_9566);
or U10240 (N_10240,N_9431,N_9057);
and U10241 (N_10241,N_9811,N_9336);
nor U10242 (N_10242,N_9126,N_9722);
and U10243 (N_10243,N_9345,N_9014);
nor U10244 (N_10244,N_9584,N_9028);
nor U10245 (N_10245,N_9891,N_9505);
nand U10246 (N_10246,N_9196,N_9293);
and U10247 (N_10247,N_9473,N_9729);
or U10248 (N_10248,N_9287,N_9745);
nand U10249 (N_10249,N_9660,N_9301);
nor U10250 (N_10250,N_9642,N_9829);
nand U10251 (N_10251,N_9368,N_9957);
or U10252 (N_10252,N_9825,N_9457);
nor U10253 (N_10253,N_9153,N_9162);
xnor U10254 (N_10254,N_9002,N_9077);
and U10255 (N_10255,N_9148,N_9091);
nor U10256 (N_10256,N_9109,N_9596);
xnor U10257 (N_10257,N_9225,N_9658);
and U10258 (N_10258,N_9810,N_9487);
nor U10259 (N_10259,N_9777,N_9390);
or U10260 (N_10260,N_9602,N_9553);
nand U10261 (N_10261,N_9118,N_9788);
nor U10262 (N_10262,N_9501,N_9204);
nor U10263 (N_10263,N_9360,N_9791);
and U10264 (N_10264,N_9842,N_9439);
nand U10265 (N_10265,N_9806,N_9800);
nor U10266 (N_10266,N_9924,N_9049);
nor U10267 (N_10267,N_9942,N_9979);
nand U10268 (N_10268,N_9008,N_9925);
and U10269 (N_10269,N_9139,N_9949);
and U10270 (N_10270,N_9037,N_9869);
and U10271 (N_10271,N_9388,N_9361);
nor U10272 (N_10272,N_9837,N_9123);
or U10273 (N_10273,N_9315,N_9015);
nor U10274 (N_10274,N_9892,N_9180);
and U10275 (N_10275,N_9959,N_9657);
nand U10276 (N_10276,N_9346,N_9420);
nor U10277 (N_10277,N_9600,N_9168);
and U10278 (N_10278,N_9734,N_9832);
xor U10279 (N_10279,N_9952,N_9946);
xnor U10280 (N_10280,N_9276,N_9779);
and U10281 (N_10281,N_9719,N_9543);
nor U10282 (N_10282,N_9095,N_9931);
xor U10283 (N_10283,N_9867,N_9894);
or U10284 (N_10284,N_9986,N_9778);
or U10285 (N_10285,N_9478,N_9890);
nand U10286 (N_10286,N_9855,N_9052);
or U10287 (N_10287,N_9761,N_9907);
and U10288 (N_10288,N_9132,N_9169);
or U10289 (N_10289,N_9760,N_9253);
nor U10290 (N_10290,N_9280,N_9317);
nor U10291 (N_10291,N_9647,N_9845);
and U10292 (N_10292,N_9878,N_9951);
nand U10293 (N_10293,N_9701,N_9396);
or U10294 (N_10294,N_9695,N_9202);
or U10295 (N_10295,N_9094,N_9386);
xnor U10296 (N_10296,N_9950,N_9440);
nand U10297 (N_10297,N_9877,N_9143);
nor U10298 (N_10298,N_9348,N_9514);
and U10299 (N_10299,N_9113,N_9234);
nand U10300 (N_10300,N_9594,N_9737);
and U10301 (N_10301,N_9407,N_9027);
and U10302 (N_10302,N_9762,N_9633);
nor U10303 (N_10303,N_9290,N_9799);
or U10304 (N_10304,N_9323,N_9798);
xnor U10305 (N_10305,N_9956,N_9302);
nor U10306 (N_10306,N_9516,N_9971);
or U10307 (N_10307,N_9058,N_9304);
or U10308 (N_10308,N_9844,N_9007);
nand U10309 (N_10309,N_9019,N_9908);
and U10310 (N_10310,N_9066,N_9145);
or U10311 (N_10311,N_9889,N_9847);
nand U10312 (N_10312,N_9980,N_9454);
and U10313 (N_10313,N_9462,N_9653);
xor U10314 (N_10314,N_9100,N_9233);
or U10315 (N_10315,N_9437,N_9018);
nand U10316 (N_10316,N_9574,N_9604);
or U10317 (N_10317,N_9561,N_9217);
xor U10318 (N_10318,N_9850,N_9404);
or U10319 (N_10319,N_9218,N_9450);
or U10320 (N_10320,N_9463,N_9307);
nor U10321 (N_10321,N_9526,N_9201);
nand U10322 (N_10322,N_9034,N_9822);
nor U10323 (N_10323,N_9427,N_9305);
or U10324 (N_10324,N_9491,N_9081);
or U10325 (N_10325,N_9726,N_9759);
nor U10326 (N_10326,N_9387,N_9648);
nand U10327 (N_10327,N_9069,N_9978);
or U10328 (N_10328,N_9887,N_9155);
nand U10329 (N_10329,N_9459,N_9379);
nor U10330 (N_10330,N_9743,N_9649);
nor U10331 (N_10331,N_9464,N_9248);
and U10332 (N_10332,N_9853,N_9413);
nand U10333 (N_10333,N_9309,N_9086);
and U10334 (N_10334,N_9862,N_9458);
and U10335 (N_10335,N_9403,N_9677);
or U10336 (N_10336,N_9641,N_9397);
nor U10337 (N_10337,N_9932,N_9898);
and U10338 (N_10338,N_9442,N_9640);
nor U10339 (N_10339,N_9236,N_9910);
nor U10340 (N_10340,N_9208,N_9886);
nor U10341 (N_10341,N_9356,N_9708);
nand U10342 (N_10342,N_9112,N_9934);
or U10343 (N_10343,N_9590,N_9030);
nand U10344 (N_10344,N_9849,N_9614);
xnor U10345 (N_10345,N_9735,N_9732);
nor U10346 (N_10346,N_9856,N_9525);
or U10347 (N_10347,N_9477,N_9483);
and U10348 (N_10348,N_9702,N_9753);
xnor U10349 (N_10349,N_9672,N_9802);
xor U10350 (N_10350,N_9636,N_9184);
nor U10351 (N_10351,N_9694,N_9377);
nor U10352 (N_10352,N_9632,N_9195);
xor U10353 (N_10353,N_9349,N_9938);
nor U10354 (N_10354,N_9451,N_9520);
and U10355 (N_10355,N_9846,N_9770);
nand U10356 (N_10356,N_9496,N_9252);
xor U10357 (N_10357,N_9206,N_9344);
xor U10358 (N_10358,N_9352,N_9953);
nand U10359 (N_10359,N_9796,N_9159);
or U10360 (N_10360,N_9101,N_9990);
or U10361 (N_10361,N_9351,N_9266);
or U10362 (N_10362,N_9272,N_9116);
and U10363 (N_10363,N_9983,N_9251);
xor U10364 (N_10364,N_9167,N_9311);
and U10365 (N_10365,N_9629,N_9772);
nand U10366 (N_10366,N_9815,N_9488);
or U10367 (N_10367,N_9668,N_9534);
or U10368 (N_10368,N_9449,N_9775);
nand U10369 (N_10369,N_9163,N_9044);
nand U10370 (N_10370,N_9961,N_9524);
or U10371 (N_10371,N_9504,N_9235);
or U10372 (N_10372,N_9723,N_9676);
nand U10373 (N_10373,N_9328,N_9964);
or U10374 (N_10374,N_9133,N_9063);
nand U10375 (N_10375,N_9230,N_9542);
nor U10376 (N_10376,N_9222,N_9216);
and U10377 (N_10377,N_9864,N_9469);
nand U10378 (N_10378,N_9797,N_9652);
or U10379 (N_10379,N_9273,N_9060);
nor U10380 (N_10380,N_9258,N_9408);
nand U10381 (N_10381,N_9395,N_9704);
and U10382 (N_10382,N_9265,N_9493);
or U10383 (N_10383,N_9364,N_9740);
and U10384 (N_10384,N_9246,N_9577);
xor U10385 (N_10385,N_9430,N_9696);
and U10386 (N_10386,N_9727,N_9374);
and U10387 (N_10387,N_9012,N_9254);
or U10388 (N_10388,N_9684,N_9175);
nor U10389 (N_10389,N_9166,N_9828);
and U10390 (N_10390,N_9913,N_9141);
nor U10391 (N_10391,N_9780,N_9340);
and U10392 (N_10392,N_9813,N_9620);
nor U10393 (N_10393,N_9067,N_9284);
xnor U10394 (N_10394,N_9746,N_9882);
or U10395 (N_10395,N_9539,N_9070);
nand U10396 (N_10396,N_9783,N_9245);
nor U10397 (N_10397,N_9506,N_9275);
or U10398 (N_10398,N_9667,N_9873);
nand U10399 (N_10399,N_9448,N_9631);
nand U10400 (N_10400,N_9698,N_9476);
or U10401 (N_10401,N_9490,N_9467);
nor U10402 (N_10402,N_9045,N_9960);
nand U10403 (N_10403,N_9807,N_9003);
nand U10404 (N_10404,N_9326,N_9426);
and U10405 (N_10405,N_9243,N_9738);
or U10406 (N_10406,N_9871,N_9160);
nor U10407 (N_10407,N_9644,N_9099);
and U10408 (N_10408,N_9029,N_9707);
nand U10409 (N_10409,N_9297,N_9940);
or U10410 (N_10410,N_9692,N_9937);
xor U10411 (N_10411,N_9948,N_9424);
and U10412 (N_10412,N_9320,N_9410);
nor U10413 (N_10413,N_9549,N_9394);
nor U10414 (N_10414,N_9861,N_9693);
nor U10415 (N_10415,N_9578,N_9901);
nor U10416 (N_10416,N_9681,N_9545);
nand U10417 (N_10417,N_9838,N_9260);
nor U10418 (N_10418,N_9758,N_9316);
nand U10419 (N_10419,N_9915,N_9926);
and U10420 (N_10420,N_9093,N_9036);
nor U10421 (N_10421,N_9747,N_9789);
or U10422 (N_10422,N_9144,N_9819);
or U10423 (N_10423,N_9572,N_9547);
and U10424 (N_10424,N_9651,N_9203);
nor U10425 (N_10425,N_9441,N_9414);
or U10426 (N_10426,N_9023,N_9784);
nand U10427 (N_10427,N_9744,N_9199);
nand U10428 (N_10428,N_9599,N_9763);
or U10429 (N_10429,N_9834,N_9573);
nand U10430 (N_10430,N_9766,N_9583);
and U10431 (N_10431,N_9687,N_9945);
and U10432 (N_10432,N_9455,N_9198);
and U10433 (N_10433,N_9017,N_9087);
nor U10434 (N_10434,N_9659,N_9662);
nor U10435 (N_10435,N_9639,N_9752);
or U10436 (N_10436,N_9337,N_9939);
and U10437 (N_10437,N_9645,N_9142);
and U10438 (N_10438,N_9105,N_9998);
nand U10439 (N_10439,N_9021,N_9076);
and U10440 (N_10440,N_9739,N_9621);
xnor U10441 (N_10441,N_9447,N_9082);
or U10442 (N_10442,N_9664,N_9146);
nor U10443 (N_10443,N_9831,N_9221);
nor U10444 (N_10444,N_9499,N_9365);
nor U10445 (N_10445,N_9725,N_9384);
or U10446 (N_10446,N_9851,N_9391);
nand U10447 (N_10447,N_9078,N_9381);
or U10448 (N_10448,N_9127,N_9480);
or U10449 (N_10449,N_9598,N_9472);
nor U10450 (N_10450,N_9125,N_9475);
and U10451 (N_10451,N_9581,N_9367);
nor U10452 (N_10452,N_9319,N_9868);
xor U10453 (N_10453,N_9250,N_9597);
nand U10454 (N_10454,N_9334,N_9025);
nor U10455 (N_10455,N_9098,N_9874);
and U10456 (N_10456,N_9554,N_9064);
and U10457 (N_10457,N_9927,N_9158);
and U10458 (N_10458,N_9419,N_9371);
xnor U10459 (N_10459,N_9354,N_9322);
or U10460 (N_10460,N_9981,N_9283);
nor U10461 (N_10461,N_9610,N_9523);
nor U10462 (N_10462,N_9703,N_9528);
nor U10463 (N_10463,N_9279,N_9129);
nor U10464 (N_10464,N_9192,N_9918);
and U10465 (N_10465,N_9935,N_9244);
or U10466 (N_10466,N_9010,N_9987);
or U10467 (N_10467,N_9568,N_9550);
nand U10468 (N_10468,N_9975,N_9080);
and U10469 (N_10469,N_9211,N_9423);
and U10470 (N_10470,N_9176,N_9551);
nor U10471 (N_10471,N_9292,N_9006);
nor U10472 (N_10472,N_9185,N_9556);
nor U10473 (N_10473,N_9880,N_9895);
nand U10474 (N_10474,N_9418,N_9298);
and U10475 (N_10475,N_9768,N_9212);
nor U10476 (N_10476,N_9854,N_9885);
or U10477 (N_10477,N_9888,N_9803);
nand U10478 (N_10478,N_9966,N_9170);
nor U10479 (N_10479,N_9330,N_9084);
nor U10480 (N_10480,N_9962,N_9466);
nand U10481 (N_10481,N_9656,N_9982);
and U10482 (N_10482,N_9615,N_9548);
or U10483 (N_10483,N_9716,N_9500);
nand U10484 (N_10484,N_9438,N_9609);
and U10485 (N_10485,N_9613,N_9612);
and U10486 (N_10486,N_9294,N_9004);
nand U10487 (N_10487,N_9879,N_9697);
xor U10488 (N_10488,N_9682,N_9443);
and U10489 (N_10489,N_9527,N_9342);
xnor U10490 (N_10490,N_9048,N_9436);
and U10491 (N_10491,N_9434,N_9511);
nor U10492 (N_10492,N_9071,N_9833);
xor U10493 (N_10493,N_9509,N_9571);
and U10494 (N_10494,N_9821,N_9786);
nor U10495 (N_10495,N_9976,N_9563);
nor U10496 (N_10496,N_9042,N_9666);
or U10497 (N_10497,N_9171,N_9068);
nor U10498 (N_10498,N_9508,N_9131);
nor U10499 (N_10499,N_9181,N_9909);
nor U10500 (N_10500,N_9968,N_9115);
and U10501 (N_10501,N_9423,N_9336);
and U10502 (N_10502,N_9197,N_9034);
and U10503 (N_10503,N_9688,N_9002);
nand U10504 (N_10504,N_9110,N_9457);
and U10505 (N_10505,N_9502,N_9274);
or U10506 (N_10506,N_9445,N_9288);
or U10507 (N_10507,N_9937,N_9773);
nand U10508 (N_10508,N_9078,N_9507);
or U10509 (N_10509,N_9039,N_9919);
nor U10510 (N_10510,N_9301,N_9735);
xnor U10511 (N_10511,N_9061,N_9545);
nor U10512 (N_10512,N_9147,N_9239);
or U10513 (N_10513,N_9542,N_9190);
and U10514 (N_10514,N_9435,N_9796);
nand U10515 (N_10515,N_9679,N_9177);
or U10516 (N_10516,N_9223,N_9631);
or U10517 (N_10517,N_9263,N_9308);
nand U10518 (N_10518,N_9619,N_9561);
xor U10519 (N_10519,N_9938,N_9333);
xor U10520 (N_10520,N_9876,N_9956);
nor U10521 (N_10521,N_9069,N_9143);
nand U10522 (N_10522,N_9226,N_9560);
nor U10523 (N_10523,N_9898,N_9902);
and U10524 (N_10524,N_9462,N_9193);
or U10525 (N_10525,N_9293,N_9598);
and U10526 (N_10526,N_9306,N_9018);
nor U10527 (N_10527,N_9383,N_9760);
and U10528 (N_10528,N_9939,N_9594);
nor U10529 (N_10529,N_9977,N_9835);
and U10530 (N_10530,N_9790,N_9078);
nor U10531 (N_10531,N_9600,N_9677);
nand U10532 (N_10532,N_9442,N_9889);
nand U10533 (N_10533,N_9081,N_9294);
nand U10534 (N_10534,N_9140,N_9972);
xor U10535 (N_10535,N_9654,N_9296);
nand U10536 (N_10536,N_9038,N_9724);
nand U10537 (N_10537,N_9462,N_9166);
and U10538 (N_10538,N_9673,N_9752);
nand U10539 (N_10539,N_9803,N_9562);
or U10540 (N_10540,N_9415,N_9302);
nor U10541 (N_10541,N_9877,N_9945);
xnor U10542 (N_10542,N_9502,N_9007);
nor U10543 (N_10543,N_9144,N_9242);
and U10544 (N_10544,N_9388,N_9828);
or U10545 (N_10545,N_9182,N_9179);
or U10546 (N_10546,N_9513,N_9102);
and U10547 (N_10547,N_9735,N_9549);
nand U10548 (N_10548,N_9662,N_9259);
or U10549 (N_10549,N_9168,N_9580);
nor U10550 (N_10550,N_9464,N_9481);
or U10551 (N_10551,N_9510,N_9164);
nand U10552 (N_10552,N_9553,N_9687);
or U10553 (N_10553,N_9979,N_9821);
nor U10554 (N_10554,N_9072,N_9451);
or U10555 (N_10555,N_9244,N_9362);
xnor U10556 (N_10556,N_9161,N_9962);
or U10557 (N_10557,N_9786,N_9489);
and U10558 (N_10558,N_9551,N_9671);
or U10559 (N_10559,N_9637,N_9859);
nor U10560 (N_10560,N_9945,N_9852);
nor U10561 (N_10561,N_9779,N_9365);
and U10562 (N_10562,N_9711,N_9976);
nor U10563 (N_10563,N_9254,N_9395);
nand U10564 (N_10564,N_9916,N_9453);
and U10565 (N_10565,N_9996,N_9004);
xor U10566 (N_10566,N_9983,N_9405);
and U10567 (N_10567,N_9783,N_9047);
or U10568 (N_10568,N_9222,N_9920);
nor U10569 (N_10569,N_9574,N_9524);
nor U10570 (N_10570,N_9032,N_9730);
and U10571 (N_10571,N_9583,N_9083);
or U10572 (N_10572,N_9568,N_9644);
or U10573 (N_10573,N_9826,N_9241);
nand U10574 (N_10574,N_9931,N_9165);
and U10575 (N_10575,N_9136,N_9955);
and U10576 (N_10576,N_9742,N_9710);
and U10577 (N_10577,N_9264,N_9407);
and U10578 (N_10578,N_9338,N_9891);
nand U10579 (N_10579,N_9674,N_9680);
nand U10580 (N_10580,N_9006,N_9637);
and U10581 (N_10581,N_9069,N_9629);
nand U10582 (N_10582,N_9157,N_9025);
nor U10583 (N_10583,N_9871,N_9814);
and U10584 (N_10584,N_9977,N_9909);
nand U10585 (N_10585,N_9984,N_9699);
nand U10586 (N_10586,N_9972,N_9616);
or U10587 (N_10587,N_9799,N_9758);
nor U10588 (N_10588,N_9530,N_9009);
and U10589 (N_10589,N_9501,N_9039);
nor U10590 (N_10590,N_9588,N_9450);
nor U10591 (N_10591,N_9382,N_9672);
nor U10592 (N_10592,N_9854,N_9237);
nor U10593 (N_10593,N_9822,N_9405);
or U10594 (N_10594,N_9728,N_9478);
or U10595 (N_10595,N_9589,N_9405);
nand U10596 (N_10596,N_9501,N_9057);
nor U10597 (N_10597,N_9473,N_9641);
xor U10598 (N_10598,N_9546,N_9965);
or U10599 (N_10599,N_9488,N_9590);
nor U10600 (N_10600,N_9833,N_9845);
xnor U10601 (N_10601,N_9851,N_9349);
nor U10602 (N_10602,N_9847,N_9455);
nand U10603 (N_10603,N_9981,N_9530);
nand U10604 (N_10604,N_9928,N_9708);
nor U10605 (N_10605,N_9480,N_9314);
xnor U10606 (N_10606,N_9383,N_9032);
and U10607 (N_10607,N_9501,N_9185);
or U10608 (N_10608,N_9023,N_9277);
or U10609 (N_10609,N_9159,N_9814);
and U10610 (N_10610,N_9622,N_9449);
xor U10611 (N_10611,N_9728,N_9518);
or U10612 (N_10612,N_9539,N_9968);
or U10613 (N_10613,N_9601,N_9573);
nand U10614 (N_10614,N_9435,N_9417);
nor U10615 (N_10615,N_9924,N_9927);
nor U10616 (N_10616,N_9231,N_9494);
nand U10617 (N_10617,N_9118,N_9967);
xor U10618 (N_10618,N_9655,N_9965);
and U10619 (N_10619,N_9042,N_9521);
and U10620 (N_10620,N_9023,N_9134);
nand U10621 (N_10621,N_9009,N_9350);
xnor U10622 (N_10622,N_9903,N_9788);
nand U10623 (N_10623,N_9065,N_9686);
nand U10624 (N_10624,N_9500,N_9447);
and U10625 (N_10625,N_9492,N_9019);
or U10626 (N_10626,N_9996,N_9009);
or U10627 (N_10627,N_9531,N_9473);
nand U10628 (N_10628,N_9336,N_9378);
nor U10629 (N_10629,N_9868,N_9728);
and U10630 (N_10630,N_9152,N_9829);
nor U10631 (N_10631,N_9247,N_9703);
and U10632 (N_10632,N_9239,N_9763);
nand U10633 (N_10633,N_9247,N_9272);
nor U10634 (N_10634,N_9490,N_9282);
nor U10635 (N_10635,N_9988,N_9362);
nor U10636 (N_10636,N_9235,N_9768);
and U10637 (N_10637,N_9461,N_9682);
nor U10638 (N_10638,N_9422,N_9090);
and U10639 (N_10639,N_9700,N_9669);
and U10640 (N_10640,N_9687,N_9463);
or U10641 (N_10641,N_9252,N_9468);
nand U10642 (N_10642,N_9000,N_9491);
or U10643 (N_10643,N_9638,N_9733);
or U10644 (N_10644,N_9044,N_9613);
or U10645 (N_10645,N_9164,N_9995);
nor U10646 (N_10646,N_9295,N_9319);
nor U10647 (N_10647,N_9501,N_9978);
or U10648 (N_10648,N_9701,N_9029);
or U10649 (N_10649,N_9971,N_9514);
nand U10650 (N_10650,N_9773,N_9027);
and U10651 (N_10651,N_9597,N_9707);
or U10652 (N_10652,N_9991,N_9657);
or U10653 (N_10653,N_9728,N_9274);
or U10654 (N_10654,N_9361,N_9632);
nor U10655 (N_10655,N_9409,N_9551);
nand U10656 (N_10656,N_9330,N_9260);
or U10657 (N_10657,N_9123,N_9212);
and U10658 (N_10658,N_9704,N_9572);
or U10659 (N_10659,N_9168,N_9420);
nand U10660 (N_10660,N_9495,N_9871);
or U10661 (N_10661,N_9918,N_9962);
nor U10662 (N_10662,N_9914,N_9511);
xnor U10663 (N_10663,N_9066,N_9881);
nand U10664 (N_10664,N_9775,N_9269);
xnor U10665 (N_10665,N_9444,N_9912);
nor U10666 (N_10666,N_9510,N_9290);
xnor U10667 (N_10667,N_9852,N_9341);
nor U10668 (N_10668,N_9164,N_9647);
or U10669 (N_10669,N_9519,N_9387);
and U10670 (N_10670,N_9549,N_9608);
or U10671 (N_10671,N_9359,N_9967);
nand U10672 (N_10672,N_9624,N_9532);
nand U10673 (N_10673,N_9889,N_9985);
nand U10674 (N_10674,N_9879,N_9936);
nor U10675 (N_10675,N_9495,N_9276);
nor U10676 (N_10676,N_9378,N_9546);
and U10677 (N_10677,N_9789,N_9596);
and U10678 (N_10678,N_9833,N_9016);
nor U10679 (N_10679,N_9214,N_9640);
nor U10680 (N_10680,N_9984,N_9765);
and U10681 (N_10681,N_9443,N_9633);
nand U10682 (N_10682,N_9641,N_9590);
nor U10683 (N_10683,N_9415,N_9849);
xnor U10684 (N_10684,N_9149,N_9227);
or U10685 (N_10685,N_9616,N_9353);
or U10686 (N_10686,N_9853,N_9547);
or U10687 (N_10687,N_9707,N_9420);
and U10688 (N_10688,N_9542,N_9720);
xnor U10689 (N_10689,N_9437,N_9899);
nor U10690 (N_10690,N_9242,N_9720);
nand U10691 (N_10691,N_9881,N_9741);
and U10692 (N_10692,N_9166,N_9620);
xnor U10693 (N_10693,N_9550,N_9464);
xor U10694 (N_10694,N_9585,N_9778);
nor U10695 (N_10695,N_9163,N_9241);
nand U10696 (N_10696,N_9689,N_9286);
nor U10697 (N_10697,N_9318,N_9543);
nand U10698 (N_10698,N_9196,N_9152);
or U10699 (N_10699,N_9878,N_9355);
nand U10700 (N_10700,N_9950,N_9214);
and U10701 (N_10701,N_9623,N_9963);
and U10702 (N_10702,N_9894,N_9076);
xor U10703 (N_10703,N_9875,N_9470);
and U10704 (N_10704,N_9252,N_9071);
or U10705 (N_10705,N_9037,N_9503);
nor U10706 (N_10706,N_9823,N_9276);
or U10707 (N_10707,N_9458,N_9715);
and U10708 (N_10708,N_9234,N_9208);
nand U10709 (N_10709,N_9486,N_9651);
or U10710 (N_10710,N_9377,N_9616);
and U10711 (N_10711,N_9663,N_9045);
nor U10712 (N_10712,N_9506,N_9311);
nor U10713 (N_10713,N_9847,N_9321);
and U10714 (N_10714,N_9016,N_9761);
and U10715 (N_10715,N_9424,N_9343);
or U10716 (N_10716,N_9137,N_9094);
and U10717 (N_10717,N_9660,N_9710);
nand U10718 (N_10718,N_9456,N_9058);
or U10719 (N_10719,N_9417,N_9140);
nor U10720 (N_10720,N_9322,N_9805);
and U10721 (N_10721,N_9769,N_9021);
and U10722 (N_10722,N_9326,N_9530);
or U10723 (N_10723,N_9263,N_9739);
nand U10724 (N_10724,N_9905,N_9225);
or U10725 (N_10725,N_9726,N_9015);
or U10726 (N_10726,N_9898,N_9528);
and U10727 (N_10727,N_9412,N_9444);
nand U10728 (N_10728,N_9557,N_9815);
nor U10729 (N_10729,N_9018,N_9781);
and U10730 (N_10730,N_9113,N_9355);
and U10731 (N_10731,N_9478,N_9624);
nor U10732 (N_10732,N_9112,N_9082);
nand U10733 (N_10733,N_9635,N_9730);
nor U10734 (N_10734,N_9763,N_9192);
nand U10735 (N_10735,N_9483,N_9489);
nor U10736 (N_10736,N_9909,N_9101);
nor U10737 (N_10737,N_9471,N_9294);
nand U10738 (N_10738,N_9182,N_9564);
nor U10739 (N_10739,N_9362,N_9130);
nor U10740 (N_10740,N_9387,N_9317);
and U10741 (N_10741,N_9138,N_9757);
xor U10742 (N_10742,N_9913,N_9121);
or U10743 (N_10743,N_9613,N_9384);
or U10744 (N_10744,N_9765,N_9449);
or U10745 (N_10745,N_9657,N_9086);
nand U10746 (N_10746,N_9632,N_9423);
or U10747 (N_10747,N_9284,N_9632);
nor U10748 (N_10748,N_9353,N_9423);
xnor U10749 (N_10749,N_9676,N_9130);
nand U10750 (N_10750,N_9339,N_9774);
xnor U10751 (N_10751,N_9018,N_9998);
or U10752 (N_10752,N_9882,N_9620);
xor U10753 (N_10753,N_9964,N_9011);
nand U10754 (N_10754,N_9402,N_9141);
and U10755 (N_10755,N_9302,N_9992);
or U10756 (N_10756,N_9200,N_9143);
nand U10757 (N_10757,N_9155,N_9896);
nor U10758 (N_10758,N_9179,N_9474);
and U10759 (N_10759,N_9663,N_9318);
and U10760 (N_10760,N_9166,N_9628);
and U10761 (N_10761,N_9583,N_9058);
and U10762 (N_10762,N_9199,N_9094);
or U10763 (N_10763,N_9752,N_9882);
or U10764 (N_10764,N_9749,N_9980);
or U10765 (N_10765,N_9797,N_9104);
or U10766 (N_10766,N_9335,N_9715);
nor U10767 (N_10767,N_9828,N_9580);
and U10768 (N_10768,N_9909,N_9177);
or U10769 (N_10769,N_9549,N_9043);
or U10770 (N_10770,N_9095,N_9271);
or U10771 (N_10771,N_9786,N_9607);
and U10772 (N_10772,N_9397,N_9823);
nand U10773 (N_10773,N_9167,N_9445);
nand U10774 (N_10774,N_9718,N_9692);
nor U10775 (N_10775,N_9049,N_9938);
nor U10776 (N_10776,N_9898,N_9877);
nand U10777 (N_10777,N_9716,N_9718);
and U10778 (N_10778,N_9026,N_9913);
and U10779 (N_10779,N_9332,N_9758);
nand U10780 (N_10780,N_9083,N_9134);
nand U10781 (N_10781,N_9407,N_9906);
or U10782 (N_10782,N_9279,N_9496);
nor U10783 (N_10783,N_9030,N_9411);
and U10784 (N_10784,N_9729,N_9722);
xor U10785 (N_10785,N_9992,N_9820);
or U10786 (N_10786,N_9949,N_9566);
and U10787 (N_10787,N_9275,N_9212);
and U10788 (N_10788,N_9676,N_9500);
xnor U10789 (N_10789,N_9167,N_9607);
nand U10790 (N_10790,N_9580,N_9606);
and U10791 (N_10791,N_9352,N_9956);
and U10792 (N_10792,N_9589,N_9551);
and U10793 (N_10793,N_9133,N_9349);
nor U10794 (N_10794,N_9444,N_9070);
and U10795 (N_10795,N_9459,N_9938);
and U10796 (N_10796,N_9018,N_9902);
nand U10797 (N_10797,N_9489,N_9879);
and U10798 (N_10798,N_9301,N_9561);
nand U10799 (N_10799,N_9261,N_9074);
nor U10800 (N_10800,N_9195,N_9700);
and U10801 (N_10801,N_9881,N_9300);
or U10802 (N_10802,N_9076,N_9844);
or U10803 (N_10803,N_9284,N_9075);
nor U10804 (N_10804,N_9498,N_9010);
and U10805 (N_10805,N_9024,N_9958);
xnor U10806 (N_10806,N_9975,N_9520);
and U10807 (N_10807,N_9962,N_9419);
or U10808 (N_10808,N_9443,N_9750);
or U10809 (N_10809,N_9310,N_9565);
nor U10810 (N_10810,N_9158,N_9287);
nor U10811 (N_10811,N_9065,N_9887);
and U10812 (N_10812,N_9049,N_9639);
or U10813 (N_10813,N_9445,N_9193);
nand U10814 (N_10814,N_9541,N_9486);
nor U10815 (N_10815,N_9214,N_9433);
and U10816 (N_10816,N_9641,N_9244);
or U10817 (N_10817,N_9772,N_9319);
xnor U10818 (N_10818,N_9605,N_9339);
nor U10819 (N_10819,N_9509,N_9674);
nand U10820 (N_10820,N_9881,N_9308);
and U10821 (N_10821,N_9901,N_9663);
nor U10822 (N_10822,N_9014,N_9142);
nand U10823 (N_10823,N_9014,N_9455);
xnor U10824 (N_10824,N_9197,N_9928);
and U10825 (N_10825,N_9455,N_9167);
and U10826 (N_10826,N_9762,N_9715);
or U10827 (N_10827,N_9842,N_9586);
xnor U10828 (N_10828,N_9818,N_9067);
nand U10829 (N_10829,N_9138,N_9063);
or U10830 (N_10830,N_9938,N_9565);
nor U10831 (N_10831,N_9953,N_9206);
nor U10832 (N_10832,N_9015,N_9533);
or U10833 (N_10833,N_9544,N_9489);
nand U10834 (N_10834,N_9446,N_9278);
or U10835 (N_10835,N_9894,N_9666);
and U10836 (N_10836,N_9457,N_9305);
nand U10837 (N_10837,N_9784,N_9668);
or U10838 (N_10838,N_9897,N_9295);
nand U10839 (N_10839,N_9877,N_9079);
nand U10840 (N_10840,N_9039,N_9432);
nor U10841 (N_10841,N_9050,N_9513);
and U10842 (N_10842,N_9993,N_9287);
and U10843 (N_10843,N_9049,N_9585);
nor U10844 (N_10844,N_9041,N_9080);
nor U10845 (N_10845,N_9225,N_9822);
xnor U10846 (N_10846,N_9900,N_9013);
xor U10847 (N_10847,N_9549,N_9226);
and U10848 (N_10848,N_9510,N_9284);
and U10849 (N_10849,N_9604,N_9239);
nand U10850 (N_10850,N_9940,N_9737);
nor U10851 (N_10851,N_9987,N_9028);
or U10852 (N_10852,N_9143,N_9271);
nor U10853 (N_10853,N_9869,N_9541);
or U10854 (N_10854,N_9589,N_9094);
or U10855 (N_10855,N_9036,N_9996);
nor U10856 (N_10856,N_9848,N_9648);
or U10857 (N_10857,N_9321,N_9286);
nor U10858 (N_10858,N_9923,N_9224);
nor U10859 (N_10859,N_9081,N_9543);
xnor U10860 (N_10860,N_9481,N_9011);
xnor U10861 (N_10861,N_9546,N_9801);
nor U10862 (N_10862,N_9875,N_9018);
and U10863 (N_10863,N_9667,N_9067);
xnor U10864 (N_10864,N_9619,N_9983);
nor U10865 (N_10865,N_9529,N_9677);
nand U10866 (N_10866,N_9891,N_9855);
xnor U10867 (N_10867,N_9322,N_9323);
nor U10868 (N_10868,N_9212,N_9013);
or U10869 (N_10869,N_9157,N_9485);
and U10870 (N_10870,N_9124,N_9314);
nand U10871 (N_10871,N_9603,N_9411);
nor U10872 (N_10872,N_9428,N_9877);
nand U10873 (N_10873,N_9841,N_9786);
nand U10874 (N_10874,N_9493,N_9007);
or U10875 (N_10875,N_9243,N_9679);
or U10876 (N_10876,N_9763,N_9925);
or U10877 (N_10877,N_9919,N_9678);
and U10878 (N_10878,N_9835,N_9281);
or U10879 (N_10879,N_9789,N_9984);
or U10880 (N_10880,N_9301,N_9167);
nand U10881 (N_10881,N_9140,N_9082);
and U10882 (N_10882,N_9159,N_9887);
nor U10883 (N_10883,N_9311,N_9607);
nor U10884 (N_10884,N_9109,N_9671);
or U10885 (N_10885,N_9789,N_9438);
nand U10886 (N_10886,N_9726,N_9875);
and U10887 (N_10887,N_9354,N_9181);
or U10888 (N_10888,N_9479,N_9845);
or U10889 (N_10889,N_9071,N_9610);
and U10890 (N_10890,N_9003,N_9890);
nor U10891 (N_10891,N_9902,N_9712);
or U10892 (N_10892,N_9869,N_9603);
and U10893 (N_10893,N_9222,N_9492);
xnor U10894 (N_10894,N_9688,N_9309);
or U10895 (N_10895,N_9786,N_9875);
xnor U10896 (N_10896,N_9704,N_9526);
nor U10897 (N_10897,N_9618,N_9852);
nand U10898 (N_10898,N_9815,N_9552);
nand U10899 (N_10899,N_9934,N_9172);
nor U10900 (N_10900,N_9711,N_9617);
nor U10901 (N_10901,N_9800,N_9811);
nor U10902 (N_10902,N_9117,N_9551);
or U10903 (N_10903,N_9925,N_9213);
nor U10904 (N_10904,N_9538,N_9953);
or U10905 (N_10905,N_9583,N_9898);
or U10906 (N_10906,N_9188,N_9931);
or U10907 (N_10907,N_9301,N_9095);
or U10908 (N_10908,N_9752,N_9289);
or U10909 (N_10909,N_9894,N_9293);
nor U10910 (N_10910,N_9947,N_9020);
or U10911 (N_10911,N_9845,N_9331);
nor U10912 (N_10912,N_9486,N_9461);
and U10913 (N_10913,N_9062,N_9099);
or U10914 (N_10914,N_9686,N_9456);
and U10915 (N_10915,N_9962,N_9511);
xnor U10916 (N_10916,N_9282,N_9967);
nand U10917 (N_10917,N_9606,N_9273);
nand U10918 (N_10918,N_9920,N_9420);
or U10919 (N_10919,N_9683,N_9385);
nand U10920 (N_10920,N_9205,N_9364);
nand U10921 (N_10921,N_9428,N_9999);
and U10922 (N_10922,N_9464,N_9929);
nor U10923 (N_10923,N_9639,N_9571);
nor U10924 (N_10924,N_9731,N_9441);
nand U10925 (N_10925,N_9337,N_9372);
nand U10926 (N_10926,N_9832,N_9902);
nand U10927 (N_10927,N_9320,N_9821);
nor U10928 (N_10928,N_9911,N_9063);
and U10929 (N_10929,N_9894,N_9423);
or U10930 (N_10930,N_9196,N_9974);
nor U10931 (N_10931,N_9930,N_9836);
nand U10932 (N_10932,N_9287,N_9819);
nor U10933 (N_10933,N_9952,N_9402);
or U10934 (N_10934,N_9279,N_9897);
and U10935 (N_10935,N_9161,N_9731);
nor U10936 (N_10936,N_9668,N_9929);
and U10937 (N_10937,N_9824,N_9494);
and U10938 (N_10938,N_9054,N_9004);
and U10939 (N_10939,N_9808,N_9935);
nand U10940 (N_10940,N_9904,N_9276);
nand U10941 (N_10941,N_9431,N_9654);
and U10942 (N_10942,N_9855,N_9106);
and U10943 (N_10943,N_9058,N_9057);
xor U10944 (N_10944,N_9376,N_9372);
nand U10945 (N_10945,N_9553,N_9658);
nand U10946 (N_10946,N_9454,N_9670);
xnor U10947 (N_10947,N_9852,N_9407);
and U10948 (N_10948,N_9107,N_9241);
nor U10949 (N_10949,N_9208,N_9603);
nand U10950 (N_10950,N_9314,N_9501);
and U10951 (N_10951,N_9935,N_9132);
or U10952 (N_10952,N_9072,N_9719);
or U10953 (N_10953,N_9652,N_9572);
xnor U10954 (N_10954,N_9636,N_9288);
or U10955 (N_10955,N_9545,N_9039);
xor U10956 (N_10956,N_9521,N_9083);
nand U10957 (N_10957,N_9240,N_9345);
nand U10958 (N_10958,N_9262,N_9259);
and U10959 (N_10959,N_9104,N_9720);
nand U10960 (N_10960,N_9442,N_9816);
nor U10961 (N_10961,N_9046,N_9773);
xnor U10962 (N_10962,N_9175,N_9423);
and U10963 (N_10963,N_9641,N_9985);
or U10964 (N_10964,N_9394,N_9920);
and U10965 (N_10965,N_9153,N_9936);
nand U10966 (N_10966,N_9914,N_9595);
and U10967 (N_10967,N_9015,N_9046);
nor U10968 (N_10968,N_9451,N_9711);
nand U10969 (N_10969,N_9974,N_9291);
nor U10970 (N_10970,N_9145,N_9711);
or U10971 (N_10971,N_9191,N_9159);
or U10972 (N_10972,N_9486,N_9744);
nand U10973 (N_10973,N_9512,N_9854);
nor U10974 (N_10974,N_9677,N_9741);
nand U10975 (N_10975,N_9067,N_9496);
xnor U10976 (N_10976,N_9382,N_9495);
nand U10977 (N_10977,N_9520,N_9738);
and U10978 (N_10978,N_9789,N_9871);
and U10979 (N_10979,N_9438,N_9204);
and U10980 (N_10980,N_9193,N_9298);
or U10981 (N_10981,N_9853,N_9552);
or U10982 (N_10982,N_9407,N_9987);
and U10983 (N_10983,N_9437,N_9014);
nand U10984 (N_10984,N_9687,N_9876);
and U10985 (N_10985,N_9098,N_9162);
and U10986 (N_10986,N_9092,N_9444);
and U10987 (N_10987,N_9771,N_9082);
or U10988 (N_10988,N_9115,N_9124);
nand U10989 (N_10989,N_9159,N_9861);
nand U10990 (N_10990,N_9438,N_9409);
and U10991 (N_10991,N_9218,N_9417);
and U10992 (N_10992,N_9173,N_9463);
nand U10993 (N_10993,N_9904,N_9169);
or U10994 (N_10994,N_9012,N_9657);
xnor U10995 (N_10995,N_9809,N_9700);
nor U10996 (N_10996,N_9142,N_9816);
and U10997 (N_10997,N_9143,N_9448);
or U10998 (N_10998,N_9599,N_9855);
and U10999 (N_10999,N_9889,N_9958);
nand U11000 (N_11000,N_10582,N_10584);
and U11001 (N_11001,N_10031,N_10300);
nand U11002 (N_11002,N_10133,N_10797);
nand U11003 (N_11003,N_10825,N_10127);
and U11004 (N_11004,N_10604,N_10730);
or U11005 (N_11005,N_10161,N_10281);
nor U11006 (N_11006,N_10726,N_10768);
xor U11007 (N_11007,N_10421,N_10263);
and U11008 (N_11008,N_10152,N_10557);
nor U11009 (N_11009,N_10747,N_10635);
and U11010 (N_11010,N_10167,N_10213);
or U11011 (N_11011,N_10120,N_10566);
or U11012 (N_11012,N_10794,N_10148);
nor U11013 (N_11013,N_10870,N_10307);
nor U11014 (N_11014,N_10625,N_10876);
and U11015 (N_11015,N_10012,N_10224);
and U11016 (N_11016,N_10991,N_10953);
nor U11017 (N_11017,N_10471,N_10862);
and U11018 (N_11018,N_10280,N_10248);
or U11019 (N_11019,N_10048,N_10312);
nand U11020 (N_11020,N_10631,N_10542);
and U11021 (N_11021,N_10569,N_10232);
nand U11022 (N_11022,N_10654,N_10922);
nor U11023 (N_11023,N_10897,N_10888);
nand U11024 (N_11024,N_10598,N_10125);
and U11025 (N_11025,N_10370,N_10196);
nor U11026 (N_11026,N_10361,N_10086);
xor U11027 (N_11027,N_10126,N_10181);
nand U11028 (N_11028,N_10366,N_10138);
nand U11029 (N_11029,N_10419,N_10273);
or U11030 (N_11030,N_10121,N_10425);
xnor U11031 (N_11031,N_10223,N_10941);
nand U11032 (N_11032,N_10387,N_10154);
or U11033 (N_11033,N_10055,N_10701);
nand U11034 (N_11034,N_10008,N_10694);
and U11035 (N_11035,N_10053,N_10347);
and U11036 (N_11036,N_10472,N_10474);
and U11037 (N_11037,N_10489,N_10191);
nor U11038 (N_11038,N_10783,N_10688);
nor U11039 (N_11039,N_10270,N_10689);
nor U11040 (N_11040,N_10993,N_10731);
or U11041 (N_11041,N_10799,N_10315);
and U11042 (N_11042,N_10013,N_10868);
nor U11043 (N_11043,N_10547,N_10195);
xor U11044 (N_11044,N_10754,N_10227);
xor U11045 (N_11045,N_10068,N_10708);
nand U11046 (N_11046,N_10554,N_10463);
or U11047 (N_11047,N_10847,N_10705);
or U11048 (N_11048,N_10653,N_10147);
and U11049 (N_11049,N_10960,N_10159);
and U11050 (N_11050,N_10518,N_10545);
nand U11051 (N_11051,N_10683,N_10549);
or U11052 (N_11052,N_10458,N_10050);
or U11053 (N_11053,N_10484,N_10795);
and U11054 (N_11054,N_10362,N_10681);
nand U11055 (N_11055,N_10771,N_10912);
or U11056 (N_11056,N_10641,N_10809);
nand U11057 (N_11057,N_10942,N_10719);
nor U11058 (N_11058,N_10402,N_10575);
and U11059 (N_11059,N_10742,N_10003);
nand U11060 (N_11060,N_10793,N_10216);
nor U11061 (N_11061,N_10913,N_10439);
and U11062 (N_11062,N_10666,N_10951);
and U11063 (N_11063,N_10811,N_10093);
xnor U11064 (N_11064,N_10643,N_10237);
nor U11065 (N_11065,N_10021,N_10269);
nand U11066 (N_11066,N_10620,N_10985);
nand U11067 (N_11067,N_10442,N_10283);
or U11068 (N_11068,N_10788,N_10473);
nand U11069 (N_11069,N_10998,N_10065);
or U11070 (N_11070,N_10395,N_10856);
nor U11071 (N_11071,N_10634,N_10408);
or U11072 (N_11072,N_10293,N_10690);
nand U11073 (N_11073,N_10578,N_10692);
nor U11074 (N_11074,N_10567,N_10679);
nand U11075 (N_11075,N_10324,N_10492);
or U11076 (N_11076,N_10657,N_10116);
nor U11077 (N_11077,N_10109,N_10864);
or U11078 (N_11078,N_10201,N_10874);
nor U11079 (N_11079,N_10958,N_10233);
nand U11080 (N_11080,N_10254,N_10556);
nor U11081 (N_11081,N_10524,N_10072);
or U11082 (N_11082,N_10215,N_10423);
xnor U11083 (N_11083,N_10606,N_10268);
nand U11084 (N_11084,N_10616,N_10267);
or U11085 (N_11085,N_10346,N_10418);
nor U11086 (N_11086,N_10735,N_10150);
nand U11087 (N_11087,N_10211,N_10710);
nand U11088 (N_11088,N_10943,N_10928);
and U11089 (N_11089,N_10308,N_10615);
or U11090 (N_11090,N_10059,N_10202);
nand U11091 (N_11091,N_10130,N_10284);
and U11092 (N_11092,N_10443,N_10949);
and U11093 (N_11093,N_10365,N_10737);
nor U11094 (N_11094,N_10781,N_10787);
xnor U11095 (N_11095,N_10400,N_10687);
nor U11096 (N_11096,N_10617,N_10818);
and U11097 (N_11097,N_10416,N_10946);
nand U11098 (N_11098,N_10626,N_10973);
nor U11099 (N_11099,N_10497,N_10672);
nand U11100 (N_11100,N_10748,N_10374);
nor U11101 (N_11101,N_10071,N_10618);
or U11102 (N_11102,N_10843,N_10565);
nand U11103 (N_11103,N_10409,N_10450);
or U11104 (N_11104,N_10822,N_10499);
and U11105 (N_11105,N_10455,N_10963);
and U11106 (N_11106,N_10983,N_10319);
and U11107 (N_11107,N_10887,N_10298);
or U11108 (N_11108,N_10774,N_10314);
nor U11109 (N_11109,N_10982,N_10173);
or U11110 (N_11110,N_10190,N_10009);
nor U11111 (N_11111,N_10453,N_10915);
or U11112 (N_11112,N_10994,N_10881);
xor U11113 (N_11113,N_10807,N_10403);
nand U11114 (N_11114,N_10430,N_10017);
and U11115 (N_11115,N_10845,N_10386);
or U11116 (N_11116,N_10686,N_10305);
or U11117 (N_11117,N_10933,N_10873);
nand U11118 (N_11118,N_10583,N_10251);
or U11119 (N_11119,N_10188,N_10790);
nor U11120 (N_11120,N_10931,N_10665);
and U11121 (N_11121,N_10144,N_10054);
and U11122 (N_11122,N_10945,N_10980);
and U11123 (N_11123,N_10066,N_10898);
xnor U11124 (N_11124,N_10350,N_10537);
nand U11125 (N_11125,N_10457,N_10630);
xor U11126 (N_11126,N_10543,N_10380);
or U11127 (N_11127,N_10860,N_10834);
nor U11128 (N_11128,N_10718,N_10494);
or U11129 (N_11129,N_10580,N_10156);
nor U11130 (N_11130,N_10971,N_10287);
or U11131 (N_11131,N_10544,N_10128);
nand U11132 (N_11132,N_10146,N_10744);
and U11133 (N_11133,N_10521,N_10548);
or U11134 (N_11134,N_10516,N_10527);
and U11135 (N_11135,N_10791,N_10288);
and U11136 (N_11136,N_10083,N_10486);
nand U11137 (N_11137,N_10610,N_10950);
or U11138 (N_11138,N_10640,N_10972);
nand U11139 (N_11139,N_10414,N_10773);
or U11140 (N_11140,N_10246,N_10883);
or U11141 (N_11141,N_10668,N_10452);
or U11142 (N_11142,N_10884,N_10675);
xnor U11143 (N_11143,N_10759,N_10658);
nand U11144 (N_11144,N_10290,N_10784);
and U11145 (N_11145,N_10096,N_10299);
nor U11146 (N_11146,N_10381,N_10798);
and U11147 (N_11147,N_10094,N_10622);
nand U11148 (N_11148,N_10422,N_10558);
nand U11149 (N_11149,N_10519,N_10424);
and U11150 (N_11150,N_10821,N_10179);
nand U11151 (N_11151,N_10377,N_10696);
and U11152 (N_11152,N_10114,N_10378);
nor U11153 (N_11153,N_10568,N_10789);
or U11154 (N_11154,N_10230,N_10820);
xnor U11155 (N_11155,N_10857,N_10770);
and U11156 (N_11156,N_10496,N_10182);
nand U11157 (N_11157,N_10741,N_10530);
and U11158 (N_11158,N_10069,N_10674);
and U11159 (N_11159,N_10670,N_10603);
nand U11160 (N_11160,N_10819,N_10392);
nor U11161 (N_11161,N_10858,N_10802);
nand U11162 (N_11162,N_10357,N_10738);
or U11163 (N_11163,N_10384,N_10602);
xor U11164 (N_11164,N_10221,N_10478);
nand U11165 (N_11165,N_10057,N_10706);
or U11166 (N_11166,N_10333,N_10174);
nor U11167 (N_11167,N_10918,N_10451);
and U11168 (N_11168,N_10662,N_10260);
nor U11169 (N_11169,N_10483,N_10212);
and U11170 (N_11170,N_10011,N_10752);
nand U11171 (N_11171,N_10728,N_10217);
xor U11172 (N_11172,N_10824,N_10029);
nand U11173 (N_11173,N_10895,N_10529);
or U11174 (N_11174,N_10398,N_10574);
and U11175 (N_11175,N_10426,N_10841);
nor U11176 (N_11176,N_10459,N_10623);
nand U11177 (N_11177,N_10515,N_10509);
and U11178 (N_11178,N_10778,N_10780);
nor U11179 (N_11179,N_10330,N_10866);
xor U11180 (N_11180,N_10326,N_10938);
or U11181 (N_11181,N_10769,N_10844);
or U11182 (N_11182,N_10647,N_10320);
or U11183 (N_11183,N_10520,N_10792);
or U11184 (N_11184,N_10231,N_10756);
nor U11185 (N_11185,N_10110,N_10240);
nand U11186 (N_11186,N_10100,N_10523);
nand U11187 (N_11187,N_10352,N_10976);
or U11188 (N_11188,N_10882,N_10732);
nand U11189 (N_11189,N_10341,N_10467);
nand U11190 (N_11190,N_10318,N_10253);
nand U11191 (N_11191,N_10045,N_10711);
and U11192 (N_11192,N_10353,N_10313);
or U11193 (N_11193,N_10061,N_10677);
nand U11194 (N_11194,N_10925,N_10908);
nor U11195 (N_11195,N_10861,N_10279);
nand U11196 (N_11196,N_10010,N_10652);
nor U11197 (N_11197,N_10228,N_10257);
nor U11198 (N_11198,N_10927,N_10644);
or U11199 (N_11199,N_10937,N_10405);
or U11200 (N_11200,N_10002,N_10812);
or U11201 (N_11201,N_10975,N_10828);
nand U11202 (N_11202,N_10389,N_10546);
or U11203 (N_11203,N_10135,N_10382);
and U11204 (N_11204,N_10241,N_10725);
nor U11205 (N_11205,N_10219,N_10225);
nand U11206 (N_11206,N_10907,N_10076);
xnor U11207 (N_11207,N_10536,N_10436);
nor U11208 (N_11208,N_10137,N_10080);
nand U11209 (N_11209,N_10921,N_10996);
nand U11210 (N_11210,N_10999,N_10619);
or U11211 (N_11211,N_10255,N_10988);
or U11212 (N_11212,N_10599,N_10169);
nor U11213 (N_11213,N_10573,N_10020);
or U11214 (N_11214,N_10676,N_10614);
or U11215 (N_11215,N_10930,N_10415);
or U11216 (N_11216,N_10208,N_10659);
nand U11217 (N_11217,N_10709,N_10296);
and U11218 (N_11218,N_10262,N_10859);
and U11219 (N_11219,N_10265,N_10707);
and U11220 (N_11220,N_10149,N_10890);
and U11221 (N_11221,N_10328,N_10823);
or U11222 (N_11222,N_10685,N_10060);
nand U11223 (N_11223,N_10244,N_10301);
or U11224 (N_11224,N_10597,N_10372);
or U11225 (N_11225,N_10981,N_10517);
or U11226 (N_11226,N_10266,N_10648);
and U11227 (N_11227,N_10295,N_10304);
xnor U11228 (N_11228,N_10902,N_10199);
and U11229 (N_11229,N_10891,N_10796);
or U11230 (N_11230,N_10838,N_10379);
or U11231 (N_11231,N_10289,N_10833);
nand U11232 (N_11232,N_10369,N_10772);
nor U11233 (N_11233,N_10691,N_10186);
xor U11234 (N_11234,N_10829,N_10349);
xnor U11235 (N_11235,N_10965,N_10183);
nor U11236 (N_11236,N_10172,N_10785);
and U11237 (N_11237,N_10826,N_10344);
nor U11238 (N_11238,N_10721,N_10562);
nand U11239 (N_11239,N_10383,N_10629);
and U11240 (N_11240,N_10175,N_10848);
nand U11241 (N_11241,N_10464,N_10206);
and U11242 (N_11242,N_10724,N_10277);
and U11243 (N_11243,N_10052,N_10892);
nand U11244 (N_11244,N_10438,N_10417);
nand U11245 (N_11245,N_10209,N_10220);
nor U11246 (N_11246,N_10952,N_10143);
or U11247 (N_11247,N_10038,N_10396);
nand U11248 (N_11248,N_10099,N_10513);
or U11249 (N_11249,N_10967,N_10385);
and U11250 (N_11250,N_10158,N_10506);
and U11251 (N_11251,N_10258,N_10024);
or U11252 (N_11252,N_10164,N_10957);
or U11253 (N_11253,N_10739,N_10118);
nand U11254 (N_11254,N_10485,N_10503);
nor U11255 (N_11255,N_10673,N_10322);
or U11256 (N_11256,N_10460,N_10786);
nand U11257 (N_11257,N_10987,N_10766);
and U11258 (N_11258,N_10663,N_10872);
or U11259 (N_11259,N_10340,N_10166);
xor U11260 (N_11260,N_10753,N_10391);
nor U11261 (N_11261,N_10292,N_10440);
and U11262 (N_11262,N_10611,N_10498);
or U11263 (N_11263,N_10302,N_10505);
nor U11264 (N_11264,N_10073,N_10758);
and U11265 (N_11265,N_10194,N_10715);
and U11266 (N_11266,N_10153,N_10348);
and U11267 (N_11267,N_10399,N_10512);
or U11268 (N_11268,N_10466,N_10388);
and U11269 (N_11269,N_10669,N_10160);
nand U11270 (N_11270,N_10555,N_10596);
nor U11271 (N_11271,N_10712,N_10016);
nor U11272 (N_11272,N_10112,N_10563);
nor U11273 (N_11273,N_10141,N_10911);
or U11274 (N_11274,N_10311,N_10041);
nand U11275 (N_11275,N_10218,N_10204);
and U11276 (N_11276,N_10810,N_10875);
nor U11277 (N_11277,N_10886,N_10782);
xor U11278 (N_11278,N_10015,N_10877);
and U11279 (N_11279,N_10334,N_10461);
nand U11280 (N_11280,N_10056,N_10222);
and U11281 (N_11281,N_10920,N_10743);
and U11282 (N_11282,N_10207,N_10282);
or U11283 (N_11283,N_10551,N_10081);
and U11284 (N_11284,N_10637,N_10085);
nand U11285 (N_11285,N_10095,N_10746);
nor U11286 (N_11286,N_10878,N_10642);
nand U11287 (N_11287,N_10944,N_10140);
nand U11288 (N_11288,N_10779,N_10363);
or U11289 (N_11289,N_10437,N_10034);
and U11290 (N_11290,N_10051,N_10074);
nor U11291 (N_11291,N_10904,N_10638);
xor U11292 (N_11292,N_10680,N_10579);
nand U11293 (N_11293,N_10919,N_10561);
xnor U11294 (N_11294,N_10197,N_10235);
nor U11295 (N_11295,N_10023,N_10343);
and U11296 (N_11296,N_10835,N_10851);
and U11297 (N_11297,N_10504,N_10502);
nand U11298 (N_11298,N_10456,N_10903);
nor U11299 (N_11299,N_10271,N_10581);
nor U11300 (N_11300,N_10410,N_10522);
nor U11301 (N_11301,N_10084,N_10462);
and U11302 (N_11302,N_10142,N_10840);
or U11303 (N_11303,N_10572,N_10560);
and U11304 (N_11304,N_10433,N_10532);
or U11305 (N_11305,N_10526,N_10699);
nand U11306 (N_11306,N_10275,N_10989);
xor U11307 (N_11307,N_10979,N_10869);
nand U11308 (N_11308,N_10853,N_10813);
nand U11309 (N_11309,N_10600,N_10808);
nor U11310 (N_11310,N_10291,N_10047);
and U11311 (N_11311,N_10087,N_10256);
or U11312 (N_11312,N_10977,N_10511);
and U11313 (N_11313,N_10645,N_10203);
nor U11314 (N_11314,N_10839,N_10624);
and U11315 (N_11315,N_10978,N_10264);
and U11316 (N_11316,N_10594,N_10803);
and U11317 (N_11317,N_10590,N_10032);
nand U11318 (N_11318,N_10553,N_10830);
nand U11319 (N_11319,N_10576,N_10805);
xnor U11320 (N_11320,N_10867,N_10088);
and U11321 (N_11321,N_10984,N_10124);
nor U11322 (N_11322,N_10577,N_10495);
nor U11323 (N_11323,N_10401,N_10661);
and U11324 (N_11324,N_10698,N_10000);
nor U11325 (N_11325,N_10633,N_10588);
or U11326 (N_11326,N_10508,N_10033);
nand U11327 (N_11327,N_10476,N_10444);
nand U11328 (N_11328,N_10815,N_10342);
or U11329 (N_11329,N_10310,N_10098);
or U11330 (N_11330,N_10354,N_10990);
and U11331 (N_11331,N_10850,N_10964);
or U11332 (N_11332,N_10490,N_10407);
xnor U11333 (N_11333,N_10373,N_10238);
or U11334 (N_11334,N_10723,N_10740);
nor U11335 (N_11335,N_10171,N_10406);
and U11336 (N_11336,N_10954,N_10356);
and U11337 (N_11337,N_10014,N_10432);
xnor U11338 (N_11338,N_10716,N_10533);
nand U11339 (N_11339,N_10760,N_10180);
nor U11340 (N_11340,N_10360,N_10170);
or U11341 (N_11341,N_10077,N_10210);
nand U11342 (N_11342,N_10046,N_10855);
and U11343 (N_11343,N_10136,N_10028);
and U11344 (N_11344,N_10193,N_10816);
nor U11345 (N_11345,N_10704,N_10935);
nor U11346 (N_11346,N_10479,N_10493);
xor U11347 (N_11347,N_10607,N_10249);
nand U11348 (N_11348,N_10037,N_10044);
and U11349 (N_11349,N_10974,N_10649);
and U11350 (N_11350,N_10157,N_10693);
xor U11351 (N_11351,N_10682,N_10684);
and U11352 (N_11352,N_10245,N_10309);
or U11353 (N_11353,N_10910,N_10286);
and U11354 (N_11354,N_10487,N_10697);
xor U11355 (N_11355,N_10132,N_10119);
nor U11356 (N_11356,N_10539,N_10940);
and U11357 (N_11357,N_10986,N_10500);
or U11358 (N_11358,N_10226,N_10700);
nand U11359 (N_11359,N_10468,N_10936);
and U11360 (N_11360,N_10660,N_10331);
or U11361 (N_11361,N_10777,N_10107);
xor U11362 (N_11362,N_10272,N_10488);
nor U11363 (N_11363,N_10108,N_10064);
or U11364 (N_11364,N_10961,N_10534);
nor U11365 (N_11365,N_10134,N_10702);
nand U11366 (N_11366,N_10062,N_10894);
and U11367 (N_11367,N_10900,N_10899);
nand U11368 (N_11368,N_10089,N_10750);
and U11369 (N_11369,N_10470,N_10703);
nor U11370 (N_11370,N_10814,N_10997);
nand U11371 (N_11371,N_10042,N_10025);
or U11372 (N_11372,N_10448,N_10541);
xnor U11373 (N_11373,N_10192,N_10454);
and U11374 (N_11374,N_10612,N_10091);
nand U11375 (N_11375,N_10429,N_10854);
and U11376 (N_11376,N_10105,N_10411);
nand U11377 (N_11377,N_10734,N_10528);
or U11378 (N_11378,N_10075,N_10906);
xor U11379 (N_11379,N_10306,N_10336);
and U11380 (N_11380,N_10278,N_10274);
xor U11381 (N_11381,N_10131,N_10200);
or U11382 (N_11382,N_10639,N_10939);
or U11383 (N_11383,N_10303,N_10355);
xnor U11384 (N_11384,N_10924,N_10259);
nand U11385 (N_11385,N_10695,N_10491);
nand U11386 (N_11386,N_10376,N_10184);
and U11387 (N_11387,N_10962,N_10205);
xor U11388 (N_11388,N_10514,N_10586);
or U11389 (N_11389,N_10004,N_10482);
nand U11390 (N_11390,N_10713,N_10501);
and U11391 (N_11391,N_10104,N_10733);
nand U11392 (N_11392,N_10510,N_10449);
or U11393 (N_11393,N_10842,N_10926);
nand U11394 (N_11394,N_10358,N_10332);
xor U11395 (N_11395,N_10956,N_10345);
nand U11396 (N_11396,N_10067,N_10880);
or U11397 (N_11397,N_10717,N_10049);
nor U11398 (N_11398,N_10837,N_10481);
nor U11399 (N_11399,N_10007,N_10764);
nand U11400 (N_11400,N_10901,N_10198);
or U11401 (N_11401,N_10595,N_10019);
and U11402 (N_11402,N_10720,N_10165);
or U11403 (N_11403,N_10585,N_10589);
xnor U11404 (N_11404,N_10564,N_10469);
nor U11405 (N_11405,N_10236,N_10090);
nand U11406 (N_11406,N_10761,N_10079);
nand U11407 (N_11407,N_10214,N_10115);
nand U11408 (N_11408,N_10187,N_10412);
and U11409 (N_11409,N_10968,N_10337);
and U11410 (N_11410,N_10621,N_10571);
and U11411 (N_11411,N_10896,N_10404);
and U11412 (N_11412,N_10832,N_10252);
and U11413 (N_11413,N_10162,N_10745);
and U11414 (N_11414,N_10992,N_10609);
nand U11415 (N_11415,N_10632,N_10168);
and U11416 (N_11416,N_10261,N_10106);
and U11417 (N_11417,N_10243,N_10005);
nand U11418 (N_11418,N_10177,N_10570);
nand U11419 (N_11419,N_10242,N_10806);
nand U11420 (N_11420,N_10397,N_10022);
nand U11421 (N_11421,N_10593,N_10755);
or U11422 (N_11422,N_10317,N_10371);
xor U11423 (N_11423,N_10664,N_10435);
or U11424 (N_11424,N_10749,N_10359);
and U11425 (N_11425,N_10827,N_10297);
and U11426 (N_11426,N_10040,N_10247);
and U11427 (N_11427,N_10036,N_10552);
nand U11428 (N_11428,N_10525,N_10917);
nor U11429 (N_11429,N_10889,N_10351);
nor U11430 (N_11430,N_10113,N_10650);
nor U11431 (N_11431,N_10947,N_10323);
or U11432 (N_11432,N_10145,N_10655);
or U11433 (N_11433,N_10364,N_10535);
nand U11434 (N_11434,N_10775,N_10285);
nand U11435 (N_11435,N_10846,N_10871);
nand U11436 (N_11436,N_10316,N_10339);
and U11437 (N_11437,N_10111,N_10018);
or U11438 (N_11438,N_10948,N_10767);
nor U11439 (N_11439,N_10959,N_10176);
nor U11440 (N_11440,N_10955,N_10420);
nand U11441 (N_11441,N_10591,N_10831);
nor U11442 (N_11442,N_10885,N_10932);
xnor U11443 (N_11443,N_10250,N_10001);
or U11444 (N_11444,N_10189,N_10276);
and U11445 (N_11445,N_10063,N_10117);
nand U11446 (N_11446,N_10367,N_10329);
nand U11447 (N_11447,N_10390,N_10656);
or U11448 (N_11448,N_10434,N_10039);
or U11449 (N_11449,N_10229,N_10646);
or U11450 (N_11450,N_10762,N_10671);
nor U11451 (N_11451,N_10027,N_10139);
and U11452 (N_11452,N_10776,N_10969);
and U11453 (N_11453,N_10628,N_10729);
nor U11454 (N_11454,N_10441,N_10605);
nor U11455 (N_11455,N_10393,N_10800);
or U11456 (N_11456,N_10129,N_10905);
nor U11457 (N_11457,N_10763,N_10587);
and U11458 (N_11458,N_10909,N_10934);
and U11459 (N_11459,N_10865,N_10078);
or U11460 (N_11460,N_10879,N_10636);
nor U11461 (N_11461,N_10338,N_10446);
nor U11462 (N_11462,N_10608,N_10092);
nand U11463 (N_11463,N_10678,N_10765);
and U11464 (N_11464,N_10540,N_10123);
or U11465 (N_11465,N_10155,N_10966);
xnor U11466 (N_11466,N_10321,N_10447);
nor U11467 (N_11467,N_10163,N_10394);
or U11468 (N_11468,N_10294,N_10714);
and U11469 (N_11469,N_10043,N_10102);
nor U11470 (N_11470,N_10058,N_10239);
xor U11471 (N_11471,N_10667,N_10801);
or U11472 (N_11472,N_10929,N_10613);
and U11473 (N_11473,N_10727,N_10465);
xor U11474 (N_11474,N_10070,N_10914);
xor U11475 (N_11475,N_10335,N_10627);
nand U11476 (N_11476,N_10559,N_10185);
xor U11477 (N_11477,N_10651,N_10916);
nor U11478 (N_11478,N_10970,N_10601);
nor U11479 (N_11479,N_10413,N_10817);
nor U11480 (N_11480,N_10101,N_10375);
nor U11481 (N_11481,N_10863,N_10428);
and U11482 (N_11482,N_10849,N_10480);
nand U11483 (N_11483,N_10757,N_10507);
nand U11484 (N_11484,N_10477,N_10006);
and U11485 (N_11485,N_10427,N_10035);
xnor U11486 (N_11486,N_10550,N_10178);
and U11487 (N_11487,N_10592,N_10475);
and U11488 (N_11488,N_10325,N_10431);
and U11489 (N_11489,N_10531,N_10327);
nor U11490 (N_11490,N_10923,N_10445);
nor U11491 (N_11491,N_10893,N_10368);
nor U11492 (N_11492,N_10852,N_10995);
or U11493 (N_11493,N_10836,N_10722);
nand U11494 (N_11494,N_10804,N_10103);
or U11495 (N_11495,N_10097,N_10751);
xnor U11496 (N_11496,N_10030,N_10026);
nand U11497 (N_11497,N_10234,N_10122);
nor U11498 (N_11498,N_10082,N_10538);
nor U11499 (N_11499,N_10151,N_10736);
nor U11500 (N_11500,N_10336,N_10032);
nor U11501 (N_11501,N_10960,N_10043);
nor U11502 (N_11502,N_10908,N_10668);
and U11503 (N_11503,N_10023,N_10068);
nor U11504 (N_11504,N_10340,N_10101);
xnor U11505 (N_11505,N_10977,N_10332);
nand U11506 (N_11506,N_10684,N_10224);
and U11507 (N_11507,N_10208,N_10745);
xor U11508 (N_11508,N_10654,N_10915);
nand U11509 (N_11509,N_10609,N_10221);
nor U11510 (N_11510,N_10796,N_10453);
or U11511 (N_11511,N_10482,N_10856);
nand U11512 (N_11512,N_10520,N_10363);
or U11513 (N_11513,N_10965,N_10970);
or U11514 (N_11514,N_10524,N_10936);
nand U11515 (N_11515,N_10170,N_10756);
and U11516 (N_11516,N_10974,N_10028);
or U11517 (N_11517,N_10028,N_10203);
nor U11518 (N_11518,N_10482,N_10922);
or U11519 (N_11519,N_10901,N_10220);
nand U11520 (N_11520,N_10134,N_10507);
nand U11521 (N_11521,N_10855,N_10832);
xor U11522 (N_11522,N_10601,N_10038);
or U11523 (N_11523,N_10836,N_10010);
and U11524 (N_11524,N_10065,N_10219);
nor U11525 (N_11525,N_10335,N_10288);
and U11526 (N_11526,N_10895,N_10914);
xor U11527 (N_11527,N_10153,N_10814);
or U11528 (N_11528,N_10208,N_10863);
xnor U11529 (N_11529,N_10349,N_10141);
and U11530 (N_11530,N_10440,N_10678);
nor U11531 (N_11531,N_10086,N_10407);
xor U11532 (N_11532,N_10733,N_10285);
nor U11533 (N_11533,N_10447,N_10362);
nand U11534 (N_11534,N_10341,N_10845);
and U11535 (N_11535,N_10546,N_10908);
xor U11536 (N_11536,N_10443,N_10919);
xnor U11537 (N_11537,N_10940,N_10466);
nor U11538 (N_11538,N_10718,N_10359);
nand U11539 (N_11539,N_10894,N_10197);
and U11540 (N_11540,N_10593,N_10071);
nand U11541 (N_11541,N_10646,N_10388);
and U11542 (N_11542,N_10250,N_10101);
or U11543 (N_11543,N_10293,N_10413);
nor U11544 (N_11544,N_10267,N_10635);
nor U11545 (N_11545,N_10992,N_10099);
and U11546 (N_11546,N_10013,N_10100);
or U11547 (N_11547,N_10187,N_10611);
nor U11548 (N_11548,N_10502,N_10901);
xnor U11549 (N_11549,N_10057,N_10672);
xnor U11550 (N_11550,N_10018,N_10760);
nand U11551 (N_11551,N_10879,N_10288);
and U11552 (N_11552,N_10549,N_10095);
nor U11553 (N_11553,N_10686,N_10145);
xor U11554 (N_11554,N_10384,N_10014);
nor U11555 (N_11555,N_10365,N_10816);
or U11556 (N_11556,N_10473,N_10932);
and U11557 (N_11557,N_10118,N_10563);
nand U11558 (N_11558,N_10180,N_10979);
or U11559 (N_11559,N_10865,N_10197);
xnor U11560 (N_11560,N_10006,N_10279);
or U11561 (N_11561,N_10278,N_10189);
and U11562 (N_11562,N_10198,N_10877);
nor U11563 (N_11563,N_10573,N_10778);
nor U11564 (N_11564,N_10072,N_10031);
xor U11565 (N_11565,N_10192,N_10682);
nand U11566 (N_11566,N_10049,N_10019);
nor U11567 (N_11567,N_10785,N_10971);
nor U11568 (N_11568,N_10981,N_10559);
and U11569 (N_11569,N_10607,N_10546);
or U11570 (N_11570,N_10022,N_10068);
xor U11571 (N_11571,N_10497,N_10259);
nor U11572 (N_11572,N_10089,N_10209);
nor U11573 (N_11573,N_10647,N_10905);
nand U11574 (N_11574,N_10372,N_10912);
or U11575 (N_11575,N_10583,N_10892);
and U11576 (N_11576,N_10586,N_10562);
nand U11577 (N_11577,N_10722,N_10352);
and U11578 (N_11578,N_10779,N_10515);
or U11579 (N_11579,N_10886,N_10358);
or U11580 (N_11580,N_10013,N_10723);
xor U11581 (N_11581,N_10652,N_10806);
nand U11582 (N_11582,N_10698,N_10482);
nand U11583 (N_11583,N_10958,N_10382);
nand U11584 (N_11584,N_10185,N_10285);
nor U11585 (N_11585,N_10992,N_10456);
nand U11586 (N_11586,N_10162,N_10387);
xor U11587 (N_11587,N_10641,N_10459);
or U11588 (N_11588,N_10570,N_10688);
or U11589 (N_11589,N_10158,N_10834);
xor U11590 (N_11590,N_10530,N_10283);
nor U11591 (N_11591,N_10413,N_10644);
nor U11592 (N_11592,N_10794,N_10189);
xor U11593 (N_11593,N_10005,N_10567);
or U11594 (N_11594,N_10007,N_10903);
or U11595 (N_11595,N_10032,N_10559);
nand U11596 (N_11596,N_10961,N_10884);
or U11597 (N_11597,N_10772,N_10926);
and U11598 (N_11598,N_10594,N_10281);
nand U11599 (N_11599,N_10616,N_10858);
and U11600 (N_11600,N_10793,N_10706);
and U11601 (N_11601,N_10701,N_10192);
and U11602 (N_11602,N_10216,N_10858);
or U11603 (N_11603,N_10886,N_10717);
nand U11604 (N_11604,N_10361,N_10543);
nor U11605 (N_11605,N_10937,N_10493);
or U11606 (N_11606,N_10416,N_10304);
nor U11607 (N_11607,N_10233,N_10099);
or U11608 (N_11608,N_10139,N_10435);
nor U11609 (N_11609,N_10178,N_10237);
xnor U11610 (N_11610,N_10934,N_10288);
xor U11611 (N_11611,N_10002,N_10897);
and U11612 (N_11612,N_10783,N_10955);
or U11613 (N_11613,N_10173,N_10253);
nor U11614 (N_11614,N_10021,N_10694);
or U11615 (N_11615,N_10406,N_10482);
nand U11616 (N_11616,N_10901,N_10995);
nand U11617 (N_11617,N_10987,N_10997);
nand U11618 (N_11618,N_10320,N_10486);
or U11619 (N_11619,N_10967,N_10949);
nand U11620 (N_11620,N_10092,N_10002);
nand U11621 (N_11621,N_10740,N_10320);
or U11622 (N_11622,N_10963,N_10006);
or U11623 (N_11623,N_10173,N_10239);
or U11624 (N_11624,N_10725,N_10550);
nor U11625 (N_11625,N_10074,N_10207);
nand U11626 (N_11626,N_10900,N_10786);
or U11627 (N_11627,N_10346,N_10072);
nand U11628 (N_11628,N_10872,N_10416);
xnor U11629 (N_11629,N_10450,N_10540);
or U11630 (N_11630,N_10893,N_10516);
xnor U11631 (N_11631,N_10786,N_10043);
or U11632 (N_11632,N_10858,N_10627);
nand U11633 (N_11633,N_10948,N_10993);
xnor U11634 (N_11634,N_10379,N_10927);
nand U11635 (N_11635,N_10872,N_10469);
nor U11636 (N_11636,N_10506,N_10839);
nand U11637 (N_11637,N_10464,N_10593);
nand U11638 (N_11638,N_10823,N_10214);
nand U11639 (N_11639,N_10681,N_10816);
or U11640 (N_11640,N_10680,N_10320);
nand U11641 (N_11641,N_10560,N_10492);
and U11642 (N_11642,N_10585,N_10282);
or U11643 (N_11643,N_10679,N_10337);
nor U11644 (N_11644,N_10027,N_10640);
or U11645 (N_11645,N_10306,N_10523);
nand U11646 (N_11646,N_10974,N_10287);
nand U11647 (N_11647,N_10869,N_10689);
nor U11648 (N_11648,N_10546,N_10665);
nand U11649 (N_11649,N_10338,N_10067);
and U11650 (N_11650,N_10957,N_10950);
nand U11651 (N_11651,N_10248,N_10840);
and U11652 (N_11652,N_10625,N_10293);
xor U11653 (N_11653,N_10677,N_10940);
or U11654 (N_11654,N_10669,N_10468);
nand U11655 (N_11655,N_10222,N_10818);
and U11656 (N_11656,N_10132,N_10840);
nor U11657 (N_11657,N_10965,N_10374);
or U11658 (N_11658,N_10846,N_10585);
nor U11659 (N_11659,N_10473,N_10984);
and U11660 (N_11660,N_10586,N_10525);
and U11661 (N_11661,N_10006,N_10292);
or U11662 (N_11662,N_10574,N_10641);
or U11663 (N_11663,N_10702,N_10034);
or U11664 (N_11664,N_10978,N_10979);
or U11665 (N_11665,N_10821,N_10168);
or U11666 (N_11666,N_10362,N_10162);
or U11667 (N_11667,N_10299,N_10930);
nor U11668 (N_11668,N_10367,N_10237);
and U11669 (N_11669,N_10543,N_10223);
nand U11670 (N_11670,N_10010,N_10409);
or U11671 (N_11671,N_10247,N_10428);
and U11672 (N_11672,N_10484,N_10014);
nand U11673 (N_11673,N_10620,N_10473);
and U11674 (N_11674,N_10556,N_10734);
and U11675 (N_11675,N_10270,N_10272);
nor U11676 (N_11676,N_10192,N_10233);
nand U11677 (N_11677,N_10852,N_10911);
nor U11678 (N_11678,N_10864,N_10072);
and U11679 (N_11679,N_10504,N_10779);
and U11680 (N_11680,N_10244,N_10277);
or U11681 (N_11681,N_10455,N_10391);
nor U11682 (N_11682,N_10417,N_10687);
nand U11683 (N_11683,N_10304,N_10440);
nor U11684 (N_11684,N_10744,N_10636);
nand U11685 (N_11685,N_10263,N_10525);
and U11686 (N_11686,N_10451,N_10466);
nor U11687 (N_11687,N_10229,N_10823);
nand U11688 (N_11688,N_10538,N_10469);
and U11689 (N_11689,N_10303,N_10412);
and U11690 (N_11690,N_10403,N_10043);
and U11691 (N_11691,N_10532,N_10116);
and U11692 (N_11692,N_10454,N_10016);
and U11693 (N_11693,N_10754,N_10276);
and U11694 (N_11694,N_10154,N_10959);
nor U11695 (N_11695,N_10711,N_10746);
or U11696 (N_11696,N_10527,N_10486);
or U11697 (N_11697,N_10896,N_10011);
or U11698 (N_11698,N_10392,N_10915);
nand U11699 (N_11699,N_10614,N_10379);
and U11700 (N_11700,N_10155,N_10529);
and U11701 (N_11701,N_10346,N_10716);
nand U11702 (N_11702,N_10557,N_10660);
or U11703 (N_11703,N_10772,N_10134);
or U11704 (N_11704,N_10694,N_10118);
nand U11705 (N_11705,N_10695,N_10582);
nor U11706 (N_11706,N_10082,N_10311);
or U11707 (N_11707,N_10326,N_10572);
and U11708 (N_11708,N_10908,N_10765);
nor U11709 (N_11709,N_10158,N_10975);
nor U11710 (N_11710,N_10305,N_10584);
nor U11711 (N_11711,N_10252,N_10019);
or U11712 (N_11712,N_10128,N_10756);
and U11713 (N_11713,N_10952,N_10901);
nand U11714 (N_11714,N_10898,N_10976);
or U11715 (N_11715,N_10034,N_10113);
or U11716 (N_11716,N_10225,N_10298);
nor U11717 (N_11717,N_10055,N_10314);
or U11718 (N_11718,N_10026,N_10813);
and U11719 (N_11719,N_10554,N_10338);
or U11720 (N_11720,N_10795,N_10091);
nor U11721 (N_11721,N_10652,N_10958);
and U11722 (N_11722,N_10611,N_10838);
or U11723 (N_11723,N_10873,N_10028);
and U11724 (N_11724,N_10534,N_10427);
or U11725 (N_11725,N_10982,N_10805);
and U11726 (N_11726,N_10160,N_10049);
nand U11727 (N_11727,N_10935,N_10954);
or U11728 (N_11728,N_10390,N_10669);
nor U11729 (N_11729,N_10926,N_10905);
xnor U11730 (N_11730,N_10064,N_10495);
and U11731 (N_11731,N_10958,N_10857);
or U11732 (N_11732,N_10491,N_10381);
xnor U11733 (N_11733,N_10526,N_10326);
or U11734 (N_11734,N_10060,N_10144);
and U11735 (N_11735,N_10285,N_10375);
and U11736 (N_11736,N_10806,N_10503);
and U11737 (N_11737,N_10669,N_10521);
nand U11738 (N_11738,N_10848,N_10581);
and U11739 (N_11739,N_10390,N_10527);
or U11740 (N_11740,N_10953,N_10983);
or U11741 (N_11741,N_10352,N_10262);
and U11742 (N_11742,N_10097,N_10535);
xor U11743 (N_11743,N_10635,N_10402);
nor U11744 (N_11744,N_10752,N_10686);
nand U11745 (N_11745,N_10050,N_10814);
xnor U11746 (N_11746,N_10626,N_10054);
and U11747 (N_11747,N_10941,N_10377);
nand U11748 (N_11748,N_10176,N_10750);
or U11749 (N_11749,N_10308,N_10941);
xnor U11750 (N_11750,N_10521,N_10067);
nand U11751 (N_11751,N_10758,N_10694);
nor U11752 (N_11752,N_10514,N_10511);
nor U11753 (N_11753,N_10523,N_10533);
or U11754 (N_11754,N_10198,N_10922);
xor U11755 (N_11755,N_10514,N_10304);
and U11756 (N_11756,N_10594,N_10976);
nand U11757 (N_11757,N_10416,N_10804);
or U11758 (N_11758,N_10806,N_10249);
and U11759 (N_11759,N_10695,N_10268);
xnor U11760 (N_11760,N_10852,N_10799);
or U11761 (N_11761,N_10682,N_10559);
nand U11762 (N_11762,N_10330,N_10927);
nand U11763 (N_11763,N_10122,N_10589);
nor U11764 (N_11764,N_10625,N_10107);
and U11765 (N_11765,N_10580,N_10421);
and U11766 (N_11766,N_10053,N_10269);
xnor U11767 (N_11767,N_10152,N_10293);
or U11768 (N_11768,N_10684,N_10819);
nand U11769 (N_11769,N_10651,N_10857);
or U11770 (N_11770,N_10627,N_10778);
and U11771 (N_11771,N_10876,N_10663);
nor U11772 (N_11772,N_10398,N_10932);
nor U11773 (N_11773,N_10450,N_10522);
or U11774 (N_11774,N_10504,N_10739);
and U11775 (N_11775,N_10356,N_10352);
nand U11776 (N_11776,N_10405,N_10527);
or U11777 (N_11777,N_10484,N_10476);
nor U11778 (N_11778,N_10621,N_10451);
nor U11779 (N_11779,N_10039,N_10758);
or U11780 (N_11780,N_10942,N_10378);
and U11781 (N_11781,N_10354,N_10847);
nor U11782 (N_11782,N_10375,N_10886);
nor U11783 (N_11783,N_10301,N_10307);
nor U11784 (N_11784,N_10557,N_10300);
nor U11785 (N_11785,N_10688,N_10803);
nor U11786 (N_11786,N_10165,N_10148);
or U11787 (N_11787,N_10877,N_10871);
nand U11788 (N_11788,N_10464,N_10273);
nand U11789 (N_11789,N_10165,N_10487);
nand U11790 (N_11790,N_10756,N_10437);
xor U11791 (N_11791,N_10709,N_10092);
and U11792 (N_11792,N_10903,N_10146);
and U11793 (N_11793,N_10558,N_10522);
and U11794 (N_11794,N_10570,N_10081);
nor U11795 (N_11795,N_10287,N_10302);
nand U11796 (N_11796,N_10631,N_10413);
nor U11797 (N_11797,N_10338,N_10086);
or U11798 (N_11798,N_10844,N_10095);
or U11799 (N_11799,N_10103,N_10655);
and U11800 (N_11800,N_10096,N_10689);
or U11801 (N_11801,N_10573,N_10510);
nand U11802 (N_11802,N_10356,N_10564);
nand U11803 (N_11803,N_10749,N_10954);
and U11804 (N_11804,N_10260,N_10162);
or U11805 (N_11805,N_10424,N_10716);
xnor U11806 (N_11806,N_10097,N_10905);
nand U11807 (N_11807,N_10875,N_10418);
and U11808 (N_11808,N_10268,N_10726);
and U11809 (N_11809,N_10647,N_10787);
xor U11810 (N_11810,N_10084,N_10187);
or U11811 (N_11811,N_10928,N_10803);
or U11812 (N_11812,N_10044,N_10511);
or U11813 (N_11813,N_10180,N_10109);
and U11814 (N_11814,N_10950,N_10243);
xor U11815 (N_11815,N_10179,N_10571);
nor U11816 (N_11816,N_10971,N_10482);
and U11817 (N_11817,N_10218,N_10061);
or U11818 (N_11818,N_10023,N_10798);
nor U11819 (N_11819,N_10001,N_10559);
xnor U11820 (N_11820,N_10592,N_10552);
and U11821 (N_11821,N_10171,N_10439);
or U11822 (N_11822,N_10007,N_10164);
nor U11823 (N_11823,N_10010,N_10988);
nor U11824 (N_11824,N_10130,N_10838);
and U11825 (N_11825,N_10542,N_10806);
and U11826 (N_11826,N_10263,N_10429);
nand U11827 (N_11827,N_10348,N_10336);
xor U11828 (N_11828,N_10148,N_10400);
nand U11829 (N_11829,N_10206,N_10466);
or U11830 (N_11830,N_10817,N_10177);
or U11831 (N_11831,N_10605,N_10248);
nor U11832 (N_11832,N_10965,N_10380);
or U11833 (N_11833,N_10658,N_10488);
nand U11834 (N_11834,N_10832,N_10968);
or U11835 (N_11835,N_10921,N_10552);
or U11836 (N_11836,N_10190,N_10629);
or U11837 (N_11837,N_10795,N_10021);
nand U11838 (N_11838,N_10140,N_10306);
xnor U11839 (N_11839,N_10050,N_10119);
nor U11840 (N_11840,N_10236,N_10058);
and U11841 (N_11841,N_10886,N_10984);
nor U11842 (N_11842,N_10783,N_10443);
or U11843 (N_11843,N_10371,N_10883);
or U11844 (N_11844,N_10391,N_10437);
and U11845 (N_11845,N_10183,N_10337);
nor U11846 (N_11846,N_10046,N_10614);
or U11847 (N_11847,N_10163,N_10600);
xor U11848 (N_11848,N_10761,N_10170);
or U11849 (N_11849,N_10584,N_10334);
or U11850 (N_11850,N_10321,N_10706);
and U11851 (N_11851,N_10394,N_10657);
xor U11852 (N_11852,N_10939,N_10544);
nor U11853 (N_11853,N_10160,N_10460);
nor U11854 (N_11854,N_10009,N_10386);
and U11855 (N_11855,N_10109,N_10349);
and U11856 (N_11856,N_10513,N_10596);
nor U11857 (N_11857,N_10111,N_10634);
nor U11858 (N_11858,N_10551,N_10864);
nor U11859 (N_11859,N_10259,N_10343);
nand U11860 (N_11860,N_10878,N_10857);
and U11861 (N_11861,N_10491,N_10882);
or U11862 (N_11862,N_10610,N_10960);
nor U11863 (N_11863,N_10790,N_10921);
and U11864 (N_11864,N_10094,N_10723);
or U11865 (N_11865,N_10025,N_10121);
xnor U11866 (N_11866,N_10416,N_10311);
nand U11867 (N_11867,N_10558,N_10901);
and U11868 (N_11868,N_10519,N_10551);
xor U11869 (N_11869,N_10045,N_10512);
and U11870 (N_11870,N_10089,N_10603);
or U11871 (N_11871,N_10275,N_10723);
nand U11872 (N_11872,N_10110,N_10079);
and U11873 (N_11873,N_10207,N_10747);
or U11874 (N_11874,N_10726,N_10161);
nor U11875 (N_11875,N_10429,N_10117);
or U11876 (N_11876,N_10453,N_10356);
nand U11877 (N_11877,N_10156,N_10840);
and U11878 (N_11878,N_10501,N_10482);
or U11879 (N_11879,N_10986,N_10359);
or U11880 (N_11880,N_10109,N_10268);
or U11881 (N_11881,N_10936,N_10907);
and U11882 (N_11882,N_10767,N_10307);
and U11883 (N_11883,N_10831,N_10703);
xnor U11884 (N_11884,N_10701,N_10243);
nor U11885 (N_11885,N_10475,N_10219);
nand U11886 (N_11886,N_10348,N_10738);
or U11887 (N_11887,N_10154,N_10104);
xor U11888 (N_11888,N_10975,N_10912);
nand U11889 (N_11889,N_10433,N_10721);
or U11890 (N_11890,N_10538,N_10608);
nand U11891 (N_11891,N_10900,N_10116);
nand U11892 (N_11892,N_10931,N_10995);
nor U11893 (N_11893,N_10130,N_10049);
nand U11894 (N_11894,N_10016,N_10437);
xor U11895 (N_11895,N_10107,N_10441);
nor U11896 (N_11896,N_10925,N_10354);
or U11897 (N_11897,N_10453,N_10461);
and U11898 (N_11898,N_10119,N_10919);
nand U11899 (N_11899,N_10894,N_10629);
xor U11900 (N_11900,N_10318,N_10312);
and U11901 (N_11901,N_10224,N_10603);
xor U11902 (N_11902,N_10788,N_10109);
or U11903 (N_11903,N_10916,N_10648);
or U11904 (N_11904,N_10611,N_10230);
nand U11905 (N_11905,N_10026,N_10501);
and U11906 (N_11906,N_10880,N_10320);
nor U11907 (N_11907,N_10443,N_10731);
or U11908 (N_11908,N_10313,N_10221);
and U11909 (N_11909,N_10197,N_10519);
nand U11910 (N_11910,N_10940,N_10001);
nor U11911 (N_11911,N_10151,N_10614);
and U11912 (N_11912,N_10255,N_10065);
xnor U11913 (N_11913,N_10398,N_10784);
nor U11914 (N_11914,N_10997,N_10881);
or U11915 (N_11915,N_10822,N_10841);
and U11916 (N_11916,N_10529,N_10468);
nand U11917 (N_11917,N_10051,N_10016);
and U11918 (N_11918,N_10762,N_10048);
or U11919 (N_11919,N_10583,N_10853);
or U11920 (N_11920,N_10783,N_10377);
nand U11921 (N_11921,N_10526,N_10755);
nand U11922 (N_11922,N_10704,N_10957);
and U11923 (N_11923,N_10923,N_10060);
nor U11924 (N_11924,N_10551,N_10675);
nand U11925 (N_11925,N_10251,N_10643);
and U11926 (N_11926,N_10106,N_10275);
or U11927 (N_11927,N_10940,N_10585);
nand U11928 (N_11928,N_10307,N_10318);
nor U11929 (N_11929,N_10019,N_10958);
nand U11930 (N_11930,N_10914,N_10485);
nand U11931 (N_11931,N_10232,N_10095);
or U11932 (N_11932,N_10163,N_10593);
or U11933 (N_11933,N_10139,N_10309);
nand U11934 (N_11934,N_10610,N_10445);
and U11935 (N_11935,N_10617,N_10829);
nor U11936 (N_11936,N_10351,N_10204);
or U11937 (N_11937,N_10869,N_10520);
xnor U11938 (N_11938,N_10955,N_10063);
or U11939 (N_11939,N_10623,N_10822);
nor U11940 (N_11940,N_10164,N_10979);
nand U11941 (N_11941,N_10780,N_10019);
nand U11942 (N_11942,N_10762,N_10506);
and U11943 (N_11943,N_10438,N_10425);
and U11944 (N_11944,N_10101,N_10674);
or U11945 (N_11945,N_10450,N_10657);
nor U11946 (N_11946,N_10073,N_10332);
nand U11947 (N_11947,N_10369,N_10428);
nand U11948 (N_11948,N_10294,N_10006);
and U11949 (N_11949,N_10388,N_10032);
and U11950 (N_11950,N_10967,N_10820);
nand U11951 (N_11951,N_10218,N_10970);
and U11952 (N_11952,N_10090,N_10315);
nand U11953 (N_11953,N_10740,N_10438);
and U11954 (N_11954,N_10987,N_10344);
and U11955 (N_11955,N_10527,N_10764);
and U11956 (N_11956,N_10896,N_10003);
nand U11957 (N_11957,N_10490,N_10380);
xnor U11958 (N_11958,N_10461,N_10520);
or U11959 (N_11959,N_10861,N_10972);
or U11960 (N_11960,N_10585,N_10437);
nand U11961 (N_11961,N_10336,N_10084);
and U11962 (N_11962,N_10222,N_10331);
and U11963 (N_11963,N_10006,N_10082);
nand U11964 (N_11964,N_10333,N_10330);
nor U11965 (N_11965,N_10307,N_10819);
nor U11966 (N_11966,N_10481,N_10166);
and U11967 (N_11967,N_10153,N_10951);
and U11968 (N_11968,N_10144,N_10332);
nand U11969 (N_11969,N_10007,N_10106);
nand U11970 (N_11970,N_10349,N_10173);
nor U11971 (N_11971,N_10439,N_10636);
nand U11972 (N_11972,N_10754,N_10896);
and U11973 (N_11973,N_10827,N_10597);
nand U11974 (N_11974,N_10769,N_10575);
nor U11975 (N_11975,N_10879,N_10389);
nand U11976 (N_11976,N_10204,N_10796);
and U11977 (N_11977,N_10806,N_10877);
nor U11978 (N_11978,N_10754,N_10104);
and U11979 (N_11979,N_10662,N_10415);
nor U11980 (N_11980,N_10269,N_10514);
nor U11981 (N_11981,N_10268,N_10882);
nand U11982 (N_11982,N_10814,N_10049);
nor U11983 (N_11983,N_10752,N_10544);
nand U11984 (N_11984,N_10260,N_10417);
nand U11985 (N_11985,N_10902,N_10755);
nor U11986 (N_11986,N_10134,N_10607);
nand U11987 (N_11987,N_10310,N_10959);
and U11988 (N_11988,N_10067,N_10498);
nand U11989 (N_11989,N_10416,N_10013);
and U11990 (N_11990,N_10682,N_10122);
xnor U11991 (N_11991,N_10673,N_10034);
xnor U11992 (N_11992,N_10983,N_10760);
xor U11993 (N_11993,N_10086,N_10502);
and U11994 (N_11994,N_10253,N_10642);
and U11995 (N_11995,N_10593,N_10372);
nor U11996 (N_11996,N_10768,N_10912);
nor U11997 (N_11997,N_10415,N_10335);
and U11998 (N_11998,N_10998,N_10012);
nand U11999 (N_11999,N_10443,N_10993);
or U12000 (N_12000,N_11280,N_11270);
and U12001 (N_12001,N_11345,N_11307);
or U12002 (N_12002,N_11153,N_11138);
or U12003 (N_12003,N_11976,N_11983);
nor U12004 (N_12004,N_11249,N_11594);
and U12005 (N_12005,N_11628,N_11181);
and U12006 (N_12006,N_11924,N_11819);
and U12007 (N_12007,N_11353,N_11070);
nand U12008 (N_12008,N_11239,N_11788);
nand U12009 (N_12009,N_11855,N_11551);
or U12010 (N_12010,N_11658,N_11154);
and U12011 (N_12011,N_11679,N_11985);
or U12012 (N_12012,N_11751,N_11499);
nand U12013 (N_12013,N_11742,N_11415);
or U12014 (N_12014,N_11895,N_11540);
and U12015 (N_12015,N_11907,N_11338);
nor U12016 (N_12016,N_11969,N_11407);
and U12017 (N_12017,N_11753,N_11128);
nand U12018 (N_12018,N_11467,N_11501);
and U12019 (N_12019,N_11411,N_11906);
or U12020 (N_12020,N_11885,N_11636);
nand U12021 (N_12021,N_11965,N_11329);
xor U12022 (N_12022,N_11993,N_11062);
and U12023 (N_12023,N_11774,N_11979);
nand U12024 (N_12024,N_11419,N_11172);
or U12025 (N_12025,N_11066,N_11022);
or U12026 (N_12026,N_11146,N_11815);
and U12027 (N_12027,N_11363,N_11629);
and U12028 (N_12028,N_11260,N_11165);
nand U12029 (N_12029,N_11125,N_11425);
nand U12030 (N_12030,N_11643,N_11040);
and U12031 (N_12031,N_11454,N_11246);
or U12032 (N_12032,N_11770,N_11341);
or U12033 (N_12033,N_11945,N_11401);
or U12034 (N_12034,N_11392,N_11351);
nand U12035 (N_12035,N_11515,N_11087);
nor U12036 (N_12036,N_11360,N_11216);
nand U12037 (N_12037,N_11612,N_11178);
xor U12038 (N_12038,N_11273,N_11086);
nand U12039 (N_12039,N_11681,N_11859);
nor U12040 (N_12040,N_11553,N_11211);
nand U12041 (N_12041,N_11085,N_11452);
nor U12042 (N_12042,N_11673,N_11768);
nor U12043 (N_12043,N_11994,N_11131);
and U12044 (N_12044,N_11269,N_11804);
xnor U12045 (N_12045,N_11206,N_11265);
nor U12046 (N_12046,N_11496,N_11326);
nand U12047 (N_12047,N_11910,N_11771);
and U12048 (N_12048,N_11013,N_11074);
xnor U12049 (N_12049,N_11990,N_11237);
xnor U12050 (N_12050,N_11310,N_11010);
and U12051 (N_12051,N_11978,N_11562);
xor U12052 (N_12052,N_11161,N_11757);
and U12053 (N_12053,N_11591,N_11396);
nand U12054 (N_12054,N_11572,N_11448);
and U12055 (N_12055,N_11199,N_11687);
nor U12056 (N_12056,N_11937,N_11881);
or U12057 (N_12057,N_11932,N_11397);
nor U12058 (N_12058,N_11322,N_11939);
nor U12059 (N_12059,N_11710,N_11474);
nor U12060 (N_12060,N_11299,N_11527);
or U12061 (N_12061,N_11221,N_11662);
or U12062 (N_12062,N_11245,N_11680);
or U12063 (N_12063,N_11488,N_11656);
or U12064 (N_12064,N_11294,N_11110);
and U12065 (N_12065,N_11974,N_11330);
xor U12066 (N_12066,N_11860,N_11875);
and U12067 (N_12067,N_11535,N_11514);
nand U12068 (N_12068,N_11275,N_11465);
and U12069 (N_12069,N_11166,N_11695);
or U12070 (N_12070,N_11926,N_11697);
or U12071 (N_12071,N_11852,N_11913);
and U12072 (N_12072,N_11879,N_11113);
nand U12073 (N_12073,N_11352,N_11207);
nand U12074 (N_12074,N_11257,N_11533);
nand U12075 (N_12075,N_11334,N_11579);
nand U12076 (N_12076,N_11048,N_11648);
nor U12077 (N_12077,N_11082,N_11016);
nand U12078 (N_12078,N_11293,N_11682);
nor U12079 (N_12079,N_11876,N_11405);
nor U12080 (N_12080,N_11067,N_11858);
nand U12081 (N_12081,N_11603,N_11027);
nor U12082 (N_12082,N_11132,N_11383);
and U12083 (N_12083,N_11469,N_11263);
xnor U12084 (N_12084,N_11343,N_11930);
or U12085 (N_12085,N_11163,N_11668);
and U12086 (N_12086,N_11830,N_11970);
xnor U12087 (N_12087,N_11327,N_11626);
or U12088 (N_12088,N_11418,N_11268);
nor U12089 (N_12089,N_11012,N_11162);
nor U12090 (N_12090,N_11802,N_11144);
or U12091 (N_12091,N_11999,N_11038);
xnor U12092 (N_12092,N_11095,N_11491);
or U12093 (N_12093,N_11349,N_11051);
nor U12094 (N_12094,N_11851,N_11692);
nor U12095 (N_12095,N_11960,N_11843);
or U12096 (N_12096,N_11097,N_11856);
or U12097 (N_12097,N_11957,N_11791);
nand U12098 (N_12098,N_11641,N_11135);
nor U12099 (N_12099,N_11309,N_11602);
nor U12100 (N_12100,N_11529,N_11019);
or U12101 (N_12101,N_11702,N_11799);
and U12102 (N_12102,N_11714,N_11773);
xnor U12103 (N_12103,N_11043,N_11244);
nor U12104 (N_12104,N_11124,N_11672);
nand U12105 (N_12105,N_11996,N_11568);
nor U12106 (N_12106,N_11348,N_11020);
or U12107 (N_12107,N_11731,N_11919);
nand U12108 (N_12108,N_11690,N_11729);
or U12109 (N_12109,N_11498,N_11747);
or U12110 (N_12110,N_11475,N_11615);
nand U12111 (N_12111,N_11806,N_11453);
nor U12112 (N_12112,N_11115,N_11992);
nand U12113 (N_12113,N_11639,N_11718);
or U12114 (N_12114,N_11549,N_11402);
xnor U12115 (N_12115,N_11505,N_11223);
nor U12116 (N_12116,N_11964,N_11446);
nor U12117 (N_12117,N_11151,N_11597);
nand U12118 (N_12118,N_11367,N_11109);
or U12119 (N_12119,N_11266,N_11106);
or U12120 (N_12120,N_11738,N_11732);
nand U12121 (N_12121,N_11767,N_11112);
nor U12122 (N_12122,N_11473,N_11780);
and U12123 (N_12123,N_11743,N_11476);
xnor U12124 (N_12124,N_11179,N_11736);
nor U12125 (N_12125,N_11619,N_11377);
and U12126 (N_12126,N_11104,N_11640);
and U12127 (N_12127,N_11036,N_11357);
nor U12128 (N_12128,N_11160,N_11882);
and U12129 (N_12129,N_11633,N_11844);
nand U12130 (N_12130,N_11061,N_11230);
and U12131 (N_12131,N_11520,N_11604);
nor U12132 (N_12132,N_11008,N_11229);
or U12133 (N_12133,N_11684,N_11168);
and U12134 (N_12134,N_11586,N_11167);
xnor U12135 (N_12135,N_11493,N_11644);
and U12136 (N_12136,N_11909,N_11721);
and U12137 (N_12137,N_11554,N_11441);
xnor U12138 (N_12138,N_11877,N_11653);
nand U12139 (N_12139,N_11276,N_11521);
nor U12140 (N_12140,N_11754,N_11796);
or U12141 (N_12141,N_11561,N_11864);
and U12142 (N_12142,N_11252,N_11047);
nand U12143 (N_12143,N_11158,N_11611);
and U12144 (N_12144,N_11825,N_11836);
or U12145 (N_12145,N_11795,N_11409);
and U12146 (N_12146,N_11443,N_11803);
and U12147 (N_12147,N_11234,N_11194);
nor U12148 (N_12148,N_11948,N_11364);
or U12149 (N_12149,N_11955,N_11426);
and U12150 (N_12150,N_11532,N_11676);
nand U12151 (N_12151,N_11437,N_11581);
or U12152 (N_12152,N_11901,N_11408);
and U12153 (N_12153,N_11654,N_11840);
nand U12154 (N_12154,N_11198,N_11526);
or U12155 (N_12155,N_11625,N_11725);
nor U12156 (N_12156,N_11421,N_11623);
and U12157 (N_12157,N_11787,N_11386);
xnor U12158 (N_12158,N_11622,N_11318);
or U12159 (N_12159,N_11776,N_11610);
and U12160 (N_12160,N_11057,N_11588);
or U12161 (N_12161,N_11303,N_11538);
nand U12162 (N_12162,N_11235,N_11140);
and U12163 (N_12163,N_11490,N_11204);
nand U12164 (N_12164,N_11321,N_11410);
or U12165 (N_12165,N_11102,N_11456);
nand U12166 (N_12166,N_11305,N_11018);
or U12167 (N_12167,N_11297,N_11208);
or U12168 (N_12168,N_11155,N_11037);
and U12169 (N_12169,N_11118,N_11370);
and U12170 (N_12170,N_11247,N_11404);
nor U12171 (N_12171,N_11482,N_11314);
nand U12172 (N_12172,N_11534,N_11372);
nand U12173 (N_12173,N_11897,N_11923);
nand U12174 (N_12174,N_11192,N_11031);
and U12175 (N_12175,N_11059,N_11849);
nand U12176 (N_12176,N_11122,N_11722);
nor U12177 (N_12177,N_11671,N_11232);
or U12178 (N_12178,N_11479,N_11333);
nand U12179 (N_12179,N_11558,N_11621);
or U12180 (N_12180,N_11084,N_11214);
and U12181 (N_12181,N_11762,N_11583);
and U12182 (N_12182,N_11393,N_11902);
xnor U12183 (N_12183,N_11137,N_11045);
nand U12184 (N_12184,N_11899,N_11127);
xor U12185 (N_12185,N_11947,N_11060);
nor U12186 (N_12186,N_11005,N_11915);
xnor U12187 (N_12187,N_11962,N_11986);
and U12188 (N_12188,N_11449,N_11023);
nand U12189 (N_12189,N_11734,N_11777);
nand U12190 (N_12190,N_11891,N_11114);
nor U12191 (N_12191,N_11359,N_11500);
nor U12192 (N_12192,N_11099,N_11093);
and U12193 (N_12193,N_11203,N_11740);
nand U12194 (N_12194,N_11279,N_11361);
nor U12195 (N_12195,N_11958,N_11820);
nand U12196 (N_12196,N_11451,N_11388);
nor U12197 (N_12197,N_11989,N_11865);
or U12198 (N_12198,N_11209,N_11130);
nor U12199 (N_12199,N_11248,N_11991);
or U12200 (N_12200,N_11033,N_11831);
nand U12201 (N_12201,N_11756,N_11778);
nor U12202 (N_12202,N_11014,N_11143);
nor U12203 (N_12203,N_11863,N_11139);
nor U12204 (N_12204,N_11355,N_11755);
or U12205 (N_12205,N_11560,N_11760);
nor U12206 (N_12206,N_11427,N_11946);
nor U12207 (N_12207,N_11555,N_11175);
or U12208 (N_12208,N_11703,N_11298);
nand U12209 (N_12209,N_11723,N_11267);
nand U12210 (N_12210,N_11727,N_11282);
and U12211 (N_12211,N_11142,N_11240);
nand U12212 (N_12212,N_11317,N_11184);
xnor U12213 (N_12213,N_11065,N_11068);
or U12214 (N_12214,N_11977,N_11663);
nand U12215 (N_12215,N_11601,N_11661);
or U12216 (N_12216,N_11458,N_11101);
nand U12217 (N_12217,N_11650,N_11573);
nor U12218 (N_12218,N_11984,N_11107);
and U12219 (N_12219,N_11278,N_11342);
nor U12220 (N_12220,N_11624,N_11570);
nand U12221 (N_12221,N_11966,N_11485);
and U12222 (N_12222,N_11823,N_11460);
nand U12223 (N_12223,N_11814,N_11827);
or U12224 (N_12224,N_11608,N_11696);
and U12225 (N_12225,N_11828,N_11116);
nand U12226 (N_12226,N_11935,N_11508);
and U12227 (N_12227,N_11373,N_11903);
or U12228 (N_12228,N_11700,N_11871);
nor U12229 (N_12229,N_11631,N_11786);
and U12230 (N_12230,N_11320,N_11949);
nand U12231 (N_12231,N_11442,N_11536);
nand U12232 (N_12232,N_11195,N_11953);
nand U12233 (N_12233,N_11782,N_11444);
nor U12234 (N_12234,N_11222,N_11685);
nor U12235 (N_12235,N_11741,N_11848);
or U12236 (N_12236,N_11826,N_11869);
or U12237 (N_12237,N_11041,N_11436);
nor U12238 (N_12238,N_11704,N_11489);
xor U12239 (N_12239,N_11921,N_11484);
nor U12240 (N_12240,N_11147,N_11792);
nor U12241 (N_12241,N_11789,N_11413);
nor U12242 (N_12242,N_11646,N_11873);
and U12243 (N_12243,N_11942,N_11618);
nor U12244 (N_12244,N_11987,N_11693);
or U12245 (N_12245,N_11576,N_11470);
or U12246 (N_12246,N_11657,N_11867);
or U12247 (N_12247,N_11034,N_11566);
nor U12248 (N_12248,N_11286,N_11254);
or U12249 (N_12249,N_11652,N_11081);
nor U12250 (N_12250,N_11001,N_11794);
and U12251 (N_12251,N_11250,N_11914);
nand U12252 (N_12252,N_11241,N_11103);
and U12253 (N_12253,N_11670,N_11660);
or U12254 (N_12254,N_11528,N_11548);
nor U12255 (N_12255,N_11758,N_11834);
or U12256 (N_12256,N_11052,N_11546);
nor U12257 (N_12257,N_11801,N_11304);
or U12258 (N_12258,N_11956,N_11088);
and U12259 (N_12259,N_11379,N_11287);
nor U12260 (N_12260,N_11542,N_11258);
and U12261 (N_12261,N_11649,N_11228);
or U12262 (N_12262,N_11417,N_11918);
nor U12263 (N_12263,N_11609,N_11455);
nor U12264 (N_12264,N_11678,N_11145);
nand U12265 (N_12265,N_11308,N_11567);
and U12266 (N_12266,N_11212,N_11058);
nor U12267 (N_12267,N_11375,N_11193);
or U12268 (N_12268,N_11032,N_11210);
nand U12269 (N_12269,N_11749,N_11183);
or U12270 (N_12270,N_11620,N_11800);
nor U12271 (N_12271,N_11177,N_11761);
nor U12272 (N_12272,N_11638,N_11812);
or U12273 (N_12273,N_11733,N_11766);
nor U12274 (N_12274,N_11784,N_11922);
or U12275 (N_12275,N_11481,N_11912);
and U12276 (N_12276,N_11691,N_11707);
nand U12277 (N_12277,N_11466,N_11988);
nor U12278 (N_12278,N_11251,N_11366);
or U12279 (N_12279,N_11226,N_11078);
nor U12280 (N_12280,N_11659,N_11862);
nor U12281 (N_12281,N_11024,N_11705);
and U12282 (N_12282,N_11215,N_11929);
or U12283 (N_12283,N_11666,N_11328);
nor U12284 (N_12284,N_11972,N_11272);
xor U12285 (N_12285,N_11587,N_11339);
and U12286 (N_12286,N_11893,N_11589);
nand U12287 (N_12287,N_11100,N_11995);
xor U12288 (N_12288,N_11874,N_11645);
nor U12289 (N_12289,N_11035,N_11471);
xor U12290 (N_12290,N_11963,N_11430);
nand U12291 (N_12291,N_11423,N_11717);
or U12292 (N_12292,N_11315,N_11982);
and U12293 (N_12293,N_11007,N_11055);
or U12294 (N_12294,N_11483,N_11818);
nor U12295 (N_12295,N_11369,N_11026);
or U12296 (N_12296,N_11651,N_11518);
or U12297 (N_12297,N_11565,N_11406);
or U12298 (N_12298,N_11332,N_11675);
and U12299 (N_12299,N_11811,N_11870);
or U12300 (N_12300,N_11997,N_11044);
xor U12301 (N_12301,N_11677,N_11916);
and U12302 (N_12302,N_11389,N_11706);
and U12303 (N_12303,N_11574,N_11779);
and U12304 (N_12304,N_11709,N_11575);
or U12305 (N_12305,N_11191,N_11072);
nor U12306 (N_12306,N_11472,N_11121);
or U12307 (N_12307,N_11447,N_11627);
nand U12308 (N_12308,N_11399,N_11853);
xnor U12309 (N_12309,N_11746,N_11769);
nor U12310 (N_12310,N_11905,N_11892);
nor U12311 (N_12311,N_11480,N_11564);
or U12312 (N_12312,N_11728,N_11711);
xor U12313 (N_12313,N_11238,N_11213);
or U12314 (N_12314,N_11790,N_11635);
and U12315 (N_12315,N_11846,N_11069);
or U12316 (N_12316,N_11833,N_11941);
and U12317 (N_12317,N_11096,N_11150);
nor U12318 (N_12318,N_11908,N_11391);
nand U12319 (N_12319,N_11841,N_11952);
nand U12320 (N_12320,N_11530,N_11816);
or U12321 (N_12321,N_11416,N_11487);
nand U12322 (N_12322,N_11464,N_11126);
or U12323 (N_12323,N_11559,N_11255);
nor U12324 (N_12324,N_11699,N_11285);
nand U12325 (N_12325,N_11933,N_11477);
xor U12326 (N_12326,N_11319,N_11064);
nand U12327 (N_12327,N_11356,N_11236);
and U12328 (N_12328,N_11003,N_11630);
nand U12329 (N_12329,N_11450,N_11382);
or U12330 (N_12330,N_11689,N_11009);
or U12331 (N_12331,N_11400,N_11385);
or U12332 (N_12332,N_11494,N_11614);
or U12333 (N_12333,N_11073,N_11950);
nand U12334 (N_12334,N_11688,N_11744);
nor U12335 (N_12335,N_11764,N_11911);
and U12336 (N_12336,N_11547,N_11539);
nand U12337 (N_12337,N_11847,N_11311);
xor U12338 (N_12338,N_11667,N_11585);
or U12339 (N_12339,N_11463,N_11878);
xor U12340 (N_12340,N_11004,N_11091);
and U12341 (N_12341,N_11961,N_11613);
xor U12342 (N_12342,N_11745,N_11599);
and U12343 (N_12343,N_11224,N_11089);
or U12344 (N_12344,N_11716,N_11071);
nor U12345 (N_12345,N_11256,N_11056);
and U12346 (N_12346,N_11511,N_11698);
and U12347 (N_12347,N_11136,N_11435);
or U12348 (N_12348,N_11092,N_11510);
nand U12349 (N_12349,N_11340,N_11550);
and U12350 (N_12350,N_11080,N_11832);
and U12351 (N_12351,N_11159,N_11824);
nand U12352 (N_12352,N_11381,N_11387);
and U12353 (N_12353,N_11884,N_11557);
nand U12354 (N_12354,N_11938,N_11927);
or U12355 (N_12355,N_11967,N_11164);
or U12356 (N_12356,N_11325,N_11459);
or U12357 (N_12357,N_11148,N_11712);
or U12358 (N_12358,N_11959,N_11556);
nor U12359 (N_12359,N_11805,N_11261);
or U12360 (N_12360,N_11701,N_11750);
nand U12361 (N_12361,N_11394,N_11998);
nand U12362 (N_12362,N_11243,N_11457);
nand U12363 (N_12363,N_11578,N_11323);
or U12364 (N_12364,N_11513,N_11607);
and U12365 (N_12365,N_11497,N_11936);
or U12366 (N_12366,N_11049,N_11202);
nor U12367 (N_12367,N_11171,N_11686);
and U12368 (N_12368,N_11904,N_11719);
and U12369 (N_12369,N_11253,N_11951);
or U12370 (N_12370,N_11015,N_11291);
nor U12371 (N_12371,N_11544,N_11090);
or U12372 (N_12372,N_11822,N_11980);
nand U12373 (N_12373,N_11420,N_11170);
or U12374 (N_12374,N_11523,N_11344);
or U12375 (N_12375,N_11123,N_11384);
nand U12376 (N_12376,N_11708,N_11200);
nand U12377 (N_12377,N_11083,N_11461);
and U12378 (N_12378,N_11730,N_11775);
or U12379 (N_12379,N_11872,N_11726);
or U12380 (N_12380,N_11288,N_11492);
xnor U12381 (N_12381,N_11346,N_11880);
nand U12382 (N_12382,N_11813,N_11900);
and U12383 (N_12383,N_11182,N_11358);
nand U12384 (N_12384,N_11647,N_11478);
and U12385 (N_12385,N_11785,N_11866);
and U12386 (N_12386,N_11502,N_11105);
nor U12387 (N_12387,N_11205,N_11075);
nor U12388 (N_12388,N_11808,N_11039);
nand U12389 (N_12389,N_11854,N_11889);
and U12390 (N_12390,N_11331,N_11694);
nor U12391 (N_12391,N_11188,N_11119);
nor U12392 (N_12392,N_11462,N_11301);
nand U12393 (N_12393,N_11220,N_11185);
nand U12394 (N_12394,N_11522,N_11431);
and U12395 (N_12395,N_11063,N_11337);
nand U12396 (N_12396,N_11887,N_11324);
or U12397 (N_12397,N_11735,N_11362);
nor U12398 (N_12398,N_11495,N_11403);
and U12399 (N_12399,N_11829,N_11422);
or U12400 (N_12400,N_11002,N_11664);
nand U12401 (N_12401,N_11637,N_11940);
or U12402 (N_12402,N_11595,N_11414);
or U12403 (N_12403,N_11634,N_11981);
or U12404 (N_12404,N_11186,N_11504);
nand U12405 (N_12405,N_11503,N_11720);
or U12406 (N_12406,N_11517,N_11316);
nor U12407 (N_12407,N_11445,N_11217);
nor U12408 (N_12408,N_11837,N_11398);
and U12409 (N_12409,N_11748,N_11606);
nor U12410 (N_12410,N_11157,N_11537);
xor U12411 (N_12411,N_11809,N_11295);
and U12412 (N_12412,N_11302,N_11134);
nor U12413 (N_12413,N_11374,N_11772);
xnor U12414 (N_12414,N_11225,N_11531);
or U12415 (N_12415,N_11838,N_11152);
and U12416 (N_12416,N_11187,N_11354);
and U12417 (N_12417,N_11582,N_11262);
or U12418 (N_12418,N_11079,N_11281);
nand U12419 (N_12419,N_11973,N_11077);
and U12420 (N_12420,N_11412,N_11429);
nand U12421 (N_12421,N_11842,N_11543);
nor U12422 (N_12422,N_11292,N_11798);
xnor U12423 (N_12423,N_11046,N_11390);
nand U12424 (N_12424,N_11665,N_11098);
nand U12425 (N_12425,N_11428,N_11432);
or U12426 (N_12426,N_11593,N_11141);
xnor U12427 (N_12427,N_11605,N_11617);
nor U12428 (N_12428,N_11076,N_11817);
or U12429 (N_12429,N_11928,N_11218);
nor U12430 (N_12430,N_11934,N_11563);
and U12431 (N_12431,N_11433,N_11283);
nand U12432 (N_12432,N_11029,N_11053);
nand U12433 (N_12433,N_11810,N_11845);
xor U12434 (N_12434,N_11737,N_11509);
and U12435 (N_12435,N_11516,N_11507);
and U12436 (N_12436,N_11821,N_11380);
nand U12437 (N_12437,N_11108,N_11642);
xnor U12438 (N_12438,N_11486,N_11368);
nor U12439 (N_12439,N_11189,N_11888);
nand U12440 (N_12440,N_11440,N_11021);
or U12441 (N_12441,N_11264,N_11219);
or U12442 (N_12442,N_11883,N_11600);
and U12443 (N_12443,N_11632,N_11519);
nor U12444 (N_12444,N_11971,N_11017);
or U12445 (N_12445,N_11752,N_11030);
nand U12446 (N_12446,N_11111,N_11577);
and U12447 (N_12447,N_11336,N_11506);
xor U12448 (N_12448,N_11149,N_11839);
nor U12449 (N_12449,N_11190,N_11028);
nor U12450 (N_12450,N_11284,N_11376);
nor U12451 (N_12451,N_11468,N_11715);
and U12452 (N_12452,N_11054,N_11042);
and U12453 (N_12453,N_11196,N_11350);
xnor U12454 (N_12454,N_11571,N_11365);
nand U12455 (N_12455,N_11835,N_11120);
or U12456 (N_12456,N_11590,N_11584);
and U12457 (N_12457,N_11674,N_11156);
nor U12458 (N_12458,N_11920,N_11783);
or U12459 (N_12459,N_11765,N_11724);
xor U12460 (N_12460,N_11763,N_11797);
nor U12461 (N_12461,N_11850,N_11006);
xor U12462 (N_12462,N_11335,N_11395);
nor U12463 (N_12463,N_11424,N_11176);
nand U12464 (N_12464,N_11868,N_11655);
xnor U12465 (N_12465,N_11306,N_11857);
nor U12466 (N_12466,N_11174,N_11592);
or U12467 (N_12467,N_11434,N_11347);
nand U12468 (N_12468,N_11886,N_11598);
nand U12469 (N_12469,N_11050,N_11201);
or U12470 (N_12470,N_11117,N_11289);
or U12471 (N_12471,N_11669,N_11944);
nand U12472 (N_12472,N_11133,N_11898);
or U12473 (N_12473,N_11683,N_11524);
or U12474 (N_12474,N_11231,N_11438);
or U12475 (N_12475,N_11277,N_11313);
nor U12476 (N_12476,N_11233,N_11439);
or U12477 (N_12477,N_11296,N_11000);
or U12478 (N_12478,N_11545,N_11807);
nor U12479 (N_12479,N_11371,N_11861);
and U12480 (N_12480,N_11274,N_11169);
or U12481 (N_12481,N_11890,N_11312);
and U12482 (N_12482,N_11242,N_11781);
or U12483 (N_12483,N_11569,N_11793);
nand U12484 (N_12484,N_11943,N_11917);
or U12485 (N_12485,N_11025,N_11129);
and U12486 (N_12486,N_11896,N_11552);
and U12487 (N_12487,N_11378,N_11925);
and U12488 (N_12488,N_11290,N_11271);
and U12489 (N_12489,N_11894,N_11975);
nor U12490 (N_12490,N_11759,N_11968);
nor U12491 (N_12491,N_11525,N_11931);
or U12492 (N_12492,N_11173,N_11094);
xnor U12493 (N_12493,N_11713,N_11596);
nand U12494 (N_12494,N_11227,N_11580);
xor U12495 (N_12495,N_11180,N_11541);
or U12496 (N_12496,N_11300,N_11197);
or U12497 (N_12497,N_11616,N_11739);
nand U12498 (N_12498,N_11011,N_11259);
and U12499 (N_12499,N_11954,N_11512);
or U12500 (N_12500,N_11646,N_11163);
nor U12501 (N_12501,N_11529,N_11909);
xnor U12502 (N_12502,N_11041,N_11235);
and U12503 (N_12503,N_11892,N_11055);
nor U12504 (N_12504,N_11236,N_11511);
and U12505 (N_12505,N_11849,N_11819);
xor U12506 (N_12506,N_11894,N_11829);
nor U12507 (N_12507,N_11441,N_11772);
and U12508 (N_12508,N_11691,N_11475);
and U12509 (N_12509,N_11860,N_11995);
and U12510 (N_12510,N_11185,N_11408);
nor U12511 (N_12511,N_11703,N_11280);
nand U12512 (N_12512,N_11351,N_11434);
nor U12513 (N_12513,N_11167,N_11934);
nor U12514 (N_12514,N_11736,N_11684);
xor U12515 (N_12515,N_11619,N_11284);
and U12516 (N_12516,N_11377,N_11851);
nor U12517 (N_12517,N_11690,N_11309);
nand U12518 (N_12518,N_11740,N_11385);
nand U12519 (N_12519,N_11533,N_11048);
nor U12520 (N_12520,N_11653,N_11564);
nand U12521 (N_12521,N_11287,N_11630);
or U12522 (N_12522,N_11188,N_11651);
and U12523 (N_12523,N_11797,N_11471);
or U12524 (N_12524,N_11015,N_11731);
and U12525 (N_12525,N_11759,N_11381);
or U12526 (N_12526,N_11377,N_11762);
nand U12527 (N_12527,N_11571,N_11034);
nand U12528 (N_12528,N_11166,N_11853);
nor U12529 (N_12529,N_11014,N_11994);
nand U12530 (N_12530,N_11015,N_11377);
xnor U12531 (N_12531,N_11764,N_11127);
or U12532 (N_12532,N_11974,N_11647);
nand U12533 (N_12533,N_11553,N_11903);
or U12534 (N_12534,N_11818,N_11386);
and U12535 (N_12535,N_11141,N_11616);
and U12536 (N_12536,N_11939,N_11185);
nor U12537 (N_12537,N_11986,N_11628);
nand U12538 (N_12538,N_11724,N_11441);
nand U12539 (N_12539,N_11624,N_11714);
or U12540 (N_12540,N_11805,N_11073);
and U12541 (N_12541,N_11000,N_11108);
or U12542 (N_12542,N_11039,N_11085);
xor U12543 (N_12543,N_11949,N_11709);
nand U12544 (N_12544,N_11573,N_11497);
or U12545 (N_12545,N_11939,N_11031);
nor U12546 (N_12546,N_11212,N_11369);
and U12547 (N_12547,N_11622,N_11641);
or U12548 (N_12548,N_11228,N_11732);
and U12549 (N_12549,N_11526,N_11639);
or U12550 (N_12550,N_11035,N_11252);
nand U12551 (N_12551,N_11541,N_11596);
or U12552 (N_12552,N_11882,N_11215);
or U12553 (N_12553,N_11708,N_11543);
nor U12554 (N_12554,N_11633,N_11379);
nand U12555 (N_12555,N_11368,N_11683);
and U12556 (N_12556,N_11614,N_11542);
or U12557 (N_12557,N_11511,N_11054);
or U12558 (N_12558,N_11249,N_11145);
nand U12559 (N_12559,N_11286,N_11731);
nand U12560 (N_12560,N_11471,N_11435);
or U12561 (N_12561,N_11224,N_11800);
or U12562 (N_12562,N_11904,N_11691);
nand U12563 (N_12563,N_11003,N_11508);
xor U12564 (N_12564,N_11143,N_11083);
or U12565 (N_12565,N_11056,N_11947);
nor U12566 (N_12566,N_11681,N_11917);
or U12567 (N_12567,N_11077,N_11645);
and U12568 (N_12568,N_11873,N_11303);
nand U12569 (N_12569,N_11404,N_11243);
or U12570 (N_12570,N_11020,N_11159);
and U12571 (N_12571,N_11414,N_11279);
nor U12572 (N_12572,N_11602,N_11499);
nand U12573 (N_12573,N_11966,N_11529);
nor U12574 (N_12574,N_11850,N_11359);
and U12575 (N_12575,N_11356,N_11713);
nor U12576 (N_12576,N_11936,N_11399);
and U12577 (N_12577,N_11779,N_11076);
nor U12578 (N_12578,N_11907,N_11529);
and U12579 (N_12579,N_11721,N_11522);
nor U12580 (N_12580,N_11921,N_11183);
or U12581 (N_12581,N_11845,N_11186);
and U12582 (N_12582,N_11431,N_11806);
and U12583 (N_12583,N_11195,N_11842);
or U12584 (N_12584,N_11494,N_11668);
nand U12585 (N_12585,N_11476,N_11731);
or U12586 (N_12586,N_11439,N_11755);
nand U12587 (N_12587,N_11356,N_11390);
or U12588 (N_12588,N_11719,N_11551);
and U12589 (N_12589,N_11805,N_11934);
xor U12590 (N_12590,N_11794,N_11760);
and U12591 (N_12591,N_11597,N_11308);
nor U12592 (N_12592,N_11452,N_11340);
nor U12593 (N_12593,N_11099,N_11247);
nand U12594 (N_12594,N_11271,N_11015);
and U12595 (N_12595,N_11635,N_11842);
and U12596 (N_12596,N_11606,N_11395);
nand U12597 (N_12597,N_11178,N_11553);
nand U12598 (N_12598,N_11968,N_11793);
or U12599 (N_12599,N_11445,N_11562);
and U12600 (N_12600,N_11278,N_11085);
xnor U12601 (N_12601,N_11495,N_11292);
nand U12602 (N_12602,N_11209,N_11224);
or U12603 (N_12603,N_11009,N_11579);
or U12604 (N_12604,N_11545,N_11922);
and U12605 (N_12605,N_11256,N_11909);
nand U12606 (N_12606,N_11923,N_11149);
and U12607 (N_12607,N_11423,N_11735);
or U12608 (N_12608,N_11274,N_11117);
and U12609 (N_12609,N_11267,N_11766);
xnor U12610 (N_12610,N_11607,N_11307);
or U12611 (N_12611,N_11038,N_11955);
and U12612 (N_12612,N_11257,N_11585);
or U12613 (N_12613,N_11762,N_11553);
nor U12614 (N_12614,N_11619,N_11707);
nand U12615 (N_12615,N_11176,N_11074);
nand U12616 (N_12616,N_11823,N_11874);
nand U12617 (N_12617,N_11997,N_11289);
nor U12618 (N_12618,N_11940,N_11041);
nor U12619 (N_12619,N_11000,N_11812);
xnor U12620 (N_12620,N_11712,N_11280);
or U12621 (N_12621,N_11831,N_11246);
or U12622 (N_12622,N_11538,N_11865);
and U12623 (N_12623,N_11040,N_11508);
nor U12624 (N_12624,N_11446,N_11426);
or U12625 (N_12625,N_11490,N_11010);
and U12626 (N_12626,N_11509,N_11099);
nand U12627 (N_12627,N_11470,N_11751);
or U12628 (N_12628,N_11099,N_11179);
and U12629 (N_12629,N_11627,N_11821);
and U12630 (N_12630,N_11708,N_11454);
or U12631 (N_12631,N_11083,N_11978);
or U12632 (N_12632,N_11426,N_11445);
or U12633 (N_12633,N_11344,N_11273);
nand U12634 (N_12634,N_11025,N_11272);
nor U12635 (N_12635,N_11753,N_11884);
nor U12636 (N_12636,N_11514,N_11003);
nor U12637 (N_12637,N_11192,N_11373);
and U12638 (N_12638,N_11592,N_11123);
and U12639 (N_12639,N_11902,N_11573);
or U12640 (N_12640,N_11980,N_11813);
nand U12641 (N_12641,N_11234,N_11418);
nor U12642 (N_12642,N_11627,N_11160);
nor U12643 (N_12643,N_11090,N_11551);
nor U12644 (N_12644,N_11378,N_11237);
or U12645 (N_12645,N_11447,N_11818);
or U12646 (N_12646,N_11817,N_11016);
or U12647 (N_12647,N_11885,N_11234);
nand U12648 (N_12648,N_11949,N_11572);
nor U12649 (N_12649,N_11695,N_11698);
or U12650 (N_12650,N_11873,N_11752);
and U12651 (N_12651,N_11399,N_11460);
nor U12652 (N_12652,N_11015,N_11118);
nand U12653 (N_12653,N_11476,N_11220);
nor U12654 (N_12654,N_11451,N_11078);
nand U12655 (N_12655,N_11658,N_11308);
or U12656 (N_12656,N_11118,N_11064);
and U12657 (N_12657,N_11432,N_11287);
xnor U12658 (N_12658,N_11629,N_11742);
or U12659 (N_12659,N_11864,N_11804);
or U12660 (N_12660,N_11912,N_11572);
nand U12661 (N_12661,N_11228,N_11362);
or U12662 (N_12662,N_11615,N_11924);
or U12663 (N_12663,N_11383,N_11817);
nand U12664 (N_12664,N_11313,N_11580);
nor U12665 (N_12665,N_11219,N_11422);
nor U12666 (N_12666,N_11418,N_11588);
or U12667 (N_12667,N_11460,N_11729);
or U12668 (N_12668,N_11281,N_11785);
nor U12669 (N_12669,N_11819,N_11529);
nor U12670 (N_12670,N_11127,N_11845);
xnor U12671 (N_12671,N_11978,N_11539);
and U12672 (N_12672,N_11418,N_11677);
nor U12673 (N_12673,N_11678,N_11222);
nor U12674 (N_12674,N_11526,N_11481);
nand U12675 (N_12675,N_11890,N_11837);
nor U12676 (N_12676,N_11875,N_11966);
or U12677 (N_12677,N_11059,N_11558);
or U12678 (N_12678,N_11437,N_11445);
or U12679 (N_12679,N_11679,N_11796);
and U12680 (N_12680,N_11256,N_11079);
nor U12681 (N_12681,N_11852,N_11594);
nand U12682 (N_12682,N_11951,N_11380);
nand U12683 (N_12683,N_11161,N_11654);
nand U12684 (N_12684,N_11490,N_11052);
xnor U12685 (N_12685,N_11158,N_11512);
nand U12686 (N_12686,N_11993,N_11057);
or U12687 (N_12687,N_11234,N_11353);
nor U12688 (N_12688,N_11643,N_11607);
xnor U12689 (N_12689,N_11432,N_11542);
or U12690 (N_12690,N_11348,N_11566);
nor U12691 (N_12691,N_11538,N_11536);
nand U12692 (N_12692,N_11389,N_11301);
nand U12693 (N_12693,N_11532,N_11708);
and U12694 (N_12694,N_11644,N_11136);
nor U12695 (N_12695,N_11040,N_11608);
xnor U12696 (N_12696,N_11312,N_11945);
nor U12697 (N_12697,N_11913,N_11020);
or U12698 (N_12698,N_11701,N_11005);
nor U12699 (N_12699,N_11337,N_11076);
or U12700 (N_12700,N_11380,N_11572);
or U12701 (N_12701,N_11248,N_11240);
or U12702 (N_12702,N_11794,N_11447);
nor U12703 (N_12703,N_11715,N_11346);
and U12704 (N_12704,N_11138,N_11568);
and U12705 (N_12705,N_11274,N_11424);
or U12706 (N_12706,N_11337,N_11049);
nand U12707 (N_12707,N_11583,N_11251);
xnor U12708 (N_12708,N_11452,N_11636);
nand U12709 (N_12709,N_11632,N_11585);
nand U12710 (N_12710,N_11514,N_11584);
xor U12711 (N_12711,N_11801,N_11698);
nand U12712 (N_12712,N_11460,N_11610);
and U12713 (N_12713,N_11039,N_11552);
or U12714 (N_12714,N_11977,N_11609);
or U12715 (N_12715,N_11729,N_11894);
nand U12716 (N_12716,N_11322,N_11913);
or U12717 (N_12717,N_11393,N_11560);
nand U12718 (N_12718,N_11515,N_11925);
or U12719 (N_12719,N_11639,N_11847);
xor U12720 (N_12720,N_11261,N_11074);
xor U12721 (N_12721,N_11367,N_11934);
and U12722 (N_12722,N_11934,N_11264);
or U12723 (N_12723,N_11908,N_11703);
or U12724 (N_12724,N_11717,N_11159);
xor U12725 (N_12725,N_11694,N_11916);
nand U12726 (N_12726,N_11941,N_11554);
or U12727 (N_12727,N_11385,N_11900);
or U12728 (N_12728,N_11104,N_11755);
nor U12729 (N_12729,N_11461,N_11445);
or U12730 (N_12730,N_11565,N_11711);
nor U12731 (N_12731,N_11076,N_11231);
and U12732 (N_12732,N_11447,N_11905);
or U12733 (N_12733,N_11337,N_11193);
and U12734 (N_12734,N_11220,N_11807);
or U12735 (N_12735,N_11803,N_11792);
nor U12736 (N_12736,N_11069,N_11780);
nand U12737 (N_12737,N_11359,N_11638);
nor U12738 (N_12738,N_11428,N_11484);
or U12739 (N_12739,N_11759,N_11992);
nand U12740 (N_12740,N_11872,N_11589);
or U12741 (N_12741,N_11724,N_11730);
nor U12742 (N_12742,N_11490,N_11012);
nor U12743 (N_12743,N_11313,N_11685);
and U12744 (N_12744,N_11312,N_11465);
nor U12745 (N_12745,N_11587,N_11424);
nor U12746 (N_12746,N_11996,N_11076);
nand U12747 (N_12747,N_11489,N_11380);
and U12748 (N_12748,N_11240,N_11695);
nor U12749 (N_12749,N_11260,N_11028);
xor U12750 (N_12750,N_11228,N_11429);
and U12751 (N_12751,N_11010,N_11739);
nor U12752 (N_12752,N_11071,N_11247);
nor U12753 (N_12753,N_11239,N_11360);
and U12754 (N_12754,N_11806,N_11014);
nand U12755 (N_12755,N_11807,N_11161);
and U12756 (N_12756,N_11362,N_11828);
nand U12757 (N_12757,N_11808,N_11032);
xor U12758 (N_12758,N_11039,N_11850);
nand U12759 (N_12759,N_11386,N_11615);
xor U12760 (N_12760,N_11847,N_11291);
and U12761 (N_12761,N_11683,N_11722);
nor U12762 (N_12762,N_11220,N_11919);
or U12763 (N_12763,N_11739,N_11756);
nand U12764 (N_12764,N_11680,N_11946);
and U12765 (N_12765,N_11976,N_11837);
nand U12766 (N_12766,N_11908,N_11773);
xor U12767 (N_12767,N_11383,N_11498);
nand U12768 (N_12768,N_11794,N_11884);
nor U12769 (N_12769,N_11208,N_11119);
and U12770 (N_12770,N_11204,N_11079);
nand U12771 (N_12771,N_11353,N_11500);
and U12772 (N_12772,N_11634,N_11919);
and U12773 (N_12773,N_11841,N_11878);
and U12774 (N_12774,N_11567,N_11415);
nand U12775 (N_12775,N_11529,N_11848);
nand U12776 (N_12776,N_11711,N_11638);
and U12777 (N_12777,N_11807,N_11031);
and U12778 (N_12778,N_11167,N_11890);
xor U12779 (N_12779,N_11689,N_11833);
xnor U12780 (N_12780,N_11663,N_11775);
and U12781 (N_12781,N_11987,N_11768);
nor U12782 (N_12782,N_11335,N_11004);
and U12783 (N_12783,N_11078,N_11805);
and U12784 (N_12784,N_11578,N_11871);
nor U12785 (N_12785,N_11978,N_11111);
or U12786 (N_12786,N_11755,N_11284);
nand U12787 (N_12787,N_11986,N_11389);
or U12788 (N_12788,N_11854,N_11103);
or U12789 (N_12789,N_11231,N_11022);
and U12790 (N_12790,N_11537,N_11898);
nor U12791 (N_12791,N_11469,N_11558);
and U12792 (N_12792,N_11853,N_11154);
or U12793 (N_12793,N_11015,N_11730);
nor U12794 (N_12794,N_11798,N_11902);
nor U12795 (N_12795,N_11160,N_11858);
nand U12796 (N_12796,N_11960,N_11966);
nor U12797 (N_12797,N_11559,N_11102);
or U12798 (N_12798,N_11171,N_11158);
xor U12799 (N_12799,N_11927,N_11065);
nand U12800 (N_12800,N_11222,N_11387);
and U12801 (N_12801,N_11551,N_11639);
or U12802 (N_12802,N_11399,N_11817);
nor U12803 (N_12803,N_11306,N_11791);
nor U12804 (N_12804,N_11220,N_11615);
nand U12805 (N_12805,N_11788,N_11473);
or U12806 (N_12806,N_11865,N_11978);
or U12807 (N_12807,N_11709,N_11490);
nor U12808 (N_12808,N_11413,N_11883);
or U12809 (N_12809,N_11266,N_11420);
and U12810 (N_12810,N_11327,N_11280);
nor U12811 (N_12811,N_11719,N_11384);
or U12812 (N_12812,N_11417,N_11642);
and U12813 (N_12813,N_11881,N_11136);
or U12814 (N_12814,N_11810,N_11319);
and U12815 (N_12815,N_11940,N_11280);
nor U12816 (N_12816,N_11829,N_11272);
nor U12817 (N_12817,N_11619,N_11913);
nand U12818 (N_12818,N_11120,N_11434);
nor U12819 (N_12819,N_11178,N_11462);
nor U12820 (N_12820,N_11882,N_11239);
nand U12821 (N_12821,N_11551,N_11692);
nor U12822 (N_12822,N_11421,N_11024);
nor U12823 (N_12823,N_11752,N_11403);
nand U12824 (N_12824,N_11901,N_11131);
or U12825 (N_12825,N_11215,N_11705);
and U12826 (N_12826,N_11715,N_11112);
or U12827 (N_12827,N_11751,N_11124);
nand U12828 (N_12828,N_11623,N_11456);
or U12829 (N_12829,N_11133,N_11816);
nand U12830 (N_12830,N_11359,N_11539);
xnor U12831 (N_12831,N_11083,N_11203);
nand U12832 (N_12832,N_11121,N_11564);
nor U12833 (N_12833,N_11742,N_11115);
or U12834 (N_12834,N_11248,N_11084);
xnor U12835 (N_12835,N_11774,N_11840);
or U12836 (N_12836,N_11441,N_11959);
nand U12837 (N_12837,N_11762,N_11215);
xnor U12838 (N_12838,N_11762,N_11445);
nor U12839 (N_12839,N_11697,N_11536);
nand U12840 (N_12840,N_11842,N_11457);
nand U12841 (N_12841,N_11196,N_11269);
nand U12842 (N_12842,N_11171,N_11297);
nor U12843 (N_12843,N_11960,N_11924);
and U12844 (N_12844,N_11998,N_11029);
nor U12845 (N_12845,N_11343,N_11926);
xor U12846 (N_12846,N_11663,N_11204);
and U12847 (N_12847,N_11676,N_11960);
and U12848 (N_12848,N_11928,N_11055);
nand U12849 (N_12849,N_11799,N_11599);
xor U12850 (N_12850,N_11742,N_11417);
or U12851 (N_12851,N_11392,N_11210);
xor U12852 (N_12852,N_11409,N_11099);
or U12853 (N_12853,N_11716,N_11528);
or U12854 (N_12854,N_11396,N_11422);
nor U12855 (N_12855,N_11668,N_11439);
nor U12856 (N_12856,N_11698,N_11517);
nand U12857 (N_12857,N_11977,N_11244);
xnor U12858 (N_12858,N_11591,N_11953);
and U12859 (N_12859,N_11736,N_11247);
xor U12860 (N_12860,N_11777,N_11095);
and U12861 (N_12861,N_11381,N_11252);
and U12862 (N_12862,N_11638,N_11194);
or U12863 (N_12863,N_11013,N_11195);
or U12864 (N_12864,N_11545,N_11052);
and U12865 (N_12865,N_11345,N_11959);
and U12866 (N_12866,N_11639,N_11737);
nor U12867 (N_12867,N_11588,N_11391);
or U12868 (N_12868,N_11124,N_11963);
nor U12869 (N_12869,N_11104,N_11058);
or U12870 (N_12870,N_11964,N_11572);
nand U12871 (N_12871,N_11887,N_11396);
or U12872 (N_12872,N_11012,N_11386);
nand U12873 (N_12873,N_11413,N_11882);
nor U12874 (N_12874,N_11000,N_11143);
nand U12875 (N_12875,N_11817,N_11551);
nand U12876 (N_12876,N_11194,N_11446);
and U12877 (N_12877,N_11973,N_11977);
nor U12878 (N_12878,N_11544,N_11500);
or U12879 (N_12879,N_11291,N_11180);
nand U12880 (N_12880,N_11211,N_11557);
and U12881 (N_12881,N_11438,N_11761);
and U12882 (N_12882,N_11530,N_11532);
and U12883 (N_12883,N_11959,N_11638);
nor U12884 (N_12884,N_11818,N_11458);
xor U12885 (N_12885,N_11832,N_11933);
and U12886 (N_12886,N_11631,N_11858);
and U12887 (N_12887,N_11461,N_11379);
and U12888 (N_12888,N_11638,N_11473);
xor U12889 (N_12889,N_11131,N_11955);
nand U12890 (N_12890,N_11358,N_11602);
nand U12891 (N_12891,N_11980,N_11725);
or U12892 (N_12892,N_11290,N_11375);
nand U12893 (N_12893,N_11409,N_11082);
or U12894 (N_12894,N_11310,N_11346);
nor U12895 (N_12895,N_11026,N_11781);
nor U12896 (N_12896,N_11310,N_11755);
nand U12897 (N_12897,N_11663,N_11132);
xnor U12898 (N_12898,N_11863,N_11901);
nand U12899 (N_12899,N_11528,N_11208);
nand U12900 (N_12900,N_11152,N_11953);
or U12901 (N_12901,N_11743,N_11177);
or U12902 (N_12902,N_11936,N_11666);
nand U12903 (N_12903,N_11869,N_11105);
and U12904 (N_12904,N_11432,N_11997);
or U12905 (N_12905,N_11226,N_11959);
nor U12906 (N_12906,N_11980,N_11173);
and U12907 (N_12907,N_11264,N_11282);
nand U12908 (N_12908,N_11492,N_11786);
or U12909 (N_12909,N_11255,N_11537);
and U12910 (N_12910,N_11432,N_11739);
nor U12911 (N_12911,N_11467,N_11964);
or U12912 (N_12912,N_11399,N_11324);
and U12913 (N_12913,N_11632,N_11735);
nand U12914 (N_12914,N_11133,N_11331);
nor U12915 (N_12915,N_11329,N_11941);
nand U12916 (N_12916,N_11664,N_11542);
nand U12917 (N_12917,N_11905,N_11752);
or U12918 (N_12918,N_11450,N_11903);
nor U12919 (N_12919,N_11384,N_11848);
and U12920 (N_12920,N_11503,N_11108);
or U12921 (N_12921,N_11815,N_11505);
xor U12922 (N_12922,N_11740,N_11576);
xor U12923 (N_12923,N_11261,N_11240);
xor U12924 (N_12924,N_11577,N_11163);
xor U12925 (N_12925,N_11346,N_11442);
nor U12926 (N_12926,N_11433,N_11343);
nor U12927 (N_12927,N_11523,N_11318);
nor U12928 (N_12928,N_11323,N_11413);
nor U12929 (N_12929,N_11732,N_11743);
nor U12930 (N_12930,N_11667,N_11405);
xor U12931 (N_12931,N_11252,N_11847);
or U12932 (N_12932,N_11522,N_11720);
nor U12933 (N_12933,N_11233,N_11223);
and U12934 (N_12934,N_11048,N_11865);
nor U12935 (N_12935,N_11802,N_11414);
and U12936 (N_12936,N_11174,N_11000);
and U12937 (N_12937,N_11199,N_11748);
and U12938 (N_12938,N_11179,N_11813);
nand U12939 (N_12939,N_11346,N_11166);
and U12940 (N_12940,N_11825,N_11505);
xor U12941 (N_12941,N_11519,N_11755);
xnor U12942 (N_12942,N_11162,N_11173);
xor U12943 (N_12943,N_11839,N_11850);
nand U12944 (N_12944,N_11496,N_11934);
nor U12945 (N_12945,N_11972,N_11904);
nand U12946 (N_12946,N_11881,N_11230);
and U12947 (N_12947,N_11599,N_11240);
nor U12948 (N_12948,N_11854,N_11670);
and U12949 (N_12949,N_11777,N_11790);
nor U12950 (N_12950,N_11982,N_11730);
or U12951 (N_12951,N_11286,N_11869);
and U12952 (N_12952,N_11612,N_11018);
nor U12953 (N_12953,N_11900,N_11744);
or U12954 (N_12954,N_11830,N_11626);
nor U12955 (N_12955,N_11508,N_11981);
and U12956 (N_12956,N_11250,N_11996);
nor U12957 (N_12957,N_11712,N_11296);
nor U12958 (N_12958,N_11420,N_11408);
or U12959 (N_12959,N_11288,N_11521);
nand U12960 (N_12960,N_11089,N_11194);
nor U12961 (N_12961,N_11635,N_11188);
and U12962 (N_12962,N_11088,N_11196);
nor U12963 (N_12963,N_11833,N_11635);
nor U12964 (N_12964,N_11733,N_11329);
nand U12965 (N_12965,N_11998,N_11269);
nor U12966 (N_12966,N_11201,N_11362);
nor U12967 (N_12967,N_11131,N_11313);
and U12968 (N_12968,N_11029,N_11024);
nand U12969 (N_12969,N_11356,N_11628);
and U12970 (N_12970,N_11897,N_11872);
nand U12971 (N_12971,N_11498,N_11788);
and U12972 (N_12972,N_11196,N_11801);
nand U12973 (N_12973,N_11213,N_11497);
and U12974 (N_12974,N_11008,N_11349);
and U12975 (N_12975,N_11489,N_11008);
xor U12976 (N_12976,N_11329,N_11893);
nand U12977 (N_12977,N_11957,N_11880);
nor U12978 (N_12978,N_11485,N_11965);
xor U12979 (N_12979,N_11567,N_11914);
nor U12980 (N_12980,N_11921,N_11344);
and U12981 (N_12981,N_11357,N_11186);
xor U12982 (N_12982,N_11866,N_11893);
nor U12983 (N_12983,N_11978,N_11582);
nor U12984 (N_12984,N_11250,N_11806);
nand U12985 (N_12985,N_11193,N_11734);
and U12986 (N_12986,N_11626,N_11925);
and U12987 (N_12987,N_11178,N_11509);
and U12988 (N_12988,N_11222,N_11992);
and U12989 (N_12989,N_11619,N_11975);
nand U12990 (N_12990,N_11158,N_11836);
or U12991 (N_12991,N_11683,N_11909);
nor U12992 (N_12992,N_11190,N_11446);
nor U12993 (N_12993,N_11127,N_11484);
nor U12994 (N_12994,N_11399,N_11560);
xnor U12995 (N_12995,N_11430,N_11894);
nor U12996 (N_12996,N_11884,N_11474);
and U12997 (N_12997,N_11998,N_11533);
xnor U12998 (N_12998,N_11564,N_11278);
or U12999 (N_12999,N_11243,N_11730);
and U13000 (N_13000,N_12000,N_12989);
nand U13001 (N_13001,N_12397,N_12217);
or U13002 (N_13002,N_12955,N_12313);
xor U13003 (N_13003,N_12156,N_12751);
and U13004 (N_13004,N_12882,N_12709);
or U13005 (N_13005,N_12515,N_12080);
or U13006 (N_13006,N_12036,N_12169);
or U13007 (N_13007,N_12807,N_12877);
nand U13008 (N_13008,N_12594,N_12719);
nand U13009 (N_13009,N_12839,N_12209);
or U13010 (N_13010,N_12282,N_12998);
xor U13011 (N_13011,N_12335,N_12402);
xnor U13012 (N_13012,N_12237,N_12454);
nand U13013 (N_13013,N_12895,N_12355);
nor U13014 (N_13014,N_12411,N_12403);
nor U13015 (N_13015,N_12983,N_12617);
nor U13016 (N_13016,N_12464,N_12950);
nor U13017 (N_13017,N_12214,N_12239);
xnor U13018 (N_13018,N_12051,N_12671);
nor U13019 (N_13019,N_12984,N_12283);
and U13020 (N_13020,N_12777,N_12910);
or U13021 (N_13021,N_12074,N_12126);
nor U13022 (N_13022,N_12363,N_12542);
nor U13023 (N_13023,N_12143,N_12798);
nand U13024 (N_13024,N_12656,N_12161);
or U13025 (N_13025,N_12177,N_12991);
nor U13026 (N_13026,N_12441,N_12623);
or U13027 (N_13027,N_12692,N_12206);
nand U13028 (N_13028,N_12852,N_12606);
and U13029 (N_13029,N_12163,N_12855);
nor U13030 (N_13030,N_12544,N_12790);
or U13031 (N_13031,N_12199,N_12257);
nor U13032 (N_13032,N_12714,N_12448);
nand U13033 (N_13033,N_12488,N_12672);
nand U13034 (N_13034,N_12121,N_12343);
nand U13035 (N_13035,N_12227,N_12001);
or U13036 (N_13036,N_12965,N_12390);
nand U13037 (N_13037,N_12788,N_12167);
xnor U13038 (N_13038,N_12532,N_12018);
xor U13039 (N_13039,N_12487,N_12136);
xor U13040 (N_13040,N_12967,N_12426);
or U13041 (N_13041,N_12974,N_12219);
nand U13042 (N_13042,N_12259,N_12383);
or U13043 (N_13043,N_12565,N_12326);
and U13044 (N_13044,N_12535,N_12596);
nand U13045 (N_13045,N_12263,N_12255);
nor U13046 (N_13046,N_12701,N_12880);
or U13047 (N_13047,N_12225,N_12869);
and U13048 (N_13048,N_12749,N_12147);
nand U13049 (N_13049,N_12871,N_12662);
nand U13050 (N_13050,N_12508,N_12850);
or U13051 (N_13051,N_12361,N_12805);
and U13052 (N_13052,N_12652,N_12058);
or U13053 (N_13053,N_12049,N_12694);
nand U13054 (N_13054,N_12182,N_12358);
and U13055 (N_13055,N_12425,N_12605);
and U13056 (N_13056,N_12584,N_12858);
nand U13057 (N_13057,N_12502,N_12884);
or U13058 (N_13058,N_12635,N_12015);
nand U13059 (N_13059,N_12248,N_12845);
nor U13060 (N_13060,N_12252,N_12600);
nor U13061 (N_13061,N_12233,N_12624);
nand U13062 (N_13062,N_12764,N_12643);
nor U13063 (N_13063,N_12585,N_12417);
or U13064 (N_13064,N_12949,N_12664);
or U13065 (N_13065,N_12538,N_12774);
and U13066 (N_13066,N_12003,N_12400);
nor U13067 (N_13067,N_12210,N_12075);
nand U13068 (N_13068,N_12513,N_12062);
xor U13069 (N_13069,N_12011,N_12149);
nand U13070 (N_13070,N_12295,N_12829);
and U13071 (N_13071,N_12653,N_12602);
nor U13072 (N_13072,N_12557,N_12471);
nor U13073 (N_13073,N_12646,N_12145);
nor U13074 (N_13074,N_12247,N_12468);
or U13075 (N_13075,N_12301,N_12945);
nand U13076 (N_13076,N_12589,N_12636);
nor U13077 (N_13077,N_12186,N_12887);
nor U13078 (N_13078,N_12530,N_12208);
and U13079 (N_13079,N_12792,N_12994);
nor U13080 (N_13080,N_12378,N_12308);
or U13081 (N_13081,N_12708,N_12319);
and U13082 (N_13082,N_12765,N_12181);
and U13083 (N_13083,N_12657,N_12506);
or U13084 (N_13084,N_12561,N_12309);
nand U13085 (N_13085,N_12689,N_12536);
nand U13086 (N_13086,N_12993,N_12386);
nor U13087 (N_13087,N_12024,N_12851);
and U13088 (N_13088,N_12615,N_12521);
nand U13089 (N_13089,N_12101,N_12682);
nand U13090 (N_13090,N_12197,N_12404);
and U13091 (N_13091,N_12514,N_12742);
nand U13092 (N_13092,N_12549,N_12666);
and U13093 (N_13093,N_12813,N_12273);
or U13094 (N_13094,N_12216,N_12595);
nor U13095 (N_13095,N_12545,N_12835);
and U13096 (N_13096,N_12930,N_12125);
or U13097 (N_13097,N_12614,N_12970);
and U13098 (N_13098,N_12838,N_12418);
nor U13099 (N_13099,N_12756,N_12999);
nor U13100 (N_13100,N_12112,N_12271);
nand U13101 (N_13101,N_12613,N_12477);
and U13102 (N_13102,N_12253,N_12429);
or U13103 (N_13103,N_12031,N_12002);
nor U13104 (N_13104,N_12598,N_12971);
and U13105 (N_13105,N_12892,N_12382);
nor U13106 (N_13106,N_12260,N_12957);
nand U13107 (N_13107,N_12913,N_12444);
nand U13108 (N_13108,N_12463,N_12604);
or U13109 (N_13109,N_12504,N_12392);
nand U13110 (N_13110,N_12572,N_12294);
nand U13111 (N_13111,N_12050,N_12582);
nor U13112 (N_13112,N_12976,N_12338);
xor U13113 (N_13113,N_12281,N_12638);
or U13114 (N_13114,N_12362,N_12391);
or U13115 (N_13115,N_12842,N_12491);
nor U13116 (N_13116,N_12238,N_12028);
nand U13117 (N_13117,N_12787,N_12927);
and U13118 (N_13118,N_12250,N_12038);
nor U13119 (N_13119,N_12469,N_12846);
or U13120 (N_13120,N_12442,N_12479);
and U13121 (N_13121,N_12127,N_12588);
xnor U13122 (N_13122,N_12017,N_12421);
and U13123 (N_13123,N_12619,N_12348);
and U13124 (N_13124,N_12223,N_12325);
nand U13125 (N_13125,N_12684,N_12909);
xnor U13126 (N_13126,N_12783,N_12826);
nand U13127 (N_13127,N_12067,N_12339);
or U13128 (N_13128,N_12629,N_12231);
and U13129 (N_13129,N_12376,N_12496);
nor U13130 (N_13130,N_12800,N_12044);
and U13131 (N_13131,N_12866,N_12990);
or U13132 (N_13132,N_12304,N_12079);
nand U13133 (N_13133,N_12303,N_12172);
or U13134 (N_13134,N_12190,N_12899);
xor U13135 (N_13135,N_12138,N_12276);
nor U13136 (N_13136,N_12921,N_12102);
and U13137 (N_13137,N_12639,N_12280);
nand U13138 (N_13138,N_12366,N_12374);
and U13139 (N_13139,N_12310,N_12739);
nand U13140 (N_13140,N_12196,N_12076);
and U13141 (N_13141,N_12558,N_12559);
and U13142 (N_13142,N_12059,N_12529);
nand U13143 (N_13143,N_12422,N_12706);
or U13144 (N_13144,N_12129,N_12878);
nor U13145 (N_13145,N_12375,N_12753);
or U13146 (N_13146,N_12071,N_12889);
nor U13147 (N_13147,N_12399,N_12410);
nand U13148 (N_13148,N_12528,N_12053);
nand U13149 (N_13149,N_12405,N_12290);
nor U13150 (N_13150,N_12262,N_12377);
or U13151 (N_13151,N_12552,N_12586);
or U13152 (N_13152,N_12801,N_12987);
and U13153 (N_13153,N_12668,N_12415);
and U13154 (N_13154,N_12320,N_12222);
nand U13155 (N_13155,N_12622,N_12816);
nand U13156 (N_13156,N_12936,N_12640);
or U13157 (N_13157,N_12898,N_12941);
xor U13158 (N_13158,N_12266,N_12499);
nand U13159 (N_13159,N_12732,N_12460);
or U13160 (N_13160,N_12010,N_12158);
nor U13161 (N_13161,N_12443,N_12857);
xor U13162 (N_13162,N_12637,N_12691);
nor U13163 (N_13163,N_12110,N_12705);
or U13164 (N_13164,N_12995,N_12799);
nand U13165 (N_13165,N_12052,N_12778);
xor U13166 (N_13166,N_12888,N_12048);
xnor U13167 (N_13167,N_12473,N_12868);
and U13168 (N_13168,N_12583,N_12235);
nand U13169 (N_13169,N_12815,N_12754);
nor U13170 (N_13170,N_12030,N_12795);
and U13171 (N_13171,N_12056,N_12771);
and U13172 (N_13172,N_12961,N_12924);
nand U13173 (N_13173,N_12342,N_12543);
or U13174 (N_13174,N_12287,N_12323);
and U13175 (N_13175,N_12457,N_12911);
nor U13176 (N_13176,N_12328,N_12091);
nor U13177 (N_13177,N_12047,N_12775);
nor U13178 (N_13178,N_12200,N_12953);
nand U13179 (N_13179,N_12943,N_12891);
xor U13180 (N_13180,N_12760,N_12834);
nand U13181 (N_13181,N_12566,N_12776);
nor U13182 (N_13182,N_12687,N_12870);
and U13183 (N_13183,N_12699,N_12420);
nand U13184 (N_13184,N_12440,N_12883);
or U13185 (N_13185,N_12370,N_12019);
or U13186 (N_13186,N_12761,N_12876);
xor U13187 (N_13187,N_12114,N_12201);
and U13188 (N_13188,N_12546,N_12485);
nor U13189 (N_13189,N_12599,N_12204);
and U13190 (N_13190,N_12937,N_12716);
and U13191 (N_13191,N_12633,N_12547);
nand U13192 (N_13192,N_12702,N_12736);
nor U13193 (N_13193,N_12180,N_12537);
nand U13194 (N_13194,N_12917,N_12864);
nand U13195 (N_13195,N_12820,N_12142);
and U13196 (N_13196,N_12134,N_12766);
nand U13197 (N_13197,N_12712,N_12312);
nand U13198 (N_13198,N_12533,N_12269);
or U13199 (N_13199,N_12213,N_12786);
or U13200 (N_13200,N_12069,N_12389);
or U13201 (N_13201,N_12236,N_12318);
or U13202 (N_13202,N_12693,N_12099);
nor U13203 (N_13203,N_12311,N_12095);
and U13204 (N_13204,N_12886,N_12187);
nor U13205 (N_13205,N_12093,N_12686);
and U13206 (N_13206,N_12008,N_12707);
and U13207 (N_13207,N_12428,N_12695);
nand U13208 (N_13208,N_12645,N_12159);
and U13209 (N_13209,N_12492,N_12986);
or U13210 (N_13210,N_12944,N_12240);
and U13211 (N_13211,N_12556,N_12352);
or U13212 (N_13212,N_12357,N_12827);
and U13213 (N_13213,N_12493,N_12450);
nor U13214 (N_13214,N_12195,N_12928);
xnor U13215 (N_13215,N_12916,N_12729);
nor U13216 (N_13216,N_12568,N_12938);
nor U13217 (N_13217,N_12804,N_12828);
nand U13218 (N_13218,N_12218,N_12371);
or U13219 (N_13219,N_12042,N_12388);
xor U13220 (N_13220,N_12670,N_12423);
nor U13221 (N_13221,N_12734,N_12202);
xnor U13222 (N_13222,N_12265,N_12717);
or U13223 (N_13223,N_12992,N_12251);
or U13224 (N_13224,N_12902,N_12368);
nand U13225 (N_13225,N_12270,N_12618);
or U13226 (N_13226,N_12580,N_12427);
nand U13227 (N_13227,N_12856,N_12905);
nand U13228 (N_13228,N_12484,N_12745);
and U13229 (N_13229,N_12948,N_12978);
xor U13230 (N_13230,N_12578,N_12661);
xor U13231 (N_13231,N_12153,N_12437);
nor U13232 (N_13232,N_12144,N_12844);
and U13233 (N_13233,N_12972,N_12497);
nand U13234 (N_13234,N_12296,N_12854);
and U13235 (N_13235,N_12184,N_12152);
nand U13236 (N_13236,N_12579,N_12193);
and U13237 (N_13237,N_12996,N_12780);
and U13238 (N_13238,N_12980,N_12413);
or U13239 (N_13239,N_12609,N_12393);
or U13240 (N_13240,N_12241,N_12525);
nand U13241 (N_13241,N_12475,N_12482);
or U13242 (N_13242,N_12726,N_12211);
nor U13243 (N_13243,N_12013,N_12244);
and U13244 (N_13244,N_12674,N_12433);
nor U13245 (N_13245,N_12680,N_12419);
or U13246 (N_13246,N_12221,N_12735);
or U13247 (N_13247,N_12486,N_12865);
nand U13248 (N_13248,N_12688,N_12249);
or U13249 (N_13249,N_12796,N_12474);
nand U13250 (N_13250,N_12246,N_12398);
and U13251 (N_13251,N_12072,N_12173);
nand U13252 (N_13252,N_12207,N_12894);
and U13253 (N_13253,N_12947,N_12785);
and U13254 (N_13254,N_12185,N_12642);
nor U13255 (N_13255,N_12171,N_12279);
and U13256 (N_13256,N_12907,N_12625);
or U13257 (N_13257,N_12942,N_12020);
nand U13258 (N_13258,N_12331,N_12356);
nand U13259 (N_13259,N_12452,N_12825);
nand U13260 (N_13260,N_12560,N_12278);
or U13261 (N_13261,N_12500,N_12490);
nor U13262 (N_13262,N_12379,N_12113);
xor U13263 (N_13263,N_12272,N_12176);
or U13264 (N_13264,N_12698,N_12453);
nand U13265 (N_13265,N_12567,N_12782);
and U13266 (N_13266,N_12063,N_12228);
nor U13267 (N_13267,N_12848,N_12954);
xnor U13268 (N_13268,N_12317,N_12344);
and U13269 (N_13269,N_12811,N_12498);
xnor U13270 (N_13270,N_12817,N_12396);
nor U13271 (N_13271,N_12025,N_12962);
nor U13272 (N_13272,N_12518,N_12931);
and U13273 (N_13273,N_12016,N_12431);
xnor U13274 (N_13274,N_12781,N_12511);
nand U13275 (N_13275,N_12060,N_12115);
or U13276 (N_13276,N_12853,N_12597);
nand U13277 (N_13277,N_12725,N_12861);
or U13278 (N_13278,N_12654,N_12300);
or U13279 (N_13279,N_12461,N_12307);
nand U13280 (N_13280,N_12906,N_12758);
xor U13281 (N_13281,N_12964,N_12098);
nor U13282 (N_13282,N_12658,N_12456);
nor U13283 (N_13283,N_12576,N_12975);
or U13284 (N_13284,N_12128,N_12258);
or U13285 (N_13285,N_12395,N_12571);
nand U13286 (N_13286,N_12243,N_12165);
or U13287 (N_13287,N_12360,N_12416);
nor U13288 (N_13288,N_12495,N_12085);
nor U13289 (N_13289,N_12007,N_12242);
and U13290 (N_13290,N_12951,N_12291);
and U13291 (N_13291,N_12824,N_12349);
or U13292 (N_13292,N_12918,N_12336);
and U13293 (N_13293,N_12430,N_12626);
nand U13294 (N_13294,N_12968,N_12522);
or U13295 (N_13295,N_12574,N_12340);
and U13296 (N_13296,N_12710,N_12759);
nor U13297 (N_13297,N_12890,N_12478);
xor U13298 (N_13298,N_12772,N_12763);
and U13299 (N_13299,N_12148,N_12057);
nand U13300 (N_13300,N_12517,N_12630);
and U13301 (N_13301,N_12934,N_12078);
nand U13302 (N_13302,N_12510,N_12324);
and U13303 (N_13303,N_12966,N_12401);
nor U13304 (N_13304,N_12347,N_12073);
and U13305 (N_13305,N_12873,N_12840);
nand U13306 (N_13306,N_12026,N_12849);
nand U13307 (N_13307,N_12818,N_12819);
and U13308 (N_13308,N_12933,N_12372);
or U13309 (N_13309,N_12192,N_12963);
or U13310 (N_13310,N_12746,N_12660);
and U13311 (N_13311,N_12224,N_12179);
nand U13312 (N_13312,N_12137,N_12956);
or U13313 (N_13313,N_12641,N_12170);
or U13314 (N_13314,N_12215,N_12897);
nand U13315 (N_13315,N_12037,N_12432);
and U13316 (N_13316,N_12744,N_12140);
nor U13317 (N_13317,N_12908,N_12256);
nor U13318 (N_13318,N_12082,N_12480);
nor U13319 (N_13319,N_12230,N_12676);
and U13320 (N_13320,N_12728,N_12133);
or U13321 (N_13321,N_12120,N_12727);
nor U13322 (N_13322,N_12822,N_12119);
nor U13323 (N_13323,N_12064,N_12472);
xor U13324 (N_13324,N_12503,N_12267);
or U13325 (N_13325,N_12178,N_12068);
and U13326 (N_13326,N_12519,N_12124);
nor U13327 (N_13327,N_12821,N_12268);
nand U13328 (N_13328,N_12040,N_12690);
and U13329 (N_13329,N_12872,N_12900);
nor U13330 (N_13330,N_12066,N_12086);
or U13331 (N_13331,N_12277,N_12446);
xor U13332 (N_13332,N_12168,N_12803);
or U13333 (N_13333,N_12647,N_12407);
nand U13334 (N_13334,N_12935,N_12683);
and U13335 (N_13335,N_12659,N_12084);
nand U13336 (N_13336,N_12679,N_12555);
or U13337 (N_13337,N_12748,N_12563);
nor U13338 (N_13338,N_12284,N_12006);
or U13339 (N_13339,N_12116,N_12959);
nand U13340 (N_13340,N_12982,N_12359);
or U13341 (N_13341,N_12554,N_12592);
nor U13342 (N_13342,N_12550,N_12203);
or U13343 (N_13343,N_12373,N_12979);
or U13344 (N_13344,N_12929,N_12154);
and U13345 (N_13345,N_12548,N_12675);
or U13346 (N_13346,N_12316,N_12245);
and U13347 (N_13347,N_12628,N_12481);
and U13348 (N_13348,N_12539,N_12737);
or U13349 (N_13349,N_12162,N_12151);
and U13350 (N_13350,N_12160,N_12194);
nand U13351 (N_13351,N_12164,N_12476);
nand U13352 (N_13352,N_12061,N_12573);
nand U13353 (N_13353,N_12593,N_12092);
or U13354 (N_13354,N_12946,N_12784);
and U13355 (N_13355,N_12105,N_12004);
nor U13356 (N_13356,N_12608,N_12205);
xor U13357 (N_13357,N_12591,N_12314);
or U13358 (N_13358,N_12723,N_12507);
and U13359 (N_13359,N_12587,N_12673);
nor U13360 (N_13360,N_12509,N_12581);
or U13361 (N_13361,N_12029,N_12449);
nand U13362 (N_13362,N_12512,N_12046);
and U13363 (N_13363,N_12770,N_12409);
and U13364 (N_13364,N_12531,N_12109);
and U13365 (N_13365,N_12229,N_12863);
or U13366 (N_13366,N_12534,N_12226);
and U13367 (N_13367,N_12436,N_12459);
nor U13368 (N_13368,N_12750,N_12081);
nor U13369 (N_13369,N_12329,N_12814);
nand U13370 (N_13370,N_12104,N_12915);
xor U13371 (N_13371,N_12090,N_12603);
nand U13372 (N_13372,N_12132,N_12885);
nand U13373 (N_13373,N_12667,N_12752);
or U13374 (N_13374,N_12035,N_12332);
or U13375 (N_13375,N_12341,N_12733);
or U13376 (N_13376,N_12741,N_12649);
or U13377 (N_13377,N_12131,N_12940);
nand U13378 (N_13378,N_12130,N_12520);
or U13379 (N_13379,N_12769,N_12054);
and U13380 (N_13380,N_12288,N_12925);
nand U13381 (N_13381,N_12569,N_12501);
and U13382 (N_13382,N_12793,N_12923);
or U13383 (N_13383,N_12997,N_12713);
nand U13384 (N_13384,N_12678,N_12087);
nor U13385 (N_13385,N_12973,N_12175);
or U13386 (N_13386,N_12191,N_12874);
or U13387 (N_13387,N_12183,N_12862);
nand U13388 (N_13388,N_12644,N_12009);
nor U13389 (N_13389,N_12135,N_12631);
xnor U13390 (N_13390,N_12330,N_12621);
xnor U13391 (N_13391,N_12097,N_12627);
or U13392 (N_13392,N_12380,N_12650);
xor U13393 (N_13393,N_12447,N_12881);
and U13394 (N_13394,N_12094,N_12364);
and U13395 (N_13395,N_12458,N_12077);
or U13396 (N_13396,N_12146,N_12802);
and U13397 (N_13397,N_12333,N_12394);
and U13398 (N_13398,N_12616,N_12740);
nor U13399 (N_13399,N_12757,N_12577);
and U13400 (N_13400,N_12789,N_12345);
nand U13401 (N_13401,N_12808,N_12860);
or U13402 (N_13402,N_12847,N_12632);
or U13403 (N_13403,N_12843,N_12832);
or U13404 (N_13404,N_12703,N_12470);
and U13405 (N_13405,N_12189,N_12141);
and U13406 (N_13406,N_12369,N_12932);
nand U13407 (N_13407,N_12292,N_12696);
nand U13408 (N_13408,N_12043,N_12424);
nand U13409 (N_13409,N_12711,N_12743);
and U13410 (N_13410,N_12065,N_12367);
nand U13411 (N_13411,N_12767,N_12232);
nor U13412 (N_13412,N_12794,N_12836);
nand U13413 (N_13413,N_12108,N_12837);
xor U13414 (N_13414,N_12715,N_12439);
nor U13415 (N_13415,N_12005,N_12286);
nand U13416 (N_13416,N_12516,N_12648);
and U13417 (N_13417,N_12264,N_12455);
or U13418 (N_13418,N_12334,N_12041);
or U13419 (N_13419,N_12540,N_12365);
and U13420 (N_13420,N_12353,N_12027);
nor U13421 (N_13421,N_12721,N_12575);
nand U13422 (N_13422,N_12022,N_12904);
nor U13423 (N_13423,N_12387,N_12350);
or U13424 (N_13424,N_12039,N_12612);
or U13425 (N_13425,N_12524,N_12275);
or U13426 (N_13426,N_12952,N_12893);
nand U13427 (N_13427,N_12155,N_12139);
nor U13428 (N_13428,N_12466,N_12327);
nand U13429 (N_13429,N_12541,N_12988);
nand U13430 (N_13430,N_12655,N_12985);
nor U13431 (N_13431,N_12111,N_12768);
or U13432 (N_13432,N_12123,N_12920);
and U13433 (N_13433,N_12730,N_12483);
nand U13434 (N_13434,N_12677,N_12914);
and U13435 (N_13435,N_12939,N_12023);
and U13436 (N_13436,N_12435,N_12188);
nand U13437 (N_13437,N_12055,N_12762);
nand U13438 (N_13438,N_12220,N_12083);
and U13439 (N_13439,N_12166,N_12285);
xor U13440 (N_13440,N_12879,N_12299);
nor U13441 (N_13441,N_12412,N_12298);
and U13442 (N_13442,N_12833,N_12354);
nor U13443 (N_13443,N_12489,N_12467);
nor U13444 (N_13444,N_12212,N_12620);
or U13445 (N_13445,N_12021,N_12823);
and U13446 (N_13446,N_12089,N_12700);
xor U13447 (N_13447,N_12032,N_12034);
nor U13448 (N_13448,N_12919,N_12505);
or U13449 (N_13449,N_12922,N_12384);
nor U13450 (N_13450,N_12969,N_12117);
or U13451 (N_13451,N_12903,N_12045);
nor U13452 (N_13452,N_12198,N_12564);
nand U13453 (N_13453,N_12070,N_12088);
or U13454 (N_13454,N_12451,N_12234);
or U13455 (N_13455,N_12526,N_12100);
and U13456 (N_13456,N_12747,N_12118);
and U13457 (N_13457,N_12681,N_12912);
nor U13458 (N_13458,N_12755,N_12590);
nand U13459 (N_13459,N_12321,N_12107);
or U13460 (N_13460,N_12305,N_12859);
xnor U13461 (N_13461,N_12663,N_12523);
nor U13462 (N_13462,N_12791,N_12926);
and U13463 (N_13463,N_12704,N_12337);
and U13464 (N_13464,N_12960,N_12669);
nand U13465 (N_13465,N_12610,N_12809);
xnor U13466 (N_13466,N_12438,N_12841);
nor U13467 (N_13467,N_12607,N_12385);
or U13468 (N_13468,N_12274,N_12651);
nor U13469 (N_13469,N_12958,N_12254);
or U13470 (N_13470,N_12896,N_12465);
nor U13471 (N_13471,N_12611,N_12977);
xnor U13472 (N_13472,N_12665,N_12601);
nand U13473 (N_13473,N_12445,N_12901);
nand U13474 (N_13474,N_12293,N_12812);
nand U13475 (N_13475,N_12875,N_12724);
xnor U13476 (N_13476,N_12014,N_12406);
or U13477 (N_13477,N_12106,N_12562);
or U13478 (N_13478,N_12346,N_12174);
or U13479 (N_13479,N_12351,N_12150);
and U13480 (N_13480,N_12830,N_12462);
nand U13481 (N_13481,N_12779,N_12831);
nand U13482 (N_13482,N_12414,N_12697);
nor U13483 (N_13483,N_12718,N_12434);
xnor U13484 (N_13484,N_12289,N_12722);
or U13485 (N_13485,N_12157,N_12306);
or U13486 (N_13486,N_12553,N_12806);
or U13487 (N_13487,N_12033,N_12867);
nor U13488 (N_13488,N_12096,N_12570);
and U13489 (N_13489,N_12797,N_12720);
nor U13490 (N_13490,N_12810,N_12634);
nor U13491 (N_13491,N_12408,N_12551);
nor U13492 (N_13492,N_12527,N_12494);
nor U13493 (N_13493,N_12981,N_12322);
or U13494 (N_13494,N_12381,N_12685);
or U13495 (N_13495,N_12297,N_12315);
or U13496 (N_13496,N_12738,N_12773);
and U13497 (N_13497,N_12261,N_12122);
nor U13498 (N_13498,N_12731,N_12012);
nor U13499 (N_13499,N_12103,N_12302);
nand U13500 (N_13500,N_12162,N_12218);
nand U13501 (N_13501,N_12310,N_12976);
or U13502 (N_13502,N_12674,N_12717);
xnor U13503 (N_13503,N_12008,N_12000);
or U13504 (N_13504,N_12679,N_12010);
or U13505 (N_13505,N_12528,N_12119);
nand U13506 (N_13506,N_12607,N_12407);
nand U13507 (N_13507,N_12073,N_12445);
nor U13508 (N_13508,N_12279,N_12457);
nand U13509 (N_13509,N_12501,N_12768);
nor U13510 (N_13510,N_12135,N_12740);
and U13511 (N_13511,N_12373,N_12564);
nor U13512 (N_13512,N_12659,N_12916);
nor U13513 (N_13513,N_12424,N_12864);
nor U13514 (N_13514,N_12710,N_12923);
nor U13515 (N_13515,N_12279,N_12807);
nand U13516 (N_13516,N_12250,N_12919);
and U13517 (N_13517,N_12753,N_12960);
nor U13518 (N_13518,N_12931,N_12933);
and U13519 (N_13519,N_12384,N_12660);
xnor U13520 (N_13520,N_12332,N_12765);
and U13521 (N_13521,N_12964,N_12598);
xor U13522 (N_13522,N_12956,N_12508);
nor U13523 (N_13523,N_12517,N_12232);
nor U13524 (N_13524,N_12037,N_12305);
nand U13525 (N_13525,N_12692,N_12140);
nand U13526 (N_13526,N_12315,N_12405);
nor U13527 (N_13527,N_12135,N_12390);
nor U13528 (N_13528,N_12386,N_12012);
nor U13529 (N_13529,N_12591,N_12859);
and U13530 (N_13530,N_12260,N_12027);
or U13531 (N_13531,N_12862,N_12220);
or U13532 (N_13532,N_12359,N_12620);
nor U13533 (N_13533,N_12396,N_12365);
nor U13534 (N_13534,N_12326,N_12468);
and U13535 (N_13535,N_12291,N_12581);
nor U13536 (N_13536,N_12523,N_12393);
nand U13537 (N_13537,N_12673,N_12147);
and U13538 (N_13538,N_12794,N_12719);
and U13539 (N_13539,N_12489,N_12523);
nor U13540 (N_13540,N_12804,N_12358);
xor U13541 (N_13541,N_12993,N_12376);
nor U13542 (N_13542,N_12874,N_12604);
nand U13543 (N_13543,N_12761,N_12854);
nand U13544 (N_13544,N_12962,N_12209);
nor U13545 (N_13545,N_12252,N_12851);
or U13546 (N_13546,N_12651,N_12042);
nor U13547 (N_13547,N_12564,N_12001);
nor U13548 (N_13548,N_12798,N_12813);
xnor U13549 (N_13549,N_12556,N_12101);
nor U13550 (N_13550,N_12497,N_12695);
nor U13551 (N_13551,N_12701,N_12381);
nand U13552 (N_13552,N_12215,N_12074);
and U13553 (N_13553,N_12583,N_12979);
nor U13554 (N_13554,N_12638,N_12654);
or U13555 (N_13555,N_12946,N_12247);
nand U13556 (N_13556,N_12543,N_12365);
and U13557 (N_13557,N_12211,N_12460);
xnor U13558 (N_13558,N_12877,N_12918);
nor U13559 (N_13559,N_12143,N_12076);
nand U13560 (N_13560,N_12323,N_12051);
nor U13561 (N_13561,N_12536,N_12835);
or U13562 (N_13562,N_12890,N_12150);
nor U13563 (N_13563,N_12394,N_12612);
nor U13564 (N_13564,N_12899,N_12282);
or U13565 (N_13565,N_12205,N_12622);
and U13566 (N_13566,N_12364,N_12515);
and U13567 (N_13567,N_12142,N_12339);
or U13568 (N_13568,N_12641,N_12227);
xor U13569 (N_13569,N_12673,N_12438);
or U13570 (N_13570,N_12820,N_12812);
nand U13571 (N_13571,N_12043,N_12462);
nor U13572 (N_13572,N_12172,N_12357);
nand U13573 (N_13573,N_12985,N_12644);
nor U13574 (N_13574,N_12953,N_12062);
or U13575 (N_13575,N_12455,N_12424);
and U13576 (N_13576,N_12986,N_12728);
and U13577 (N_13577,N_12235,N_12066);
nor U13578 (N_13578,N_12000,N_12928);
nor U13579 (N_13579,N_12443,N_12185);
nand U13580 (N_13580,N_12636,N_12312);
or U13581 (N_13581,N_12556,N_12900);
or U13582 (N_13582,N_12031,N_12799);
and U13583 (N_13583,N_12525,N_12958);
xnor U13584 (N_13584,N_12412,N_12305);
xnor U13585 (N_13585,N_12058,N_12659);
and U13586 (N_13586,N_12579,N_12268);
nor U13587 (N_13587,N_12230,N_12177);
nand U13588 (N_13588,N_12192,N_12602);
nand U13589 (N_13589,N_12049,N_12278);
nand U13590 (N_13590,N_12831,N_12165);
or U13591 (N_13591,N_12150,N_12571);
nor U13592 (N_13592,N_12375,N_12334);
or U13593 (N_13593,N_12580,N_12141);
nor U13594 (N_13594,N_12863,N_12692);
and U13595 (N_13595,N_12710,N_12645);
nand U13596 (N_13596,N_12586,N_12423);
nand U13597 (N_13597,N_12976,N_12809);
nand U13598 (N_13598,N_12927,N_12287);
nor U13599 (N_13599,N_12914,N_12882);
nor U13600 (N_13600,N_12187,N_12671);
and U13601 (N_13601,N_12241,N_12253);
nor U13602 (N_13602,N_12663,N_12213);
xnor U13603 (N_13603,N_12003,N_12683);
and U13604 (N_13604,N_12600,N_12400);
and U13605 (N_13605,N_12159,N_12334);
nand U13606 (N_13606,N_12978,N_12310);
nand U13607 (N_13607,N_12968,N_12564);
or U13608 (N_13608,N_12668,N_12259);
nand U13609 (N_13609,N_12534,N_12073);
or U13610 (N_13610,N_12967,N_12358);
or U13611 (N_13611,N_12866,N_12989);
and U13612 (N_13612,N_12310,N_12426);
and U13613 (N_13613,N_12688,N_12947);
nor U13614 (N_13614,N_12657,N_12109);
xnor U13615 (N_13615,N_12184,N_12499);
xor U13616 (N_13616,N_12272,N_12044);
and U13617 (N_13617,N_12402,N_12088);
or U13618 (N_13618,N_12999,N_12992);
and U13619 (N_13619,N_12852,N_12829);
nand U13620 (N_13620,N_12526,N_12493);
nor U13621 (N_13621,N_12618,N_12296);
or U13622 (N_13622,N_12262,N_12555);
nor U13623 (N_13623,N_12564,N_12652);
or U13624 (N_13624,N_12537,N_12349);
or U13625 (N_13625,N_12244,N_12052);
nand U13626 (N_13626,N_12772,N_12624);
and U13627 (N_13627,N_12159,N_12065);
nand U13628 (N_13628,N_12704,N_12147);
nor U13629 (N_13629,N_12368,N_12522);
xor U13630 (N_13630,N_12710,N_12605);
and U13631 (N_13631,N_12894,N_12925);
nand U13632 (N_13632,N_12558,N_12376);
nor U13633 (N_13633,N_12339,N_12448);
or U13634 (N_13634,N_12571,N_12721);
and U13635 (N_13635,N_12926,N_12434);
or U13636 (N_13636,N_12618,N_12393);
nor U13637 (N_13637,N_12748,N_12098);
or U13638 (N_13638,N_12901,N_12350);
or U13639 (N_13639,N_12826,N_12745);
or U13640 (N_13640,N_12630,N_12455);
nand U13641 (N_13641,N_12608,N_12373);
and U13642 (N_13642,N_12016,N_12951);
nand U13643 (N_13643,N_12047,N_12951);
nor U13644 (N_13644,N_12763,N_12452);
nor U13645 (N_13645,N_12554,N_12327);
nor U13646 (N_13646,N_12802,N_12064);
or U13647 (N_13647,N_12816,N_12499);
and U13648 (N_13648,N_12532,N_12035);
and U13649 (N_13649,N_12275,N_12990);
nand U13650 (N_13650,N_12540,N_12938);
or U13651 (N_13651,N_12839,N_12246);
and U13652 (N_13652,N_12763,N_12001);
nand U13653 (N_13653,N_12145,N_12514);
nand U13654 (N_13654,N_12781,N_12069);
nand U13655 (N_13655,N_12426,N_12610);
nand U13656 (N_13656,N_12608,N_12708);
and U13657 (N_13657,N_12248,N_12934);
nand U13658 (N_13658,N_12781,N_12627);
or U13659 (N_13659,N_12906,N_12428);
nor U13660 (N_13660,N_12407,N_12656);
nor U13661 (N_13661,N_12300,N_12663);
or U13662 (N_13662,N_12420,N_12150);
and U13663 (N_13663,N_12686,N_12759);
xor U13664 (N_13664,N_12142,N_12029);
or U13665 (N_13665,N_12736,N_12590);
nand U13666 (N_13666,N_12706,N_12229);
nor U13667 (N_13667,N_12247,N_12764);
xnor U13668 (N_13668,N_12295,N_12924);
and U13669 (N_13669,N_12633,N_12148);
or U13670 (N_13670,N_12033,N_12318);
or U13671 (N_13671,N_12655,N_12122);
and U13672 (N_13672,N_12036,N_12502);
nand U13673 (N_13673,N_12266,N_12694);
nor U13674 (N_13674,N_12170,N_12242);
nor U13675 (N_13675,N_12899,N_12238);
nor U13676 (N_13676,N_12295,N_12596);
nor U13677 (N_13677,N_12190,N_12576);
or U13678 (N_13678,N_12772,N_12766);
xnor U13679 (N_13679,N_12071,N_12165);
or U13680 (N_13680,N_12112,N_12932);
nand U13681 (N_13681,N_12212,N_12708);
nand U13682 (N_13682,N_12231,N_12538);
or U13683 (N_13683,N_12905,N_12560);
nand U13684 (N_13684,N_12083,N_12792);
or U13685 (N_13685,N_12958,N_12161);
nand U13686 (N_13686,N_12798,N_12384);
and U13687 (N_13687,N_12439,N_12474);
or U13688 (N_13688,N_12022,N_12765);
and U13689 (N_13689,N_12383,N_12649);
nor U13690 (N_13690,N_12687,N_12151);
nor U13691 (N_13691,N_12316,N_12498);
and U13692 (N_13692,N_12388,N_12928);
nor U13693 (N_13693,N_12700,N_12079);
nor U13694 (N_13694,N_12115,N_12304);
and U13695 (N_13695,N_12039,N_12342);
nand U13696 (N_13696,N_12387,N_12216);
nor U13697 (N_13697,N_12266,N_12766);
xnor U13698 (N_13698,N_12720,N_12873);
nand U13699 (N_13699,N_12338,N_12510);
nor U13700 (N_13700,N_12769,N_12561);
and U13701 (N_13701,N_12837,N_12978);
and U13702 (N_13702,N_12888,N_12508);
nor U13703 (N_13703,N_12019,N_12710);
nand U13704 (N_13704,N_12146,N_12955);
nand U13705 (N_13705,N_12035,N_12014);
nor U13706 (N_13706,N_12708,N_12481);
xnor U13707 (N_13707,N_12561,N_12393);
or U13708 (N_13708,N_12068,N_12421);
or U13709 (N_13709,N_12004,N_12824);
nor U13710 (N_13710,N_12443,N_12384);
nand U13711 (N_13711,N_12500,N_12019);
and U13712 (N_13712,N_12431,N_12894);
or U13713 (N_13713,N_12370,N_12955);
nor U13714 (N_13714,N_12416,N_12233);
and U13715 (N_13715,N_12302,N_12446);
nor U13716 (N_13716,N_12469,N_12920);
and U13717 (N_13717,N_12345,N_12104);
or U13718 (N_13718,N_12515,N_12712);
nand U13719 (N_13719,N_12565,N_12186);
nand U13720 (N_13720,N_12992,N_12412);
xor U13721 (N_13721,N_12322,N_12369);
nand U13722 (N_13722,N_12525,N_12704);
nor U13723 (N_13723,N_12299,N_12514);
or U13724 (N_13724,N_12839,N_12069);
xnor U13725 (N_13725,N_12244,N_12484);
and U13726 (N_13726,N_12229,N_12286);
and U13727 (N_13727,N_12863,N_12116);
xor U13728 (N_13728,N_12820,N_12681);
xor U13729 (N_13729,N_12467,N_12218);
nand U13730 (N_13730,N_12518,N_12832);
xnor U13731 (N_13731,N_12180,N_12063);
xor U13732 (N_13732,N_12167,N_12459);
or U13733 (N_13733,N_12509,N_12056);
or U13734 (N_13734,N_12220,N_12830);
nand U13735 (N_13735,N_12309,N_12945);
and U13736 (N_13736,N_12460,N_12797);
xnor U13737 (N_13737,N_12977,N_12503);
or U13738 (N_13738,N_12805,N_12122);
nand U13739 (N_13739,N_12136,N_12879);
or U13740 (N_13740,N_12665,N_12998);
nand U13741 (N_13741,N_12826,N_12055);
or U13742 (N_13742,N_12781,N_12366);
xor U13743 (N_13743,N_12257,N_12852);
nand U13744 (N_13744,N_12387,N_12043);
nor U13745 (N_13745,N_12128,N_12293);
xor U13746 (N_13746,N_12493,N_12784);
nand U13747 (N_13747,N_12270,N_12263);
nand U13748 (N_13748,N_12817,N_12866);
nor U13749 (N_13749,N_12263,N_12215);
and U13750 (N_13750,N_12336,N_12293);
and U13751 (N_13751,N_12764,N_12557);
nor U13752 (N_13752,N_12048,N_12864);
nor U13753 (N_13753,N_12410,N_12969);
or U13754 (N_13754,N_12023,N_12696);
nand U13755 (N_13755,N_12071,N_12934);
or U13756 (N_13756,N_12236,N_12260);
or U13757 (N_13757,N_12196,N_12849);
nand U13758 (N_13758,N_12479,N_12436);
or U13759 (N_13759,N_12502,N_12648);
and U13760 (N_13760,N_12127,N_12619);
or U13761 (N_13761,N_12730,N_12658);
and U13762 (N_13762,N_12563,N_12424);
nand U13763 (N_13763,N_12055,N_12658);
nor U13764 (N_13764,N_12235,N_12323);
nand U13765 (N_13765,N_12583,N_12856);
xor U13766 (N_13766,N_12163,N_12739);
nor U13767 (N_13767,N_12438,N_12601);
nor U13768 (N_13768,N_12359,N_12703);
or U13769 (N_13769,N_12293,N_12821);
and U13770 (N_13770,N_12459,N_12189);
nand U13771 (N_13771,N_12591,N_12256);
nand U13772 (N_13772,N_12759,N_12693);
nand U13773 (N_13773,N_12502,N_12604);
nand U13774 (N_13774,N_12589,N_12808);
nor U13775 (N_13775,N_12707,N_12954);
nand U13776 (N_13776,N_12692,N_12802);
nand U13777 (N_13777,N_12329,N_12785);
nand U13778 (N_13778,N_12317,N_12840);
and U13779 (N_13779,N_12831,N_12606);
nor U13780 (N_13780,N_12321,N_12030);
nor U13781 (N_13781,N_12994,N_12389);
nor U13782 (N_13782,N_12237,N_12519);
xnor U13783 (N_13783,N_12966,N_12315);
and U13784 (N_13784,N_12976,N_12111);
nor U13785 (N_13785,N_12911,N_12391);
nor U13786 (N_13786,N_12243,N_12338);
and U13787 (N_13787,N_12175,N_12232);
and U13788 (N_13788,N_12649,N_12160);
and U13789 (N_13789,N_12201,N_12691);
xnor U13790 (N_13790,N_12371,N_12392);
nand U13791 (N_13791,N_12109,N_12364);
nand U13792 (N_13792,N_12363,N_12865);
nor U13793 (N_13793,N_12065,N_12590);
and U13794 (N_13794,N_12091,N_12019);
nor U13795 (N_13795,N_12329,N_12382);
or U13796 (N_13796,N_12698,N_12077);
nand U13797 (N_13797,N_12481,N_12154);
nor U13798 (N_13798,N_12667,N_12262);
nand U13799 (N_13799,N_12872,N_12144);
xnor U13800 (N_13800,N_12828,N_12131);
and U13801 (N_13801,N_12883,N_12540);
xor U13802 (N_13802,N_12411,N_12732);
or U13803 (N_13803,N_12955,N_12321);
or U13804 (N_13804,N_12058,N_12823);
nor U13805 (N_13805,N_12566,N_12267);
and U13806 (N_13806,N_12960,N_12394);
nand U13807 (N_13807,N_12245,N_12962);
nor U13808 (N_13808,N_12228,N_12619);
nor U13809 (N_13809,N_12235,N_12060);
nand U13810 (N_13810,N_12053,N_12509);
xor U13811 (N_13811,N_12278,N_12299);
or U13812 (N_13812,N_12664,N_12396);
or U13813 (N_13813,N_12911,N_12055);
nor U13814 (N_13814,N_12633,N_12191);
nand U13815 (N_13815,N_12335,N_12264);
and U13816 (N_13816,N_12412,N_12165);
or U13817 (N_13817,N_12957,N_12116);
nor U13818 (N_13818,N_12128,N_12965);
nor U13819 (N_13819,N_12246,N_12734);
nand U13820 (N_13820,N_12047,N_12364);
nand U13821 (N_13821,N_12279,N_12025);
nand U13822 (N_13822,N_12585,N_12430);
xnor U13823 (N_13823,N_12481,N_12864);
nor U13824 (N_13824,N_12732,N_12303);
or U13825 (N_13825,N_12309,N_12512);
and U13826 (N_13826,N_12959,N_12530);
and U13827 (N_13827,N_12078,N_12481);
and U13828 (N_13828,N_12384,N_12755);
and U13829 (N_13829,N_12062,N_12571);
or U13830 (N_13830,N_12356,N_12431);
nor U13831 (N_13831,N_12770,N_12081);
nor U13832 (N_13832,N_12464,N_12106);
nor U13833 (N_13833,N_12046,N_12343);
or U13834 (N_13834,N_12441,N_12615);
and U13835 (N_13835,N_12142,N_12683);
and U13836 (N_13836,N_12935,N_12603);
and U13837 (N_13837,N_12464,N_12628);
and U13838 (N_13838,N_12031,N_12124);
nand U13839 (N_13839,N_12432,N_12213);
and U13840 (N_13840,N_12405,N_12288);
xor U13841 (N_13841,N_12817,N_12111);
and U13842 (N_13842,N_12906,N_12488);
and U13843 (N_13843,N_12599,N_12865);
and U13844 (N_13844,N_12234,N_12696);
or U13845 (N_13845,N_12955,N_12135);
and U13846 (N_13846,N_12179,N_12080);
and U13847 (N_13847,N_12056,N_12472);
xor U13848 (N_13848,N_12922,N_12553);
nor U13849 (N_13849,N_12370,N_12870);
nor U13850 (N_13850,N_12958,N_12231);
or U13851 (N_13851,N_12498,N_12834);
or U13852 (N_13852,N_12452,N_12801);
and U13853 (N_13853,N_12654,N_12914);
nor U13854 (N_13854,N_12200,N_12438);
nand U13855 (N_13855,N_12822,N_12379);
nand U13856 (N_13856,N_12609,N_12936);
nor U13857 (N_13857,N_12772,N_12571);
nand U13858 (N_13858,N_12465,N_12079);
nor U13859 (N_13859,N_12222,N_12933);
nor U13860 (N_13860,N_12478,N_12422);
and U13861 (N_13861,N_12923,N_12412);
nand U13862 (N_13862,N_12645,N_12079);
xor U13863 (N_13863,N_12144,N_12828);
and U13864 (N_13864,N_12023,N_12649);
and U13865 (N_13865,N_12616,N_12609);
xnor U13866 (N_13866,N_12903,N_12467);
nor U13867 (N_13867,N_12003,N_12985);
xnor U13868 (N_13868,N_12709,N_12120);
nand U13869 (N_13869,N_12998,N_12430);
or U13870 (N_13870,N_12829,N_12859);
and U13871 (N_13871,N_12184,N_12379);
xor U13872 (N_13872,N_12862,N_12096);
or U13873 (N_13873,N_12409,N_12721);
nand U13874 (N_13874,N_12170,N_12110);
and U13875 (N_13875,N_12154,N_12875);
or U13876 (N_13876,N_12163,N_12790);
nand U13877 (N_13877,N_12400,N_12042);
nor U13878 (N_13878,N_12856,N_12647);
or U13879 (N_13879,N_12866,N_12638);
nor U13880 (N_13880,N_12667,N_12906);
nor U13881 (N_13881,N_12520,N_12683);
nor U13882 (N_13882,N_12207,N_12063);
or U13883 (N_13883,N_12270,N_12703);
nand U13884 (N_13884,N_12816,N_12007);
or U13885 (N_13885,N_12216,N_12541);
nand U13886 (N_13886,N_12749,N_12809);
nor U13887 (N_13887,N_12551,N_12851);
or U13888 (N_13888,N_12094,N_12526);
xor U13889 (N_13889,N_12655,N_12412);
nand U13890 (N_13890,N_12867,N_12627);
or U13891 (N_13891,N_12234,N_12829);
nand U13892 (N_13892,N_12478,N_12988);
nor U13893 (N_13893,N_12108,N_12761);
xor U13894 (N_13894,N_12544,N_12607);
or U13895 (N_13895,N_12372,N_12424);
nand U13896 (N_13896,N_12076,N_12384);
and U13897 (N_13897,N_12812,N_12044);
xor U13898 (N_13898,N_12937,N_12361);
nand U13899 (N_13899,N_12842,N_12879);
or U13900 (N_13900,N_12800,N_12940);
nand U13901 (N_13901,N_12932,N_12491);
nor U13902 (N_13902,N_12771,N_12382);
nor U13903 (N_13903,N_12591,N_12991);
nor U13904 (N_13904,N_12031,N_12974);
nand U13905 (N_13905,N_12691,N_12781);
or U13906 (N_13906,N_12533,N_12298);
and U13907 (N_13907,N_12973,N_12516);
and U13908 (N_13908,N_12209,N_12359);
or U13909 (N_13909,N_12405,N_12843);
nor U13910 (N_13910,N_12492,N_12647);
or U13911 (N_13911,N_12116,N_12835);
and U13912 (N_13912,N_12410,N_12434);
or U13913 (N_13913,N_12083,N_12897);
nand U13914 (N_13914,N_12469,N_12563);
and U13915 (N_13915,N_12891,N_12287);
nor U13916 (N_13916,N_12773,N_12502);
nor U13917 (N_13917,N_12957,N_12492);
or U13918 (N_13918,N_12102,N_12271);
nand U13919 (N_13919,N_12692,N_12828);
nand U13920 (N_13920,N_12525,N_12050);
nor U13921 (N_13921,N_12243,N_12709);
nor U13922 (N_13922,N_12817,N_12347);
nand U13923 (N_13923,N_12446,N_12627);
nand U13924 (N_13924,N_12484,N_12606);
nor U13925 (N_13925,N_12980,N_12788);
xor U13926 (N_13926,N_12154,N_12801);
nand U13927 (N_13927,N_12549,N_12326);
xor U13928 (N_13928,N_12238,N_12451);
and U13929 (N_13929,N_12773,N_12386);
xnor U13930 (N_13930,N_12744,N_12310);
and U13931 (N_13931,N_12318,N_12602);
nor U13932 (N_13932,N_12940,N_12726);
and U13933 (N_13933,N_12948,N_12788);
nand U13934 (N_13934,N_12727,N_12016);
nand U13935 (N_13935,N_12277,N_12223);
or U13936 (N_13936,N_12847,N_12174);
nor U13937 (N_13937,N_12232,N_12011);
and U13938 (N_13938,N_12896,N_12933);
or U13939 (N_13939,N_12096,N_12362);
nor U13940 (N_13940,N_12937,N_12951);
and U13941 (N_13941,N_12334,N_12510);
nand U13942 (N_13942,N_12483,N_12957);
nor U13943 (N_13943,N_12031,N_12132);
nand U13944 (N_13944,N_12971,N_12917);
nand U13945 (N_13945,N_12910,N_12619);
xnor U13946 (N_13946,N_12706,N_12892);
nor U13947 (N_13947,N_12553,N_12274);
xor U13948 (N_13948,N_12145,N_12251);
and U13949 (N_13949,N_12697,N_12735);
nor U13950 (N_13950,N_12062,N_12231);
xor U13951 (N_13951,N_12347,N_12082);
or U13952 (N_13952,N_12310,N_12846);
nand U13953 (N_13953,N_12625,N_12066);
nand U13954 (N_13954,N_12071,N_12078);
or U13955 (N_13955,N_12876,N_12012);
and U13956 (N_13956,N_12933,N_12599);
nor U13957 (N_13957,N_12802,N_12797);
or U13958 (N_13958,N_12697,N_12674);
and U13959 (N_13959,N_12476,N_12210);
and U13960 (N_13960,N_12466,N_12221);
or U13961 (N_13961,N_12372,N_12588);
and U13962 (N_13962,N_12658,N_12770);
and U13963 (N_13963,N_12588,N_12882);
and U13964 (N_13964,N_12559,N_12063);
nor U13965 (N_13965,N_12368,N_12878);
nor U13966 (N_13966,N_12953,N_12517);
xnor U13967 (N_13967,N_12524,N_12190);
nand U13968 (N_13968,N_12656,N_12716);
or U13969 (N_13969,N_12953,N_12268);
and U13970 (N_13970,N_12415,N_12074);
or U13971 (N_13971,N_12650,N_12788);
or U13972 (N_13972,N_12580,N_12668);
nand U13973 (N_13973,N_12414,N_12261);
nor U13974 (N_13974,N_12184,N_12491);
xor U13975 (N_13975,N_12941,N_12101);
and U13976 (N_13976,N_12209,N_12397);
nor U13977 (N_13977,N_12959,N_12750);
or U13978 (N_13978,N_12485,N_12066);
or U13979 (N_13979,N_12110,N_12824);
nor U13980 (N_13980,N_12768,N_12179);
nor U13981 (N_13981,N_12611,N_12087);
xor U13982 (N_13982,N_12035,N_12963);
and U13983 (N_13983,N_12547,N_12361);
nand U13984 (N_13984,N_12629,N_12280);
xor U13985 (N_13985,N_12173,N_12890);
or U13986 (N_13986,N_12055,N_12604);
nand U13987 (N_13987,N_12583,N_12199);
or U13988 (N_13988,N_12491,N_12274);
or U13989 (N_13989,N_12423,N_12972);
and U13990 (N_13990,N_12811,N_12299);
nor U13991 (N_13991,N_12928,N_12507);
nor U13992 (N_13992,N_12543,N_12396);
and U13993 (N_13993,N_12845,N_12665);
or U13994 (N_13994,N_12114,N_12069);
and U13995 (N_13995,N_12650,N_12576);
nor U13996 (N_13996,N_12572,N_12594);
xnor U13997 (N_13997,N_12523,N_12829);
nor U13998 (N_13998,N_12102,N_12928);
nor U13999 (N_13999,N_12584,N_12448);
nand U14000 (N_14000,N_13488,N_13098);
nand U14001 (N_14001,N_13354,N_13036);
and U14002 (N_14002,N_13486,N_13523);
nand U14003 (N_14003,N_13765,N_13821);
and U14004 (N_14004,N_13651,N_13965);
and U14005 (N_14005,N_13095,N_13740);
nor U14006 (N_14006,N_13876,N_13730);
nor U14007 (N_14007,N_13463,N_13238);
and U14008 (N_14008,N_13737,N_13469);
and U14009 (N_14009,N_13418,N_13173);
nor U14010 (N_14010,N_13636,N_13849);
nand U14011 (N_14011,N_13243,N_13580);
nor U14012 (N_14012,N_13624,N_13249);
xor U14013 (N_14013,N_13426,N_13809);
or U14014 (N_14014,N_13402,N_13177);
xnor U14015 (N_14015,N_13917,N_13033);
nand U14016 (N_14016,N_13604,N_13495);
and U14017 (N_14017,N_13029,N_13622);
nor U14018 (N_14018,N_13091,N_13387);
or U14019 (N_14019,N_13712,N_13031);
or U14020 (N_14020,N_13168,N_13052);
nor U14021 (N_14021,N_13422,N_13760);
xnor U14022 (N_14022,N_13151,N_13562);
xnor U14023 (N_14023,N_13334,N_13817);
nor U14024 (N_14024,N_13159,N_13648);
or U14025 (N_14025,N_13076,N_13181);
and U14026 (N_14026,N_13815,N_13374);
nand U14027 (N_14027,N_13125,N_13278);
nor U14028 (N_14028,N_13135,N_13072);
or U14029 (N_14029,N_13451,N_13943);
nor U14030 (N_14030,N_13048,N_13642);
and U14031 (N_14031,N_13211,N_13128);
nor U14032 (N_14032,N_13365,N_13573);
or U14033 (N_14033,N_13319,N_13529);
nor U14034 (N_14034,N_13873,N_13621);
and U14035 (N_14035,N_13681,N_13153);
nor U14036 (N_14036,N_13443,N_13901);
or U14037 (N_14037,N_13596,N_13263);
nand U14038 (N_14038,N_13942,N_13617);
or U14039 (N_14039,N_13685,N_13498);
nor U14040 (N_14040,N_13741,N_13096);
nand U14041 (N_14041,N_13259,N_13574);
nor U14042 (N_14042,N_13919,N_13613);
or U14043 (N_14043,N_13522,N_13215);
nand U14044 (N_14044,N_13021,N_13951);
or U14045 (N_14045,N_13851,N_13814);
and U14046 (N_14046,N_13258,N_13708);
and U14047 (N_14047,N_13588,N_13466);
and U14048 (N_14048,N_13534,N_13736);
or U14049 (N_14049,N_13755,N_13081);
and U14050 (N_14050,N_13936,N_13510);
nand U14051 (N_14051,N_13302,N_13930);
xor U14052 (N_14052,N_13692,N_13360);
and U14053 (N_14053,N_13179,N_13246);
and U14054 (N_14054,N_13967,N_13801);
or U14055 (N_14055,N_13117,N_13050);
nor U14056 (N_14056,N_13137,N_13156);
xor U14057 (N_14057,N_13183,N_13370);
and U14058 (N_14058,N_13652,N_13390);
or U14059 (N_14059,N_13524,N_13442);
or U14060 (N_14060,N_13157,N_13892);
and U14061 (N_14061,N_13269,N_13414);
nor U14062 (N_14062,N_13499,N_13615);
and U14063 (N_14063,N_13541,N_13823);
nor U14064 (N_14064,N_13417,N_13966);
and U14065 (N_14065,N_13436,N_13010);
or U14066 (N_14066,N_13092,N_13280);
nand U14067 (N_14067,N_13663,N_13424);
nand U14068 (N_14068,N_13839,N_13282);
and U14069 (N_14069,N_13535,N_13607);
nand U14070 (N_14070,N_13716,N_13078);
and U14071 (N_14071,N_13608,N_13399);
or U14072 (N_14072,N_13080,N_13467);
nand U14073 (N_14073,N_13266,N_13083);
or U14074 (N_14074,N_13700,N_13361);
or U14075 (N_14075,N_13165,N_13518);
nor U14076 (N_14076,N_13514,N_13383);
and U14077 (N_14077,N_13353,N_13471);
and U14078 (N_14078,N_13500,N_13074);
and U14079 (N_14079,N_13493,N_13688);
nor U14080 (N_14080,N_13233,N_13234);
and U14081 (N_14081,N_13998,N_13643);
and U14082 (N_14082,N_13844,N_13953);
or U14083 (N_14083,N_13237,N_13551);
or U14084 (N_14084,N_13475,N_13497);
nand U14085 (N_14085,N_13980,N_13971);
or U14086 (N_14086,N_13411,N_13767);
and U14087 (N_14087,N_13579,N_13589);
and U14088 (N_14088,N_13987,N_13232);
and U14089 (N_14089,N_13837,N_13556);
nor U14090 (N_14090,N_13576,N_13264);
and U14091 (N_14091,N_13056,N_13062);
nand U14092 (N_14092,N_13047,N_13388);
nor U14093 (N_14093,N_13777,N_13260);
nand U14094 (N_14094,N_13400,N_13057);
and U14095 (N_14095,N_13061,N_13447);
and U14096 (N_14096,N_13526,N_13199);
nand U14097 (N_14097,N_13216,N_13188);
nor U14098 (N_14098,N_13315,N_13275);
nand U14099 (N_14099,N_13537,N_13582);
and U14100 (N_14100,N_13875,N_13401);
nor U14101 (N_14101,N_13931,N_13207);
nand U14102 (N_14102,N_13060,N_13727);
and U14103 (N_14103,N_13271,N_13673);
nor U14104 (N_14104,N_13833,N_13569);
and U14105 (N_14105,N_13182,N_13605);
nand U14106 (N_14106,N_13515,N_13889);
nand U14107 (N_14107,N_13940,N_13894);
or U14108 (N_14108,N_13783,N_13077);
and U14109 (N_14109,N_13542,N_13472);
nand U14110 (N_14110,N_13773,N_13295);
and U14111 (N_14111,N_13881,N_13070);
nor U14112 (N_14112,N_13300,N_13960);
nor U14113 (N_14113,N_13085,N_13464);
or U14114 (N_14114,N_13208,N_13650);
nand U14115 (N_14115,N_13598,N_13709);
nand U14116 (N_14116,N_13570,N_13540);
or U14117 (N_14117,N_13364,N_13553);
nand U14118 (N_14118,N_13481,N_13721);
xnor U14119 (N_14119,N_13593,N_13735);
and U14120 (N_14120,N_13776,N_13880);
and U14121 (N_14121,N_13140,N_13016);
and U14122 (N_14122,N_13385,N_13254);
or U14123 (N_14123,N_13143,N_13867);
nor U14124 (N_14124,N_13004,N_13274);
nor U14125 (N_14125,N_13158,N_13829);
nand U14126 (N_14126,N_13206,N_13185);
and U14127 (N_14127,N_13398,N_13819);
nand U14128 (N_14128,N_13090,N_13338);
nor U14129 (N_14129,N_13386,N_13419);
xor U14130 (N_14130,N_13119,N_13903);
nor U14131 (N_14131,N_13792,N_13668);
nor U14132 (N_14132,N_13494,N_13743);
and U14133 (N_14133,N_13732,N_13267);
and U14134 (N_14134,N_13192,N_13214);
xor U14135 (N_14135,N_13797,N_13381);
or U14136 (N_14136,N_13150,N_13152);
and U14137 (N_14137,N_13926,N_13883);
nor U14138 (N_14138,N_13321,N_13130);
nand U14139 (N_14139,N_13439,N_13154);
nor U14140 (N_14140,N_13195,N_13590);
or U14141 (N_14141,N_13440,N_13291);
nor U14142 (N_14142,N_13898,N_13812);
nand U14143 (N_14143,N_13788,N_13799);
and U14144 (N_14144,N_13123,N_13629);
and U14145 (N_14145,N_13226,N_13209);
nand U14146 (N_14146,N_13028,N_13093);
or U14147 (N_14147,N_13508,N_13184);
or U14148 (N_14148,N_13944,N_13670);
and U14149 (N_14149,N_13476,N_13908);
xor U14150 (N_14150,N_13307,N_13539);
and U14151 (N_14151,N_13311,N_13979);
nor U14152 (N_14152,N_13552,N_13240);
or U14153 (N_14153,N_13148,N_13661);
or U14154 (N_14154,N_13798,N_13477);
xnor U14155 (N_14155,N_13759,N_13733);
nand U14156 (N_14156,N_13363,N_13671);
and U14157 (N_14157,N_13020,N_13546);
or U14158 (N_14158,N_13836,N_13606);
xnor U14159 (N_14159,N_13772,N_13714);
or U14160 (N_14160,N_13581,N_13170);
nand U14161 (N_14161,N_13236,N_13230);
xor U14162 (N_14162,N_13748,N_13039);
nand U14163 (N_14163,N_13262,N_13927);
xnor U14164 (N_14164,N_13647,N_13468);
nor U14165 (N_14165,N_13102,N_13501);
nor U14166 (N_14166,N_13599,N_13502);
nand U14167 (N_14167,N_13100,N_13174);
xnor U14168 (N_14168,N_13774,N_13923);
nor U14169 (N_14169,N_13887,N_13068);
or U14170 (N_14170,N_13686,N_13838);
or U14171 (N_14171,N_13832,N_13133);
or U14172 (N_14172,N_13255,N_13909);
nor U14173 (N_14173,N_13678,N_13425);
and U14174 (N_14174,N_13884,N_13828);
and U14175 (N_14175,N_13084,N_13664);
or U14176 (N_14176,N_13164,N_13089);
and U14177 (N_14177,N_13640,N_13391);
nand U14178 (N_14178,N_13509,N_13726);
nor U14179 (N_14179,N_13974,N_13283);
or U14180 (N_14180,N_13566,N_13403);
and U14181 (N_14181,N_13413,N_13348);
nand U14182 (N_14182,N_13322,N_13024);
or U14183 (N_14183,N_13253,N_13620);
nand U14184 (N_14184,N_13793,N_13830);
nor U14185 (N_14185,N_13227,N_13231);
xor U14186 (N_14186,N_13059,N_13749);
nor U14187 (N_14187,N_13891,N_13101);
and U14188 (N_14188,N_13323,N_13674);
or U14189 (N_14189,N_13934,N_13122);
nor U14190 (N_14190,N_13108,N_13454);
or U14191 (N_14191,N_13392,N_13519);
or U14192 (N_14192,N_13790,N_13571);
or U14193 (N_14193,N_13308,N_13000);
nand U14194 (N_14194,N_13742,N_13795);
or U14195 (N_14195,N_13693,N_13657);
nor U14196 (N_14196,N_13032,N_13022);
nor U14197 (N_14197,N_13228,N_13775);
nor U14198 (N_14198,N_13985,N_13450);
xnor U14199 (N_14199,N_13958,N_13146);
xor U14200 (N_14200,N_13666,N_13705);
nor U14201 (N_14201,N_13452,N_13223);
nor U14202 (N_14202,N_13166,N_13899);
nor U14203 (N_14203,N_13310,N_13327);
and U14204 (N_14204,N_13339,N_13530);
or U14205 (N_14205,N_13860,N_13470);
nor U14206 (N_14206,N_13583,N_13396);
xnor U14207 (N_14207,N_13707,N_13252);
nand U14208 (N_14208,N_13268,N_13446);
nor U14209 (N_14209,N_13432,N_13644);
nand U14210 (N_14210,N_13811,N_13715);
or U14211 (N_14211,N_13538,N_13285);
nor U14212 (N_14212,N_13191,N_13438);
nor U14213 (N_14213,N_13366,N_13554);
and U14214 (N_14214,N_13895,N_13284);
and U14215 (N_14215,N_13852,N_13001);
and U14216 (N_14216,N_13196,N_13684);
or U14217 (N_14217,N_13752,N_13754);
nor U14218 (N_14218,N_13568,N_13279);
nor U14219 (N_14219,N_13136,N_13332);
nor U14220 (N_14220,N_13505,N_13969);
nor U14221 (N_14221,N_13299,N_13210);
xor U14222 (N_14222,N_13993,N_13005);
nand U14223 (N_14223,N_13026,N_13572);
xnor U14224 (N_14224,N_13789,N_13296);
xnor U14225 (N_14225,N_13197,N_13487);
nand U14226 (N_14226,N_13456,N_13637);
xor U14227 (N_14227,N_13378,N_13171);
and U14228 (N_14228,N_13764,N_13990);
and U14229 (N_14229,N_13806,N_13030);
and U14230 (N_14230,N_13954,N_13563);
and U14231 (N_14231,N_13659,N_13914);
nor U14232 (N_14232,N_13127,N_13324);
nand U14233 (N_14233,N_13453,N_13982);
and U14234 (N_14234,N_13846,N_13646);
nand U14235 (N_14235,N_13784,N_13961);
nand U14236 (N_14236,N_13097,N_13328);
or U14237 (N_14237,N_13762,N_13303);
or U14238 (N_14238,N_13369,N_13087);
and U14239 (N_14239,N_13750,N_13680);
nand U14240 (N_14240,N_13293,N_13461);
nor U14241 (N_14241,N_13445,N_13169);
nor U14242 (N_14242,N_13297,N_13229);
and U14243 (N_14243,N_13618,N_13532);
nor U14244 (N_14244,N_13935,N_13910);
nor U14245 (N_14245,N_13513,N_13485);
nor U14246 (N_14246,N_13920,N_13858);
or U14247 (N_14247,N_13198,N_13602);
nor U14248 (N_14248,N_13932,N_13594);
or U14249 (N_14249,N_13675,N_13907);
or U14250 (N_14250,N_13110,N_13325);
and U14251 (N_14251,N_13067,N_13614);
nor U14252 (N_14252,N_13444,N_13273);
nand U14253 (N_14253,N_13746,N_13999);
nand U14254 (N_14254,N_13781,N_13729);
nand U14255 (N_14255,N_13318,N_13616);
and U14256 (N_14256,N_13835,N_13739);
and U14257 (N_14257,N_13992,N_13433);
and U14258 (N_14258,N_13088,N_13531);
nand U14259 (N_14259,N_13972,N_13193);
or U14260 (N_14260,N_13724,N_13769);
and U14261 (N_14261,N_13561,N_13957);
or U14262 (N_14262,N_13866,N_13843);
nor U14263 (N_14263,N_13118,N_13009);
or U14264 (N_14264,N_13771,N_13950);
and U14265 (N_14265,N_13483,N_13528);
xor U14266 (N_14266,N_13905,N_13782);
nor U14267 (N_14267,N_13288,N_13114);
or U14268 (N_14268,N_13035,N_13863);
or U14269 (N_14269,N_13977,N_13458);
xnor U14270 (N_14270,N_13014,N_13995);
nand U14271 (N_14271,N_13371,N_13350);
nand U14272 (N_14272,N_13660,N_13794);
xnor U14273 (N_14273,N_13820,N_13725);
nor U14274 (N_14274,N_13698,N_13430);
and U14275 (N_14275,N_13272,N_13343);
and U14276 (N_14276,N_13054,N_13879);
or U14277 (N_14277,N_13219,N_13803);
nand U14278 (N_14278,N_13601,N_13994);
or U14279 (N_14279,N_13455,N_13393);
nand U14280 (N_14280,N_13722,N_13111);
and U14281 (N_14281,N_13065,N_13710);
or U14282 (N_14282,N_13527,N_13241);
nor U14283 (N_14283,N_13691,N_13217);
and U14284 (N_14284,N_13560,N_13718);
and U14285 (N_14285,N_13989,N_13897);
or U14286 (N_14286,N_13073,N_13239);
nand U14287 (N_14287,N_13521,N_13802);
xnor U14288 (N_14288,N_13204,N_13753);
or U14289 (N_14289,N_13679,N_13224);
nor U14290 (N_14290,N_13827,N_13298);
nor U14291 (N_14291,N_13479,N_13921);
and U14292 (N_14292,N_13677,N_13115);
and U14293 (N_14293,N_13149,N_13690);
nand U14294 (N_14294,N_13341,N_13906);
or U14295 (N_14295,N_13359,N_13952);
and U14296 (N_14296,N_13431,N_13492);
nand U14297 (N_14297,N_13704,N_13034);
nor U14298 (N_14298,N_13877,N_13409);
and U14299 (N_14299,N_13706,N_13094);
or U14300 (N_14300,N_13825,N_13517);
nand U14301 (N_14301,N_13956,N_13862);
nor U14302 (N_14302,N_13728,N_13147);
or U14303 (N_14303,N_13547,N_13981);
and U14304 (N_14304,N_13018,N_13808);
nand U14305 (N_14305,N_13747,N_13203);
nand U14306 (N_14306,N_13397,N_13536);
and U14307 (N_14307,N_13305,N_13058);
xnor U14308 (N_14308,N_13603,N_13548);
and U14309 (N_14309,N_13745,N_13482);
and U14310 (N_14310,N_13558,N_13326);
and U14311 (N_14311,N_13429,N_13516);
xnor U14312 (N_14312,N_13352,N_13213);
nand U14313 (N_14313,N_13962,N_13333);
and U14314 (N_14314,N_13201,N_13012);
or U14315 (N_14315,N_13449,N_13612);
and U14316 (N_14316,N_13405,N_13941);
and U14317 (N_14317,N_13427,N_13929);
nor U14318 (N_14318,N_13856,N_13007);
nor U14319 (N_14319,N_13375,N_13027);
nor U14320 (N_14320,N_13874,N_13126);
nor U14321 (N_14321,N_13973,N_13428);
and U14322 (N_14322,N_13404,N_13242);
xor U14323 (N_14323,N_13888,N_13701);
or U14324 (N_14324,N_13770,N_13038);
nand U14325 (N_14325,N_13623,N_13002);
nor U14326 (N_14326,N_13842,N_13609);
and U14327 (N_14327,N_13565,N_13633);
nor U14328 (N_14328,N_13682,N_13225);
nor U14329 (N_14329,N_13768,N_13578);
nor U14330 (N_14330,N_13786,N_13356);
xnor U14331 (N_14331,N_13340,N_13787);
and U14332 (N_14332,N_13306,N_13313);
nor U14333 (N_14333,N_13379,N_13460);
nor U14334 (N_14334,N_13329,N_13006);
nor U14335 (N_14335,N_13362,N_13544);
or U14336 (N_14336,N_13473,N_13855);
and U14337 (N_14337,N_13129,N_13893);
nor U14338 (N_14338,N_13702,N_13778);
or U14339 (N_14339,N_13367,N_13996);
xor U14340 (N_14340,N_13176,N_13758);
or U14341 (N_14341,N_13635,N_13695);
nand U14342 (N_14342,N_13885,N_13053);
and U14343 (N_14343,N_13330,N_13800);
nor U14344 (N_14344,N_13281,N_13896);
nor U14345 (N_14345,N_13490,N_13864);
or U14346 (N_14346,N_13964,N_13421);
and U14347 (N_14347,N_13949,N_13567);
nor U14348 (N_14348,N_13848,N_13116);
nor U14349 (N_14349,N_13703,N_13577);
nand U14350 (N_14350,N_13756,N_13845);
nor U14351 (N_14351,N_13902,N_13984);
and U14352 (N_14352,N_13112,N_13160);
nor U14353 (N_14353,N_13395,N_13407);
nand U14354 (N_14354,N_13172,N_13983);
or U14355 (N_14355,N_13945,N_13653);
nand U14356 (N_14356,N_13286,N_13441);
nand U14357 (N_14357,N_13040,N_13478);
nand U14358 (N_14358,N_13412,N_13069);
xnor U14359 (N_14359,N_13459,N_13457);
and U14360 (N_14360,N_13109,N_13595);
nor U14361 (N_14361,N_13290,N_13861);
or U14362 (N_14362,N_13520,N_13947);
nand U14363 (N_14363,N_13187,N_13638);
nor U14364 (N_14364,N_13186,N_13420);
or U14365 (N_14365,N_13344,N_13857);
nor U14366 (N_14366,N_13766,N_13063);
and U14367 (N_14367,N_13744,N_13336);
or U14368 (N_14368,N_13878,N_13654);
nand U14369 (N_14369,N_13731,N_13627);
or U14370 (N_14370,N_13051,N_13003);
nor U14371 (N_14371,N_13669,N_13320);
and U14372 (N_14372,N_13667,N_13448);
and U14373 (N_14373,N_13550,N_13506);
and U14374 (N_14374,N_13155,N_13625);
or U14375 (N_14375,N_13918,N_13355);
or U14376 (N_14376,N_13377,N_13824);
xor U14377 (N_14377,N_13872,N_13549);
nand U14378 (N_14378,N_13585,N_13854);
xor U14379 (N_14379,N_13346,N_13631);
nand U14380 (N_14380,N_13840,N_13946);
nand U14381 (N_14381,N_13289,N_13317);
nand U14382 (N_14382,N_13304,N_13041);
xor U14383 (N_14383,N_13955,N_13376);
and U14384 (N_14384,N_13959,N_13103);
and U14385 (N_14385,N_13434,N_13277);
and U14386 (N_14386,N_13312,N_13805);
and U14387 (N_14387,N_13256,N_13301);
and U14388 (N_14388,N_13345,N_13504);
nor U14389 (N_14389,N_13121,N_13435);
nand U14390 (N_14390,N_13222,N_13751);
xor U14391 (N_14391,N_13496,N_13804);
nand U14392 (N_14392,N_13105,N_13120);
xor U14393 (N_14393,N_13139,N_13900);
xor U14394 (N_14394,N_13757,N_13813);
and U14395 (N_14395,N_13489,N_13437);
nor U14396 (N_14396,N_13968,N_13584);
nor U14397 (N_14397,N_13079,N_13904);
nand U14398 (N_14398,N_13064,N_13106);
or U14399 (N_14399,N_13847,N_13720);
xor U14400 (N_14400,N_13592,N_13132);
nor U14401 (N_14401,N_13017,N_13124);
and U14402 (N_14402,N_13525,N_13415);
nor U14403 (N_14403,N_13066,N_13591);
nand U14404 (N_14404,N_13694,N_13406);
and U14405 (N_14405,N_13928,N_13630);
or U14406 (N_14406,N_13503,N_13865);
and U14407 (N_14407,N_13978,N_13948);
and U14408 (N_14408,N_13408,N_13372);
and U14409 (N_14409,N_13717,N_13351);
and U14410 (N_14410,N_13976,N_13075);
or U14411 (N_14411,N_13632,N_13575);
and U14412 (N_14412,N_13221,N_13316);
or U14413 (N_14413,N_13373,N_13134);
or U14414 (N_14414,N_13349,N_13251);
and U14415 (N_14415,N_13175,N_13697);
nand U14416 (N_14416,N_13142,N_13939);
nand U14417 (N_14417,N_13723,N_13086);
nor U14418 (N_14418,N_13719,N_13416);
nor U14419 (N_14419,N_13816,N_13480);
and U14420 (N_14420,N_13818,N_13465);
nor U14421 (N_14421,N_13015,N_13911);
and U14422 (N_14422,N_13104,N_13099);
nand U14423 (N_14423,N_13394,N_13082);
and U14424 (N_14424,N_13212,N_13055);
xor U14425 (N_14425,N_13190,N_13025);
nor U14426 (N_14426,N_13358,N_13368);
xor U14427 (N_14427,N_13975,N_13662);
or U14428 (N_14428,N_13997,N_13382);
nor U14429 (N_14429,N_13042,N_13113);
nand U14430 (N_14430,N_13761,N_13597);
and U14431 (N_14431,N_13335,N_13194);
or U14432 (N_14432,N_13167,N_13261);
nor U14433 (N_14433,N_13970,N_13826);
or U14434 (N_14434,N_13559,N_13886);
nor U14435 (N_14435,N_13071,N_13163);
and U14436 (N_14436,N_13141,N_13220);
and U14437 (N_14437,N_13810,N_13045);
or U14438 (N_14438,N_13850,N_13347);
or U14439 (N_14439,N_13161,N_13734);
or U14440 (N_14440,N_13922,N_13107);
xor U14441 (N_14441,N_13831,N_13250);
nand U14442 (N_14442,N_13988,N_13871);
nand U14443 (N_14443,N_13144,N_13138);
or U14444 (N_14444,N_13244,N_13711);
and U14445 (N_14445,N_13389,N_13131);
nand U14446 (N_14446,N_13683,N_13342);
nor U14447 (N_14447,N_13023,N_13564);
nor U14448 (N_14448,N_13779,N_13145);
or U14449 (N_14449,N_13628,N_13986);
or U14450 (N_14450,N_13247,N_13933);
or U14451 (N_14451,N_13915,N_13796);
nor U14452 (N_14452,N_13859,N_13043);
nand U14453 (N_14453,N_13462,N_13410);
nand U14454 (N_14454,N_13357,N_13011);
nor U14455 (N_14455,N_13019,N_13511);
or U14456 (N_14456,N_13276,N_13763);
nand U14457 (N_14457,N_13655,N_13870);
nand U14458 (N_14458,N_13314,N_13557);
and U14459 (N_14459,N_13780,N_13491);
and U14460 (N_14460,N_13205,N_13738);
nand U14461 (N_14461,N_13868,N_13543);
nor U14462 (N_14462,N_13937,N_13218);
or U14463 (N_14463,N_13991,N_13555);
nand U14464 (N_14464,N_13507,N_13665);
nor U14465 (N_14465,N_13248,N_13634);
or U14466 (N_14466,N_13046,N_13337);
or U14467 (N_14467,N_13912,N_13245);
and U14468 (N_14468,N_13639,N_13785);
nand U14469 (N_14469,N_13587,N_13013);
nor U14470 (N_14470,N_13309,N_13044);
and U14471 (N_14471,N_13645,N_13586);
nand U14472 (N_14472,N_13641,N_13512);
or U14473 (N_14473,N_13687,N_13423);
and U14474 (N_14474,N_13202,N_13611);
and U14475 (N_14475,N_13882,N_13699);
or U14476 (N_14476,N_13474,N_13925);
or U14477 (N_14477,N_13834,N_13869);
and U14478 (N_14478,N_13619,N_13807);
nor U14479 (N_14479,N_13689,N_13841);
or U14480 (N_14480,N_13656,N_13257);
and U14481 (N_14481,N_13270,N_13484);
or U14482 (N_14482,N_13676,N_13626);
nor U14483 (N_14483,N_13963,N_13890);
or U14484 (N_14484,N_13200,N_13294);
nand U14485 (N_14485,N_13610,N_13853);
or U14486 (N_14486,N_13162,N_13292);
nand U14487 (N_14487,N_13049,N_13235);
or U14488 (N_14488,N_13938,N_13180);
nor U14489 (N_14489,N_13696,N_13178);
nor U14490 (N_14490,N_13791,N_13189);
nor U14491 (N_14491,N_13649,N_13913);
nand U14492 (N_14492,N_13916,N_13822);
nor U14493 (N_14493,N_13380,N_13672);
and U14494 (N_14494,N_13008,N_13600);
or U14495 (N_14495,N_13384,N_13037);
nand U14496 (N_14496,N_13924,N_13545);
xor U14497 (N_14497,N_13265,N_13533);
nor U14498 (N_14498,N_13658,N_13287);
or U14499 (N_14499,N_13331,N_13713);
and U14500 (N_14500,N_13158,N_13449);
nand U14501 (N_14501,N_13388,N_13780);
nand U14502 (N_14502,N_13986,N_13515);
and U14503 (N_14503,N_13118,N_13399);
xor U14504 (N_14504,N_13215,N_13933);
nand U14505 (N_14505,N_13276,N_13442);
nor U14506 (N_14506,N_13462,N_13033);
nor U14507 (N_14507,N_13584,N_13738);
nand U14508 (N_14508,N_13491,N_13223);
or U14509 (N_14509,N_13332,N_13679);
and U14510 (N_14510,N_13233,N_13126);
nand U14511 (N_14511,N_13973,N_13937);
or U14512 (N_14512,N_13960,N_13587);
and U14513 (N_14513,N_13679,N_13538);
xnor U14514 (N_14514,N_13752,N_13305);
and U14515 (N_14515,N_13189,N_13515);
nor U14516 (N_14516,N_13375,N_13846);
nor U14517 (N_14517,N_13591,N_13108);
and U14518 (N_14518,N_13672,N_13444);
nor U14519 (N_14519,N_13949,N_13243);
nand U14520 (N_14520,N_13388,N_13279);
or U14521 (N_14521,N_13908,N_13100);
or U14522 (N_14522,N_13007,N_13158);
and U14523 (N_14523,N_13272,N_13957);
or U14524 (N_14524,N_13678,N_13167);
and U14525 (N_14525,N_13957,N_13412);
nor U14526 (N_14526,N_13294,N_13026);
nor U14527 (N_14527,N_13171,N_13119);
nor U14528 (N_14528,N_13664,N_13493);
nand U14529 (N_14529,N_13773,N_13286);
nand U14530 (N_14530,N_13833,N_13322);
xor U14531 (N_14531,N_13852,N_13664);
nor U14532 (N_14532,N_13182,N_13835);
or U14533 (N_14533,N_13636,N_13318);
xnor U14534 (N_14534,N_13750,N_13069);
nand U14535 (N_14535,N_13776,N_13113);
and U14536 (N_14536,N_13194,N_13528);
nor U14537 (N_14537,N_13149,N_13133);
or U14538 (N_14538,N_13346,N_13054);
or U14539 (N_14539,N_13120,N_13856);
or U14540 (N_14540,N_13179,N_13842);
xnor U14541 (N_14541,N_13366,N_13412);
and U14542 (N_14542,N_13181,N_13020);
or U14543 (N_14543,N_13168,N_13559);
or U14544 (N_14544,N_13838,N_13833);
or U14545 (N_14545,N_13378,N_13688);
or U14546 (N_14546,N_13452,N_13095);
nor U14547 (N_14547,N_13885,N_13477);
nand U14548 (N_14548,N_13293,N_13956);
nand U14549 (N_14549,N_13746,N_13814);
or U14550 (N_14550,N_13355,N_13762);
xnor U14551 (N_14551,N_13851,N_13528);
or U14552 (N_14552,N_13111,N_13485);
nor U14553 (N_14553,N_13106,N_13785);
xnor U14554 (N_14554,N_13239,N_13269);
nor U14555 (N_14555,N_13570,N_13838);
nand U14556 (N_14556,N_13450,N_13672);
xor U14557 (N_14557,N_13698,N_13965);
and U14558 (N_14558,N_13525,N_13882);
or U14559 (N_14559,N_13597,N_13018);
nor U14560 (N_14560,N_13804,N_13056);
nor U14561 (N_14561,N_13157,N_13430);
and U14562 (N_14562,N_13809,N_13319);
and U14563 (N_14563,N_13402,N_13747);
nand U14564 (N_14564,N_13312,N_13619);
nand U14565 (N_14565,N_13580,N_13117);
or U14566 (N_14566,N_13848,N_13705);
or U14567 (N_14567,N_13091,N_13639);
and U14568 (N_14568,N_13346,N_13300);
nor U14569 (N_14569,N_13055,N_13628);
nand U14570 (N_14570,N_13234,N_13823);
and U14571 (N_14571,N_13522,N_13542);
and U14572 (N_14572,N_13549,N_13536);
or U14573 (N_14573,N_13128,N_13641);
or U14574 (N_14574,N_13261,N_13276);
and U14575 (N_14575,N_13450,N_13036);
or U14576 (N_14576,N_13124,N_13935);
or U14577 (N_14577,N_13268,N_13183);
nand U14578 (N_14578,N_13594,N_13589);
or U14579 (N_14579,N_13667,N_13808);
and U14580 (N_14580,N_13064,N_13417);
nor U14581 (N_14581,N_13308,N_13083);
and U14582 (N_14582,N_13119,N_13340);
nand U14583 (N_14583,N_13571,N_13832);
xor U14584 (N_14584,N_13326,N_13114);
xor U14585 (N_14585,N_13610,N_13167);
nand U14586 (N_14586,N_13917,N_13481);
nand U14587 (N_14587,N_13109,N_13705);
and U14588 (N_14588,N_13067,N_13694);
nor U14589 (N_14589,N_13628,N_13770);
nor U14590 (N_14590,N_13372,N_13367);
nor U14591 (N_14591,N_13503,N_13903);
xnor U14592 (N_14592,N_13203,N_13746);
and U14593 (N_14593,N_13970,N_13305);
and U14594 (N_14594,N_13076,N_13649);
nand U14595 (N_14595,N_13280,N_13104);
or U14596 (N_14596,N_13416,N_13893);
and U14597 (N_14597,N_13183,N_13650);
nor U14598 (N_14598,N_13044,N_13705);
nor U14599 (N_14599,N_13837,N_13704);
nand U14600 (N_14600,N_13656,N_13960);
or U14601 (N_14601,N_13235,N_13263);
or U14602 (N_14602,N_13685,N_13203);
or U14603 (N_14603,N_13921,N_13884);
and U14604 (N_14604,N_13710,N_13169);
xnor U14605 (N_14605,N_13615,N_13218);
nor U14606 (N_14606,N_13350,N_13057);
and U14607 (N_14607,N_13426,N_13436);
xor U14608 (N_14608,N_13497,N_13599);
nand U14609 (N_14609,N_13774,N_13341);
nor U14610 (N_14610,N_13467,N_13479);
nor U14611 (N_14611,N_13438,N_13294);
nor U14612 (N_14612,N_13692,N_13113);
and U14613 (N_14613,N_13267,N_13157);
and U14614 (N_14614,N_13179,N_13987);
nor U14615 (N_14615,N_13065,N_13836);
and U14616 (N_14616,N_13855,N_13739);
nor U14617 (N_14617,N_13213,N_13575);
xnor U14618 (N_14618,N_13630,N_13786);
or U14619 (N_14619,N_13273,N_13146);
nor U14620 (N_14620,N_13017,N_13804);
and U14621 (N_14621,N_13117,N_13654);
or U14622 (N_14622,N_13240,N_13674);
nand U14623 (N_14623,N_13295,N_13836);
nor U14624 (N_14624,N_13106,N_13364);
xor U14625 (N_14625,N_13021,N_13961);
nand U14626 (N_14626,N_13190,N_13835);
nand U14627 (N_14627,N_13729,N_13089);
xnor U14628 (N_14628,N_13372,N_13505);
and U14629 (N_14629,N_13340,N_13175);
xnor U14630 (N_14630,N_13999,N_13933);
and U14631 (N_14631,N_13454,N_13244);
or U14632 (N_14632,N_13016,N_13949);
and U14633 (N_14633,N_13531,N_13174);
nor U14634 (N_14634,N_13783,N_13569);
nor U14635 (N_14635,N_13166,N_13996);
nor U14636 (N_14636,N_13024,N_13421);
or U14637 (N_14637,N_13459,N_13443);
nor U14638 (N_14638,N_13919,N_13055);
and U14639 (N_14639,N_13207,N_13383);
nor U14640 (N_14640,N_13755,N_13215);
nand U14641 (N_14641,N_13617,N_13065);
or U14642 (N_14642,N_13413,N_13983);
xnor U14643 (N_14643,N_13220,N_13994);
xor U14644 (N_14644,N_13416,N_13329);
or U14645 (N_14645,N_13869,N_13359);
or U14646 (N_14646,N_13026,N_13199);
xnor U14647 (N_14647,N_13207,N_13630);
or U14648 (N_14648,N_13327,N_13091);
xnor U14649 (N_14649,N_13725,N_13219);
nor U14650 (N_14650,N_13085,N_13124);
and U14651 (N_14651,N_13526,N_13087);
or U14652 (N_14652,N_13035,N_13125);
nand U14653 (N_14653,N_13843,N_13003);
and U14654 (N_14654,N_13404,N_13561);
and U14655 (N_14655,N_13001,N_13152);
nor U14656 (N_14656,N_13977,N_13031);
and U14657 (N_14657,N_13596,N_13311);
and U14658 (N_14658,N_13974,N_13741);
nor U14659 (N_14659,N_13330,N_13411);
xor U14660 (N_14660,N_13963,N_13269);
and U14661 (N_14661,N_13243,N_13596);
xor U14662 (N_14662,N_13274,N_13462);
xor U14663 (N_14663,N_13171,N_13859);
and U14664 (N_14664,N_13826,N_13325);
nand U14665 (N_14665,N_13080,N_13333);
nand U14666 (N_14666,N_13678,N_13834);
nor U14667 (N_14667,N_13346,N_13718);
or U14668 (N_14668,N_13862,N_13865);
or U14669 (N_14669,N_13245,N_13683);
nand U14670 (N_14670,N_13947,N_13189);
nand U14671 (N_14671,N_13085,N_13721);
nor U14672 (N_14672,N_13678,N_13149);
and U14673 (N_14673,N_13788,N_13107);
nand U14674 (N_14674,N_13158,N_13530);
and U14675 (N_14675,N_13351,N_13651);
nor U14676 (N_14676,N_13291,N_13917);
or U14677 (N_14677,N_13536,N_13555);
or U14678 (N_14678,N_13452,N_13774);
and U14679 (N_14679,N_13540,N_13301);
xor U14680 (N_14680,N_13420,N_13710);
nor U14681 (N_14681,N_13909,N_13350);
nand U14682 (N_14682,N_13391,N_13724);
or U14683 (N_14683,N_13120,N_13521);
or U14684 (N_14684,N_13920,N_13567);
and U14685 (N_14685,N_13388,N_13786);
and U14686 (N_14686,N_13511,N_13790);
or U14687 (N_14687,N_13976,N_13146);
or U14688 (N_14688,N_13153,N_13195);
or U14689 (N_14689,N_13772,N_13671);
xnor U14690 (N_14690,N_13542,N_13507);
or U14691 (N_14691,N_13135,N_13083);
xnor U14692 (N_14692,N_13321,N_13412);
nor U14693 (N_14693,N_13835,N_13408);
or U14694 (N_14694,N_13610,N_13948);
nand U14695 (N_14695,N_13489,N_13668);
or U14696 (N_14696,N_13411,N_13119);
nand U14697 (N_14697,N_13851,N_13920);
and U14698 (N_14698,N_13893,N_13566);
nand U14699 (N_14699,N_13517,N_13544);
or U14700 (N_14700,N_13521,N_13716);
nand U14701 (N_14701,N_13202,N_13786);
nand U14702 (N_14702,N_13266,N_13342);
and U14703 (N_14703,N_13448,N_13421);
or U14704 (N_14704,N_13368,N_13396);
nand U14705 (N_14705,N_13254,N_13666);
nand U14706 (N_14706,N_13111,N_13219);
nand U14707 (N_14707,N_13919,N_13588);
nor U14708 (N_14708,N_13871,N_13424);
and U14709 (N_14709,N_13008,N_13804);
and U14710 (N_14710,N_13893,N_13249);
nand U14711 (N_14711,N_13347,N_13059);
or U14712 (N_14712,N_13606,N_13853);
or U14713 (N_14713,N_13914,N_13918);
nor U14714 (N_14714,N_13562,N_13833);
and U14715 (N_14715,N_13385,N_13811);
or U14716 (N_14716,N_13796,N_13649);
xnor U14717 (N_14717,N_13673,N_13739);
or U14718 (N_14718,N_13903,N_13249);
nand U14719 (N_14719,N_13876,N_13896);
nand U14720 (N_14720,N_13766,N_13488);
nor U14721 (N_14721,N_13954,N_13425);
nor U14722 (N_14722,N_13901,N_13131);
nor U14723 (N_14723,N_13488,N_13494);
xnor U14724 (N_14724,N_13272,N_13534);
and U14725 (N_14725,N_13035,N_13773);
and U14726 (N_14726,N_13095,N_13935);
nand U14727 (N_14727,N_13603,N_13233);
or U14728 (N_14728,N_13147,N_13572);
nor U14729 (N_14729,N_13843,N_13291);
and U14730 (N_14730,N_13290,N_13156);
nor U14731 (N_14731,N_13881,N_13512);
and U14732 (N_14732,N_13166,N_13681);
nand U14733 (N_14733,N_13447,N_13738);
and U14734 (N_14734,N_13222,N_13481);
nor U14735 (N_14735,N_13165,N_13760);
nor U14736 (N_14736,N_13240,N_13119);
nor U14737 (N_14737,N_13613,N_13155);
nand U14738 (N_14738,N_13225,N_13777);
and U14739 (N_14739,N_13258,N_13733);
and U14740 (N_14740,N_13798,N_13372);
nor U14741 (N_14741,N_13907,N_13240);
nand U14742 (N_14742,N_13222,N_13398);
nand U14743 (N_14743,N_13777,N_13201);
xor U14744 (N_14744,N_13457,N_13018);
nand U14745 (N_14745,N_13549,N_13803);
nor U14746 (N_14746,N_13837,N_13240);
and U14747 (N_14747,N_13156,N_13467);
and U14748 (N_14748,N_13400,N_13530);
or U14749 (N_14749,N_13479,N_13900);
nand U14750 (N_14750,N_13328,N_13262);
or U14751 (N_14751,N_13088,N_13682);
nor U14752 (N_14752,N_13101,N_13464);
nor U14753 (N_14753,N_13430,N_13681);
nand U14754 (N_14754,N_13384,N_13063);
nor U14755 (N_14755,N_13649,N_13167);
or U14756 (N_14756,N_13306,N_13842);
and U14757 (N_14757,N_13915,N_13671);
xor U14758 (N_14758,N_13261,N_13786);
nand U14759 (N_14759,N_13699,N_13103);
nand U14760 (N_14760,N_13587,N_13885);
nand U14761 (N_14761,N_13219,N_13526);
and U14762 (N_14762,N_13006,N_13390);
or U14763 (N_14763,N_13208,N_13788);
xor U14764 (N_14764,N_13486,N_13077);
nor U14765 (N_14765,N_13830,N_13119);
xor U14766 (N_14766,N_13742,N_13474);
and U14767 (N_14767,N_13847,N_13700);
nand U14768 (N_14768,N_13878,N_13160);
nand U14769 (N_14769,N_13449,N_13566);
and U14770 (N_14770,N_13952,N_13691);
nor U14771 (N_14771,N_13175,N_13716);
or U14772 (N_14772,N_13273,N_13628);
nor U14773 (N_14773,N_13868,N_13020);
and U14774 (N_14774,N_13530,N_13585);
and U14775 (N_14775,N_13705,N_13690);
xnor U14776 (N_14776,N_13972,N_13275);
xor U14777 (N_14777,N_13287,N_13672);
xnor U14778 (N_14778,N_13730,N_13022);
nor U14779 (N_14779,N_13035,N_13761);
xor U14780 (N_14780,N_13304,N_13515);
nor U14781 (N_14781,N_13667,N_13628);
nand U14782 (N_14782,N_13088,N_13272);
nand U14783 (N_14783,N_13369,N_13923);
and U14784 (N_14784,N_13089,N_13524);
xnor U14785 (N_14785,N_13165,N_13370);
xor U14786 (N_14786,N_13408,N_13314);
and U14787 (N_14787,N_13979,N_13253);
nand U14788 (N_14788,N_13013,N_13958);
and U14789 (N_14789,N_13873,N_13858);
nor U14790 (N_14790,N_13822,N_13562);
nand U14791 (N_14791,N_13298,N_13637);
nor U14792 (N_14792,N_13848,N_13867);
nor U14793 (N_14793,N_13550,N_13637);
and U14794 (N_14794,N_13003,N_13111);
nor U14795 (N_14795,N_13160,N_13551);
or U14796 (N_14796,N_13551,N_13323);
nand U14797 (N_14797,N_13486,N_13515);
nor U14798 (N_14798,N_13822,N_13258);
or U14799 (N_14799,N_13908,N_13200);
nor U14800 (N_14800,N_13879,N_13692);
nor U14801 (N_14801,N_13192,N_13290);
xnor U14802 (N_14802,N_13040,N_13614);
nor U14803 (N_14803,N_13478,N_13508);
or U14804 (N_14804,N_13190,N_13339);
and U14805 (N_14805,N_13424,N_13920);
and U14806 (N_14806,N_13184,N_13613);
nor U14807 (N_14807,N_13231,N_13041);
or U14808 (N_14808,N_13579,N_13100);
nand U14809 (N_14809,N_13026,N_13292);
or U14810 (N_14810,N_13316,N_13528);
or U14811 (N_14811,N_13635,N_13579);
or U14812 (N_14812,N_13855,N_13896);
or U14813 (N_14813,N_13474,N_13493);
nand U14814 (N_14814,N_13761,N_13530);
and U14815 (N_14815,N_13471,N_13865);
or U14816 (N_14816,N_13601,N_13116);
and U14817 (N_14817,N_13866,N_13932);
nand U14818 (N_14818,N_13023,N_13410);
and U14819 (N_14819,N_13526,N_13816);
nor U14820 (N_14820,N_13866,N_13134);
nor U14821 (N_14821,N_13795,N_13754);
nand U14822 (N_14822,N_13835,N_13969);
or U14823 (N_14823,N_13582,N_13664);
nand U14824 (N_14824,N_13025,N_13151);
and U14825 (N_14825,N_13521,N_13871);
nor U14826 (N_14826,N_13481,N_13543);
and U14827 (N_14827,N_13107,N_13874);
nand U14828 (N_14828,N_13631,N_13909);
nand U14829 (N_14829,N_13315,N_13515);
nor U14830 (N_14830,N_13415,N_13744);
nor U14831 (N_14831,N_13891,N_13362);
nand U14832 (N_14832,N_13375,N_13754);
xor U14833 (N_14833,N_13166,N_13299);
or U14834 (N_14834,N_13382,N_13064);
and U14835 (N_14835,N_13802,N_13229);
nand U14836 (N_14836,N_13925,N_13138);
and U14837 (N_14837,N_13392,N_13821);
xnor U14838 (N_14838,N_13357,N_13738);
and U14839 (N_14839,N_13318,N_13151);
nand U14840 (N_14840,N_13017,N_13572);
and U14841 (N_14841,N_13170,N_13709);
and U14842 (N_14842,N_13858,N_13119);
nor U14843 (N_14843,N_13092,N_13737);
xor U14844 (N_14844,N_13868,N_13075);
nor U14845 (N_14845,N_13652,N_13734);
or U14846 (N_14846,N_13735,N_13970);
nor U14847 (N_14847,N_13979,N_13842);
and U14848 (N_14848,N_13500,N_13836);
nand U14849 (N_14849,N_13898,N_13666);
nand U14850 (N_14850,N_13749,N_13796);
nor U14851 (N_14851,N_13650,N_13528);
or U14852 (N_14852,N_13210,N_13845);
xnor U14853 (N_14853,N_13792,N_13130);
and U14854 (N_14854,N_13578,N_13554);
nor U14855 (N_14855,N_13447,N_13147);
and U14856 (N_14856,N_13424,N_13712);
nand U14857 (N_14857,N_13250,N_13341);
and U14858 (N_14858,N_13639,N_13310);
nor U14859 (N_14859,N_13020,N_13790);
nand U14860 (N_14860,N_13368,N_13667);
and U14861 (N_14861,N_13758,N_13156);
nand U14862 (N_14862,N_13112,N_13349);
or U14863 (N_14863,N_13499,N_13425);
nand U14864 (N_14864,N_13105,N_13213);
or U14865 (N_14865,N_13214,N_13305);
or U14866 (N_14866,N_13410,N_13885);
nor U14867 (N_14867,N_13713,N_13428);
and U14868 (N_14868,N_13165,N_13759);
and U14869 (N_14869,N_13997,N_13089);
nor U14870 (N_14870,N_13719,N_13806);
or U14871 (N_14871,N_13211,N_13327);
or U14872 (N_14872,N_13398,N_13418);
nand U14873 (N_14873,N_13153,N_13491);
nand U14874 (N_14874,N_13345,N_13068);
nor U14875 (N_14875,N_13812,N_13062);
nand U14876 (N_14876,N_13001,N_13681);
nand U14877 (N_14877,N_13151,N_13584);
nor U14878 (N_14878,N_13015,N_13751);
nand U14879 (N_14879,N_13750,N_13366);
nor U14880 (N_14880,N_13853,N_13755);
nand U14881 (N_14881,N_13373,N_13632);
xnor U14882 (N_14882,N_13825,N_13392);
nand U14883 (N_14883,N_13715,N_13823);
nor U14884 (N_14884,N_13176,N_13894);
nor U14885 (N_14885,N_13471,N_13278);
nor U14886 (N_14886,N_13749,N_13964);
or U14887 (N_14887,N_13362,N_13063);
xor U14888 (N_14888,N_13197,N_13294);
nor U14889 (N_14889,N_13948,N_13996);
nand U14890 (N_14890,N_13533,N_13514);
nor U14891 (N_14891,N_13214,N_13797);
nor U14892 (N_14892,N_13129,N_13677);
nand U14893 (N_14893,N_13236,N_13613);
and U14894 (N_14894,N_13824,N_13807);
or U14895 (N_14895,N_13804,N_13807);
nor U14896 (N_14896,N_13476,N_13799);
nor U14897 (N_14897,N_13154,N_13097);
xor U14898 (N_14898,N_13802,N_13528);
nor U14899 (N_14899,N_13447,N_13904);
xor U14900 (N_14900,N_13365,N_13706);
and U14901 (N_14901,N_13427,N_13540);
nand U14902 (N_14902,N_13273,N_13586);
xor U14903 (N_14903,N_13482,N_13004);
xor U14904 (N_14904,N_13556,N_13966);
nor U14905 (N_14905,N_13574,N_13914);
and U14906 (N_14906,N_13959,N_13756);
nor U14907 (N_14907,N_13344,N_13644);
nor U14908 (N_14908,N_13196,N_13367);
xor U14909 (N_14909,N_13323,N_13868);
nand U14910 (N_14910,N_13004,N_13020);
nand U14911 (N_14911,N_13698,N_13921);
and U14912 (N_14912,N_13764,N_13942);
xnor U14913 (N_14913,N_13975,N_13559);
and U14914 (N_14914,N_13907,N_13876);
and U14915 (N_14915,N_13804,N_13894);
and U14916 (N_14916,N_13051,N_13305);
or U14917 (N_14917,N_13970,N_13273);
xor U14918 (N_14918,N_13985,N_13610);
nor U14919 (N_14919,N_13064,N_13583);
nor U14920 (N_14920,N_13422,N_13374);
and U14921 (N_14921,N_13640,N_13803);
nor U14922 (N_14922,N_13718,N_13278);
and U14923 (N_14923,N_13610,N_13218);
nand U14924 (N_14924,N_13731,N_13450);
nand U14925 (N_14925,N_13507,N_13866);
or U14926 (N_14926,N_13593,N_13104);
nand U14927 (N_14927,N_13944,N_13734);
nand U14928 (N_14928,N_13856,N_13334);
or U14929 (N_14929,N_13559,N_13634);
xor U14930 (N_14930,N_13888,N_13854);
or U14931 (N_14931,N_13058,N_13051);
nor U14932 (N_14932,N_13702,N_13300);
xnor U14933 (N_14933,N_13355,N_13296);
nor U14934 (N_14934,N_13344,N_13127);
or U14935 (N_14935,N_13274,N_13016);
xnor U14936 (N_14936,N_13523,N_13383);
nor U14937 (N_14937,N_13858,N_13583);
nor U14938 (N_14938,N_13816,N_13575);
nand U14939 (N_14939,N_13259,N_13682);
or U14940 (N_14940,N_13927,N_13246);
nor U14941 (N_14941,N_13869,N_13884);
nor U14942 (N_14942,N_13641,N_13183);
nand U14943 (N_14943,N_13035,N_13305);
or U14944 (N_14944,N_13475,N_13980);
nor U14945 (N_14945,N_13894,N_13650);
or U14946 (N_14946,N_13685,N_13874);
and U14947 (N_14947,N_13936,N_13437);
and U14948 (N_14948,N_13793,N_13498);
nand U14949 (N_14949,N_13839,N_13460);
nor U14950 (N_14950,N_13077,N_13190);
nor U14951 (N_14951,N_13411,N_13061);
nor U14952 (N_14952,N_13551,N_13726);
nor U14953 (N_14953,N_13015,N_13769);
or U14954 (N_14954,N_13436,N_13140);
nor U14955 (N_14955,N_13189,N_13010);
and U14956 (N_14956,N_13163,N_13687);
and U14957 (N_14957,N_13484,N_13564);
nand U14958 (N_14958,N_13535,N_13747);
or U14959 (N_14959,N_13210,N_13395);
or U14960 (N_14960,N_13323,N_13519);
nand U14961 (N_14961,N_13416,N_13927);
and U14962 (N_14962,N_13953,N_13852);
and U14963 (N_14963,N_13693,N_13246);
or U14964 (N_14964,N_13477,N_13647);
xor U14965 (N_14965,N_13821,N_13292);
xor U14966 (N_14966,N_13833,N_13310);
nand U14967 (N_14967,N_13020,N_13256);
and U14968 (N_14968,N_13908,N_13542);
or U14969 (N_14969,N_13663,N_13847);
nor U14970 (N_14970,N_13724,N_13185);
xor U14971 (N_14971,N_13180,N_13904);
nand U14972 (N_14972,N_13851,N_13953);
nor U14973 (N_14973,N_13676,N_13983);
xnor U14974 (N_14974,N_13559,N_13009);
nor U14975 (N_14975,N_13433,N_13346);
xnor U14976 (N_14976,N_13728,N_13923);
or U14977 (N_14977,N_13167,N_13528);
and U14978 (N_14978,N_13912,N_13097);
and U14979 (N_14979,N_13539,N_13624);
xor U14980 (N_14980,N_13135,N_13254);
nor U14981 (N_14981,N_13096,N_13791);
or U14982 (N_14982,N_13089,N_13067);
or U14983 (N_14983,N_13116,N_13795);
nor U14984 (N_14984,N_13972,N_13662);
or U14985 (N_14985,N_13282,N_13599);
or U14986 (N_14986,N_13459,N_13197);
or U14987 (N_14987,N_13897,N_13393);
nor U14988 (N_14988,N_13143,N_13922);
and U14989 (N_14989,N_13059,N_13110);
nor U14990 (N_14990,N_13540,N_13750);
or U14991 (N_14991,N_13888,N_13782);
nand U14992 (N_14992,N_13761,N_13648);
nand U14993 (N_14993,N_13371,N_13356);
or U14994 (N_14994,N_13337,N_13220);
and U14995 (N_14995,N_13730,N_13480);
nor U14996 (N_14996,N_13109,N_13201);
nand U14997 (N_14997,N_13124,N_13459);
nor U14998 (N_14998,N_13207,N_13391);
nand U14999 (N_14999,N_13402,N_13277);
xor UO_0 (O_0,N_14161,N_14565);
and UO_1 (O_1,N_14517,N_14152);
nor UO_2 (O_2,N_14809,N_14531);
nand UO_3 (O_3,N_14770,N_14082);
xor UO_4 (O_4,N_14042,N_14114);
nor UO_5 (O_5,N_14244,N_14110);
nand UO_6 (O_6,N_14991,N_14045);
or UO_7 (O_7,N_14941,N_14858);
and UO_8 (O_8,N_14599,N_14625);
and UO_9 (O_9,N_14254,N_14654);
or UO_10 (O_10,N_14894,N_14495);
nor UO_11 (O_11,N_14125,N_14060);
and UO_12 (O_12,N_14791,N_14111);
or UO_13 (O_13,N_14198,N_14616);
nand UO_14 (O_14,N_14221,N_14689);
nor UO_15 (O_15,N_14106,N_14996);
and UO_16 (O_16,N_14573,N_14799);
or UO_17 (O_17,N_14721,N_14231);
nand UO_18 (O_18,N_14930,N_14609);
nand UO_19 (O_19,N_14406,N_14031);
nand UO_20 (O_20,N_14344,N_14168);
nand UO_21 (O_21,N_14132,N_14300);
nand UO_22 (O_22,N_14632,N_14690);
or UO_23 (O_23,N_14462,N_14157);
xnor UO_24 (O_24,N_14897,N_14141);
and UO_25 (O_25,N_14765,N_14054);
and UO_26 (O_26,N_14988,N_14435);
nor UO_27 (O_27,N_14730,N_14960);
xnor UO_28 (O_28,N_14425,N_14171);
nand UO_29 (O_29,N_14493,N_14744);
or UO_30 (O_30,N_14113,N_14541);
or UO_31 (O_31,N_14257,N_14685);
nor UO_32 (O_32,N_14698,N_14888);
xnor UO_33 (O_33,N_14557,N_14306);
and UO_34 (O_34,N_14145,N_14269);
nor UO_35 (O_35,N_14592,N_14128);
and UO_36 (O_36,N_14445,N_14709);
nor UO_37 (O_37,N_14334,N_14240);
or UO_38 (O_38,N_14547,N_14696);
xor UO_39 (O_39,N_14562,N_14749);
nand UO_40 (O_40,N_14478,N_14933);
and UO_41 (O_41,N_14922,N_14348);
and UO_42 (O_42,N_14188,N_14220);
and UO_43 (O_43,N_14838,N_14475);
nand UO_44 (O_44,N_14309,N_14596);
nor UO_45 (O_45,N_14326,N_14673);
or UO_46 (O_46,N_14852,N_14041);
or UO_47 (O_47,N_14528,N_14539);
nor UO_48 (O_48,N_14232,N_14661);
or UO_49 (O_49,N_14426,N_14669);
and UO_50 (O_50,N_14787,N_14369);
xor UO_51 (O_51,N_14663,N_14280);
and UO_52 (O_52,N_14999,N_14164);
and UO_53 (O_53,N_14259,N_14497);
and UO_54 (O_54,N_14238,N_14359);
and UO_55 (O_55,N_14830,N_14252);
nor UO_56 (O_56,N_14291,N_14849);
xor UO_57 (O_57,N_14627,N_14750);
or UO_58 (O_58,N_14071,N_14803);
nand UO_59 (O_59,N_14078,N_14525);
nor UO_60 (O_60,N_14199,N_14590);
nand UO_61 (O_61,N_14962,N_14030);
nand UO_62 (O_62,N_14467,N_14998);
or UO_63 (O_63,N_14835,N_14583);
and UO_64 (O_64,N_14024,N_14346);
nor UO_65 (O_65,N_14647,N_14239);
xor UO_66 (O_66,N_14226,N_14107);
nor UO_67 (O_67,N_14969,N_14453);
nand UO_68 (O_68,N_14458,N_14289);
nor UO_69 (O_69,N_14368,N_14470);
xnor UO_70 (O_70,N_14247,N_14190);
and UO_71 (O_71,N_14511,N_14405);
and UO_72 (O_72,N_14800,N_14595);
xnor UO_73 (O_73,N_14513,N_14354);
and UO_74 (O_74,N_14544,N_14575);
nor UO_75 (O_75,N_14092,N_14299);
nand UO_76 (O_76,N_14798,N_14169);
and UO_77 (O_77,N_14938,N_14095);
nand UO_78 (O_78,N_14964,N_14695);
nand UO_79 (O_79,N_14755,N_14260);
nand UO_80 (O_80,N_14437,N_14452);
or UO_81 (O_81,N_14454,N_14699);
nand UO_82 (O_82,N_14570,N_14811);
or UO_83 (O_83,N_14841,N_14913);
nand UO_84 (O_84,N_14711,N_14653);
and UO_85 (O_85,N_14408,N_14372);
or UO_86 (O_86,N_14958,N_14485);
nand UO_87 (O_87,N_14498,N_14973);
and UO_88 (O_88,N_14006,N_14477);
nor UO_89 (O_89,N_14449,N_14637);
xnor UO_90 (O_90,N_14923,N_14581);
or UO_91 (O_91,N_14831,N_14754);
nand UO_92 (O_92,N_14196,N_14651);
and UO_93 (O_93,N_14481,N_14116);
nand UO_94 (O_94,N_14055,N_14277);
nand UO_95 (O_95,N_14182,N_14777);
nand UO_96 (O_96,N_14068,N_14314);
and UO_97 (O_97,N_14223,N_14686);
nor UO_98 (O_98,N_14212,N_14717);
and UO_99 (O_99,N_14684,N_14812);
nand UO_100 (O_100,N_14332,N_14615);
nor UO_101 (O_101,N_14605,N_14586);
or UO_102 (O_102,N_14619,N_14568);
nor UO_103 (O_103,N_14886,N_14965);
and UO_104 (O_104,N_14028,N_14139);
or UO_105 (O_105,N_14476,N_14856);
and UO_106 (O_106,N_14402,N_14211);
and UO_107 (O_107,N_14648,N_14644);
xor UO_108 (O_108,N_14026,N_14771);
and UO_109 (O_109,N_14207,N_14620);
or UO_110 (O_110,N_14558,N_14526);
nor UO_111 (O_111,N_14967,N_14303);
nor UO_112 (O_112,N_14316,N_14392);
or UO_113 (O_113,N_14665,N_14455);
nand UO_114 (O_114,N_14482,N_14763);
and UO_115 (O_115,N_14912,N_14708);
nand UO_116 (O_116,N_14639,N_14117);
xnor UO_117 (O_117,N_14086,N_14154);
and UO_118 (O_118,N_14155,N_14379);
and UO_119 (O_119,N_14694,N_14712);
xnor UO_120 (O_120,N_14138,N_14726);
nor UO_121 (O_121,N_14178,N_14918);
or UO_122 (O_122,N_14889,N_14255);
nor UO_123 (O_123,N_14412,N_14905);
or UO_124 (O_124,N_14384,N_14347);
nand UO_125 (O_125,N_14263,N_14275);
nand UO_126 (O_126,N_14911,N_14807);
or UO_127 (O_127,N_14735,N_14268);
and UO_128 (O_128,N_14075,N_14725);
nand UO_129 (O_129,N_14954,N_14740);
xor UO_130 (O_130,N_14772,N_14366);
xnor UO_131 (O_131,N_14414,N_14782);
xor UO_132 (O_132,N_14785,N_14003);
nor UO_133 (O_133,N_14465,N_14135);
nand UO_134 (O_134,N_14457,N_14992);
and UO_135 (O_135,N_14084,N_14046);
or UO_136 (O_136,N_14410,N_14939);
and UO_137 (O_137,N_14025,N_14192);
nand UO_138 (O_138,N_14503,N_14404);
nor UO_139 (O_139,N_14707,N_14146);
and UO_140 (O_140,N_14950,N_14987);
nand UO_141 (O_141,N_14387,N_14403);
xnor UO_142 (O_142,N_14191,N_14201);
nor UO_143 (O_143,N_14472,N_14824);
or UO_144 (O_144,N_14937,N_14052);
and UO_145 (O_145,N_14716,N_14091);
nor UO_146 (O_146,N_14446,N_14459);
and UO_147 (O_147,N_14500,N_14502);
nand UO_148 (O_148,N_14050,N_14140);
or UO_149 (O_149,N_14027,N_14608);
nand UO_150 (O_150,N_14242,N_14471);
xnor UO_151 (O_151,N_14622,N_14243);
nor UO_152 (O_152,N_14509,N_14837);
nor UO_153 (O_153,N_14752,N_14534);
and UO_154 (O_154,N_14090,N_14222);
or UO_155 (O_155,N_14401,N_14442);
and UO_156 (O_156,N_14460,N_14951);
or UO_157 (O_157,N_14900,N_14056);
nor UO_158 (O_158,N_14853,N_14331);
or UO_159 (O_159,N_14600,N_14943);
nor UO_160 (O_160,N_14370,N_14448);
or UO_161 (O_161,N_14217,N_14133);
and UO_162 (O_162,N_14876,N_14416);
nand UO_163 (O_163,N_14642,N_14013);
or UO_164 (O_164,N_14183,N_14640);
and UO_165 (O_165,N_14432,N_14645);
and UO_166 (O_166,N_14591,N_14746);
and UO_167 (O_167,N_14248,N_14739);
nor UO_168 (O_168,N_14934,N_14336);
nand UO_169 (O_169,N_14868,N_14990);
nor UO_170 (O_170,N_14779,N_14670);
or UO_171 (O_171,N_14241,N_14767);
and UO_172 (O_172,N_14319,N_14044);
or UO_173 (O_173,N_14165,N_14284);
or UO_174 (O_174,N_14884,N_14400);
nand UO_175 (O_175,N_14680,N_14451);
and UO_176 (O_176,N_14820,N_14548);
or UO_177 (O_177,N_14743,N_14313);
nand UO_178 (O_178,N_14096,N_14293);
nand UO_179 (O_179,N_14015,N_14066);
and UO_180 (O_180,N_14560,N_14649);
xnor UO_181 (O_181,N_14098,N_14235);
or UO_182 (O_182,N_14143,N_14993);
and UO_183 (O_183,N_14479,N_14216);
xnor UO_184 (O_184,N_14104,N_14792);
nor UO_185 (O_185,N_14508,N_14234);
nor UO_186 (O_186,N_14163,N_14974);
or UO_187 (O_187,N_14335,N_14524);
and UO_188 (O_188,N_14904,N_14441);
nor UO_189 (O_189,N_14315,N_14345);
nand UO_190 (O_190,N_14643,N_14397);
nand UO_191 (O_191,N_14340,N_14433);
nand UO_192 (O_192,N_14775,N_14688);
and UO_193 (O_193,N_14563,N_14129);
xor UO_194 (O_194,N_14351,N_14093);
or UO_195 (O_195,N_14523,N_14109);
nor UO_196 (O_196,N_14363,N_14396);
nor UO_197 (O_197,N_14839,N_14288);
or UO_198 (O_198,N_14295,N_14122);
nand UO_199 (O_199,N_14720,N_14323);
nor UO_200 (O_200,N_14488,N_14983);
and UO_201 (O_201,N_14603,N_14519);
and UO_202 (O_202,N_14421,N_14959);
or UO_203 (O_203,N_14383,N_14944);
and UO_204 (O_204,N_14758,N_14692);
and UO_205 (O_205,N_14701,N_14832);
or UO_206 (O_206,N_14034,N_14736);
or UO_207 (O_207,N_14979,N_14444);
and UO_208 (O_208,N_14167,N_14099);
or UO_209 (O_209,N_14415,N_14774);
or UO_210 (O_210,N_14039,N_14549);
and UO_211 (O_211,N_14579,N_14567);
nand UO_212 (O_212,N_14607,N_14817);
nor UO_213 (O_213,N_14806,N_14863);
nor UO_214 (O_214,N_14174,N_14762);
nor UO_215 (O_215,N_14976,N_14977);
or UO_216 (O_216,N_14819,N_14724);
nand UO_217 (O_217,N_14337,N_14995);
or UO_218 (O_218,N_14759,N_14963);
or UO_219 (O_219,N_14147,N_14008);
xor UO_220 (O_220,N_14434,N_14826);
and UO_221 (O_221,N_14290,N_14058);
xnor UO_222 (O_222,N_14483,N_14864);
xnor UO_223 (O_223,N_14891,N_14131);
or UO_224 (O_224,N_14660,N_14679);
nor UO_225 (O_225,N_14776,N_14360);
nand UO_226 (O_226,N_14343,N_14678);
or UO_227 (O_227,N_14468,N_14287);
nand UO_228 (O_228,N_14450,N_14081);
and UO_229 (O_229,N_14009,N_14957);
nand UO_230 (O_230,N_14173,N_14907);
nand UO_231 (O_231,N_14658,N_14474);
xor UO_232 (O_232,N_14593,N_14874);
nand UO_233 (O_233,N_14816,N_14386);
nor UO_234 (O_234,N_14624,N_14885);
xnor UO_235 (O_235,N_14283,N_14267);
or UO_236 (O_236,N_14916,N_14875);
or UO_237 (O_237,N_14896,N_14333);
nand UO_238 (O_238,N_14810,N_14598);
and UO_239 (O_239,N_14076,N_14512);
and UO_240 (O_240,N_14361,N_14048);
or UO_241 (O_241,N_14120,N_14516);
nor UO_242 (O_242,N_14804,N_14394);
xnor UO_243 (O_243,N_14953,N_14317);
and UO_244 (O_244,N_14738,N_14773);
and UO_245 (O_245,N_14641,N_14245);
or UO_246 (O_246,N_14466,N_14158);
nor UO_247 (O_247,N_14200,N_14978);
and UO_248 (O_248,N_14022,N_14691);
or UO_249 (O_249,N_14342,N_14589);
and UO_250 (O_250,N_14718,N_14229);
nor UO_251 (O_251,N_14456,N_14873);
and UO_252 (O_252,N_14505,N_14321);
or UO_253 (O_253,N_14862,N_14438);
nand UO_254 (O_254,N_14029,N_14311);
and UO_255 (O_255,N_14703,N_14757);
or UO_256 (O_256,N_14538,N_14655);
nand UO_257 (O_257,N_14552,N_14714);
nor UO_258 (O_258,N_14903,N_14697);
nor UO_259 (O_259,N_14797,N_14910);
nand UO_260 (O_260,N_14422,N_14683);
nand UO_261 (O_261,N_14064,N_14909);
nor UO_262 (O_262,N_14914,N_14710);
nand UO_263 (O_263,N_14439,N_14705);
nand UO_264 (O_264,N_14845,N_14393);
nor UO_265 (O_265,N_14310,N_14742);
or UO_266 (O_266,N_14796,N_14023);
or UO_267 (O_267,N_14072,N_14399);
and UO_268 (O_268,N_14318,N_14413);
nand UO_269 (O_269,N_14206,N_14429);
or UO_270 (O_270,N_14588,N_14427);
nand UO_271 (O_271,N_14121,N_14085);
or UO_272 (O_272,N_14919,N_14365);
nor UO_273 (O_273,N_14582,N_14205);
nand UO_274 (O_274,N_14423,N_14391);
or UO_275 (O_275,N_14584,N_14224);
nor UO_276 (O_276,N_14840,N_14431);
or UO_277 (O_277,N_14985,N_14219);
and UO_278 (O_278,N_14606,N_14926);
nor UO_279 (O_279,N_14123,N_14704);
nand UO_280 (O_280,N_14002,N_14305);
nor UO_281 (O_281,N_14677,N_14080);
xor UO_282 (O_282,N_14428,N_14601);
nor UO_283 (O_283,N_14307,N_14371);
or UO_284 (O_284,N_14051,N_14713);
nand UO_285 (O_285,N_14324,N_14376);
or UO_286 (O_286,N_14265,N_14367);
nand UO_287 (O_287,N_14971,N_14251);
nor UO_288 (O_288,N_14823,N_14156);
and UO_289 (O_289,N_14902,N_14160);
nor UO_290 (O_290,N_14948,N_14870);
and UO_291 (O_291,N_14626,N_14970);
and UO_292 (O_292,N_14017,N_14322);
nor UO_293 (O_293,N_14860,N_14550);
and UO_294 (O_294,N_14297,N_14294);
or UO_295 (O_295,N_14892,N_14915);
nand UO_296 (O_296,N_14228,N_14920);
and UO_297 (O_297,N_14529,N_14233);
and UO_298 (O_298,N_14530,N_14186);
nor UO_299 (O_299,N_14036,N_14753);
xor UO_300 (O_300,N_14170,N_14733);
or UO_301 (O_301,N_14153,N_14927);
nor UO_302 (O_302,N_14543,N_14952);
xor UO_303 (O_303,N_14955,N_14214);
or UO_304 (O_304,N_14610,N_14877);
and UO_305 (O_305,N_14040,N_14264);
nor UO_306 (O_306,N_14989,N_14793);
xor UO_307 (O_307,N_14225,N_14180);
or UO_308 (O_308,N_14230,N_14004);
and UO_309 (O_309,N_14646,N_14364);
or UO_310 (O_310,N_14671,N_14499);
and UO_311 (O_311,N_14652,N_14781);
xor UO_312 (O_312,N_14702,N_14181);
nand UO_313 (O_313,N_14866,N_14067);
and UO_314 (O_314,N_14802,N_14270);
nand UO_315 (O_315,N_14822,N_14330);
or UO_316 (O_316,N_14148,N_14623);
nor UO_317 (O_317,N_14256,N_14063);
and UO_318 (O_318,N_14633,N_14202);
or UO_319 (O_319,N_14079,N_14302);
nand UO_320 (O_320,N_14571,N_14184);
xor UO_321 (O_321,N_14341,N_14489);
or UO_322 (O_322,N_14732,N_14828);
nor UO_323 (O_323,N_14005,N_14278);
nand UO_324 (O_324,N_14159,N_14818);
or UO_325 (O_325,N_14246,N_14890);
and UO_326 (O_326,N_14966,N_14859);
nor UO_327 (O_327,N_14298,N_14846);
nor UO_328 (O_328,N_14813,N_14795);
and UO_329 (O_329,N_14836,N_14921);
and UO_330 (O_330,N_14491,N_14577);
nor UO_331 (O_331,N_14578,N_14301);
or UO_332 (O_332,N_14177,N_14790);
nand UO_333 (O_333,N_14204,N_14127);
or UO_334 (O_334,N_14038,N_14536);
nand UO_335 (O_335,N_14424,N_14878);
or UO_336 (O_336,N_14150,N_14968);
nand UO_337 (O_337,N_14358,N_14101);
nand UO_338 (O_338,N_14418,N_14855);
nand UO_339 (O_339,N_14001,N_14018);
nor UO_340 (O_340,N_14561,N_14010);
nor UO_341 (O_341,N_14355,N_14554);
and UO_342 (O_342,N_14994,N_14585);
or UO_343 (O_343,N_14597,N_14215);
and UO_344 (O_344,N_14674,N_14057);
nor UO_345 (O_345,N_14764,N_14357);
nor UO_346 (O_346,N_14869,N_14576);
or UO_347 (O_347,N_14440,N_14115);
or UO_348 (O_348,N_14069,N_14848);
nand UO_349 (O_349,N_14077,N_14566);
or UO_350 (O_350,N_14327,N_14484);
and UO_351 (O_351,N_14266,N_14794);
and UO_352 (O_352,N_14532,N_14043);
xor UO_353 (O_353,N_14356,N_14843);
and UO_354 (O_354,N_14162,N_14033);
nor UO_355 (O_355,N_14533,N_14666);
xnor UO_356 (O_356,N_14636,N_14786);
or UO_357 (O_357,N_14634,N_14882);
nand UO_358 (O_358,N_14087,N_14144);
xnor UO_359 (O_359,N_14880,N_14377);
nand UO_360 (O_360,N_14844,N_14602);
nor UO_361 (O_361,N_14325,N_14388);
and UO_362 (O_362,N_14016,N_14789);
nand UO_363 (O_363,N_14827,N_14706);
nand UO_364 (O_364,N_14469,N_14631);
nand UO_365 (O_365,N_14172,N_14203);
and UO_366 (O_366,N_14981,N_14961);
nand UO_367 (O_367,N_14700,N_14527);
and UO_368 (O_368,N_14374,N_14847);
nand UO_369 (O_369,N_14094,N_14540);
or UO_370 (O_370,N_14137,N_14715);
xnor UO_371 (O_371,N_14942,N_14865);
nor UO_372 (O_372,N_14766,N_14286);
nand UO_373 (O_373,N_14719,N_14741);
and UO_374 (O_374,N_14282,N_14729);
or UO_375 (O_375,N_14893,N_14731);
and UO_376 (O_376,N_14805,N_14630);
and UO_377 (O_377,N_14105,N_14014);
nand UO_378 (O_378,N_14667,N_14515);
or UO_379 (O_379,N_14854,N_14185);
xor UO_380 (O_380,N_14271,N_14788);
and UO_381 (O_381,N_14194,N_14100);
or UO_382 (O_382,N_14520,N_14130);
or UO_383 (O_383,N_14629,N_14821);
nor UO_384 (O_384,N_14208,N_14166);
nor UO_385 (O_385,N_14542,N_14409);
nand UO_386 (O_386,N_14492,N_14501);
nor UO_387 (O_387,N_14769,N_14521);
and UO_388 (O_388,N_14748,N_14136);
xnor UO_389 (O_389,N_14447,N_14569);
or UO_390 (O_390,N_14681,N_14984);
and UO_391 (O_391,N_14047,N_14308);
or UO_392 (O_392,N_14430,N_14473);
nand UO_393 (O_393,N_14258,N_14751);
nand UO_394 (O_394,N_14236,N_14611);
and UO_395 (O_395,N_14518,N_14693);
nand UO_396 (O_396,N_14021,N_14124);
or UO_397 (O_397,N_14825,N_14149);
nand UO_398 (O_398,N_14572,N_14249);
or UO_399 (O_399,N_14980,N_14612);
and UO_400 (O_400,N_14037,N_14722);
and UO_401 (O_401,N_14176,N_14420);
and UO_402 (O_402,N_14443,N_14975);
nor UO_403 (O_403,N_14352,N_14328);
xor UO_404 (O_404,N_14879,N_14378);
nor UO_405 (O_405,N_14553,N_14020);
xor UO_406 (O_406,N_14761,N_14373);
nand UO_407 (O_407,N_14019,N_14353);
and UO_408 (O_408,N_14936,N_14285);
nor UO_409 (O_409,N_14778,N_14947);
nor UO_410 (O_410,N_14908,N_14676);
nand UO_411 (O_411,N_14556,N_14834);
nand UO_412 (O_412,N_14102,N_14175);
or UO_413 (O_413,N_14850,N_14279);
or UO_414 (O_414,N_14768,N_14949);
and UO_415 (O_415,N_14972,N_14931);
nor UO_416 (O_416,N_14296,N_14545);
or UO_417 (O_417,N_14514,N_14281);
and UO_418 (O_418,N_14062,N_14119);
and UO_419 (O_419,N_14253,N_14083);
or UO_420 (O_420,N_14312,N_14380);
and UO_421 (O_421,N_14675,N_14338);
nand UO_422 (O_422,N_14756,N_14407);
xor UO_423 (O_423,N_14329,N_14049);
nand UO_424 (O_424,N_14898,N_14261);
or UO_425 (O_425,N_14638,N_14237);
nand UO_426 (O_426,N_14881,N_14925);
or UO_427 (O_427,N_14618,N_14664);
xnor UO_428 (O_428,N_14000,N_14461);
and UO_429 (O_429,N_14871,N_14389);
and UO_430 (O_430,N_14070,N_14932);
nor UO_431 (O_431,N_14734,N_14381);
or UO_432 (O_432,N_14375,N_14035);
nand UO_433 (O_433,N_14385,N_14486);
or UO_434 (O_434,N_14189,N_14103);
nor UO_435 (O_435,N_14580,N_14535);
nand UO_436 (O_436,N_14350,N_14614);
or UO_437 (O_437,N_14780,N_14728);
or UO_438 (O_438,N_14929,N_14872);
or UO_439 (O_439,N_14887,N_14662);
nand UO_440 (O_440,N_14179,N_14982);
or UO_441 (O_441,N_14842,N_14808);
nor UO_442 (O_442,N_14564,N_14272);
and UO_443 (O_443,N_14760,N_14851);
xor UO_444 (O_444,N_14463,N_14411);
nand UO_445 (O_445,N_14213,N_14906);
nor UO_446 (O_446,N_14537,N_14073);
and UO_447 (O_447,N_14928,N_14395);
or UO_448 (O_448,N_14011,N_14506);
nand UO_449 (O_449,N_14339,N_14727);
xor UO_450 (O_450,N_14089,N_14012);
or UO_451 (O_451,N_14197,N_14895);
and UO_452 (O_452,N_14747,N_14587);
xor UO_453 (O_453,N_14917,N_14682);
or UO_454 (O_454,N_14901,N_14436);
and UO_455 (O_455,N_14659,N_14945);
nand UO_456 (O_456,N_14250,N_14007);
or UO_457 (O_457,N_14883,N_14650);
or UO_458 (O_458,N_14059,N_14657);
and UO_459 (O_459,N_14053,N_14118);
and UO_460 (O_460,N_14097,N_14604);
and UO_461 (O_461,N_14126,N_14559);
xnor UO_462 (O_462,N_14551,N_14480);
and UO_463 (O_463,N_14108,N_14490);
or UO_464 (O_464,N_14362,N_14262);
or UO_465 (O_465,N_14074,N_14274);
and UO_466 (O_466,N_14861,N_14801);
xor UO_467 (O_467,N_14494,N_14510);
or UO_468 (O_468,N_14784,N_14273);
or UO_469 (O_469,N_14574,N_14737);
or UO_470 (O_470,N_14187,N_14815);
and UO_471 (O_471,N_14594,N_14555);
nand UO_472 (O_472,N_14419,N_14507);
nor UO_473 (O_473,N_14924,N_14276);
and UO_474 (O_474,N_14814,N_14867);
and UO_475 (O_475,N_14061,N_14151);
nand UO_476 (O_476,N_14656,N_14617);
nor UO_477 (O_477,N_14745,N_14504);
and UO_478 (O_478,N_14956,N_14134);
or UO_479 (O_479,N_14496,N_14320);
or UO_480 (O_480,N_14522,N_14210);
or UO_481 (O_481,N_14672,N_14464);
nand UO_482 (O_482,N_14304,N_14546);
nor UO_483 (O_483,N_14635,N_14783);
nor UO_484 (O_484,N_14829,N_14668);
nor UO_485 (O_485,N_14613,N_14142);
or UO_486 (O_486,N_14899,N_14227);
or UO_487 (O_487,N_14032,N_14292);
or UO_488 (O_488,N_14209,N_14349);
nor UO_489 (O_489,N_14195,N_14628);
and UO_490 (O_490,N_14382,N_14986);
nand UO_491 (O_491,N_14193,N_14946);
nor UO_492 (O_492,N_14857,N_14935);
and UO_493 (O_493,N_14997,N_14398);
nor UO_494 (O_494,N_14088,N_14940);
and UO_495 (O_495,N_14687,N_14065);
nand UO_496 (O_496,N_14112,N_14723);
nand UO_497 (O_497,N_14417,N_14218);
nand UO_498 (O_498,N_14487,N_14390);
nand UO_499 (O_499,N_14621,N_14833);
nand UO_500 (O_500,N_14421,N_14703);
nor UO_501 (O_501,N_14554,N_14512);
or UO_502 (O_502,N_14292,N_14048);
and UO_503 (O_503,N_14181,N_14771);
or UO_504 (O_504,N_14158,N_14785);
or UO_505 (O_505,N_14947,N_14883);
nor UO_506 (O_506,N_14506,N_14368);
nand UO_507 (O_507,N_14226,N_14998);
or UO_508 (O_508,N_14521,N_14709);
or UO_509 (O_509,N_14181,N_14584);
and UO_510 (O_510,N_14955,N_14628);
nor UO_511 (O_511,N_14127,N_14736);
xor UO_512 (O_512,N_14087,N_14743);
xnor UO_513 (O_513,N_14655,N_14316);
nand UO_514 (O_514,N_14302,N_14471);
and UO_515 (O_515,N_14976,N_14569);
nor UO_516 (O_516,N_14604,N_14300);
nand UO_517 (O_517,N_14622,N_14483);
or UO_518 (O_518,N_14773,N_14741);
or UO_519 (O_519,N_14328,N_14150);
or UO_520 (O_520,N_14016,N_14911);
and UO_521 (O_521,N_14985,N_14478);
or UO_522 (O_522,N_14456,N_14883);
and UO_523 (O_523,N_14488,N_14570);
nor UO_524 (O_524,N_14103,N_14517);
or UO_525 (O_525,N_14498,N_14423);
xnor UO_526 (O_526,N_14649,N_14030);
and UO_527 (O_527,N_14823,N_14293);
nor UO_528 (O_528,N_14626,N_14913);
xor UO_529 (O_529,N_14091,N_14619);
or UO_530 (O_530,N_14469,N_14421);
and UO_531 (O_531,N_14447,N_14385);
nand UO_532 (O_532,N_14009,N_14870);
nor UO_533 (O_533,N_14764,N_14209);
or UO_534 (O_534,N_14634,N_14737);
and UO_535 (O_535,N_14641,N_14769);
nand UO_536 (O_536,N_14262,N_14626);
or UO_537 (O_537,N_14506,N_14742);
and UO_538 (O_538,N_14649,N_14555);
nor UO_539 (O_539,N_14195,N_14435);
nand UO_540 (O_540,N_14319,N_14495);
nand UO_541 (O_541,N_14004,N_14423);
nand UO_542 (O_542,N_14843,N_14641);
nor UO_543 (O_543,N_14360,N_14089);
or UO_544 (O_544,N_14973,N_14533);
or UO_545 (O_545,N_14155,N_14045);
or UO_546 (O_546,N_14133,N_14474);
nand UO_547 (O_547,N_14156,N_14738);
nand UO_548 (O_548,N_14609,N_14852);
or UO_549 (O_549,N_14032,N_14481);
nand UO_550 (O_550,N_14925,N_14084);
nor UO_551 (O_551,N_14449,N_14902);
and UO_552 (O_552,N_14344,N_14292);
nand UO_553 (O_553,N_14313,N_14853);
nand UO_554 (O_554,N_14210,N_14053);
xor UO_555 (O_555,N_14075,N_14215);
and UO_556 (O_556,N_14569,N_14729);
or UO_557 (O_557,N_14448,N_14127);
nand UO_558 (O_558,N_14382,N_14169);
nor UO_559 (O_559,N_14401,N_14713);
nor UO_560 (O_560,N_14908,N_14409);
and UO_561 (O_561,N_14739,N_14303);
or UO_562 (O_562,N_14290,N_14509);
and UO_563 (O_563,N_14157,N_14591);
nand UO_564 (O_564,N_14366,N_14936);
and UO_565 (O_565,N_14925,N_14330);
nand UO_566 (O_566,N_14707,N_14251);
nor UO_567 (O_567,N_14865,N_14530);
or UO_568 (O_568,N_14376,N_14397);
nor UO_569 (O_569,N_14558,N_14397);
nor UO_570 (O_570,N_14038,N_14994);
nand UO_571 (O_571,N_14051,N_14919);
nand UO_572 (O_572,N_14413,N_14095);
nor UO_573 (O_573,N_14772,N_14032);
nand UO_574 (O_574,N_14629,N_14208);
xor UO_575 (O_575,N_14283,N_14228);
nand UO_576 (O_576,N_14975,N_14452);
and UO_577 (O_577,N_14090,N_14770);
nand UO_578 (O_578,N_14743,N_14074);
xnor UO_579 (O_579,N_14226,N_14649);
xnor UO_580 (O_580,N_14471,N_14809);
and UO_581 (O_581,N_14147,N_14935);
nand UO_582 (O_582,N_14742,N_14810);
and UO_583 (O_583,N_14354,N_14597);
nor UO_584 (O_584,N_14001,N_14014);
nand UO_585 (O_585,N_14258,N_14245);
and UO_586 (O_586,N_14144,N_14573);
nor UO_587 (O_587,N_14865,N_14042);
nor UO_588 (O_588,N_14174,N_14192);
or UO_589 (O_589,N_14455,N_14830);
nor UO_590 (O_590,N_14696,N_14414);
and UO_591 (O_591,N_14812,N_14477);
and UO_592 (O_592,N_14634,N_14492);
or UO_593 (O_593,N_14008,N_14272);
or UO_594 (O_594,N_14373,N_14776);
xor UO_595 (O_595,N_14685,N_14858);
nor UO_596 (O_596,N_14314,N_14250);
nand UO_597 (O_597,N_14293,N_14387);
nand UO_598 (O_598,N_14846,N_14977);
and UO_599 (O_599,N_14803,N_14744);
nand UO_600 (O_600,N_14347,N_14548);
or UO_601 (O_601,N_14453,N_14818);
or UO_602 (O_602,N_14660,N_14058);
nand UO_603 (O_603,N_14143,N_14645);
xor UO_604 (O_604,N_14795,N_14938);
or UO_605 (O_605,N_14371,N_14508);
or UO_606 (O_606,N_14533,N_14488);
or UO_607 (O_607,N_14983,N_14329);
and UO_608 (O_608,N_14044,N_14212);
nand UO_609 (O_609,N_14690,N_14089);
nor UO_610 (O_610,N_14017,N_14871);
nand UO_611 (O_611,N_14493,N_14521);
or UO_612 (O_612,N_14899,N_14231);
xnor UO_613 (O_613,N_14485,N_14280);
or UO_614 (O_614,N_14664,N_14904);
nor UO_615 (O_615,N_14711,N_14831);
nand UO_616 (O_616,N_14063,N_14156);
xor UO_617 (O_617,N_14265,N_14198);
and UO_618 (O_618,N_14516,N_14599);
nor UO_619 (O_619,N_14229,N_14654);
or UO_620 (O_620,N_14141,N_14452);
nor UO_621 (O_621,N_14268,N_14037);
or UO_622 (O_622,N_14713,N_14953);
and UO_623 (O_623,N_14511,N_14966);
or UO_624 (O_624,N_14913,N_14560);
or UO_625 (O_625,N_14439,N_14236);
nor UO_626 (O_626,N_14832,N_14970);
or UO_627 (O_627,N_14928,N_14892);
nor UO_628 (O_628,N_14563,N_14821);
or UO_629 (O_629,N_14052,N_14854);
or UO_630 (O_630,N_14597,N_14741);
and UO_631 (O_631,N_14948,N_14105);
or UO_632 (O_632,N_14216,N_14251);
nor UO_633 (O_633,N_14194,N_14483);
or UO_634 (O_634,N_14092,N_14039);
nor UO_635 (O_635,N_14361,N_14493);
nand UO_636 (O_636,N_14504,N_14832);
and UO_637 (O_637,N_14673,N_14882);
nor UO_638 (O_638,N_14528,N_14232);
nand UO_639 (O_639,N_14753,N_14001);
xnor UO_640 (O_640,N_14355,N_14445);
nor UO_641 (O_641,N_14392,N_14991);
nand UO_642 (O_642,N_14919,N_14665);
or UO_643 (O_643,N_14365,N_14736);
or UO_644 (O_644,N_14414,N_14292);
and UO_645 (O_645,N_14472,N_14391);
and UO_646 (O_646,N_14453,N_14809);
and UO_647 (O_647,N_14160,N_14715);
xnor UO_648 (O_648,N_14555,N_14120);
and UO_649 (O_649,N_14294,N_14986);
nand UO_650 (O_650,N_14019,N_14436);
nor UO_651 (O_651,N_14521,N_14931);
or UO_652 (O_652,N_14863,N_14226);
and UO_653 (O_653,N_14329,N_14913);
or UO_654 (O_654,N_14710,N_14301);
nand UO_655 (O_655,N_14606,N_14564);
nor UO_656 (O_656,N_14028,N_14365);
or UO_657 (O_657,N_14834,N_14741);
nand UO_658 (O_658,N_14236,N_14741);
nor UO_659 (O_659,N_14061,N_14199);
nor UO_660 (O_660,N_14976,N_14216);
nor UO_661 (O_661,N_14986,N_14009);
and UO_662 (O_662,N_14299,N_14221);
nand UO_663 (O_663,N_14988,N_14225);
nand UO_664 (O_664,N_14933,N_14485);
nand UO_665 (O_665,N_14142,N_14140);
or UO_666 (O_666,N_14036,N_14478);
nor UO_667 (O_667,N_14710,N_14666);
or UO_668 (O_668,N_14679,N_14780);
nand UO_669 (O_669,N_14125,N_14485);
nor UO_670 (O_670,N_14188,N_14139);
and UO_671 (O_671,N_14952,N_14550);
and UO_672 (O_672,N_14704,N_14478);
or UO_673 (O_673,N_14655,N_14143);
xnor UO_674 (O_674,N_14426,N_14560);
or UO_675 (O_675,N_14238,N_14956);
nand UO_676 (O_676,N_14390,N_14502);
or UO_677 (O_677,N_14556,N_14331);
and UO_678 (O_678,N_14716,N_14252);
xor UO_679 (O_679,N_14952,N_14937);
nor UO_680 (O_680,N_14666,N_14874);
nand UO_681 (O_681,N_14974,N_14726);
xor UO_682 (O_682,N_14912,N_14748);
and UO_683 (O_683,N_14378,N_14566);
xnor UO_684 (O_684,N_14436,N_14508);
xor UO_685 (O_685,N_14880,N_14226);
nor UO_686 (O_686,N_14197,N_14835);
and UO_687 (O_687,N_14310,N_14210);
and UO_688 (O_688,N_14713,N_14995);
or UO_689 (O_689,N_14145,N_14530);
xor UO_690 (O_690,N_14906,N_14310);
xor UO_691 (O_691,N_14234,N_14247);
xor UO_692 (O_692,N_14897,N_14959);
and UO_693 (O_693,N_14973,N_14965);
and UO_694 (O_694,N_14373,N_14588);
xnor UO_695 (O_695,N_14668,N_14806);
xor UO_696 (O_696,N_14863,N_14836);
nor UO_697 (O_697,N_14185,N_14996);
nand UO_698 (O_698,N_14509,N_14985);
or UO_699 (O_699,N_14988,N_14507);
and UO_700 (O_700,N_14406,N_14396);
and UO_701 (O_701,N_14326,N_14632);
xor UO_702 (O_702,N_14145,N_14142);
xnor UO_703 (O_703,N_14676,N_14448);
and UO_704 (O_704,N_14025,N_14176);
nand UO_705 (O_705,N_14613,N_14636);
nor UO_706 (O_706,N_14820,N_14008);
xor UO_707 (O_707,N_14631,N_14194);
and UO_708 (O_708,N_14232,N_14198);
nor UO_709 (O_709,N_14803,N_14682);
and UO_710 (O_710,N_14286,N_14550);
nor UO_711 (O_711,N_14497,N_14616);
or UO_712 (O_712,N_14379,N_14876);
nor UO_713 (O_713,N_14753,N_14649);
nor UO_714 (O_714,N_14015,N_14596);
or UO_715 (O_715,N_14862,N_14780);
xor UO_716 (O_716,N_14604,N_14277);
nand UO_717 (O_717,N_14388,N_14166);
or UO_718 (O_718,N_14452,N_14714);
or UO_719 (O_719,N_14462,N_14943);
nor UO_720 (O_720,N_14781,N_14827);
and UO_721 (O_721,N_14822,N_14602);
nor UO_722 (O_722,N_14556,N_14046);
and UO_723 (O_723,N_14328,N_14148);
nor UO_724 (O_724,N_14248,N_14196);
nor UO_725 (O_725,N_14538,N_14281);
and UO_726 (O_726,N_14774,N_14500);
and UO_727 (O_727,N_14482,N_14158);
xnor UO_728 (O_728,N_14532,N_14045);
or UO_729 (O_729,N_14129,N_14460);
and UO_730 (O_730,N_14911,N_14235);
nor UO_731 (O_731,N_14568,N_14912);
nor UO_732 (O_732,N_14618,N_14394);
xnor UO_733 (O_733,N_14517,N_14238);
nand UO_734 (O_734,N_14492,N_14620);
and UO_735 (O_735,N_14102,N_14568);
or UO_736 (O_736,N_14103,N_14042);
and UO_737 (O_737,N_14530,N_14458);
nand UO_738 (O_738,N_14398,N_14465);
and UO_739 (O_739,N_14386,N_14825);
nor UO_740 (O_740,N_14030,N_14337);
nor UO_741 (O_741,N_14707,N_14838);
and UO_742 (O_742,N_14371,N_14735);
and UO_743 (O_743,N_14126,N_14256);
and UO_744 (O_744,N_14201,N_14037);
or UO_745 (O_745,N_14035,N_14602);
nand UO_746 (O_746,N_14321,N_14779);
or UO_747 (O_747,N_14616,N_14713);
or UO_748 (O_748,N_14049,N_14145);
or UO_749 (O_749,N_14739,N_14990);
and UO_750 (O_750,N_14569,N_14662);
and UO_751 (O_751,N_14186,N_14238);
and UO_752 (O_752,N_14054,N_14849);
nand UO_753 (O_753,N_14433,N_14704);
or UO_754 (O_754,N_14685,N_14798);
nor UO_755 (O_755,N_14599,N_14963);
or UO_756 (O_756,N_14590,N_14346);
nand UO_757 (O_757,N_14636,N_14911);
and UO_758 (O_758,N_14120,N_14735);
or UO_759 (O_759,N_14168,N_14431);
or UO_760 (O_760,N_14211,N_14441);
nand UO_761 (O_761,N_14787,N_14658);
nor UO_762 (O_762,N_14931,N_14031);
nand UO_763 (O_763,N_14574,N_14988);
nand UO_764 (O_764,N_14480,N_14921);
xnor UO_765 (O_765,N_14192,N_14124);
nand UO_766 (O_766,N_14538,N_14935);
nor UO_767 (O_767,N_14088,N_14738);
nor UO_768 (O_768,N_14243,N_14835);
or UO_769 (O_769,N_14608,N_14612);
nor UO_770 (O_770,N_14305,N_14677);
nor UO_771 (O_771,N_14766,N_14077);
and UO_772 (O_772,N_14636,N_14900);
or UO_773 (O_773,N_14732,N_14226);
or UO_774 (O_774,N_14778,N_14597);
or UO_775 (O_775,N_14408,N_14912);
nor UO_776 (O_776,N_14641,N_14724);
or UO_777 (O_777,N_14815,N_14009);
nand UO_778 (O_778,N_14522,N_14390);
nand UO_779 (O_779,N_14351,N_14390);
or UO_780 (O_780,N_14819,N_14562);
or UO_781 (O_781,N_14121,N_14633);
xnor UO_782 (O_782,N_14036,N_14333);
nor UO_783 (O_783,N_14960,N_14140);
nor UO_784 (O_784,N_14171,N_14019);
nand UO_785 (O_785,N_14118,N_14863);
nand UO_786 (O_786,N_14395,N_14164);
nand UO_787 (O_787,N_14422,N_14530);
or UO_788 (O_788,N_14486,N_14304);
and UO_789 (O_789,N_14845,N_14983);
nor UO_790 (O_790,N_14138,N_14234);
and UO_791 (O_791,N_14308,N_14925);
nor UO_792 (O_792,N_14525,N_14750);
xor UO_793 (O_793,N_14373,N_14236);
or UO_794 (O_794,N_14817,N_14645);
and UO_795 (O_795,N_14833,N_14894);
and UO_796 (O_796,N_14023,N_14210);
nand UO_797 (O_797,N_14133,N_14846);
nor UO_798 (O_798,N_14911,N_14132);
nand UO_799 (O_799,N_14419,N_14787);
nand UO_800 (O_800,N_14566,N_14895);
or UO_801 (O_801,N_14097,N_14341);
nor UO_802 (O_802,N_14840,N_14876);
nor UO_803 (O_803,N_14064,N_14800);
or UO_804 (O_804,N_14008,N_14808);
and UO_805 (O_805,N_14016,N_14439);
and UO_806 (O_806,N_14836,N_14057);
xor UO_807 (O_807,N_14283,N_14435);
nand UO_808 (O_808,N_14912,N_14233);
nor UO_809 (O_809,N_14485,N_14591);
and UO_810 (O_810,N_14008,N_14266);
nor UO_811 (O_811,N_14638,N_14975);
or UO_812 (O_812,N_14530,N_14945);
and UO_813 (O_813,N_14367,N_14622);
nor UO_814 (O_814,N_14114,N_14169);
nor UO_815 (O_815,N_14774,N_14297);
xnor UO_816 (O_816,N_14542,N_14443);
or UO_817 (O_817,N_14385,N_14602);
nand UO_818 (O_818,N_14854,N_14728);
nor UO_819 (O_819,N_14359,N_14513);
nor UO_820 (O_820,N_14419,N_14260);
nand UO_821 (O_821,N_14570,N_14522);
or UO_822 (O_822,N_14081,N_14456);
nand UO_823 (O_823,N_14885,N_14620);
and UO_824 (O_824,N_14594,N_14476);
or UO_825 (O_825,N_14768,N_14194);
and UO_826 (O_826,N_14856,N_14537);
nor UO_827 (O_827,N_14678,N_14619);
nor UO_828 (O_828,N_14297,N_14554);
or UO_829 (O_829,N_14307,N_14107);
and UO_830 (O_830,N_14774,N_14521);
nand UO_831 (O_831,N_14138,N_14631);
nand UO_832 (O_832,N_14463,N_14912);
or UO_833 (O_833,N_14159,N_14960);
or UO_834 (O_834,N_14146,N_14467);
nor UO_835 (O_835,N_14148,N_14850);
nor UO_836 (O_836,N_14759,N_14571);
xor UO_837 (O_837,N_14768,N_14502);
nand UO_838 (O_838,N_14137,N_14127);
and UO_839 (O_839,N_14767,N_14193);
nor UO_840 (O_840,N_14954,N_14044);
nor UO_841 (O_841,N_14933,N_14777);
or UO_842 (O_842,N_14725,N_14492);
or UO_843 (O_843,N_14774,N_14729);
xor UO_844 (O_844,N_14484,N_14824);
nor UO_845 (O_845,N_14831,N_14301);
nor UO_846 (O_846,N_14447,N_14522);
nor UO_847 (O_847,N_14273,N_14971);
and UO_848 (O_848,N_14352,N_14381);
or UO_849 (O_849,N_14470,N_14066);
nor UO_850 (O_850,N_14511,N_14872);
and UO_851 (O_851,N_14056,N_14129);
and UO_852 (O_852,N_14047,N_14776);
nand UO_853 (O_853,N_14026,N_14544);
and UO_854 (O_854,N_14974,N_14851);
nand UO_855 (O_855,N_14412,N_14868);
nor UO_856 (O_856,N_14385,N_14079);
and UO_857 (O_857,N_14706,N_14329);
xnor UO_858 (O_858,N_14189,N_14104);
or UO_859 (O_859,N_14964,N_14971);
nor UO_860 (O_860,N_14249,N_14055);
nor UO_861 (O_861,N_14115,N_14648);
and UO_862 (O_862,N_14117,N_14290);
nand UO_863 (O_863,N_14787,N_14037);
nand UO_864 (O_864,N_14023,N_14911);
or UO_865 (O_865,N_14114,N_14787);
nor UO_866 (O_866,N_14541,N_14183);
nor UO_867 (O_867,N_14007,N_14427);
nor UO_868 (O_868,N_14509,N_14029);
nand UO_869 (O_869,N_14395,N_14384);
nand UO_870 (O_870,N_14350,N_14812);
and UO_871 (O_871,N_14383,N_14332);
nor UO_872 (O_872,N_14739,N_14600);
nor UO_873 (O_873,N_14157,N_14898);
nand UO_874 (O_874,N_14994,N_14643);
nor UO_875 (O_875,N_14142,N_14847);
nand UO_876 (O_876,N_14271,N_14658);
xor UO_877 (O_877,N_14254,N_14201);
nor UO_878 (O_878,N_14435,N_14093);
nor UO_879 (O_879,N_14874,N_14683);
or UO_880 (O_880,N_14195,N_14550);
and UO_881 (O_881,N_14732,N_14444);
and UO_882 (O_882,N_14468,N_14120);
and UO_883 (O_883,N_14555,N_14414);
or UO_884 (O_884,N_14455,N_14332);
or UO_885 (O_885,N_14941,N_14363);
nand UO_886 (O_886,N_14521,N_14857);
and UO_887 (O_887,N_14868,N_14484);
nand UO_888 (O_888,N_14635,N_14732);
or UO_889 (O_889,N_14763,N_14296);
and UO_890 (O_890,N_14842,N_14229);
nand UO_891 (O_891,N_14199,N_14619);
nor UO_892 (O_892,N_14768,N_14818);
xor UO_893 (O_893,N_14515,N_14303);
and UO_894 (O_894,N_14169,N_14049);
and UO_895 (O_895,N_14145,N_14615);
and UO_896 (O_896,N_14718,N_14748);
xor UO_897 (O_897,N_14987,N_14310);
and UO_898 (O_898,N_14412,N_14840);
or UO_899 (O_899,N_14839,N_14763);
nand UO_900 (O_900,N_14684,N_14578);
or UO_901 (O_901,N_14290,N_14628);
or UO_902 (O_902,N_14972,N_14779);
or UO_903 (O_903,N_14843,N_14287);
nor UO_904 (O_904,N_14171,N_14044);
and UO_905 (O_905,N_14270,N_14168);
and UO_906 (O_906,N_14040,N_14204);
and UO_907 (O_907,N_14241,N_14355);
and UO_908 (O_908,N_14535,N_14443);
nor UO_909 (O_909,N_14105,N_14371);
xnor UO_910 (O_910,N_14790,N_14842);
nand UO_911 (O_911,N_14569,N_14879);
nor UO_912 (O_912,N_14931,N_14207);
or UO_913 (O_913,N_14860,N_14309);
xor UO_914 (O_914,N_14384,N_14294);
or UO_915 (O_915,N_14715,N_14503);
nand UO_916 (O_916,N_14921,N_14318);
nor UO_917 (O_917,N_14226,N_14949);
and UO_918 (O_918,N_14035,N_14689);
nand UO_919 (O_919,N_14277,N_14383);
or UO_920 (O_920,N_14398,N_14339);
xor UO_921 (O_921,N_14322,N_14833);
and UO_922 (O_922,N_14275,N_14227);
or UO_923 (O_923,N_14951,N_14445);
xnor UO_924 (O_924,N_14053,N_14980);
nand UO_925 (O_925,N_14641,N_14548);
and UO_926 (O_926,N_14533,N_14597);
and UO_927 (O_927,N_14637,N_14398);
nor UO_928 (O_928,N_14422,N_14176);
or UO_929 (O_929,N_14629,N_14519);
and UO_930 (O_930,N_14221,N_14962);
or UO_931 (O_931,N_14195,N_14173);
and UO_932 (O_932,N_14314,N_14034);
nor UO_933 (O_933,N_14476,N_14458);
nand UO_934 (O_934,N_14760,N_14216);
nor UO_935 (O_935,N_14019,N_14696);
nor UO_936 (O_936,N_14248,N_14275);
or UO_937 (O_937,N_14288,N_14633);
or UO_938 (O_938,N_14494,N_14483);
xor UO_939 (O_939,N_14379,N_14008);
nor UO_940 (O_940,N_14385,N_14330);
and UO_941 (O_941,N_14491,N_14319);
and UO_942 (O_942,N_14552,N_14290);
nand UO_943 (O_943,N_14207,N_14357);
xor UO_944 (O_944,N_14908,N_14533);
nor UO_945 (O_945,N_14033,N_14361);
or UO_946 (O_946,N_14568,N_14223);
and UO_947 (O_947,N_14532,N_14802);
xnor UO_948 (O_948,N_14905,N_14282);
and UO_949 (O_949,N_14162,N_14789);
xnor UO_950 (O_950,N_14594,N_14883);
or UO_951 (O_951,N_14527,N_14814);
or UO_952 (O_952,N_14628,N_14522);
nand UO_953 (O_953,N_14946,N_14690);
or UO_954 (O_954,N_14771,N_14515);
or UO_955 (O_955,N_14216,N_14905);
nand UO_956 (O_956,N_14140,N_14882);
and UO_957 (O_957,N_14092,N_14499);
and UO_958 (O_958,N_14387,N_14231);
or UO_959 (O_959,N_14256,N_14030);
nor UO_960 (O_960,N_14910,N_14912);
nand UO_961 (O_961,N_14985,N_14170);
nand UO_962 (O_962,N_14015,N_14036);
nor UO_963 (O_963,N_14046,N_14609);
xnor UO_964 (O_964,N_14554,N_14123);
xor UO_965 (O_965,N_14359,N_14817);
and UO_966 (O_966,N_14779,N_14667);
xor UO_967 (O_967,N_14436,N_14481);
or UO_968 (O_968,N_14442,N_14810);
and UO_969 (O_969,N_14767,N_14300);
and UO_970 (O_970,N_14866,N_14700);
nor UO_971 (O_971,N_14142,N_14766);
and UO_972 (O_972,N_14328,N_14973);
and UO_973 (O_973,N_14420,N_14748);
nand UO_974 (O_974,N_14444,N_14798);
xor UO_975 (O_975,N_14789,N_14784);
nor UO_976 (O_976,N_14595,N_14351);
nor UO_977 (O_977,N_14014,N_14046);
or UO_978 (O_978,N_14867,N_14810);
or UO_979 (O_979,N_14860,N_14253);
xnor UO_980 (O_980,N_14887,N_14810);
nor UO_981 (O_981,N_14704,N_14703);
and UO_982 (O_982,N_14921,N_14346);
nand UO_983 (O_983,N_14029,N_14506);
or UO_984 (O_984,N_14703,N_14958);
and UO_985 (O_985,N_14310,N_14832);
or UO_986 (O_986,N_14932,N_14714);
nand UO_987 (O_987,N_14210,N_14117);
xnor UO_988 (O_988,N_14737,N_14975);
nor UO_989 (O_989,N_14167,N_14249);
nand UO_990 (O_990,N_14471,N_14392);
or UO_991 (O_991,N_14552,N_14113);
nand UO_992 (O_992,N_14683,N_14951);
xor UO_993 (O_993,N_14043,N_14992);
and UO_994 (O_994,N_14524,N_14879);
nand UO_995 (O_995,N_14957,N_14970);
or UO_996 (O_996,N_14764,N_14417);
nand UO_997 (O_997,N_14212,N_14066);
nor UO_998 (O_998,N_14725,N_14998);
and UO_999 (O_999,N_14903,N_14382);
or UO_1000 (O_1000,N_14018,N_14273);
xor UO_1001 (O_1001,N_14409,N_14208);
nor UO_1002 (O_1002,N_14008,N_14998);
or UO_1003 (O_1003,N_14289,N_14180);
nor UO_1004 (O_1004,N_14664,N_14062);
nand UO_1005 (O_1005,N_14635,N_14139);
and UO_1006 (O_1006,N_14197,N_14412);
xor UO_1007 (O_1007,N_14909,N_14490);
or UO_1008 (O_1008,N_14206,N_14289);
or UO_1009 (O_1009,N_14706,N_14434);
nor UO_1010 (O_1010,N_14012,N_14351);
or UO_1011 (O_1011,N_14224,N_14420);
nand UO_1012 (O_1012,N_14981,N_14424);
nand UO_1013 (O_1013,N_14547,N_14330);
and UO_1014 (O_1014,N_14661,N_14008);
nand UO_1015 (O_1015,N_14937,N_14124);
and UO_1016 (O_1016,N_14735,N_14124);
nor UO_1017 (O_1017,N_14703,N_14750);
or UO_1018 (O_1018,N_14198,N_14803);
or UO_1019 (O_1019,N_14570,N_14365);
xor UO_1020 (O_1020,N_14240,N_14950);
nor UO_1021 (O_1021,N_14939,N_14229);
or UO_1022 (O_1022,N_14036,N_14778);
xnor UO_1023 (O_1023,N_14678,N_14928);
xnor UO_1024 (O_1024,N_14197,N_14619);
xor UO_1025 (O_1025,N_14213,N_14160);
xor UO_1026 (O_1026,N_14194,N_14777);
or UO_1027 (O_1027,N_14936,N_14202);
or UO_1028 (O_1028,N_14217,N_14286);
nor UO_1029 (O_1029,N_14037,N_14497);
nand UO_1030 (O_1030,N_14179,N_14065);
nor UO_1031 (O_1031,N_14595,N_14213);
or UO_1032 (O_1032,N_14444,N_14559);
and UO_1033 (O_1033,N_14209,N_14751);
nand UO_1034 (O_1034,N_14418,N_14948);
or UO_1035 (O_1035,N_14720,N_14161);
nand UO_1036 (O_1036,N_14122,N_14526);
or UO_1037 (O_1037,N_14852,N_14274);
nand UO_1038 (O_1038,N_14135,N_14502);
nand UO_1039 (O_1039,N_14304,N_14858);
and UO_1040 (O_1040,N_14626,N_14621);
and UO_1041 (O_1041,N_14210,N_14765);
and UO_1042 (O_1042,N_14410,N_14783);
nand UO_1043 (O_1043,N_14356,N_14309);
or UO_1044 (O_1044,N_14235,N_14191);
nand UO_1045 (O_1045,N_14658,N_14996);
nand UO_1046 (O_1046,N_14879,N_14964);
and UO_1047 (O_1047,N_14431,N_14201);
nand UO_1048 (O_1048,N_14634,N_14322);
nand UO_1049 (O_1049,N_14785,N_14826);
and UO_1050 (O_1050,N_14387,N_14295);
and UO_1051 (O_1051,N_14166,N_14449);
nand UO_1052 (O_1052,N_14877,N_14568);
or UO_1053 (O_1053,N_14248,N_14041);
xnor UO_1054 (O_1054,N_14532,N_14451);
nor UO_1055 (O_1055,N_14185,N_14632);
nand UO_1056 (O_1056,N_14957,N_14298);
or UO_1057 (O_1057,N_14448,N_14707);
or UO_1058 (O_1058,N_14012,N_14679);
xnor UO_1059 (O_1059,N_14510,N_14898);
or UO_1060 (O_1060,N_14981,N_14223);
nor UO_1061 (O_1061,N_14366,N_14667);
or UO_1062 (O_1062,N_14288,N_14418);
nand UO_1063 (O_1063,N_14456,N_14681);
nand UO_1064 (O_1064,N_14862,N_14005);
xnor UO_1065 (O_1065,N_14874,N_14984);
xnor UO_1066 (O_1066,N_14563,N_14746);
nand UO_1067 (O_1067,N_14243,N_14285);
nor UO_1068 (O_1068,N_14490,N_14283);
xnor UO_1069 (O_1069,N_14368,N_14073);
or UO_1070 (O_1070,N_14272,N_14101);
xnor UO_1071 (O_1071,N_14545,N_14672);
or UO_1072 (O_1072,N_14784,N_14951);
or UO_1073 (O_1073,N_14015,N_14930);
and UO_1074 (O_1074,N_14378,N_14670);
nand UO_1075 (O_1075,N_14950,N_14940);
and UO_1076 (O_1076,N_14146,N_14554);
xor UO_1077 (O_1077,N_14924,N_14090);
and UO_1078 (O_1078,N_14414,N_14760);
or UO_1079 (O_1079,N_14739,N_14925);
nand UO_1080 (O_1080,N_14908,N_14929);
nand UO_1081 (O_1081,N_14366,N_14910);
xnor UO_1082 (O_1082,N_14958,N_14314);
and UO_1083 (O_1083,N_14945,N_14708);
nor UO_1084 (O_1084,N_14024,N_14380);
or UO_1085 (O_1085,N_14017,N_14007);
nand UO_1086 (O_1086,N_14303,N_14436);
or UO_1087 (O_1087,N_14947,N_14177);
nor UO_1088 (O_1088,N_14597,N_14942);
nor UO_1089 (O_1089,N_14642,N_14703);
and UO_1090 (O_1090,N_14978,N_14051);
and UO_1091 (O_1091,N_14147,N_14754);
and UO_1092 (O_1092,N_14454,N_14031);
nor UO_1093 (O_1093,N_14382,N_14199);
nand UO_1094 (O_1094,N_14561,N_14090);
nor UO_1095 (O_1095,N_14197,N_14908);
or UO_1096 (O_1096,N_14778,N_14455);
nor UO_1097 (O_1097,N_14946,N_14190);
nand UO_1098 (O_1098,N_14254,N_14063);
nand UO_1099 (O_1099,N_14240,N_14203);
and UO_1100 (O_1100,N_14794,N_14136);
nand UO_1101 (O_1101,N_14028,N_14043);
and UO_1102 (O_1102,N_14113,N_14454);
xnor UO_1103 (O_1103,N_14243,N_14993);
or UO_1104 (O_1104,N_14219,N_14856);
nor UO_1105 (O_1105,N_14629,N_14782);
nor UO_1106 (O_1106,N_14551,N_14174);
or UO_1107 (O_1107,N_14144,N_14921);
or UO_1108 (O_1108,N_14200,N_14253);
and UO_1109 (O_1109,N_14366,N_14240);
nor UO_1110 (O_1110,N_14683,N_14331);
nor UO_1111 (O_1111,N_14970,N_14341);
or UO_1112 (O_1112,N_14963,N_14580);
nor UO_1113 (O_1113,N_14515,N_14587);
or UO_1114 (O_1114,N_14614,N_14440);
nor UO_1115 (O_1115,N_14454,N_14851);
and UO_1116 (O_1116,N_14717,N_14363);
xor UO_1117 (O_1117,N_14133,N_14852);
nor UO_1118 (O_1118,N_14988,N_14384);
xnor UO_1119 (O_1119,N_14539,N_14678);
and UO_1120 (O_1120,N_14738,N_14162);
or UO_1121 (O_1121,N_14039,N_14791);
nor UO_1122 (O_1122,N_14762,N_14459);
nor UO_1123 (O_1123,N_14746,N_14955);
nand UO_1124 (O_1124,N_14235,N_14749);
and UO_1125 (O_1125,N_14976,N_14092);
nand UO_1126 (O_1126,N_14888,N_14693);
and UO_1127 (O_1127,N_14285,N_14629);
and UO_1128 (O_1128,N_14134,N_14805);
and UO_1129 (O_1129,N_14954,N_14729);
nor UO_1130 (O_1130,N_14762,N_14221);
or UO_1131 (O_1131,N_14159,N_14464);
and UO_1132 (O_1132,N_14342,N_14925);
xor UO_1133 (O_1133,N_14929,N_14149);
nor UO_1134 (O_1134,N_14896,N_14533);
and UO_1135 (O_1135,N_14653,N_14707);
nand UO_1136 (O_1136,N_14001,N_14816);
nand UO_1137 (O_1137,N_14221,N_14474);
nand UO_1138 (O_1138,N_14431,N_14327);
or UO_1139 (O_1139,N_14729,N_14917);
or UO_1140 (O_1140,N_14352,N_14753);
and UO_1141 (O_1141,N_14365,N_14089);
and UO_1142 (O_1142,N_14245,N_14921);
nor UO_1143 (O_1143,N_14397,N_14979);
or UO_1144 (O_1144,N_14370,N_14064);
nor UO_1145 (O_1145,N_14598,N_14299);
and UO_1146 (O_1146,N_14563,N_14742);
or UO_1147 (O_1147,N_14360,N_14591);
or UO_1148 (O_1148,N_14609,N_14309);
nor UO_1149 (O_1149,N_14756,N_14539);
and UO_1150 (O_1150,N_14177,N_14313);
or UO_1151 (O_1151,N_14104,N_14524);
nand UO_1152 (O_1152,N_14340,N_14606);
nand UO_1153 (O_1153,N_14859,N_14254);
nand UO_1154 (O_1154,N_14470,N_14265);
nor UO_1155 (O_1155,N_14642,N_14735);
nor UO_1156 (O_1156,N_14771,N_14613);
nor UO_1157 (O_1157,N_14760,N_14853);
and UO_1158 (O_1158,N_14228,N_14270);
and UO_1159 (O_1159,N_14766,N_14541);
or UO_1160 (O_1160,N_14273,N_14174);
nor UO_1161 (O_1161,N_14503,N_14056);
xor UO_1162 (O_1162,N_14625,N_14919);
and UO_1163 (O_1163,N_14528,N_14150);
xor UO_1164 (O_1164,N_14276,N_14406);
or UO_1165 (O_1165,N_14573,N_14465);
nand UO_1166 (O_1166,N_14740,N_14796);
nor UO_1167 (O_1167,N_14660,N_14210);
nand UO_1168 (O_1168,N_14712,N_14348);
nand UO_1169 (O_1169,N_14634,N_14043);
or UO_1170 (O_1170,N_14878,N_14285);
or UO_1171 (O_1171,N_14642,N_14127);
or UO_1172 (O_1172,N_14412,N_14959);
nor UO_1173 (O_1173,N_14232,N_14055);
and UO_1174 (O_1174,N_14800,N_14241);
nor UO_1175 (O_1175,N_14498,N_14750);
or UO_1176 (O_1176,N_14901,N_14394);
and UO_1177 (O_1177,N_14267,N_14974);
nor UO_1178 (O_1178,N_14187,N_14276);
nand UO_1179 (O_1179,N_14092,N_14349);
and UO_1180 (O_1180,N_14904,N_14887);
or UO_1181 (O_1181,N_14203,N_14211);
and UO_1182 (O_1182,N_14819,N_14919);
and UO_1183 (O_1183,N_14601,N_14019);
xor UO_1184 (O_1184,N_14587,N_14055);
or UO_1185 (O_1185,N_14148,N_14298);
nor UO_1186 (O_1186,N_14325,N_14838);
nand UO_1187 (O_1187,N_14091,N_14109);
nor UO_1188 (O_1188,N_14202,N_14888);
and UO_1189 (O_1189,N_14421,N_14231);
or UO_1190 (O_1190,N_14732,N_14343);
nor UO_1191 (O_1191,N_14052,N_14905);
and UO_1192 (O_1192,N_14099,N_14896);
and UO_1193 (O_1193,N_14119,N_14491);
xor UO_1194 (O_1194,N_14440,N_14842);
and UO_1195 (O_1195,N_14980,N_14376);
or UO_1196 (O_1196,N_14784,N_14018);
and UO_1197 (O_1197,N_14449,N_14689);
nor UO_1198 (O_1198,N_14652,N_14621);
and UO_1199 (O_1199,N_14279,N_14480);
nor UO_1200 (O_1200,N_14934,N_14452);
nor UO_1201 (O_1201,N_14238,N_14007);
nand UO_1202 (O_1202,N_14121,N_14506);
nand UO_1203 (O_1203,N_14392,N_14555);
nand UO_1204 (O_1204,N_14862,N_14308);
or UO_1205 (O_1205,N_14374,N_14008);
and UO_1206 (O_1206,N_14921,N_14355);
or UO_1207 (O_1207,N_14109,N_14143);
or UO_1208 (O_1208,N_14818,N_14797);
or UO_1209 (O_1209,N_14539,N_14625);
nor UO_1210 (O_1210,N_14502,N_14173);
nor UO_1211 (O_1211,N_14221,N_14139);
and UO_1212 (O_1212,N_14297,N_14836);
or UO_1213 (O_1213,N_14197,N_14553);
or UO_1214 (O_1214,N_14091,N_14265);
and UO_1215 (O_1215,N_14717,N_14490);
and UO_1216 (O_1216,N_14655,N_14889);
or UO_1217 (O_1217,N_14330,N_14278);
nand UO_1218 (O_1218,N_14717,N_14664);
and UO_1219 (O_1219,N_14904,N_14929);
or UO_1220 (O_1220,N_14764,N_14311);
or UO_1221 (O_1221,N_14333,N_14682);
or UO_1222 (O_1222,N_14437,N_14383);
nand UO_1223 (O_1223,N_14022,N_14510);
and UO_1224 (O_1224,N_14083,N_14448);
nor UO_1225 (O_1225,N_14017,N_14268);
nor UO_1226 (O_1226,N_14690,N_14670);
nor UO_1227 (O_1227,N_14900,N_14046);
nor UO_1228 (O_1228,N_14458,N_14805);
and UO_1229 (O_1229,N_14598,N_14799);
and UO_1230 (O_1230,N_14555,N_14093);
nor UO_1231 (O_1231,N_14837,N_14664);
and UO_1232 (O_1232,N_14548,N_14291);
xnor UO_1233 (O_1233,N_14453,N_14260);
and UO_1234 (O_1234,N_14599,N_14960);
nand UO_1235 (O_1235,N_14443,N_14363);
nand UO_1236 (O_1236,N_14911,N_14954);
nand UO_1237 (O_1237,N_14235,N_14054);
or UO_1238 (O_1238,N_14701,N_14861);
and UO_1239 (O_1239,N_14987,N_14288);
nor UO_1240 (O_1240,N_14751,N_14178);
nor UO_1241 (O_1241,N_14993,N_14145);
and UO_1242 (O_1242,N_14264,N_14480);
and UO_1243 (O_1243,N_14424,N_14163);
nand UO_1244 (O_1244,N_14256,N_14647);
nor UO_1245 (O_1245,N_14321,N_14871);
nand UO_1246 (O_1246,N_14749,N_14537);
and UO_1247 (O_1247,N_14693,N_14110);
or UO_1248 (O_1248,N_14272,N_14631);
or UO_1249 (O_1249,N_14201,N_14106);
nand UO_1250 (O_1250,N_14802,N_14376);
nor UO_1251 (O_1251,N_14841,N_14371);
or UO_1252 (O_1252,N_14495,N_14553);
nor UO_1253 (O_1253,N_14766,N_14182);
and UO_1254 (O_1254,N_14079,N_14958);
xnor UO_1255 (O_1255,N_14638,N_14185);
nand UO_1256 (O_1256,N_14970,N_14508);
nor UO_1257 (O_1257,N_14875,N_14047);
nor UO_1258 (O_1258,N_14682,N_14581);
nor UO_1259 (O_1259,N_14111,N_14494);
xor UO_1260 (O_1260,N_14181,N_14441);
nor UO_1261 (O_1261,N_14984,N_14937);
nand UO_1262 (O_1262,N_14659,N_14279);
or UO_1263 (O_1263,N_14387,N_14492);
nor UO_1264 (O_1264,N_14754,N_14542);
nor UO_1265 (O_1265,N_14306,N_14288);
or UO_1266 (O_1266,N_14542,N_14256);
and UO_1267 (O_1267,N_14238,N_14750);
nor UO_1268 (O_1268,N_14234,N_14323);
nand UO_1269 (O_1269,N_14267,N_14657);
or UO_1270 (O_1270,N_14314,N_14151);
and UO_1271 (O_1271,N_14703,N_14561);
and UO_1272 (O_1272,N_14689,N_14290);
and UO_1273 (O_1273,N_14108,N_14262);
nand UO_1274 (O_1274,N_14512,N_14398);
and UO_1275 (O_1275,N_14355,N_14046);
or UO_1276 (O_1276,N_14059,N_14506);
and UO_1277 (O_1277,N_14962,N_14650);
xnor UO_1278 (O_1278,N_14138,N_14408);
or UO_1279 (O_1279,N_14713,N_14764);
or UO_1280 (O_1280,N_14961,N_14631);
or UO_1281 (O_1281,N_14700,N_14917);
and UO_1282 (O_1282,N_14860,N_14147);
and UO_1283 (O_1283,N_14183,N_14699);
nand UO_1284 (O_1284,N_14793,N_14893);
and UO_1285 (O_1285,N_14086,N_14529);
nand UO_1286 (O_1286,N_14901,N_14932);
nor UO_1287 (O_1287,N_14599,N_14819);
or UO_1288 (O_1288,N_14870,N_14425);
nand UO_1289 (O_1289,N_14786,N_14480);
nand UO_1290 (O_1290,N_14146,N_14733);
or UO_1291 (O_1291,N_14433,N_14010);
or UO_1292 (O_1292,N_14843,N_14490);
nor UO_1293 (O_1293,N_14848,N_14045);
nor UO_1294 (O_1294,N_14928,N_14140);
nor UO_1295 (O_1295,N_14884,N_14285);
and UO_1296 (O_1296,N_14444,N_14551);
or UO_1297 (O_1297,N_14067,N_14830);
nand UO_1298 (O_1298,N_14923,N_14784);
nand UO_1299 (O_1299,N_14086,N_14710);
xor UO_1300 (O_1300,N_14666,N_14164);
or UO_1301 (O_1301,N_14568,N_14864);
nor UO_1302 (O_1302,N_14361,N_14423);
nor UO_1303 (O_1303,N_14464,N_14730);
nor UO_1304 (O_1304,N_14203,N_14538);
or UO_1305 (O_1305,N_14336,N_14025);
or UO_1306 (O_1306,N_14303,N_14910);
nand UO_1307 (O_1307,N_14443,N_14084);
or UO_1308 (O_1308,N_14163,N_14885);
or UO_1309 (O_1309,N_14314,N_14698);
nand UO_1310 (O_1310,N_14472,N_14894);
nor UO_1311 (O_1311,N_14629,N_14193);
and UO_1312 (O_1312,N_14318,N_14356);
xor UO_1313 (O_1313,N_14301,N_14113);
or UO_1314 (O_1314,N_14383,N_14213);
nor UO_1315 (O_1315,N_14950,N_14131);
nand UO_1316 (O_1316,N_14021,N_14116);
and UO_1317 (O_1317,N_14805,N_14757);
nor UO_1318 (O_1318,N_14200,N_14450);
nand UO_1319 (O_1319,N_14094,N_14276);
and UO_1320 (O_1320,N_14353,N_14697);
and UO_1321 (O_1321,N_14761,N_14553);
xor UO_1322 (O_1322,N_14052,N_14538);
nand UO_1323 (O_1323,N_14642,N_14793);
or UO_1324 (O_1324,N_14059,N_14353);
and UO_1325 (O_1325,N_14344,N_14314);
or UO_1326 (O_1326,N_14277,N_14273);
nor UO_1327 (O_1327,N_14665,N_14289);
and UO_1328 (O_1328,N_14323,N_14859);
nand UO_1329 (O_1329,N_14903,N_14898);
and UO_1330 (O_1330,N_14539,N_14698);
nor UO_1331 (O_1331,N_14693,N_14461);
or UO_1332 (O_1332,N_14840,N_14144);
or UO_1333 (O_1333,N_14720,N_14396);
nand UO_1334 (O_1334,N_14170,N_14803);
nand UO_1335 (O_1335,N_14977,N_14268);
nor UO_1336 (O_1336,N_14021,N_14043);
nor UO_1337 (O_1337,N_14157,N_14620);
and UO_1338 (O_1338,N_14370,N_14289);
and UO_1339 (O_1339,N_14657,N_14581);
or UO_1340 (O_1340,N_14263,N_14480);
nand UO_1341 (O_1341,N_14739,N_14999);
or UO_1342 (O_1342,N_14257,N_14827);
xor UO_1343 (O_1343,N_14891,N_14569);
nor UO_1344 (O_1344,N_14247,N_14889);
nand UO_1345 (O_1345,N_14531,N_14723);
or UO_1346 (O_1346,N_14658,N_14049);
xor UO_1347 (O_1347,N_14052,N_14795);
and UO_1348 (O_1348,N_14443,N_14541);
nand UO_1349 (O_1349,N_14605,N_14516);
and UO_1350 (O_1350,N_14603,N_14516);
nand UO_1351 (O_1351,N_14488,N_14263);
xor UO_1352 (O_1352,N_14926,N_14935);
nand UO_1353 (O_1353,N_14680,N_14016);
and UO_1354 (O_1354,N_14526,N_14950);
and UO_1355 (O_1355,N_14303,N_14773);
nor UO_1356 (O_1356,N_14662,N_14524);
nand UO_1357 (O_1357,N_14765,N_14642);
nor UO_1358 (O_1358,N_14229,N_14745);
nor UO_1359 (O_1359,N_14604,N_14756);
nor UO_1360 (O_1360,N_14763,N_14894);
nand UO_1361 (O_1361,N_14607,N_14645);
and UO_1362 (O_1362,N_14117,N_14006);
nor UO_1363 (O_1363,N_14560,N_14826);
nor UO_1364 (O_1364,N_14364,N_14801);
and UO_1365 (O_1365,N_14548,N_14838);
nor UO_1366 (O_1366,N_14154,N_14773);
nand UO_1367 (O_1367,N_14430,N_14204);
and UO_1368 (O_1368,N_14304,N_14344);
nand UO_1369 (O_1369,N_14322,N_14676);
or UO_1370 (O_1370,N_14721,N_14073);
nand UO_1371 (O_1371,N_14444,N_14518);
xor UO_1372 (O_1372,N_14373,N_14431);
nor UO_1373 (O_1373,N_14473,N_14718);
nand UO_1374 (O_1374,N_14800,N_14051);
or UO_1375 (O_1375,N_14621,N_14655);
nor UO_1376 (O_1376,N_14796,N_14876);
and UO_1377 (O_1377,N_14272,N_14017);
and UO_1378 (O_1378,N_14809,N_14593);
nand UO_1379 (O_1379,N_14067,N_14489);
nor UO_1380 (O_1380,N_14625,N_14717);
and UO_1381 (O_1381,N_14668,N_14110);
nand UO_1382 (O_1382,N_14555,N_14396);
or UO_1383 (O_1383,N_14130,N_14373);
and UO_1384 (O_1384,N_14508,N_14075);
or UO_1385 (O_1385,N_14714,N_14644);
or UO_1386 (O_1386,N_14011,N_14901);
nor UO_1387 (O_1387,N_14920,N_14187);
nor UO_1388 (O_1388,N_14255,N_14538);
nand UO_1389 (O_1389,N_14383,N_14036);
or UO_1390 (O_1390,N_14624,N_14935);
nand UO_1391 (O_1391,N_14551,N_14467);
nor UO_1392 (O_1392,N_14965,N_14808);
or UO_1393 (O_1393,N_14777,N_14374);
or UO_1394 (O_1394,N_14819,N_14893);
nor UO_1395 (O_1395,N_14846,N_14124);
nor UO_1396 (O_1396,N_14082,N_14837);
nor UO_1397 (O_1397,N_14750,N_14986);
and UO_1398 (O_1398,N_14695,N_14131);
or UO_1399 (O_1399,N_14593,N_14436);
xnor UO_1400 (O_1400,N_14120,N_14923);
nor UO_1401 (O_1401,N_14472,N_14862);
xor UO_1402 (O_1402,N_14333,N_14456);
nand UO_1403 (O_1403,N_14164,N_14143);
or UO_1404 (O_1404,N_14735,N_14381);
nor UO_1405 (O_1405,N_14774,N_14487);
nor UO_1406 (O_1406,N_14179,N_14612);
or UO_1407 (O_1407,N_14643,N_14850);
or UO_1408 (O_1408,N_14236,N_14946);
and UO_1409 (O_1409,N_14352,N_14966);
nand UO_1410 (O_1410,N_14515,N_14960);
nor UO_1411 (O_1411,N_14090,N_14510);
nor UO_1412 (O_1412,N_14126,N_14616);
or UO_1413 (O_1413,N_14733,N_14942);
and UO_1414 (O_1414,N_14154,N_14156);
nor UO_1415 (O_1415,N_14951,N_14371);
and UO_1416 (O_1416,N_14411,N_14611);
or UO_1417 (O_1417,N_14336,N_14156);
xnor UO_1418 (O_1418,N_14034,N_14133);
and UO_1419 (O_1419,N_14952,N_14651);
nor UO_1420 (O_1420,N_14427,N_14262);
nor UO_1421 (O_1421,N_14042,N_14643);
or UO_1422 (O_1422,N_14915,N_14465);
or UO_1423 (O_1423,N_14073,N_14015);
xor UO_1424 (O_1424,N_14623,N_14521);
and UO_1425 (O_1425,N_14352,N_14138);
xor UO_1426 (O_1426,N_14258,N_14262);
xor UO_1427 (O_1427,N_14392,N_14172);
or UO_1428 (O_1428,N_14163,N_14285);
nand UO_1429 (O_1429,N_14312,N_14755);
nand UO_1430 (O_1430,N_14649,N_14852);
and UO_1431 (O_1431,N_14811,N_14507);
and UO_1432 (O_1432,N_14213,N_14751);
nand UO_1433 (O_1433,N_14548,N_14859);
nand UO_1434 (O_1434,N_14419,N_14650);
and UO_1435 (O_1435,N_14881,N_14219);
nor UO_1436 (O_1436,N_14012,N_14241);
and UO_1437 (O_1437,N_14702,N_14025);
xor UO_1438 (O_1438,N_14687,N_14652);
or UO_1439 (O_1439,N_14722,N_14270);
xnor UO_1440 (O_1440,N_14051,N_14157);
nor UO_1441 (O_1441,N_14769,N_14807);
or UO_1442 (O_1442,N_14264,N_14530);
nor UO_1443 (O_1443,N_14735,N_14751);
nand UO_1444 (O_1444,N_14084,N_14586);
or UO_1445 (O_1445,N_14071,N_14103);
nand UO_1446 (O_1446,N_14382,N_14530);
nand UO_1447 (O_1447,N_14722,N_14163);
or UO_1448 (O_1448,N_14369,N_14289);
or UO_1449 (O_1449,N_14559,N_14632);
and UO_1450 (O_1450,N_14284,N_14114);
and UO_1451 (O_1451,N_14720,N_14823);
nand UO_1452 (O_1452,N_14540,N_14793);
and UO_1453 (O_1453,N_14183,N_14125);
nor UO_1454 (O_1454,N_14514,N_14494);
and UO_1455 (O_1455,N_14115,N_14906);
or UO_1456 (O_1456,N_14840,N_14444);
nand UO_1457 (O_1457,N_14511,N_14454);
or UO_1458 (O_1458,N_14565,N_14297);
nor UO_1459 (O_1459,N_14563,N_14264);
and UO_1460 (O_1460,N_14760,N_14285);
and UO_1461 (O_1461,N_14781,N_14072);
nand UO_1462 (O_1462,N_14673,N_14500);
nor UO_1463 (O_1463,N_14709,N_14679);
nand UO_1464 (O_1464,N_14027,N_14028);
nand UO_1465 (O_1465,N_14758,N_14254);
nand UO_1466 (O_1466,N_14877,N_14964);
xor UO_1467 (O_1467,N_14860,N_14841);
nand UO_1468 (O_1468,N_14411,N_14157);
nor UO_1469 (O_1469,N_14642,N_14087);
xor UO_1470 (O_1470,N_14003,N_14918);
and UO_1471 (O_1471,N_14218,N_14585);
or UO_1472 (O_1472,N_14918,N_14649);
nor UO_1473 (O_1473,N_14485,N_14149);
nor UO_1474 (O_1474,N_14982,N_14222);
or UO_1475 (O_1475,N_14610,N_14069);
and UO_1476 (O_1476,N_14889,N_14654);
nor UO_1477 (O_1477,N_14048,N_14008);
or UO_1478 (O_1478,N_14525,N_14488);
or UO_1479 (O_1479,N_14724,N_14405);
or UO_1480 (O_1480,N_14427,N_14152);
nand UO_1481 (O_1481,N_14300,N_14183);
nor UO_1482 (O_1482,N_14991,N_14720);
nand UO_1483 (O_1483,N_14991,N_14248);
nor UO_1484 (O_1484,N_14831,N_14104);
nand UO_1485 (O_1485,N_14363,N_14015);
xnor UO_1486 (O_1486,N_14499,N_14051);
nor UO_1487 (O_1487,N_14939,N_14244);
nor UO_1488 (O_1488,N_14654,N_14624);
or UO_1489 (O_1489,N_14630,N_14135);
and UO_1490 (O_1490,N_14642,N_14528);
and UO_1491 (O_1491,N_14867,N_14618);
xor UO_1492 (O_1492,N_14132,N_14226);
nor UO_1493 (O_1493,N_14947,N_14437);
nand UO_1494 (O_1494,N_14511,N_14613);
or UO_1495 (O_1495,N_14909,N_14561);
or UO_1496 (O_1496,N_14670,N_14032);
and UO_1497 (O_1497,N_14311,N_14183);
nor UO_1498 (O_1498,N_14049,N_14163);
nor UO_1499 (O_1499,N_14739,N_14956);
and UO_1500 (O_1500,N_14094,N_14708);
and UO_1501 (O_1501,N_14344,N_14169);
and UO_1502 (O_1502,N_14780,N_14544);
or UO_1503 (O_1503,N_14861,N_14170);
and UO_1504 (O_1504,N_14498,N_14055);
nand UO_1505 (O_1505,N_14697,N_14350);
nor UO_1506 (O_1506,N_14939,N_14928);
and UO_1507 (O_1507,N_14933,N_14091);
nor UO_1508 (O_1508,N_14019,N_14899);
or UO_1509 (O_1509,N_14193,N_14386);
and UO_1510 (O_1510,N_14021,N_14130);
or UO_1511 (O_1511,N_14704,N_14649);
xor UO_1512 (O_1512,N_14380,N_14521);
and UO_1513 (O_1513,N_14452,N_14372);
and UO_1514 (O_1514,N_14195,N_14810);
nand UO_1515 (O_1515,N_14559,N_14466);
or UO_1516 (O_1516,N_14350,N_14603);
and UO_1517 (O_1517,N_14827,N_14334);
nor UO_1518 (O_1518,N_14362,N_14880);
nor UO_1519 (O_1519,N_14400,N_14595);
nor UO_1520 (O_1520,N_14250,N_14495);
nand UO_1521 (O_1521,N_14988,N_14329);
nor UO_1522 (O_1522,N_14171,N_14281);
xor UO_1523 (O_1523,N_14891,N_14089);
nor UO_1524 (O_1524,N_14699,N_14003);
and UO_1525 (O_1525,N_14504,N_14614);
nor UO_1526 (O_1526,N_14579,N_14388);
nand UO_1527 (O_1527,N_14770,N_14824);
xor UO_1528 (O_1528,N_14070,N_14116);
and UO_1529 (O_1529,N_14535,N_14751);
nand UO_1530 (O_1530,N_14774,N_14068);
nor UO_1531 (O_1531,N_14797,N_14245);
nor UO_1532 (O_1532,N_14692,N_14970);
nand UO_1533 (O_1533,N_14075,N_14191);
or UO_1534 (O_1534,N_14851,N_14086);
nand UO_1535 (O_1535,N_14210,N_14609);
and UO_1536 (O_1536,N_14536,N_14531);
and UO_1537 (O_1537,N_14483,N_14678);
nand UO_1538 (O_1538,N_14188,N_14606);
nand UO_1539 (O_1539,N_14342,N_14056);
nor UO_1540 (O_1540,N_14067,N_14496);
xnor UO_1541 (O_1541,N_14979,N_14671);
xnor UO_1542 (O_1542,N_14274,N_14133);
xor UO_1543 (O_1543,N_14203,N_14300);
nor UO_1544 (O_1544,N_14522,N_14324);
and UO_1545 (O_1545,N_14607,N_14217);
nand UO_1546 (O_1546,N_14471,N_14615);
nand UO_1547 (O_1547,N_14857,N_14617);
and UO_1548 (O_1548,N_14247,N_14421);
nand UO_1549 (O_1549,N_14695,N_14765);
or UO_1550 (O_1550,N_14341,N_14047);
or UO_1551 (O_1551,N_14456,N_14002);
and UO_1552 (O_1552,N_14035,N_14805);
xnor UO_1553 (O_1553,N_14835,N_14899);
or UO_1554 (O_1554,N_14021,N_14721);
or UO_1555 (O_1555,N_14391,N_14171);
nor UO_1556 (O_1556,N_14601,N_14431);
and UO_1557 (O_1557,N_14492,N_14997);
nand UO_1558 (O_1558,N_14131,N_14897);
and UO_1559 (O_1559,N_14188,N_14621);
xor UO_1560 (O_1560,N_14438,N_14131);
and UO_1561 (O_1561,N_14578,N_14431);
or UO_1562 (O_1562,N_14069,N_14813);
nor UO_1563 (O_1563,N_14537,N_14306);
nor UO_1564 (O_1564,N_14993,N_14337);
xnor UO_1565 (O_1565,N_14476,N_14673);
xor UO_1566 (O_1566,N_14098,N_14950);
nand UO_1567 (O_1567,N_14116,N_14690);
and UO_1568 (O_1568,N_14931,N_14176);
nand UO_1569 (O_1569,N_14149,N_14616);
nor UO_1570 (O_1570,N_14486,N_14050);
or UO_1571 (O_1571,N_14731,N_14968);
or UO_1572 (O_1572,N_14638,N_14235);
xnor UO_1573 (O_1573,N_14923,N_14275);
or UO_1574 (O_1574,N_14686,N_14111);
nand UO_1575 (O_1575,N_14151,N_14505);
nand UO_1576 (O_1576,N_14962,N_14239);
nor UO_1577 (O_1577,N_14842,N_14360);
nand UO_1578 (O_1578,N_14780,N_14003);
or UO_1579 (O_1579,N_14086,N_14202);
nor UO_1580 (O_1580,N_14694,N_14097);
and UO_1581 (O_1581,N_14358,N_14670);
and UO_1582 (O_1582,N_14421,N_14245);
or UO_1583 (O_1583,N_14208,N_14769);
nor UO_1584 (O_1584,N_14961,N_14750);
or UO_1585 (O_1585,N_14441,N_14262);
xor UO_1586 (O_1586,N_14364,N_14691);
nor UO_1587 (O_1587,N_14641,N_14339);
nand UO_1588 (O_1588,N_14574,N_14484);
nand UO_1589 (O_1589,N_14592,N_14621);
or UO_1590 (O_1590,N_14374,N_14539);
nand UO_1591 (O_1591,N_14463,N_14663);
or UO_1592 (O_1592,N_14533,N_14454);
or UO_1593 (O_1593,N_14522,N_14967);
xnor UO_1594 (O_1594,N_14887,N_14338);
or UO_1595 (O_1595,N_14263,N_14634);
nand UO_1596 (O_1596,N_14374,N_14280);
or UO_1597 (O_1597,N_14738,N_14172);
or UO_1598 (O_1598,N_14455,N_14341);
or UO_1599 (O_1599,N_14095,N_14456);
nor UO_1600 (O_1600,N_14132,N_14171);
nand UO_1601 (O_1601,N_14690,N_14984);
xor UO_1602 (O_1602,N_14900,N_14345);
nand UO_1603 (O_1603,N_14338,N_14917);
nor UO_1604 (O_1604,N_14019,N_14270);
nand UO_1605 (O_1605,N_14784,N_14684);
nor UO_1606 (O_1606,N_14747,N_14609);
or UO_1607 (O_1607,N_14651,N_14318);
or UO_1608 (O_1608,N_14072,N_14712);
nor UO_1609 (O_1609,N_14088,N_14884);
nor UO_1610 (O_1610,N_14242,N_14427);
and UO_1611 (O_1611,N_14029,N_14573);
and UO_1612 (O_1612,N_14989,N_14796);
xor UO_1613 (O_1613,N_14907,N_14194);
nor UO_1614 (O_1614,N_14367,N_14868);
nand UO_1615 (O_1615,N_14726,N_14155);
nor UO_1616 (O_1616,N_14945,N_14051);
and UO_1617 (O_1617,N_14451,N_14311);
nand UO_1618 (O_1618,N_14772,N_14846);
nand UO_1619 (O_1619,N_14151,N_14228);
or UO_1620 (O_1620,N_14376,N_14144);
nand UO_1621 (O_1621,N_14073,N_14486);
nor UO_1622 (O_1622,N_14439,N_14004);
or UO_1623 (O_1623,N_14381,N_14003);
nand UO_1624 (O_1624,N_14431,N_14794);
xor UO_1625 (O_1625,N_14740,N_14913);
or UO_1626 (O_1626,N_14764,N_14801);
xor UO_1627 (O_1627,N_14335,N_14984);
nand UO_1628 (O_1628,N_14186,N_14485);
and UO_1629 (O_1629,N_14839,N_14571);
nand UO_1630 (O_1630,N_14150,N_14291);
or UO_1631 (O_1631,N_14928,N_14715);
nor UO_1632 (O_1632,N_14976,N_14999);
nand UO_1633 (O_1633,N_14065,N_14456);
nor UO_1634 (O_1634,N_14841,N_14282);
nor UO_1635 (O_1635,N_14960,N_14338);
and UO_1636 (O_1636,N_14698,N_14628);
and UO_1637 (O_1637,N_14220,N_14291);
nand UO_1638 (O_1638,N_14399,N_14286);
nand UO_1639 (O_1639,N_14163,N_14680);
and UO_1640 (O_1640,N_14016,N_14263);
xnor UO_1641 (O_1641,N_14848,N_14584);
nand UO_1642 (O_1642,N_14291,N_14806);
nand UO_1643 (O_1643,N_14321,N_14654);
or UO_1644 (O_1644,N_14029,N_14478);
xor UO_1645 (O_1645,N_14762,N_14228);
nand UO_1646 (O_1646,N_14208,N_14296);
or UO_1647 (O_1647,N_14470,N_14659);
nor UO_1648 (O_1648,N_14038,N_14766);
nand UO_1649 (O_1649,N_14080,N_14522);
or UO_1650 (O_1650,N_14678,N_14536);
nor UO_1651 (O_1651,N_14658,N_14883);
or UO_1652 (O_1652,N_14184,N_14445);
nor UO_1653 (O_1653,N_14733,N_14411);
nand UO_1654 (O_1654,N_14373,N_14483);
xnor UO_1655 (O_1655,N_14127,N_14858);
nand UO_1656 (O_1656,N_14495,N_14538);
or UO_1657 (O_1657,N_14323,N_14803);
nand UO_1658 (O_1658,N_14982,N_14589);
and UO_1659 (O_1659,N_14808,N_14228);
nor UO_1660 (O_1660,N_14990,N_14786);
nand UO_1661 (O_1661,N_14959,N_14852);
nor UO_1662 (O_1662,N_14866,N_14387);
nor UO_1663 (O_1663,N_14524,N_14186);
and UO_1664 (O_1664,N_14422,N_14292);
and UO_1665 (O_1665,N_14184,N_14592);
xor UO_1666 (O_1666,N_14255,N_14686);
nand UO_1667 (O_1667,N_14749,N_14442);
and UO_1668 (O_1668,N_14307,N_14354);
nand UO_1669 (O_1669,N_14937,N_14272);
nor UO_1670 (O_1670,N_14124,N_14160);
or UO_1671 (O_1671,N_14913,N_14599);
or UO_1672 (O_1672,N_14508,N_14507);
nor UO_1673 (O_1673,N_14597,N_14415);
nor UO_1674 (O_1674,N_14469,N_14270);
nand UO_1675 (O_1675,N_14336,N_14861);
or UO_1676 (O_1676,N_14736,N_14562);
or UO_1677 (O_1677,N_14532,N_14746);
and UO_1678 (O_1678,N_14422,N_14549);
nor UO_1679 (O_1679,N_14169,N_14176);
nand UO_1680 (O_1680,N_14989,N_14790);
xnor UO_1681 (O_1681,N_14538,N_14225);
and UO_1682 (O_1682,N_14319,N_14750);
or UO_1683 (O_1683,N_14540,N_14817);
nor UO_1684 (O_1684,N_14072,N_14017);
nor UO_1685 (O_1685,N_14494,N_14822);
or UO_1686 (O_1686,N_14166,N_14397);
and UO_1687 (O_1687,N_14934,N_14365);
or UO_1688 (O_1688,N_14782,N_14057);
or UO_1689 (O_1689,N_14085,N_14904);
nand UO_1690 (O_1690,N_14363,N_14597);
nand UO_1691 (O_1691,N_14414,N_14097);
or UO_1692 (O_1692,N_14693,N_14993);
and UO_1693 (O_1693,N_14478,N_14687);
nor UO_1694 (O_1694,N_14031,N_14038);
nor UO_1695 (O_1695,N_14612,N_14630);
nand UO_1696 (O_1696,N_14977,N_14908);
or UO_1697 (O_1697,N_14574,N_14227);
or UO_1698 (O_1698,N_14061,N_14774);
nand UO_1699 (O_1699,N_14957,N_14762);
nor UO_1700 (O_1700,N_14461,N_14408);
and UO_1701 (O_1701,N_14865,N_14958);
and UO_1702 (O_1702,N_14432,N_14613);
nor UO_1703 (O_1703,N_14054,N_14004);
nor UO_1704 (O_1704,N_14338,N_14769);
xnor UO_1705 (O_1705,N_14811,N_14677);
nor UO_1706 (O_1706,N_14133,N_14514);
or UO_1707 (O_1707,N_14824,N_14479);
nor UO_1708 (O_1708,N_14144,N_14092);
and UO_1709 (O_1709,N_14788,N_14019);
xor UO_1710 (O_1710,N_14228,N_14969);
or UO_1711 (O_1711,N_14217,N_14810);
or UO_1712 (O_1712,N_14752,N_14268);
and UO_1713 (O_1713,N_14644,N_14256);
or UO_1714 (O_1714,N_14852,N_14012);
nor UO_1715 (O_1715,N_14384,N_14064);
nand UO_1716 (O_1716,N_14541,N_14515);
nor UO_1717 (O_1717,N_14520,N_14005);
or UO_1718 (O_1718,N_14334,N_14749);
nor UO_1719 (O_1719,N_14835,N_14365);
nand UO_1720 (O_1720,N_14861,N_14130);
nand UO_1721 (O_1721,N_14239,N_14401);
xnor UO_1722 (O_1722,N_14759,N_14053);
nor UO_1723 (O_1723,N_14747,N_14857);
nor UO_1724 (O_1724,N_14990,N_14138);
nor UO_1725 (O_1725,N_14442,N_14014);
or UO_1726 (O_1726,N_14307,N_14296);
nor UO_1727 (O_1727,N_14664,N_14449);
nor UO_1728 (O_1728,N_14977,N_14278);
nor UO_1729 (O_1729,N_14298,N_14104);
or UO_1730 (O_1730,N_14941,N_14895);
or UO_1731 (O_1731,N_14831,N_14439);
or UO_1732 (O_1732,N_14017,N_14539);
or UO_1733 (O_1733,N_14693,N_14296);
nand UO_1734 (O_1734,N_14943,N_14877);
nand UO_1735 (O_1735,N_14713,N_14724);
nor UO_1736 (O_1736,N_14930,N_14142);
and UO_1737 (O_1737,N_14331,N_14974);
and UO_1738 (O_1738,N_14106,N_14020);
and UO_1739 (O_1739,N_14482,N_14094);
and UO_1740 (O_1740,N_14184,N_14303);
or UO_1741 (O_1741,N_14750,N_14450);
or UO_1742 (O_1742,N_14278,N_14405);
nor UO_1743 (O_1743,N_14690,N_14583);
nand UO_1744 (O_1744,N_14360,N_14644);
or UO_1745 (O_1745,N_14264,N_14832);
and UO_1746 (O_1746,N_14450,N_14615);
and UO_1747 (O_1747,N_14764,N_14559);
or UO_1748 (O_1748,N_14829,N_14915);
nand UO_1749 (O_1749,N_14976,N_14663);
and UO_1750 (O_1750,N_14680,N_14902);
xnor UO_1751 (O_1751,N_14968,N_14949);
and UO_1752 (O_1752,N_14854,N_14563);
and UO_1753 (O_1753,N_14895,N_14354);
and UO_1754 (O_1754,N_14049,N_14773);
nor UO_1755 (O_1755,N_14872,N_14304);
and UO_1756 (O_1756,N_14533,N_14028);
nand UO_1757 (O_1757,N_14260,N_14421);
nand UO_1758 (O_1758,N_14469,N_14303);
or UO_1759 (O_1759,N_14324,N_14508);
or UO_1760 (O_1760,N_14627,N_14906);
xor UO_1761 (O_1761,N_14992,N_14638);
or UO_1762 (O_1762,N_14390,N_14934);
or UO_1763 (O_1763,N_14613,N_14104);
and UO_1764 (O_1764,N_14711,N_14691);
xnor UO_1765 (O_1765,N_14885,N_14712);
and UO_1766 (O_1766,N_14592,N_14023);
nand UO_1767 (O_1767,N_14649,N_14566);
nor UO_1768 (O_1768,N_14513,N_14677);
xnor UO_1769 (O_1769,N_14795,N_14392);
or UO_1770 (O_1770,N_14768,N_14871);
and UO_1771 (O_1771,N_14545,N_14096);
or UO_1772 (O_1772,N_14999,N_14188);
nand UO_1773 (O_1773,N_14425,N_14423);
nor UO_1774 (O_1774,N_14471,N_14139);
or UO_1775 (O_1775,N_14029,N_14921);
nand UO_1776 (O_1776,N_14556,N_14272);
nand UO_1777 (O_1777,N_14221,N_14754);
and UO_1778 (O_1778,N_14428,N_14285);
nand UO_1779 (O_1779,N_14541,N_14552);
and UO_1780 (O_1780,N_14423,N_14907);
nand UO_1781 (O_1781,N_14484,N_14727);
nor UO_1782 (O_1782,N_14862,N_14545);
and UO_1783 (O_1783,N_14642,N_14757);
and UO_1784 (O_1784,N_14121,N_14104);
or UO_1785 (O_1785,N_14338,N_14640);
and UO_1786 (O_1786,N_14914,N_14625);
and UO_1787 (O_1787,N_14351,N_14368);
or UO_1788 (O_1788,N_14093,N_14070);
and UO_1789 (O_1789,N_14012,N_14864);
xor UO_1790 (O_1790,N_14042,N_14797);
nand UO_1791 (O_1791,N_14215,N_14826);
or UO_1792 (O_1792,N_14371,N_14222);
or UO_1793 (O_1793,N_14174,N_14178);
or UO_1794 (O_1794,N_14424,N_14481);
nor UO_1795 (O_1795,N_14036,N_14663);
nand UO_1796 (O_1796,N_14357,N_14263);
xor UO_1797 (O_1797,N_14705,N_14599);
nor UO_1798 (O_1798,N_14402,N_14077);
and UO_1799 (O_1799,N_14336,N_14877);
xnor UO_1800 (O_1800,N_14571,N_14713);
nand UO_1801 (O_1801,N_14620,N_14178);
and UO_1802 (O_1802,N_14612,N_14848);
or UO_1803 (O_1803,N_14199,N_14643);
nor UO_1804 (O_1804,N_14809,N_14533);
xor UO_1805 (O_1805,N_14181,N_14231);
nand UO_1806 (O_1806,N_14309,N_14003);
and UO_1807 (O_1807,N_14622,N_14055);
or UO_1808 (O_1808,N_14962,N_14414);
nand UO_1809 (O_1809,N_14338,N_14828);
nor UO_1810 (O_1810,N_14005,N_14789);
xor UO_1811 (O_1811,N_14429,N_14364);
nor UO_1812 (O_1812,N_14952,N_14117);
nand UO_1813 (O_1813,N_14204,N_14947);
nand UO_1814 (O_1814,N_14032,N_14569);
and UO_1815 (O_1815,N_14115,N_14069);
nand UO_1816 (O_1816,N_14186,N_14310);
and UO_1817 (O_1817,N_14991,N_14077);
or UO_1818 (O_1818,N_14632,N_14815);
nor UO_1819 (O_1819,N_14017,N_14350);
nor UO_1820 (O_1820,N_14520,N_14100);
or UO_1821 (O_1821,N_14349,N_14577);
nor UO_1822 (O_1822,N_14382,N_14582);
or UO_1823 (O_1823,N_14483,N_14752);
or UO_1824 (O_1824,N_14493,N_14813);
nor UO_1825 (O_1825,N_14967,N_14147);
nand UO_1826 (O_1826,N_14597,N_14416);
or UO_1827 (O_1827,N_14779,N_14268);
or UO_1828 (O_1828,N_14543,N_14226);
and UO_1829 (O_1829,N_14955,N_14285);
nor UO_1830 (O_1830,N_14695,N_14887);
nor UO_1831 (O_1831,N_14348,N_14694);
xor UO_1832 (O_1832,N_14571,N_14883);
nor UO_1833 (O_1833,N_14954,N_14189);
xor UO_1834 (O_1834,N_14938,N_14397);
xnor UO_1835 (O_1835,N_14965,N_14240);
and UO_1836 (O_1836,N_14448,N_14455);
or UO_1837 (O_1837,N_14616,N_14304);
nor UO_1838 (O_1838,N_14041,N_14317);
or UO_1839 (O_1839,N_14771,N_14180);
nand UO_1840 (O_1840,N_14272,N_14920);
and UO_1841 (O_1841,N_14262,N_14063);
and UO_1842 (O_1842,N_14086,N_14643);
and UO_1843 (O_1843,N_14598,N_14793);
or UO_1844 (O_1844,N_14944,N_14612);
nand UO_1845 (O_1845,N_14693,N_14656);
nand UO_1846 (O_1846,N_14971,N_14871);
nand UO_1847 (O_1847,N_14476,N_14591);
or UO_1848 (O_1848,N_14187,N_14280);
or UO_1849 (O_1849,N_14209,N_14777);
and UO_1850 (O_1850,N_14792,N_14551);
and UO_1851 (O_1851,N_14854,N_14382);
nor UO_1852 (O_1852,N_14752,N_14766);
and UO_1853 (O_1853,N_14785,N_14850);
or UO_1854 (O_1854,N_14232,N_14867);
xor UO_1855 (O_1855,N_14964,N_14731);
and UO_1856 (O_1856,N_14956,N_14303);
nor UO_1857 (O_1857,N_14322,N_14020);
xnor UO_1858 (O_1858,N_14424,N_14362);
nor UO_1859 (O_1859,N_14765,N_14288);
and UO_1860 (O_1860,N_14221,N_14657);
or UO_1861 (O_1861,N_14449,N_14730);
xor UO_1862 (O_1862,N_14899,N_14277);
nor UO_1863 (O_1863,N_14306,N_14631);
nand UO_1864 (O_1864,N_14255,N_14376);
nor UO_1865 (O_1865,N_14776,N_14061);
and UO_1866 (O_1866,N_14356,N_14106);
or UO_1867 (O_1867,N_14209,N_14597);
nand UO_1868 (O_1868,N_14085,N_14227);
nor UO_1869 (O_1869,N_14547,N_14839);
or UO_1870 (O_1870,N_14191,N_14493);
and UO_1871 (O_1871,N_14723,N_14978);
nand UO_1872 (O_1872,N_14733,N_14949);
and UO_1873 (O_1873,N_14414,N_14130);
and UO_1874 (O_1874,N_14910,N_14332);
nand UO_1875 (O_1875,N_14061,N_14233);
or UO_1876 (O_1876,N_14211,N_14908);
and UO_1877 (O_1877,N_14460,N_14736);
or UO_1878 (O_1878,N_14263,N_14569);
nor UO_1879 (O_1879,N_14250,N_14109);
and UO_1880 (O_1880,N_14837,N_14602);
nor UO_1881 (O_1881,N_14686,N_14697);
and UO_1882 (O_1882,N_14876,N_14129);
and UO_1883 (O_1883,N_14598,N_14998);
and UO_1884 (O_1884,N_14352,N_14237);
nor UO_1885 (O_1885,N_14651,N_14955);
nor UO_1886 (O_1886,N_14225,N_14933);
nand UO_1887 (O_1887,N_14944,N_14442);
nand UO_1888 (O_1888,N_14892,N_14704);
and UO_1889 (O_1889,N_14703,N_14896);
nand UO_1890 (O_1890,N_14373,N_14847);
nand UO_1891 (O_1891,N_14009,N_14952);
nor UO_1892 (O_1892,N_14492,N_14318);
and UO_1893 (O_1893,N_14585,N_14659);
and UO_1894 (O_1894,N_14780,N_14220);
or UO_1895 (O_1895,N_14220,N_14517);
and UO_1896 (O_1896,N_14404,N_14937);
and UO_1897 (O_1897,N_14693,N_14554);
xnor UO_1898 (O_1898,N_14581,N_14954);
nor UO_1899 (O_1899,N_14732,N_14397);
and UO_1900 (O_1900,N_14973,N_14636);
or UO_1901 (O_1901,N_14723,N_14696);
nand UO_1902 (O_1902,N_14514,N_14145);
or UO_1903 (O_1903,N_14087,N_14161);
nor UO_1904 (O_1904,N_14704,N_14449);
nor UO_1905 (O_1905,N_14255,N_14475);
nand UO_1906 (O_1906,N_14013,N_14220);
or UO_1907 (O_1907,N_14421,N_14983);
or UO_1908 (O_1908,N_14521,N_14270);
or UO_1909 (O_1909,N_14804,N_14763);
nand UO_1910 (O_1910,N_14397,N_14710);
or UO_1911 (O_1911,N_14574,N_14787);
and UO_1912 (O_1912,N_14085,N_14122);
or UO_1913 (O_1913,N_14109,N_14119);
nor UO_1914 (O_1914,N_14821,N_14363);
or UO_1915 (O_1915,N_14610,N_14633);
or UO_1916 (O_1916,N_14395,N_14234);
xor UO_1917 (O_1917,N_14335,N_14479);
nor UO_1918 (O_1918,N_14311,N_14222);
xor UO_1919 (O_1919,N_14955,N_14602);
xnor UO_1920 (O_1920,N_14704,N_14100);
and UO_1921 (O_1921,N_14733,N_14561);
and UO_1922 (O_1922,N_14175,N_14100);
or UO_1923 (O_1923,N_14068,N_14144);
nor UO_1924 (O_1924,N_14807,N_14592);
nor UO_1925 (O_1925,N_14872,N_14376);
nor UO_1926 (O_1926,N_14125,N_14601);
nor UO_1927 (O_1927,N_14967,N_14796);
nor UO_1928 (O_1928,N_14853,N_14686);
and UO_1929 (O_1929,N_14811,N_14625);
nor UO_1930 (O_1930,N_14348,N_14789);
nand UO_1931 (O_1931,N_14682,N_14663);
nand UO_1932 (O_1932,N_14990,N_14438);
and UO_1933 (O_1933,N_14384,N_14522);
nand UO_1934 (O_1934,N_14203,N_14168);
nand UO_1935 (O_1935,N_14918,N_14920);
nand UO_1936 (O_1936,N_14022,N_14524);
and UO_1937 (O_1937,N_14258,N_14368);
or UO_1938 (O_1938,N_14743,N_14167);
nor UO_1939 (O_1939,N_14733,N_14094);
nand UO_1940 (O_1940,N_14487,N_14601);
or UO_1941 (O_1941,N_14642,N_14504);
or UO_1942 (O_1942,N_14722,N_14074);
nand UO_1943 (O_1943,N_14658,N_14023);
or UO_1944 (O_1944,N_14688,N_14429);
nand UO_1945 (O_1945,N_14334,N_14456);
nand UO_1946 (O_1946,N_14594,N_14319);
or UO_1947 (O_1947,N_14249,N_14404);
or UO_1948 (O_1948,N_14769,N_14304);
nor UO_1949 (O_1949,N_14952,N_14190);
nand UO_1950 (O_1950,N_14180,N_14822);
nand UO_1951 (O_1951,N_14865,N_14650);
or UO_1952 (O_1952,N_14940,N_14253);
nor UO_1953 (O_1953,N_14660,N_14560);
xnor UO_1954 (O_1954,N_14081,N_14588);
nor UO_1955 (O_1955,N_14543,N_14086);
nor UO_1956 (O_1956,N_14682,N_14107);
and UO_1957 (O_1957,N_14050,N_14962);
nor UO_1958 (O_1958,N_14013,N_14854);
nand UO_1959 (O_1959,N_14254,N_14663);
nor UO_1960 (O_1960,N_14848,N_14970);
or UO_1961 (O_1961,N_14801,N_14373);
nor UO_1962 (O_1962,N_14403,N_14136);
xnor UO_1963 (O_1963,N_14784,N_14661);
and UO_1964 (O_1964,N_14317,N_14485);
and UO_1965 (O_1965,N_14006,N_14924);
nor UO_1966 (O_1966,N_14497,N_14753);
nand UO_1967 (O_1967,N_14820,N_14045);
nor UO_1968 (O_1968,N_14827,N_14024);
or UO_1969 (O_1969,N_14782,N_14668);
nand UO_1970 (O_1970,N_14823,N_14559);
nor UO_1971 (O_1971,N_14420,N_14282);
and UO_1972 (O_1972,N_14697,N_14399);
nand UO_1973 (O_1973,N_14729,N_14838);
xnor UO_1974 (O_1974,N_14788,N_14380);
and UO_1975 (O_1975,N_14585,N_14065);
nand UO_1976 (O_1976,N_14385,N_14125);
or UO_1977 (O_1977,N_14355,N_14707);
nand UO_1978 (O_1978,N_14826,N_14416);
xor UO_1979 (O_1979,N_14626,N_14798);
or UO_1980 (O_1980,N_14298,N_14788);
nor UO_1981 (O_1981,N_14200,N_14130);
nor UO_1982 (O_1982,N_14303,N_14748);
and UO_1983 (O_1983,N_14646,N_14591);
xnor UO_1984 (O_1984,N_14506,N_14126);
nand UO_1985 (O_1985,N_14828,N_14574);
nor UO_1986 (O_1986,N_14972,N_14887);
nand UO_1987 (O_1987,N_14418,N_14959);
nand UO_1988 (O_1988,N_14617,N_14681);
nor UO_1989 (O_1989,N_14846,N_14262);
or UO_1990 (O_1990,N_14090,N_14638);
and UO_1991 (O_1991,N_14342,N_14902);
nor UO_1992 (O_1992,N_14649,N_14829);
xnor UO_1993 (O_1993,N_14051,N_14987);
and UO_1994 (O_1994,N_14618,N_14082);
or UO_1995 (O_1995,N_14883,N_14916);
nor UO_1996 (O_1996,N_14118,N_14116);
nor UO_1997 (O_1997,N_14162,N_14989);
or UO_1998 (O_1998,N_14511,N_14576);
or UO_1999 (O_1999,N_14627,N_14599);
endmodule